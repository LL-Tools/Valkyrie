

module b17_C_AntiSAT_k_256_10 ( P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, 
        DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, 
        DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, 
        DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, 
        DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, 
        DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, 
        HOLD, NA, BS16, READY1, READY2, P1_READREQUEST_REG_SCAN_IN, 
        P1_ADS_N_REG_SCAN_IN, P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, 
        P1_D_C_N_REG_SCAN_IN, P1_REQUESTPENDING_REG_SCAN_IN, 
        P1_STATEBS16_REG_SCAN_IN, P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, 
        P1_W_R_N_REG_SCAN_IN, P1_BYTEENABLE_REG_0__SCAN_IN, 
        P1_BYTEENABLE_REG_1__SCAN_IN, P1_BYTEENABLE_REG_2__SCAN_IN, 
        P1_BYTEENABLE_REG_3__SCAN_IN, P1_REIP_REG_31__SCAN_IN, 
        P1_REIP_REG_30__SCAN_IN, P1_REIP_REG_29__SCAN_IN, 
        P1_REIP_REG_28__SCAN_IN, P1_REIP_REG_27__SCAN_IN, 
        P1_REIP_REG_26__SCAN_IN, P1_REIP_REG_25__SCAN_IN, 
        P1_REIP_REG_24__SCAN_IN, P1_REIP_REG_23__SCAN_IN, 
        P1_REIP_REG_22__SCAN_IN, P1_REIP_REG_21__SCAN_IN, 
        P1_REIP_REG_20__SCAN_IN, P1_REIP_REG_19__SCAN_IN, 
        P1_REIP_REG_18__SCAN_IN, P1_REIP_REG_17__SCAN_IN, 
        P1_REIP_REG_16__SCAN_IN, P1_REIP_REG_15__SCAN_IN, 
        P1_REIP_REG_14__SCAN_IN, P1_REIP_REG_13__SCAN_IN, 
        P1_REIP_REG_12__SCAN_IN, P1_REIP_REG_11__SCAN_IN, 
        P1_REIP_REG_10__SCAN_IN, P1_REIP_REG_9__SCAN_IN, 
        P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN, 
        P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, P1_REIP_REG_3__SCAN_IN, 
        P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN, 
        P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, P1_EBX_REG_29__SCAN_IN, 
        P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN, 
        P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, P1_EBX_REG_23__SCAN_IN, 
        P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN, 
        P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, P1_EBX_REG_17__SCAN_IN, 
        P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN, 
        P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, P1_EBX_REG_11__SCAN_IN, 
        P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, P1_EBX_REG_8__SCAN_IN, 
        P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, P1_EBX_REG_5__SCAN_IN, 
        P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, P1_EBX_REG_2__SCAN_IN, 
        P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, P1_EAX_REG_31__SCAN_IN, 
        P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN, 
        P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, P1_EAX_REG_25__SCAN_IN, 
        P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN, 
        P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, P1_EAX_REG_19__SCAN_IN, 
        P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN, 
        P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, P1_EAX_REG_13__SCAN_IN, 
        P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, 
        P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, 
        P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, 
        P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, 
        P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, 
        keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, 
        keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, 
        keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, 
        keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, 
        keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, 
        keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, 
        keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, 
        keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, 
        keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, 
        keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, 
        keyinput60, keyinput61, keyinput62, keyinput63, keyinput64, keyinput65, 
        keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, keyinput71, 
        keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, keyinput77, 
        keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, keyinput83, 
        keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, keyinput89, 
        keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, keyinput95, 
        keyinput96, keyinput97, keyinput98, keyinput99, keyinput100, 
        keyinput101, keyinput102, keyinput103, keyinput104, keyinput105, 
        keyinput106, keyinput107, keyinput108, keyinput109, keyinput110, 
        keyinput111, keyinput112, keyinput113, keyinput114, keyinput115, 
        keyinput116, keyinput117, keyinput118, keyinput119, keyinput120, 
        keyinput121, keyinput122, keyinput123, keyinput124, keyinput125, 
        keyinput126, keyinput127, keyinput128, keyinput129, keyinput130, 
        keyinput131, keyinput132, keyinput133, keyinput134, keyinput135, 
        keyinput136, keyinput137, keyinput138, keyinput139, keyinput140, 
        keyinput141, keyinput142, keyinput143, keyinput144, keyinput145, 
        keyinput146, keyinput147, keyinput148, keyinput149, keyinput150, 
        keyinput151, keyinput152, keyinput153, keyinput154, keyinput155, 
        keyinput156, keyinput157, keyinput158, keyinput159, keyinput160, 
        keyinput161, keyinput162, keyinput163, keyinput164, keyinput165, 
        keyinput166, keyinput167, keyinput168, keyinput169, keyinput170, 
        keyinput171, keyinput172, keyinput173, keyinput174, keyinput175, 
        keyinput176, keyinput177, keyinput178, keyinput179, keyinput180, 
        keyinput181, keyinput182, keyinput183, keyinput184, keyinput185, 
        keyinput186, keyinput187, keyinput188, keyinput189, keyinput190, 
        keyinput191, keyinput192, keyinput193, keyinput194, keyinput195, 
        keyinput196, keyinput197, keyinput198, keyinput199, keyinput200, 
        keyinput201, keyinput202, keyinput203, keyinput204, keyinput205, 
        keyinput206, keyinput207, keyinput208, keyinput209, keyinput210, 
        keyinput211, keyinput212, keyinput213, keyinput214, keyinput215, 
        keyinput216, keyinput217, keyinput218, keyinput219, keyinput220, 
        keyinput221, keyinput222, keyinput223, keyinput224, keyinput225, 
        keyinput226, keyinput227, keyinput228, keyinput229, keyinput230, 
        keyinput231, keyinput232, keyinput233, keyinput234, keyinput235, 
        keyinput236, keyinput237, keyinput238, keyinput239, keyinput240, 
        keyinput241, keyinput242, keyinput243, keyinput244, keyinput245, 
        keyinput246, keyinput247, keyinput248, keyinput249, keyinput250, 
        keyinput251, keyinput252, keyinput253, keyinput254, keyinput255, U355, 
        U356, U357, U358, U359, U360, U361, U362, U363, U364, U366, U367, U368, 
        U369, U370, U371, U372, U373, U374, U375, U347, U348, U349, U350, U351, 
        U352, U353, U354, U365, U376, U247, U246, U245, U244, U243, U242, U241, 
        U240, U239, U238, U237, U236, U235, U234, U233, U232, U231, U230, U229, 
        U228, U227, U226, U225, U224, U223, U222, U221, U220, U219, U218, U217, 
        U216, U251, U252, U253, U254, U255, U256, U257, U258, U259, U260, U261, 
        U262, U263, U264, U265, U266, U267, U268, U269, U270, U271, U272, U273, 
        U274, U275, U276, U277, U278, U279, U280, U281, U282, U212, U215, U213, 
        U214, P3_U3274, P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, 
        P3_U3059, P3_U3058, P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, 
        P3_U3052, P3_U3051, P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, 
        P3_U3045, P3_U3044, P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, 
        P3_U3038, P3_U3037, P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, 
        P3_U3031, P3_U3030, P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, 
        P3_U3026, P3_U3025, P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, 
        P3_U3019, P3_U3018, P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, 
        P3_U3012, P3_U3011, P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, 
        P3_U3005, P3_U3004, P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, 
        P3_U3282, P3_U2998, P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, 
        P3_U2992, P3_U2991, P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, 
        P3_U2985, P3_U2984, P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, 
        P3_U2978, P3_U2977, P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, 
        P3_U2971, P3_U2970, P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, 
        P3_U2964, P3_U2963, P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, 
        P3_U2957, P3_U2956, P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, 
        P3_U2950, P3_U2949, P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, 
        P3_U2943, P3_U2942, P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, 
        P3_U2936, P3_U2935, P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, 
        P3_U2929, P3_U2928, P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, 
        P3_U2922, P3_U2921, P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, 
        P3_U2915, P3_U2914, P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, 
        P3_U2908, P3_U2907, P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, 
        P3_U2901, P3_U2900, P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, 
        P3_U2894, P3_U2893, P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, 
        P3_U2887, P3_U2886, P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, 
        P3_U2880, P3_U2879, P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, 
        P3_U2873, P3_U2872, P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, 
        P3_U3285, P3_U3288, P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, 
        P3_U2864, P3_U2863, P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, 
        P3_U2857, P3_U2856, P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, 
        P3_U2850, P3_U2849, P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, 
        P3_U2843, P3_U2842, P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, 
        P3_U2836, P3_U2835, P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, 
        P3_U2829, P3_U2828, P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, 
        P3_U2822, P3_U2821, P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, 
        P3_U2815, P3_U2814, P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, 
        P3_U2808, P3_U2807, P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, 
        P3_U2801, P3_U2800, P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, 
        P3_U2794, P3_U2793, P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, 
        P3_U2787, P3_U2786, P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, 
        P3_U2780, P3_U2779, P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, 
        P3_U2773, P3_U2772, P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, 
        P3_U2766, P3_U2765, P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, 
        P3_U2759, P3_U2758, P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, 
        P3_U2752, P3_U2751, P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, 
        P3_U2745, P3_U2744, P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, 
        P3_U2738, P3_U2737, P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, 
        P3_U2731, P3_U2730, P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, 
        P3_U2724, P3_U2723, P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, 
        P3_U2717, P3_U2716, P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, 
        P3_U2710, P3_U2709, P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, 
        P3_U2703, P3_U2702, P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, 
        P3_U2696, P3_U2695, P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, 
        P3_U2689, P3_U2688, P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, 
        P3_U2682, P3_U2681, P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, 
        P3_U2675, P3_U2674, P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, 
        P3_U2668, P3_U2667, P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, 
        P3_U2661, P3_U2660, P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, 
        P3_U2654, P3_U2653, P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, 
        P3_U2647, P3_U2646, P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, 
        P3_U2640, P3_U2639, P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, 
        P3_U3295, P3_U2636, P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, 
        P3_U3298, P3_U3299, P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, 
        P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, 
        P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, 
        P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, 
        P2_U3179, P2_U3593, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, 
        P2_U3173, P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, 
        P2_U3166, P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, 
        P2_U3159, P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, 
        P2_U3152, P2_U3151, P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, 
        P2_U3145, P2_U3144, P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, 
        P2_U3138, P2_U3137, P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, 
        P2_U3131, P2_U3130, P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, 
        P2_U3124, P2_U3123, P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, 
        P2_U3117, P2_U3116, P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, 
        P2_U3110, P2_U3109, P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, 
        P2_U3103, P2_U3102, P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, 
        P2_U3096, P2_U3095, P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, 
        P2_U3089, P2_U3088, P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, 
        P2_U3082, P2_U3081, P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, 
        P2_U3075, P2_U3074, P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, 
        P2_U3068, P2_U3067, P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, 
        P2_U3061, P2_U3060, P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, 
        P2_U3054, P2_U3053, P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, 
        P2_U3595, P2_U3596, P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, 
        P2_U3603, P2_U3604, P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, 
        P2_U3042, P2_U3041, P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, 
        P2_U3035, P2_U3034, P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, 
        P2_U3028, P2_U3027, P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, 
        P2_U3021, P2_U3020, P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, 
        P2_U3014, P2_U3013, P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, 
        P2_U3007, P2_U3006, P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, 
        P2_U3000, P2_U2999, P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, 
        P2_U2993, P2_U2992, P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, 
        P2_U2986, P2_U2985, P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, 
        P2_U2979, P2_U2978, P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, 
        P2_U2972, P2_U2971, P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, 
        P2_U2965, P2_U2964, P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, 
        P2_U2958, P2_U2957, P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, 
        P2_U2951, P2_U2950, P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, 
        P2_U2944, P2_U2943, P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, 
        P2_U2937, P2_U2936, P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, 
        P2_U2930, P2_U2929, P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, 
        P2_U2923, P2_U2922, P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, 
        P2_U2916, P2_U2915, P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, 
        P2_U2909, P2_U2908, P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, 
        P2_U2902, P2_U2901, P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, 
        P2_U2895, P2_U2894, P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, 
        P2_U2888, P2_U2887, P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, 
        P2_U2881, P2_U2880, P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, 
        P2_U2874, P2_U2873, P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, 
        P2_U2867, P2_U2866, P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, 
        P2_U2860, P2_U2859, P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, 
        P2_U2853, P2_U2852, P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, 
        P2_U2846, P2_U2845, P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, 
        P2_U2839, P2_U2838, P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, 
        P2_U2832, P2_U2831, P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, 
        P2_U2825, P2_U2824, P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, 
        P2_U2819, P2_U3609, P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, 
        P2_U2815, P2_U3612, P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, 
        P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, 
        P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, 
        P1_U3212, P1_U3211, P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, 
        P1_U3205, P1_U3204, P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, 
        P1_U3198, P1_U3197, P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, 
        P1_U3193, P1_U3192, P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, 
        P1_U3186, P1_U3185, P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, 
        P1_U3179, P1_U3178, P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, 
        P1_U3172, P1_U3171, P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, 
        P1_U3165, P1_U3164, P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, 
        P1_U3159, P1_U3158, P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, 
        P1_U3152, P1_U3151, P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, 
        P1_U3145, P1_U3144, P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, 
        P1_U3138, P1_U3137, P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, 
        P1_U3131, P1_U3130, P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, 
        P1_U3124, P1_U3123, P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, 
        P1_U3117, P1_U3116, P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, 
        P1_U3110, P1_U3109, P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, 
        P1_U3103, P1_U3102, P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, 
        P1_U3096, P1_U3095, P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, 
        P1_U3089, P1_U3088, P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, 
        P1_U3082, P1_U3081, P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, 
        P1_U3075, P1_U3074, P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, 
        P1_U3068, P1_U3067, P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, 
        P1_U3061, P1_U3060, P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, 
        P1_U3054, P1_U3053, P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, 
        P1_U3047, P1_U3046, P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, 
        P1_U3040, P1_U3039, P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, 
        P1_U3033, P1_U3468, P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, 
        P1_U3475, P1_U3476, P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, 
        P1_U3028, P1_U3027, P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, 
        P1_U3021, P1_U3020, P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, 
        P1_U3014, P1_U3013, P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, 
        P1_U3007, P1_U3006, P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, 
        P1_U3000, P1_U2999, P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, 
        P1_U2993, P1_U2992, P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, 
        P1_U2986, P1_U2985, P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, 
        P1_U2979, P1_U2978, P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, 
        P1_U2972, P1_U2971, P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, 
        P1_U2965, P1_U2964, P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, 
        P1_U2958, P1_U2957, P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, 
        P1_U2951, P1_U2950, P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, 
        P1_U2944, P1_U2943, P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, 
        P1_U2937, P1_U2936, P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, 
        P1_U2930, P1_U2929, P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, 
        P1_U2923, P1_U2922, P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, 
        P1_U2916, P1_U2915, P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, 
        P1_U2909, P1_U2908, P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, 
        P1_U2902, P1_U2901, P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, 
        P1_U2895, P1_U2894, P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, 
        P1_U2888, P1_U2887, P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, 
        P1_U2881, P1_U2880, P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, 
        P1_U2874, P1_U2873, P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, 
        P1_U2867, P1_U2866, P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, 
        P1_U2860, P1_U2859, P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, 
        P1_U2853, P1_U2852, P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, 
        P1_U2846, P1_U2845, P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, 
        P1_U2839, P1_U2838, P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, 
        P1_U2832, P1_U2831, P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, 
        P1_U2825, P1_U2824, P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, 
        P1_U2818, P1_U2817, P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, 
        P1_U2811, P1_U2810, P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, 
        P1_U3483, P1_U2806, P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, 
        P1_U2803, P1_U2802, P1_U3487, P1_U2801 );
  input P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_,
         DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_,
         DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_,
         DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_,
         DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_,
         DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2,
         P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
         P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
         P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
         P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
         P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
         P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
         P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
         P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
         P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
         P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
         P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
         P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
         P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
         P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
         P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
         P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
         P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
         P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN,
         P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
         P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
         P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN,
         P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN,
         P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
         P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
         P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN,
         P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
         P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
         P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN,
         P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
         P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
         P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN,
         P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
         P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
         P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
         P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
         P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
         P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
         P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN,
         P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
         P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
         P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN,
         P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
         P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
         P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN,
         P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
         P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
         P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
         P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
         P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
         P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN, keyinput0, keyinput1, keyinput2,
         keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8,
         keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127, keyinput128, keyinput129,
         keyinput130, keyinput131, keyinput132, keyinput133, keyinput134,
         keyinput135, keyinput136, keyinput137, keyinput138, keyinput139,
         keyinput140, keyinput141, keyinput142, keyinput143, keyinput144,
         keyinput145, keyinput146, keyinput147, keyinput148, keyinput149,
         keyinput150, keyinput151, keyinput152, keyinput153, keyinput154,
         keyinput155, keyinput156, keyinput157, keyinput158, keyinput159,
         keyinput160, keyinput161, keyinput162, keyinput163, keyinput164,
         keyinput165, keyinput166, keyinput167, keyinput168, keyinput169,
         keyinput170, keyinput171, keyinput172, keyinput173, keyinput174,
         keyinput175, keyinput176, keyinput177, keyinput178, keyinput179,
         keyinput180, keyinput181, keyinput182, keyinput183, keyinput184,
         keyinput185, keyinput186, keyinput187, keyinput188, keyinput189,
         keyinput190, keyinput191, keyinput192, keyinput193, keyinput194,
         keyinput195, keyinput196, keyinput197, keyinput198, keyinput199,
         keyinput200, keyinput201, keyinput202, keyinput203, keyinput204,
         keyinput205, keyinput206, keyinput207, keyinput208, keyinput209,
         keyinput210, keyinput211, keyinput212, keyinput213, keyinput214,
         keyinput215, keyinput216, keyinput217, keyinput218, keyinput219,
         keyinput220, keyinput221, keyinput222, keyinput223, keyinput224,
         keyinput225, keyinput226, keyinput227, keyinput228, keyinput229,
         keyinput230, keyinput231, keyinput232, keyinput233, keyinput234,
         keyinput235, keyinput236, keyinput237, keyinput238, keyinput239,
         keyinput240, keyinput241, keyinput242, keyinput243, keyinput244,
         keyinput245, keyinput246, keyinput247, keyinput248, keyinput249,
         keyinput250, keyinput251, keyinput252, keyinput253, keyinput254,
         keyinput255;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825,
         n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835,
         n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845,
         n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855,
         n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865,
         n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875,
         n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885,
         n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895,
         n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905,
         n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915,
         n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925,
         n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935,
         n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945,
         n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955,
         n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965,
         n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975,
         n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985,
         n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995,
         n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004,
         n10005, n10006, n10007, n10008, n10009, n10010, n10011, n10012,
         n10013, n10014, n10015, n10016, n10017, n10018, n10019, n10020,
         n10021, n10022, n10023, n10024, n10025, n10026, n10027, n10028,
         n10029, n10030, n10031, n10032, n10033, n10034, n10035, n10036,
         n10037, n10038, n10039, n10040, n10041, n10042, n10043, n10044,
         n10045, n10046, n10047, n10048, n10049, n10050, n10051, n10052,
         n10053, n10054, n10055, n10056, n10057, n10058, n10059, n10060,
         n10061, n10062, n10063, n10064, n10065, n10066, n10067, n10068,
         n10069, n10070, n10071, n10072, n10073, n10074, n10075, n10076,
         n10077, n10078, n10079, n10080, n10081, n10082, n10083, n10084,
         n10085, n10086, n10087, n10088, n10089, n10090, n10091, n10092,
         n10093, n10094, n10095, n10096, n10097, n10098, n10099, n10100,
         n10101, n10102, n10103, n10104, n10105, n10106, n10107, n10108,
         n10109, n10110, n10111, n10112, n10113, n10114, n10115, n10116,
         n10117, n10118, n10119, n10120, n10121, n10122, n10123, n10124,
         n10125, n10126, n10127, n10128, n10129, n10130, n10131, n10132,
         n10133, n10134, n10135, n10136, n10137, n10138, n10139, n10140,
         n10141, n10142, n10143, n10144, n10145, n10146, n10147, n10148,
         n10149, n10150, n10151, n10152, n10153, n10154, n10155, n10156,
         n10157, n10158, n10159, n10160, n10161, n10162, n10163, n10164,
         n10165, n10166, n10167, n10168, n10169, n10170, n10171, n10172,
         n10173, n10174, n10175, n10176, n10177, n10178, n10179, n10180,
         n10181, n10182, n10183, n10184, n10185, n10186, n10187, n10188,
         n10189, n10190, n10191, n10192, n10193, n10194, n10195, n10196,
         n10197, n10198, n10199, n10200, n10201, n10202, n10203, n10204,
         n10205, n10206, n10207, n10208, n10209, n10210, n10211, n10212,
         n10213, n10214, n10215, n10216, n10217, n10218, n10219, n10220,
         n10221, n10222, n10223, n10224, n10225, n10226, n10227, n10228,
         n10229, n10230, n10231, n10232, n10233, n10234, n10235, n10236,
         n10237, n10238, n10239, n10240, n10241, n10242, n10243, n10244,
         n10245, n10246, n10247, n10248, n10249, n10250, n10251, n10252,
         n10253, n10254, n10255, n10256, n10257, n10258, n10259, n10260,
         n10261, n10262, n10263, n10264, n10265, n10266, n10267, n10268,
         n10269, n10270, n10271, n10272, n10273, n10274, n10275, n10276,
         n10277, n10278, n10279, n10280, n10281, n10282, n10283, n10284,
         n10285, n10286, n10287, n10288, n10289, n10290, n10291, n10292,
         n10293, n10294, n10295, n10296, n10297, n10298, n10299, n10300,
         n10301, n10302, n10303, n10304, n10305, n10306, n10307, n10308,
         n10309, n10310, n10311, n10312, n10313, n10314, n10315, n10316,
         n10317, n10318, n10319, n10320, n10321, n10322, n10323, n10324,
         n10325, n10326, n10327, n10328, n10329, n10330, n10331, n10332,
         n10333, n10334, n10335, n10336, n10337, n10338, n10339, n10340,
         n10341, n10342, n10343, n10344, n10345, n10346, n10347, n10348,
         n10349, n10350, n10351, n10352, n10353, n10354, n10355, n10356,
         n10357, n10358, n10359, n10360, n10361, n10362, n10363, n10364,
         n10365, n10366, n10367, n10368, n10369, n10370, n10371, n10372,
         n10373, n10374, n10375, n10376, n10377, n10378, n10379, n10380,
         n10381, n10382, n10383, n10384, n10385, n10386, n10387, n10388,
         n10389, n10390, n10391, n10392, n10393, n10394, n10395, n10396,
         n10397, n10398, n10399, n10400, n10401, n10402, n10403, n10404,
         n10405, n10406, n10407, n10408, n10409, n10410, n10411, n10412,
         n10413, n10414, n10415, n10416, n10417, n10418, n10419, n10420,
         n10421, n10422, n10423, n10424, n10425, n10426, n10427, n10428,
         n10429, n10430, n10431, n10432, n10433, n10434, n10435, n10436,
         n10437, n10438, n10439, n10440, n10441, n10442, n10443, n10444,
         n10445, n10446, n10447, n10448, n10449, n10450, n10451, n10452,
         n10453, n10454, n10455, n10456, n10457, n10458, n10459, n10460,
         n10461, n10462, n10463, n10464, n10465, n10466, n10467, n10468,
         n10469, n10470, n10471, n10472, n10473, n10474, n10475, n10476,
         n10477, n10478, n10479, n10480, n10481, n10482, n10483, n10484,
         n10485, n10486, n10487, n10488, n10489, n10490, n10491, n10492,
         n10493, n10494, n10495, n10496, n10497, n10498, n10499, n10500,
         n10501, n10502, n10503, n10504, n10505, n10506, n10507, n10508,
         n10509, n10510, n10511, n10512, n10513, n10514, n10515, n10516,
         n10517, n10518, n10519, n10520, n10521, n10522, n10523, n10524,
         n10525, n10526, n10527, n10528, n10529, n10530, n10531, n10532,
         n10533, n10534, n10535, n10536, n10537, n10538, n10539, n10540,
         n10541, n10542, n10543, n10544, n10545, n10546, n10547, n10548,
         n10549, n10550, n10551, n10552, n10553, n10554, n10555, n10556,
         n10557, n10558, n10559, n10560, n10561, n10562, n10563, n10564,
         n10565, n10566, n10567, n10568, n10569, n10570, n10571, n10572,
         n10573, n10574, n10575, n10576, n10577, n10578, n10579, n10580,
         n10581, n10582, n10583, n10584, n10585, n10586, n10587, n10588,
         n10589, n10590, n10591, n10592, n10593, n10594, n10595, n10596,
         n10597, n10598, n10599, n10600, n10601, n10602, n10603, n10604,
         n10605, n10606, n10607, n10608, n10609, n10610, n10611, n10612,
         n10613, n10614, n10615, n10616, n10617, n10618, n10619, n10620,
         n10621, n10622, n10623, n10624, n10625, n10626, n10627, n10628,
         n10629, n10630, n10631, n10632, n10633, n10634, n10635, n10636,
         n10637, n10638, n10639, n10640, n10641, n10642, n10643, n10644,
         n10645, n10646, n10647, n10648, n10649, n10650, n10651, n10652,
         n10653, n10654, n10655, n10656, n10657, n10658, n10659, n10660,
         n10661, n10662, n10663, n10664, n10665, n10666, n10667, n10668,
         n10669, n10670, n10671, n10672, n10673, n10674, n10675, n10676,
         n10677, n10678, n10679, n10680, n10681, n10682, n10683, n10684,
         n10685, n10686, n10687, n10688, n10689, n10690, n10691, n10692,
         n10693, n10694, n10695, n10696, n10697, n10698, n10699, n10700,
         n10701, n10702, n10703, n10704, n10705, n10706, n10707, n10708,
         n10709, n10710, n10711, n10712, n10713, n10714, n10715, n10716,
         n10717, n10718, n10719, n10720, n10721, n10722, n10723, n10724,
         n10725, n10726, n10727, n10728, n10729, n10730, n10731, n10732,
         n10733, n10734, n10735, n10736, n10737, n10738, n10739, n10740,
         n10741, n10742, n10743, n10744, n10745, n10746, n10747, n10748,
         n10749, n10750, n10751, n10752, n10753, n10754, n10755, n10756,
         n10757, n10758, n10759, n10760, n10761, n10762, n10763, n10764,
         n10765, n10766, n10767, n10768, n10769, n10770, n10771, n10772,
         n10773, n10774, n10775, n10776, n10777, n10778, n10779, n10780,
         n10781, n10782, n10783, n10784, n10785, n10786, n10787, n10788,
         n10789, n10790, n10791, n10792, n10793, n10794, n10795, n10796,
         n10797, n10798, n10799, n10800, n10801, n10802, n10803, n10804,
         n10805, n10806, n10807, n10808, n10809, n10810, n10811, n10812,
         n10813, n10814, n10815, n10816, n10817, n10818, n10819, n10820,
         n10821, n10822, n10823, n10824, n10825, n10826, n10827, n10828,
         n10829, n10830, n10831, n10832, n10833, n10834, n10835, n10836,
         n10837, n10838, n10839, n10840, n10841, n10842, n10843, n10844,
         n10845, n10846, n10847, n10848, n10849, n10850, n10851, n10852,
         n10853, n10854, n10855, n10856, n10857, n10858, n10859, n10860,
         n10861, n10862, n10863, n10864, n10865, n10866, n10867, n10868,
         n10869, n10870, n10871, n10872, n10873, n10874, n10875, n10876,
         n10877, n10878, n10879, n10880, n10881, n10882, n10883, n10884,
         n10885, n10886, n10887, n10888, n10889, n10890, n10891, n10892,
         n10893, n10894, n10895, n10896, n10897, n10898, n10899, n10900,
         n10901, n10902, n10903, n10904, n10905, n10906, n10907, n10908,
         n10909, n10910, n10911, n10912, n10913, n10914, n10915, n10916,
         n10917, n10918, n10919, n10920, n10921, n10922, n10923, n10924,
         n10925, n10926, n10927, n10928, n10929, n10930, n10931, n10932,
         n10933, n10934, n10935, n10936, n10937, n10938, n10939, n10940,
         n10941, n10942, n10943, n10944, n10945, n10946, n10947, n10948,
         n10949, n10950, n10951, n10952, n10953, n10954, n10955, n10956,
         n10957, n10958, n10959, n10960, n10961, n10962, n10963, n10964,
         n10965, n10966, n10967, n10968, n10969, n10970, n10971, n10972,
         n10973, n10974, n10975, n10976, n10977, n10978, n10979, n10980,
         n10981, n10982, n10983, n10984, n10985, n10986, n10987, n10988,
         n10989, n10990, n10991, n10992, n10993, n10994, n10995, n10996,
         n10997, n10998, n10999, n11000, n11001, n11002, n11003, n11004,
         n11005, n11006, n11007, n11008, n11009, n11010, n11011, n11012,
         n11013, n11014, n11015, n11016, n11017, n11018, n11019, n11020,
         n11021, n11022, n11023, n11024, n11025, n11026, n11027, n11028,
         n11029, n11030, n11031, n11032, n11033, n11034, n11035, n11036,
         n11037, n11038, n11039, n11040, n11041, n11042, n11043, n11044,
         n11045, n11046, n11047, n11048, n11049, n11050, n11051, n11052,
         n11053, n11054, n11055, n11056, n11057, n11058, n11059, n11060,
         n11061, n11062, n11063, n11064, n11065, n11066, n11067, n11068,
         n11069, n11070, n11071, n11072, n11073, n11074, n11075, n11076,
         n11077, n11078, n11079, n11080, n11081, n11082, n11083, n11084,
         n11085, n11086, n11087, n11088, n11089, n11090, n11091, n11092,
         n11093, n11094, n11095, n11096, n11097, n11098, n11099, n11100,
         n11101, n11102, n11103, n11104, n11105, n11106, n11107, n11108,
         n11109, n11110, n11111, n11112, n11113, n11114, n11115, n11116,
         n11117, n11118, n11119, n11120, n11121, n11122, n11123, n11124,
         n11125, n11126, n11127, n11128, n11129, n11130, n11131, n11132,
         n11133, n11134, n11135, n11136, n11137, n11138, n11139, n11140,
         n11141, n11142, n11143, n11144, n11145, n11146, n11147, n11148,
         n11149, n11150, n11151, n11152, n11153, n11154, n11155, n11156,
         n11157, n11158, n11159, n11160, n11161, n11162, n11163, n11164,
         n11165, n11166, n11167, n11168, n11169, n11170, n11171, n11172,
         n11173, n11174, n11175, n11176, n11177, n11178, n11179, n11180,
         n11181, n11182, n11183, n11184, n11185, n11186, n11187, n11188,
         n11189, n11190, n11191, n11192, n11193, n11194, n11195, n11196,
         n11197, n11198, n11199, n11200, n11201, n11202, n11203, n11204,
         n11205, n11206, n11207, n11208, n11209, n11210, n11211, n11212,
         n11213, n11214, n11215, n11216, n11217, n11218, n11219, n11220,
         n11221, n11222, n11223, n11224, n11225, n11226, n11227, n11228,
         n11229, n11230, n11231, n11232, n11233, n11234, n11235, n11236,
         n11237, n11238, n11239, n11240, n11241, n11242, n11243, n11244,
         n11245, n11246, n11247, n11248, n11249, n11250, n11251, n11252,
         n11253, n11254, n11255, n11256, n11257, n11258, n11259, n11260,
         n11261, n11262, n11263, n11264, n11265, n11266, n11267, n11268,
         n11269, n11270, n11271, n11272, n11273, n11274, n11275, n11276,
         n11277, n11278, n11279, n11280, n11281, n11282, n11283, n11284,
         n11285, n11286, n11287, n11288, n11289, n11290, n11291, n11292,
         n11293, n11294, n11295, n11296, n11297, n11298, n11299, n11300,
         n11301, n11302, n11303, n11304, n11305, n11306, n11307, n11308,
         n11309, n11310, n11311, n11312, n11313, n11314, n11315, n11316,
         n11317, n11318, n11319, n11320, n11321, n11322, n11323, n11324,
         n11325, n11326, n11327, n11328, n11329, n11330, n11331, n11332,
         n11333, n11334, n11335, n11336, n11337, n11338, n11339, n11340,
         n11341, n11342, n11343, n11344, n11345, n11346, n11347, n11348,
         n11349, n11350, n11351, n11352, n11353, n11354, n11355, n11356,
         n11357, n11358, n11359, n11360, n11361, n11362, n11363, n11364,
         n11365, n11366, n11367, n11368, n11369, n11370, n11371, n11372,
         n11373, n11374, n11375, n11376, n11377, n11378, n11379, n11380,
         n11381, n11382, n11383, n11384, n11385, n11386, n11387, n11388,
         n11389, n11390, n11391, n11392, n11393, n11394, n11395, n11396,
         n11397, n11398, n11399, n11400, n11401, n11402, n11403, n11404,
         n11405, n11406, n11407, n11408, n11409, n11410, n11411, n11412,
         n11413, n11414, n11415, n11416, n11417, n11418, n11419, n11420,
         n11421, n11422, n11423, n11424, n11425, n11426, n11427, n11428,
         n11429, n11430, n11431, n11432, n11433, n11434, n11435, n11436,
         n11437, n11438, n11439, n11440, n11441, n11442, n11443, n11444,
         n11445, n11446, n11447, n11448, n11449, n11450, n11451, n11452,
         n11453, n11454, n11455, n11456, n11457, n11458, n11459, n11460,
         n11461, n11462, n11463, n11464, n11465, n11466, n11467, n11468,
         n11469, n11470, n11471, n11472, n11473, n11474, n11475, n11476,
         n11477, n11478, n11479, n11480, n11481, n11482, n11483, n11484,
         n11485, n11486, n11487, n11488, n11489, n11490, n11491, n11492,
         n11493, n11494, n11495, n11496, n11497, n11498, n11499, n11500,
         n11501, n11502, n11503, n11504, n11505, n11506, n11507, n11508,
         n11509, n11510, n11511, n11512, n11513, n11514, n11515, n11516,
         n11517, n11518, n11519, n11520, n11521, n11522, n11523, n11524,
         n11525, n11526, n11527, n11528, n11529, n11530, n11531, n11532,
         n11533, n11534, n11535, n11536, n11537, n11538, n11539, n11540,
         n11541, n11542, n11543, n11544, n11545, n11546, n11547, n11548,
         n11549, n11550, n11551, n11552, n11553, n11554, n11555, n11556,
         n11557, n11558, n11559, n11560, n11561, n11562, n11563, n11564,
         n11565, n11566, n11567, n11568, n11569, n11570, n11571, n11572,
         n11573, n11574, n11575, n11576, n11577, n11578, n11579, n11580,
         n11581, n11582, n11583, n11584, n11585, n11586, n11587, n11588,
         n11589, n11590, n11591, n11592, n11593, n11594, n11595, n11596,
         n11597, n11598, n11599, n11600, n11601, n11602, n11603, n11604,
         n11605, n11606, n11607, n11608, n11609, n11610, n11611, n11612,
         n11613, n11614, n11615, n11616, n11617, n11618, n11619, n11620,
         n11621, n11622, n11623, n11624, n11625, n11626, n11627, n11628,
         n11629, n11630, n11631, n11632, n11633, n11634, n11635, n11636,
         n11637, n11638, n11639, n11640, n11641, n11642, n11643, n11644,
         n11645, n11646, n11647, n11648, n11649, n11650, n11651, n11652,
         n11653, n11654, n11655, n11656, n11657, n11658, n11659, n11660,
         n11661, n11662, n11663, n11664, n11665, n11666, n11667, n11668,
         n11669, n11670, n11671, n11672, n11673, n11674, n11675, n11676,
         n11677, n11678, n11679, n11680, n11681, n11682, n11683, n11684,
         n11685, n11686, n11687, n11688, n11689, n11690, n11691, n11692,
         n11693, n11694, n11695, n11696, n11697, n11698, n11699, n11700,
         n11701, n11702, n11703, n11704, n11705, n11706, n11707, n11708,
         n11709, n11710, n11711, n11712, n11713, n11714, n11715, n11716,
         n11717, n11718, n11719, n11720, n11721, n11722, n11723, n11724,
         n11725, n11726, n11727, n11728, n11729, n11730, n11731, n11732,
         n11733, n11734, n11735, n11736, n11737, n11738, n11739, n11740,
         n11741, n11742, n11743, n11744, n11745, n11746, n11747, n11748,
         n11749, n11750, n11751, n11752, n11753, n11754, n11755, n11756,
         n11757, n11758, n11759, n11760, n11761, n11762, n11763, n11764,
         n11765, n11766, n11767, n11768, n11769, n11770, n11771, n11772,
         n11773, n11774, n11775, n11776, n11777, n11778, n11779, n11780,
         n11781, n11782, n11783, n11784, n11785, n11786, n11787, n11788,
         n11789, n11790, n11791, n11792, n11793, n11794, n11795, n11796,
         n11797, n11798, n11799, n11800, n11801, n11802, n11803, n11804,
         n11805, n11806, n11807, n11808, n11809, n11810, n11811, n11812,
         n11813, n11814, n11815, n11816, n11817, n11818, n11819, n11820,
         n11821, n11822, n11823, n11824, n11825, n11826, n11827, n11828,
         n11829, n11830, n11831, n11832, n11833, n11834, n11835, n11836,
         n11837, n11838, n11839, n11840, n11841, n11842, n11843, n11844,
         n11845, n11846, n11847, n11848, n11849, n11850, n11851, n11852,
         n11853, n11854, n11855, n11856, n11857, n11858, n11859, n11860,
         n11861, n11862, n11863, n11864, n11865, n11866, n11867, n11868,
         n11869, n11870, n11871, n11872, n11873, n11874, n11875, n11876,
         n11877, n11878, n11879, n11880, n11881, n11882, n11883, n11884,
         n11885, n11886, n11887, n11888, n11889, n11890, n11891, n11892,
         n11893, n11894, n11895, n11896, n11897, n11898, n11899, n11900,
         n11901, n11902, n11903, n11904, n11905, n11906, n11907, n11908,
         n11909, n11910, n11911, n11912, n11913, n11914, n11915, n11916,
         n11917, n11918, n11919, n11920, n11921, n11922, n11923, n11924,
         n11925, n11926, n11927, n11928, n11929, n11930, n11931, n11932,
         n11933, n11934, n11935, n11936, n11937, n11938, n11939, n11940,
         n11941, n11942, n11943, n11944, n11945, n11946, n11947, n11948,
         n11949, n11950, n11951, n11952, n11953, n11954, n11955, n11956,
         n11957, n11958, n11959, n11960, n11961, n11962, n11963, n11964,
         n11965, n11966, n11967, n11968, n11969, n11970, n11971, n11972,
         n11973, n11974, n11975, n11976, n11977, n11978, n11979, n11980,
         n11981, n11982, n11983, n11984, n11985, n11986, n11987, n11988,
         n11989, n11990, n11991, n11992, n11993, n11994, n11995, n11996,
         n11997, n11998, n11999, n12000, n12001, n12002, n12003, n12004,
         n12005, n12006, n12007, n12008, n12009, n12010, n12011, n12012,
         n12013, n12014, n12015, n12016, n12017, n12018, n12019, n12020,
         n12021, n12022, n12023, n12024, n12025, n12026, n12027, n12028,
         n12029, n12030, n12031, n12032, n12033, n12034, n12035, n12036,
         n12037, n12038, n12039, n12040, n12041, n12042, n12043, n12044,
         n12045, n12046, n12047, n12048, n12049, n12050, n12051, n12052,
         n12053, n12054, n12055, n12056, n12057, n12058, n12059, n12060,
         n12061, n12062, n12063, n12064, n12065, n12066, n12067, n12068,
         n12069, n12070, n12071, n12072, n12073, n12074, n12075, n12076,
         n12077, n12078, n12079, n12080, n12081, n12082, n12083, n12084,
         n12085, n12086, n12087, n12088, n12089, n12090, n12091, n12092,
         n12093, n12094, n12095, n12096, n12097, n12098, n12099, n12100,
         n12101, n12102, n12103, n12104, n12105, n12106, n12107, n12108,
         n12109, n12110, n12111, n12112, n12113, n12114, n12115, n12116,
         n12117, n12118, n12119, n12120, n12121, n12122, n12123, n12124,
         n12125, n12126, n12127, n12128, n12129, n12130, n12131, n12132,
         n12133, n12134, n12135, n12136, n12137, n12138, n12139, n12140,
         n12141, n12142, n12143, n12144, n12145, n12146, n12147, n12148,
         n12149, n12150, n12151, n12152, n12153, n12154, n12155, n12156,
         n12157, n12158, n12159, n12160, n12161, n12162, n12163, n12164,
         n12165, n12166, n12167, n12168, n12169, n12170, n12171, n12172,
         n12173, n12174, n12175, n12176, n12177, n12178, n12179, n12180,
         n12181, n12182, n12183, n12184, n12185, n12186, n12187, n12188,
         n12189, n12190, n12191, n12192, n12193, n12194, n12195, n12196,
         n12197, n12198, n12199, n12200, n12201, n12202, n12203, n12204,
         n12205, n12206, n12207, n12208, n12209, n12210, n12211, n12212,
         n12213, n12214, n12215, n12216, n12217, n12218, n12219, n12220,
         n12221, n12222, n12223, n12224, n12225, n12226, n12227, n12228,
         n12229, n12230, n12231, n12232, n12233, n12234, n12235, n12236,
         n12237, n12238, n12239, n12240, n12241, n12242, n12243, n12244,
         n12245, n12246, n12247, n12248, n12249, n12250, n12251, n12252,
         n12253, n12254, n12255, n12256, n12257, n12258, n12259, n12260,
         n12261, n12262, n12263, n12264, n12265, n12266, n12267, n12268,
         n12269, n12270, n12271, n12272, n12273, n12274, n12275, n12276,
         n12277, n12278, n12279, n12280, n12281, n12282, n12283, n12284,
         n12285, n12286, n12287, n12288, n12289, n12290, n12291, n12292,
         n12293, n12294, n12295, n12296, n12297, n12298, n12299, n12300,
         n12301, n12302, n12303, n12304, n12305, n12306, n12307, n12308,
         n12309, n12310, n12311, n12312, n12313, n12314, n12315, n12316,
         n12317, n12318, n12319, n12320, n12321, n12322, n12323, n12324,
         n12325, n12326, n12327, n12328, n12329, n12330, n12331, n12332,
         n12333, n12334, n12335, n12336, n12337, n12338, n12339, n12340,
         n12341, n12342, n12343, n12344, n12345, n12346, n12347, n12348,
         n12349, n12350, n12351, n12352, n12353, n12354, n12355, n12356,
         n12357, n12358, n12359, n12360, n12361, n12362, n12363, n12364,
         n12365, n12366, n12367, n12368, n12369, n12370, n12371, n12372,
         n12373, n12374, n12375, n12376, n12377, n12378, n12379, n12380,
         n12381, n12382, n12383, n12384, n12385, n12386, n12387, n12388,
         n12389, n12390, n12391, n12392, n12393, n12394, n12395, n12396,
         n12397, n12398, n12399, n12400, n12401, n12402, n12403, n12404,
         n12405, n12406, n12407, n12408, n12409, n12410, n12411, n12412,
         n12413, n12414, n12415, n12416, n12417, n12418, n12419, n12420,
         n12421, n12422, n12423, n12424, n12425, n12426, n12427, n12428,
         n12429, n12430, n12431, n12432, n12433, n12434, n12435, n12436,
         n12437, n12438, n12439, n12440, n12441, n12442, n12443, n12444,
         n12445, n12446, n12447, n12448, n12449, n12450, n12451, n12452,
         n12453, n12454, n12455, n12456, n12457, n12458, n12459, n12460,
         n12461, n12462, n12463, n12464, n12465, n12466, n12467, n12468,
         n12469, n12470, n12471, n12472, n12473, n12474, n12475, n12476,
         n12477, n12478, n12479, n12480, n12481, n12482, n12483, n12484,
         n12485, n12486, n12487, n12488, n12489, n12490, n12491, n12492,
         n12493, n12494, n12495, n12496, n12497, n12498, n12499, n12500,
         n12501, n12502, n12503, n12504, n12505, n12506, n12507, n12508,
         n12509, n12510, n12511, n12512, n12513, n12514, n12515, n12516,
         n12517, n12518, n12519, n12520, n12521, n12522, n12523, n12524,
         n12525, n12526, n12527, n12528, n12529, n12530, n12531, n12532,
         n12533, n12534, n12535, n12536, n12537, n12538, n12539, n12540,
         n12541, n12542, n12543, n12544, n12545, n12546, n12547, n12548,
         n12549, n12550, n12551, n12552, n12553, n12554, n12555, n12556,
         n12557, n12558, n12559, n12560, n12561, n12562, n12563, n12564,
         n12565, n12566, n12567, n12568, n12569, n12570, n12571, n12572,
         n12573, n12574, n12575, n12576, n12577, n12578, n12579, n12580,
         n12581, n12582, n12583, n12584, n12585, n12586, n12587, n12588,
         n12589, n12590, n12591, n12592, n12593, n12594, n12595, n12596,
         n12597, n12598, n12599, n12600, n12601, n12602, n12603, n12604,
         n12605, n12606, n12607, n12608, n12609, n12610, n12611, n12612,
         n12613, n12614, n12615, n12616, n12617, n12618, n12619, n12620,
         n12621, n12622, n12623, n12624, n12625, n12626, n12627, n12628,
         n12629, n12630, n12631, n12632, n12633, n12634, n12635, n12636,
         n12637, n12638, n12639, n12640, n12641, n12642, n12643, n12644,
         n12645, n12646, n12647, n12648, n12649, n12650, n12651, n12652,
         n12653, n12654, n12655, n12656, n12657, n12658, n12659, n12660,
         n12661, n12662, n12663, n12664, n12665, n12666, n12667, n12668,
         n12669, n12670, n12671, n12672, n12673, n12674, n12675, n12676,
         n12677, n12678, n12679, n12680, n12681, n12682, n12683, n12684,
         n12685, n12686, n12687, n12688, n12689, n12690, n12691, n12692,
         n12693, n12694, n12695, n12696, n12697, n12698, n12699, n12700,
         n12701, n12702, n12703, n12704, n12705, n12706, n12707, n12708,
         n12709, n12710, n12711, n12712, n12713, n12714, n12715, n12716,
         n12717, n12718, n12719, n12720, n12721, n12722, n12723, n12724,
         n12725, n12726, n12727, n12728, n12729, n12730, n12731, n12732,
         n12733, n12734, n12735, n12736, n12737, n12738, n12739, n12740,
         n12741, n12742, n12743, n12744, n12745, n12746, n12747, n12748,
         n12749, n12750, n12751, n12752, n12753, n12754, n12755, n12756,
         n12757, n12758, n12759, n12760, n12761, n12762, n12763, n12764,
         n12765, n12766, n12767, n12768, n12769, n12770, n12771, n12772,
         n12773, n12774, n12775, n12776, n12777, n12778, n12779, n12780,
         n12781, n12782, n12783, n12784, n12785, n12786, n12787, n12788,
         n12789, n12790, n12791, n12792, n12793, n12794, n12795, n12796,
         n12797, n12798, n12799, n12800, n12801, n12802, n12803, n12804,
         n12805, n12806, n12807, n12808, n12809, n12810, n12811, n12812,
         n12813, n12814, n12815, n12816, n12817, n12818, n12819, n12820,
         n12821, n12822, n12823, n12824, n12825, n12826, n12827, n12828,
         n12829, n12830, n12831, n12832, n12833, n12834, n12835, n12836,
         n12837, n12838, n12839, n12840, n12841, n12842, n12843, n12844,
         n12845, n12846, n12847, n12848, n12849, n12850, n12851, n12852,
         n12853, n12854, n12855, n12856, n12857, n12858, n12859, n12860,
         n12861, n12862, n12863, n12864, n12865, n12866, n12867, n12868,
         n12869, n12870, n12871, n12872, n12873, n12874, n12875, n12876,
         n12877, n12878, n12879, n12880, n12881, n12882, n12883, n12884,
         n12885, n12886, n12887, n12888, n12889, n12890, n12891, n12892,
         n12893, n12894, n12895, n12896, n12897, n12898, n12899, n12900,
         n12901, n12902, n12903, n12904, n12905, n12906, n12907, n12908,
         n12909, n12910, n12911, n12912, n12913, n12914, n12915, n12916,
         n12917, n12918, n12919, n12920, n12921, n12922, n12923, n12924,
         n12925, n12926, n12927, n12928, n12929, n12930, n12931, n12932,
         n12933, n12934, n12935, n12936, n12937, n12938, n12939, n12940,
         n12941, n12942, n12943, n12944, n12945, n12946, n12947, n12948,
         n12949, n12950, n12951, n12952, n12953, n12954, n12955, n12956,
         n12957, n12958, n12959, n12960, n12961, n12962, n12963, n12964,
         n12965, n12966, n12967, n12968, n12969, n12970, n12971, n12972,
         n12973, n12974, n12975, n12976, n12977, n12978, n12979, n12980,
         n12981, n12982, n12983, n12984, n12985, n12986, n12987, n12988,
         n12989, n12990, n12991, n12992, n12993, n12994, n12995, n12996,
         n12997, n12998, n12999, n13000, n13001, n13002, n13003, n13004,
         n13005, n13006, n13007, n13008, n13009, n13010, n13011, n13012,
         n13013, n13014, n13015, n13016, n13017, n13018, n13019, n13020,
         n13021, n13022, n13023, n13024, n13025, n13026, n13027, n13028,
         n13029, n13030, n13031, n13032, n13033, n13034, n13035, n13036,
         n13037, n13038, n13039, n13040, n13041, n13042, n13043, n13044,
         n13045, n13046, n13047, n13048, n13049, n13050, n13051, n13052,
         n13053, n13054, n13055, n13056, n13057, n13058, n13059, n13060,
         n13061, n13062, n13063, n13064, n13065, n13066, n13067, n13068,
         n13069, n13070, n13071, n13072, n13073, n13074, n13075, n13076,
         n13077, n13078, n13079, n13080, n13081, n13082, n13083, n13084,
         n13085, n13086, n13087, n13088, n13089, n13090, n13091, n13092,
         n13093, n13094, n13095, n13096, n13097, n13098, n13099, n13100,
         n13101, n13102, n13103, n13104, n13105, n13106, n13107, n13108,
         n13109, n13110, n13111, n13112, n13113, n13114, n13115, n13116,
         n13117, n13118, n13119, n13120, n13121, n13122, n13123, n13124,
         n13125, n13126, n13127, n13128, n13129, n13130, n13131, n13132,
         n13133, n13134, n13135, n13136, n13137, n13138, n13139, n13140,
         n13141, n13142, n13143, n13144, n13145, n13146, n13147, n13148,
         n13149, n13150, n13151, n13152, n13153, n13154, n13155, n13156,
         n13157, n13158, n13159, n13160, n13161, n13162, n13163, n13164,
         n13165, n13166, n13167, n13168, n13169, n13170, n13171, n13172,
         n13173, n13174, n13175, n13176, n13177, n13178, n13179, n13180,
         n13181, n13182, n13183, n13184, n13185, n13186, n13187, n13188,
         n13189, n13190, n13191, n13192, n13193, n13194, n13195, n13196,
         n13197, n13198, n13199, n13200, n13201, n13202, n13203, n13204,
         n13205, n13206, n13207, n13208, n13209, n13210, n13211, n13212,
         n13213, n13214, n13215, n13216, n13217, n13218, n13219, n13220,
         n13221, n13222, n13223, n13224, n13225, n13226, n13227, n13228,
         n13229, n13230, n13231, n13232, n13233, n13234, n13235, n13236,
         n13237, n13238, n13239, n13240, n13241, n13242, n13243, n13244,
         n13245, n13246, n13247, n13248, n13249, n13250, n13251, n13252,
         n13253, n13254, n13255, n13256, n13257, n13258, n13259, n13260,
         n13261, n13262, n13263, n13264, n13265, n13266, n13267, n13268,
         n13269, n13270, n13271, n13272, n13273, n13274, n13275, n13276,
         n13277, n13278, n13279, n13280, n13281, n13282, n13283, n13284,
         n13285, n13286, n13287, n13288, n13289, n13290, n13291, n13292,
         n13293, n13294, n13295, n13296, n13297, n13298, n13299, n13300,
         n13301, n13302, n13303, n13304, n13305, n13306, n13307, n13308,
         n13309, n13310, n13311, n13312, n13313, n13314, n13315, n13316,
         n13317, n13318, n13319, n13320, n13321, n13322, n13323, n13324,
         n13325, n13326, n13327, n13328, n13329, n13330, n13331, n13332,
         n13333, n13334, n13335, n13336, n13337, n13338, n13339, n13340,
         n13341, n13342, n13343, n13344, n13345, n13346, n13347, n13348,
         n13349, n13350, n13351, n13352, n13353, n13354, n13355, n13356,
         n13357, n13358, n13359, n13360, n13361, n13362, n13363, n13364,
         n13365, n13366, n13367, n13368, n13369, n13370, n13371, n13372,
         n13373, n13374, n13375, n13376, n13377, n13378, n13379, n13380,
         n13381, n13382, n13383, n13384, n13385, n13386, n13387, n13388,
         n13389, n13390, n13391, n13392, n13393, n13394, n13395, n13396,
         n13397, n13398, n13399, n13400, n13401, n13402, n13403, n13404,
         n13405, n13406, n13407, n13408, n13409, n13410, n13411, n13412,
         n13413, n13414, n13415, n13416, n13417, n13418, n13419, n13420,
         n13421, n13422, n13423, n13424, n13425, n13426, n13427, n13428,
         n13429, n13430, n13431, n13432, n13433, n13434, n13435, n13436,
         n13437, n13438, n13439, n13440, n13441, n13442, n13443, n13444,
         n13445, n13446, n13447, n13448, n13449, n13450, n13451, n13452,
         n13453, n13454, n13455, n13456, n13457, n13458, n13459, n13460,
         n13461, n13462, n13463, n13464, n13465, n13466, n13467, n13468,
         n13469, n13470, n13471, n13472, n13473, n13474, n13475, n13476,
         n13477, n13478, n13479, n13480, n13481, n13482, n13483, n13484,
         n13485, n13486, n13487, n13488, n13489, n13490, n13491, n13492,
         n13493, n13494, n13495, n13496, n13497, n13498, n13499, n13500,
         n13501, n13502, n13503, n13504, n13505, n13506, n13507, n13508,
         n13509, n13510, n13511, n13512, n13513, n13514, n13515, n13516,
         n13517, n13518, n13519, n13520, n13521, n13522, n13523, n13524,
         n13525, n13526, n13527, n13528, n13529, n13530, n13531, n13532,
         n13533, n13534, n13535, n13536, n13537, n13538, n13539, n13540,
         n13541, n13542, n13543, n13544, n13545, n13546, n13547, n13548,
         n13549, n13550, n13551, n13552, n13553, n13554, n13555, n13556,
         n13557, n13558, n13559, n13560, n13561, n13562, n13563, n13564,
         n13565, n13566, n13567, n13568, n13569, n13570, n13571, n13572,
         n13573, n13574, n13575, n13576, n13577, n13578, n13579, n13580,
         n13581, n13582, n13583, n13584, n13585, n13586, n13587, n13588,
         n13589, n13590, n13591, n13592, n13593, n13594, n13595, n13596,
         n13597, n13598, n13599, n13600, n13601, n13602, n13603, n13604,
         n13605, n13606, n13607, n13608, n13609, n13610, n13611, n13612,
         n13613, n13614, n13615, n13616, n13617, n13618, n13619, n13620,
         n13621, n13622, n13623, n13624, n13625, n13626, n13627, n13628,
         n13629, n13630, n13631, n13632, n13633, n13634, n13635, n13636,
         n13637, n13638, n13639, n13640, n13641, n13642, n13643, n13644,
         n13645, n13646, n13647, n13648, n13649, n13650, n13651, n13652,
         n13653, n13654, n13655, n13656, n13657, n13658, n13659, n13660,
         n13661, n13662, n13663, n13664, n13665, n13666, n13667, n13668,
         n13669, n13670, n13671, n13672, n13673, n13674, n13675, n13676,
         n13677, n13678, n13679, n13680, n13681, n13682, n13683, n13684,
         n13685, n13686, n13687, n13688, n13689, n13690, n13691, n13692,
         n13693, n13694, n13695, n13696, n13697, n13698, n13699, n13700,
         n13701, n13702, n13703, n13704, n13705, n13706, n13707, n13708,
         n13709, n13710, n13711, n13712, n13713, n13714, n13715, n13716,
         n13717, n13718, n13719, n13720, n13721, n13722, n13723, n13724,
         n13725, n13726, n13727, n13728, n13729, n13730, n13731, n13732,
         n13733, n13734, n13735, n13736, n13737, n13738, n13739, n13740,
         n13741, n13742, n13743, n13744, n13745, n13746, n13747, n13748,
         n13749, n13750, n13751, n13752, n13753, n13754, n13755, n13756,
         n13757, n13758, n13759, n13760, n13761, n13762, n13763, n13764,
         n13765, n13766, n13767, n13768, n13769, n13770, n13771, n13772,
         n13773, n13774, n13775, n13776, n13777, n13778, n13779, n13780,
         n13781, n13782, n13783, n13784, n13785, n13786, n13787, n13788,
         n13789, n13790, n13791, n13792, n13793, n13794, n13795, n13796,
         n13797, n13798, n13799, n13800, n13801, n13802, n13803, n13804,
         n13805, n13806, n13807, n13808, n13809, n13810, n13811, n13812,
         n13813, n13814, n13815, n13816, n13817, n13818, n13819, n13820,
         n13821, n13822, n13823, n13824, n13825, n13826, n13827, n13828,
         n13829, n13830, n13831, n13832, n13833, n13834, n13835, n13836,
         n13837, n13838, n13839, n13840, n13841, n13842, n13843, n13844,
         n13845, n13846, n13847, n13848, n13849, n13850, n13851, n13852,
         n13853, n13854, n13855, n13856, n13857, n13858, n13859, n13860,
         n13861, n13862, n13863, n13864, n13865, n13866, n13867, n13868,
         n13869, n13870, n13871, n13872, n13873, n13874, n13875, n13876,
         n13877, n13878, n13879, n13880, n13881, n13882, n13883, n13884,
         n13885, n13886, n13887, n13888, n13889, n13890, n13891, n13892,
         n13893, n13894, n13895, n13896, n13897, n13898, n13899, n13900,
         n13901, n13902, n13903, n13904, n13905, n13906, n13907, n13908,
         n13909, n13910, n13911, n13912, n13913, n13914, n13915, n13916,
         n13917, n13918, n13919, n13920, n13921, n13922, n13923, n13924,
         n13925, n13926, n13927, n13928, n13929, n13930, n13931, n13932,
         n13933, n13934, n13935, n13936, n13937, n13938, n13939, n13940,
         n13941, n13942, n13943, n13944, n13945, n13946, n13947, n13948,
         n13949, n13950, n13951, n13952, n13953, n13954, n13955, n13956,
         n13957, n13958, n13959, n13960, n13961, n13962, n13963, n13964,
         n13965, n13966, n13967, n13968, n13969, n13970, n13971, n13972,
         n13973, n13974, n13975, n13976, n13977, n13978, n13979, n13980,
         n13981, n13982, n13983, n13984, n13985, n13986, n13987, n13988,
         n13989, n13990, n13991, n13992, n13993, n13994, n13995, n13996,
         n13997, n13998, n13999, n14000, n14001, n14002, n14003, n14004,
         n14005, n14006, n14007, n14008, n14009, n14010, n14011, n14012,
         n14013, n14014, n14015, n14016, n14017, n14018, n14019, n14020,
         n14021, n14022, n14023, n14024, n14025, n14026, n14027, n14028,
         n14029, n14030, n14031, n14032, n14033, n14034, n14035, n14036,
         n14037, n14038, n14039, n14040, n14041, n14042, n14043, n14044,
         n14045, n14046, n14047, n14048, n14049, n14050, n14051, n14052,
         n14053, n14054, n14055, n14056, n14057, n14058, n14059, n14060,
         n14061, n14062, n14063, n14064, n14065, n14066, n14067, n14068,
         n14069, n14070, n14071, n14072, n14073, n14074, n14075, n14076,
         n14077, n14078, n14079, n14080, n14081, n14082, n14083, n14084,
         n14085, n14086, n14087, n14088, n14089, n14090, n14091, n14092,
         n14093, n14094, n14095, n14096, n14097, n14098, n14099, n14100,
         n14101, n14102, n14103, n14104, n14105, n14106, n14107, n14108,
         n14109, n14110, n14111, n14112, n14113, n14114, n14115, n14116,
         n14117, n14118, n14119, n14120, n14121, n14122, n14123, n14124,
         n14125, n14126, n14127, n14128, n14129, n14130, n14131, n14132,
         n14133, n14134, n14135, n14136, n14137, n14138, n14139, n14140,
         n14141, n14142, n14143, n14144, n14145, n14146, n14147, n14148,
         n14149, n14150, n14151, n14152, n14153, n14154, n14155, n14156,
         n14157, n14158, n14159, n14160, n14161, n14162, n14163, n14164,
         n14165, n14166, n14167, n14168, n14169, n14170, n14171, n14172,
         n14173, n14174, n14175, n14176, n14177, n14178, n14179, n14180,
         n14181, n14182, n14183, n14184, n14185, n14186, n14187, n14188,
         n14189, n14190, n14191, n14192, n14193, n14194, n14195, n14196,
         n14197, n14198, n14199, n14200, n14201, n14202, n14203, n14204,
         n14205, n14206, n14207, n14208, n14209, n14210, n14211, n14212,
         n14213, n14214, n14215, n14216, n14217, n14218, n14219, n14220,
         n14221, n14222, n14223, n14224, n14225, n14226, n14227, n14228,
         n14229, n14230, n14231, n14232, n14233, n14234, n14235, n14236,
         n14237, n14238, n14239, n14240, n14241, n14242, n14243, n14244,
         n14245, n14246, n14247, n14248, n14249, n14250, n14251, n14252,
         n14253, n14254, n14255, n14256, n14257, n14258, n14259, n14260,
         n14261, n14262, n14263, n14264, n14265, n14266, n14267, n14268,
         n14269, n14270, n14271, n14272, n14273, n14274, n14275, n14276,
         n14277, n14278, n14279, n14280, n14281, n14282, n14283, n14284,
         n14285, n14286, n14287, n14288, n14289, n14290, n14291, n14292,
         n14293, n14294, n14295, n14296, n14297, n14298, n14299, n14300,
         n14301, n14302, n14303, n14304, n14305, n14306, n14307, n14308,
         n14309, n14310, n14311, n14312, n14313, n14314, n14315, n14316,
         n14317, n14318, n14319, n14320, n14321, n14322, n14323, n14324,
         n14325, n14326, n14327, n14328, n14329, n14330, n14331, n14332,
         n14333, n14334, n14335, n14336, n14337, n14338, n14339, n14340,
         n14341, n14342, n14343, n14344, n14345, n14346, n14347, n14348,
         n14349, n14350, n14351, n14352, n14353, n14354, n14355, n14356,
         n14357, n14358, n14359, n14360, n14361, n14362, n14363, n14364,
         n14365, n14366, n14367, n14368, n14369, n14370, n14371, n14372,
         n14373, n14374, n14375, n14376, n14377, n14378, n14379, n14380,
         n14381, n14382, n14383, n14384, n14385, n14386, n14387, n14388,
         n14389, n14390, n14391, n14392, n14393, n14394, n14395, n14396,
         n14397, n14398, n14399, n14400, n14401, n14402, n14403, n14404,
         n14405, n14406, n14407, n14408, n14409, n14410, n14411, n14412,
         n14413, n14414, n14415, n14416, n14417, n14418, n14419, n14420,
         n14421, n14422, n14423, n14424, n14425, n14426, n14427, n14428,
         n14429, n14430, n14431, n14432, n14433, n14434, n14435, n14436,
         n14437, n14438, n14439, n14440, n14441, n14442, n14443, n14444,
         n14445, n14446, n14447, n14448, n14449, n14450, n14451, n14452,
         n14453, n14454, n14455, n14456, n14457, n14458, n14459, n14460,
         n14461, n14462, n14463, n14464, n14465, n14466, n14467, n14468,
         n14469, n14470, n14471, n14472, n14473, n14474, n14475, n14476,
         n14477, n14478, n14479, n14480, n14481, n14482, n14483, n14484,
         n14485, n14486, n14487, n14488, n14489, n14490, n14491, n14492,
         n14493, n14494, n14495, n14496, n14497, n14498, n14499, n14500,
         n14501, n14502, n14503, n14504, n14505, n14506, n14507, n14508,
         n14509, n14510, n14511, n14512, n14513, n14514, n14515, n14516,
         n14517, n14518, n14519, n14520, n14521, n14522, n14523, n14524,
         n14525, n14526, n14527, n14528, n14529, n14530, n14531, n14532,
         n14533, n14534, n14535, n14536, n14537, n14538, n14539, n14540,
         n14541, n14542, n14543, n14544, n14545, n14546, n14547, n14548,
         n14549, n14550, n14551, n14552, n14553, n14554, n14555, n14556,
         n14557, n14558, n14559, n14560, n14561, n14562, n14563, n14564,
         n14565, n14566, n14567, n14568, n14569, n14570, n14571, n14572,
         n14573, n14574, n14575, n14576, n14577, n14578, n14579, n14580,
         n14581, n14582, n14583, n14584, n14585, n14586, n14587, n14588,
         n14589, n14590, n14591, n14592, n14593, n14594, n14595, n14596,
         n14597, n14598, n14599, n14600, n14601, n14602, n14603, n14604,
         n14605, n14606, n14607, n14608, n14609, n14610, n14611, n14612,
         n14613, n14614, n14615, n14616, n14617, n14618, n14619, n14620,
         n14621, n14622, n14623, n14624, n14625, n14626, n14627, n14628,
         n14629, n14630, n14631, n14632, n14633, n14634, n14635, n14636,
         n14637, n14638, n14639, n14640, n14641, n14642, n14643, n14644,
         n14645, n14646, n14647, n14648, n14649, n14650, n14651, n14652,
         n14653, n14654, n14655, n14656, n14657, n14658, n14659, n14660,
         n14661, n14662, n14663, n14664, n14665, n14666, n14667, n14668,
         n14669, n14670, n14671, n14672, n14673, n14674, n14675, n14676,
         n14677, n14678, n14679, n14680, n14681, n14682, n14683, n14684,
         n14685, n14686, n14687, n14688, n14689, n14690, n14691, n14692,
         n14693, n14694, n14695, n14696, n14697, n14698, n14699, n14700,
         n14701, n14702, n14703, n14704, n14705, n14706, n14707, n14708,
         n14709, n14710, n14711, n14712, n14713, n14714, n14715, n14716,
         n14717, n14718, n14719, n14720, n14721, n14722, n14723, n14724,
         n14725, n14726, n14727, n14728, n14729, n14730, n14731, n14732,
         n14733, n14734, n14735, n14736, n14737, n14738, n14739, n14740,
         n14741, n14742, n14743, n14744, n14745, n14746, n14747, n14748,
         n14749, n14750, n14751, n14752, n14753, n14754, n14755, n14756,
         n14757, n14758, n14759, n14760, n14761, n14762, n14763, n14764,
         n14765, n14766, n14767, n14768, n14769, n14770, n14771, n14772,
         n14773, n14774, n14775, n14776, n14777, n14778, n14779, n14780,
         n14781, n14782, n14783, n14784, n14785, n14786, n14787, n14788,
         n14789, n14790, n14791, n14792, n14793, n14794, n14795, n14796,
         n14797, n14798, n14799, n14800, n14801, n14802, n14803, n14804,
         n14805, n14806, n14808, n14809, n14810, n14811, n14812, n14813,
         n14814, n14815, n14816, n14817, n14818, n14819, n14820, n14821,
         n14822, n14823, n14824, n14825, n14826, n14827, n14828, n14829,
         n14830, n14831, n14832, n14833, n14834, n14835, n14836, n14837,
         n14838, n14839, n14840, n14841, n14842, n14843, n14844, n14845,
         n14846, n14847, n14848, n14849, n14850, n14851, n14852, n14853,
         n14854, n14855, n14856, n14857, n14858, n14859, n14860, n14861,
         n14862, n14863, n14864, n14865, n14866, n14867, n14868, n14869,
         n14870, n14871, n14872, n14873, n14874, n14875, n14876, n14877,
         n14878, n14879, n14880, n14881, n14882, n14883, n14884, n14885,
         n14886, n14887, n14888, n14889, n14890, n14891, n14892, n14893,
         n14894, n14895, n14896, n14897, n14898, n14899, n14900, n14901,
         n14902, n14903, n14904, n14905, n14906, n14907, n14908, n14909,
         n14910, n14911, n14912, n14913, n14914, n14915, n14916, n14917,
         n14918, n14919, n14920, n14921, n14922, n14923, n14924, n14925,
         n14926, n14927, n14928, n14929, n14930, n14931, n14932, n14933,
         n14934, n14935, n14936, n14937, n14938, n14939, n14940, n14941,
         n14942, n14943, n14944, n14945, n14946, n14947, n14948, n14949,
         n14950, n14951, n14952, n14953, n14954, n14955, n14956, n14957,
         n14958, n14959, n14960, n14961, n14962, n14963, n14964, n14965,
         n14966, n14967, n14968, n14969, n14970, n14971, n14972, n14973,
         n14974, n14975, n14976, n14977, n14978, n14979, n14980, n14981,
         n14982, n14983, n14984, n14985, n14986, n14987, n14988, n14989,
         n14990, n14991, n14992, n14993, n14994, n14995, n14996, n14997,
         n14998, n14999, n15000, n15001, n15002, n15003, n15004, n15005,
         n15006, n15007, n15008, n15009, n15010, n15011, n15012, n15013,
         n15014, n15015, n15016, n15017, n15018, n15019, n15020, n15021,
         n15022, n15023, n15024, n15025, n15026, n15027, n15028, n15029,
         n15030, n15031, n15032, n15033, n15034, n15035, n15036, n15037,
         n15038, n15039, n15040, n15041, n15042, n15043, n15044, n15045,
         n15046, n15047, n15048, n15049, n15050, n15051, n15052, n15053,
         n15054, n15055, n15056, n15057, n15058, n15059, n15060, n15061,
         n15062, n15063, n15064, n15065, n15066, n15067, n15068, n15069,
         n15070, n15071, n15072, n15073, n15074, n15075, n15076, n15077,
         n15078, n15079, n15080, n15081, n15082, n15083, n15084, n15085,
         n15086, n15087, n15088, n15089, n15090, n15091, n15092, n15093,
         n15094, n15095, n15096, n15097, n15098, n15099, n15100, n15101,
         n15102, n15103, n15104, n15105, n15106, n15107, n15108, n15109,
         n15110, n15111, n15112, n15113, n15114, n15115, n15116, n15117,
         n15118, n15119, n15120, n15121, n15122, n15123, n15124, n15125,
         n15126, n15127, n15128, n15129, n15130, n15131, n15132, n15133,
         n15134, n15135, n15136, n15137, n15138, n15139, n15140, n15141,
         n15142, n15143, n15144, n15145, n15146, n15147, n15148, n15149,
         n15150, n15151, n15152, n15153, n15154, n15155, n15156, n15157,
         n15158, n15159, n15160, n15161, n15162, n15163, n15164, n15165,
         n15166, n15167, n15168, n15169, n15170, n15171, n15172, n15173,
         n15174, n15175, n15176, n15177, n15178, n15179, n15180, n15181,
         n15182, n15183, n15184, n15185, n15186, n15187, n15188, n15189,
         n15190, n15191, n15192, n15193, n15194, n15195, n15196, n15197,
         n15198, n15199, n15200, n15201, n15202, n15203, n15204, n15205,
         n15206, n15207, n15208, n15209, n15210, n15211, n15212, n15213,
         n15214, n15215, n15216, n15217, n15218, n15219, n15220, n15221,
         n15222, n15223, n15224, n15225, n15226, n15227, n15228, n15229,
         n15230, n15231, n15232, n15233, n15234, n15235, n15236, n15237,
         n15238, n15239, n15240, n15241, n15242, n15243, n15244, n15245,
         n15246, n15247, n15248, n15249, n15250, n15251, n15252, n15253,
         n15254, n15255, n15256, n15257, n15258, n15259, n15260, n15261,
         n15262, n15263, n15264, n15265, n15266, n15267, n15268, n15269,
         n15270, n15271, n15272, n15273, n15274, n15275, n15276, n15277,
         n15278, n15279, n15280, n15281, n15282, n15283, n15284, n15285,
         n15286, n15287, n15288, n15289, n15290, n15291, n15292, n15293,
         n15294, n15295, n15296, n15297, n15298, n15299, n15300, n15301,
         n15302, n15303, n15304, n15305, n15306, n15307, n15308, n15309,
         n15310, n15311, n15312, n15313, n15314, n15315, n15316, n15317,
         n15318, n15319, n15320, n15321, n15322, n15323, n15324, n15325,
         n15326, n15327, n15328, n15329, n15330, n15331, n15332, n15333,
         n15334, n15335, n15336, n15337, n15338, n15339, n15340, n15341,
         n15342, n15343, n15344, n15345, n15346, n15347, n15348, n15349,
         n15350, n15351, n15352, n15353, n15354, n15355, n15356, n15357,
         n15358, n15359, n15360, n15361, n15362, n15363, n15364, n15365,
         n15366, n15367, n15368, n15369, n15370, n15371, n15372, n15373,
         n15374, n15375, n15376, n15377, n15378, n15379, n15380, n15381,
         n15382, n15383, n15384, n15385, n15386, n15387, n15388, n15389,
         n15390, n15391, n15392, n15393, n15394, n15395, n15396, n15397,
         n15398, n15399, n15400, n15401, n15402, n15403, n15404, n15405,
         n15406, n15407, n15408, n15409, n15410, n15411, n15412, n15413,
         n15414, n15415, n15416, n15417, n15418, n15419, n15420, n15421,
         n15422, n15423, n15424, n15425, n15426, n15427, n15428, n15429,
         n15430, n15431, n15432, n15433, n15434, n15435, n15436, n15437,
         n15438, n15439, n15440, n15441, n15442, n15443, n15444, n15445,
         n15446, n15447, n15448, n15449, n15450, n15451, n15452, n15453,
         n15454, n15455, n15456, n15457, n15458, n15459, n15460, n15461,
         n15462, n15463, n15464, n15465, n15466, n15467, n15468, n15469,
         n15470, n15471, n15472, n15473, n15474, n15475, n15476, n15477,
         n15478, n15479, n15480, n15481, n15482, n15483, n15484, n15485,
         n15486, n15487, n15488, n15489, n15490, n15491, n15492, n15493,
         n15494, n15495, n15496, n15497, n15498, n15499, n15500, n15501,
         n15502, n15503, n15504, n15505, n15506, n15507, n15508, n15509,
         n15510, n15511, n15512, n15513, n15514, n15515, n15516, n15517,
         n15518, n15519, n15520, n15521, n15522, n15523, n15524, n15525,
         n15526, n15527, n15528, n15529, n15530, n15531, n15532, n15533,
         n15534, n15535, n15536, n15537, n15538, n15539, n15540, n15541,
         n15542, n15543, n15544, n15545, n15546, n15547, n15548, n15549,
         n15550, n15551, n15552, n15553, n15554, n15555, n15556, n15557,
         n15558, n15559, n15560, n15561, n15562, n15563, n15564, n15565,
         n15566, n15567, n15568, n15569, n15570, n15571, n15572, n15573,
         n15574, n15575, n15576, n15577, n15578, n15579, n15580, n15581,
         n15582, n15583, n15584, n15585, n15586, n15587, n15588, n15589,
         n15590, n15591, n15592, n15593, n15594, n15595, n15596, n15597,
         n15598, n15599, n15600, n15601, n15602, n15603, n15604, n15605,
         n15606, n15607, n15608, n15609, n15610, n15611, n15612, n15613,
         n15614, n15615, n15616, n15617, n15618, n15619, n15620, n15621,
         n15622, n15623, n15624, n15625, n15626, n15627, n15628, n15629,
         n15630, n15631, n15632, n15633, n15634, n15635, n15636, n15637,
         n15638, n15639, n15640, n15641, n15642, n15643, n15644, n15645,
         n15646, n15647, n15648, n15649, n15650, n15651, n15652, n15653,
         n15654, n15655, n15656, n15657, n15658, n15659, n15660, n15661,
         n15662, n15663, n15664, n15665, n15666, n15667, n15668, n15669,
         n15670, n15671, n15672, n15673, n15674, n15675, n15676, n15677,
         n15678, n15679, n15680, n15681, n15682, n15683, n15684, n15685,
         n15686, n15687, n15688, n15689, n15690, n15691, n15692, n15693,
         n15694, n15695, n15696, n15697, n15698, n15699, n15700, n15701,
         n15702, n15703, n15704, n15705, n15706, n15707, n15708, n15709,
         n15710, n15711, n15712, n15713, n15714, n15715, n15716, n15717,
         n15718, n15719, n15720, n15721, n15722, n15723, n15724, n15725,
         n15726, n15727, n15728, n15729, n15730, n15731, n15732, n15733,
         n15734, n15735, n15736, n15737, n15738, n15739, n15740, n15741,
         n15742, n15743, n15744, n15745, n15746, n15747, n15748, n15749,
         n15750, n15751, n15752, n15753, n15754, n15755, n15756, n15757,
         n15758, n15759, n15760, n15761, n15762, n15763, n15764, n15765,
         n15766, n15767, n15768, n15769, n15770, n15771, n15772, n15773,
         n15774, n15775, n15776, n15777, n15778, n15779, n15780, n15781,
         n15782, n15783, n15784, n15785, n15786, n15787, n15788, n15789,
         n15790, n15791, n15792, n15793, n15794, n15795, n15796, n15797,
         n15798, n15799, n15800, n15801, n15802, n15803, n15804, n15805,
         n15806, n15807, n15808, n15809, n15810, n15811, n15812, n15813,
         n15814, n15815, n15816, n15817, n15818, n15819, n15820, n15821,
         n15822, n15823, n15824, n15825, n15826, n15827, n15828, n15829,
         n15830, n15831, n15832, n15833, n15834, n15835, n15836, n15837,
         n15838, n15839, n15840, n15841, n15842, n15843, n15844, n15845,
         n15846, n15847, n15848, n15849, n15850, n15851, n15852, n15853,
         n15854, n15855, n15856, n15857, n15858, n15859, n15860, n15861,
         n15862, n15863, n15864, n15865, n15866, n15867, n15868, n15869,
         n15870, n15871, n15872, n15873, n15874, n15875, n15876, n15877,
         n15878, n15879, n15880, n15881, n15882, n15883, n15884, n15885,
         n15886, n15887, n15888, n15889, n15890, n15891, n15892, n15893,
         n15894, n15895, n15896, n15897, n15898, n15899, n15900, n15901,
         n15902, n15903, n15904, n15905, n15906, n15907, n15908, n15909,
         n15910, n15911, n15912, n15913, n15914, n15915, n15916, n15917,
         n15918, n15919, n15920, n15921, n15922, n15923, n15924, n15925,
         n15926, n15927, n15928, n15929, n15930, n15931, n15932, n15933,
         n15934, n15935, n15936, n15937, n15938, n15939, n15940, n15941,
         n15942, n15943, n15944, n15945, n15946, n15947, n15948, n15949,
         n15950, n15951, n15952, n15953, n15954, n15955, n15956, n15957,
         n15958, n15959, n15960, n15961, n15962, n15963, n15964, n15965,
         n15966, n15967, n15968, n15969, n15970, n15971, n15972, n15973,
         n15974, n15975, n15976, n15977, n15978, n15979, n15980, n15981,
         n15982, n15983, n15984, n15985, n15986, n15987, n15988, n15989,
         n15990, n15991, n15992, n15993, n15994, n15995, n15996, n15997,
         n15998, n15999, n16000, n16001, n16002, n16003, n16004, n16005,
         n16006, n16007, n16008, n16009, n16010, n16011, n16012, n16013,
         n16014, n16015, n16016, n16017, n16018, n16019, n16020, n16021,
         n16022, n16023, n16024, n16025, n16026, n16027, n16028, n16029,
         n16030, n16031, n16032, n16033, n16034, n16035, n16036, n16037,
         n16038, n16039, n16040, n16041, n16042, n16043, n16044, n16045,
         n16046, n16047, n16048, n16049, n16050, n16051, n16052, n16053,
         n16054, n16055, n16056, n16057, n16058, n16059, n16060, n16061,
         n16062, n16063, n16064, n16065, n16066, n16067, n16068, n16069,
         n16070, n16071, n16072, n16073, n16074, n16075, n16076, n16077,
         n16078, n16079, n16080, n16081, n16082, n16083, n16084, n16085,
         n16086, n16087, n16088, n16089, n16090, n16091, n16092, n16093,
         n16094, n16095, n16096, n16097, n16098, n16099, n16100, n16101,
         n16102, n16103, n16104, n16105, n16106, n16107, n16108, n16109,
         n16110, n16111, n16112, n16113, n16114, n16115, n16116, n16117,
         n16118, n16119, n16120, n16121, n16122, n16123, n16124, n16126,
         n16127, n16128, n16129, n16130, n16131, n16132, n16133, n16134,
         n16135, n16136, n16137, n16138, n16139, n16140, n16141, n16142,
         n16143, n16144, n16145, n16146, n16147, n16148, n16149, n16150,
         n16151, n16152, n16153, n16154, n16155, n16156, n16157, n16158,
         n16159, n16160, n16161, n16162, n16163, n16164, n16165, n16166,
         n16167, n16168, n16169, n16170, n16171, n16172, n16173, n16174,
         n16175, n16176, n16177, n16178, n16179, n16180, n16181, n16182,
         n16183, n16184, n16185, n16186, n16187, n16188, n16189, n16190,
         n16191, n16192, n16193, n16194, n16195, n16196, n16197, n16198,
         n16199, n16200, n16201, n16202, n16203, n16204, n16205, n16206,
         n16207, n16208, n16209, n16210, n16211, n16212, n16213, n16214,
         n16215, n16216, n16217, n16218, n16219, n16220, n16221, n16222,
         n16223, n16224, n16225, n16226, n16227, n16228, n16229, n16230,
         n16231, n16232, n16233, n16234, n16235, n16236, n16237, n16238,
         n16239, n16240, n16241, n16242, n16243, n16244, n16245, n16246,
         n16247, n16248, n16249, n16250, n16251, n16252, n16253, n16254,
         n16255, n16256, n16257, n16258, n16259, n16260, n16261, n16262,
         n16263, n16264, n16265, n16266, n16267, n16268, n16269, n16270,
         n16271, n16272, n16273, n16274, n16275, n16276, n16277, n16278,
         n16279, n16280, n16281, n16282, n16283, n16284, n16285, n16286,
         n16287, n16288, n16289, n16290, n16291, n16292, n16293, n16294,
         n16295, n16296, n16297, n16298, n16299, n16300, n16301, n16302,
         n16303, n16304, n16305, n16306, n16307, n16308, n16309, n16310,
         n16311, n16312, n16313, n16314, n16315, n16316, n16317, n16318,
         n16319, n16320, n16321, n16322, n16323, n16324, n16325, n16326,
         n16327, n16328, n16329, n16330, n16331, n16332, n16333, n16334,
         n16335, n16336, n16337, n16338, n16339, n16340, n16341, n16342,
         n16343, n16344, n16345, n16346, n16347, n16348, n16349, n16350,
         n16351, n16352, n16353, n16354, n16355, n16356, n16357, n16358,
         n16359, n16360, n16361, n16362, n16363, n16364, n16365, n16366,
         n16367, n16368, n16369, n16370, n16371, n16372, n16373, n16374,
         n16375, n16376, n16377, n16378, n16379, n16380, n16381, n16382,
         n16383, n16384, n16385, n16386, n16387, n16388, n16389, n16390,
         n16391, n16392, n16393, n16394, n16395, n16396, n16397, n16398,
         n16399, n16400, n16401, n16402, n16403, n16404, n16405, n16406,
         n16407, n16408, n16409, n16410, n16411, n16412, n16413, n16414,
         n16415, n16416, n16417, n16418, n16419, n16420, n16421, n16422,
         n16423, n16424, n16425, n16426, n16427, n16428, n16429, n16430,
         n16431, n16432, n16433, n16434, n16435, n16436, n16437, n16438,
         n16439, n16440, n16441, n16442, n16443, n16444, n16445, n16446,
         n16447, n16448, n16449, n16450, n16451, n16452, n16453, n16454,
         n16455, n16456, n16457, n16458, n16459, n16460, n16461, n16462,
         n16463, n16464, n16465, n16466, n16467, n16468, n16469, n16470,
         n16471, n16472, n16473, n16474, n16475, n16476, n16477, n16478,
         n16479, n16480, n16481, n16482, n16483, n16484, n16485, n16486,
         n16487, n16488, n16489, n16490, n16491, n16492, n16493, n16494,
         n16495, n16496, n16497, n16498, n16499, n16500, n16501, n16502,
         n16503, n16504, n16505, n16506, n16507, n16508, n16509, n16510,
         n16511, n16512, n16513, n16514, n16515, n16516, n16517, n16518,
         n16519, n16520, n16521, n16522, n16523, n16524, n16525, n16526,
         n16527, n16528, n16529, n16530, n16531, n16532, n16533, n16534,
         n16535, n16536, n16537, n16538, n16539, n16540, n16541, n16542,
         n16543, n16544, n16545, n16546, n16547, n16548, n16549, n16550,
         n16551, n16552, n16553, n16554, n16555, n16556, n16557, n16558,
         n16559, n16560, n16561, n16562, n16563, n16564, n16565, n16566,
         n16567, n16568, n16569, n16570, n16571, n16572, n16573, n16574,
         n16575, n16576, n16577, n16578, n16579, n16580, n16581, n16582,
         n16583, n16584, n16585, n16586, n16587, n16588, n16589, n16590,
         n16591, n16592, n16593, n16594, n16595, n16596, n16597, n16598,
         n16599, n16600, n16601, n16602, n16603, n16604, n16605, n16606,
         n16607, n16608, n16609, n16610, n16611, n16612, n16613, n16614,
         n16615, n16616, n16617, n16618, n16619, n16620, n16621, n16622,
         n16623, n16624, n16625, n16626, n16627, n16628, n16629, n16630,
         n16631, n16632, n16633, n16634, n16635, n16636, n16637, n16638,
         n16639, n16640, n16641, n16642, n16643, n16644, n16645, n16646,
         n16647, n16648, n16649, n16650, n16651, n16652, n16653, n16654,
         n16655, n16656, n16657, n16658, n16659, n16660, n16661, n16662,
         n16663, n16664, n16665, n16666, n16667, n16668, n16669, n16670,
         n16671, n16672, n16673, n16674, n16675, n16676, n16677, n16678,
         n16679, n16680, n16681, n16682, n16683, n16684, n16685, n16686,
         n16687, n16688, n16689, n16690, n16691, n16692, n16693, n16694,
         n16695, n16696, n16697, n16698, n16699, n16700, n16701, n16702,
         n16703, n16704, n16705, n16706, n16707, n16708, n16709, n16710,
         n16711, n16712, n16713, n16714, n16715, n16716, n16717, n16718,
         n16719, n16720, n16721, n16722, n16723, n16724, n16725, n16726,
         n16727, n16728, n16729, n16730, n16731, n16732, n16733, n16734,
         n16735, n16736, n16737, n16738, n16739, n16740, n16741, n16742,
         n16743, n16744, n16745, n16746, n16747, n16748, n16749, n16750,
         n16751, n16752, n16753, n16754, n16755, n16756, n16757, n16758,
         n16759, n16760, n16761, n16762, n16763, n16764, n16765, n16766,
         n16767, n16768, n16769, n16770, n16771, n16772, n16773, n16774,
         n16775, n16776, n16777, n16778, n16779, n16780, n16781, n16782,
         n16783, n16784, n16785, n16786, n16787, n16788, n16789, n16790,
         n16791, n16792, n16793, n16794, n16795, n16796, n16797, n16798,
         n16799, n16800, n16801, n16802, n16803, n16804, n16805, n16806,
         n16807, n16808, n16809, n16810, n16811, n16812, n16813, n16814,
         n16815, n16816, n16817, n16818, n16819, n16820, n16821, n16822,
         n16823, n16824, n16825, n16826, n16827, n16828, n16829, n16830,
         n16831, n16832, n16833, n16834, n16835, n16836, n16837, n16838,
         n16839, n16840, n16841, n16842, n16843, n16844, n16845, n16846,
         n16847, n16848, n16849, n16850, n16851, n16852, n16853, n16854,
         n16855, n16856, n16857, n16858, n16859, n16860, n16861, n16862,
         n16863, n16864, n16865, n16866, n16867, n16868, n16869, n16870,
         n16871, n16872, n16873, n16874, n16875, n16876, n16877, n16878,
         n16879, n16880, n16881, n16882, n16883, n16884, n16885, n16886,
         n16887, n16888, n16889, n16890, n16891, n16892, n16893, n16894,
         n16895, n16896, n16897, n16898, n16899, n16900, n16901, n16902,
         n16903, n16904, n16905, n16906, n16907, n16908, n16909, n16910,
         n16911, n16912, n16913, n16914, n16915, n16916, n16917, n16918,
         n16919, n16920, n16921, n16922, n16923, n16924, n16925, n16926,
         n16927, n16928, n16929, n16930, n16931, n16932, n16933, n16934,
         n16935, n16936, n16937, n16938, n16939, n16940, n16941, n16942,
         n16943, n16944, n16945, n16946, n16947, n16948, n16949, n16950,
         n16951, n16952, n16953, n16954, n16955, n16956, n16957, n16958,
         n16959, n16960, n16961, n16962, n16963, n16964, n16965, n16966,
         n16967, n16968, n16969, n16970, n16971, n16972, n16973, n16974,
         n16975, n16976, n16977, n16978, n16979, n16980, n16981, n16982,
         n16983, n16984, n16985, n16986, n16987, n16988, n16989, n16990,
         n16991, n16992, n16993, n16994, n16995, n16996, n16997, n16998,
         n16999, n17000, n17001, n17002, n17003, n17004, n17005, n17006,
         n17007, n17008, n17009, n17010, n17011, n17012, n17013, n17014,
         n17015, n17016, n17017, n17018, n17019, n17020, n17021, n17022,
         n17023, n17024, n17025, n17026, n17027, n17028, n17029, n17030,
         n17031, n17032, n17033, n17034, n17035, n17036, n17037, n17038,
         n17039, n17040, n17041, n17042, n17043, n17044, n17045, n17046,
         n17047, n17048, n17049, n17050, n17051, n17052, n17053, n17054,
         n17055, n17056, n17057, n17058, n17059, n17060, n17061, n17062,
         n17063, n17064, n17065, n17066, n17067, n17068, n17069, n17070,
         n17071, n17072, n17073, n17074, n17075, n17076, n17077, n17078,
         n17079, n17080, n17081, n17082, n17083, n17084, n17085, n17086,
         n17087, n17088, n17089, n17090, n17091, n17092, n17093, n17094,
         n17095, n17096, n17097, n17098, n17099, n17100, n17101, n17102,
         n17103, n17104, n17105, n17106, n17107, n17108, n17109, n17110,
         n17111, n17112, n17113, n17114, n17115, n17116, n17117, n17118,
         n17119, n17120, n17121, n17122, n17123, n17124, n17125, n17126,
         n17127, n17128, n17129, n17130, n17131, n17132, n17133, n17134,
         n17135, n17136, n17137, n17138, n17139, n17140, n17141, n17142,
         n17143, n17144, n17145, n17146, n17147, n17148, n17149, n17150,
         n17151, n17152, n17153, n17154, n17155, n17156, n17157, n17158,
         n17159, n17160, n17161, n17162, n17163, n17164, n17165, n17166,
         n17167, n17168, n17169, n17170, n17171, n17172, n17173, n17174,
         n17175, n17176, n17177, n17178, n17179, n17180, n17181, n17182,
         n17183, n17184, n17185, n17186, n17187, n17188, n17189, n17190,
         n17191, n17192, n17193, n17194, n17195, n17196, n17197, n17198,
         n17199, n17200, n17201, n17202, n17203, n17204, n17205, n17206,
         n17207, n17208, n17209, n17210, n17211, n17212, n17213, n17214,
         n17215, n17216, n17217, n17218, n17219, n17220, n17221, n17222,
         n17223, n17224, n17225, n17226, n17227, n17228, n17229, n17230,
         n17231, n17232, n17233, n17234, n17235, n17236, n17237, n17238,
         n17239, n17240, n17241, n17242, n17243, n17244, n17245, n17246,
         n17247, n17248, n17249, n17250, n17251, n17252, n17253, n17254,
         n17255, n17256, n17257, n17258, n17259, n17260, n17261, n17262,
         n17263, n17264, n17265, n17266, n17267, n17268, n17269, n17270,
         n17271, n17272, n17273, n17274, n17275, n17276, n17277, n17278,
         n17279, n17280, n17281, n17282, n17283, n17284, n17285, n17286,
         n17287, n17288, n17289, n17290, n17291, n17292, n17293, n17294,
         n17295, n17296, n17297, n17298, n17299, n17300, n17301, n17302,
         n17303, n17304, n17305, n17306, n17307, n17308, n17309, n17310,
         n17311, n17312, n17313, n17314, n17315, n17316, n17317, n17318,
         n17319, n17320, n17321, n17322, n17323, n17324, n17325, n17326,
         n17327, n17328, n17329, n17330, n17331, n17332, n17333, n17334,
         n17335, n17336, n17337, n17338, n17339, n17340, n17341, n17342,
         n17343, n17344, n17345, n17346, n17347, n17348, n17349, n17350,
         n17351, n17352, n17353, n17354, n17355, n17356, n17357, n17358,
         n17359, n17360, n17361, n17362, n17363, n17364, n17365, n17366,
         n17367, n17368, n17369, n17370, n17371, n17372, n17373, n17374,
         n17375, n17376, n17377, n17378, n17379, n17380, n17381, n17382,
         n17383, n17384, n17385, n17386, n17387, n17388, n17389, n17390,
         n17391, n17392, n17393, n17394, n17395, n17396, n17397, n17398,
         n17399, n17400, n17401, n17402, n17403, n17404, n17405, n17406,
         n17407, n17408, n17409, n17410, n17411, n17412, n17413, n17414,
         n17415, n17416, n17417, n17418, n17419, n17420, n17421, n17422,
         n17423, n17424, n17425, n17426, n17427, n17428, n17429, n17430,
         n17431, n17432, n17433, n17434, n17435, n17436, n17437, n17438,
         n17439, n17440, n17441, n17442, n17443, n17444, n17445, n17446,
         n17447, n17448, n17449, n17450, n17451, n17452, n17453, n17454,
         n17455, n17456, n17457, n17458, n17459, n17460, n17461, n17462,
         n17463, n17464, n17465, n17466, n17467, n17468, n17469, n17470,
         n17471, n17472, n17473, n17474, n17475, n17476, n17477, n17478,
         n17479, n17480, n17481, n17482, n17483, n17484, n17485, n17486,
         n17487, n17488, n17489, n17490, n17491, n17492, n17493, n17494,
         n17495, n17496, n17497, n17498, n17499, n17500, n17501, n17502,
         n17503, n17504, n17505, n17506, n17507, n17508, n17509, n17510,
         n17511, n17512, n17513, n17514, n17515, n17516, n17517, n17518,
         n17519, n17520, n17521, n17522, n17523, n17524, n17525, n17526,
         n17527, n17528, n17529, n17530, n17531, n17532, n17533, n17534,
         n17535, n17536, n17537, n17538, n17539, n17540, n17541, n17542,
         n17543, n17544, n17545, n17546, n17547, n17548, n17549, n17550,
         n17551, n17552, n17553, n17554, n17555, n17556, n17557, n17558,
         n17559, n17560, n17561, n17562, n17563, n17564, n17565, n17566,
         n17567, n17568, n17569, n17570, n17571, n17572, n17573, n17574,
         n17575, n17576, n17577, n17578, n17579, n17580, n17581, n17582,
         n17583, n17584, n17585, n17586, n17587, n17588, n17589, n17590,
         n17591, n17592, n17593, n17594, n17595, n17596, n17597, n17598,
         n17599, n17600, n17601, n17602, n17603, n17604, n17605, n17606,
         n17607, n17608, n17609, n17610, n17611, n17612, n17613, n17614,
         n17615, n17616, n17617, n17618, n17619, n17620, n17621, n17622,
         n17623, n17624, n17625, n17626, n17627, n17628, n17629, n17630,
         n17631, n17632, n17633, n17634, n17635, n17636, n17637, n17638,
         n17639, n17640, n17641, n17642, n17643, n17644, n17645, n17646,
         n17647, n17648, n17649, n17650, n17651, n17652, n17653, n17654,
         n17655, n17656, n17657, n17658, n17659, n17660, n17661, n17662,
         n17663, n17664, n17665, n17666, n17667, n17668, n17669, n17670,
         n17671, n17672, n17673, n17674, n17675, n17676, n17677, n17678,
         n17679, n17680, n17681, n17682, n17683, n17684, n17685, n17686,
         n17687, n17688, n17689, n17690, n17691, n17692, n17693, n17694,
         n17695, n17696, n17697, n17698, n17699, n17700, n17701, n17702,
         n17703, n17704, n17705, n17706, n17707, n17708, n17709, n17710,
         n17711, n17712, n17713, n17714, n17715, n17716, n17717, n17718,
         n17719, n17720, n17721, n17722, n17723, n17724, n17725, n17726,
         n17727, n17728, n17729, n17730, n17731, n17732, n17733, n17734,
         n17735, n17736, n17737, n17738, n17739, n17740, n17741, n17742,
         n17743, n17744, n17745, n17746, n17747, n17748, n17749, n17750,
         n17751, n17752, n17753, n17754, n17755, n17756, n17757, n17758,
         n17759, n17760, n17761, n17762, n17763, n17764, n17765, n17766,
         n17767, n17768, n17769, n17770, n17771, n17772, n17773, n17774,
         n17775, n17776, n17777, n17778, n17779, n17780, n17781, n17782,
         n17783, n17784, n17785, n17786, n17787, n17788, n17789, n17790,
         n17791, n17792, n17793, n17794, n17795, n17796, n17797, n17798,
         n17799, n17800, n17801, n17802, n17803, n17804, n17805, n17806,
         n17807, n17808, n17809, n17810, n17811, n17812, n17813, n17814,
         n17815, n17816, n17817, n17818, n17819, n17820, n17821, n17822,
         n17823, n17824, n17825, n17826, n17827, n17828, n17829, n17830,
         n17831, n17832, n17833, n17834, n17835, n17836, n17837, n17838,
         n17839, n17840, n17841, n17842, n17843, n17844, n17845, n17846,
         n17847, n17848, n17849, n17850, n17851, n17852, n17853, n17854,
         n17855, n17856, n17857, n17858, n17859, n17860, n17861, n17862,
         n17863, n17864, n17865, n17866, n17867, n17868, n17869, n17870,
         n17871, n17872, n17873, n17874, n17875, n17876, n17877, n17878,
         n17879, n17880, n17881, n17882, n17883, n17884, n17885, n17886,
         n17887, n17888, n17889, n17890, n17891, n17892, n17893, n17894,
         n17895, n17896, n17897, n17898, n17899, n17900, n17901, n17902,
         n17903, n17904, n17905, n17906, n17907, n17908, n17909, n17910,
         n17911, n17912, n17913, n17914, n17915, n17916, n17917, n17918,
         n17919, n17920, n17921, n17922, n17923, n17924, n17925, n17926,
         n17927, n17928, n17929, n17930, n17931, n17932, n17933, n17934,
         n17935, n17936, n17937, n17938, n17939, n17940, n17941, n17942,
         n17943, n17944, n17945, n17946, n17947, n17948, n17949, n17950,
         n17951, n17952, n17953, n17954, n17955, n17956, n17957, n17958,
         n17959, n17960, n17961, n17962, n17963, n17964, n17965, n17966,
         n17967, n17968, n17969, n17970, n17971, n17972, n17973, n17974,
         n17975, n17976, n17977, n17978, n17979, n17980, n17981, n17982,
         n17983, n17984, n17985, n17986, n17987, n17988, n17989, n17990,
         n17991, n17992, n17993, n17994, n17995, n17996, n17997, n17998,
         n17999, n18000, n18001, n18002, n18003, n18004, n18005, n18006,
         n18007, n18008, n18009, n18010, n18011, n18012, n18013, n18014,
         n18015, n18016, n18017, n18018, n18019, n18020, n18021, n18022,
         n18023, n18024, n18025, n18026, n18027, n18028, n18029, n18030,
         n18031, n18032, n18033, n18034, n18035, n18036, n18037, n18038,
         n18039, n18040, n18041, n18042, n18043, n18044, n18045, n18046,
         n18047, n18048, n18049, n18050, n18051, n18052, n18053, n18054,
         n18055, n18056, n18057, n18058, n18059, n18060, n18061, n18062,
         n18063, n18064, n18065, n18066, n18067, n18068, n18069, n18070,
         n18071, n18072, n18073, n18074, n18075, n18076, n18077, n18078,
         n18079, n18080, n18081, n18082, n18083, n18084, n18085, n18086,
         n18087, n18088, n18089, n18090, n18091, n18092, n18093, n18094,
         n18095, n18096, n18097, n18098, n18099, n18100, n18101, n18102,
         n18103, n18104, n18105, n18106, n18107, n18108, n18109, n18110,
         n18111, n18112, n18113, n18114, n18115, n18116, n18117, n18118,
         n18119, n18120, n18121, n18122, n18123, n18124, n18125, n18126,
         n18127, n18128, n18129, n18130, n18131, n18132, n18133, n18134,
         n18135, n18136, n18137, n18138, n18139, n18140, n18141, n18142,
         n18143, n18144, n18145, n18146, n18147, n18148, n18149, n18150,
         n18151, n18152, n18153, n18154, n18155, n18156, n18157, n18158,
         n18159, n18160, n18161, n18162, n18163, n18164, n18165, n18166,
         n18167, n18168, n18169, n18170, n18171, n18172, n18173, n18174,
         n18175, n18176, n18177, n18178, n18179, n18180, n18181, n18182,
         n18183, n18184, n18185, n18186, n18187, n18188, n18189, n18190,
         n18191, n18192, n18193, n18194, n18195, n18196, n18197, n18198,
         n18199, n18200, n18201, n18202, n18203, n18204, n18205, n18206,
         n18207, n18208, n18209, n18210, n18211, n18212, n18213, n18214,
         n18215, n18216, n18217, n18218, n18219, n18220, n18221, n18222,
         n18223, n18224, n18225, n18226, n18227, n18228, n18229, n18230,
         n18231, n18232, n18233, n18234, n18235, n18236, n18237, n18238,
         n18239, n18240, n18241, n18242, n18243, n18244, n18245, n18246,
         n18247, n18248, n18249, n18250, n18251, n18252, n18253, n18254,
         n18255, n18256, n18257, n18258, n18259, n18260, n18261, n18262,
         n18263, n18264, n18265, n18266, n18267, n18268, n18269, n18270,
         n18271, n18272, n18273, n18274, n18275, n18276, n18277, n18278,
         n18279, n18280, n18281, n18282, n18283, n18284, n18285, n18286,
         n18287, n18288, n18289, n18290, n18291, n18292, n18293, n18294,
         n18295, n18296, n18297, n18298, n18299, n18300, n18301, n18302,
         n18303, n18304, n18305, n18306, n18307, n18308, n18309, n18310,
         n18311, n18312, n18313, n18314, n18315, n18316, n18317, n18318,
         n18319, n18320, n18321, n18322, n18323, n18324, n18325, n18326,
         n18327, n18328, n18329, n18330, n18331, n18332, n18333, n18334,
         n18335, n18336, n18337, n18338, n18339, n18340, n18341, n18342,
         n18343, n18344, n18345, n18346, n18347, n18348, n18349, n18350,
         n18351, n18352, n18353, n18354, n18355, n18356, n18357, n18358,
         n18359, n18360, n18361, n18362, n18363, n18364, n18365, n18366,
         n18367, n18368, n18369, n18370, n18371, n18372, n18373, n18374,
         n18375, n18376, n18377, n18378, n18379, n18380, n18381, n18382,
         n18383, n18384, n18385, n18386, n18387, n18388, n18389, n18390,
         n18391, n18392, n18393, n18394, n18395, n18396, n18397, n18398,
         n18399, n18400, n18401, n18402, n18403, n18404, n18405, n18406,
         n18407, n18408, n18409, n18410, n18411, n18412, n18413, n18414,
         n18415, n18416, n18417, n18418, n18419, n18420, n18421, n18422,
         n18423, n18424, n18425, n18426, n18427, n18428, n18429, n18430,
         n18431, n18432, n18433, n18434, n18435, n18436, n18437, n18438,
         n18439, n18440, n18441, n18442, n18443, n18444, n18445, n18446,
         n18447, n18448, n18449, n18450, n18451, n18452, n18453, n18454,
         n18455, n18456, n18457, n18458, n18459, n18460, n18461, n18462,
         n18463, n18464, n18465, n18466, n18467, n18468, n18469, n18470,
         n18471, n18472, n18473, n18474, n18475, n18476, n18477, n18478,
         n18479, n18480, n18481, n18482, n18483, n18484, n18485, n18486,
         n18487, n18488, n18489, n18490, n18491, n18492, n18493, n18494,
         n18495, n18496, n18497, n18498, n18499, n18500, n18501, n18502,
         n18503, n18504, n18505, n18506, n18507, n18508, n18509, n18510,
         n18511, n18512, n18513, n18514, n18515, n18516, n18517, n18518,
         n18519, n18520, n18521, n18522, n18523, n18524, n18525, n18526,
         n18527, n18528, n18529, n18530, n18531, n18532, n18533, n18534,
         n18535, n18536, n18537, n18538, n18539, n18540, n18541, n18542,
         n18543, n18544, n18545, n18546, n18547, n18548, n18549, n18550,
         n18551, n18552, n18553, n18554, n18555, n18556, n18557, n18558,
         n18559, n18560, n18561, n18562, n18563, n18564, n18565, n18566,
         n18567, n18568, n18569, n18570, n18571, n18572, n18573, n18574,
         n18575, n18576, n18577, n18578, n18579, n18580, n18581, n18582,
         n18583, n18584, n18585, n18586, n18587, n18588, n18589, n18590,
         n18591, n18592, n18593, n18594, n18595, n18596, n18597, n18598,
         n18599, n18600, n18601, n18602, n18603, n18604, n18605, n18606,
         n18607, n18608, n18609, n18610, n18611, n18612, n18613, n18614,
         n18615, n18616, n18617, n18618, n18619, n18620, n18621, n18622,
         n18623, n18624, n18625, n18626, n18627, n18628, n18629, n18630,
         n18631, n18632, n18633, n18634, n18635, n18636, n18637, n18638,
         n18639, n18640, n18641, n18642, n18643, n18644, n18645, n18646,
         n18647, n18648, n18649, n18650, n18651, n18652, n18653, n18654,
         n18655, n18656, n18657, n18658, n18659, n18660, n18661, n18662,
         n18663, n18664, n18665, n18666, n18667, n18668, n18669, n18670,
         n18671, n18672, n18673, n18674, n18675, n18676, n18677, n18678,
         n18679, n18680, n18681, n18682, n18683, n18684, n18685, n18686,
         n18687, n18688, n18689, n18690, n18691, n18692, n18693, n18694,
         n18695, n18696, n18697, n18698, n18699, n18700, n18701, n18702,
         n18703, n18704, n18705, n18706, n18707, n18708, n18709, n18710,
         n18711, n18712, n18713, n18714, n18715, n18716, n18717, n18718,
         n18719, n18720, n18721, n18722, n18723, n18724, n18725, n18726,
         n18727, n18728, n18729, n18730, n18731, n18732, n18733, n18734,
         n18735, n18736, n18737, n18738, n18739, n18740, n18741, n18742,
         n18743, n18744, n18745, n18746, n18747, n18748, n18749, n18750,
         n18751, n18752, n18753, n18754, n18755, n18756, n18757, n18758,
         n18759, n18760, n18761, n18762, n18763, n18764, n18765, n18766,
         n18767, n18768, n18769, n18770, n18771, n18772, n18773, n18774,
         n18775, n18776, n18777, n18778, n18779, n18780, n18781, n18782,
         n18783, n18784, n18785, n18786, n18787, n18788, n18789, n18790,
         n18791, n18792, n18793, n18794, n18795, n18796, n18797, n18798,
         n18799, n18800, n18801, n18802, n18803, n18804, n18805, n18806,
         n18807, n18808, n18809, n18810, n18811, n18812, n18813, n18814,
         n18815, n18816, n18817, n18818, n18819, n18820, n18821, n18822,
         n18823, n18824, n18825, n18826, n18827, n18828, n18829, n18830,
         n18831, n18832, n18833, n18834, n18835, n18836, n18837, n18838,
         n18839, n18840, n18841, n18842, n18843, n18844, n18845, n18846,
         n18847, n18848, n18849, n18850, n18851, n18852, n18853, n18854,
         n18855, n18856, n18857, n18858, n18859, n18860, n18861, n18862,
         n18863, n18864, n18865, n18866, n18867, n18868, n18869, n18870,
         n18871, n18872, n18873, n18874, n18875, n18876, n18877, n18878,
         n18879, n18880, n18881, n18882, n18883, n18884, n18885, n18886,
         n18887, n18888, n18889, n18890, n18891, n18892, n18893, n18894,
         n18895, n18896, n18897, n18898, n18899, n18900, n18901, n18902,
         n18903, n18904, n18905, n18906, n18907, n18908, n18909, n18910,
         n18911, n18912, n18913, n18914, n18915, n18916, n18917, n18918,
         n18919, n18920, n18921, n18922, n18923, n18924, n18925, n18926,
         n18927, n18928, n18929, n18930, n18931, n18932, n18933, n18934,
         n18935, n18936, n18937, n18938, n18939, n18940, n18941, n18942,
         n18943, n18944, n18945, n18946, n18947, n18948, n18949, n18950,
         n18951, n18952, n18953, n18954, n18955, n18956, n18957, n18958,
         n18959, n18960, n18961, n18962, n18963, n18964, n18965, n18966,
         n18967, n18968, n18969, n18970, n18971, n18972, n18973, n18974,
         n18975, n18976, n18977, n18978, n18979, n18980, n18981, n18982,
         n18983, n18984, n18985, n18986, n18987, n18988, n18989, n18990,
         n18991, n18992, n18993, n18994, n18995, n18996, n18997, n18998,
         n18999, n19000, n19001, n19002, n19003, n19004, n19005, n19006,
         n19007, n19008, n19009, n19010, n19011, n19012, n19013, n19014,
         n19015, n19016, n19017, n19018, n19019, n19020, n19021, n19022,
         n19023, n19024, n19025, n19026, n19027, n19028, n19029, n19030,
         n19031, n19032, n19033, n19034, n19035, n19036, n19037, n19038,
         n19039, n19040, n19041, n19042, n19043, n19044, n19045, n19046,
         n19047, n19048, n19049, n19050, n19051, n19052, n19053, n19054,
         n19055, n19056, n19057, n19058, n19059, n19060, n19061, n19062,
         n19063, n19064, n19065, n19066, n19067, n19068, n19069, n19070,
         n19071, n19072, n19073, n19074, n19075, n19076, n19077, n19078,
         n19079, n19080, n19081, n19082, n19083, n19084, n19085, n19086,
         n19087, n19088, n19089, n19090, n19091, n19092, n19093, n19094,
         n19095, n19096, n19097, n19098, n19099, n19100, n19101, n19102,
         n19103, n19104, n19105, n19106, n19107, n19108, n19109, n19110,
         n19111, n19112, n19113, n19114, n19115, n19116, n19117, n19118,
         n19119, n19120, n19121, n19122, n19123, n19124, n19125, n19126,
         n19127, n19128, n19129, n19130, n19131, n19132, n19133, n19134,
         n19135, n19136, n19137, n19138, n19139, n19140, n19141, n19142,
         n19143, n19144, n19145, n19146, n19147, n19148, n19149, n19150,
         n19151, n19152, n19153, n19154, n19155, n19156, n19157, n19158,
         n19159, n19160, n19161, n19162, n19163, n19164, n19165, n19166,
         n19167, n19168, n19169, n19170, n19171, n19172, n19173, n19174,
         n19175, n19176, n19177, n19178, n19179, n19180, n19181, n19182,
         n19183, n19184, n19185, n19186, n19187, n19188, n19189, n19190,
         n19191, n19192, n19193, n19194, n19195, n19196, n19197, n19198,
         n19199, n19200, n19201, n19202, n19203, n19204, n19205, n19206,
         n19207, n19208, n19209, n19210, n19211, n19212, n19213, n19214,
         n19215, n19216, n19217, n19218, n19219, n19220, n19221, n19222,
         n19223, n19224, n19225, n19226, n19227, n19228, n19229, n19230,
         n19231, n19232, n19233, n19234, n19235, n19236, n19237, n19238,
         n19239, n19240, n19241, n19242, n19243, n19244, n19245, n19246,
         n19247, n19248, n19249, n19250, n19251, n19252, n19253, n19254,
         n19255, n19256, n19257, n19258, n19259, n19260, n19261, n19262,
         n19263, n19264, n19265, n19266, n19267, n19268, n19269, n19270,
         n19271, n19272, n19273, n19274, n19275, n19276, n19277, n19278,
         n19279, n19280, n19281, n19282, n19283, n19284, n19285, n19286,
         n19287, n19288, n19289, n19290, n19291, n19292, n19293, n19294,
         n19295, n19296, n19297, n19298, n19299, n19300, n19301, n19302,
         n19303, n19304, n19305, n19306, n19307, n19308, n19309, n19310,
         n19311, n19312, n19313, n19314, n19315, n19316, n19317, n19318,
         n19319, n19320, n19321, n19322, n19323, n19324, n19325, n19326,
         n19327, n19328, n19329, n19330, n19331, n19332, n19333, n19334,
         n19335, n19336, n19337, n19338, n19339, n19340, n19341, n19342,
         n19343, n19344, n19345, n19346, n19347, n19348, n19349, n19350,
         n19351, n19352, n19353, n19354, n19355, n19356, n19357, n19358,
         n19359, n19360, n19361, n19362, n19363, n19364, n19365, n19366,
         n19367, n19368, n19369, n19370, n19371, n19372, n19373, n19374,
         n19375, n19376, n19377, n19378, n19379, n19380, n19381, n19382,
         n19383, n19384, n19385, n19386, n19387, n19388, n19389, n19390,
         n19391, n19392, n19393, n19394, n19395, n19396, n19397, n19398,
         n19399, n19400, n19401, n19402, n19403, n19404, n19405, n19406,
         n19407, n19408, n19409, n19410, n19411, n19412, n19413, n19414,
         n19415, n19416, n19417, n19418, n19419, n19420, n19421, n19422,
         n19423, n19424, n19425, n19426, n19427, n19428, n19429, n19430,
         n19431, n19432, n19433, n19434, n19435, n19436, n19437, n19438,
         n19439, n19440, n19441, n19442, n19443, n19444, n19445, n19446,
         n19447, n19448, n19449, n19450, n19451, n19452, n19453, n19454,
         n19455, n19456, n19457, n19458, n19459, n19460, n19461, n19462,
         n19463, n19464, n19465, n19466, n19467, n19468, n19469, n19470,
         n19471, n19472, n19473, n19474, n19475, n19476, n19477, n19478,
         n19479, n19480, n19481, n19482, n19483, n19484, n19485, n19486,
         n19487, n19488, n19489, n19490, n19491, n19492, n19493, n19494,
         n19495, n19496, n19497, n19498, n19499, n19500, n19501, n19502,
         n19503, n19504, n19505, n19506, n19507, n19508, n19509, n19510,
         n19511, n19512, n19513, n19514, n19515, n19516, n19517, n19518,
         n19519, n19520, n19521, n19522, n19523, n19524, n19525, n19526,
         n19527, n19528, n19529, n19530, n19531, n19532, n19533, n19534,
         n19535, n19536, n19537, n19538, n19539, n19540, n19541, n19542,
         n19543, n19544, n19545, n19546, n19547, n19548, n19549, n19550,
         n19551, n19552, n19553, n19554, n19555, n19556, n19557, n19558,
         n19559, n19560, n19561, n19562, n19563, n19564, n19565, n19566,
         n19567, n19568, n19569, n19570, n19571, n19572, n19573, n19574,
         n19575, n19576, n19577, n19578, n19579, n19580, n19581, n19582,
         n19583, n19584, n19585, n19586, n19587, n19588, n19589, n19590,
         n19591, n19592, n19593, n19594, n19595, n19596, n19597, n19598,
         n19599, n19600, n19601, n19602, n19603, n19604, n19605, n19606,
         n19607, n19608, n19609, n19610, n19611, n19612, n19613, n19614,
         n19615, n19616, n19617, n19618, n19619, n19620, n19621, n19622,
         n19623, n19624, n19625, n19626, n19627, n19628, n19629, n19630,
         n19631, n19632, n19633, n19634, n19635, n19636, n19637, n19638,
         n19639, n19640, n19641, n19642, n19643, n19644, n19645, n19646,
         n19647, n19648, n19649, n19650, n19651, n19652, n19653, n19654,
         n19655, n19656, n19657, n19658, n19659, n19660, n19661, n19662,
         n19663, n19664, n19665, n19666, n19667, n19668, n19669, n19670,
         n19671, n19672, n19673, n19674, n19675, n19676, n19677, n19678,
         n19679, n19680, n19681, n19682, n19683, n19684, n19685, n19686,
         n19687, n19688, n19689, n19690, n19691, n19692, n19693, n19694,
         n19695, n19696, n19697, n19698, n19699, n19700, n19701, n19702,
         n19703, n19704, n19705, n19706, n19707, n19708, n19709, n19710,
         n19711, n19712, n19713, n19714, n19715, n19716, n19717, n19718,
         n19719, n19720, n19721, n19722, n19723, n19724, n19725, n19726,
         n19727, n19728, n19729, n19730, n19731, n19732, n19733, n19734,
         n19735, n19736, n19737, n19738, n19739, n19740, n19741, n19742,
         n19743, n19744, n19745, n19746, n19747, n19748, n19749, n19750,
         n19751, n19752, n19753, n19754, n19755, n19756, n19757, n19758,
         n19759, n19760, n19761, n19762, n19763, n19764, n19765, n19766,
         n19767, n19768, n19769, n19770, n19771, n19772, n19773, n19774,
         n19775, n19776, n19777, n19778, n19779, n19780, n19781, n19782,
         n19783, n19784, n19785, n19786, n19787, n19788, n19789, n19790,
         n19791, n19792, n19793, n19794, n19795, n19796, n19797, n19798,
         n19799, n19800, n19801, n19802, n19803, n19804, n19805, n19806,
         n19807, n19808, n19809, n19810, n19811, n19812, n19813, n19814,
         n19815, n19816, n19817, n19818, n19819, n19820, n19821, n19822,
         n19823, n19824, n19825, n19826, n19827, n19828, n19829, n19830,
         n19831, n19832, n19833, n19834, n19835, n19836, n19837, n19838,
         n19839, n19840, n19841, n19842, n19843, n19844, n19845, n19846,
         n19847, n19848, n19849, n19850, n19851, n19852, n19853, n19854,
         n19855, n19856, n19857, n19858, n19859, n19860, n19861, n19862,
         n19863, n19864, n19865, n19866, n19867, n19868, n19869, n19870,
         n19871, n19872, n19873, n19874, n19875, n19876, n19877, n19878,
         n19879, n19880, n19881, n19882, n19883, n19884, n19885, n19886,
         n19887, n19888, n19889, n19890, n19891, n19892, n19893, n19894,
         n19895, n19896, n19897, n19898, n19899, n19900, n19901, n19902,
         n19903, n19904, n19905, n19906, n19907, n19908, n19909, n19910,
         n19911, n19912, n19913, n19914, n19915, n19916, n19917, n19918,
         n19919, n19920, n19921, n19922, n19923, n19924, n19925, n19926,
         n19927, n19928, n19929, n19930, n19931, n19932, n19933, n19934,
         n19935, n19936, n19937, n19938, n19939, n19940, n19941, n19942,
         n19943, n19944, n19945, n19946, n19947, n19948, n19949, n19950,
         n19951, n19952, n19953, n19954, n19955, n19956, n19957, n19958,
         n19959, n19960, n19961, n19962, n19963, n19964, n19965, n19966,
         n19967, n19968, n19969, n19970, n19971, n19972, n19973, n19974,
         n19975, n19976, n19977, n19978, n19979, n19980, n19981, n19982,
         n19983, n19984, n19985, n19986, n19987, n19988, n19989, n19990,
         n19991, n19992, n19993, n19994, n19995, n19996, n19997, n19998,
         n19999, n20000, n20001, n20002, n20003, n20004, n20005, n20006,
         n20007, n20008, n20009, n20010, n20011, n20012, n20013, n20014,
         n20015, n20016, n20017, n20018, n20019, n20020, n20021, n20022,
         n20023, n20024, n20025, n20026, n20027, n20028, n20029, n20030,
         n20031, n20032, n20033, n20034, n20035, n20036, n20037, n20038,
         n20039, n20040, n20041, n20042, n20043, n20044, n20045, n20046,
         n20047, n20048, n20049, n20050, n20051, n20052, n20053, n20054,
         n20055, n20056, n20057, n20058, n20059, n20060, n20061, n20062,
         n20063, n20064, n20065, n20066, n20067, n20068, n20069, n20070,
         n20071, n20072, n20073, n20074, n20075, n20076, n20077, n20078,
         n20079, n20080, n20081, n20082, n20083, n20084, n20085, n20086,
         n20087, n20088, n20089, n20090, n20091, n20092, n20093, n20094,
         n20095, n20096, n20097, n20098, n20099, n20100, n20101, n20102,
         n20103, n20104, n20105, n20106, n20107, n20108, n20109, n20110,
         n20111, n20112, n20113, n20114, n20115, n20116, n20117, n20118,
         n20119, n20120, n20121, n20122, n20123, n20124, n20125, n20126,
         n20127, n20128, n20129, n20130, n20131, n20132, n20133, n20134,
         n20135, n20136, n20137, n20138, n20139, n20140, n20141, n20142,
         n20143, n20144, n20145, n20146, n20147, n20148, n20149, n20150,
         n20151, n20152, n20153, n20154, n20155, n20156, n20157, n20158,
         n20159, n20160, n20161, n20162, n20163, n20164, n20165, n20166,
         n20167, n20168, n20169, n20170, n20171, n20172, n20173, n20174,
         n20175, n20176, n20177, n20178, n20179, n20180, n20181, n20182,
         n20183, n20184, n20185, n20186, n20187, n20188, n20189, n20190,
         n20191, n20192, n20193, n20194, n20195, n20196, n20197, n20198,
         n20199, n20200, n20201, n20202, n20203, n20204, n20205, n20206,
         n20207, n20208, n20209, n20210, n20211, n20212, n20213, n20214,
         n20215, n20216, n20217, n20218, n20219, n20220, n20221, n20222,
         n20223, n20224, n20225, n20226, n20227, n20228, n20229, n20230,
         n20231, n20232, n20233, n20234, n20235, n20236, n20237, n20238,
         n20239, n20240, n20241, n20242, n20243, n20244, n20245, n20246,
         n20247, n20248, n20249, n20250, n20251, n20252, n20253, n20254,
         n20255, n20256, n20257, n20258, n20259, n20260, n20261, n20262,
         n20263, n20264, n20265, n20266, n20267, n20268, n20269, n20270,
         n20271, n20272, n20273, n20274, n20275, n20276, n20277, n20278,
         n20279, n20280, n20281, n20282, n20283, n20284, n20285, n20286,
         n20287, n20288, n20289, n20290, n20291, n20292, n20293, n20294,
         n20295, n20296, n20297, n20298, n20299, n20300, n20301, n20302,
         n20303, n20304, n20305, n20306, n20307, n20308, n20309, n20310,
         n20311, n20312, n20313, n20314, n20315, n20316, n20317, n20318,
         n20319, n20320, n20321, n20322, n20323, n20324, n20325, n20326,
         n20327, n20328, n20329, n20330, n20331, n20332, n20333, n20334,
         n20335, n20336, n20337, n20338, n20339, n20340, n20341, n20342,
         n20343, n20344, n20345, n20346, n20347, n20348, n20349, n20350,
         n20351, n20352, n20353, n20354, n20355, n20356, n20357, n20358,
         n20359, n20360, n20361, n20362, n20363, n20364, n20365, n20366,
         n20367, n20368, n20369, n20370, n20371, n20372, n20373, n20374,
         n20375, n20376, n20377, n20378, n20379, n20380, n20381, n20382,
         n20383, n20384, n20385, n20386, n20387, n20388, n20389, n20390,
         n20391, n20392, n20393, n20394, n20395, n20396, n20397, n20398,
         n20399, n20400, n20401, n20402, n20403, n20404, n20405, n20406,
         n20407, n20408, n20409, n20410, n20411, n20412, n20413, n20414,
         n20415, n20416, n20417, n20418, n20419, n20420, n20421, n20422,
         n20423, n20424, n20425, n20426, n20427, n20428, n20429, n20430,
         n20431, n20432, n20433, n20434, n20435, n20436, n20437, n20438,
         n20439, n20440, n20441, n20442, n20443, n20444, n20445, n20446,
         n20447, n20448, n20449, n20450, n20451, n20452, n20453, n20454,
         n20455, n20456, n20457, n20458, n20459, n20460, n20461, n20462,
         n20463, n20464, n20465, n20466, n20467, n20468, n20469, n20470,
         n20471, n20472, n20473, n20474, n20475, n20476, n20477, n20478,
         n20479, n20480, n20481, n20482, n20483, n20484, n20485, n20486,
         n20487, n20488, n20489, n20490, n20491, n20492, n20493, n20494,
         n20495, n20496, n20497, n20498, n20499, n20500, n20501, n20502,
         n20503, n20504, n20505, n20506, n20507, n20508, n20509, n20510,
         n20511, n20512, n20513, n20514, n20515, n20516, n20517, n20518,
         n20519, n20520, n20521, n20522, n20523, n20524, n20525, n20526,
         n20527, n20528, n20529, n20530, n20531, n20532, n20533, n20534,
         n20535, n20536, n20537, n20538, n20539, n20540, n20541, n20542,
         n20543, n20544, n20545, n20546, n20547, n20548, n20549, n20550,
         n20551, n20552, n20553, n20554, n20555, n20556, n20557, n20558,
         n20559, n20560, n20561, n20562, n20563, n20564, n20565, n20566,
         n20567, n20568, n20569, n20570, n20571, n20572, n20573, n20574,
         n20575, n20576, n20577, n20578, n20579, n20580, n20581, n20582,
         n20583, n20584, n20585, n20586, n20587, n20588, n20589, n20590,
         n20591, n20592, n20593, n20594, n20595, n20596, n20597, n20598,
         n20599, n20600, n20601, n20602, n20603, n20604, n20605, n20606,
         n20607, n20608, n20609, n20610, n20611, n20612, n20613, n20614,
         n20615, n20616, n20617, n20618, n20619, n20620, n20621, n20622,
         n20623, n20624, n20625, n20626, n20627, n20628, n20629, n20630,
         n20631, n20632, n20633, n20634, n20635, n20636, n20637, n20638,
         n20639, n20640, n20641, n20642, n20643, n20644, n20645, n20646,
         n20647, n20648, n20649, n20650, n20651, n20652, n20653, n20654,
         n20655, n20656, n20657, n20658, n20659, n20660, n20661, n20662,
         n20663, n20664, n20665, n20666, n20667, n20668, n20669, n20670,
         n20671, n20672, n20673, n20674, n20675, n20676, n20677, n20678,
         n20679, n20680, n20681, n20682, n20683, n20684, n20685, n20686,
         n20687, n20688, n20689, n20690, n20691, n20692, n20693, n20694,
         n20695, n20696, n20697, n20698, n20699, n20700, n20701, n20702,
         n20703, n20704, n20705, n20706, n20707, n20708, n20709, n20710,
         n20711, n20712, n20713, n20714, n20715, n20716, n20717, n20718,
         n20719, n20720, n20721, n20722, n20723, n20724, n20725, n20726,
         n20727, n20728, n20729, n20730, n20731, n20732, n20733, n20734,
         n20735, n20736, n20737, n20738, n20739, n20740, n20741, n20742,
         n20743, n20744, n20745, n20746, n20747, n20748, n20749, n20750,
         n20751, n20752, n20753, n20754, n20755, n20756, n20757, n20758,
         n20759, n20760, n20761, n20762, n20763, n20764, n20765, n20766,
         n20767, n20768, n20769, n20770, n20771, n20772, n20773, n20774,
         n20775, n20776, n20777, n20778, n20779, n20780, n20781, n20782,
         n20783, n20784, n20785, n20786, n20787, n20788, n20789, n20790,
         n20791, n20792, n20793, n20794, n20795, n20796, n20797, n20798,
         n20799, n20800, n20801, n20802, n20803, n20804, n20805, n20806,
         n20807, n20808, n20809, n20810, n20811, n20812, n20813, n20814,
         n20815, n20816, n20817, n20818, n20819, n20820, n20821, n20822,
         n20823, n20824, n20825, n20826, n20827, n20828, n20829, n20830,
         n20831, n20832, n20833, n20834, n20835, n20836, n20837, n20838,
         n20839, n20840, n20841, n20842, n20843, n20844, n20845, n20846,
         n20847, n20848, n20849, n20850, n20851, n20852, n20853, n20854,
         n20855, n20856, n20857, n20858, n20859, n20860, n20861, n20862,
         n20863, n20864, n20865, n20866, n20867, n20868, n20869, n20870,
         n20871, n20872, n20873, n20874, n20875, n20876, n20877, n20878,
         n20879, n20880, n20881, n20882, n20883, n20884, n20885, n20886,
         n20887, n20888, n20889, n20890, n20891, n20892, n20893, n20894,
         n20895, n20896, n20897, n20898, n20899, n20900, n20901, n20902,
         n20903, n20904, n20905, n20906, n20907, n20908, n20909, n20910,
         n20911, n20912, n20913, n20914, n20915, n20916, n20917, n20918,
         n20919, n20920, n20921, n20922, n20923, n20924, n20925, n20926,
         n20927, n20928, n20929, n20930, n20931, n20932, n20933, n20934,
         n20935, n20936, n20937, n20938, n20939, n20940, n20941, n20942,
         n20943, n20944, n20945, n20946, n20947, n20948, n20949, n20950,
         n20951, n20952, n20953, n20954, n20955, n20956, n20957, n20958,
         n20959, n20960, n20961, n20962, n20963, n20964, n20965, n20966,
         n20967, n20968, n20969, n20970, n20971, n20972, n20973, n20974,
         n20975, n20976, n20977, n20978, n20979, n20980, n20981, n20982,
         n20983, n20984, n20985, n20986, n20987, n20988, n20989, n20990,
         n20991, n20992, n20993, n20994, n20995, n20996, n20997, n20998,
         n20999, n21000, n21001, n21002, n21003, n21004, n21005, n21006,
         n21007, n21008, n21009, n21010, n21011, n21012, n21013, n21014,
         n21015, n21016, n21017, n21018, n21019, n21020, n21021, n21022,
         n21023, n21024, n21025, n21026, n21027, n21028, n21029, n21030,
         n21031, n21032, n21033, n21034, n21035, n21036, n21037, n21038,
         n21039, n21040, n21041, n21042, n21043, n21044, n21045, n21046,
         n21047, n21048, n21049, n21050, n21051, n21052, n21053, n21054,
         n21055, n21056, n21057, n21058, n21059, n21060, n21061, n21062,
         n21063, n21064, n21065, n21066, n21067, n21068, n21069, n21070,
         n21071, n21072, n21073, n21074, n21075, n21076, n21077, n21078,
         n21079, n21080, n21081, n21082, n21083, n21084, n21085, n21086,
         n21087, n21088, n21089, n21090, n21091, n21092, n21093, n21094,
         n21095, n21096, n21097, n21098, n21099, n21100, n21101, n21102,
         n21103, n21104, n21105, n21106, n21107, n21108, n21109, n21110,
         n21111, n21112, n21113, n21114, n21115, n21116, n21117, n21118,
         n21119, n21120, n21121, n21122, n21123, n21124, n21125, n21126,
         n21127, n21128, n21129, n21130, n21131, n21132, n21133, n21134,
         n21135, n21136, n21137, n21138, n21139, n21140, n21141, n21142,
         n21143, n21144, n21145, n21146, n21147, n21148, n21149, n21150,
         n21151, n21152, n21153, n21154, n21155, n21156, n21157, n21158,
         n21159, n21160, n21161, n21162, n21163, n21164, n21165, n21166,
         n21167, n21168, n21169, n21170, n21171, n21172, n21173, n21174,
         n21175, n21176, n21177, n21178, n21179, n21180, n21181, n21182,
         n21183, n21184, n21185, n21186, n21187, n21188, n21189, n21190,
         n21191, n21192, n21193, n21194, n21195, n21196, n21197, n21198,
         n21199, n21200, n21201, n21202, n21203, n21204, n21205, n21206,
         n21207, n21208, n21209, n21210, n21211, n21212, n21213, n21214,
         n21215, n21216, n21217, n21218, n21219, n21220, n21221, n21222,
         n21223, n21224, n21225, n21226, n21227, n21228, n21229, n21230,
         n21231, n21232, n21233, n21234, n21235, n21236, n21237, n21238,
         n21239, n21240, n21241, n21242, n21243, n21244, n21245, n21246,
         n21247, n21248, n21249, n21250, n21251, n21252, n21253, n21254,
         n21255, n21256, n21257, n21258, n21259, n21260, n21261, n21262,
         n21263, n21264, n21265, n21266, n21267, n21268, n21269, n21270,
         n21271, n21272, n21273, n21274, n21275, n21276, n21277, n21278,
         n21279, n21280, n21281, n21282, n21283, n21284, n21285, n21286,
         n21287, n21288, n21289, n21290, n21291, n21292, n21293, n21294,
         n21295, n21296, n21297, n21298, n21299, n21300, n21301, n21302,
         n21303, n21304, n21305, n21306, n21307, n21308, n21309, n21310,
         n21311, n21312, n21313, n21314, n21315, n21316, n21317, n21318,
         n21319, n21320, n21321, n21322, n21323, n21324, n21325, n21326,
         n21327, n21328, n21329, n21330, n21331, n21332, n21333, n21334,
         n21335, n21336, n21337, n21338, n21339, n21340, n21341, n21342,
         n21343, n21344, n21345, n21346, n21347, n21348, n21349, n21350,
         n21351, n21352, n21353, n21354, n21355, n21356, n21357, n21358,
         n21359, n21360, n21361, n21362, n21363, n21364, n21365, n21366,
         n21367, n21368, n21369, n21370, n21371, n21372, n21373, n21374,
         n21375, n21376, n21377, n21378, n21379, n21380, n21381, n21382,
         n21383, n21384, n21385, n21386, n21387, n21388, n21389, n21390,
         n21391, n21392, n21393, n21394, n21395, n21396, n21397, n21398,
         n21399, n21400, n21401;

  NAND2_X1 U11260 ( .A1(n18195), .A2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n18194) );
  INV_X1 U11261 ( .A(n18050), .ZN(n18039) );
  AND2_X1 U11262 ( .A1(n10130), .A2(n10135), .ZN(n15519) );
  NOR2_X2 U11263 ( .A1(n9996), .A2(n18864), .ZN(n17432) );
  INV_X1 U11264 ( .A(n19159), .ZN(n10135) );
  CLKBUF_X2 U11265 ( .A(n11907), .Z(n9844) );
  AND4_X1 U11267 ( .A1(n11221), .A2(n11220), .A3(n11219), .A4(n11218), .ZN(
        n11228) );
  AND2_X2 U11268 ( .A1(n11177), .A2(n19354), .ZN(n11222) );
  CLKBUF_X2 U11269 ( .A(n12651), .Z(n17327) );
  NAND2_X1 U11270 ( .A1(n11144), .A2(n11145), .ZN(n11168) );
  INV_X1 U11271 ( .A(n14610), .ZN(n10663) );
  AND2_X1 U11272 ( .A1(n14624), .A2(n10435), .ZN(n14598) );
  AND2_X1 U11273 ( .A1(n9823), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10667) );
  INV_X1 U11274 ( .A(n10549), .ZN(n14579) );
  INV_X1 U11275 ( .A(n10351), .ZN(n14618) );
  NAND2_X1 U11276 ( .A1(n14770), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n14603) );
  CLKBUF_X1 U11277 ( .A(n11622), .Z(n12356) );
  INV_X2 U11278 ( .A(n16201), .ZN(n11633) );
  CLKBUF_X2 U11279 ( .A(n11599), .Z(n9850) );
  MUX2_X1 U11280 ( .A(n10625), .B(n10624), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n19391) );
  INV_X1 U11281 ( .A(n11816), .ZN(n11641) );
  NAND2_X1 U11282 ( .A1(n10209), .A2(n10607), .ZN(n10208) );
  AND2_X2 U11283 ( .A1(n10435), .A2(n9840), .ZN(n10644) );
  AND2_X2 U11284 ( .A1(n11527), .A2(n13946), .ZN(n11612) );
  AND2_X1 U11285 ( .A1(n11536), .A2(n13945), .ZN(n11766) );
  NOR2_X2 U11286 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10425) );
  INV_X1 U11287 ( .A(n12730), .ZN(n9816) );
  INV_X2 U11288 ( .A(n9816), .ZN(n9817) );
  INV_X1 U11289 ( .A(n14601), .ZN(n10664) );
  AND2_X2 U11290 ( .A1(n11527), .A2(n10328), .ZN(n11599) );
  BUF_X1 U11291 ( .A(n9825), .Z(n9852) );
  CLKBUF_X3 U11292 ( .A(n10648), .Z(n14770) );
  INV_X1 U11293 ( .A(n10352), .ZN(n14599) );
  NOR2_X1 U11294 ( .A1(n10077), .A2(n10076), .ZN(n10994) );
  AND2_X1 U11295 ( .A1(n11162), .A2(n14805), .ZN(n19715) );
  INV_X2 U11296 ( .A(n17344), .ZN(n17363) );
  OR2_X1 U11298 ( .A1(n11583), .A2(n11582), .ZN(n11640) );
  OR2_X1 U11299 ( .A1(n14250), .A2(n14403), .ZN(n14432) );
  AND2_X1 U11300 ( .A1(n11160), .A2(n14805), .ZN(n19672) );
  INV_X2 U11301 ( .A(n12537), .ZN(n17245) );
  OR2_X2 U11302 ( .A1(n11549), .A2(n11548), .ZN(n11979) );
  XNOR2_X1 U11303 ( .A(n11843), .B(n14501), .ZN(n13733) );
  XNOR2_X1 U11305 ( .A(n13471), .B(n20460), .ZN(n20597) );
  NOR2_X1 U11306 ( .A1(n15519), .A2(n15786), .ZN(n15518) );
  NAND2_X1 U11307 ( .A1(n11299), .A2(n10960), .ZN(n12460) );
  NOR2_X1 U11308 ( .A1(n16631), .A2(n16610), .ZN(n16609) );
  OR4_X1 U11309 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A4(n12516), .ZN(n13050) );
  INV_X1 U11310 ( .A(n20122), .ZN(n20147) );
  NAND2_X1 U11311 ( .A1(n14853), .A2(n14854), .ZN(n14833) );
  CLKBUF_X3 U11312 ( .A(n13002), .Z(n15174) );
  NAND2_X1 U11313 ( .A1(n13354), .A2(n13353), .ZN(n16107) );
  INV_X1 U11314 ( .A(n9919), .ZN(n17386) );
  INV_X1 U11315 ( .A(n18413), .ZN(n17547) );
  NAND2_X1 U11316 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n18189), .ZN(
        n18188) );
  INV_X1 U11317 ( .A(n18031), .ZN(n17763) );
  NAND2_X1 U11318 ( .A1(n18222), .A2(n18821), .ZN(n18276) );
  INV_X2 U11319 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n12516) );
  AND2_X1 U11320 ( .A1(n12515), .A2(n18972), .ZN(n9818) );
  BUF_X1 U11321 ( .A(n10971), .Z(n9839) );
  NAND2_X4 U11322 ( .A1(n9855), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n14601) );
  AND2_X2 U11323 ( .A1(n15263), .A2(n11901), .ZN(n9837) );
  NOR2_X4 U11324 ( .A1(n11466), .A2(n15566), .ZN(n15553) );
  INV_X2 U11325 ( .A(n13214), .ZN(n17581) );
  NAND3_X2 U11326 ( .A1(n13096), .A2(n13095), .A3(n13094), .ZN(n13214) );
  AND2_X2 U11327 ( .A1(n11168), .A2(n11148), .ZN(n14093) );
  INV_X2 U11328 ( .A(n11644), .ZN(n13775) );
  AND2_X1 U11329 ( .A1(n13958), .A2(n11528), .ZN(n9819) );
  AND2_X1 U11330 ( .A1(n13958), .A2(n11528), .ZN(n9820) );
  AND2_X2 U11331 ( .A1(n13958), .A2(n11528), .ZN(n12392) );
  AND4_X2 U11332 ( .A1(n11553), .A2(n11552), .A3(n11551), .A4(n11550), .ZN(
        n11561) );
  NAND2_X4 U11333 ( .A1(n10210), .A2(n10208), .ZN(n19420) );
  XNOR2_X2 U11334 ( .A(n11871), .B(n16430), .ZN(n16341) );
  NAND2_X1 U11335 ( .A1(n13734), .A2(n13733), .ZN(n13735) );
  AND2_X1 U11336 ( .A1(n13958), .A2(n13946), .ZN(n9821) );
  AND2_X1 U11337 ( .A1(n13958), .A2(n13946), .ZN(n12723) );
  INV_X1 U11338 ( .A(n17379), .ZN(n17360) );
  NOR2_X2 U11339 ( .A1(n10399), .A2(n16506), .ZN(n10400) );
  AND2_X1 U11340 ( .A1(n10435), .A2(n9840), .ZN(n9822) );
  AND2_X2 U11341 ( .A1(n10435), .A2(n9840), .ZN(n9823) );
  OR2_X4 U11342 ( .A1(n11632), .A2(n11631), .ZN(n16201) );
  AND2_X2 U11343 ( .A1(n10647), .A2(n10607), .ZN(n10485) );
  CLKBUF_X1 U11344 ( .A(n11573), .Z(n9824) );
  BUF_X4 U11345 ( .A(n11573), .Z(n9825) );
  BUF_X4 U11346 ( .A(n11573), .Z(n9826) );
  INV_X2 U11347 ( .A(n9818), .ZN(n9827) );
  AND2_X4 U11348 ( .A1(n13946), .A2(n15472), .ZN(n11716) );
  AND2_X4 U11349 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n15472) );
  NOR2_X2 U11350 ( .A1(n11559), .A2(n11558), .ZN(n11560) );
  CLKBUF_X1 U11351 ( .A(n15180), .Z(n15181) );
  NOR2_X1 U11352 ( .A1(n14727), .A2(n14726), .ZN(n14730) );
  AND2_X1 U11353 ( .A1(n14727), .A2(n14726), .ZN(n14728) );
  NAND2_X1 U11354 ( .A1(n15263), .A2(n11901), .ZN(n15219) );
  NOR3_X1 U11355 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17957), .A3(
        n17709), .ZN(n16164) );
  NOR2_X1 U11356 ( .A1(n17697), .A2(n17696), .ZN(n17695) );
  INV_X2 U11357 ( .A(n9845), .ZN(n16302) );
  NAND2_X1 U11358 ( .A1(n11885), .A2(n11818), .ZN(n11907) );
  NAND2_X1 U11359 ( .A1(n18215), .A2(n18228), .ZN(n18221) );
  NAND2_X1 U11360 ( .A1(n13161), .A2(n17795), .ZN(n17829) );
  AND2_X1 U11361 ( .A1(n13662), .A2(n10148), .ZN(n13811) );
  AND2_X1 U11362 ( .A1(n11158), .A2(n14805), .ZN(n19433) );
  AND2_X1 U11363 ( .A1(n9979), .A2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n13224) );
  AND2_X1 U11364 ( .A1(n11169), .A2(n19342), .ZN(n11178) );
  AND2_X1 U11365 ( .A1(n11161), .A2(n14805), .ZN(n11208) );
  AND2_X1 U11366 ( .A1(n11158), .A2(n19342), .ZN(n11207) );
  OR2_X1 U11367 ( .A1(n17976), .A2(n17977), .ZN(n9979) );
  AOI21_X1 U11368 ( .B1(n17969), .B2(n13150), .A(n18283), .ZN(n17896) );
  NAND2_X2 U11369 ( .A1(n17432), .A2(n18413), .ZN(n17571) );
  CLKBUF_X2 U11370 ( .A(n13564), .Z(n19342) );
  CLKBUF_X2 U11371 ( .A(n13415), .Z(n9860) );
  NAND2_X1 U11372 ( .A1(n14302), .A2(n14304), .ZN(n19424) );
  NAND2_X1 U11373 ( .A1(n11019), .A2(n11018), .ZN(n11141) );
  AND2_X1 U11374 ( .A1(n11318), .A2(n9938), .ZN(n11338) );
  AOI21_X1 U11375 ( .B1(n13174), .B2(n13175), .A(n13185), .ZN(n13290) );
  NAND3_X1 U11376 ( .A1(n13176), .A2(n13172), .A3(n18378), .ZN(n16732) );
  NOR2_X2 U11377 ( .A1(n11277), .A2(n11276), .ZN(n11301) );
  AOI22_X1 U11378 ( .A1(n14090), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(n14129), 
        .B2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n10964) );
  AND2_X1 U11379 ( .A1(n11258), .A2(n11264), .ZN(n11271) );
  CLKBUF_X3 U11380 ( .A(n11021), .Z(n12812) );
  NOR2_X1 U11381 ( .A1(n18393), .A2(n12617), .ZN(n13198) );
  AND2_X1 U11382 ( .A1(n11597), .A2(n11596), .ZN(n11649) );
  NAND2_X1 U11383 ( .A1(n12579), .A2(n9902), .ZN(n18405) );
  NAND2_X1 U11384 ( .A1(n18413), .A2(n16232), .ZN(n13173) );
  INV_X1 U11385 ( .A(n12755), .ZN(n21001) );
  AOI211_X1 U11386 ( .C1(n17378), .C2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A(
        n13048), .B(n13047), .ZN(n17557) );
  NAND2_X1 U11387 ( .A1(n11633), .A2(n11644), .ZN(n12755) );
  AND2_X1 U11389 ( .A1(n11636), .A2(n11979), .ZN(n11650) );
  CLKBUF_X2 U11390 ( .A(n10689), .Z(n12819) );
  INV_X4 U11391 ( .A(n10960), .ZN(n10543) );
  INV_X1 U11392 ( .A(n10959), .ZN(n10971) );
  NAND2_X1 U11393 ( .A1(n20331), .A2(n16201), .ZN(n12848) );
  NAND2_X1 U11394 ( .A1(n10075), .A2(n10456), .ZN(n10959) );
  OAI21_X1 U11395 ( .B1(n10455), .B2(n10454), .A(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10075) );
  INV_X2 U11396 ( .A(n14603), .ZN(n10672) );
  INV_X4 U11397 ( .A(n17395), .ZN(n13080) );
  INV_X4 U11398 ( .A(n9827), .ZN(n13089) );
  BUF_X2 U11399 ( .A(n11692), .Z(n12732) );
  CLKBUF_X2 U11400 ( .A(n11697), .Z(n12729) );
  BUF_X2 U11401 ( .A(n11684), .Z(n12286) );
  CLKBUF_X2 U11402 ( .A(n11715), .Z(n12731) );
  CLKBUF_X2 U11403 ( .A(n11766), .Z(n12250) );
  INV_X1 U11404 ( .A(n14609), .ZN(n10666) );
  INV_X2 U11405 ( .A(n13079), .ZN(n12551) );
  BUF_X2 U11406 ( .A(n10649), .Z(n9855) );
  INV_X4 U11407 ( .A(n17283), .ZN(n12552) );
  NAND2_X1 U11408 ( .A1(n10646), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n14609) );
  NOR2_X1 U11409 ( .A1(n12507), .A2(n12516), .ZN(n12515) );
  INV_X4 U11410 ( .A(n17306), .ZN(n17365) );
  INV_X4 U11411 ( .A(n13050), .ZN(n17361) );
  NOR2_X4 U11412 ( .A1(n12508), .A2(n18840), .ZN(n17379) );
  INV_X4 U11413 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n18982) );
  NOR2_X4 U11414 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10328) );
  NOR2_X4 U11415 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13958) );
  NOR2_X1 U11417 ( .A1(n12831), .A2(n12830), .ZN(n12832) );
  OR2_X1 U11418 ( .A1(n12997), .A2(n16553), .ZN(n12981) );
  OR2_X1 U11419 ( .A1(n12997), .A2(n19363), .ZN(n12998) );
  NOR2_X1 U11420 ( .A1(n15154), .A2(n15348), .ZN(n9986) );
  NAND2_X1 U11421 ( .A1(n14821), .A2(n12410), .ZN(n14516) );
  INV_X1 U11422 ( .A(n13001), .ZN(n11911) );
  XNOR2_X1 U11423 ( .A(n12751), .B(n12750), .ZN(n13010) );
  NOR2_X1 U11424 ( .A1(n14730), .A2(n14728), .ZN(n15637) );
  OR2_X1 U11425 ( .A1(n14833), .A2(n10346), .ZN(n12751) );
  NOR2_X1 U11426 ( .A1(n14531), .A2(n16072), .ZN(n15859) );
  AND2_X1 U11427 ( .A1(n11130), .A2(n11129), .ZN(n11131) );
  NOR2_X2 U11428 ( .A1(n14858), .A2(n14860), .ZN(n14853) );
  XNOR2_X1 U11429 ( .A(n14706), .B(n14703), .ZN(n15647) );
  AND2_X1 U11430 ( .A1(n11906), .A2(n9989), .ZN(n9988) );
  AOI21_X1 U11431 ( .B1(n15873), .B2(n19341), .A(n15872), .ZN(n15876) );
  XNOR2_X1 U11432 ( .A(n12817), .B(n12816), .ZN(n15624) );
  NAND2_X1 U11433 ( .A1(n15650), .A2(n10378), .ZN(n14706) );
  NAND2_X1 U11434 ( .A1(n14469), .A2(n11899), .ZN(n10300) );
  AND2_X1 U11435 ( .A1(n9914), .A2(n11456), .ZN(n10081) );
  NAND2_X1 U11436 ( .A1(n9981), .A2(n16330), .ZN(n14469) );
  OR2_X1 U11437 ( .A1(n13316), .A2(n13319), .ZN(n15889) );
  OR2_X1 U11438 ( .A1(n15222), .A2(n15220), .ZN(n10049) );
  AND2_X1 U11439 ( .A1(n16301), .A2(n10294), .ZN(n10293) );
  OR2_X1 U11440 ( .A1(n15644), .A2(n13317), .ZN(n16452) );
  NOR2_X1 U11441 ( .A1(n10089), .A2(n10086), .ZN(n10085) );
  OR2_X1 U11442 ( .A1(n16538), .A2(n11476), .ZN(n10086) );
  AND2_X1 U11443 ( .A1(n15224), .A2(n15221), .ZN(n16301) );
  OR2_X1 U11444 ( .A1(n14470), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11899) );
  NOR2_X1 U11445 ( .A1(n10306), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n10089) );
  NAND2_X1 U11446 ( .A1(n15235), .A2(n11902), .ZN(n15248) );
  AND2_X1 U11447 ( .A1(n16312), .A2(n16311), .ZN(n15224) );
  NOR2_X1 U11448 ( .A1(n14020), .A2(n10332), .ZN(n10331) );
  AND2_X1 U11449 ( .A1(n9844), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n13006) );
  INV_X1 U11450 ( .A(n14290), .ZN(n10333) );
  OR2_X1 U11451 ( .A1(n11459), .A2(n11458), .ZN(n11461) );
  NAND2_X1 U11452 ( .A1(n13850), .A2(n13849), .ZN(n13848) );
  AOI21_X1 U11453 ( .B1(n12037), .B2(n12154), .A(n12036), .ZN(n14290) );
  NAND2_X1 U11454 ( .A1(n10330), .A2(n10329), .ZN(n10332) );
  AND2_X1 U11455 ( .A1(n15510), .A2(n12490), .ZN(n12492) );
  NOR2_X1 U11456 ( .A1(n18194), .A2(n17729), .ZN(n17734) );
  NAND2_X1 U11457 ( .A1(n11815), .A2(n11814), .ZN(n11885) );
  NOR2_X1 U11458 ( .A1(n9886), .A2(n15509), .ZN(n15510) );
  AND2_X1 U11459 ( .A1(n11252), .A2(n11251), .ZN(n11450) );
  NAND4_X1 U11460 ( .A1(n11182), .A2(n11181), .A3(n11180), .A4(n11179), .ZN(
        n11185) );
  INV_X2 U11461 ( .A(n16293), .ZN(n15090) );
  AND2_X1 U11462 ( .A1(n11190), .A2(n11189), .ZN(n11191) );
  NOR2_X1 U11463 ( .A1(n13826), .A2(n13997), .ZN(n11061) );
  NAND2_X1 U11464 ( .A1(n18045), .A2(n18006), .ZN(n18041) );
  INV_X2 U11465 ( .A(n20178), .ZN(n9828) );
  NAND2_X1 U11466 ( .A1(n11990), .A2(n11989), .ZN(n13542) );
  NAND2_X1 U11467 ( .A1(n13592), .A2(n13593), .ZN(n13624) );
  OAI21_X2 U11468 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n19019), .A(n16733), 
        .ZN(n18045) );
  AND2_X1 U11469 ( .A1(n11161), .A2(n19342), .ZN(n19605) );
  CLKBUF_X1 U11470 ( .A(n13973), .Z(n9853) );
  NAND2_X1 U11471 ( .A1(n19012), .A2(n13232), .ZN(n18050) );
  AND2_X1 U11472 ( .A1(n10135), .A2(n10133), .ZN(n15550) );
  AOI21_X2 U11473 ( .B1(n13574), .B2(n13573), .A(n13572), .ZN(n13619) );
  NAND2_X1 U11474 ( .A1(n10147), .A2(n9907), .ZN(n13660) );
  NAND2_X1 U11475 ( .A1(n11778), .A2(n11777), .ZN(n13972) );
  NAND2_X1 U11476 ( .A1(n17969), .A2(n9905), .ZN(n13199) );
  INV_X1 U11477 ( .A(n11820), .ZN(n9983) );
  NAND2_X1 U11478 ( .A1(n17970), .A2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n17969) );
  NOR2_X1 U11479 ( .A1(n14171), .A2(n14172), .ZN(n16075) );
  NAND2_X1 U11480 ( .A1(n13744), .A2(n13223), .ZN(n17976) );
  AND2_X1 U11481 ( .A1(n17375), .A2(n9882), .ZN(n13981) );
  XNOR2_X1 U11482 ( .A(n16107), .B(n13570), .ZN(n13573) );
  NAND2_X1 U11483 ( .A1(n10264), .A2(n9903), .ZN(n10263) );
  INV_X1 U11484 ( .A(n9860), .ZN(n19354) );
  AOI21_X1 U11485 ( .B1(n13415), .B2(n13587), .A(n13414), .ZN(n13574) );
  AND2_X1 U11486 ( .A1(n9896), .A2(n13668), .ZN(n9907) );
  NAND2_X1 U11487 ( .A1(n9993), .A2(n11691), .ZN(n11831) );
  AND2_X1 U11488 ( .A1(n10150), .A2(n10149), .ZN(n10148) );
  NAND2_X1 U11489 ( .A1(n11747), .A2(n11746), .ZN(n13471) );
  AND2_X1 U11490 ( .A1(n10151), .A2(n13707), .ZN(n10150) );
  NAND2_X1 U11491 ( .A1(n11741), .A2(n11740), .ZN(n11747) );
  CLKBUF_X3 U11492 ( .A(n10415), .Z(n19159) );
  NAND2_X1 U11493 ( .A1(n11678), .A2(n20423), .ZN(n11741) );
  NAND2_X1 U11494 ( .A1(n11014), .A2(n11015), .ZN(n11019) );
  NOR2_X1 U11495 ( .A1(n13723), .A2(n10152), .ZN(n10151) );
  CLKBUF_X1 U11496 ( .A(n11993), .Z(n20422) );
  NAND2_X1 U11497 ( .A1(n9970), .A2(n9969), .ZN(n13743) );
  XNOR2_X1 U11498 ( .A(n11662), .B(n11735), .ZN(n20423) );
  NAND2_X1 U11499 ( .A1(n13290), .A2(n13289), .ZN(n18824) );
  AND2_X1 U11500 ( .A1(n11038), .A2(n11037), .ZN(n13661) );
  AND2_X1 U11501 ( .A1(n11044), .A2(n11043), .ZN(n13723) );
  OAI211_X1 U11502 ( .C1(n20318), .C2(n11745), .A(n11744), .B(n11743), .ZN(
        n11746) );
  NAND2_X1 U11503 ( .A1(n10965), .A2(n10964), .ZN(n10993) );
  NAND2_X1 U11504 ( .A1(n16231), .A2(n10128), .ZN(n17425) );
  INV_X1 U11505 ( .A(n11053), .ZN(n12815) );
  NAND3_X1 U11506 ( .A1(n10215), .A2(n10988), .A3(n10214), .ZN(n11013) );
  NAND2_X1 U11507 ( .A1(n9968), .A2(n13139), .ZN(n13140) );
  NAND2_X1 U11508 ( .A1(n10079), .A2(n10078), .ZN(n10077) );
  AND3_X1 U11509 ( .A1(n10990), .A2(n10989), .A3(n10361), .ZN(n10991) );
  NAND2_X1 U11510 ( .A1(n10043), .A2(n10042), .ZN(n10363) );
  NOR2_X1 U11511 ( .A1(n17557), .A2(n13143), .ZN(n13144) );
  AND3_X1 U11512 ( .A1(n10973), .A2(n14073), .A3(n10972), .ZN(n10974) );
  AND2_X1 U11513 ( .A1(n13367), .A2(n13368), .ZN(n13366) );
  AND2_X1 U11514 ( .A1(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n10383), .ZN(
        n10396) );
  INV_X1 U11515 ( .A(n12757), .ZN(n11634) );
  INV_X1 U11516 ( .A(n14388), .ZN(n10329) );
  NOR2_X1 U11517 ( .A1(n11266), .A2(n11265), .ZN(n11264) );
  CLKBUF_X1 U11518 ( .A(n12849), .Z(n13630) );
  OR2_X1 U11519 ( .A1(n11470), .A2(n11384), .ZN(n10988) );
  NAND2_X1 U11520 ( .A1(n10975), .A2(n10941), .ZN(n10983) );
  AND2_X1 U11521 ( .A1(n10362), .A2(n13380), .ZN(n11469) );
  AND2_X1 U11522 ( .A1(n16156), .A2(n11481), .ZN(n11492) );
  AND2_X1 U11523 ( .A1(n10976), .A2(n14723), .ZN(n11022) );
  NOR2_X1 U11524 ( .A1(n18405), .A2(n17433), .ZN(n12617) );
  AND3_X1 U11525 ( .A1(n9995), .A2(n11639), .A3(n9994), .ZN(n11597) );
  AND2_X1 U11526 ( .A1(n16196), .A2(n12848), .ZN(n13420) );
  NOR2_X2 U11527 ( .A1(n11640), .A2(n20331), .ZN(n13943) );
  NAND2_X1 U11528 ( .A1(n11654), .A2(n11585), .ZN(n11657) );
  AND2_X1 U11529 ( .A1(n11408), .A2(n10657), .ZN(n10976) );
  OR2_X1 U11530 ( .A1(n13078), .A2(n13077), .ZN(n17568) );
  OAI211_X2 U11531 ( .C1(n12561), .C2(n21152), .A(n12524), .B(n12523), .ZN(
        n18413) );
  AND3_X2 U11532 ( .A1(n10679), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n20062), 
        .ZN(n14723) );
  INV_X1 U11533 ( .A(n11640), .ZN(n13762) );
  AND3_X1 U11534 ( .A1(n13133), .A2(n13132), .A3(n13131), .ZN(n10364) );
  NAND2_X1 U11535 ( .A1(n10679), .A2(n10680), .ZN(n10968) );
  AND2_X1 U11536 ( .A1(n13063), .A2(n10360), .ZN(n17564) );
  OAI211_X1 U11537 ( .C1(n13050), .C2(n21306), .A(n12591), .B(n12590), .ZN(
        n18393) );
  AND2_X1 U11538 ( .A1(n13351), .A2(n19420), .ZN(n13389) );
  INV_X1 U11539 ( .A(n19384), .ZN(n11487) );
  NAND2_X1 U11540 ( .A1(n10959), .A2(n10657), .ZN(n11379) );
  CLKBUF_X1 U11541 ( .A(n11635), .Z(n11679) );
  OR2_X1 U11542 ( .A1(n10490), .A2(n10489), .ZN(n10707) );
  CLKBUF_X3 U11543 ( .A(n10959), .Z(n20062) );
  AND2_X1 U11544 ( .A1(n10935), .A2(n10679), .ZN(n10966) );
  OR2_X2 U11545 ( .A1(n11595), .A2(n11594), .ZN(n20331) );
  NAND2_X1 U11546 ( .A1(n10615), .A2(n10614), .ZN(n19384) );
  NAND2_X2 U11547 ( .A1(n10273), .A2(n10272), .ZN(n10657) );
  CLKBUF_X1 U11548 ( .A(n11651), .Z(n11652) );
  AND4_X1 U11549 ( .A1(n11616), .A2(n11615), .A3(n11614), .A4(n11613), .ZN(
        n11617) );
  NAND3_X1 U11550 ( .A1(n11539), .A2(n10382), .A3(n11538), .ZN(n11651) );
  NAND2_X2 U11551 ( .A1(n11571), .A2(n11570), .ZN(n11816) );
  AND4_X1 U11552 ( .A1(n11611), .A2(n11610), .A3(n11609), .A4(n11608), .ZN(
        n11618) );
  AND4_X1 U11553 ( .A1(n11607), .A2(n11606), .A3(n11605), .A4(n11604), .ZN(
        n11619) );
  CLKBUF_X3 U11554 ( .A(n11599), .Z(n9851) );
  AND4_X1 U11555 ( .A1(n11534), .A2(n11533), .A3(n11532), .A4(n11531), .ZN(
        n10382) );
  AND4_X1 U11556 ( .A1(n10606), .A2(n10605), .A3(n10604), .A4(n10603), .ZN(
        n10608) );
  AND4_X1 U11557 ( .A1(n11569), .A2(n11568), .A3(n11567), .A4(n11566), .ZN(
        n11570) );
  OR2_X2 U11558 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n13326), .ZN(n19345) );
  AND4_X1 U11559 ( .A1(n11565), .A2(n11564), .A3(n11563), .A4(n11562), .ZN(
        n11571) );
  NAND2_X2 U11560 ( .A1(n18720), .A2(n16145), .ZN(n18418) );
  AND3_X1 U11561 ( .A1(n11525), .A2(n11524), .A3(n11523), .ZN(n11539) );
  AOI22_X1 U11562 ( .A1(n11766), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12722), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11554) );
  NAND2_X2 U11563 ( .A1(n18960), .A2(n18897), .ZN(n18946) );
  BUF_X4 U11564 ( .A(n12043), .Z(n9838) );
  AND3_X1 U11565 ( .A1(n10598), .A2(n10597), .A3(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10599) );
  AND2_X1 U11566 ( .A1(n10593), .A2(n10607), .ZN(n10594) );
  INV_X2 U11567 ( .A(n12561), .ZN(n9829) );
  AND2_X1 U11568 ( .A1(n10633), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10634) );
  AND3_X1 U11569 ( .A1(n10630), .A2(n10629), .A3(n10628), .ZN(n10631) );
  INV_X2 U11570 ( .A(n9919), .ZN(n17357) );
  INV_X2 U11571 ( .A(n12651), .ZN(n17384) );
  INV_X2 U11572 ( .A(n16722), .ZN(n16724) );
  BUF_X2 U11573 ( .A(n10462), .Z(n9857) );
  CLKBUF_X3 U11574 ( .A(n10462), .Z(n9859) );
  AND3_X1 U11575 ( .A1(n10407), .A2(n10138), .A3(n10136), .ZN(n10409) );
  OR2_X1 U11576 ( .A1(n12514), .A2(n9980), .ZN(n12537) );
  BUF_X2 U11577 ( .A(n10462), .Z(n9858) );
  OR2_X1 U11578 ( .A1(n12513), .A2(n12514), .ZN(n9884) );
  AND2_X2 U11579 ( .A1(n11528), .A2(n15472), .ZN(n12043) );
  NAND2_X1 U11580 ( .A1(n18972), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12508) );
  NAND3_X1 U11581 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n17099), .ZN(n17283) );
  AND2_X2 U11582 ( .A1(n10190), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11528) );
  AND3_X2 U11583 ( .A1(n10438), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10647) );
  AND2_X1 U11584 ( .A1(n11526), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11530) );
  AND3_X2 U11585 ( .A1(n9840), .A2(n10438), .A3(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10646) );
  AND3_X2 U11586 ( .A1(n10144), .A2(n10438), .A3(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n9847) );
  AND2_X4 U11587 ( .A1(n13958), .A2(n10328), .ZN(n11573) );
  AND3_X2 U11588 ( .A1(n10438), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n9854) );
  NOR2_X2 U11589 ( .A1(n10405), .A2(n14064), .ZN(n10407) );
  INV_X1 U11590 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n14064) );
  INV_X4 U11591 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10438) );
  AND2_X2 U11592 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10436) );
  NOR2_X2 U11593 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20769) );
  NOR2_X1 U11594 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n17099) );
  INV_X1 U11595 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13554) );
  NOR2_X1 U11596 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11537) );
  AND2_X1 U11597 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13945) );
  OAI21_X2 U11598 ( .B1(n10315), .B2(n10314), .A(n10312), .ZN(n15935) );
  NOR2_X2 U11599 ( .A1(n15689), .A2(n10155), .ZN(n10159) );
  OR2_X1 U11600 ( .A1(n14432), .A2(n14431), .ZN(n15689) );
  NOR2_X2 U11601 ( .A1(n16019), .A2(n16034), .ZN(n16000) );
  AND2_X1 U11602 ( .A1(n11171), .A2(n11172), .ZN(n19461) );
  OAI21_X1 U11603 ( .B1(n11006), .B2(n11499), .A(n11002), .ZN(n11137) );
  OAI211_X1 U11604 ( .C1(n11006), .C2(n16105), .A(n10992), .B(n10991), .ZN(
        n11145) );
  NOR2_X2 U11605 ( .A1(n15023), .A2(n15026), .ZN(n14962) );
  NOR2_X2 U11606 ( .A1(n14387), .A2(n14494), .ZN(n14456) );
  INV_X1 U11607 ( .A(n10268), .ZN(n9830) );
  AND2_X2 U11608 ( .A1(n9831), .A2(n13702), .ZN(n13829) );
  NOR2_X1 U11609 ( .A1(n13814), .A2(n9830), .ZN(n9831) );
  NOR2_X1 U11610 ( .A1(n14730), .A2(n14728), .ZN(n9832) );
  CLKBUF_X1 U11611 ( .A(n20243), .Z(n9833) );
  AND2_X1 U11612 ( .A1(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n13006), .ZN(
        n9835) );
  INV_X1 U11613 ( .A(n15128), .ZN(n9834) );
  NAND2_X1 U11614 ( .A1(n9834), .A2(n13006), .ZN(n9836) );
  NAND2_X1 U11615 ( .A1(n20245), .A2(n20244), .ZN(n20243) );
  NAND2_X1 U11616 ( .A1(n9982), .A2(n11881), .ZN(n16329) );
  AND2_X2 U11617 ( .A1(n14363), .A2(n14434), .ZN(n9947) );
  XNOR2_X1 U11618 ( .A(n11852), .B(n20273), .ZN(n13850) );
  AND3_X1 U11619 ( .A1(n13003), .A2(n9937), .A3(n15146), .ZN(n15129) );
  INV_X1 U11620 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n9840) );
  AND2_X4 U11621 ( .A1(n10308), .A2(n14088), .ZN(n10649) );
  NAND2_X2 U11622 ( .A1(n10963), .A2(n10973), .ZN(n14090) );
  NAND2_X2 U11623 ( .A1(n13578), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13579) );
  XNOR2_X2 U11624 ( .A(n11840), .B(n11841), .ZN(n13578) );
  INV_X2 U11625 ( .A(n10657), .ZN(n20064) );
  AND2_X1 U11626 ( .A1(n10435), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n9841) );
  INV_X1 U11627 ( .A(n9841), .ZN(n9842) );
  NAND2_X2 U11628 ( .A1(n13533), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n11840) );
  AND2_X2 U11629 ( .A1(n10436), .A2(n14088), .ZN(n9843) );
  NAND2_X2 U11630 ( .A1(n13579), .A2(n11842), .ZN(n11843) );
  INV_X1 U11631 ( .A(n11654), .ZN(n11670) );
  AND3_X1 U11632 ( .A1(n10144), .A2(n10438), .A3(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n9846) );
  AND2_X1 U11633 ( .A1(n11710), .A2(n11708), .ZN(n11678) );
  INV_X1 U11634 ( .A(n13564), .ZN(n14805) );
  OR2_X1 U11635 ( .A1(n13002), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15155) );
  AND2_X2 U11636 ( .A1(n11530), .A2(n15472), .ZN(n12724) );
  AND2_X2 U11637 ( .A1(n11530), .A2(n15472), .ZN(n9849) );
  NAND2_X1 U11638 ( .A1(n15137), .A2(n15314), .ZN(n15128) );
  NAND2_X1 U11639 ( .A1(n13848), .A2(n11853), .ZN(n20245) );
  NOR2_X2 U11640 ( .A1(n11653), .A2(n11652), .ZN(n11669) );
  NAND2_X2 U11641 ( .A1(n11635), .A2(n11816), .ZN(n11598) );
  AND2_X2 U11642 ( .A1(n11530), .A2(n15472), .ZN(n9848) );
  NAND4_X2 U11643 ( .A1(n13598), .A2(n13597), .A3(n13623), .A4(n13596), .ZN(
        n13702) );
  AND2_X4 U11644 ( .A1(n10328), .A2(n15472), .ZN(n11622) );
  XNOR2_X2 U11645 ( .A(n11295), .B(n14488), .ZN(n14484) );
  OAI21_X2 U11646 ( .B1(n11447), .B2(n12808), .A(n19153), .ZN(n11295) );
  NOR2_X4 U11647 ( .A1(n15796), .A2(n15922), .ZN(n15771) );
  AOI21_X2 U11648 ( .B1(n14822), .B2(n14821), .A(n14820), .ZN(n15134) );
  NOR2_X1 U11649 ( .A1(n14833), .A2(n10348), .ZN(n14820) );
  AND3_X1 U11650 ( .A1(n11172), .A2(n14805), .A3(n19354), .ZN(n11188) );
  AND2_X1 U11651 ( .A1(n11172), .A2(n19342), .ZN(n11177) );
  AOI21_X2 U11652 ( .B1(n10087), .B2(n10085), .A(n10084), .ZN(n16019) );
  NAND2_X2 U11653 ( .A1(n14478), .A2(n10081), .ZN(n10087) );
  NAND2_X2 U11654 ( .A1(n11297), .A2(n11296), .ZN(n14410) );
  NAND2_X2 U11655 ( .A1(n13735), .A2(n11844), .ZN(n11852) );
  NOR2_X2 U11656 ( .A1(n15645), .A2(n14707), .ZN(n14727) );
  NAND2_X2 U11657 ( .A1(n10300), .A2(n10299), .ZN(n15263) );
  AND2_X1 U11658 ( .A1(n13627), .A2(n19198), .ZN(n11169) );
  NOR2_X1 U11659 ( .A1(n13627), .A2(n14093), .ZN(n11172) );
  NAND3_X2 U11660 ( .A1(n10265), .A2(n10263), .A3(n11143), .ZN(n13627) );
  NAND2_X2 U11661 ( .A1(n11725), .A2(n11724), .ZN(n10282) );
  NOR2_X4 U11662 ( .A1(n13660), .A2(n13661), .ZN(n13662) );
  AND2_X2 U11663 ( .A1(n13829), .A2(n13831), .ZN(n14030) );
  INV_X2 U11664 ( .A(n10936), .ZN(n10938) );
  NAND2_X2 U11665 ( .A1(n10639), .A2(n10638), .ZN(n10936) );
  INV_X4 U11666 ( .A(n11006), .ZN(n11053) );
  NOR2_X2 U11667 ( .A1(n15678), .A2(n15679), .ZN(n15672) );
  INV_X2 U11668 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n14088) );
  AND2_X4 U11669 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10435) );
  XNOR2_X1 U11670 ( .A(n11168), .B(n11167), .ZN(n13415) );
  INV_X2 U11671 ( .A(n14287), .ZN(n15661) );
  NOR2_X1 U11672 ( .A1(n10058), .A2(n10061), .ZN(n10059) );
  NAND2_X1 U11673 ( .A1(n11652), .A2(n11644), .ZN(n11765) );
  NAND2_X1 U11674 ( .A1(n12516), .A2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12514) );
  INV_X1 U11675 ( .A(n19040), .ZN(n13386) );
  CLKBUF_X1 U11676 ( .A(n12038), .Z(n12116) );
  BUF_X1 U11677 ( .A(n11612), .Z(n12374) );
  NAND2_X1 U11678 ( .A1(n12752), .A2(n12941), .ZN(n10044) );
  NAND4_X1 U11679 ( .A1(n10041), .A2(n10040), .A3(n11659), .A4(n13518), .ZN(
        n10039) );
  AND2_X1 U11680 ( .A1(n11675), .A2(n9916), .ZN(n10041) );
  NAND2_X1 U11681 ( .A1(n11661), .A2(n10038), .ZN(n10037) );
  INV_X1 U11682 ( .A(n12978), .ZN(n10174) );
  INV_X1 U11683 ( .A(n10321), .ZN(n10320) );
  NOR2_X1 U11684 ( .A1(n10959), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n10712) );
  NOR2_X1 U11685 ( .A1(n9869), .A2(n10005), .ZN(n10004) );
  INV_X1 U11686 ( .A(n10295), .ZN(n10294) );
  OAI21_X1 U11687 ( .B1(n9845), .B2(n10297), .A(n10296), .ZN(n10295) );
  NAND2_X1 U11688 ( .A1(n16302), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n10297) );
  AND2_X1 U11689 ( .A1(n9845), .A2(n15432), .ZN(n10298) );
  NOR2_X2 U11690 ( .A1(n16195), .A2(n12934), .ZN(n12923) );
  NAND2_X1 U11691 ( .A1(n11645), .A2(n11644), .ZN(n12929) );
  NAND2_X1 U11692 ( .A1(n12929), .A2(n12848), .ZN(n12849) );
  NAND2_X1 U11693 ( .A1(n11705), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11959) );
  AND2_X1 U11694 ( .A1(n9933), .A2(n11896), .ZN(n11817) );
  NAND2_X1 U11695 ( .A1(n10262), .A2(n10261), .ZN(n13592) );
  NAND2_X1 U11696 ( .A1(n9862), .A2(n13350), .ZN(n10261) );
  NAND2_X1 U11697 ( .A1(n11481), .A2(n10072), .ZN(n10071) );
  INV_X1 U11698 ( .A(n11379), .ZN(n10072) );
  NAND2_X1 U11699 ( .A1(n10064), .A2(n10062), .ZN(n11324) );
  AOI21_X1 U11700 ( .B1(n10067), .B2(n10065), .A(n10063), .ZN(n10062) );
  INV_X1 U11701 ( .A(n16514), .ZN(n10063) );
  INV_X1 U11702 ( .A(n11291), .ZN(n10074) );
  OAI21_X1 U11703 ( .B1(n10957), .B2(n14112), .A(n10956), .ZN(n11470) );
  NAND2_X1 U11704 ( .A1(n10712), .A2(n10680), .ZN(n10890) );
  AOI21_X1 U11705 ( .B1(n12610), .B2(n12609), .A(n12608), .ZN(n13188) );
  AOI21_X1 U11706 ( .B1(n18847), .B2(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(
        n12613), .ZN(n13192) );
  NAND2_X1 U11707 ( .A1(n13762), .A2(n20331), .ZN(n13774) );
  NOR2_X1 U11708 ( .A1(n10387), .A2(n12790), .ZN(n10386) );
  OR2_X1 U11709 ( .A1(n14108), .A2(n14106), .ZN(n13689) );
  AND2_X1 U11710 ( .A1(n12490), .A2(n10923), .ZN(n10218) );
  OR2_X1 U11711 ( .A1(n19216), .A2(n19327), .ZN(n10219) );
  AND2_X1 U11712 ( .A1(n11089), .A2(n11088), .ZN(n11467) );
  NAND2_X1 U11713 ( .A1(n15988), .A2(n15987), .ZN(n15828) );
  NAND2_X1 U11714 ( .A1(n19431), .A2(n19207), .ZN(n19568) );
  OR2_X1 U11715 ( .A1(n19431), .A2(n19207), .ZN(n19782) );
  OR2_X1 U11716 ( .A1(n19431), .A2(n20040), .ZN(n19802) );
  NOR2_X1 U11717 ( .A1(n16153), .A2(n12516), .ZN(n12651) );
  INV_X1 U11718 ( .A(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n21140) );
  NAND2_X1 U11719 ( .A1(n18972), .A2(n18982), .ZN(n9980) );
  OAI21_X1 U11720 ( .B1(n16149), .B2(n16150), .A(n9911), .ZN(n16231) );
  AND2_X1 U11721 ( .A1(n17742), .A2(n10356), .ZN(n13165) );
  NAND2_X1 U11722 ( .A1(n13164), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n9974) );
  INV_X1 U11723 ( .A(n17551), .ZN(n16624) );
  NAND2_X1 U11724 ( .A1(n18409), .A2(n18405), .ZN(n13246) );
  NAND2_X1 U11725 ( .A1(n18838), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n16153) );
  NAND2_X1 U11726 ( .A1(n12786), .A2(n12785), .ZN(n19042) );
  NAND2_X1 U11727 ( .A1(P3_EAX_REG_24__SCAN_IN), .A2(P3_EAX_REG_25__SCAN_IN), 
        .ZN(n10006) );
  NAND2_X1 U11728 ( .A1(n17432), .A2(P3_EAX_REG_0__SCAN_IN), .ZN(n17576) );
  NAND2_X1 U11729 ( .A1(n16234), .A2(n17432), .ZN(n17580) );
  NAND3_X1 U11730 ( .A1(n16624), .A2(n18804), .A3(n18359), .ZN(n18211) );
  AOI21_X1 U11731 ( .B1(n12729), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A(
        n10031), .ZN(n11785) );
  AND2_X1 U11732 ( .A1(n10016), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n10031) );
  NAND2_X1 U11733 ( .A1(n11021), .A2(P2_EBX_REG_1__SCAN_IN), .ZN(n10079) );
  NAND2_X1 U11734 ( .A1(n10947), .A2(n11485), .ZN(n10217) );
  AND2_X1 U11735 ( .A1(n10016), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n10027) );
  AND2_X1 U11736 ( .A1(n10016), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n10035) );
  AND2_X1 U11737 ( .A1(n10016), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n10025) );
  CLKBUF_X1 U11738 ( .A(n12392), .Z(n12730) );
  AOI21_X1 U11739 ( .B1(n9838), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .A(
        n10018), .ZN(n11805) );
  AND2_X1 U11740 ( .A1(n10016), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n10018) );
  OR2_X1 U11741 ( .A1(n11690), .A2(n11689), .ZN(n11834) );
  OR2_X1 U11742 ( .A1(n11776), .A2(n11775), .ZN(n11865) );
  NOR2_X1 U11743 ( .A1(n13554), .A2(n20310), .ZN(n10038) );
  INV_X1 U11744 ( .A(n11959), .ZN(n11968) );
  AND2_X1 U11745 ( .A1(n10492), .A2(n10491), .ZN(n10494) );
  NOR2_X1 U11746 ( .A1(n11325), .A2(n10188), .ZN(n10187) );
  NOR2_X1 U11747 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n14624) );
  NOR2_X1 U11748 ( .A1(n10225), .A2(n10224), .ZN(n10223) );
  INV_X1 U11749 ( .A(n10668), .ZN(n10225) );
  OAI21_X1 U11750 ( .B1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(n15753), .ZN(n12473) );
  OR2_X1 U11751 ( .A1(n10443), .A2(n10442), .ZN(n11439) );
  OR2_X1 U11752 ( .A1(n11153), .A2(n11137), .ZN(n11138) );
  OR2_X1 U11753 ( .A1(n11432), .A2(n10182), .ZN(n11205) );
  AND2_X1 U11754 ( .A1(n13627), .A2(n11156), .ZN(n11162) );
  NOR2_X1 U11755 ( .A1(n10364), .A2(n17581), .ZN(n13210) );
  AOI21_X1 U11756 ( .B1(n18620), .B2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n12604), .ZN(n12610) );
  OAI22_X1 U11757 ( .A1(n18982), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B1(
        n18845), .B2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n12609) );
  OR2_X1 U11758 ( .A1(n12757), .A2(n16192), .ZN(n12938) );
  NOR2_X1 U11759 ( .A1(n9879), .A2(n10339), .ZN(n10337) );
  INV_X1 U11760 ( .A(n10342), .ZN(n10341) );
  OR2_X1 U11761 ( .A1(n11722), .A2(n11721), .ZN(n11833) );
  NAND2_X1 U11762 ( .A1(n10201), .A2(n14520), .ZN(n10200) );
  INV_X1 U11763 ( .A(n14845), .ZN(n10201) );
  NOR2_X1 U11764 ( .A1(n10196), .A2(n14917), .ZN(n10195) );
  INV_X1 U11765 ( .A(n14934), .ZN(n10196) );
  NAND2_X1 U11766 ( .A1(n12905), .A2(n10205), .ZN(n10204) );
  INV_X1 U11767 ( .A(n14985), .ZN(n10205) );
  INV_X1 U11768 ( .A(n15248), .ZN(n10050) );
  NAND2_X1 U11769 ( .A1(n13548), .A2(n12934), .ZN(n12927) );
  OR2_X1 U11770 ( .A1(n11703), .A2(n11702), .ZN(n11896) );
  NAND2_X1 U11771 ( .A1(n11734), .A2(n11733), .ZN(n11819) );
  OR2_X1 U11772 ( .A1(n11831), .A2(n11732), .ZN(n11733) );
  XNOR2_X1 U11773 ( .A(n10056), .B(n11760), .ZN(n11820) );
  OAI211_X1 U11774 ( .C1(n11747), .C2(n10053), .A(n10054), .B(n10052), .ZN(
        n10056) );
  INV_X1 U11775 ( .A(n10013), .ZN(n11779) );
  NAND2_X1 U11776 ( .A1(n11764), .A2(n11763), .ZN(n20460) );
  OR2_X1 U11777 ( .A1(n11742), .A2(n11535), .ZN(n11764) );
  AND2_X1 U11778 ( .A1(n20732), .A2(n20696), .ZN(n20656) );
  OAI21_X1 U11779 ( .B1(n13964), .B2(n13963), .A(n15481), .ZN(n20309) );
  AND2_X1 U11780 ( .A1(n10543), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n11343) );
  AND2_X1 U11781 ( .A1(n10543), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n11329) );
  AND2_X1 U11782 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10437) );
  INV_X1 U11783 ( .A(n15523), .ZN(n10258) );
  NAND2_X1 U11784 ( .A1(n9949), .A2(n15657), .ZN(n10271) );
  AND2_X1 U11785 ( .A1(n14561), .A2(n10371), .ZN(n10278) );
  INV_X1 U11786 ( .A(n14413), .ZN(n10234) );
  OAI21_X1 U11787 ( .B1(n11429), .B2(n10890), .A(n10683), .ZN(n13367) );
  NOR2_X1 U11788 ( .A1(n15765), .A2(n10143), .ZN(n10142) );
  INV_X1 U11789 ( .A(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n10143) );
  NOR2_X1 U11790 ( .A1(n15845), .A2(n10141), .ZN(n10140) );
  INV_X1 U11791 ( .A(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n10141) );
  NOR2_X1 U11792 ( .A1(n15862), .A2(n10132), .ZN(n10131) );
  INV_X1 U11793 ( .A(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n10132) );
  OR2_X1 U11794 ( .A1(n11254), .A2(n16573), .ZN(n11458) );
  INV_X1 U11795 ( .A(n12432), .ZN(n10247) );
  AND2_X1 U11796 ( .A1(n16015), .A2(n10238), .ZN(n10237) );
  NAND2_X1 U11797 ( .A1(n10239), .A2(n10240), .ZN(n10238) );
  INV_X1 U11798 ( .A(n10244), .ZN(n10239) );
  AOI21_X1 U11799 ( .B1(n10318), .B2(n10320), .A(n10069), .ZN(n10068) );
  INV_X1 U11800 ( .A(n15865), .ZN(n10069) );
  INV_X1 U11801 ( .A(n13819), .ZN(n10152) );
  OAI21_X1 U11802 ( .B1(n11291), .B2(n11290), .A(n10310), .ZN(n11253) );
  NAND2_X1 U11803 ( .A1(n11438), .A2(n11437), .ZN(n11441) );
  AOI21_X1 U11804 ( .B1(n11013), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n11012), .ZN(n11015) );
  AND2_X1 U11805 ( .A1(n11019), .A2(n13609), .ZN(n10146) );
  INV_X1 U11806 ( .A(n10706), .ZN(n10249) );
  AND2_X1 U11807 ( .A1(n13627), .A2(n11151), .ZN(n11160) );
  AND2_X1 U11808 ( .A1(n14805), .A2(n9860), .ZN(n11171) );
  NAND2_X1 U11809 ( .A1(n10448), .A2(n10607), .ZN(n10456) );
  INV_X1 U11810 ( .A(n10450), .ZN(n10455) );
  NAND2_X1 U11811 ( .A1(n12506), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12507) );
  INV_X1 U11812 ( .A(n17340), .ZN(n13068) );
  NOR2_X1 U11813 ( .A1(n17283), .A2(n13091), .ZN(n13092) );
  AND2_X1 U11814 ( .A1(n17343), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n13088) );
  OAI211_X1 U11815 ( .C1(n12537), .C2(n9977), .A(n9976), .B(n9912), .ZN(n9975)
         );
  INV_X1 U11816 ( .A(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n9977) );
  NAND2_X1 U11817 ( .A1(n17386), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n9976) );
  AND2_X1 U11818 ( .A1(n17378), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n12545) );
  NAND2_X1 U11819 ( .A1(n18621), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13190) );
  OR2_X1 U11820 ( .A1(n13179), .A2(n16731), .ZN(n16146) );
  NOR2_X1 U11821 ( .A1(n17857), .A2(n10114), .ZN(n10113) );
  INV_X1 U11822 ( .A(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n10114) );
  INV_X1 U11823 ( .A(n16908), .ZN(n16896) );
  NAND2_X1 U11824 ( .A1(n17846), .A2(n13160), .ZN(n13161) );
  AND2_X1 U11825 ( .A1(n10001), .A2(n10000), .ZN(n13186) );
  NAND2_X1 U11826 ( .A1(n13183), .A2(n18397), .ZN(n10000) );
  NOR2_X1 U11827 ( .A1(n13244), .A2(n13243), .ZN(n10001) );
  XNOR2_X1 U11828 ( .A(n17581), .B(n17568), .ZN(n13135) );
  XNOR2_X1 U11829 ( .A(n13210), .B(n17568), .ZN(n13211) );
  OAI22_X1 U11830 ( .A1(n12506), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B1(
        n18620), .B2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13191) );
  NAND2_X1 U11831 ( .A1(n13128), .A2(n10355), .ZN(n13129) );
  NAND2_X1 U11832 ( .A1(n17379), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n13128) );
  NAND2_X1 U11833 ( .A1(n17379), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n10125) );
  NOR2_X1 U11834 ( .A1(n9901), .A2(n10122), .ZN(n10121) );
  OAI211_X1 U11835 ( .C1(n13050), .C2(n21237), .A(n10124), .B(n10123), .ZN(
        n10122) );
  NAND2_X1 U11836 ( .A1(n12552), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n10123) );
  INV_X1 U11837 ( .A(n12005), .ZN(n12748) );
  AND2_X1 U11838 ( .A1(n12698), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12699) );
  NAND2_X1 U11839 ( .A1(n12699), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12845) );
  NAND2_X1 U11840 ( .A1(n12328), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n12368) );
  NAND2_X1 U11841 ( .A1(n12247), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12281) );
  INV_X1 U11842 ( .A(n15120), .ZN(n13005) );
  NAND2_X1 U11843 ( .A1(n15129), .A2(n15315), .ZN(n15120) );
  NOR3_X1 U11844 ( .A1(n14861), .A2(n10199), .A3(n10200), .ZN(n14819) );
  OR2_X1 U11845 ( .A1(n14837), .A2(n14817), .ZN(n10199) );
  NOR2_X1 U11846 ( .A1(n14903), .A2(n14891), .ZN(n14892) );
  AND2_X1 U11847 ( .A1(n15398), .A2(n15290), .ZN(n15367) );
  AND2_X1 U11848 ( .A1(n12917), .A2(n12916), .ZN(n14905) );
  NOR2_X1 U11849 ( .A1(n9887), .A2(n15007), .ZN(n15009) );
  NAND2_X1 U11850 ( .A1(n9837), .A2(n9988), .ZN(n9990) );
  INV_X1 U11851 ( .A(n10298), .ZN(n9989) );
  AND2_X1 U11852 ( .A1(n10359), .A2(n11900), .ZN(n10299) );
  NAND2_X1 U11853 ( .A1(n10057), .A2(n11885), .ZN(n11879) );
  INV_X1 U11854 ( .A(n11861), .ZN(n10289) );
  NAND2_X1 U11855 ( .A1(n13780), .A2(n20298), .ZN(n16400) );
  INV_X1 U11856 ( .A(n13514), .ZN(n10043) );
  INV_X1 U11857 ( .A(n11668), .ZN(n11647) );
  OR2_X1 U11858 ( .A1(n13774), .A2(n16195), .ZN(n13458) );
  AND2_X1 U11859 ( .A1(n13769), .A2(n13768), .ZN(n13795) );
  OR2_X1 U11860 ( .A1(n12757), .A2(n11633), .ZN(n15468) );
  INV_X1 U11861 ( .A(n20086), .ZN(n13768) );
  NOR2_X1 U11862 ( .A1(n20657), .A2(n20469), .ZN(n20803) );
  INV_X1 U11863 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20846) );
  NAND2_X1 U11864 ( .A1(n20310), .A2(n20309), .ZN(n20469) );
  INV_X1 U11865 ( .A(n20652), .ZN(n20794) );
  OR2_X1 U11866 ( .A1(n20593), .A2(n13974), .ZN(n20855) );
  AOI21_X1 U11867 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n20767), .A(n20469), 
        .ZN(n20856) );
  AND2_X1 U11868 ( .A1(n11977), .A2(n11976), .ZN(n16193) );
  NAND2_X1 U11869 ( .A1(n11939), .A2(n12758), .ZN(n11977) );
  OAI21_X1 U11870 ( .B1(n10182), .B2(n11379), .A(n10181), .ZN(n11400) );
  NAND2_X1 U11871 ( .A1(n11379), .A2(n11373), .ZN(n10181) );
  NOR2_X1 U11872 ( .A1(n12470), .A2(n12471), .ZN(n12469) );
  NAND2_X1 U11873 ( .A1(n12804), .A2(n12466), .ZN(n12470) );
  NOR2_X1 U11874 ( .A1(n15549), .A2(n19159), .ZN(n15532) );
  OR2_X1 U11875 ( .A1(n15532), .A2(n15533), .ZN(n10130) );
  NAND2_X1 U11876 ( .A1(n11135), .A2(n10184), .ZN(n15536) );
  NAND2_X1 U11877 ( .A1(n10256), .A2(n16060), .ZN(n10255) );
  INV_X1 U11878 ( .A(n15620), .ZN(n10256) );
  AND2_X1 U11879 ( .A1(n15569), .A2(n15570), .ZN(n15572) );
  AND2_X1 U11880 ( .A1(n10897), .A2(n10254), .ZN(n10253) );
  INV_X1 U11881 ( .A(n14381), .ZN(n10254) );
  AND3_X1 U11882 ( .A1(n10744), .A2(n10743), .A3(n10742), .ZN(n14160) );
  INV_X1 U11883 ( .A(n10719), .ZN(n14481) );
  XNOR2_X1 U11884 ( .A(n10384), .B(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n12834) );
  AOI21_X1 U11885 ( .B1(n15842), .B2(n15841), .A(n11347), .ZN(n15988) );
  AND2_X1 U11886 ( .A1(n11052), .A2(n11051), .ZN(n13812) );
  INV_X1 U11887 ( .A(n14408), .ZN(n10306) );
  XNOR2_X1 U11888 ( .A(n10170), .B(n12810), .ZN(n12839) );
  NAND2_X1 U11889 ( .A1(n10154), .A2(n10153), .ZN(n12817) );
  INV_X1 U11890 ( .A(n11124), .ZN(n10153) );
  AND2_X1 U11891 ( .A1(n10161), .A2(n9951), .ZN(n10160) );
  INV_X1 U11892 ( .A(n15522), .ZN(n10161) );
  AND2_X1 U11893 ( .A1(n10313), .A2(n15950), .ZN(n10312) );
  OR2_X1 U11894 ( .A1(n12440), .A2(n10314), .ZN(n10313) );
  INV_X1 U11895 ( .A(n15951), .ZN(n10314) );
  NOR2_X1 U11896 ( .A1(n10302), .A2(n15990), .ZN(n10096) );
  NAND2_X1 U11897 ( .A1(n10303), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n10302) );
  INV_X1 U11898 ( .A(n10305), .ZN(n10303) );
  NAND2_X1 U11899 ( .A1(n10157), .A2(n10156), .ZN(n10155) );
  INV_X1 U11900 ( .A(n15688), .ZN(n10156) );
  NOR2_X1 U11901 ( .A1(n11467), .A2(n10158), .ZN(n10157) );
  NAND2_X1 U11903 ( .A1(n16075), .A2(n16076), .ZN(n16074) );
  AOI21_X1 U11904 ( .B1(n11313), .B2(n11306), .A(n9913), .ZN(n10321) );
  NOR2_X1 U11905 ( .A1(n13868), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10230) );
  NAND2_X1 U11906 ( .A1(n11259), .A2(n10231), .ZN(n10229) );
  AOI21_X1 U11907 ( .B1(n13868), .B2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        n10232), .ZN(n10231) );
  INV_X1 U11908 ( .A(n14068), .ZN(n10232) );
  NAND2_X1 U11909 ( .A1(n11155), .A2(n11003), .ZN(n11004) );
  OAI21_X1 U11910 ( .B1(n11155), .B2(n11003), .A(n11152), .ZN(n11005) );
  NAND2_X1 U11911 ( .A1(n10147), .A2(n10146), .ZN(n13612) );
  AND3_X1 U11912 ( .A1(n19332), .A2(n11507), .A3(n19349), .ZN(n14054) );
  AND2_X1 U11913 ( .A1(n11426), .A2(n13386), .ZN(n11505) );
  OR2_X1 U11914 ( .A1(n10706), .A2(n10703), .ZN(n13914) );
  AOI21_X1 U11915 ( .B1(n13451), .B2(n10702), .A(n10701), .ZN(n10706) );
  AOI21_X1 U11916 ( .B1(n13582), .B2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n13352), .ZN(n13353) );
  NAND2_X1 U11917 ( .A1(n14093), .A2(n13587), .ZN(n13354) );
  INV_X1 U11918 ( .A(n20002), .ZN(n20006) );
  OR2_X1 U11919 ( .A1(n19364), .A2(n20029), .ZN(n19667) );
  INV_X1 U11920 ( .A(n11217), .ZN(n14295) );
  OR2_X1 U11921 ( .A1(n19364), .A2(n20026), .ZN(n20004) );
  NAND2_X1 U11922 ( .A1(n19364), .A2(n20026), .ZN(n19781) );
  NAND2_X1 U11923 ( .A1(n11386), .A2(n11385), .ZN(n14108) );
  INV_X1 U11924 ( .A(n11387), .ZN(n11386) );
  NOR4_X1 U11925 ( .A1(n18401), .A2(n18397), .A3(n13246), .A4(n13173), .ZN(
        n13184) );
  NOR2_X1 U11926 ( .A1(n17100), .A2(n17083), .ZN(n16909) );
  INV_X1 U11927 ( .A(n18409), .ZN(n17433) );
  NAND2_X1 U11928 ( .A1(n17099), .A2(n12510), .ZN(n17252) );
  NOR2_X1 U11929 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n12510) );
  NOR2_X1 U11930 ( .A1(n12561), .A2(n21208), .ZN(n13056) );
  AOI21_X1 U11931 ( .B1(n13080), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A(
        n10169), .ZN(n13049) );
  AND2_X1 U11932 ( .A1(n17344), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n10169) );
  OR2_X1 U11933 ( .A1(n17921), .A2(n17924), .ZN(n17900) );
  NOR2_X1 U11934 ( .A1(n18008), .A2(n13142), .ZN(n17995) );
  NOR2_X2 U11935 ( .A1(n18811), .A2(n18864), .ZN(n13232) );
  NAND2_X1 U11936 ( .A1(n13144), .A2(n17553), .ZN(n16638) );
  NAND2_X1 U11937 ( .A1(n10165), .A2(n13151), .ZN(n10163) );
  AOI22_X1 U11938 ( .A1(n13153), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B1(
        n17957), .B2(n18181), .ZN(n9973) );
  NOR2_X1 U11939 ( .A1(n13251), .A2(n13245), .ZN(n18804) );
  OR3_X1 U11940 ( .A1(n12754), .A2(n20086), .A3(n16210), .ZN(n13637) );
  AND2_X1 U11941 ( .A1(n13837), .A2(n13836), .ZN(n20154) );
  CLKBUF_X1 U11942 ( .A(n13971), .Z(n20593) );
  INV_X1 U11943 ( .A(n20465), .ZN(n20490) );
  OR2_X1 U11944 ( .A1(n14115), .A2(n10655), .ZN(n13421) );
  NAND2_X1 U11945 ( .A1(n13421), .A2(n19208), .ZN(n20056) );
  XNOR2_X1 U11946 ( .A(n13626), .B(n13625), .ZN(n19431) );
  AND2_X1 U11947 ( .A1(n13624), .A2(n13623), .ZN(n13625) );
  OAI21_X1 U11948 ( .B1(n13622), .B2(n13621), .A(n13620), .ZN(n13626) );
  XNOR2_X1 U11949 ( .A(n12823), .B(n12822), .ZN(n19216) );
  NAND2_X1 U11950 ( .A1(n12823), .A2(n10926), .ZN(n14786) );
  INV_X1 U11951 ( .A(n19274), .ZN(n19257) );
  NAND2_X1 U11952 ( .A1(n19042), .A2(n12787), .ZN(n16559) );
  AND2_X1 U11953 ( .A1(n16559), .A2(n20024), .ZN(n19315) );
  XNOR2_X1 U11954 ( .A(n12798), .B(n12797), .ZN(n12844) );
  XNOR2_X1 U11955 ( .A(n10221), .B(n10220), .ZN(n15814) );
  INV_X1 U11956 ( .A(n11362), .ZN(n10220) );
  OAI21_X1 U11957 ( .B1(n15816), .B2(n12430), .A(n15817), .ZN(n10221) );
  INV_X1 U11958 ( .A(n19353), .ZN(n16561) );
  INV_X1 U11959 ( .A(n19331), .ZN(n19363) );
  INV_X1 U11960 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20043) );
  INV_X1 U11961 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n20034) );
  INV_X1 U11962 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20033) );
  INV_X1 U11963 ( .A(n20029), .ZN(n20026) );
  INV_X1 U11964 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20017) );
  NAND2_X1 U11965 ( .A1(n19364), .A2(n20029), .ZN(n20001) );
  XNOR2_X1 U11966 ( .A(n13621), .B(n13619), .ZN(n19364) );
  AND2_X1 U11967 ( .A1(n13584), .A2(n13583), .ZN(n19643) );
  NOR2_X1 U11968 ( .A1(n17175), .A2(n10126), .ZN(n17160) );
  OR3_X1 U11969 ( .A1(n10127), .A2(n17121), .A3(n17120), .ZN(n10126) );
  NOR2_X1 U11970 ( .A1(n19012), .A2(n10129), .ZN(n10128) );
  NAND2_X1 U11971 ( .A1(n18378), .A2(n19020), .ZN(n10129) );
  NOR2_X2 U11972 ( .A1(n17547), .A2(n17425), .ZN(n17426) );
  AND2_X1 U11973 ( .A1(n17454), .A2(P3_EAX_REG_27__SCAN_IN), .ZN(n17447) );
  NOR2_X1 U11974 ( .A1(n21227), .A2(n9885), .ZN(n17454) );
  NOR2_X2 U11975 ( .A1(n18405), .A2(n17571), .ZN(n17500) );
  NOR2_X1 U11976 ( .A1(n17514), .A2(n17688), .ZN(n17510) );
  AOI22_X1 U11977 ( .A1(n13089), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17385), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12524) );
  AOI211_X1 U11978 ( .C1(n13079), .C2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A(
        n12522), .B(n12521), .ZN(n12523) );
  NOR2_X1 U11979 ( .A1(n17616), .A2(n17549), .ZN(n17542) );
  AOI211_X2 U11980 ( .C1(n17378), .C2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A(
        n13037), .B(n13036), .ZN(n17551) );
  INV_X1 U11981 ( .A(n17571), .ZN(n17575) );
  NOR2_X1 U11982 ( .A1(n18802), .A2(n9998), .ZN(n9997) );
  INV_X1 U11983 ( .A(n17567), .ZN(n17578) );
  NAND2_X1 U11984 ( .A1(n10177), .A2(n10180), .ZN(n17709) );
  INV_X1 U11985 ( .A(n18211), .ZN(n18287) );
  AOI21_X2 U11986 ( .B1(n16148), .B2(n13255), .A(n18864), .ZN(n18359) );
  AND2_X1 U11987 ( .A1(n20767), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11944) );
  AOI21_X1 U11988 ( .B1(n12286), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .A(
        n10026), .ZN(n12358) );
  AND2_X1 U11989 ( .A1(n10016), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n10026) );
  AOI21_X1 U11990 ( .B1(n12286), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .A(
        n10023), .ZN(n11797) );
  AND2_X1 U11991 ( .A1(n10016), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n10023) );
  AOI21_X1 U11992 ( .B1(n12286), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .A(
        n10021), .ZN(n11753) );
  AND2_X1 U11993 ( .A1(n9821), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(
        n10021) );
  NAND2_X1 U11994 ( .A1(n11584), .A2(n11643), .ZN(n11639) );
  AOI21_X1 U11995 ( .B1(n12286), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .A(
        n10022), .ZN(n11772) );
  AND2_X1 U11996 ( .A1(n10016), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n10022) );
  NOR2_X1 U11997 ( .A1(n11964), .A2(n11963), .ZN(n12762) );
  AND4_X1 U11998 ( .A1(n11214), .A2(n11213), .A3(n11212), .A4(n11211), .ZN(
        n11229) );
  OAI21_X1 U11999 ( .B1(n11238), .B2(n11170), .A(n10309), .ZN(n11176) );
  NAND2_X1 U12000 ( .A1(n11217), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n10309) );
  AOI21_X1 U12001 ( .B1(n9852), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A(n10019), .ZN(n12256) );
  AND2_X1 U12002 ( .A1(n10016), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n10019) );
  AOI21_X1 U12003 ( .B1(n12729), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .A(
        n10034), .ZN(n12216) );
  AND2_X1 U12004 ( .A1(n10016), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n10034) );
  AOI21_X1 U12005 ( .B1(n9848), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A(
        n10030), .ZN(n12170) );
  AND2_X1 U12006 ( .A1(n10016), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n10030) );
  AOI21_X1 U12007 ( .B1(n12729), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .A(
        n10033), .ZN(n12151) );
  AND2_X1 U12008 ( .A1(n10016), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n10033) );
  AOI21_X1 U12009 ( .B1(n12729), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .A(
        n10032), .ZN(n12108) );
  AND2_X1 U12010 ( .A1(n10016), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n10032) );
  AOI21_X1 U12011 ( .B1(n12732), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .A(
        n10028), .ZN(n12061) );
  AND2_X1 U12012 ( .A1(n10016), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n10028) );
  AOI21_X1 U12013 ( .B1(n12286), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A(
        n10020), .ZN(n11718) );
  AND2_X1 U12014 ( .A1(n12723), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n10020) );
  NAND2_X1 U12015 ( .A1(n16302), .A2(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n10296) );
  OR2_X1 U12016 ( .A1(n11789), .A2(n11788), .ZN(n11864) );
  AOI21_X1 U12017 ( .B1(n11599), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A(
        n10017), .ZN(n11701) );
  AND2_X1 U12018 ( .A1(n9821), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n10017) );
  NAND2_X1 U12019 ( .A1(n9933), .A2(n10055), .ZN(n10054) );
  INV_X1 U12020 ( .A(n11846), .ZN(n10055) );
  NAND2_X1 U12021 ( .A1(n11651), .A2(n11979), .ZN(n11584) );
  AOI22_X1 U12022 ( .A1(n11766), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12722), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11566) );
  NAND2_X1 U12023 ( .A1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n13478), .ZN(
        n11963) );
  OR2_X1 U12024 ( .A1(n14601), .A2(n10505), .ZN(n10508) );
  AND2_X1 U12025 ( .A1(n10438), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10424) );
  NOR2_X1 U12026 ( .A1(n10438), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10426) );
  OR2_X1 U12027 ( .A1(n15752), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n10373) );
  AND4_X1 U12028 ( .A1(n11237), .A2(n11236), .A3(n11235), .A4(n11234), .ZN(
        n11249) );
  OR2_X1 U12029 ( .A1(n10542), .A2(n10541), .ZN(n11230) );
  AOI22_X1 U12030 ( .A1(n11022), .A2(P2_REIP_REG_3__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11007) );
  AND2_X1 U12031 ( .A1(n11021), .A2(P2_EBX_REG_3__SCAN_IN), .ZN(n11009) );
  AND2_X1 U12032 ( .A1(n10301), .A2(n9942), .ZN(n10076) );
  AOI21_X1 U12033 ( .B1(n11022), .B2(P2_REIP_REG_1__SCAN_IN), .A(n9935), .ZN(
        n10078) );
  OR2_X1 U12034 ( .A1(n10494), .A2(n10493), .ZN(n11375) );
  NAND2_X1 U12035 ( .A1(n11021), .A2(P2_EBX_REG_0__SCAN_IN), .ZN(n10989) );
  NAND2_X1 U12036 ( .A1(n10982), .A2(n10216), .ZN(n10214) );
  NOR2_X1 U12037 ( .A1(n11379), .A2(n14298), .ZN(n10216) );
  NAND2_X1 U12038 ( .A1(n10967), .A2(n10951), .ZN(n10970) );
  NAND2_X1 U12039 ( .A1(n17344), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n10124) );
  AND2_X1 U12040 ( .A1(n13461), .A2(n11644), .ZN(n12752) );
  AOI21_X1 U12041 ( .B1(n12286), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A(
        n10024), .ZN(n12118) );
  AND2_X1 U12042 ( .A1(n10016), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n10024) );
  OR2_X1 U12043 ( .A1(n10349), .A2(n14822), .ZN(n10348) );
  NAND2_X1 U12044 ( .A1(n10350), .A2(n12409), .ZN(n10349) );
  INV_X1 U12045 ( .A(n14834), .ZN(n10350) );
  AOI21_X1 U12046 ( .B1(n12286), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A(
        n10027), .ZN(n12231) );
  AOI21_X1 U12047 ( .B1(n12732), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .A(
        n10029), .ZN(n12197) );
  AND2_X1 U12048 ( .A1(n10016), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n10029) );
  INV_X1 U12049 ( .A(n12717), .ZN(n12744) );
  AOI21_X1 U12050 ( .B1(n9817), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .A(
        n10035), .ZN(n12187) );
  AOI21_X1 U12051 ( .B1(n12286), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .A(
        n10025), .ZN(n12131) );
  NAND2_X1 U12052 ( .A1(n9878), .A2(n9956), .ZN(n10342) );
  INV_X1 U12053 ( .A(n14249), .ZN(n10330) );
  XNOR2_X1 U12054 ( .A(n11885), .B(n11884), .ZN(n12037) );
  NAND2_X1 U12055 ( .A1(n11665), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12143) );
  INV_X1 U12056 ( .A(n12143), .ZN(n12154) );
  NAND2_X1 U12057 ( .A1(n10014), .A2(n9986), .ZN(n13003) );
  AOI21_X1 U12058 ( .B1(n10293), .B2(n10298), .A(n10292), .ZN(n10291) );
  INV_X1 U12059 ( .A(n15214), .ZN(n10292) );
  NAND2_X1 U12060 ( .A1(n10287), .A2(n11872), .ZN(n10286) );
  OR2_X1 U12061 ( .A1(n11813), .A2(n11812), .ZN(n11888) );
  OAI22_X1 U12062 ( .A1(n11598), .A2(n12848), .B1(n13775), .B2(n13762), .ZN(
        n11668) );
  AND2_X1 U12063 ( .A1(n11707), .A2(n11706), .ZN(n11731) );
  INV_X1 U12064 ( .A(n11819), .ZN(n9984) );
  CLKBUF_X1 U12065 ( .A(n13461), .Z(n13462) );
  NAND2_X1 U12066 ( .A1(n20597), .A2(n20310), .ZN(n11778) );
  NAND2_X1 U12067 ( .A1(n9821), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n11604) );
  NAND2_X1 U12068 ( .A1(n10039), .A2(n10038), .ZN(n10036) );
  AND2_X1 U12069 ( .A1(n11765), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11939) );
  NOR2_X1 U12070 ( .A1(n11959), .A2(n11929), .ZN(n11962) );
  AND2_X1 U12071 ( .A1(n11928), .A2(n11963), .ZN(n12758) );
  OR2_X1 U12072 ( .A1(n11964), .A2(n11927), .ZN(n11928) );
  AND2_X1 U12073 ( .A1(n20302), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n11927) );
  AOI21_X1 U12074 ( .B1(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n20017), .A(
        n10494), .ZN(n10588) );
  NOR2_X1 U12075 ( .A1(n12448), .A2(n10185), .ZN(n10184) );
  INV_X1 U12076 ( .A(n11329), .ZN(n10186) );
  AND2_X1 U12077 ( .A1(n10543), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n11325) );
  NAND2_X1 U12078 ( .A1(n11318), .A2(n10187), .ZN(n11330) );
  NAND2_X1 U12079 ( .A1(n11318), .A2(n11319), .ZN(n11326) );
  NOR2_X1 U12080 ( .A1(n15542), .A2(n10260), .ZN(n10259) );
  INV_X1 U12081 ( .A(n15556), .ZN(n10260) );
  INV_X1 U12082 ( .A(n15602), .ZN(n10897) );
  NAND2_X1 U12083 ( .A1(n10280), .A2(n14241), .ZN(n10279) );
  AND2_X1 U12084 ( .A1(n14206), .A2(n10281), .ZN(n10280) );
  INV_X1 U12085 ( .A(n14255), .ZN(n10281) );
  AND2_X1 U12086 ( .A1(n10358), .A2(n10563), .ZN(n11250) );
  AND2_X1 U12087 ( .A1(n14723), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n13589) );
  NAND2_X1 U12088 ( .A1(n10657), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11384) );
  AND2_X1 U12089 ( .A1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n10138) );
  INV_X1 U12090 ( .A(n13601), .ZN(n10145) );
  XNOR2_X1 U12091 ( .A(n10993), .B(n10994), .ZN(n11149) );
  NOR2_X1 U12092 ( .A1(n10226), .A2(n10222), .ZN(n11429) );
  NAND2_X1 U12093 ( .A1(n10670), .A2(n10669), .ZN(n10226) );
  INV_X1 U12094 ( .A(n12481), .ZN(n10173) );
  NAND2_X1 U12095 ( .A1(n10174), .A2(n9870), .ZN(n10171) );
  AND2_X1 U12096 ( .A1(n15895), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n10307) );
  NOR2_X1 U12097 ( .A1(n15773), .A2(n10327), .ZN(n10326) );
  INV_X1 U12098 ( .A(n15780), .ZN(n10327) );
  OR2_X1 U12099 ( .A1(n15530), .A2(n11254), .ZN(n12478) );
  NAND2_X1 U12100 ( .A1(n10376), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n10305) );
  AND2_X1 U12101 ( .A1(n11335), .A2(n10245), .ZN(n10244) );
  INV_X1 U12102 ( .A(n16023), .ZN(n10245) );
  INV_X1 U12103 ( .A(n16038), .ZN(n10246) );
  OR2_X1 U12104 ( .A1(n11290), .A2(n11283), .ZN(n11282) );
  AND2_X1 U12105 ( .A1(n9929), .A2(n11439), .ZN(n10080) );
  XNOR2_X1 U12106 ( .A(n11290), .B(n11291), .ZN(n11446) );
  NOR2_X1 U12107 ( .A1(n11446), .A2(n14270), .ZN(n11449) );
  NAND2_X1 U12108 ( .A1(n11011), .A2(n11010), .ZN(n11016) );
  NOR2_X1 U12109 ( .A1(n11009), .A2(n11008), .ZN(n11010) );
  NAND2_X1 U12110 ( .A1(n11053), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11011) );
  INV_X1 U12111 ( .A(n11007), .ZN(n11008) );
  INV_X1 U12112 ( .A(n11155), .ZN(n10264) );
  NAND2_X1 U12113 ( .A1(n11141), .A2(n11139), .ZN(n10267) );
  NAND2_X1 U12114 ( .A1(n10073), .A2(n11138), .ZN(n10266) );
  NAND2_X1 U12115 ( .A1(n11185), .A2(n11184), .ZN(n10213) );
  NAND2_X1 U12116 ( .A1(n11206), .A2(n11205), .ZN(n10212) );
  INV_X1 U12117 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n11499) );
  NAND2_X1 U12118 ( .A1(n13590), .A2(n20013), .ZN(n13582) );
  NAND2_X1 U12119 ( .A1(n14723), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n13570) );
  NAND2_X1 U12120 ( .A1(n11177), .A2(n9860), .ZN(n19572) );
  AOI21_X1 U12121 ( .B1(n10645), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A(
        n10632), .ZN(n10637) );
  NAND2_X1 U12122 ( .A1(n10645), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n10598) );
  NOR2_X1 U12123 ( .A1(n19610), .A2(n20028), .ZN(n14304) );
  NOR2_X1 U12124 ( .A1(n13250), .A2(n12593), .ZN(n13183) );
  NOR2_X1 U12125 ( .A1(n12508), .A2(n12514), .ZN(n13082) );
  NAND2_X1 U12126 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n18982), .ZN(
        n12513) );
  INV_X1 U12127 ( .A(n17099), .ZN(n12509) );
  AND2_X1 U12128 ( .A1(n17920), .A2(n18258), .ZN(n10168) );
  OR2_X1 U12129 ( .A1(n13181), .A2(n18378), .ZN(n10002) );
  NOR3_X1 U12130 ( .A1(n10004), .A2(n13178), .A3(n13177), .ZN(n10003) );
  NOR2_X1 U12131 ( .A1(n12581), .A2(n10012), .ZN(n10011) );
  NOR2_X1 U12132 ( .A1(n13051), .A2(n17201), .ZN(n10012) );
  NAND2_X1 U12133 ( .A1(n17379), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n10010) );
  AOI21_X1 U12134 ( .B1(n18367), .B2(n19016), .A(n18988), .ZN(n18377) );
  NAND2_X1 U12135 ( .A1(n13172), .A2(n18816), .ZN(n16149) );
  INV_X1 U12136 ( .A(n12938), .ZN(n16194) );
  CLKBUF_X1 U12137 ( .A(n12752), .Z(n12753) );
  INV_X1 U12138 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n14951) );
  AND2_X1 U12139 ( .A1(n16264), .A2(n14956), .ZN(n16237) );
  INV_X1 U12140 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n20104) );
  OR2_X1 U12141 ( .A1(n12054), .A2(n14392), .ZN(n12079) );
  AND2_X1 U12142 ( .A1(n12926), .A2(n12925), .ZN(n14845) );
  NAND2_X1 U12143 ( .A1(n13631), .A2(n13548), .ZN(n10197) );
  NAND2_X1 U12144 ( .A1(n13549), .A2(n13548), .ZN(n13551) );
  XNOR2_X1 U12145 ( .A(n10198), .B(n13631), .ZN(n13549) );
  OAI21_X1 U12146 ( .B1(n12938), .B2(n12765), .A(n12764), .ZN(n13460) );
  OR2_X1 U12147 ( .A1(n13792), .A2(n16210), .ZN(n12764) );
  NAND2_X1 U12148 ( .A1(n15090), .A2(n10042), .ZN(n14002) );
  NAND2_X1 U12149 ( .A1(n10347), .A2(n13015), .ZN(n10346) );
  INV_X1 U12150 ( .A(n10348), .ZN(n10347) );
  NAND2_X1 U12151 ( .A1(n12370), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n12697) );
  NOR2_X1 U12152 ( .A1(n12327), .A2(n15167), .ZN(n12328) );
  OR2_X1 U12153 ( .A1(n15160), .A2(n12742), .ZN(n12349) );
  CLKBUF_X1 U12154 ( .A(n14858), .Z(n14859) );
  OR2_X1 U12155 ( .A1(n12281), .A2(n15185), .ZN(n12319) );
  NOR2_X1 U12156 ( .A1(n12246), .A2(n15202), .ZN(n12247) );
  AND2_X1 U12157 ( .A1(n12265), .A2(n12264), .ZN(n14914) );
  AND2_X1 U12158 ( .A1(n12210), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n12211) );
  NOR2_X1 U12159 ( .A1(n15005), .A2(n10345), .ZN(n10343) );
  NAND2_X1 U12160 ( .A1(n12180), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12194) );
  NAND2_X1 U12161 ( .A1(n12145), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12162) );
  CLKBUF_X1 U12162 ( .A(n15023), .Z(n15024) );
  INV_X1 U12163 ( .A(n12127), .ZN(n12102) );
  AND2_X1 U12164 ( .A1(n12083), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n12084) );
  NAND2_X1 U12165 ( .A1(n12084), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n12127) );
  NAND2_X1 U12166 ( .A1(n12032), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12054) );
  NOR2_X1 U12167 ( .A1(n12019), .A2(n21092), .ZN(n12026) );
  INV_X1 U12168 ( .A(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n21092) );
  AND2_X1 U12169 ( .A1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n12000), .ZN(
        n12010) );
  AOI21_X1 U12170 ( .B1(n11983), .B2(n12143), .A(n10335), .ZN(n10334) );
  INV_X1 U12171 ( .A(n11999), .ZN(n10335) );
  NAND2_X1 U12172 ( .A1(n13971), .A2(n11983), .ZN(n10336) );
  NAND2_X1 U12173 ( .A1(n13542), .A2(n13541), .ZN(n13729) );
  NOR3_X1 U12174 ( .A1(n14861), .A2(n14837), .A3(n14845), .ZN(n14835) );
  NOR2_X1 U12175 ( .A1(n14861), .A2(n14845), .ZN(n14846) );
  NAND2_X1 U12176 ( .A1(n15146), .A2(n13003), .ZN(n15137) );
  NAND2_X1 U12177 ( .A1(n13002), .A2(n15344), .ZN(n10014) );
  NAND2_X1 U12178 ( .A1(n15009), .A2(n9955), .ZN(n14903) );
  INV_X1 U12179 ( .A(n14905), .ZN(n10194) );
  AOI21_X1 U12180 ( .B1(n15191), .B2(n11910), .A(n9844), .ZN(n15182) );
  NAND2_X1 U12181 ( .A1(n15009), .A2(n10195), .ZN(n14919) );
  NAND2_X1 U12182 ( .A1(n15009), .A2(n14934), .ZN(n14933) );
  INV_X1 U12183 ( .A(n15013), .ZN(n10206) );
  INV_X1 U12184 ( .A(n10204), .ZN(n10203) );
  NAND2_X1 U12185 ( .A1(n10048), .A2(n10045), .ZN(n16300) );
  NOR2_X1 U12186 ( .A1(n10047), .A2(n10046), .ZN(n10045) );
  INV_X1 U12187 ( .A(n15226), .ZN(n10046) );
  AND2_X1 U12188 ( .A1(n12903), .A2(n12902), .ZN(n14965) );
  NOR3_X1 U12189 ( .A1(n15039), .A2(n10207), .A3(n14985), .ZN(n14966) );
  OR2_X1 U12190 ( .A1(n15044), .A2(n15037), .ZN(n15039) );
  NOR2_X1 U12191 ( .A1(n15039), .A2(n14985), .ZN(n15030) );
  AND2_X1 U12192 ( .A1(n12883), .A2(n12882), .ZN(n15042) );
  AND2_X1 U12193 ( .A1(n16410), .A2(n12879), .ZN(n15040) );
  AND2_X1 U12194 ( .A1(n11817), .A2(n11886), .ZN(n11818) );
  NOR2_X1 U12195 ( .A1(n16408), .A2(n16407), .ZN(n16410) );
  NOR2_X1 U12196 ( .A1(n10192), .A2(n16422), .ZN(n10191) );
  INV_X1 U12197 ( .A(n14044), .ZN(n10192) );
  OR2_X1 U12198 ( .A1(n16424), .A2(n14259), .ZN(n16408) );
  NOR2_X1 U12199 ( .A1(n13858), .A2(n13859), .ZN(n14045) );
  NAND2_X1 U12200 ( .A1(n14045), .A2(n14044), .ZN(n10193) );
  OR2_X1 U12201 ( .A1(n13754), .A2(n13753), .ZN(n13858) );
  INV_X1 U12202 ( .A(n15284), .ZN(n20277) );
  INV_X1 U12203 ( .A(n13521), .ZN(n15466) );
  CLKBUF_X1 U12204 ( .A(n13473), .Z(n13474) );
  OR2_X1 U12205 ( .A1(n9853), .A2(n11991), .ZN(n20631) );
  INV_X1 U12206 ( .A(n20350), .ZN(n20341) );
  OR2_X1 U12207 ( .A1(n20704), .A2(n20631), .ZN(n20653) );
  NAND2_X1 U12208 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20696) );
  OR2_X1 U12209 ( .A1(n20594), .A2(n11822), .ZN(n20704) );
  OR2_X1 U12210 ( .A1(n9853), .A2(n20307), .ZN(n20725) );
  NOR2_X2 U12211 ( .A1(n20306), .A2(n20305), .ZN(n20345) );
  NAND3_X1 U12212 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n20310), .A3(n20309), 
        .ZN(n20350) );
  NAND2_X1 U12213 ( .A1(n11372), .A2(n11379), .ZN(n13380) );
  NOR2_X1 U12214 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n14129) );
  OR2_X1 U12215 ( .A1(n11480), .A2(n11479), .ZN(n14105) );
  AOI221_X1 U12216 ( .B1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(n10588), 
        .C1(n11383), .C2(n10588), .A(n10587), .ZN(n11402) );
  NOR2_X1 U12217 ( .A1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n16228), .ZN(
        n10587) );
  NAND2_X1 U12218 ( .A1(n9889), .A2(n12460), .ZN(n12804) );
  AND2_X1 U12219 ( .A1(n10543), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n12471) );
  AND2_X1 U12220 ( .A1(n11135), .A2(n9953), .ZN(n12457) );
  NAND2_X1 U12221 ( .A1(n15561), .A2(n16484), .ZN(n10133) );
  OR2_X1 U12222 ( .A1(n10415), .A2(n10134), .ZN(n15561) );
  NOR2_X1 U12223 ( .A1(n15585), .A2(n15805), .ZN(n10134) );
  AND2_X1 U12224 ( .A1(n9875), .A2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n10139) );
  NAND2_X1 U12225 ( .A1(n10517), .A2(n10516), .ZN(n11266) );
  NAND2_X1 U12226 ( .A1(n11400), .A2(n10960), .ZN(n10517) );
  INV_X1 U12227 ( .A(n19180), .ZN(n19166) );
  AND2_X1 U12228 ( .A1(n15553), .A2(n15554), .ZN(n15537) );
  NAND2_X1 U12229 ( .A1(n13702), .A2(n10268), .ZN(n13813) );
  AND2_X1 U12230 ( .A1(n13701), .A2(n13705), .ZN(n10268) );
  NAND2_X1 U12231 ( .A1(n13569), .A2(n13589), .ZN(n13620) );
  NAND2_X1 U12232 ( .A1(n15572), .A2(n9957), .ZN(n15717) );
  AND2_X1 U12233 ( .A1(n15572), .A2(n9952), .ZN(n15719) );
  XNOR2_X1 U12234 ( .A(n14686), .B(n14682), .ZN(n15652) );
  NAND2_X1 U12235 ( .A1(n15572), .A2(n10259), .ZN(n15544) );
  NAND2_X1 U12236 ( .A1(n15572), .A2(n15556), .ZN(n15541) );
  XNOR2_X1 U12237 ( .A(n14642), .B(n14665), .ZN(n15665) );
  AND2_X1 U12238 ( .A1(n10898), .A2(n9958), .ZN(n15569) );
  INV_X1 U12239 ( .A(n14242), .ZN(n10898) );
  AND2_X1 U12240 ( .A1(n10900), .A2(n10899), .ZN(n14381) );
  NAND2_X1 U12241 ( .A1(n10898), .A2(n10897), .ZN(n15604) );
  OR2_X1 U12242 ( .A1(n10722), .A2(n10234), .ZN(n14415) );
  INV_X1 U12243 ( .A(n19420), .ZN(n10937) );
  INV_X1 U12244 ( .A(n13285), .ZN(n14302) );
  NAND2_X1 U12245 ( .A1(n10393), .A2(n9881), .ZN(n10387) );
  NAND2_X1 U12246 ( .A1(n10393), .A2(n10142), .ZN(n10390) );
  NAND2_X1 U12247 ( .A1(n10393), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n10392) );
  AND2_X1 U12248 ( .A1(n11082), .A2(n11081), .ZN(n15688) );
  NAND2_X1 U12249 ( .A1(n10400), .A2(n9875), .ZN(n10413) );
  INV_X1 U12250 ( .A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n15845) );
  NAND2_X1 U12251 ( .A1(n10400), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n10412) );
  AND2_X1 U12252 ( .A1(n10404), .A2(n9873), .ZN(n10411) );
  AND3_X1 U12253 ( .A1(n11064), .A2(n11063), .A3(n11062), .ZN(n14028) );
  AND3_X1 U12254 ( .A1(n11060), .A2(n11059), .A3(n11058), .ZN(n13997) );
  NAND2_X1 U12255 ( .A1(n10404), .A2(n9866), .ZN(n10410) );
  NAND2_X1 U12256 ( .A1(n13662), .A2(n13819), .ZN(n13818) );
  NOR2_X1 U12257 ( .A1(n14424), .A2(n10137), .ZN(n10136) );
  INV_X1 U12258 ( .A(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n10137) );
  NAND2_X1 U12259 ( .A1(n10407), .A2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10406) );
  INV_X1 U12260 ( .A(n10154), .ZN(n12489) );
  NAND2_X1 U12261 ( .A1(n12801), .A2(n12800), .ZN(n12975) );
  NOR2_X1 U12262 ( .A1(n13315), .A2(n11254), .ZN(n15752) );
  NOR2_X1 U12263 ( .A1(n12472), .A2(n11254), .ZN(n15753) );
  AOI21_X1 U12264 ( .B1(n15782), .B2(n10326), .A(n15749), .ZN(n15750) );
  INV_X1 U12265 ( .A(n12422), .ZN(n15763) );
  AND2_X1 U12266 ( .A1(n11107), .A2(n11106), .ZN(n15642) );
  AND2_X1 U12267 ( .A1(n11103), .A2(n11102), .ZN(n15522) );
  NAND2_X1 U12268 ( .A1(n15553), .A2(n9951), .ZN(n15540) );
  OR2_X1 U12269 ( .A1(n15955), .A2(n12484), .ZN(n15910) );
  OR2_X1 U12270 ( .A1(n12478), .A2(n15912), .ZN(n15781) );
  XNOR2_X1 U12271 ( .A(n12451), .B(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15936) );
  AND3_X1 U12272 ( .A1(n11092), .A2(n11091), .A3(n11090), .ZN(n15566) );
  NOR2_X1 U12273 ( .A1(n12441), .A2(n10317), .ZN(n10316) );
  INV_X1 U12274 ( .A(n11323), .ZN(n10317) );
  NOR2_X1 U12275 ( .A1(n15828), .A2(n11358), .ZN(n15816) );
  INV_X1 U12276 ( .A(n15834), .ZN(n10304) );
  OR2_X1 U12277 ( .A1(n11512), .A2(n16052), .ZN(n15976) );
  AND2_X1 U12278 ( .A1(n11079), .A2(n11078), .ZN(n14431) );
  AND3_X1 U12279 ( .A1(n11075), .A2(n11074), .A3(n11073), .ZN(n14403) );
  AOI21_X1 U12280 ( .B1(n10237), .B2(n10241), .A(n9934), .ZN(n10236) );
  AND2_X1 U12281 ( .A1(n14442), .A2(n14443), .ZN(n14445) );
  NAND2_X1 U12282 ( .A1(n16041), .A2(n10244), .ZN(n10242) );
  NAND2_X1 U12283 ( .A1(n10246), .A2(n10245), .ZN(n10243) );
  AOI21_X1 U12284 ( .B1(n16041), .B2(n11335), .A(n10246), .ZN(n16022) );
  NOR2_X1 U12285 ( .A1(n11461), .A2(n11476), .ZN(n10084) );
  AOI21_X1 U12286 ( .B1(n10068), .B2(n10319), .A(n10066), .ZN(n10065) );
  AND2_X1 U12287 ( .A1(n9868), .A2(n10322), .ZN(n10066) );
  NOR2_X1 U12288 ( .A1(n10068), .A2(n9868), .ZN(n10067) );
  INV_X1 U12289 ( .A(n13812), .ZN(n10149) );
  AND3_X1 U12290 ( .A1(n10827), .A2(n10826), .A3(n10825), .ZN(n15620) );
  INV_X1 U12291 ( .A(n14532), .ZN(n10233) );
  NAND2_X1 U12292 ( .A1(n10087), .A2(n10083), .ZN(n10082) );
  NOR2_X1 U12293 ( .A1(n16538), .A2(n10089), .ZN(n10083) );
  INV_X1 U12294 ( .A(n14410), .ZN(n10324) );
  INV_X1 U12295 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n16573) );
  NOR2_X1 U12296 ( .A1(n13915), .A2(n10250), .ZN(n14272) );
  NAND2_X1 U12297 ( .A1(n10249), .A2(n10248), .ZN(n10250) );
  AND2_X1 U12298 ( .A1(n10251), .A2(n13874), .ZN(n10248) );
  INV_X1 U12299 ( .A(n14037), .ZN(n10251) );
  INV_X1 U12300 ( .A(n11442), .ZN(n11443) );
  XNOR2_X1 U12301 ( .A(n13366), .B(n10693), .ZN(n13453) );
  NAND2_X1 U12302 ( .A1(n10249), .A2(n13874), .ZN(n10252) );
  NAND2_X1 U12303 ( .A1(n13588), .A2(n13620), .ZN(n13621) );
  INV_X1 U12304 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n16105) );
  NAND2_X1 U12305 ( .A1(n10971), .A2(n20064), .ZN(n11372) );
  AND2_X1 U12306 ( .A1(n10680), .A2(n10936), .ZN(n10954) );
  NAND2_X1 U12307 ( .A1(n19431), .A2(n20040), .ZN(n19615) );
  OR2_X1 U12308 ( .A1(n19782), .A2(n19781), .ZN(n19803) );
  NAND2_X1 U12309 ( .A1(n10608), .A2(n10607), .ZN(n10615) );
  NAND2_X1 U12310 ( .A1(n14304), .A2(n14303), .ZN(n19422) );
  INV_X1 U12311 ( .A(n19412), .ZN(n19419) );
  NOR2_X1 U12312 ( .A1(n20034), .A2(n13362), .ZN(n13694) );
  NOR2_X1 U12313 ( .A1(n13183), .A2(n13195), .ZN(n13172) );
  INV_X1 U12314 ( .A(n18405), .ZN(n13176) );
  NOR2_X1 U12315 ( .A1(n16776), .A2(n16775), .ZN(n16774) );
  NOR2_X1 U12316 ( .A1(n16795), .A2(n16794), .ZN(n16793) );
  INV_X1 U12317 ( .A(n17083), .ZN(n17104) );
  NAND2_X1 U12318 ( .A1(n19030), .A2(n18378), .ZN(n13305) );
  NAND2_X1 U12319 ( .A1(n17215), .A2(P3_EBX_REG_20__SCAN_IN), .ZN(n17198) );
  NOR2_X1 U12320 ( .A1(n17322), .A2(n10119), .ZN(n10118) );
  INV_X1 U12321 ( .A(P3_EBX_REG_10__SCAN_IN), .ZN(n10119) );
  INV_X1 U12322 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n17022) );
  INV_X1 U12323 ( .A(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n17217) );
  INV_X1 U12324 ( .A(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n21152) );
  INV_X1 U12325 ( .A(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n17211) );
  OR3_X1 U12326 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n18840), .ZN(n17306) );
  INV_X1 U12327 ( .A(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n17359) );
  INV_X1 U12328 ( .A(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n21237) );
  INV_X1 U12329 ( .A(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n21277) );
  NOR2_X1 U12330 ( .A1(n13088), .A2(n9975), .ZN(n13095) );
  NOR2_X1 U12331 ( .A1(n13093), .A2(n13092), .ZN(n13094) );
  AND2_X1 U12332 ( .A1(n12549), .A2(n12548), .ZN(n16232) );
  NOR2_X1 U12333 ( .A1(n17395), .A2(n13127), .ZN(n12546) );
  NAND2_X1 U12334 ( .A1(n16152), .A2(n9999), .ZN(n16229) );
  OR2_X1 U12335 ( .A1(n16732), .A2(n19012), .ZN(n9999) );
  AOI21_X1 U12336 ( .B1(n16146), .B2(n18857), .A(n19011), .ZN(n17582) );
  INV_X1 U12337 ( .A(n16732), .ZN(n17632) );
  AND2_X1 U12338 ( .A1(n17722), .A2(n9880), .ZN(n16614) );
  NAND2_X1 U12339 ( .A1(n17722), .A2(n9874), .ZN(n13235) );
  NOR2_X1 U12340 ( .A1(n17703), .A2(n10098), .ZN(n10097) );
  NAND2_X1 U12341 ( .A1(n17722), .A2(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n17702) );
  NOR2_X1 U12342 ( .A1(n17736), .A2(n17737), .ZN(n17722) );
  NOR2_X1 U12343 ( .A1(n10115), .A2(n10112), .ZN(n10111) );
  INV_X1 U12344 ( .A(n10113), .ZN(n10112) );
  NAND2_X1 U12345 ( .A1(n17882), .A2(n10111), .ZN(n17785) );
  NAND2_X1 U12346 ( .A1(n17882), .A2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n17856) );
  NOR2_X1 U12347 ( .A1(n17900), .A2(n17902), .ZN(n17882) );
  AOI21_X1 U12348 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n17806), .A(
        n18748), .ZN(n17901) );
  NAND2_X1 U12349 ( .A1(n16994), .A2(n9931), .ZN(n17921) );
  INV_X1 U12350 ( .A(n16994), .ZN(n17945) );
  NOR2_X1 U12351 ( .A1(n17971), .A2(n17989), .ZN(n17954) );
  NAND2_X1 U12352 ( .A1(n17996), .A2(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n9969) );
  NAND2_X1 U12353 ( .A1(n17995), .A2(n9971), .ZN(n9970) );
  OR2_X1 U12354 ( .A1(n17996), .A2(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n9971) );
  NAND2_X1 U12355 ( .A1(n18003), .A2(n13219), .ZN(n17991) );
  NAND2_X1 U12356 ( .A1(n17991), .A2(n17992), .ZN(n17990) );
  INV_X1 U12357 ( .A(n18007), .ZN(n17052) );
  AND2_X1 U12358 ( .A1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n18007) );
  AOI21_X1 U12359 ( .B1(n16217), .B2(n17957), .A(n16603), .ZN(n13166) );
  NAND2_X1 U12360 ( .A1(n16165), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16217) );
  AND2_X1 U12361 ( .A1(n16623), .A2(n9972), .ZN(n16165) );
  NOR2_X1 U12362 ( .A1(n13160), .A2(n17693), .ZN(n9972) );
  NOR2_X1 U12363 ( .A1(n13159), .A2(n17811), .ZN(n17757) );
  NAND2_X1 U12364 ( .A1(n17757), .A2(n18098), .ZN(n17756) );
  INV_X1 U12365 ( .A(n13161), .ZN(n17811) );
  INV_X1 U12366 ( .A(n17853), .ZN(n16637) );
  NAND2_X1 U12367 ( .A1(n10167), .A2(n10168), .ZN(n17910) );
  INV_X1 U12368 ( .A(n17933), .ZN(n10167) );
  NAND2_X1 U12369 ( .A1(n13186), .A2(n13184), .ZN(n13289) );
  NOR2_X1 U12370 ( .A1(n13199), .A2(n17957), .ZN(n17942) );
  XNOR2_X1 U12371 ( .A(n13148), .B(n13147), .ZN(n17970) );
  INV_X1 U12372 ( .A(n13149), .ZN(n13147) );
  XNOR2_X1 U12373 ( .A(n13217), .B(n9978), .ZN(n18004) );
  INV_X1 U12374 ( .A(n13218), .ZN(n9978) );
  NAND2_X1 U12375 ( .A1(n18004), .A2(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n18003) );
  INV_X1 U12376 ( .A(n18831), .ZN(n18807) );
  XNOR2_X1 U12377 ( .A(n13135), .B(n13118), .ZN(n18029) );
  AOI211_X1 U12378 ( .C1(n12616), .C2(n12615), .A(n13188), .B(n12614), .ZN(
        n18808) );
  NOR2_X1 U12379 ( .A1(n13130), .A2(n13129), .ZN(n13131) );
  NOR2_X2 U12380 ( .A1(n19029), .A2(n16149), .ZN(n18831) );
  NAND2_X1 U12381 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n18840) );
  AND2_X1 U12382 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n18838) );
  INV_X1 U12383 ( .A(n16232), .ZN(n18378) );
  OAI211_X1 U12384 ( .C1(n12537), .C2(n21140), .A(n12603), .B(n12602), .ZN(
        n18397) );
  AOI211_X1 U12385 ( .C1(n17344), .C2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A(
        n12601), .B(n12600), .ZN(n12602) );
  NOR2_X1 U12386 ( .A1(n12564), .A2(n12563), .ZN(n12565) );
  AND2_X1 U12387 ( .A1(n17357), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n12563) );
  INV_X1 U12388 ( .A(n12571), .ZN(n10120) );
  INV_X1 U12389 ( .A(n18720), .ZN(n18415) );
  INV_X1 U12390 ( .A(n18864), .ZN(n19020) );
  OR2_X1 U12391 ( .A1(n20910), .A2(n20310), .ZN(n20086) );
  NAND2_X1 U12392 ( .A1(READY11_REG_SCAN_IN), .A2(READY1), .ZN(n21010) );
  INV_X1 U12393 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n16258) );
  OR2_X1 U12394 ( .A1(n16280), .A2(n14957), .ZN(n16260) );
  NAND2_X1 U12395 ( .A1(n20117), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20158) );
  NAND2_X1 U12396 ( .A1(n12955), .A2(n12953), .ZN(n20151) );
  INV_X1 U12397 ( .A(n14988), .ZN(n20131) );
  INV_X1 U12398 ( .A(n20124), .ZN(n20149) );
  NAND2_X1 U12399 ( .A1(n12955), .A2(n12954), .ZN(n20122) );
  INV_X1 U12400 ( .A(n20158), .ZN(n20140) );
  AND2_X1 U12401 ( .A1(n20182), .A2(n11979), .ZN(n20178) );
  INV_X1 U12402 ( .A(n20182), .ZN(n15032) );
  AND2_X1 U12403 ( .A1(n20182), .A2(n20349), .ZN(n20171) );
  AND2_X2 U12404 ( .A1(n13547), .A2(n13768), .ZN(n20182) );
  INV_X1 U12405 ( .A(n20171), .ZN(n20175) );
  NAND2_X1 U12406 ( .A1(n15090), .A2(n13020), .ZN(n15091) );
  INV_X1 U12407 ( .A(n15103), .ZN(n16295) );
  INV_X1 U12408 ( .A(n16299), .ZN(n15105) );
  AND2_X1 U12409 ( .A1(n15091), .A2(n14002), .ZN(n15116) );
  AND2_X1 U12410 ( .A1(n13639), .A2(n13638), .ZN(n20187) );
  OAI22_X1 U12411 ( .A1(n13637), .A2(n16201), .B1(n15468), .B2(n13636), .ZN(
        n13639) );
  INV_X2 U12412 ( .A(n13808), .ZN(n20238) );
  OR2_X1 U12413 ( .A1(n12845), .A2(n15124), .ZN(n12846) );
  INV_X1 U12414 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n15202) );
  NAND2_X1 U12415 ( .A1(n9833), .A2(n11861), .ZN(n16342) );
  INV_X1 U12416 ( .A(n20248), .ZN(n20088) );
  INV_X1 U12417 ( .A(n20252), .ZN(n16316) );
  INV_X1 U12418 ( .A(n15228), .ZN(n20242) );
  XNOR2_X1 U12419 ( .A(n12937), .B(n12936), .ZN(n15274) );
  XNOR2_X1 U12420 ( .A(n13009), .B(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n15303) );
  NAND2_X1 U12421 ( .A1(n13008), .A2(n13007), .ZN(n13009) );
  OR2_X1 U12422 ( .A1(n14819), .A2(n14818), .ZN(n15322) );
  AND2_X1 U12423 ( .A1(n15367), .A2(n15292), .ZN(n15356) );
  OAI21_X1 U12424 ( .B1(n9833), .B2(n10287), .A(n10283), .ZN(n16337) );
  AOI21_X1 U12425 ( .B1(n16341), .B2(n10289), .A(n10288), .ZN(n10283) );
  NOR2_X1 U12426 ( .A1(n16399), .A2(n20258), .ZN(n16431) );
  AND2_X1 U12427 ( .A1(n13795), .A2(n13794), .ZN(n20278) );
  NAND2_X1 U12428 ( .A1(n13795), .A2(n16175), .ZN(n20298) );
  AND2_X1 U12429 ( .A1(n13795), .A2(n13779), .ZN(n20288) );
  INV_X1 U12430 ( .A(n20256), .ZN(n20296) );
  AND2_X1 U12431 ( .A1(n13795), .A2(n13770), .ZN(n20289) );
  INV_X1 U12432 ( .A(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n20302) );
  OAI21_X1 U12433 ( .B1(n13965), .B2(n16443), .A(n20469), .ZN(n20301) );
  INV_X1 U12434 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13523) );
  INV_X1 U12435 ( .A(n15468), .ZN(n16175) );
  NOR2_X1 U12436 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n20080) );
  NAND2_X1 U12437 ( .A1(n16193), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n15481) );
  OAI211_X1 U12438 ( .C1(n20461), .C2(n20999), .A(n20663), .B(n20315), .ZN(
        n20355) );
  OAI221_X1 U12439 ( .B1(n20488), .B2(n20738), .C1(n20488), .C2(n20470), .A(
        n20803), .ZN(n20491) );
  INV_X1 U12440 ( .A(n20560), .ZN(n20515) );
  OAI211_X1 U12441 ( .C1(n10375), .C2(n20738), .A(n20663), .B(n20605), .ZN(
        n20622) );
  INV_X1 U12442 ( .A(n20586), .ZN(n20621) );
  INV_X1 U12443 ( .A(n20653), .ZN(n20689) );
  OAI211_X1 U12444 ( .C1(n10377), .C2(n20738), .A(n20803), .B(n20737), .ZN(
        n20761) );
  NOR2_X2 U12445 ( .A1(n20704), .A2(n20703), .ZN(n20760) );
  OAI21_X1 U12446 ( .B1(n20773), .B2(n20772), .A(n20856), .ZN(n20791) );
  OAI211_X1 U12447 ( .C1(n20834), .C2(n20804), .A(n20803), .B(n20802), .ZN(
        n20838) );
  INV_X1 U12448 ( .A(n20659), .ZN(n20853) );
  INV_X1 U12449 ( .A(n20744), .ZN(n20863) );
  INV_X1 U12450 ( .A(n20671), .ZN(n20869) );
  INV_X1 U12451 ( .A(n20675), .ZN(n20876) );
  INV_X1 U12452 ( .A(n20753), .ZN(n20881) );
  AND2_X1 U12453 ( .A1(n20353), .A2(n20338), .ZN(n20888) );
  AND2_X1 U12454 ( .A1(n20353), .A2(n20342), .ZN(n20894) );
  NOR2_X2 U12455 ( .A1(n20855), .A2(n20703), .ZN(n20904) );
  OAI21_X1 U12456 ( .B1(n20858), .B2(n20857), .A(n20856), .ZN(n20905) );
  AND2_X1 U12457 ( .A1(n20353), .A2(n20352), .ZN(n20902) );
  INV_X1 U12458 ( .A(n16193), .ZN(n16210) );
  INV_X1 U12459 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n16442) );
  NAND2_X1 U12460 ( .A1(n16442), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20910) );
  INV_X2 U12461 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n20999) );
  OR2_X1 U12462 ( .A1(n12492), .A2(n12491), .ZN(n15697) );
  INV_X1 U12463 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n15765) );
  INV_X1 U12464 ( .A(n10130), .ZN(n15531) );
  INV_X1 U12465 ( .A(n10133), .ZN(n15564) );
  NAND2_X1 U12466 ( .A1(n11349), .A2(n9876), .ZN(n11133) );
  INV_X1 U12467 ( .A(n19211), .ZN(n19180) );
  OR2_X1 U12468 ( .A1(n16074), .A2(n10255), .ZN(n16051) );
  INV_X1 U12469 ( .A(n19197), .ZN(n19179) );
  AND2_X1 U12470 ( .A1(n11126), .A2(n10658), .ZN(n19186) );
  OR2_X1 U12471 ( .A1(n14115), .A2(n13359), .ZN(n19208) );
  NOR2_X1 U12472 ( .A1(n19210), .A2(n20036), .ZN(n19211) );
  INV_X1 U12473 ( .A(n14205), .ZN(n14281) );
  NAND2_X1 U12474 ( .A1(n13689), .A2(n13677), .ZN(n13349) );
  INV_X1 U12475 ( .A(n19258), .ZN(n19270) );
  INV_X1 U12476 ( .A(n19229), .ZN(n19265) );
  OR2_X1 U12477 ( .A1(n13687), .A2(n13385), .ZN(n13387) );
  OR2_X1 U12478 ( .A1(n16107), .A2(n13356), .ZN(n19207) );
  NAND2_X1 U12479 ( .A1(n19274), .A2(n13391), .ZN(n19258) );
  INV_X1 U12480 ( .A(n19312), .ZN(n19303) );
  AND2_X1 U12481 ( .A1(n13361), .A2(n13360), .ZN(n19310) );
  OR2_X1 U12482 ( .A1(n19310), .A2(n20057), .ZN(n19312) );
  OAI21_X1 U12483 ( .B1(n9839), .B2(n20069), .A(n13422), .ZN(n13447) );
  NOR2_X2 U12484 ( .A1(n13421), .A2(n20062), .ZN(n13527) );
  INV_X1 U12485 ( .A(n13527), .ZN(n13657) );
  INV_X1 U12486 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n15788) );
  INV_X1 U12487 ( .A(n15666), .ZN(n16476) );
  OAI21_X1 U12488 ( .B1(n19325), .B2(n16484), .A(n16483), .ZN(n10093) );
  INV_X1 U12489 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n15808) );
  INV_X1 U12490 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n15862) );
  INV_X1 U12491 ( .A(n10089), .ZN(n10088) );
  INV_X1 U12492 ( .A(n16550), .ZN(n19325) );
  INV_X1 U12493 ( .A(n16559), .ZN(n19313) );
  NAND2_X1 U12494 ( .A1(n12829), .A2(n9892), .ZN(n12830) );
  NAND2_X1 U12495 ( .A1(n15624), .A2(n19341), .ZN(n12829) );
  NOR2_X1 U12496 ( .A1(n10365), .A2(n12827), .ZN(n12828) );
  AOI21_X1 U12497 ( .B1(n12993), .B2(n19347), .A(n12992), .ZN(n12994) );
  INV_X1 U12498 ( .A(n14786), .ZN(n12993) );
  NAND2_X1 U12499 ( .A1(n15948), .A2(n10094), .ZN(n16480) );
  NAND2_X1 U12500 ( .A1(n10095), .A2(n15938), .ZN(n10094) );
  NAND2_X1 U12501 ( .A1(n14410), .A2(n11313), .ZN(n10070) );
  AND2_X1 U12502 ( .A1(n16574), .A2(n11511), .ZN(n16047) );
  INV_X1 U12503 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n16072) );
  NOR2_X1 U12504 ( .A1(n16580), .A2(n14412), .ZN(n16073) );
  INV_X1 U12505 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n14421) );
  CLKBUF_X1 U12506 ( .A(n14478), .Z(n14479) );
  AND2_X1 U12507 ( .A1(n10229), .A2(n10227), .ZN(n14052) );
  INV_X1 U12508 ( .A(n10230), .ZN(n10227) );
  AND2_X1 U12509 ( .A1(n10147), .A2(n11019), .ZN(n13610) );
  NAND2_X1 U12510 ( .A1(n11259), .A2(n14068), .ZN(n13870) );
  AND2_X1 U12511 ( .A1(n19336), .A2(n19333), .ZN(n19353) );
  AND2_X1 U12512 ( .A1(n11505), .A2(n20050), .ZN(n19331) );
  INV_X1 U12513 ( .A(n19207), .ZN(n20040) );
  OR2_X1 U12514 ( .A1(n20002), .A2(n20061), .ZN(n20028) );
  INV_X1 U12515 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n16228) );
  INV_X1 U12517 ( .A(n11372), .ZN(n16156) );
  INV_X1 U12518 ( .A(n19468), .ZN(n19488) );
  OR2_X1 U12519 ( .A1(n19615), .A2(n20004), .ZN(n19530) );
  INV_X1 U12520 ( .A(n19530), .ZN(n19535) );
  OAI21_X1 U12521 ( .B1(n14322), .B2(n20002), .A(n14321), .ZN(n19534) );
  INV_X1 U12522 ( .A(n19561), .ZN(n19563) );
  OAI21_X1 U12523 ( .B1(n19546), .B2(n19545), .A(n19544), .ZN(n19564) );
  OAI21_X1 U12524 ( .B1(n19546), .B2(n19543), .A(n19542), .ZN(n19565) );
  INV_X1 U12525 ( .A(n19603), .ZN(n19583) );
  INV_X1 U12526 ( .A(n19587), .ZN(n19600) );
  NOR2_X1 U12527 ( .A1(n20001), .A2(n19568), .ZN(n19604) );
  OAI21_X1 U12528 ( .B1(n19643), .B2(n20036), .A(n19614), .ZN(n19631) );
  OR2_X1 U12529 ( .A1(n19802), .A2(n19667), .ZN(n19697) );
  OAI21_X1 U12530 ( .B1(n19675), .B2(n19674), .A(n19673), .ZN(n19693) );
  OAI21_X1 U12531 ( .B1(n19717), .B2(n19579), .A(n14305), .ZN(n19709) );
  INV_X1 U12532 ( .A(n14301), .ZN(n19714) );
  NOR2_X2 U12533 ( .A1(n19802), .A2(n20004), .ZN(n19737) );
  NOR2_X1 U12534 ( .A1(n19802), .A2(n19781), .ZN(n19760) );
  INV_X1 U12535 ( .A(n19769), .ZN(n19763) );
  INV_X1 U12536 ( .A(n19780), .ZN(n19798) );
  OAI22_X1 U12537 ( .A1(n19390), .A2(n19424), .B1(n19389), .B2(n19422), .ZN(
        n19826) );
  OAI22_X1 U12538 ( .A1(n19398), .A2(n19424), .B1(n19397), .B2(n19422), .ZN(
        n19830) );
  OAI22_X1 U12539 ( .A1(n19405), .A2(n19422), .B1(n19404), .B2(n19424), .ZN(
        n19834) );
  OAI22_X1 U12540 ( .A1(n19411), .A2(n19422), .B1(n19410), .B2(n19424), .ZN(
        n19838) );
  INV_X1 U12541 ( .A(n19912), .ZN(n19845) );
  INV_X1 U12542 ( .A(n19803), .ZN(n19844) );
  OAI22_X1 U12543 ( .A1(n20347), .A2(n19424), .B1(n19418), .B2(n19422), .ZN(
        n19843) );
  AND2_X1 U12544 ( .A1(n10657), .A2(n19419), .ZN(n19855) );
  AND2_X1 U12545 ( .A1(n20062), .A2(n19419), .ZN(n19867) );
  INV_X1 U12546 ( .A(n19821), .ZN(n19868) );
  INV_X1 U12547 ( .A(n19825), .ZN(n19874) );
  INV_X1 U12548 ( .A(n19826), .ZN(n19884) );
  INV_X1 U12549 ( .A(n19833), .ZN(n19886) );
  INV_X1 U12550 ( .A(n19837), .ZN(n19892) );
  INV_X1 U12551 ( .A(n19834), .ZN(n19896) );
  OR2_X1 U12552 ( .A1(n19802), .A2(n20001), .ZN(n19912) );
  INV_X1 U12553 ( .A(n19370), .ZN(n19908) );
  AND2_X1 U12554 ( .A1(n14108), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n16589) );
  CLKBUF_X1 U12555 ( .A(n10416), .Z(n19175) );
  NAND2_X1 U12556 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n20069) );
  INV_X1 U12557 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n19027) );
  INV_X1 U12558 ( .A(n17051), .ZN(n19030) );
  OR2_X1 U12559 ( .A1(n16772), .A2(P3_EBX_REG_30__SCAN_IN), .ZN(n10105) );
  NOR2_X1 U12560 ( .A1(n10104), .A2(n10103), .ZN(n10102) );
  NOR2_X1 U12561 ( .A1(n17102), .A2(n16769), .ZN(n10104) );
  INV_X1 U12562 ( .A(n16768), .ZN(n10103) );
  NAND2_X1 U12563 ( .A1(n10107), .A2(P3_EBX_REG_30__SCAN_IN), .ZN(n10106) );
  OR2_X1 U12564 ( .A1(n16766), .A2(n17059), .ZN(n10107) );
  NOR2_X1 U12565 ( .A1(n17104), .A2(n16752), .ZN(n16798) );
  NAND2_X1 U12566 ( .A1(n17101), .A2(n10366), .ZN(n16868) );
  NAND2_X1 U12567 ( .A1(n16868), .A2(n17807), .ZN(n16867) );
  AND2_X1 U12568 ( .A1(n17965), .A2(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n16994) );
  INV_X1 U12569 ( .A(n17101), .ZN(n17068) );
  INV_X1 U12570 ( .A(n17110), .ZN(n17086) );
  INV_X1 U12571 ( .A(n17114), .ZN(n17100) );
  INV_X1 U12572 ( .A(n17059), .ZN(n17111) );
  NOR3_X1 U12573 ( .A1(n17175), .A2(n21285), .A3(n16807), .ZN(n17174) );
  NOR2_X1 U12574 ( .A1(n17175), .A2(n21285), .ZN(n17178) );
  NOR2_X1 U12575 ( .A1(n17197), .A2(n17118), .ZN(n17179) );
  NAND2_X1 U12576 ( .A1(n17212), .A2(P3_EBX_REG_21__SCAN_IN), .ZN(n17197) );
  NOR2_X1 U12577 ( .A1(n17198), .A2(n18413), .ZN(n17212) );
  NOR2_X1 U12578 ( .A1(n17239), .A2(n21148), .ZN(n17215) );
  INV_X1 U12579 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n21148) );
  NOR2_X1 U12580 ( .A1(n16904), .A2(n17257), .ZN(n17271) );
  NOR2_X1 U12581 ( .A1(n10117), .A2(n9963), .ZN(n10116) );
  INV_X1 U12582 ( .A(n10118), .ZN(n10117) );
  NAND2_X1 U12583 ( .A1(n17375), .A2(P3_EBX_REG_10__SCAN_IN), .ZN(n17354) );
  NOR2_X1 U12584 ( .A1(n16996), .A2(n17374), .ZN(n17375) );
  NOR3_X1 U12585 ( .A1(n17404), .A2(n17022), .A3(n21274), .ZN(n17403) );
  INV_X1 U12586 ( .A(P3_EBX_REG_6__SCAN_IN), .ZN(n21274) );
  NOR4_X1 U12587 ( .A1(n17425), .A2(n12619), .A3(n17410), .A4(n17079), .ZN(
        n17413) );
  INV_X1 U12588 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n21090) );
  NOR2_X1 U12589 ( .A1(n17446), .A2(n17587), .ZN(n17440) );
  NAND2_X1 U12590 ( .A1(n17447), .A2(P3_EAX_REG_28__SCAN_IN), .ZN(n17446) );
  NOR3_X1 U12591 ( .A1(n17468), .A2(n18413), .A3(n10007), .ZN(n17459) );
  NOR3_X1 U12592 ( .A1(n17509), .A2(n17475), .A3(n17431), .ZN(n17469) );
  NOR2_X1 U12593 ( .A1(n17640), .A2(n17496), .ZN(n17491) );
  NAND2_X1 U12594 ( .A1(P3_EAX_REG_16__SCAN_IN), .A2(n17510), .ZN(n17509) );
  NAND2_X1 U12595 ( .A1(n17574), .A2(n10008), .ZN(n17514) );
  AND2_X1 U12596 ( .A1(n17520), .A2(n10009), .ZN(n10008) );
  NOR2_X1 U12597 ( .A1(n9960), .A2(n17430), .ZN(n10009) );
  AOI21_X1 U12598 ( .B1(n12552), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A(
        n13056), .ZN(n13061) );
  INV_X1 U12599 ( .A(n17580), .ZN(n17569) );
  NAND2_X1 U12600 ( .A1(n17631), .A2(n17582), .ZN(n17629) );
  INV_X1 U12601 ( .A(n17687), .ZN(n17678) );
  INV_X1 U12602 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n17688) );
  CLKBUF_X1 U12603 ( .A(n17677), .Z(n17684) );
  NOR2_X2 U12604 ( .A1(n19012), .A2(n17684), .ZN(n17685) );
  NAND3_X1 U12605 ( .A1(n19012), .A2(n17632), .A3(n17631), .ZN(n17687) );
  AND2_X1 U12606 ( .A1(n17882), .A2(n10109), .ZN(n17766) );
  AND2_X1 U12607 ( .A1(n10111), .A2(n10110), .ZN(n10109) );
  INV_X1 U12608 ( .A(n17786), .ZN(n10110) );
  INV_X1 U12609 ( .A(n17895), .ZN(n17919) );
  INV_X1 U12610 ( .A(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n17924) );
  AND2_X1 U12611 ( .A1(n17954), .A2(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n17965) );
  INV_X1 U12612 ( .A(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n17989) );
  AND2_X1 U12613 ( .A1(n18007), .A2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n17993) );
  NAND2_X1 U12614 ( .A1(n17995), .A2(n17996), .ZN(n17994) );
  INV_X1 U12615 ( .A(n16623), .ZN(n17708) );
  AND2_X1 U12616 ( .A1(n13163), .A2(n9974), .ZN(n17728) );
  INV_X1 U12617 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n18098) );
  AND2_X1 U12618 ( .A1(n10162), .A2(n9973), .ZN(n17848) );
  NAND2_X1 U12619 ( .A1(n18316), .A2(n18349), .ZN(n18350) );
  INV_X1 U12620 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n18283) );
  INV_X1 U12621 ( .A(n18824), .ZN(n18837) );
  INV_X1 U12622 ( .A(n18326), .ZN(n18364) );
  INV_X1 U12623 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18621) );
  INV_X1 U12624 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n18620) );
  INV_X1 U12625 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18845) );
  INV_X1 U12626 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n18847) );
  AOI22_X1 U12627 ( .A1(n18823), .A2(n12516), .B1(n18824), .B2(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n18992) );
  NAND2_X1 U12628 ( .A1(n18414), .A2(n18387), .ZN(n18758) );
  NAND2_X1 U12629 ( .A1(n18414), .A2(n18405), .ZN(n18782) );
  NAND2_X1 U12630 ( .A1(n18414), .A2(n18413), .ZN(n18799) );
  NAND2_X1 U12631 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n18877), .ZN(n18873) );
  OAI211_X1 U12632 ( .C1(P3_STATE_REG_1__SCAN_IN), .C2(P3_STATE_REG_2__SCAN_IN), .A(n18894), .B(n18954), .ZN(n19011) );
  INV_X1 U12633 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n18894) );
  NAND2_X1 U12634 ( .A1(n18894), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n19025) );
  AND2_X2 U12635 ( .A1(n12779), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n20303)
         );
  NOR2_X1 U12636 ( .A1(n14303), .A2(n13288), .ZN(n16647) );
  AOI21_X1 U12637 ( .B1(n10417), .B2(n12971), .A(n19214), .ZN(n10418) );
  AOI21_X1 U12638 ( .B1(n15624), .B2(n19315), .A(n12838), .ZN(n12843) );
  OAI21_X1 U12639 ( .B1(n16480), .B2(n19319), .A(n10090), .ZN(P2_U2992) );
  AOI21_X1 U12640 ( .B1(n16482), .B2(n12840), .A(n10091), .ZN(n10090) );
  INV_X1 U12641 ( .A(n10092), .ZN(n10091) );
  AOI21_X1 U12642 ( .B1(n16481), .B2(n19315), .A(n10093), .ZN(n10092) );
  OAI21_X1 U12643 ( .B1(n15809), .B2(n19356), .A(n11519), .ZN(n11520) );
  OAI21_X1 U12644 ( .B1(n10108), .B2(n18873), .A(n10100), .ZN(P3_U2641) );
  XNOR2_X1 U12645 ( .A(n16764), .B(n16765), .ZN(n10108) );
  AND2_X1 U12646 ( .A1(n10106), .A2(n10101), .ZN(n10100) );
  AND2_X1 U12647 ( .A1(n10105), .A2(n10102), .ZN(n10101) );
  OAI21_X1 U12648 ( .B1(n12694), .B2(P3_EBX_REG_28__SCAN_IN), .A(n12693), .ZN(
        n12695) );
  INV_X1 U12649 ( .A(n17447), .ZN(n17450) );
  NAND2_X1 U12650 ( .A1(n17574), .A2(n17520), .ZN(n17543) );
  AOI21_X1 U12651 ( .B1(n13271), .B2(n17926), .A(n13240), .ZN(n13241) );
  OAI21_X1 U12652 ( .B1(n13269), .B2(n18050), .A(n13239), .ZN(n13240) );
  AOI21_X1 U12653 ( .B1(n13271), .B2(n18288), .A(n13270), .ZN(n13272) );
  OAI21_X1 U12654 ( .B1(n13269), .B2(n18326), .A(n13268), .ZN(n13270) );
  AOI221_X1 U12655 ( .B1(n16643), .B2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), 
        .C1(n16642), .C2(n17693), .A(n16641), .ZN(n16644) );
  NAND2_X1 U12656 ( .A1(n16647), .A2(U214), .ZN(U212) );
  INV_X4 U12657 ( .A(n17252), .ZN(n13120) );
  NAND2_X1 U12658 ( .A1(n20358), .A2(n11741), .ZN(n13838) );
  AND2_X2 U12659 ( .A1(n16000), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n9861) );
  AND2_X1 U12660 ( .A1(n13586), .A2(n14341), .ZN(n9862) );
  NAND2_X1 U12661 ( .A1(n10404), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n10401) );
  NAND2_X1 U12662 ( .A1(n10304), .A2(n10376), .ZN(n15822) );
  NAND2_X1 U12663 ( .A1(n15782), .A2(n15780), .ZN(n15772) );
  OR3_X1 U12664 ( .A1(n15689), .A2(n15688), .A3(n10158), .ZN(n9863) );
  NAND2_X1 U12665 ( .A1(n15771), .A2(n15895), .ZN(n9864) );
  NOR2_X1 U12666 ( .A1(n16074), .A2(n9924), .ZN(n9865) );
  NAND2_X1 U12667 ( .A1(n11299), .A2(n9893), .ZN(n11307) );
  AND2_X1 U12668 ( .A1(n10131), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n9866) );
  OR3_X1 U12669 ( .A1(n14861), .A2(n10200), .A3(n14837), .ZN(n9867) );
  AND2_X1 U12670 ( .A1(n10321), .A2(n16080), .ZN(n9868) );
  AND2_X1 U12671 ( .A1(n18413), .A2(n13246), .ZN(n9869) );
  AND2_X1 U12672 ( .A1(n12800), .A2(n15749), .ZN(n9870) );
  NOR2_X1 U12673 ( .A1(n16074), .A2(n9932), .ZN(n14442) );
  NOR2_X1 U12674 ( .A1(n15663), .A2(n14644), .ZN(n15656) );
  INV_X1 U12675 ( .A(n11306), .ZN(n10323) );
  AND2_X1 U12676 ( .A1(n10898), .A2(n9948), .ZN(n9871) );
  AND2_X1 U12677 ( .A1(n13541), .A2(n10334), .ZN(n9872) );
  AND2_X1 U12678 ( .A1(n9866), .A2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n9873) );
  NAND2_X1 U12679 ( .A1(n9947), .A2(n10371), .ZN(n14543) );
  OAI21_X1 U12680 ( .B1(n13194), .B2(n13193), .A(n13192), .ZN(n18802) );
  AND2_X1 U12681 ( .A1(n10097), .A2(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n9874) );
  NAND2_X1 U12682 ( .A1(n13662), .A2(n10150), .ZN(n13709) );
  AND2_X1 U12683 ( .A1(n10140), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n9875) );
  AND2_X1 U12684 ( .A1(n9926), .A2(n10585), .ZN(n9876) );
  NOR2_X1 U12685 ( .A1(n10722), .A2(n9925), .ZN(n9877) );
  AND2_X1 U12686 ( .A1(n14979), .A2(n15035), .ZN(n9878) );
  INV_X1 U12687 ( .A(n10241), .ZN(n10240) );
  NAND2_X1 U12688 ( .A1(n10243), .A2(n12436), .ZN(n10241) );
  OR2_X1 U12689 ( .A1(n14875), .A2(n14888), .ZN(n9879) );
  AND2_X1 U12690 ( .A1(n9874), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n9880) );
  NAND2_X1 U12691 ( .A1(n11020), .A2(n10073), .ZN(n10147) );
  INV_X1 U12692 ( .A(n19356), .ZN(n16577) );
  AND2_X1 U12693 ( .A1(n10142), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n9881) );
  AND2_X1 U12694 ( .A1(n10116), .A2(P3_EBX_REG_15__SCAN_IN), .ZN(n9882) );
  AND2_X1 U12695 ( .A1(n10307), .A2(n9965), .ZN(n9883) );
  INV_X1 U12696 ( .A(n12561), .ZN(n13064) );
  INV_X1 U12697 ( .A(n13082), .ZN(n12561) );
  OR3_X1 U12698 ( .A1(n17468), .A2(n18413), .A3(n10006), .ZN(n9885) );
  NAND2_X1 U12699 ( .A1(n10999), .A2(n10998), .ZN(n11153) );
  OR2_X1 U12700 ( .A1(n15717), .A2(n13320), .ZN(n9886) );
  OR2_X1 U12701 ( .A1(n15039), .A2(n10202), .ZN(n9887) );
  OR2_X1 U12702 ( .A1(n11341), .A2(n10584), .ZN(n9888) );
  NAND2_X1 U12703 ( .A1(n14915), .A2(n10338), .ZN(n14873) );
  NAND2_X1 U12704 ( .A1(n10082), .A2(n11461), .ZN(n14530) );
  INV_X1 U12705 ( .A(n10935), .ZN(n10680) );
  OR2_X1 U12706 ( .A1(P2_EBX_REG_26__SCAN_IN), .A2(n12462), .ZN(n9889) );
  AND2_X1 U12707 ( .A1(n14943), .A2(n14942), .ZN(n14944) );
  NAND2_X1 U12708 ( .A1(n11299), .A2(n11298), .ZN(n9890) );
  AND2_X1 U12709 ( .A1(n11463), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15934) );
  NOR2_X1 U12710 ( .A1(n15834), .A2(n10305), .ZN(n11464) );
  NOR2_X4 U12711 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n16153), .ZN(
        n13079) );
  NOR2_X1 U12712 ( .A1(n10403), .A2(n16529), .ZN(n10404) );
  AND2_X1 U12713 ( .A1(n10407), .A2(n10138), .ZN(n9891) );
  AND2_X1 U12714 ( .A1(n10219), .A2(n12828), .ZN(n9892) );
  AND2_X1 U12715 ( .A1(n11298), .A2(n10583), .ZN(n9893) );
  OR2_X1 U12716 ( .A1(n14833), .A2(n10349), .ZN(n14821) );
  AND2_X1 U12717 ( .A1(n14915), .A2(n14914), .ZN(n14900) );
  OR2_X1 U12718 ( .A1(n11449), .A2(n11447), .ZN(n9894) );
  OR2_X1 U12719 ( .A1(n17175), .A2(n10127), .ZN(n9895) );
  NOR2_X1 U12720 ( .A1(n18840), .A2(n12513), .ZN(n13083) );
  INV_X1 U12721 ( .A(n13083), .ZN(n13051) );
  OAI21_X1 U12722 ( .B1(n14410), .B2(n10067), .A(n10065), .ZN(n16513) );
  NAND2_X1 U12723 ( .A1(n10315), .A2(n12440), .ZN(n15949) );
  NAND2_X1 U12724 ( .A1(n10087), .A2(n10088), .ZN(n16537) );
  AND2_X1 U12725 ( .A1(n10146), .A2(n10145), .ZN(n9896) );
  AND2_X1 U12726 ( .A1(n9893), .A2(n10175), .ZN(n9897) );
  INV_X1 U12727 ( .A(n10095), .ZN(n11463) );
  AND2_X1 U12728 ( .A1(n10242), .A2(n10240), .ZN(n9898) );
  AND4_X1 U12729 ( .A1(n12429), .A2(n16015), .A3(n12428), .A4(n15841), .ZN(
        n9899) );
  AND2_X1 U12730 ( .A1(n11440), .A2(n11256), .ZN(n9900) );
  AND2_X1 U12731 ( .A1(n11178), .A2(n9860), .ZN(n11223) );
  INV_X1 U12732 ( .A(n11651), .ZN(n11635) );
  NAND2_X1 U12733 ( .A1(n9990), .A2(n10293), .ZN(n15213) );
  AND2_X1 U12734 ( .A1(n11169), .A2(n11171), .ZN(n11217) );
  AND2_X1 U12735 ( .A1(n13089), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n9901) );
  AND3_X1 U12736 ( .A1(n10011), .A2(n12580), .A3(n10010), .ZN(n9902) );
  NAND3_X1 U12737 ( .A1(n11185), .A2(n11206), .A3(n10080), .ZN(n11291) );
  XNOR2_X1 U12738 ( .A(n11831), .B(n11731), .ZN(n11984) );
  INV_X1 U12739 ( .A(n10162), .ZN(n13155) );
  NAND2_X1 U12740 ( .A1(n10324), .A2(n10323), .ZN(n14538) );
  NAND2_X1 U12741 ( .A1(n14943), .A2(n10344), .ZN(n15004) );
  AND2_X1 U12742 ( .A1(n11141), .A2(n11138), .ZN(n9903) );
  AND3_X1 U12743 ( .A1(n16232), .A2(n19012), .A3(n16231), .ZN(n9904) );
  INV_X1 U12744 ( .A(n10319), .ZN(n10318) );
  OAI21_X1 U12745 ( .B1(n11313), .B2(n10320), .A(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n10319) );
  AND2_X1 U12746 ( .A1(n13150), .A2(n18283), .ZN(n9905) );
  AND2_X1 U12747 ( .A1(n10242), .A2(n10243), .ZN(n9906) );
  NAND2_X1 U12748 ( .A1(n11253), .A2(n11457), .ZN(n11447) );
  INV_X1 U12749 ( .A(n11872), .ZN(n10288) );
  NOR2_X1 U12750 ( .A1(n15643), .A2(n15642), .ZN(n13317) );
  AND3_X1 U12751 ( .A1(n11169), .A2(n14805), .A3(n19354), .ZN(n11216) );
  AND4_X1 U12752 ( .A1(n10125), .A2(n10121), .A3(n12570), .A4(n12569), .ZN(
        n9908) );
  INV_X1 U12753 ( .A(n11141), .ZN(n10073) );
  INV_X1 U12754 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10607) );
  INV_X1 U12755 ( .A(n11290), .ZN(n10311) );
  NAND2_X1 U12756 ( .A1(n11233), .A2(n11232), .ZN(n11290) );
  AND2_X1 U12757 ( .A1(n10014), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n9909) );
  NAND2_X1 U12758 ( .A1(n10473), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9910) );
  NAND2_X1 U12759 ( .A1(n10940), .A2(n10939), .ZN(n10942) );
  NAND2_X1 U12760 ( .A1(n10951), .A2(n19384), .ZN(n11486) );
  OR2_X1 U12761 ( .A1(n13171), .A2(n12618), .ZN(n9911) );
  OR2_X1 U12762 ( .A1(n17306), .A2(n17261), .ZN(n9912) );
  NAND2_X1 U12763 ( .A1(n16093), .A2(n16090), .ZN(n9913) );
  NAND2_X1 U12764 ( .A1(n9861), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n15834) );
  NAND2_X1 U12766 ( .A1(n9861), .A2(n10096), .ZN(n10095) );
  NAND2_X1 U12767 ( .A1(n10340), .A2(n12089), .ZN(n14976) );
  INV_X1 U12768 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n18972) );
  OR2_X1 U12769 ( .A1(n14408), .A2(n14421), .ZN(n9914) );
  AND2_X1 U12770 ( .A1(n13317), .A2(n13318), .ZN(n13316) );
  AND3_X1 U12771 ( .A1(n18982), .A2(n12506), .A3(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n9915) );
  OAI21_X1 U12772 ( .B1(n12426), .B2(n11254), .A(n12425), .ZN(n12800) );
  AND2_X1 U12773 ( .A1(n11648), .A2(n13839), .ZN(n9916) );
  NOR2_X1 U12774 ( .A1(n15246), .A2(n15243), .ZN(n9917) );
  AND2_X1 U12775 ( .A1(n9897), .A2(n19122), .ZN(n9918) );
  INV_X1 U12776 ( .A(n11313), .ZN(n10322) );
  INV_X1 U12777 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10144) );
  INV_X1 U12778 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n12506) );
  AND2_X2 U12779 ( .A1(n10959), .A2(n20013), .ZN(n10690) );
  OAI21_X1 U12780 ( .B1(n11747), .B2(n11746), .A(n13471), .ZN(n13553) );
  OR2_X1 U12781 ( .A1(n12509), .A2(n12508), .ZN(n9919) );
  AND2_X1 U12782 ( .A1(n17375), .A2(n10118), .ZN(n9920) );
  NOR2_X1 U12783 ( .A1(n9871), .A2(n15591), .ZN(n9921) );
  AND2_X1 U12784 ( .A1(n17882), .A2(n10113), .ZN(n9922) );
  INV_X1 U12785 ( .A(n11643), .ZN(n10042) );
  NOR2_X1 U12786 ( .A1(n14027), .A2(n14028), .ZN(n14026) );
  AND2_X1 U12787 ( .A1(n14962), .A2(n12179), .ZN(n14943) );
  NOR2_X1 U12788 ( .A1(n14457), .A2(n10342), .ZN(n14980) );
  NOR2_X2 U12789 ( .A1(n17551), .A2(n16638), .ZN(n17957) );
  NOR2_X1 U12790 ( .A1(n17933), .A2(n10164), .ZN(n17868) );
  NOR2_X1 U12791 ( .A1(n10414), .A2(n15808), .ZN(n10397) );
  AND2_X1 U12792 ( .A1(n10404), .A2(n10131), .ZN(n10402) );
  AND2_X1 U12793 ( .A1(n10400), .A2(n10140), .ZN(n9923) );
  NAND2_X1 U12794 ( .A1(n12566), .A2(n12565), .ZN(n18401) );
  INV_X1 U12795 ( .A(n18401), .ZN(n10005) );
  INV_X1 U12796 ( .A(n11854), .ZN(n10058) );
  NOR2_X1 U12797 ( .A1(n14878), .A2(n14862), .ZN(n12922) );
  XNOR2_X1 U12798 ( .A(n11984), .B(n11985), .ZN(n13973) );
  NAND2_X1 U12799 ( .A1(n14281), .A2(n14206), .ZN(n14254) );
  NAND2_X1 U12800 ( .A1(n10333), .A2(n14289), .ZN(n14288) );
  OR2_X1 U12801 ( .A1(n10255), .A2(n16050), .ZN(n9924) );
  OR2_X1 U12802 ( .A1(n10234), .A2(n14160), .ZN(n9925) );
  NAND2_X1 U12803 ( .A1(n14478), .A2(n11456), .ZN(n14407) );
  NAND2_X1 U12804 ( .A1(n10300), .A2(n11900), .ZN(n14499) );
  NAND2_X1 U12805 ( .A1(n10070), .A2(n10321), .ZN(n15864) );
  AND2_X1 U12806 ( .A1(n14026), .A2(n14282), .ZN(n14251) );
  NOR2_X1 U12807 ( .A1(n16074), .A2(n15620), .ZN(n15619) );
  AND2_X1 U12808 ( .A1(n11353), .A2(n11348), .ZN(n9926) );
  INV_X1 U12809 ( .A(n16310), .ZN(n10047) );
  INV_X1 U12810 ( .A(n19012), .ZN(n18387) );
  OAI211_X1 U12811 ( .C1(n11448), .C2(n9894), .A(n11452), .B(n11451), .ZN(
        n14477) );
  OR3_X1 U12812 ( .A1(n15039), .A2(n10204), .A3(n10207), .ZN(n9927) );
  AND2_X1 U12813 ( .A1(n10400), .A2(n10139), .ZN(n10398) );
  NOR2_X1 U12814 ( .A1(n15656), .A2(n15657), .ZN(n9928) );
  AND2_X1 U12815 ( .A1(n11205), .A2(n11184), .ZN(n9929) );
  NOR2_X1 U12816 ( .A1(n10890), .A2(n11254), .ZN(n9930) );
  INV_X1 U12817 ( .A(n13511), .ZN(n10040) );
  INV_X1 U12818 ( .A(n10182), .ZN(n11433) );
  OR3_X1 U12819 ( .A1(n10512), .A2(n10511), .A3(n10357), .ZN(n10182) );
  INV_X1 U12820 ( .A(n12436), .ZN(n16025) );
  AND2_X1 U12821 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n9931) );
  INV_X1 U12822 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n19111) );
  INV_X1 U12823 ( .A(n10345), .ZN(n10344) );
  NAND2_X1 U12824 ( .A1(n15012), .A2(n14942), .ZN(n10345) );
  INV_X1 U12825 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n20310) );
  INV_X1 U12826 ( .A(n10339), .ZN(n10338) );
  NAND2_X1 U12827 ( .A1(n14914), .A2(n14901), .ZN(n10339) );
  NOR2_X1 U12828 ( .A1(n14020), .A2(n14249), .ZN(n14289) );
  OR2_X1 U12829 ( .A1(n9924), .A2(n10257), .ZN(n9932) );
  AND2_X1 U12830 ( .A1(n11679), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n9933) );
  AND2_X1 U12831 ( .A1(n10247), .A2(n12808), .ZN(n9934) );
  AND2_X1 U12832 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n9935) );
  AND2_X1 U12833 ( .A1(n15028), .A2(n10341), .ZN(n9936) );
  NOR2_X1 U12834 ( .A1(n9845), .A2(n15331), .ZN(n9937) );
  AND2_X1 U12835 ( .A1(n10187), .A2(n10186), .ZN(n9938) );
  NOR2_X1 U12836 ( .A1(n10890), .A2(n11250), .ZN(n9939) );
  NAND2_X1 U12837 ( .A1(n11299), .A2(n9897), .ZN(n9940) );
  AND2_X1 U12838 ( .A1(n10898), .A2(n10253), .ZN(n9941) );
  AND2_X1 U12839 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n9942) );
  AND2_X1 U12840 ( .A1(n9876), .A2(n10189), .ZN(n9943) );
  INV_X1 U12841 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n19064) );
  OR2_X1 U12842 ( .A1(n9925), .A2(n10233), .ZN(n9944) );
  AOI22_X1 U12843 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_31__SCAN_IN), .B1(n12834), .B2(n14298), .ZN(
        n10415) );
  INV_X1 U12844 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n13362) );
  INV_X1 U12845 ( .A(n19355), .ZN(n19341) );
  NAND2_X1 U12846 ( .A1(n11505), .A2(n11472), .ZN(n19327) );
  OR2_X1 U12847 ( .A1(n13915), .A2(n10252), .ZN(n13872) );
  AND2_X1 U12848 ( .A1(n14281), .A2(n10280), .ZN(n9945) );
  OR2_X1 U12849 ( .A1(n10722), .A2(n9944), .ZN(n14171) );
  NAND2_X1 U12850 ( .A1(n13702), .A2(n13701), .ZN(n13703) );
  NAND2_X1 U12851 ( .A1(n9992), .A2(n9991), .ZN(n20358) );
  AND2_X1 U12852 ( .A1(n10147), .A2(n9896), .ZN(n13602) );
  NOR2_X1 U12853 ( .A1(n20597), .A2(n20313), .ZN(n9946) );
  AND2_X1 U12854 ( .A1(n10253), .A2(n15590), .ZN(n9948) );
  INV_X1 U12855 ( .A(n19319), .ZN(n16539) );
  OR2_X1 U12856 ( .A1(n19042), .A2(n20062), .ZN(n19319) );
  OR3_X1 U12857 ( .A1(n14665), .A2(n14664), .A3(n15659), .ZN(n9949) );
  NAND2_X1 U12858 ( .A1(n13662), .A2(n10151), .ZN(n9950) );
  AND2_X1 U12859 ( .A1(n15538), .A2(n15554), .ZN(n9951) );
  AND2_X1 U12860 ( .A1(n10259), .A2(n10258), .ZN(n9952) );
  AND2_X1 U12861 ( .A1(n10184), .A2(n10183), .ZN(n9953) );
  INV_X1 U12862 ( .A(n11319), .ZN(n10188) );
  INV_X1 U12863 ( .A(n12443), .ZN(n10185) );
  AND2_X1 U12864 ( .A1(n17375), .A2(n10116), .ZN(n9954) );
  NAND2_X1 U12865 ( .A1(n10336), .A2(n10334), .ZN(n13728) );
  AND2_X1 U12866 ( .A1(n10195), .A2(n10194), .ZN(n9955) );
  OR2_X1 U12867 ( .A1(n12089), .A2(n12101), .ZN(n9956) );
  AND2_X1 U12868 ( .A1(n9952), .A2(n15718), .ZN(n9957) );
  INV_X1 U12869 ( .A(n13350), .ZN(n13587) );
  NAND2_X1 U12870 ( .A1(n14298), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n13350) );
  NAND2_X1 U12871 ( .A1(n13461), .A2(n13548), .ZN(n13464) );
  AND2_X1 U12872 ( .A1(n9948), .A2(n11473), .ZN(n9958) );
  AND2_X1 U12873 ( .A1(n9953), .A2(n15653), .ZN(n9959) );
  INV_X1 U12874 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n14270) );
  NAND3_X1 U12875 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(P3_EAX_REG_8__SCAN_IN), 
        .A3(P3_EAX_REG_12__SCAN_IN), .ZN(n9960) );
  NAND2_X1 U12876 ( .A1(READY22_REG_SCAN_IN), .A2(READY2), .ZN(n18858) );
  INV_X1 U12877 ( .A(n18858), .ZN(n9998) );
  XOR2_X1 U12878 ( .A(n11273), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .Z(n9961) );
  INV_X1 U12879 ( .A(n11254), .ZN(n12808) );
  INV_X1 U12880 ( .A(n12763), .ZN(n16196) );
  AND2_X1 U12881 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13946) );
  AND2_X1 U12882 ( .A1(n17722), .A2(n10097), .ZN(n9962) );
  INV_X1 U12883 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16080) );
  NAND3_X1 U12884 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(P3_EBX_REG_12__SCAN_IN), 
        .A3(P3_EBX_REG_13__SCAN_IN), .ZN(n9963) );
  INV_X1 U12885 ( .A(n10165), .ZN(n10164) );
  AND2_X1 U12886 ( .A1(n10168), .A2(n10166), .ZN(n10165) );
  INV_X1 U12887 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n18295) );
  INV_X1 U12888 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n10180) );
  INV_X1 U12889 ( .A(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n10098) );
  INV_X1 U12890 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15963) );
  INV_X1 U12891 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n16923) );
  AND2_X1 U12892 ( .A1(n9883), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n9964) );
  INV_X1 U12893 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n10166) );
  INV_X1 U12894 ( .A(P2_EBX_REG_24__SCAN_IN), .ZN(n10183) );
  AND2_X1 U12895 ( .A1(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n9965) );
  INV_X1 U12896 ( .A(P2_EBX_REG_10__SCAN_IN), .ZN(n10175) );
  INV_X1 U12897 ( .A(P2_EBX_REG_21__SCAN_IN), .ZN(n10189) );
  OAI21_X1 U12898 ( .B1(n19646), .B2(n19661), .A(n19861), .ZN(n19663) );
  NAND2_X1 U12899 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19861), .ZN(n19412) );
  INV_X1 U12900 ( .A(n19861), .ZN(n19610) );
  AOI22_X1 U12901 ( .A1(n18996), .A2(n18997), .B1(n12516), .B2(n18998), .ZN(
        P3_U3290) );
  CLKBUF_X1 U12902 ( .A(n19873), .Z(n9966) );
  NAND2_X1 U12903 ( .A1(n9968), .A2(n9967), .ZN(n18332) );
  OR2_X1 U12904 ( .A1(n18017), .A2(n18018), .ZN(n9967) );
  NAND2_X1 U12905 ( .A1(n18017), .A2(n18018), .ZN(n9968) );
  NAND3_X1 U12906 ( .A1(n10162), .A2(n9973), .A3(n17847), .ZN(n17846) );
  NAND3_X1 U12907 ( .A1(n13163), .A2(n18054), .A3(n9974), .ZN(n17727) );
  NAND3_X1 U12908 ( .A1(n17756), .A2(n17760), .A3(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n13164) );
  INV_X1 U12909 ( .A(n9979), .ZN(n17975) );
  NAND2_X1 U12910 ( .A1(n13745), .A2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13744) );
  NOR2_X2 U12911 ( .A1(n18221), .A2(n13230), .ZN(n18195) );
  NAND2_X2 U12912 ( .A1(n17958), .A2(n13229), .ZN(n18215) );
  NAND2_X1 U12913 ( .A1(n16329), .A2(n16331), .ZN(n9981) );
  NAND3_X1 U12914 ( .A1(n10284), .A2(n10286), .A3(n11880), .ZN(n9982) );
  NAND2_X1 U12915 ( .A1(n11821), .A2(n10013), .ZN(n13971) );
  NAND2_X2 U12916 ( .A1(n9984), .A2(n9983), .ZN(n10013) );
  OR3_X2 U12917 ( .A1(n13002), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        n13000), .ZN(n9985) );
  NAND2_X2 U12918 ( .A1(n9985), .A2(n16302), .ZN(n15146) );
  NAND2_X1 U12919 ( .A1(n9987), .A2(n10293), .ZN(n10290) );
  NAND2_X1 U12920 ( .A1(n9837), .A2(n11906), .ZN(n9987) );
  INV_X1 U12921 ( .A(n11678), .ZN(n9992) );
  INV_X1 U12922 ( .A(n20423), .ZN(n9991) );
  NAND3_X1 U12923 ( .A1(n20358), .A2(n20310), .A3(n11741), .ZN(n9993) );
  NAND3_X1 U12924 ( .A1(n13762), .A2(n11816), .A3(n12766), .ZN(n9994) );
  NAND2_X1 U12925 ( .A1(n11979), .A2(n12766), .ZN(n11643) );
  NAND2_X1 U12926 ( .A1(n11598), .A2(n11640), .ZN(n9995) );
  AOI21_X1 U12927 ( .B1(n16229), .B2(n9997), .A(n9904), .ZN(n9996) );
  NAND3_X1 U12928 ( .A1(n13180), .A2(n10003), .A3(n10002), .ZN(n13244) );
  NOR2_X1 U12929 ( .A1(n17468), .A2(n18413), .ZN(n17464) );
  INV_X1 U12930 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n10007) );
  INV_X1 U12931 ( .A(n17459), .ZN(n17463) );
  NAND2_X1 U12932 ( .A1(n10013), .A2(n13974), .ZN(n11845) );
  NAND2_X2 U12933 ( .A1(n10015), .A2(n11911), .ZN(n13002) );
  INV_X1 U12934 ( .A(n15182), .ZN(n10015) );
  CLKBUF_X1 U12935 ( .A(n12723), .Z(n10016) );
  OAI21_X2 U12936 ( .B1(n11661), .B2(n10039), .A(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n11742) );
  NAND3_X1 U12937 ( .A1(n10037), .A2(n11660), .A3(n10036), .ZN(n11662) );
  NAND2_X1 U12938 ( .A1(n11656), .A2(n11658), .ZN(n13518) );
  NAND3_X2 U12939 ( .A1(n13793), .A2(n10044), .A3(n10363), .ZN(n11661) );
  AND2_X2 U12940 ( .A1(n13473), .A2(n13464), .ZN(n13793) );
  XNOR2_X1 U12941 ( .A(n16302), .B(n16359), .ZN(n15226) );
  NAND2_X1 U12942 ( .A1(n10049), .A2(n15224), .ZN(n10048) );
  NAND2_X1 U12943 ( .A1(n10050), .A2(n9917), .ZN(n15220) );
  NOR2_X1 U12944 ( .A1(n11746), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10051) );
  NAND2_X1 U12945 ( .A1(n11747), .A2(n10051), .ZN(n10052) );
  NAND2_X1 U12946 ( .A1(n11746), .A2(n20310), .ZN(n10053) );
  AND2_X1 U12947 ( .A1(n12031), .A2(n11886), .ZN(n10057) );
  INV_X1 U12948 ( .A(n11855), .ZN(n10060) );
  NAND2_X1 U12949 ( .A1(n10060), .A2(n10059), .ZN(n11874) );
  OR2_X2 U12950 ( .A1(n11855), .A2(n10058), .ZN(n11863) );
  INV_X1 U12951 ( .A(n11862), .ZN(n10061) );
  NAND2_X1 U12952 ( .A1(n14410), .A2(n10065), .ZN(n10064) );
  NOR2_X2 U12953 ( .A1(n10975), .A2(n10071), .ZN(n11496) );
  NAND3_X1 U12954 ( .A1(n10311), .A2(n11450), .A3(n10074), .ZN(n11457) );
  NAND2_X2 U12955 ( .A1(n12456), .A2(n15793), .ZN(n15782) );
  NOR2_X1 U12956 ( .A1(n13627), .A2(n11157), .ZN(n11158) );
  NOR2_X1 U12957 ( .A1(n13627), .A2(n11159), .ZN(n11161) );
  NAND2_X1 U12958 ( .A1(n10974), .A2(n13676), .ZN(n10301) );
  NAND2_X2 U12959 ( .A1(n10301), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11006) );
  AND2_X2 U12960 ( .A1(n11496), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11021) );
  NAND3_X1 U12961 ( .A1(n11185), .A2(n11206), .A3(n9929), .ZN(n11440) );
  INV_X1 U12962 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n10099) );
  INV_X1 U12963 ( .A(n13296), .ZN(n10115) );
  XNOR2_X2 U12964 ( .A(n13233), .B(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n17101) );
  NAND3_X1 U12965 ( .A1(n12572), .A2(n9908), .A3(n10120), .ZN(n18409) );
  NAND3_X1 U12966 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(P3_EBX_REG_26__SCAN_IN), 
        .A3(P3_EBX_REG_25__SCAN_IN), .ZN(n10127) );
  NAND2_X1 U12967 ( .A1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n10405) );
  NAND3_X1 U12968 ( .A1(n10407), .A2(n10138), .A3(
        P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n10408) );
  NOR2_X2 U12969 ( .A1(n12486), .A2(n12487), .ZN(n10154) );
  NOR2_X1 U12970 ( .A1(n15689), .A2(n15688), .ZN(n15691) );
  INV_X1 U12971 ( .A(n15588), .ZN(n10158) );
  INV_X1 U12972 ( .A(n10159), .ZN(n11466) );
  NAND2_X1 U12973 ( .A1(n15553), .A2(n10160), .ZN(n15643) );
  OAI21_X1 U12974 ( .B1(n17933), .B2(n10163), .A(n13160), .ZN(n10162) );
  NOR2_X1 U12975 ( .A1(n17933), .A2(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n17927) );
  AND2_X2 U12976 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n9915), .ZN(
        n17344) );
  NAND3_X1 U12977 ( .A1(n10172), .A2(n10171), .A3(n10369), .ZN(n10170) );
  NAND3_X1 U12978 ( .A1(n10174), .A2(n12800), .A3(n10173), .ZN(n10172) );
  NAND2_X1 U12979 ( .A1(n11299), .A2(n9918), .ZN(n11320) );
  NAND3_X1 U12980 ( .A1(n17727), .A2(n13165), .A3(n10179), .ZN(n10176) );
  NAND2_X1 U12981 ( .A1(n10176), .A2(n10178), .ZN(n17697) );
  AND3_X1 U12982 ( .A1(n17727), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A3(
        n13165), .ZN(n16623) );
  NAND2_X1 U12983 ( .A1(n17727), .A2(n13165), .ZN(n10177) );
  NAND2_X1 U12984 ( .A1(n13160), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n10178) );
  NAND2_X1 U12985 ( .A1(n17957), .A2(n10180), .ZN(n10179) );
  NAND2_X1 U12986 ( .A1(n11135), .A2(n9959), .ZN(n12462) );
  NAND2_X1 U12987 ( .A1(n11135), .A2(n12443), .ZN(n12449) );
  NAND2_X1 U12988 ( .A1(n11349), .A2(n9943), .ZN(n12444) );
  AND2_X1 U12989 ( .A1(n11349), .A2(n9926), .ZN(n11352) );
  AND2_X1 U12990 ( .A1(n11349), .A2(n11348), .ZN(n11354) );
  NAND2_X1 U12991 ( .A1(n13743), .A2(n13742), .ZN(n13741) );
  INV_X1 U12992 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10190) );
  NAND2_X1 U12993 ( .A1(n14045), .A2(n10191), .ZN(n16424) );
  NAND2_X1 U12994 ( .A1(n10193), .A2(n16422), .ZN(n16423) );
  NAND2_X1 U12995 ( .A1(n14046), .A2(n10193), .ZN(n20257) );
  NAND2_X1 U12996 ( .A1(n12854), .A2(n12853), .ZN(n10198) );
  NAND2_X1 U12997 ( .A1(n10198), .A2(n10197), .ZN(n13754) );
  NAND3_X1 U12998 ( .A1(n10203), .A2(n10206), .A3(n12899), .ZN(n10202) );
  INV_X1 U12999 ( .A(n12899), .ZN(n10207) );
  NAND4_X1 U13000 ( .A1(n10640), .A2(n10641), .A3(n10642), .A4(n10643), .ZN(
        n10209) );
  NAND2_X1 U13001 ( .A1(n10211), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10210) );
  NAND4_X1 U13002 ( .A1(n10650), .A2(n10652), .A3(n10651), .A4(n10653), .ZN(
        n10211) );
  NAND2_X1 U13003 ( .A1(n10213), .A2(n10212), .ZN(n11256) );
  AND2_X2 U13004 ( .A1(n19342), .A2(n11162), .ZN(n11210) );
  NAND2_X2 U13005 ( .A1(n10266), .A2(n10267), .ZN(n10265) );
  NAND2_X1 U13006 ( .A1(n10217), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10215) );
  INV_X1 U13007 ( .A(n10217), .ZN(n10981) );
  NAND2_X1 U13008 ( .A1(n15510), .A2(n10218), .ZN(n12823) );
  NAND3_X1 U13009 ( .A1(n10676), .A2(n10671), .A3(n10223), .ZN(n10222) );
  NAND3_X1 U13010 ( .A1(n10677), .A2(n10675), .A3(n10678), .ZN(n10224) );
  NAND2_X1 U13011 ( .A1(n10229), .A2(n10228), .ZN(n11275) );
  NOR2_X1 U13012 ( .A1(n10230), .A2(n9961), .ZN(n10228) );
  INV_X1 U13013 ( .A(n10722), .ZN(n14414) );
  NAND2_X1 U13014 ( .A1(n16041), .A2(n10237), .ZN(n10235) );
  NAND2_X1 U13015 ( .A1(n10235), .A2(n10236), .ZN(n15842) );
  NOR2_X1 U13016 ( .A1(n13914), .A2(n13913), .ZN(n13915) );
  NOR2_X1 U13017 ( .A1(n13915), .A2(n10706), .ZN(n13873) );
  INV_X1 U13018 ( .A(n16028), .ZN(n10257) );
  NAND4_X1 U13019 ( .A1(n10263), .A2(n10265), .A3(n9862), .A4(n11143), .ZN(
        n10262) );
  INV_X1 U13020 ( .A(n14644), .ZN(n10269) );
  NAND2_X1 U13021 ( .A1(n10269), .A2(n9949), .ZN(n10270) );
  OAI21_X2 U13022 ( .B1(n15663), .B2(n10270), .A(n10271), .ZN(n14686) );
  NAND2_X1 U13023 ( .A1(n10467), .A2(n10607), .ZN(n10272) );
  NAND2_X1 U13024 ( .A1(n10461), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10273) );
  OAI21_X2 U13025 ( .B1(n10277), .B2(n9910), .A(n10274), .ZN(n10935) );
  NAND3_X1 U13026 ( .A1(n10367), .A2(n10607), .A3(n10370), .ZN(n10274) );
  NAND2_X1 U13027 ( .A1(n10966), .A2(n20064), .ZN(n10967) );
  NAND2_X2 U13028 ( .A1(n10276), .A2(n10275), .ZN(n10679) );
  NAND4_X1 U13029 ( .A1(n10599), .A2(n10600), .A3(n10601), .A4(n10602), .ZN(
        n10275) );
  NAND3_X1 U13030 ( .A1(n10596), .A2(n10594), .A3(n10595), .ZN(n10276) );
  NAND3_X1 U13031 ( .A1(n10474), .A2(n10475), .A3(n10476), .ZN(n10277) );
  NAND2_X1 U13032 ( .A1(n9947), .A2(n10278), .ZN(n15678) );
  NOR2_X2 U13033 ( .A1(n14205), .A2(n10279), .ZN(n14363) );
  AOI21_X1 U13034 ( .B1(n10282), .B2(n11827), .A(n11817), .ZN(n11985) );
  XNOR2_X2 U13035 ( .A(n10282), .B(n11827), .ZN(n11991) );
  NAND2_X1 U13036 ( .A1(n20243), .A2(n10285), .ZN(n10284) );
  INV_X1 U13037 ( .A(n16341), .ZN(n10287) );
  NOR2_X1 U13038 ( .A1(n10288), .A2(n10289), .ZN(n10285) );
  NAND2_X1 U13039 ( .A1(n16342), .A2(n16341), .ZN(n16340) );
  NAND2_X1 U13040 ( .A1(n10290), .A2(n10291), .ZN(n15180) );
  AND2_X1 U13041 ( .A1(n10301), .A2(n9839), .ZN(n11468) );
  NAND3_X1 U13042 ( .A1(n11256), .A2(n11440), .A3(n13871), .ZN(n11438) );
  NAND2_X1 U13043 ( .A1(n9900), .A2(n11254), .ZN(n11259) );
  AND2_X1 U13044 ( .A1(n15771), .A2(n9883), .ZN(n12968) );
  NAND2_X1 U13045 ( .A1(n15771), .A2(n9964), .ZN(n12798) );
  NAND2_X1 U13046 ( .A1(n15771), .A2(n10307), .ZN(n12422) );
  NOR2_X1 U13047 ( .A1(n10436), .A2(n10308), .ZN(n14077) );
  INV_X1 U13048 ( .A(n10679), .ZN(n13351) );
  MUX2_X1 U13049 ( .A(n10935), .B(n10938), .S(n10679), .Z(n10940) );
  INV_X1 U13050 ( .A(n11450), .ZN(n10310) );
  NAND2_X1 U13051 ( .A1(n12481), .A2(n12480), .ZN(n12801) );
  NAND2_X1 U13052 ( .A1(n11324), .A2(n11323), .ZN(n12442) );
  NAND2_X1 U13053 ( .A1(n11324), .A2(n10316), .ZN(n10315) );
  NAND2_X1 U13054 ( .A1(n12473), .A2(n10325), .ZN(n12477) );
  NAND3_X1 U13055 ( .A1(n15782), .A2(n10326), .A3(n10373), .ZN(n10325) );
  AND2_X2 U13056 ( .A1(n11529), .A2(n10328), .ZN(n11715) );
  MUX2_X1 U13057 ( .A(n10328), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n15472), .Z(n13947) );
  NAND2_X1 U13058 ( .A1(n10333), .A2(n10331), .ZN(n14387) );
  NAND3_X1 U13059 ( .A1(n13542), .A2(n10336), .A3(n9872), .ZN(n13727) );
  NAND2_X1 U13060 ( .A1(n14915), .A2(n10337), .ZN(n14858) );
  INV_X1 U13061 ( .A(n14457), .ZN(n10340) );
  NAND2_X1 U13062 ( .A1(n10340), .A2(n9936), .ZN(n15023) );
  NAND2_X1 U13063 ( .A1(n14943), .A2(n10343), .ZN(n14929) );
  NOR2_X1 U13064 ( .A1(n14833), .A2(n14834), .ZN(n12408) );
  AND2_X1 U13065 ( .A1(n12755), .A2(n20919), .ZN(n12756) );
  INV_X1 U13066 ( .A(n11216), .ZN(n11238) );
  NOR2_X1 U13067 ( .A1(n12503), .A2(n12502), .ZN(n12504) );
  CLKBUF_X1 U13068 ( .A(n15678), .Z(n15682) );
  NAND2_X1 U13069 ( .A1(n11444), .A2(n11443), .ZN(n14050) );
  NOR2_X1 U13070 ( .A1(n19384), .A2(n19412), .ZN(n19873) );
  AND2_X1 U13071 ( .A1(n19384), .A2(n19391), .ZN(n10955) );
  INV_X1 U13072 ( .A(n11441), .ZN(n11444) );
  AOI21_X1 U13073 ( .B1(n10646), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A(
        n10449), .ZN(n10450) );
  NAND2_X1 U13074 ( .A1(n10975), .A2(n10951), .ZN(n10952) );
  NOR2_X1 U13075 ( .A1(n11141), .A2(n11140), .ZN(n11142) );
  AND2_X1 U13076 ( .A1(n19391), .A2(n19419), .ZN(n19879) );
  NAND2_X1 U13077 ( .A1(n10968), .A2(n19391), .ZN(n10969) );
  INV_X1 U13078 ( .A(n19391), .ZN(n10951) );
  AND2_X1 U13079 ( .A1(n19420), .A2(n19419), .ZN(n19904) );
  NAND2_X1 U13080 ( .A1(n19420), .A2(n14287), .ZN(n15694) );
  NAND2_X1 U13081 ( .A1(n10938), .A2(n10937), .ZN(n10939) );
  NAND2_X1 U13082 ( .A1(n10937), .A2(n19274), .ZN(n19229) );
  AOI22_X1 U13083 ( .A1(n12043), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12723), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11563) );
  OR3_X1 U13084 ( .A1(n13544), .A2(n13543), .A3(n16195), .ZN(n13545) );
  NOR2_X1 U13085 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n13554), .ZN(
        n11529) );
  AOI22_X1 U13086 ( .A1(n10649), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n10648), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10470) );
  AOI22_X1 U13087 ( .A1(n9847), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n10645), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10471) );
  AOI21_X1 U13088 ( .B1(n12038), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A(
        n11572), .ZN(n11577) );
  NAND2_X1 U13089 ( .A1(n13727), .A2(n11999), .ZN(n13853) );
  AOI22_X1 U13090 ( .A1(n13678), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n10644), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10643) );
  NAND2_X1 U13091 ( .A1(n13678), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n10628) );
  NAND2_X1 U13092 ( .A1(n13678), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n10597) );
  AND2_X2 U13093 ( .A1(n11528), .A2(n11529), .ZN(n11697) );
  AOI22_X1 U13094 ( .A1(n11692), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n11715), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11581) );
  INV_X1 U13095 ( .A(n10645), .ZN(n14626) );
  INV_X1 U13096 ( .A(n17957), .ZN(n13160) );
  NAND2_X1 U13097 ( .A1(n14624), .A2(n10426), .ZN(n10351) );
  NAND2_X1 U13098 ( .A1(n10425), .A2(n14624), .ZN(n10352) );
  NOR2_X1 U13099 ( .A1(n12509), .A2(n12513), .ZN(n12631) );
  AND2_X1 U13100 ( .A1(n10938), .A2(n19420), .ZN(n10353) );
  AND2_X1 U13101 ( .A1(n10887), .A2(n10886), .ZN(n14280) );
  INV_X1 U13102 ( .A(n14280), .ZN(n14206) );
  AND2_X1 U13103 ( .A1(n10987), .A2(n10986), .ZN(n10354) );
  OR2_X1 U13104 ( .A1(n17283), .A2(n13127), .ZN(n10355) );
  OR2_X1 U13105 ( .A1(n13160), .A2(n17694), .ZN(n10356) );
  INV_X1 U13106 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n13867) );
  INV_X1 U13107 ( .A(n13910), .ZN(n20189) );
  NAND3_X1 U13108 ( .A1(n10499), .A2(n10498), .A3(n10497), .ZN(n10357) );
  AND2_X1 U13109 ( .A1(n10782), .A2(n10781), .ZN(n13704) );
  AND3_X1 U13110 ( .A1(n10548), .A2(n10547), .A3(n10546), .ZN(n10358) );
  OR2_X1 U13111 ( .A1(n9845), .A2(n16390), .ZN(n10359) );
  AND3_X1 U13112 ( .A1(n13062), .A2(n13061), .A3(n13060), .ZN(n10360) );
  AND2_X1 U13113 ( .A1(n10988), .A2(n10354), .ZN(n10361) );
  AND3_X1 U13114 ( .A1(n10353), .A2(n10970), .A3(n10969), .ZN(n10362) );
  AND4_X1 U13115 ( .A1(n12985), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n12984), .A4(n12797), .ZN(n10365) );
  INV_X2 U13116 ( .A(n20075), .ZN(n19994) );
  NAND2_X1 U13117 ( .A1(n13349), .A2(n13386), .ZN(n15667) );
  OR2_X1 U13118 ( .A1(n16897), .A2(n17805), .ZN(n10366) );
  AND3_X1 U13119 ( .A1(n10470), .A2(n10469), .A3(n10468), .ZN(n10367) );
  AND2_X1 U13120 ( .A1(n15105), .A2(BUF1_REG_30__SCAN_IN), .ZN(n10368) );
  INV_X2 U13121 ( .A(n19025), .ZN(n18960) );
  NOR2_X1 U13122 ( .A1(n11979), .A2(n20999), .ZN(n12025) );
  AND2_X1 U13123 ( .A1(n12976), .A2(n12974), .ZN(n10369) );
  AND2_X1 U13124 ( .A1(n20769), .A2(n12411), .ZN(n16325) );
  NAND2_X1 U13125 ( .A1(n11816), .A2(n16201), .ZN(n11929) );
  AND2_X1 U13126 ( .A1(n10472), .A2(n10471), .ZN(n10370) );
  OR2_X1 U13127 ( .A1(n18994), .A2(n18046), .ZN(n19021) );
  INV_X1 U13128 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n20036) );
  AND2_X1 U13129 ( .A1(n12414), .A2(n20999), .ZN(n20280) );
  INV_X1 U13130 ( .A(n20280), .ZN(n20256) );
  INV_X1 U13131 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n13004) );
  OR2_X1 U13132 ( .A1(n14380), .A2(n14379), .ZN(n10371) );
  INV_X1 U13133 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n13478) );
  NOR2_X1 U13134 ( .A1(n17806), .A2(n17895), .ZN(n18031) );
  AND2_X1 U13135 ( .A1(n10627), .A2(n10626), .ZN(n10372) );
  INV_X1 U13136 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15990) );
  OR2_X1 U13137 ( .A1(n13630), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n10374) );
  INV_X2 U13138 ( .A(n17426), .ZN(n17418) );
  NAND2_X2 U13139 ( .A1(n15090), .A2(n13018), .ZN(n15118) );
  INV_X1 U13140 ( .A(n15118), .ZN(n13019) );
  NOR2_X1 U13141 ( .A1(n20732), .A2(n20695), .ZN(n10375) );
  AND2_X1 U13142 ( .A1(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n10376) );
  NOR2_X1 U13143 ( .A1(n20732), .A2(n20845), .ZN(n10377) );
  INV_X1 U13144 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n20061) );
  INV_X1 U13145 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n14298) );
  INV_X1 U13146 ( .A(n14705), .ZN(n14703) );
  OR2_X1 U13147 ( .A1(n14686), .A2(n14685), .ZN(n10378) );
  INV_X1 U13148 ( .A(n15771), .ZN(n15798) );
  INV_X1 U13149 ( .A(n12742), .ZN(n12847) );
  AND2_X1 U13150 ( .A1(n14387), .A2(n14494), .ZN(n10379) );
  OR2_X1 U13151 ( .A1(n19042), .A2(n9839), .ZN(n16553) );
  INV_X1 U13152 ( .A(n16553), .ZN(n12840) );
  OR2_X1 U13153 ( .A1(n12795), .A2(n16553), .ZN(n10380) );
  AND2_X1 U13154 ( .A1(n13519), .A2(n11666), .ZN(n10381) );
  NAND2_X1 U13155 ( .A1(n11188), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11189) );
  AOI22_X1 U13156 ( .A1(n11684), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n12723), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11534) );
  AND2_X1 U13157 ( .A1(n9819), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11572) );
  NAND2_X1 U13158 ( .A1(n13678), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n10468) );
  OR2_X1 U13159 ( .A1(n11801), .A2(n11800), .ZN(n11887) );
  INV_X1 U13160 ( .A(n11833), .ZN(n11727) );
  AND2_X1 U13161 ( .A1(n10968), .A2(n10971), .ZN(n10941) );
  NOR2_X1 U13162 ( .A1(n11535), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11536) );
  INV_X1 U13163 ( .A(n13774), .ZN(n11835) );
  NAND2_X1 U13164 ( .A1(n12849), .A2(n13774), .ZN(n11646) );
  INV_X1 U13165 ( .A(n11765), .ZN(n11705) );
  AND2_X1 U13166 ( .A1(n10648), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n10449) );
  AND2_X1 U13167 ( .A1(n9846), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10632) );
  AOI22_X1 U13168 ( .A1(n12038), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n9820), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11545) );
  INV_X1 U13169 ( .A(n14963), .ZN(n12179) );
  OR2_X1 U13170 ( .A1(n9844), .A2(n15392), .ZN(n11909) );
  INV_X1 U13171 ( .A(n11929), .ZN(n11886) );
  NOR2_X1 U13172 ( .A1(n11757), .A2(n11756), .ZN(n11846) );
  AND2_X1 U13173 ( .A1(n10543), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n10584) );
  NAND2_X1 U13174 ( .A1(n11153), .A2(n11137), .ZN(n11139) );
  INV_X1 U13175 ( .A(n10673), .ZN(n10530) );
  AND2_X1 U13176 ( .A1(n14706), .A2(n14703), .ZN(n14707) );
  AND2_X1 U13177 ( .A1(n15673), .A2(n14643), .ZN(n14644) );
  INV_X1 U13178 ( .A(n12987), .ZN(n12988) );
  NAND2_X1 U13179 ( .A1(n10543), .A2(P2_EBX_REG_2__SCAN_IN), .ZN(n10516) );
  OR2_X1 U13180 ( .A1(n10908), .A2(n19934), .ZN(n10692) );
  INV_X1 U13181 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n11383) );
  INV_X1 U13182 ( .A(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n13127) );
  NAND2_X1 U13183 ( .A1(n10381), .A2(n11677), .ZN(n11708) );
  INV_X1 U13184 ( .A(n14977), .ZN(n12089) );
  NAND2_X1 U13185 ( .A1(n12763), .A2(n11642), .ZN(n13514) );
  AND2_X1 U13186 ( .A1(n12369), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12370) );
  NAND2_X1 U13187 ( .A1(n15466), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12717) );
  NOR2_X1 U13188 ( .A1(n12194), .A2(n14951), .ZN(n12210) );
  NAND2_X1 U13189 ( .A1(n12102), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n12140) );
  INV_X1 U13190 ( .A(n12025), .ZN(n12005) );
  NAND2_X1 U13191 ( .A1(n13853), .A2(n13852), .ZN(n13851) );
  OAI21_X1 U13192 ( .B1(n16302), .B2(n11912), .A(n15174), .ZN(n11913) );
  AND2_X1 U13193 ( .A1(n15244), .A2(n15242), .ZN(n15221) );
  INV_X1 U13194 ( .A(n13464), .ZN(n13465) );
  OAI21_X1 U13195 ( .B1(n11959), .B2(n11730), .A(n11729), .ZN(n11827) );
  AND2_X1 U13196 ( .A1(n10714), .A2(n10545), .ZN(n11276) );
  INV_X1 U13197 ( .A(n11022), .ZN(n11116) );
  NAND2_X1 U13198 ( .A1(n13568), .A2(n13567), .ZN(n13569) );
  AOI22_X1 U13199 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n9859), .B1(
        n10647), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n10642) );
  INV_X1 U13200 ( .A(n15684), .ZN(n14561) );
  INV_X1 U13201 ( .A(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n12790) );
  OAI22_X1 U13202 ( .A1(n11013), .A2(n10977), .B1(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n11021), .ZN(n10980) );
  OR2_X1 U13203 ( .A1(n14267), .A2(n11450), .ZN(n11451) );
  AND2_X1 U13204 ( .A1(n10936), .A2(n19420), .ZN(n10654) );
  INV_X1 U13205 ( .A(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n17383) );
  INV_X1 U13206 ( .A(n18804), .ZN(n16626) );
  OAI21_X1 U13207 ( .B1(n17852), .B2(n17755), .A(n13157), .ZN(n13158) );
  INV_X1 U13208 ( .A(n12543), .ZN(n12544) );
  INV_X1 U13209 ( .A(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n17201) );
  INV_X1 U13210 ( .A(n11708), .ZN(n11709) );
  AND4_X1 U13211 ( .A1(n11603), .A2(n11602), .A3(n11601), .A4(n11600), .ZN(
        n11620) );
  AOI21_X1 U13212 ( .B1(n15122), .B2(n12847), .A(n12746), .ZN(n13015) );
  NOR2_X1 U13213 ( .A1(n12140), .A2(n14983), .ZN(n12145) );
  AND2_X1 U13214 ( .A1(n20999), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n12747) );
  OR2_X1 U13215 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n12742) );
  INV_X1 U13216 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20387) );
  INV_X1 U13217 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20598) );
  OR2_X1 U13218 ( .A1(n9853), .A2(n21000), .ZN(n20628) );
  NAND2_X1 U13219 ( .A1(n11975), .A2(n11974), .ZN(n11976) );
  NAND2_X1 U13220 ( .A1(n10958), .A2(n10972), .ZN(n14104) );
  INV_X1 U13221 ( .A(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n15756) );
  INV_X1 U13222 ( .A(n10935), .ZN(n10960) );
  NAND2_X1 U13223 ( .A1(n16157), .A2(n20064), .ZN(n10972) );
  OR2_X1 U13224 ( .A1(n13569), .A2(n13589), .ZN(n13588) );
  INV_X1 U13225 ( .A(n10908), .ZN(n12818) );
  AND2_X1 U13226 ( .A1(n11030), .A2(n11029), .ZN(n13601) );
  AND2_X1 U13227 ( .A1(n16054), .A2(n11462), .ZN(n16004) );
  OR2_X1 U13228 ( .A1(n15615), .A2(n11254), .ZN(n11322) );
  INV_X1 U13229 ( .A(n14105), .ZN(n13379) );
  AND2_X2 U13230 ( .A1(n11178), .A2(n19354), .ZN(n11225) );
  INV_X1 U13231 ( .A(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n21208) );
  AOI21_X1 U13232 ( .B1(n17327), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A(
        n13069), .ZN(n13070) );
  INV_X1 U13233 ( .A(n17776), .ZN(n17806) );
  NOR2_X1 U13234 ( .A1(n16627), .A2(n16626), .ZN(n16628) );
  NOR2_X1 U13235 ( .A1(n13152), .A2(n18177), .ZN(n17853) );
  NOR2_X1 U13236 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n18009), .ZN(
        n18008) );
  NOR4_X1 U13237 ( .A1(n12547), .A2(n12546), .A3(n12545), .A4(n12544), .ZN(
        n12548) );
  INV_X1 U13238 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n14890) );
  INV_X1 U13239 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n14983) );
  INV_X1 U13240 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n14392) );
  OR2_X1 U13241 ( .A1(n21008), .A2(n12943), .ZN(n20117) );
  AND2_X1 U13242 ( .A1(n20151), .A2(n20117), .ZN(n14958) );
  OR2_X1 U13243 ( .A1(n14002), .A2(n20303), .ZN(n15103) );
  OAI21_X1 U13244 ( .B1(n13460), .B2(n12767), .A(n13768), .ZN(n12768) );
  INV_X1 U13245 ( .A(n12416), .ZN(n12417) );
  INV_X1 U13246 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n15167) );
  NAND2_X1 U13247 ( .A1(n12211), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n12246) );
  NOR2_X1 U13248 ( .A1(n12162), .A2(n16258), .ZN(n12180) );
  NOR2_X1 U13249 ( .A1(n12079), .A2(n20104), .ZN(n12083) );
  AND3_X1 U13250 ( .A1(n12053), .A2(n12052), .A3(n12051), .ZN(n14388) );
  NOR2_X1 U13251 ( .A1(n11919), .A2(n11920), .ZN(n13791) );
  AND2_X1 U13252 ( .A1(n12897), .A2(n12896), .ZN(n15029) );
  AND2_X1 U13253 ( .A1(n20080), .A2(n20310), .ZN(n12414) );
  NAND2_X1 U13254 ( .A1(n16400), .A2(n20275), .ZN(n20258) );
  AND2_X1 U13255 ( .A1(n13783), .A2(n13782), .ZN(n15284) );
  INV_X1 U13256 ( .A(n11991), .ZN(n20307) );
  OR2_X1 U13257 ( .A1(n20593), .A2(n13972), .ZN(n20496) );
  AND2_X1 U13258 ( .A1(n20796), .A2(n20353), .ZN(n20663) );
  INV_X1 U13259 ( .A(n13838), .ZN(n20799) );
  INV_X1 U13260 ( .A(n20769), .ZN(n20848) );
  NOR2_X1 U13261 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n16442), .ZN(n21002) );
  NOR2_X1 U13262 ( .A1(n19925), .A2(n20063), .ZN(n14113) );
  INV_X1 U13263 ( .A(n10972), .ZN(n13686) );
  AND2_X1 U13264 ( .A1(n11119), .A2(n11118), .ZN(n12487) );
  AND2_X1 U13265 ( .A1(n14658), .A2(n14657), .ZN(n14663) );
  AND2_X1 U13266 ( .A1(n10802), .A2(n10801), .ZN(n13814) );
  AND3_X1 U13267 ( .A1(n10662), .A2(n10661), .A3(n10660), .ZN(n14037) );
  OAI21_X1 U13268 ( .B1(n13284), .B2(n13283), .A(P2_ADDRESS_REG_29__SCAN_IN), 
        .ZN(n13285) );
  INV_X1 U13269 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n14424) );
  INV_X1 U13270 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15922) );
  AND3_X1 U13271 ( .A1(n10785), .A2(n10784), .A3(n10783), .ZN(n14172) );
  AND2_X1 U13272 ( .A1(n14054), .A2(n11510), .ZN(n16574) );
  XNOR2_X1 U13273 ( .A(n11436), .B(n13867), .ZN(n13871) );
  NAND2_X1 U13274 ( .A1(n11505), .A2(n11468), .ZN(n19355) );
  INV_X1 U13275 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n20013) );
  NAND2_X1 U13276 ( .A1(n20034), .A2(n20013), .ZN(n20002) );
  AND2_X1 U13277 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n13584) );
  OR2_X1 U13278 ( .A1(n14315), .A2(n20002), .ZN(n19579) );
  INV_X1 U13279 ( .A(n19720), .ZN(n19717) );
  OR2_X1 U13280 ( .A1(n16589), .A2(n14297), .ZN(n14299) );
  OR2_X1 U13281 ( .A1(n19782), .A2(n20001), .ZN(n19370) );
  INV_X1 U13282 ( .A(n13188), .ZN(n13193) );
  NOR2_X1 U13283 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n16903), .ZN(n16887) );
  INV_X1 U13284 ( .A(n16876), .ZN(n16934) );
  INV_X1 U13285 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n17069) );
  INV_X1 U13286 ( .A(P3_EBX_REG_22__SCAN_IN), .ZN(n17118) );
  INV_X1 U13287 ( .A(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n17308) );
  INV_X1 U13288 ( .A(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n21308) );
  NOR2_X1 U13289 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n19027), .ZN(n17892) );
  NAND2_X1 U13290 ( .A1(n17892), .A2(n18045), .ZN(n17776) );
  INV_X1 U13291 ( .A(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n17804) );
  OAI21_X1 U13292 ( .B1(n16629), .B2(n17551), .A(n16628), .ZN(n16633) );
  INV_X1 U13293 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n17828) );
  INV_X1 U13294 ( .A(n17836), .ZN(n18161) );
  NOR2_X1 U13295 ( .A1(n17957), .A2(n17960), .ZN(n17956) );
  INV_X1 U13296 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n13118) );
  NOR2_X1 U13297 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18377), .ZN(n18720) );
  INV_X1 U13298 ( .A(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n21306) );
  AOI22_X1 U13299 ( .A1(n18808), .A2(n18244), .B1(n18800), .B2(n18804), .ZN(
        n18811) );
  NAND2_X1 U13300 ( .A1(n13396), .A2(n13637), .ZN(n21008) );
  OAI21_X1 U13301 ( .B1(n15274), .B2(n20124), .A(n12964), .ZN(n12965) );
  OR2_X1 U13302 ( .A1(n12319), .A2(n14890), .ZN(n12327) );
  XNOR2_X1 U13303 ( .A(n12846), .B(n12956), .ZN(n13837) );
  INV_X1 U13304 ( .A(n20151), .ZN(n20137) );
  AND2_X1 U13305 ( .A1(n13809), .A2(n12768), .ZN(n16293) );
  INV_X1 U13306 ( .A(n15076), .ZN(n20342) );
  INV_X1 U13307 ( .A(n15071), .ZN(n20352) );
  INV_X1 U13308 ( .A(n13809), .ZN(n20224) );
  AND2_X1 U13309 ( .A1(n14929), .A2(n15006), .ZN(n16296) );
  AND2_X1 U13310 ( .A1(n12026), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12032) );
  OR2_X1 U13311 ( .A1(n20248), .A2(n12412), .ZN(n15228) );
  AND3_X1 U13312 ( .A1(n13791), .A2(n16193), .A3(n11978), .ZN(n20248) );
  AND2_X1 U13313 ( .A1(n15378), .A2(n15279), .ZN(n15340) );
  AND2_X1 U13314 ( .A1(n15431), .A2(n15278), .ZN(n15378) );
  INV_X1 U13315 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n15453) );
  INV_X1 U13316 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n16390) );
  NAND2_X1 U13317 ( .A1(n15366), .A2(n15385), .ZN(n15431) );
  AND2_X1 U13318 ( .A1(n13795), .A2(n13772), .ZN(n20282) );
  OR2_X1 U13319 ( .A1(n16400), .A2(n20289), .ZN(n20276) );
  INV_X1 U13320 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13561) );
  OAI22_X1 U13321 ( .A1(n20322), .A2(n20321), .B1(n20601), .B2(n20320), .ZN(
        n20354) );
  INV_X1 U13322 ( .A(n20418), .ZN(n20375) );
  OAI22_X1 U13323 ( .A1(n20391), .A2(n20390), .B1(n20601), .B2(n20527), .ZN(
        n20414) );
  NAND2_X1 U13324 ( .A1(n9853), .A2(n20307), .ZN(n20703) );
  NAND2_X1 U13325 ( .A1(n20594), .A2(n20593), .ZN(n20425) );
  INV_X1 U13326 ( .A(n20478), .ZN(n20488) );
  OAI22_X1 U13327 ( .A1(n20529), .A2(n20528), .B1(n20527), .B2(n20796), .ZN(
        n20556) );
  INV_X1 U13328 ( .A(n20496), .ZN(n20570) );
  INV_X1 U13329 ( .A(n20725), .ZN(n20595) );
  OAI211_X1 U13330 ( .C1(n20666), .C2(n20665), .A(n20664), .B(n20663), .ZN(
        n20691) );
  NAND2_X1 U13331 ( .A1(n9853), .A2(n11991), .ZN(n20652) );
  INV_X1 U13332 ( .A(n20469), .ZN(n20353) );
  NOR2_X2 U13333 ( .A1(n20855), .A2(n20725), .ZN(n20790) );
  INV_X1 U13334 ( .A(n20631), .ZN(n20766) );
  INV_X1 U13335 ( .A(n20805), .ZN(n20837) );
  INV_X1 U13336 ( .A(n20741), .ZN(n20852) );
  INV_X1 U13337 ( .A(n20750), .ZN(n20875) );
  INV_X1 U13338 ( .A(n20684), .ZN(n20893) );
  INV_X1 U13339 ( .A(n20855), .ZN(n20795) );
  NOR2_X1 U13340 ( .A1(n16442), .A2(n20999), .ZN(n13963) );
  INV_X1 U13341 ( .A(n21010), .ZN(n20919) );
  INV_X1 U13342 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n20928) );
  INV_X1 U13343 ( .A(n20970), .ZN(n20977) );
  OR2_X1 U13344 ( .A1(n14789), .A2(n19197), .ZN(n11129) );
  AND2_X1 U13345 ( .A1(n13527), .A2(n14128), .ZN(n19183) );
  OR2_X1 U13346 ( .A1(n11402), .A2(n10590), .ZN(n14115) );
  INV_X1 U13347 ( .A(n15694), .ZN(n15685) );
  OR2_X1 U13348 ( .A1(n19221), .A2(n13390), .ZN(n19266) );
  INV_X1 U13349 ( .A(n13655), .ZN(n13526) );
  AND2_X1 U13350 ( .A1(n16559), .A2(n13346), .ZN(n16550) );
  NOR2_X1 U13351 ( .A1(n12795), .A2(n19363), .ZN(n12503) );
  OR2_X1 U13352 ( .A1(n15953), .A2(n12497), .ZN(n15930) );
  AND2_X1 U13353 ( .A1(n15689), .A2(n14433), .ZN(n16486) );
  INV_X1 U13354 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n16034) );
  INV_X1 U13355 ( .A(n19327), .ZN(n19347) );
  AND2_X1 U13356 ( .A1(n14112), .A2(n20060), .ZN(n20049) );
  INV_X1 U13357 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n19348) );
  XNOR2_X1 U13358 ( .A(n13573), .B(n13574), .ZN(n20029) );
  INV_X1 U13359 ( .A(n19372), .ZN(n19421) );
  NOR2_X2 U13360 ( .A1(n19667), .A2(n19568), .ZN(n19454) );
  NOR2_X1 U13361 ( .A1(n19667), .A2(n19615), .ZN(n19487) );
  OAI21_X1 U13362 ( .B1(n19498), .B2(n19497), .A(n19496), .ZN(n19515) );
  NAND2_X1 U13363 ( .A1(n14320), .A2(n14319), .ZN(n19536) );
  OAI21_X1 U13364 ( .B1(n19539), .B2(n19579), .A(n19578), .ZN(n19599) );
  NOR2_X2 U13365 ( .A1(n19615), .A2(n20001), .ZN(n19662) );
  INV_X1 U13366 ( .A(n19697), .ZN(n19680) );
  INV_X1 U13367 ( .A(n19683), .ZN(n19710) );
  AND2_X1 U13368 ( .A1(n19723), .A2(n19721), .ZN(n19745) );
  NOR2_X1 U13369 ( .A1(n19782), .A2(n20004), .ZN(n19769) );
  NOR2_X1 U13370 ( .A1(n19776), .A2(n19775), .ZN(n19797) );
  AND2_X1 U13371 ( .A1(n14299), .A2(n14298), .ZN(n19861) );
  INV_X1 U13372 ( .A(n19817), .ZN(n19856) );
  INV_X1 U13373 ( .A(n19829), .ZN(n19880) );
  INV_X1 U13374 ( .A(n19841), .ZN(n19898) );
  NAND2_X1 U13375 ( .A1(n20034), .A2(n13362), .ZN(n16225) );
  INV_X1 U13376 ( .A(n20069), .ZN(n19925) );
  INV_X1 U13377 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n19933) );
  NAND2_X1 U13378 ( .A1(n17631), .A2(n18801), .ZN(n17051) );
  INV_X1 U13379 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n17120) );
  NOR2_X1 U13380 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n16874), .ZN(n16862) );
  NOR2_X1 U13381 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n16922), .ZN(n16912) );
  NOR3_X1 U13382 ( .A1(n17104), .A2(n16942), .A3(n16827), .ZN(n16927) );
  NOR2_X1 U13383 ( .A1(n18856), .A2(n13305), .ZN(n17083) );
  INV_X1 U13384 ( .A(n17102), .ZN(n17070) );
  NAND4_X1 U13385 ( .A1(n18316), .A2(n17051), .A3(n18873), .A4(n18862), .ZN(
        n17114) );
  INV_X1 U13386 ( .A(P3_EBX_REG_24__SCAN_IN), .ZN(n21285) );
  INV_X1 U13387 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n16904) );
  INV_X1 U13388 ( .A(P3_EBX_REG_4__SCAN_IN), .ZN(n12619) );
  NOR3_X1 U13389 ( .A1(n18413), .A2(n17509), .A3(n17636), .ZN(n17501) );
  NOR2_X2 U13390 ( .A1(n17433), .A2(n17571), .ZN(n17508) );
  INV_X2 U13391 ( .A(n13051), .ZN(n17378) );
  INV_X1 U13392 ( .A(n17629), .ZN(n17584) );
  INV_X1 U13393 ( .A(n17892), .ZN(n18046) );
  OAI211_X1 U13394 ( .C1(n19012), .C2(n18858), .A(n17632), .B(n17631), .ZN(
        n17677) );
  INV_X1 U13395 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n18094) );
  NOR2_X1 U13396 ( .A1(n18994), .A2(n18041), .ZN(n17895) );
  INV_X1 U13397 ( .A(n18418), .ZN(n18748) );
  INV_X1 U13398 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n18040) );
  INV_X1 U13399 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n17693) );
  INV_X1 U13400 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n19017) );
  NOR2_X1 U13401 ( .A1(n17729), .A2(n18188), .ZN(n17741) );
  INV_X1 U13402 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n18115) );
  NOR2_X1 U13403 ( .A1(n18250), .A2(n18237), .ZN(n18228) );
  NOR2_X2 U13404 ( .A1(n18387), .A2(n18276), .ZN(n18244) );
  INV_X1 U13405 ( .A(n18350), .ZN(n18344) );
  INV_X1 U13406 ( .A(n18359), .ZN(n18349) );
  NOR3_X1 U13407 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(P3_STATE2_REG_3__SCAN_IN), .A3(n19013), .ZN(n16145) );
  NOR2_X1 U13408 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18967), .ZN(
        n18988) );
  INV_X1 U13409 ( .A(n18741), .ZN(n18721) );
  INV_X1 U13410 ( .A(n18422), .ZN(n18482) );
  INV_X1 U13411 ( .A(n18509), .ZN(n18550) );
  INV_X1 U13412 ( .A(n18507), .ZN(n18572) );
  INV_X1 U13413 ( .A(n18532), .ZN(n18594) );
  INV_X1 U13414 ( .A(n18554), .ZN(n18615) );
  INV_X1 U13415 ( .A(n18598), .ZN(n18663) );
  INV_X1 U13416 ( .A(n18622), .ZN(n18685) );
  INV_X1 U13417 ( .A(n18644), .ZN(n18709) );
  INV_X1 U13418 ( .A(n18667), .ZN(n18737) );
  NOR2_X1 U13419 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n19017), .ZN(n18870) );
  INV_X1 U13420 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n18897) );
  INV_X2 U13421 ( .A(n14302), .ZN(n14303) );
  INV_X1 U13422 ( .A(n21008), .ZN(n13840) );
  INV_X1 U13423 ( .A(n12965), .ZN(n12966) );
  NAND2_X1 U13424 ( .A1(n12955), .A2(n12939), .ZN(n20124) );
  OR2_X1 U13425 ( .A1(n13837), .A2(n13835), .ZN(n14988) );
  INV_X1 U13426 ( .A(n20154), .ZN(n20143) );
  OR2_X1 U13427 ( .A1(n14002), .A2(n20305), .ZN(n16299) );
  AND2_X1 U13428 ( .A1(n13717), .A2(n13716), .ZN(n15071) );
  AND2_X1 U13429 ( .A1(n14012), .A2(n14011), .ZN(n20328) );
  NAND2_X1 U13430 ( .A1(n20187), .A2(n11644), .ZN(n13912) );
  INV_X1 U13431 ( .A(n20187), .ZN(n20208) );
  NOR2_X1 U13432 ( .A1(n13637), .A2(n12756), .ZN(n13808) );
  NAND2_X1 U13433 ( .A1(n13808), .A2(n16201), .ZN(n13809) );
  OAI21_X1 U13434 ( .B1(n14932), .B2(n14931), .A(n14930), .ZN(n15207) );
  NAND2_X1 U13435 ( .A1(n15228), .A2(n13537), .ZN(n20252) );
  INV_X1 U13436 ( .A(n16325), .ZN(n20306) );
  XNOR2_X1 U13437 ( .A(n11918), .B(n15327), .ZN(n15334) );
  INV_X1 U13438 ( .A(n20282), .ZN(n20292) );
  INV_X1 U13439 ( .A(n20278), .ZN(n20293) );
  INV_X1 U13440 ( .A(n15431), .ZN(n16421) );
  INV_X1 U13441 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n20267) );
  INV_X1 U13442 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20767) );
  AND2_X1 U13443 ( .A1(n13476), .A2(n13470), .ZN(n15484) );
  OR2_X1 U13444 ( .A1(n20425), .A2(n20725), .ZN(n20378) );
  OR2_X1 U13445 ( .A1(n20425), .A2(n20631), .ZN(n20418) );
  OR2_X1 U13446 ( .A1(n20425), .A2(n20703), .ZN(n20465) );
  OR2_X1 U13447 ( .A1(n20425), .A2(n20652), .ZN(n20459) );
  NAND2_X1 U13448 ( .A1(n20570), .A2(n20595), .ZN(n20519) );
  NAND2_X1 U13449 ( .A1(n20570), .A2(n20766), .ZN(n20560) );
  NAND2_X1 U13450 ( .A1(n20570), .A2(n20794), .ZN(n20592) );
  NAND2_X1 U13451 ( .A1(n20596), .A2(n20595), .ZN(n20651) );
  AOI22_X1 U13452 ( .A1(n20661), .A2(n20665), .B1(n20658), .B2(n20657), .ZN(
        n20694) );
  OR2_X1 U13453 ( .A1(n20704), .A2(n20652), .ZN(n20724) );
  AOI22_X1 U13454 ( .A1(n20736), .A2(n20733), .B1(n20731), .B2(n20730), .ZN(
        n20765) );
  NAND2_X1 U13455 ( .A1(n20795), .A2(n20766), .ZN(n20805) );
  NAND2_X1 U13456 ( .A1(n20795), .A2(n20794), .ZN(n20908) );
  INV_X1 U13457 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n20738) );
  AOI21_X1 U13458 ( .B1(P1_STATE_REG_0__SCAN_IN), .B2(n20918), .A(n21013), 
        .ZN(n20989) );
  INV_X1 U13459 ( .A(P1_ADDRESS_REG_2__SCAN_IN), .ZN(n20931) );
  NAND2_X1 U13460 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n21013), .ZN(n20970) );
  OR2_X1 U13461 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n20077), .ZN(n20997) );
  INV_X1 U13462 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n21257) );
  INV_X1 U13463 ( .A(n15624), .ZN(n15494) );
  OR2_X1 U13464 ( .A1(n11128), .A2(n11127), .ZN(n19197) );
  INV_X1 U13465 ( .A(n19186), .ZN(n19202) );
  INV_X1 U13466 ( .A(n19210), .ZN(n19181) );
  INV_X1 U13467 ( .A(n19183), .ZN(n19200) );
  INV_X1 U13468 ( .A(n19175), .ZN(n19214) );
  AND2_X1 U13469 ( .A1(n19258), .A2(n19229), .ZN(n19264) );
  AND2_X1 U13470 ( .A1(n13387), .A2(n13386), .ZN(n19274) );
  NAND2_X1 U13471 ( .A1(n19310), .A2(n13363), .ZN(n19276) );
  INV_X1 U13472 ( .A(n19310), .ZN(n19308) );
  INV_X1 U13473 ( .A(n13447), .ZN(n13655) );
  NAND2_X1 U13474 ( .A1(n12841), .A2(n12840), .ZN(n12842) );
  INV_X1 U13475 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n16506) );
  INV_X1 U13476 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n16529) );
  INV_X1 U13477 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n16558) );
  INV_X1 U13478 ( .A(n19315), .ZN(n16545) );
  INV_X1 U13479 ( .A(n11520), .ZN(n11521) );
  INV_X1 U13480 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n16491) );
  INV_X1 U13481 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n16570) );
  NAND2_X1 U13482 ( .A1(n11505), .A2(n20049), .ZN(n19356) );
  INV_X1 U13483 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20023) );
  AOI21_X1 U13484 ( .B1(n19371), .B2(n19375), .A(n19369), .ZN(n19429) );
  INV_X1 U13485 ( .A(n19487), .ZN(n19462) );
  OR2_X1 U13486 ( .A1(n19568), .A2(n20004), .ZN(n19519) );
  INV_X1 U13487 ( .A(n19536), .ZN(n19523) );
  OR2_X1 U13488 ( .A1(n19568), .A2(n19781), .ZN(n19561) );
  AND2_X1 U13489 ( .A1(n19577), .A2(n19576), .ZN(n19587) );
  OR2_X1 U13490 ( .A1(n19615), .A2(n19781), .ZN(n19603) );
  INV_X1 U13491 ( .A(n19604), .ZN(n19634) );
  OAI21_X1 U13492 ( .B1(n19642), .B2(P2_STATE2_REG_2__SCAN_IN), .A(n19641), 
        .ZN(n19666) );
  OR2_X1 U13493 ( .A1(n19782), .A2(n19667), .ZN(n19683) );
  INV_X1 U13494 ( .A(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n19713) );
  INV_X1 U13495 ( .A(n19737), .ZN(n19749) );
  INV_X1 U13496 ( .A(n19875), .ZN(n19755) );
  INV_X1 U13497 ( .A(n19899), .ZN(n19766) );
  INV_X1 U13498 ( .A(n19760), .ZN(n19801) );
  AOI21_X1 U13499 ( .B1(n19809), .B2(n19813), .A(n19807), .ZN(n19850) );
  INV_X1 U13500 ( .A(n19830), .ZN(n19890) );
  OR2_X1 U13501 ( .A1(n10928), .A2(n20034), .ZN(n19040) );
  INV_X1 U13502 ( .A(n20000), .ZN(n19914) );
  OAI21_X1 U13503 ( .B1(n21257), .B2(n19922), .A(n19919), .ZN(n20000) );
  NOR2_X1 U13504 ( .A1(n18864), .A2(n18802), .ZN(n17631) );
  INV_X1 U13505 ( .A(n13232), .ZN(n16733) );
  INV_X1 U13506 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n17322) );
  NAND2_X1 U13507 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n17114), .ZN(n17102) );
  INV_X1 U13508 ( .A(P3_EBX_REG_3__SCAN_IN), .ZN(n17079) );
  NOR2_X1 U13509 ( .A1(n17127), .A2(n17126), .ZN(n17154) );
  NOR2_X1 U13510 ( .A1(n16950), .A2(n16137), .ZN(n17301) );
  INV_X1 U13511 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n17401) );
  AND2_X1 U13512 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n17528), .ZN(n17531) );
  INV_X1 U13513 ( .A(n17537), .ZN(n17541) );
  AND2_X1 U13514 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(n17566), .ZN(n17562) );
  INV_X1 U13515 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n17583) );
  NAND2_X1 U13516 ( .A1(n17584), .A2(n18378), .ZN(n17604) );
  INV_X1 U13517 ( .A(n17602), .ZN(n17609) );
  INV_X1 U13518 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n21127) );
  INV_X1 U13519 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n17659) );
  INV_X1 U13520 ( .A(n17685), .ZN(n17680) );
  INV_X1 U13521 ( .A(n17849), .ZN(n17864) );
  INV_X1 U13522 ( .A(n17963), .ZN(n17889) );
  INV_X1 U13523 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n18269) );
  INV_X1 U13524 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16610) );
  INV_X1 U13525 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n18127) );
  INV_X1 U13526 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n18156) );
  INV_X1 U13527 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n18237) );
  INV_X1 U13528 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n18308) );
  INV_X1 U13529 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18846) );
  AOI211_X1 U13530 ( .C1(n19020), .C2(n18842), .A(n16151), .B(n18375), .ZN(
        n18998) );
  INV_X1 U13531 ( .A(n18503), .ZN(n18443) );
  INV_X1 U13532 ( .A(n18793), .ZN(n18713) );
  NAND2_X1 U13533 ( .A1(n18414), .A2(n18378), .ZN(n18752) );
  NAND2_X1 U13534 ( .A1(n18414), .A2(n18401), .ZN(n18776) );
  NAND2_X1 U13535 ( .A1(n18870), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n18864) );
  INV_X1 U13536 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n18967) );
  INV_X1 U13537 ( .A(n18964), .ZN(n18879) );
  INV_X1 U13538 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n18903) );
  INV_X1 U13539 ( .A(BUF2_REG_27__SCAN_IN), .ZN(n19389) );
  INV_X1 U13540 ( .A(BUF2_REG_19__SCAN_IN), .ZN(n19392) );
  INV_X1 U13541 ( .A(n16690), .ZN(n16686) );
  INV_X1 U13542 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n19939) );
  OAI21_X1 U13543 ( .B1(n15334), .B2(n20088), .A(n12421), .ZN(P1_U2971) );
  OAI21_X1 U13544 ( .B1(n15814), .B2(n19363), .A(n11521), .ZN(P2_U3025) );
  OR4_X1 U13545 ( .A1(n13311), .A2(n13310), .A3(n13309), .A4(n13308), .ZN(
        P3_U2645) );
  NAND4_X1 U13546 ( .A1(n20303), .A2(P1_M_IO_N_REG_SCAN_IN), .A3(n13275), .A4(
        n13274), .ZN(U214) );
  NAND2_X1 U13547 ( .A1(n10409), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10403) );
  NAND2_X1 U13548 ( .A1(n10411), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n10399) );
  NAND2_X1 U13549 ( .A1(n10398), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n10414) );
  NAND2_X1 U13550 ( .A1(n10397), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n10395) );
  INV_X1 U13551 ( .A(n10395), .ZN(n10383) );
  NAND2_X1 U13552 ( .A1(n10396), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n10394) );
  NOR2_X2 U13553 ( .A1(n10394), .A2(n15788), .ZN(n10393) );
  INV_X1 U13554 ( .A(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n12969) );
  XNOR2_X1 U13555 ( .A(n10386), .B(n12969), .ZN(n12971) );
  NAND2_X1 U13556 ( .A1(n10386), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10384) );
  AND2_X1 U13557 ( .A1(n10387), .A2(n12790), .ZN(n10385) );
  NOR2_X1 U13558 ( .A1(n10386), .A2(n10385), .ZN(n15500) );
  INV_X1 U13559 ( .A(n10387), .ZN(n10388) );
  AOI21_X1 U13560 ( .B1(n15756), .B2(n10390), .A(n10388), .ZN(n15758) );
  NAND2_X1 U13561 ( .A1(n10392), .A2(n15765), .ZN(n10389) );
  AND2_X1 U13562 ( .A1(n10390), .A2(n10389), .ZN(n15767) );
  OR2_X1 U13563 ( .A1(n10393), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n10391) );
  NAND2_X1 U13564 ( .A1(n10392), .A2(n10391), .ZN(n15776) );
  INV_X1 U13565 ( .A(n15776), .ZN(n16446) );
  AOI21_X1 U13566 ( .B1(n15788), .B2(n10394), .A(n10393), .ZN(n15786) );
  OAI21_X1 U13567 ( .B1(n10396), .B2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n10394), .ZN(n15800) );
  INV_X1 U13568 ( .A(n15800), .ZN(n15533) );
  INV_X1 U13569 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n16479) );
  AOI21_X1 U13570 ( .B1(n16479), .B2(n10395), .A(n10396), .ZN(n16472) );
  OAI21_X1 U13571 ( .B1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n10397), .A(
        n10395), .ZN(n16484) );
  AOI21_X1 U13572 ( .B1(n15808), .B2(n10414), .A(n10397), .ZN(n15805) );
  AOI21_X1 U13573 ( .B1(n10413), .B2(n19064), .A(n10398), .ZN(n19063) );
  AOI21_X1 U13574 ( .B1(n15845), .B2(n10412), .A(n9923), .ZN(n19076) );
  AOI21_X1 U13575 ( .B1(n16506), .B2(n10399), .A(n10400), .ZN(n19087) );
  AOI21_X1 U13576 ( .B1(n19111), .B2(n10410), .A(n10411), .ZN(n15854) );
  AOI21_X1 U13577 ( .B1(n15862), .B2(n10401), .A(n10402), .ZN(n19126) );
  AOI21_X1 U13578 ( .B1(n16529), .B2(n10403), .A(n10404), .ZN(n19132) );
  AOI21_X1 U13579 ( .B1(n14424), .B2(n10408), .A(n10409), .ZN(n19143) );
  AOI21_X1 U13580 ( .B1(n16558), .B2(n10406), .A(n9891), .ZN(n19173) );
  AOI21_X1 U13581 ( .B1(n14064), .B2(n10405), .A(n10407), .ZN(n14062) );
  OAI22_X1 U13582 ( .A1(n14298), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(P2_STATE2_REG_0__SCAN_IN), .ZN(
        n19215) );
  INV_X1 U13583 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n19191) );
  OAI22_X1 U13584 ( .A1(n14298), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(
        n19191), .B2(P2_STATE2_REG_0__SCAN_IN), .ZN(n16114) );
  AND2_X1 U13585 ( .A1(n19215), .A2(n16114), .ZN(n14195) );
  OAI21_X1 U13586 ( .B1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n10405), .ZN(n14796) );
  NAND2_X1 U13587 ( .A1(n14195), .A2(n14796), .ZN(n14060) );
  NOR2_X1 U13588 ( .A1(n14062), .A2(n14060), .ZN(n14181) );
  OAI21_X1 U13589 ( .B1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n10407), .A(
        n10406), .ZN(n19324) );
  NAND2_X1 U13590 ( .A1(n14181), .A2(n19324), .ZN(n19171) );
  NOR2_X1 U13591 ( .A1(n19173), .A2(n19171), .ZN(n19158) );
  OAI21_X1 U13592 ( .B1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n9891), .A(
        n10408), .ZN(n19160) );
  NAND2_X1 U13593 ( .A1(n19158), .A2(n19160), .ZN(n19142) );
  NOR2_X1 U13594 ( .A1(n19143), .A2(n19142), .ZN(n14156) );
  OAI21_X1 U13595 ( .B1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n10409), .A(
        n10403), .ZN(n16542) );
  NAND2_X1 U13596 ( .A1(n14156), .A2(n16542), .ZN(n19131) );
  NOR2_X1 U13597 ( .A1(n19132), .A2(n19131), .ZN(n14168) );
  OAI21_X1 U13598 ( .B1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n10404), .A(
        n10401), .ZN(n16523) );
  NAND2_X1 U13599 ( .A1(n14168), .A2(n16523), .ZN(n19124) );
  NOR2_X1 U13600 ( .A1(n19126), .A2(n19124), .ZN(n15611) );
  OAI21_X1 U13601 ( .B1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n10402), .A(
        n10410), .ZN(n16517) );
  NAND2_X1 U13602 ( .A1(n15611), .A2(n16517), .ZN(n19107) );
  NOR2_X1 U13603 ( .A1(n15854), .A2(n19107), .ZN(n19096) );
  OAI21_X1 U13604 ( .B1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n10411), .A(
        n10399), .ZN(n19097) );
  NAND2_X1 U13605 ( .A1(n19096), .A2(n19097), .ZN(n19086) );
  NOR2_X1 U13606 ( .A1(n19087), .A2(n19086), .ZN(n14440) );
  OAI21_X1 U13607 ( .B1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n10400), .A(
        n10412), .ZN(n16499) );
  NAND2_X1 U13608 ( .A1(n14440), .A2(n16499), .ZN(n19074) );
  NOR2_X1 U13609 ( .A1(n19076), .A2(n19074), .ZN(n15599) );
  OAI21_X1 U13610 ( .B1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n9923), .A(
        n10413), .ZN(n16490) );
  NAND2_X1 U13611 ( .A1(n15599), .A2(n16490), .ZN(n19061) );
  NOR2_X1 U13612 ( .A1(n19063), .A2(n19061), .ZN(n15587) );
  OAI21_X1 U13613 ( .B1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n10398), .A(
        n10414), .ZN(n15823) );
  NAND2_X1 U13614 ( .A1(n15587), .A2(n15823), .ZN(n15585) );
  NOR2_X1 U13615 ( .A1(n16472), .A2(n15550), .ZN(n15549) );
  NOR2_X1 U13616 ( .A1(n19159), .A2(n15518), .ZN(n16445) );
  NOR2_X1 U13617 ( .A1(n16446), .A2(n16445), .ZN(n16444) );
  NOR2_X1 U13618 ( .A1(n19159), .A2(n16444), .ZN(n13313) );
  NOR2_X1 U13619 ( .A1(n15767), .A2(n13313), .ZN(n13312) );
  NOR2_X1 U13620 ( .A1(n19159), .A2(n13312), .ZN(n15507) );
  NOR2_X1 U13621 ( .A1(n15758), .A2(n15507), .ZN(n15506) );
  NOR2_X1 U13622 ( .A1(n19159), .A2(n15506), .ZN(n15499) );
  NOR2_X1 U13623 ( .A1(n15500), .A2(n15499), .ZN(n15498) );
  NOR2_X1 U13624 ( .A1(n19159), .A2(n15498), .ZN(n10417) );
  NOR2_X1 U13625 ( .A1(n12971), .A2(n10417), .ZN(n15486) );
  INV_X1 U13626 ( .A(n15486), .ZN(n10419) );
  NOR4_X1 U13627 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(P2_STATEBS16_REG_SCAN_IN), .A4(n13362), .ZN(n10416) );
  NAND2_X1 U13628 ( .A1(n10419), .A2(n10418), .ZN(n11132) );
  MUX2_X1 U13629 ( .A(n20033), .B(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .S(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .Z(n11397) );
  NAND2_X1 U13630 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n20043), .ZN(
        n11260) );
  INV_X1 U13631 ( .A(n11260), .ZN(n10420) );
  NAND2_X1 U13632 ( .A1(n11397), .A2(n10420), .ZN(n10422) );
  NAND2_X1 U13633 ( .A1(n20033), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10421) );
  NAND2_X1 U13634 ( .A1(n10422), .A2(n10421), .ZN(n10515) );
  XNOR2_X1 U13635 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n10514) );
  NAND2_X1 U13636 ( .A1(n10515), .A2(n10514), .ZN(n10513) );
  NAND2_X1 U13637 ( .A1(n20023), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10423) );
  NAND2_X1 U13638 ( .A1(n10513), .A2(n10423), .ZN(n10492) );
  MUX2_X1 U13639 ( .A(n20017), .B(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n10491) );
  NAND3_X1 U13640 ( .A1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n10588), .A3(
        n11383), .ZN(n11363) );
  AND2_X4 U13641 ( .A1(n10425), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10648) );
  NAND2_X2 U13642 ( .A1(n14770), .A2(n10607), .ZN(n14610) );
  AOI22_X1 U13643 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n10663), .B1(
        n10672), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10434) );
  AOI22_X1 U13644 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n10664), .B1(
        n10666), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n10433) );
  NAND2_X1 U13645 ( .A1(n14624), .A2(n10424), .ZN(n10549) );
  NAND2_X1 U13646 ( .A1(n14579), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n10430) );
  NAND2_X1 U13647 ( .A1(n14599), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n10429) );
  NAND2_X1 U13648 ( .A1(n14598), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n10428) );
  NAND2_X1 U13649 ( .A1(n14618), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n10427) );
  AND4_X1 U13650 ( .A1(n10430), .A2(n10429), .A3(n10428), .A4(n10427), .ZN(
        n10432) );
  AND2_X4 U13651 ( .A1(n10436), .A2(n14088), .ZN(n10645) );
  AND2_X2 U13652 ( .A1(n9843), .A2(n10607), .ZN(n14614) );
  AND2_X4 U13653 ( .A1(n10435), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13678) );
  AND2_X2 U13654 ( .A1(n9841), .A2(n10607), .ZN(n14613) );
  AOI22_X1 U13655 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n14614), .B1(
        n14613), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10431) );
  NAND4_X1 U13656 ( .A1(n10434), .A2(n10433), .A3(n10432), .A4(n10431), .ZN(
        n10443) );
  AND2_X2 U13657 ( .A1(n10645), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10674) );
  AOI22_X1 U13658 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n10667), .B1(
        n10674), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10441) );
  AND3_X2 U13659 ( .A1(n10144), .A2(n14088), .A3(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10462) );
  AND2_X2 U13660 ( .A1(n9858), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10665) );
  INV_X1 U13661 ( .A(n10436), .ZN(n13681) );
  AND2_X1 U13662 ( .A1(n10436), .A2(n10437), .ZN(n10673) );
  AOI22_X1 U13663 ( .A1(n10665), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__4__SCAN_IN), .B2(n10673), .ZN(n10440) );
  AND2_X2 U13664 ( .A1(n10647), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10496) );
  AOI22_X1 U13665 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n10485), .B1(
        n10496), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10439) );
  NAND3_X1 U13666 ( .A1(n10441), .A2(n10440), .A3(n10439), .ZN(n10442) );
  AOI22_X1 U13667 ( .A1(n9857), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(n9854), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10447) );
  AOI22_X1 U13668 ( .A1(n10649), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n9847), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10446) );
  AOI22_X1 U13669 ( .A1(n10648), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n10645), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10445) );
  AOI22_X1 U13670 ( .A1(n13678), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n9823), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10444) );
  NAND4_X1 U13671 ( .A1(n10447), .A2(n10446), .A3(n10445), .A4(n10444), .ZN(
        n10448) );
  AOI22_X1 U13672 ( .A1(n9857), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n9854), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10453) );
  AOI22_X1 U13673 ( .A1(n9841), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n10644), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10452) );
  AOI22_X1 U13674 ( .A1(n10649), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n9843), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10451) );
  NAND3_X1 U13675 ( .A1(n10453), .A2(n10452), .A3(n10451), .ZN(n10454) );
  AOI22_X1 U13676 ( .A1(n9858), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n10647), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10460) );
  AOI22_X1 U13677 ( .A1(n10649), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n10646), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10459) );
  AOI22_X1 U13678 ( .A1(n10648), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n9843), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10458) );
  AOI22_X1 U13679 ( .A1(n13678), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n9823), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10457) );
  NAND4_X1 U13680 ( .A1(n10460), .A2(n10459), .A3(n10458), .A4(n10457), .ZN(
        n10461) );
  AOI22_X1 U13681 ( .A1(n9858), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(n9854), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10466) );
  AOI22_X1 U13682 ( .A1(n10649), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n9847), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10465) );
  AOI22_X1 U13683 ( .A1(n10648), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n9843), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10464) );
  AOI22_X1 U13684 ( .A1(n13678), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n10644), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10463) );
  NAND4_X1 U13685 ( .A1(n10466), .A2(n10465), .A3(n10464), .A4(n10463), .ZN(
        n10467) );
  MUX2_X1 U13686 ( .A(n11363), .B(n11439), .S(n10072), .Z(n11366) );
  INV_X1 U13687 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n14188) );
  NAND2_X1 U13688 ( .A1(n10644), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n10469) );
  AOI22_X1 U13689 ( .A1(n9858), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n10647), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10472) );
  AOI22_X1 U13690 ( .A1(n9847), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(n9843), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10476) );
  AOI22_X1 U13691 ( .A1(n9841), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n9823), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10475) );
  AOI22_X1 U13692 ( .A1(n9859), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n9854), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10474) );
  AOI22_X1 U13693 ( .A1(n10649), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10648), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10473) );
  MUX2_X1 U13694 ( .A(n11366), .B(n14188), .S(n10543), .Z(n11272) );
  AOI22_X1 U13695 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n10664), .B1(
        n10666), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10484) );
  AOI22_X1 U13696 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n10663), .B1(
        n10672), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10483) );
  NAND2_X1 U13697 ( .A1(n14579), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n10480) );
  NAND2_X1 U13698 ( .A1(n14599), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n10479) );
  NAND2_X1 U13699 ( .A1(n14598), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(
        n10478) );
  NAND2_X1 U13700 ( .A1(n14618), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(
        n10477) );
  AND4_X1 U13701 ( .A1(n10480), .A2(n10479), .A3(n10478), .A4(n10477), .ZN(
        n10482) );
  AOI22_X1 U13702 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n10667), .B1(
        n10674), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10481) );
  NAND4_X1 U13703 ( .A1(n10484), .A2(n10483), .A3(n10482), .A4(n10481), .ZN(
        n10490) );
  AOI22_X1 U13704 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n14614), .B1(
        n14613), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10488) );
  AOI22_X1 U13705 ( .A1(n10496), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__3__SCAN_IN), .B2(n10673), .ZN(n10487) );
  AOI22_X1 U13706 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n10665), .B1(
        n10485), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10486) );
  NAND3_X1 U13707 ( .A1(n10488), .A2(n10487), .A3(n10486), .ZN(n10489) );
  NOR2_X1 U13708 ( .A1(n10492), .A2(n10491), .ZN(n10493) );
  INV_X1 U13709 ( .A(n11375), .ZN(n10495) );
  MUX2_X1 U13710 ( .A(n10707), .B(n10495), .S(n11379), .Z(n11365) );
  INV_X1 U13711 ( .A(P2_EBX_REG_3__SCAN_IN), .ZN(n13628) );
  MUX2_X1 U13712 ( .A(n11365), .B(n13628), .S(n10543), .Z(n11258) );
  AOI22_X1 U13713 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n10667), .B1(
        n10674), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10499) );
  AOI22_X1 U13714 ( .A1(n10485), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__2__SCAN_IN), .B2(n10673), .ZN(n10498) );
  AOI22_X1 U13715 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n10665), .B1(
        n10496), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10497) );
  INV_X1 U13716 ( .A(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10500) );
  OR2_X1 U13717 ( .A1(n14603), .A2(n10500), .ZN(n10504) );
  INV_X1 U13718 ( .A(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n10769) );
  OR2_X1 U13719 ( .A1(n14609), .A2(n10769), .ZN(n10503) );
  NAND2_X1 U13720 ( .A1(n14613), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n10502) );
  NAND2_X1 U13721 ( .A1(n14614), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n10501) );
  NAND4_X1 U13722 ( .A1(n10504), .A2(n10503), .A3(n10502), .A4(n10501), .ZN(
        n10512) );
  AOI22_X1 U13723 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n14598), .B1(
        n14618), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10510) );
  AOI22_X1 U13724 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n14599), .B1(
        n14579), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10509) );
  INV_X1 U13725 ( .A(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10505) );
  INV_X1 U13726 ( .A(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10506) );
  OR2_X1 U13727 ( .A1(n14610), .A2(n10506), .ZN(n10507) );
  NAND4_X1 U13728 ( .A1(n10510), .A2(n10509), .A3(n10508), .A4(n10507), .ZN(
        n10511) );
  OAI21_X1 U13729 ( .B1(n10515), .B2(n10514), .A(n10513), .ZN(n11373) );
  AOI22_X1 U13730 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n10496), .B1(
        n10485), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10521) );
  AOI22_X1 U13731 ( .A1(n10672), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_11__1__SCAN_IN), .B2(n10665), .ZN(n10520) );
  AOI22_X1 U13732 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n10663), .B1(
        n10666), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10519) );
  AOI22_X1 U13733 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n10667), .B1(
        n10674), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10518) );
  NAND4_X1 U13734 ( .A1(n10521), .A2(n10520), .A3(n10519), .A4(n10518), .ZN(
        n10527) );
  AOI22_X1 U13735 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n14598), .B1(
        n14579), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10525) );
  AOI22_X1 U13736 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n14599), .B1(
        n14618), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10524) );
  AOI22_X1 U13737 ( .A1(n10664), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__1__SCAN_IN), .B2(n10673), .ZN(n10523) );
  AOI22_X1 U13738 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n14614), .B1(
        n14613), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10522) );
  NAND4_X1 U13739 ( .A1(n10525), .A2(n10524), .A3(n10523), .A4(n10522), .ZN(
        n10526) );
  NOR2_X1 U13740 ( .A1(n10527), .A2(n10526), .ZN(n11428) );
  OR2_X1 U13741 ( .A1(P2_EBX_REG_0__SCAN_IN), .A2(P2_EBX_REG_1__SCAN_IN), .ZN(
        n10528) );
  MUX2_X1 U13742 ( .A(n11428), .B(n10528), .S(n10543), .Z(n11265) );
  NAND2_X1 U13743 ( .A1(n11272), .A2(n11271), .ZN(n11277) );
  AOI22_X1 U13744 ( .A1(n10664), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10663), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10537) );
  AOI22_X1 U13745 ( .A1(n10672), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n10666), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10536) );
  INV_X1 U13746 ( .A(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10529) );
  INV_X1 U13747 ( .A(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11215) );
  OAI22_X1 U13748 ( .A1(n10351), .A2(n10529), .B1(n10549), .B2(n11215), .ZN(
        n10533) );
  INV_X1 U13749 ( .A(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10531) );
  INV_X1 U13750 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13669) );
  OAI22_X1 U13751 ( .A1(n10352), .A2(n10531), .B1(n10530), .B2(n13669), .ZN(
        n10532) );
  NOR2_X1 U13752 ( .A1(n10533), .A2(n10532), .ZN(n10535) );
  AOI22_X1 U13753 ( .A1(n10667), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n14613), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10534) );
  NAND4_X1 U13754 ( .A1(n10537), .A2(n10536), .A3(n10535), .A4(n10534), .ZN(
        n10542) );
  AOI22_X1 U13755 ( .A1(n10674), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n14614), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10540) );
  AOI22_X1 U13756 ( .A1(n10665), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n14598), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10539) );
  AOI22_X1 U13757 ( .A1(n10485), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10496), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10538) );
  NAND3_X1 U13758 ( .A1(n10540), .A2(n10539), .A3(n10538), .ZN(n10541) );
  NAND2_X1 U13759 ( .A1(n10960), .A2(n11230), .ZN(n10714) );
  INV_X1 U13760 ( .A(P2_EBX_REG_5__SCAN_IN), .ZN(n10544) );
  NAND2_X1 U13761 ( .A1(n10543), .A2(n10544), .ZN(n10545) );
  AOI22_X1 U13762 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n10667), .B1(
        n10674), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10548) );
  AOI22_X1 U13763 ( .A1(n10665), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n14618), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10547) );
  AOI22_X1 U13764 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n10485), .B1(
        n10496), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10546) );
  AOI22_X1 U13765 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n14598), .B1(
        n14599), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10555) );
  AOI22_X1 U13766 ( .A1(n14579), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n10673), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10554) );
  INV_X1 U13767 ( .A(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10550) );
  OR2_X1 U13768 ( .A1(n14601), .A2(n10550), .ZN(n10553) );
  INV_X1 U13769 ( .A(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10551) );
  OR2_X1 U13770 ( .A1(n14603), .A2(n10551), .ZN(n10552) );
  NAND4_X1 U13771 ( .A1(n10555), .A2(n10554), .A3(n10553), .A4(n10552), .ZN(
        n10562) );
  INV_X1 U13772 ( .A(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10556) );
  OR2_X1 U13773 ( .A1(n14610), .A2(n10556), .ZN(n10560) );
  INV_X1 U13774 ( .A(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11242) );
  OR2_X1 U13775 ( .A1(n14609), .A2(n11242), .ZN(n10559) );
  NAND2_X1 U13776 ( .A1(n14614), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n10558) );
  NAND2_X1 U13777 ( .A1(n14613), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n10557) );
  NAND4_X1 U13778 ( .A1(n10560), .A2(n10559), .A3(n10558), .A4(n10557), .ZN(
        n10561) );
  NOR2_X1 U13779 ( .A1(n10562), .A2(n10561), .ZN(n10563) );
  MUX2_X1 U13780 ( .A(n11250), .B(P2_EBX_REG_6__SCAN_IN), .S(n10543), .Z(
        n11255) );
  AOI22_X1 U13781 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n10667), .B1(
        n10674), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10566) );
  AOI22_X1 U13782 ( .A1(n10665), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n14618), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10565) );
  AOI22_X1 U13783 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n10485), .B1(
        n10496), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10564) );
  AND3_X1 U13784 ( .A1(n10566), .A2(n10565), .A3(n10564), .ZN(n10581) );
  AOI22_X1 U13785 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n14598), .B1(
        n14599), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10572) );
  AOI22_X1 U13786 ( .A1(n14579), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n10673), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10571) );
  INV_X1 U13787 ( .A(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n10567) );
  OR2_X1 U13788 ( .A1(n14601), .A2(n10567), .ZN(n10570) );
  INV_X1 U13789 ( .A(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10568) );
  OR2_X1 U13790 ( .A1(n14603), .A2(n10568), .ZN(n10569) );
  NAND4_X1 U13791 ( .A1(n10572), .A2(n10571), .A3(n10570), .A4(n10569), .ZN(
        n10579) );
  INV_X1 U13792 ( .A(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n10573) );
  OR2_X1 U13793 ( .A1(n14610), .A2(n10573), .ZN(n10577) );
  OR2_X1 U13794 ( .A1(n14609), .A2(n19713), .ZN(n10576) );
  NAND2_X1 U13795 ( .A1(n14614), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n10575) );
  NAND2_X1 U13796 ( .A1(n14613), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n10574) );
  NAND4_X1 U13797 ( .A1(n10577), .A2(n10576), .A3(n10575), .A4(n10574), .ZN(
        n10578) );
  NOR2_X1 U13798 ( .A1(n10579), .A2(n10578), .ZN(n10580) );
  AND2_X2 U13799 ( .A1(n10581), .A2(n10580), .ZN(n11254) );
  MUX2_X1 U13800 ( .A(n11254), .B(P2_EBX_REG_7__SCAN_IN), .S(n10543), .Z(
        n11302) );
  NOR2_X1 U13801 ( .A1(n11255), .A2(n11302), .ZN(n10582) );
  AND2_X2 U13802 ( .A1(n11301), .A2(n10582), .ZN(n11299) );
  INV_X1 U13803 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n19122) );
  NAND2_X1 U13804 ( .A1(n10543), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n11298) );
  INV_X1 U13805 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n10583) );
  NAND2_X1 U13806 ( .A1(n12460), .A2(n11320), .ZN(n11318) );
  NAND2_X1 U13807 ( .A1(n10543), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n11319) );
  NAND2_X1 U13808 ( .A1(n10543), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n11336) );
  NAND2_X1 U13809 ( .A1(n11338), .A2(n11336), .ZN(n11341) );
  NOR2_X2 U13810 ( .A1(n9888), .A2(n11343), .ZN(n11349) );
  NAND2_X1 U13811 ( .A1(n10543), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n11348) );
  NAND2_X1 U13812 ( .A1(n10543), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n11353) );
  INV_X1 U13813 ( .A(P2_EBX_REG_20__SCAN_IN), .ZN(n10585) );
  NAND2_X1 U13814 ( .A1(n12444), .A2(n12460), .ZN(n11135) );
  NAND2_X1 U13815 ( .A1(n10543), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n12443) );
  AND2_X1 U13816 ( .A1(n10543), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n12448) );
  INV_X1 U13817 ( .A(P2_EBX_REG_25__SCAN_IN), .ZN(n15653) );
  NAND2_X1 U13818 ( .A1(n10543), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n12466) );
  NAND2_X1 U13819 ( .A1(n10543), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n12424) );
  NAND2_X1 U13820 ( .A1(n12469), .A2(n12424), .ZN(n12805) );
  NAND2_X1 U13821 ( .A1(n10543), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n10586) );
  XNOR2_X1 U13822 ( .A(n12805), .B(n10586), .ZN(n12803) );
  XNOR2_X1 U13823 ( .A(n11397), .B(n11260), .ZN(n11368) );
  INV_X1 U13824 ( .A(n11363), .ZN(n10589) );
  NOR3_X1 U13825 ( .A1(n11375), .A2(n11373), .A3(n10589), .ZN(n11389) );
  AND2_X1 U13826 ( .A1(n11368), .A2(n11389), .ZN(n10590) );
  AOI22_X1 U13827 ( .A1(n9857), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(n9854), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10592) );
  AOI22_X1 U13828 ( .A1(n9843), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(n9823), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10591) );
  AND2_X1 U13829 ( .A1(n10592), .A2(n10591), .ZN(n10596) );
  AOI22_X1 U13830 ( .A1(n10649), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n13678), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10595) );
  AOI22_X1 U13831 ( .A1(n10646), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n10648), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10593) );
  AOI22_X1 U13832 ( .A1(n10649), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n10648), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10602) );
  AOI22_X1 U13833 ( .A1(n10646), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n10644), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10601) );
  AOI22_X1 U13834 ( .A1(n9857), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n10647), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10600) );
  AOI22_X1 U13835 ( .A1(n10649), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n10648), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10606) );
  AOI22_X1 U13836 ( .A1(n9858), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n10647), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10605) );
  AOI22_X1 U13837 ( .A1(n10646), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n9843), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10604) );
  AOI22_X1 U13838 ( .A1(n9841), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(n9822), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10603) );
  AOI22_X1 U13839 ( .A1(n10649), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n10648), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10613) );
  AOI22_X1 U13840 ( .A1(n9857), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n9854), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10612) );
  AOI22_X1 U13841 ( .A1(n9841), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n9823), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10610) );
  AOI22_X1 U13842 ( .A1(n10646), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n9843), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10609) );
  AND3_X1 U13843 ( .A1(n10610), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(
        n10609), .ZN(n10611) );
  NAND3_X1 U13844 ( .A1(n10613), .A2(n10612), .A3(n10611), .ZN(n10614) );
  AOI22_X1 U13845 ( .A1(n10649), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n10648), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10619) );
  AOI22_X1 U13846 ( .A1(n9859), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n10647), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10618) );
  AOI22_X1 U13847 ( .A1(n10646), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n10645), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10617) );
  AOI22_X1 U13848 ( .A1(n13678), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n10644), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10616) );
  NAND4_X1 U13849 ( .A1(n10619), .A2(n10618), .A3(n10617), .A4(n10616), .ZN(
        n10625) );
  AOI22_X1 U13850 ( .A1(n10646), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n10645), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10623) );
  AOI22_X1 U13851 ( .A1(n13678), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n10644), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10622) );
  AOI22_X1 U13852 ( .A1(n9858), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n10647), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10621) );
  AOI22_X1 U13853 ( .A1(n10649), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n10648), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10620) );
  NAND4_X1 U13854 ( .A1(n10623), .A2(n10622), .A3(n10621), .A4(n10620), .ZN(
        n10624) );
  AOI22_X1 U13855 ( .A1(n9859), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(n9854), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10627) );
  AOI22_X1 U13856 ( .A1(n9847), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n10645), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10626) );
  AOI22_X1 U13857 ( .A1(n10649), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n10648), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10630) );
  NAND2_X1 U13858 ( .A1(n10644), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n10629) );
  NAND3_X1 U13859 ( .A1(n10372), .A2(n10607), .A3(n10631), .ZN(n10639) );
  AOI22_X1 U13860 ( .A1(n13678), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n9823), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n10636) );
  AOI22_X1 U13861 ( .A1(n9857), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n9854), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10635) );
  AOI22_X1 U13862 ( .A1(n10649), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n10648), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10633) );
  NAND4_X1 U13863 ( .A1(n10637), .A2(n10636), .A3(n10635), .A4(n10634), .ZN(
        n10638) );
  AOI22_X1 U13864 ( .A1(n10646), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n10645), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n10641) );
  AOI22_X1 U13865 ( .A1(n10649), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n10648), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10640) );
  AOI22_X1 U13866 ( .A1(n13678), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n9822), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n10653) );
  AOI22_X1 U13867 ( .A1(n10646), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n10645), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10652) );
  AOI22_X1 U13868 ( .A1(n9859), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n10647), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10651) );
  AOI22_X1 U13869 ( .A1(n10649), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n10648), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n10650) );
  AND3_X2 U13870 ( .A1(n10966), .A2(n10955), .A3(n10654), .ZN(n11408) );
  NAND2_X1 U13871 ( .A1(n13362), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10928) );
  NAND2_X1 U13872 ( .A1(n10976), .A2(n13386), .ZN(n10655) );
  AND2_X1 U13873 ( .A1(n10951), .A2(n11487), .ZN(n10656) );
  AND3_X2 U13874 ( .A1(n10656), .A2(n10954), .A3(n13389), .ZN(n16157) );
  NAND2_X1 U13875 ( .A1(n13686), .A2(n13386), .ZN(n13359) );
  AND2_X1 U13876 ( .A1(n20056), .A2(n10072), .ZN(n11126) );
  NAND2_X1 U13877 ( .A1(n20061), .A2(n20069), .ZN(n11127) );
  AND2_X1 U13878 ( .A1(P2_EBX_REG_31__SCAN_IN), .A2(n11127), .ZN(n10658) );
  AND2_X1 U13879 ( .A1(n10935), .A2(n19420), .ZN(n13388) );
  NAND2_X1 U13880 ( .A1(n13388), .A2(n10712), .ZN(n10908) );
  NAND2_X1 U13881 ( .A1(n12818), .A2(P2_REIP_REG_4__SCAN_IN), .ZN(n10662) );
  NOR2_X1 U13882 ( .A1(n19420), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n10689) );
  AOI22_X1 U13883 ( .A1(n12819), .A2(P2_EAX_REG_4__SCAN_IN), .B1(n10690), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n10661) );
  INV_X1 U13884 ( .A(n11439), .ZN(n10659) );
  OR2_X1 U13885 ( .A1(n10890), .A2(n10659), .ZN(n10660) );
  AOI22_X1 U13886 ( .A1(n14614), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n10496), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10671) );
  AOI22_X1 U13887 ( .A1(n10664), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10663), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10670) );
  AOI22_X1 U13888 ( .A1(n10666), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n10665), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10669) );
  AOI22_X1 U13889 ( .A1(n10667), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n14613), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10668) );
  AOI22_X1 U13890 ( .A1(n14579), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n14599), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10678) );
  AOI22_X1 U13891 ( .A1(n14618), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n14598), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10677) );
  AOI22_X1 U13892 ( .A1(n10672), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10485), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10676) );
  AOI22_X1 U13893 ( .A1(n10674), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n10673), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10675) );
  INV_X1 U13894 ( .A(n10968), .ZN(n13391) );
  NAND2_X1 U13895 ( .A1(n13391), .A2(n10690), .ZN(n10699) );
  OAI22_X1 U13896 ( .A1(n19420), .A2(P2_STATE2_REG_3__SCAN_IN), .B1(n20043), 
        .B2(n20013), .ZN(n10681) );
  INV_X1 U13897 ( .A(n10681), .ZN(n10682) );
  AND2_X1 U13898 ( .A1(n10699), .A2(n10682), .ZN(n10683) );
  INV_X1 U13899 ( .A(n10908), .ZN(n10684) );
  NAND2_X1 U13900 ( .A1(n10684), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n10688) );
  INV_X1 U13901 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n13658) );
  NAND2_X1 U13902 ( .A1(n20062), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n10685) );
  OAI211_X1 U13903 ( .C1(n19420), .C2(n13658), .A(n10685), .B(n20013), .ZN(
        n10686) );
  INV_X1 U13904 ( .A(n10686), .ZN(n10687) );
  NAND2_X1 U13905 ( .A1(n10688), .A2(n10687), .ZN(n13368) );
  INV_X1 U13906 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n19934) );
  AOI22_X1 U13907 ( .A1(n10689), .A2(P2_EAX_REG_1__SCAN_IN), .B1(n10690), .B2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n10691) );
  NAND2_X1 U13908 ( .A1(n10692), .A2(n10691), .ZN(n10698) );
  INV_X1 U13909 ( .A(n10698), .ZN(n10693) );
  OR2_X1 U13910 ( .A1(n11428), .A2(n10890), .ZN(n10697) );
  AND2_X1 U13911 ( .A1(n19420), .A2(n20036), .ZN(n10695) );
  NOR2_X1 U13912 ( .A1(n20036), .A2(n20033), .ZN(n10694) );
  AOI21_X1 U13913 ( .B1(n10968), .B2(n10695), .A(n10694), .ZN(n10696) );
  AND2_X1 U13914 ( .A1(n10697), .A2(n10696), .ZN(n13452) );
  NAND2_X1 U13915 ( .A1(n13453), .A2(n13452), .ZN(n13451) );
  OR2_X1 U13916 ( .A1(n13366), .A2(n10698), .ZN(n10702) );
  OR2_X1 U13917 ( .A1(n10890), .A2(n11433), .ZN(n10700) );
  OAI211_X1 U13918 ( .C1(n20013), .C2(n20023), .A(n10700), .B(n10699), .ZN(
        n10701) );
  AND3_X1 U13919 ( .A1(n13451), .A2(n10702), .A3(n10701), .ZN(n10703) );
  NAND2_X1 U13920 ( .A1(n12818), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n10705) );
  AOI22_X1 U13921 ( .A1(n12819), .A2(P2_EAX_REG_2__SCAN_IN), .B1(n10690), .B2(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n10704) );
  NAND2_X1 U13922 ( .A1(n10705), .A2(n10704), .ZN(n13913) );
  INV_X1 U13923 ( .A(n10707), .ZN(n11183) );
  NAND2_X1 U13924 ( .A1(n12818), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n10711) );
  AOI22_X1 U13925 ( .A1(n10690), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B1(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n10709) );
  NAND2_X1 U13926 ( .A1(n12819), .A2(P2_EAX_REG_3__SCAN_IN), .ZN(n10708) );
  AND2_X1 U13927 ( .A1(n10709), .A2(n10708), .ZN(n10710) );
  OAI211_X1 U13928 ( .C1(n10890), .C2(n11183), .A(n10711), .B(n10710), .ZN(
        n13874) );
  NAND2_X1 U13929 ( .A1(n12818), .A2(P2_REIP_REG_5__SCAN_IN), .ZN(n10718) );
  INV_X1 U13930 ( .A(n10712), .ZN(n10713) );
  OR2_X1 U13931 ( .A1(n10714), .A2(n10713), .ZN(n10717) );
  NAND2_X1 U13932 ( .A1(n12819), .A2(P2_EAX_REG_5__SCAN_IN), .ZN(n10716) );
  NAND2_X1 U13933 ( .A1(n10690), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10715) );
  NAND4_X1 U13934 ( .A1(n10718), .A2(n10717), .A3(n10716), .A4(n10715), .ZN(
        n14273) );
  AOI21_X1 U13935 ( .B1(n14272), .B2(n14273), .A(n9939), .ZN(n10719) );
  NAND2_X1 U13936 ( .A1(n12818), .A2(P2_REIP_REG_6__SCAN_IN), .ZN(n10721) );
  AOI22_X1 U13937 ( .A1(n12819), .A2(P2_EAX_REG_6__SCAN_IN), .B1(n10690), .B2(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n10720) );
  NAND2_X1 U13938 ( .A1(n10721), .A2(n10720), .ZN(n14480) );
  AOI21_X1 U13939 ( .B1(n14481), .B2(n14480), .A(n9930), .ZN(n10722) );
  NAND2_X1 U13940 ( .A1(n12818), .A2(P2_REIP_REG_7__SCAN_IN), .ZN(n10724) );
  AOI22_X1 U13941 ( .A1(n12819), .A2(P2_EAX_REG_7__SCAN_IN), .B1(n10690), .B2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n10723) );
  NAND2_X1 U13942 ( .A1(n10724), .A2(n10723), .ZN(n14413) );
  NAND2_X1 U13943 ( .A1(n12818), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n10744) );
  AOI22_X1 U13944 ( .A1(n12819), .A2(P2_EAX_REG_8__SCAN_IN), .B1(n10690), .B2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n10743) );
  AOI22_X1 U13945 ( .A1(n14579), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n14598), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10728) );
  AOI22_X1 U13946 ( .A1(n14618), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n14599), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10727) );
  INV_X1 U13947 ( .A(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n14312) );
  OR2_X1 U13948 ( .A1(n14601), .A2(n14312), .ZN(n10726) );
  INV_X1 U13949 ( .A(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n19582) );
  OR2_X1 U13950 ( .A1(n14610), .A2(n19582), .ZN(n10725) );
  AND4_X1 U13951 ( .A1(n10728), .A2(n10727), .A3(n10726), .A4(n10725), .ZN(
        n10741) );
  AOI22_X1 U13952 ( .A1(n10667), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n14614), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10740) );
  NAND2_X1 U13953 ( .A1(n10665), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n10732) );
  NAND2_X1 U13954 ( .A1(n10485), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n10731) );
  NAND2_X1 U13955 ( .A1(n10496), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n10730) );
  NAND2_X1 U13956 ( .A1(n10673), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n10729) );
  AND4_X1 U13957 ( .A1(n10732), .A2(n10731), .A3(n10730), .A4(n10729), .ZN(
        n10739) );
  INV_X1 U13958 ( .A(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10733) );
  OR2_X1 U13959 ( .A1(n14603), .A2(n10733), .ZN(n10737) );
  INV_X1 U13960 ( .A(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n14207) );
  OR2_X1 U13961 ( .A1(n14609), .A2(n14207), .ZN(n10736) );
  NAND2_X1 U13962 ( .A1(n14613), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n10735) );
  NAND2_X1 U13963 ( .A1(n10674), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n10734) );
  AND4_X1 U13964 ( .A1(n10737), .A2(n10736), .A3(n10735), .A4(n10734), .ZN(
        n10738) );
  NAND4_X1 U13965 ( .A1(n10741), .A2(n10740), .A3(n10739), .A4(n10738), .ZN(
        n13699) );
  INV_X1 U13966 ( .A(n13699), .ZN(n13822) );
  OR2_X1 U13967 ( .A1(n10890), .A2(n13822), .ZN(n10742) );
  AOI22_X1 U13968 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n14598), .B1(
        n14599), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10749) );
  AOI22_X1 U13969 ( .A1(n14579), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n10673), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10748) );
  INV_X1 U13970 ( .A(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n14309) );
  OR2_X1 U13971 ( .A1(n14601), .A2(n14309), .ZN(n10747) );
  INV_X1 U13972 ( .A(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10745) );
  OR2_X1 U13973 ( .A1(n14603), .A2(n10745), .ZN(n10746) );
  AND4_X1 U13974 ( .A1(n10749), .A2(n10748), .A3(n10747), .A4(n10746), .ZN(
        n10761) );
  AOI22_X1 U13975 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n10674), .B1(
        n10667), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10760) );
  OR2_X1 U13976 ( .A1(n14610), .A2(n19586), .ZN(n10753) );
  INV_X1 U13977 ( .A(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n14223) );
  OR2_X1 U13978 ( .A1(n14609), .A2(n14223), .ZN(n10752) );
  NAND2_X1 U13979 ( .A1(n14614), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n10751) );
  NAND2_X1 U13980 ( .A1(n14613), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n10750) );
  AND4_X1 U13981 ( .A1(n10753), .A2(n10752), .A3(n10751), .A4(n10750), .ZN(
        n10759) );
  NAND2_X1 U13982 ( .A1(n10665), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n10757) );
  NAND2_X1 U13983 ( .A1(n10485), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n10756) );
  NAND2_X1 U13984 ( .A1(n10496), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n10755) );
  NAND2_X1 U13985 ( .A1(n14618), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n10754) );
  AND4_X1 U13986 ( .A1(n10757), .A2(n10756), .A3(n10755), .A4(n10754), .ZN(
        n10758) );
  NAND4_X1 U13987 ( .A1(n10761), .A2(n10760), .A3(n10759), .A4(n10758), .ZN(
        n13722) );
  INV_X1 U13988 ( .A(n13722), .ZN(n10764) );
  NAND2_X1 U13989 ( .A1(n12818), .A2(P2_REIP_REG_9__SCAN_IN), .ZN(n10763) );
  AOI22_X1 U13990 ( .A1(n12819), .A2(P2_EAX_REG_9__SCAN_IN), .B1(n10690), .B2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n10762) );
  OAI211_X1 U13991 ( .C1(n10890), .C2(n10764), .A(n10763), .B(n10762), .ZN(
        n14532) );
  NAND2_X1 U13992 ( .A1(n12818), .A2(P2_REIP_REG_10__SCAN_IN), .ZN(n10785) );
  AOI22_X1 U13993 ( .A1(n12819), .A2(P2_EAX_REG_10__SCAN_IN), .B1(n10690), 
        .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n10784) );
  AOI22_X1 U13994 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n10674), .B1(
        n10667), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10767) );
  AOI22_X1 U13995 ( .A1(n10485), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__2__SCAN_IN), .B2(n10673), .ZN(n10766) );
  AOI22_X1 U13996 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n10665), .B1(
        n10496), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10765) );
  AND3_X1 U13997 ( .A1(n10767), .A2(n10766), .A3(n10765), .ZN(n10782) );
  AOI22_X1 U13998 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n14598), .B1(
        n14579), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10773) );
  AOI22_X1 U13999 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n14618), .B1(
        n14599), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10772) );
  INV_X1 U14000 ( .A(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10768) );
  OR2_X1 U14001 ( .A1(n14603), .A2(n10768), .ZN(n10771) );
  OR2_X1 U14002 ( .A1(n14601), .A2(n10769), .ZN(n10770) );
  NAND4_X1 U14003 ( .A1(n10773), .A2(n10772), .A3(n10771), .A4(n10770), .ZN(
        n10780) );
  INV_X1 U14004 ( .A(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10774) );
  OR2_X1 U14005 ( .A1(n14610), .A2(n10774), .ZN(n10778) );
  INV_X1 U14006 ( .A(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n14345) );
  OR2_X1 U14007 ( .A1(n14609), .A2(n14345), .ZN(n10777) );
  NAND2_X1 U14008 ( .A1(n14613), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n10776) );
  NAND2_X1 U14009 ( .A1(n14614), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n10775) );
  NAND4_X1 U14010 ( .A1(n10778), .A2(n10777), .A3(n10776), .A4(n10775), .ZN(
        n10779) );
  NOR2_X1 U14011 ( .A1(n10780), .A2(n10779), .ZN(n10781) );
  OR2_X1 U14012 ( .A1(n10890), .A2(n13704), .ZN(n10783) );
  AOI22_X1 U14013 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n10674), .B1(
        n10667), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10788) );
  AOI22_X1 U14014 ( .A1(n10665), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n14618), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10787) );
  AOI22_X1 U14015 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n10485), .B1(
        n10496), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10786) );
  AND3_X1 U14016 ( .A1(n10788), .A2(n10787), .A3(n10786), .ZN(n10802) );
  AOI22_X1 U14017 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n14598), .B1(
        n14599), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10793) );
  AOI22_X1 U14018 ( .A1(n14579), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n10673), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10792) );
  INV_X1 U14019 ( .A(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n21213) );
  OR2_X1 U14020 ( .A1(n14601), .A2(n21213), .ZN(n10791) );
  INV_X1 U14021 ( .A(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10789) );
  OR2_X1 U14022 ( .A1(n14603), .A2(n10789), .ZN(n10790) );
  NAND4_X1 U14023 ( .A1(n10793), .A2(n10792), .A3(n10791), .A4(n10790), .ZN(
        n10800) );
  INV_X1 U14024 ( .A(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10794) );
  OR2_X1 U14025 ( .A1(n14610), .A2(n10794), .ZN(n10798) );
  INV_X1 U14026 ( .A(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n14364) );
  OR2_X1 U14027 ( .A1(n14609), .A2(n14364), .ZN(n10797) );
  NAND2_X1 U14028 ( .A1(n14614), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(
        n10796) );
  NAND2_X1 U14029 ( .A1(n14613), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n10795) );
  NAND4_X1 U14030 ( .A1(n10798), .A2(n10797), .A3(n10796), .A4(n10795), .ZN(
        n10799) );
  NOR2_X1 U14031 ( .A1(n10800), .A2(n10799), .ZN(n10801) );
  NAND2_X1 U14032 ( .A1(n12818), .A2(P2_REIP_REG_11__SCAN_IN), .ZN(n10804) );
  AOI22_X1 U14033 ( .A1(n12819), .A2(P2_EAX_REG_11__SCAN_IN), .B1(n10690), 
        .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n10803) );
  OAI211_X1 U14034 ( .C1(n13814), .C2(n10890), .A(n10804), .B(n10803), .ZN(
        n16076) );
  NAND2_X1 U14035 ( .A1(n12818), .A2(P2_REIP_REG_12__SCAN_IN), .ZN(n10827) );
  AOI22_X1 U14036 ( .A1(n12819), .A2(P2_EAX_REG_12__SCAN_IN), .B1(n10690), 
        .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n10826) );
  AOI22_X1 U14037 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n14618), .B1(
        n14579), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10809) );
  AOI22_X1 U14038 ( .A1(n14599), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n10673), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10808) );
  INV_X1 U14039 ( .A(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n14544) );
  OR2_X1 U14040 ( .A1(n14609), .A2(n14544), .ZN(n10807) );
  INV_X1 U14041 ( .A(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n10805) );
  OR2_X1 U14042 ( .A1(n14601), .A2(n10805), .ZN(n10806) );
  AND4_X1 U14043 ( .A1(n10809), .A2(n10808), .A3(n10807), .A4(n10806), .ZN(
        n10823) );
  AOI22_X1 U14044 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n10674), .B1(
        n10667), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10822) );
  INV_X1 U14045 ( .A(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10810) );
  OR2_X1 U14046 ( .A1(n14610), .A2(n10810), .ZN(n10815) );
  INV_X1 U14047 ( .A(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10811) );
  OR2_X1 U14048 ( .A1(n14603), .A2(n10811), .ZN(n10814) );
  NAND2_X1 U14049 ( .A1(n14614), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n10813) );
  NAND2_X1 U14050 ( .A1(n14613), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n10812) );
  AND4_X1 U14051 ( .A1(n10815), .A2(n10814), .A3(n10813), .A4(n10812), .ZN(
        n10821) );
  NAND2_X1 U14052 ( .A1(n10485), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n10819) );
  NAND2_X1 U14053 ( .A1(n10665), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n10818) );
  NAND2_X1 U14054 ( .A1(n10496), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n10817) );
  NAND2_X1 U14055 ( .A1(n14598), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n10816) );
  AND4_X1 U14056 ( .A1(n10819), .A2(n10818), .A3(n10817), .A4(n10816), .ZN(
        n10820) );
  NAND4_X1 U14057 ( .A1(n10823), .A2(n10822), .A3(n10821), .A4(n10820), .ZN(
        n13831) );
  INV_X1 U14058 ( .A(n13831), .ZN(n10824) );
  OR2_X1 U14059 ( .A1(n10890), .A2(n10824), .ZN(n10825) );
  INV_X1 U14060 ( .A(n10890), .ZN(n10870) );
  AOI22_X1 U14061 ( .A1(n14599), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n14598), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10833) );
  AOI22_X1 U14062 ( .A1(n14579), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n10673), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10832) );
  INV_X1 U14063 ( .A(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10828) );
  OR2_X1 U14064 ( .A1(n14601), .A2(n10828), .ZN(n10831) );
  INV_X1 U14065 ( .A(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10829) );
  OR2_X1 U14066 ( .A1(n14603), .A2(n10829), .ZN(n10830) );
  AND4_X1 U14067 ( .A1(n10833), .A2(n10832), .A3(n10831), .A4(n10830), .ZN(
        n10846) );
  AOI22_X1 U14068 ( .A1(n10674), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n10667), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10845) );
  INV_X1 U14069 ( .A(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10834) );
  OR2_X1 U14070 ( .A1(n14610), .A2(n10834), .ZN(n10838) );
  INV_X1 U14071 ( .A(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n14562) );
  OR2_X1 U14072 ( .A1(n14609), .A2(n14562), .ZN(n10837) );
  NAND2_X1 U14073 ( .A1(n14614), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n10836) );
  NAND2_X1 U14074 ( .A1(n14613), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n10835) );
  AND4_X1 U14075 ( .A1(n10838), .A2(n10837), .A3(n10836), .A4(n10835), .ZN(
        n10844) );
  NAND2_X1 U14076 ( .A1(n10665), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n10842) );
  NAND2_X1 U14077 ( .A1(n10485), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n10841) );
  NAND2_X1 U14078 ( .A1(n10496), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n10840) );
  NAND2_X1 U14079 ( .A1(n14618), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n10839) );
  AND4_X1 U14080 ( .A1(n10842), .A2(n10841), .A3(n10840), .A4(n10839), .ZN(
        n10843) );
  NAND4_X1 U14081 ( .A1(n10846), .A2(n10845), .A3(n10844), .A4(n10843), .ZN(
        n14032) );
  AOI22_X1 U14082 ( .A1(n10870), .A2(n14032), .B1(n12818), .B2(
        P2_REIP_REG_13__SCAN_IN), .ZN(n10848) );
  AOI22_X1 U14083 ( .A1(n12819), .A2(P2_EAX_REG_13__SCAN_IN), .B1(n10690), 
        .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n10847) );
  NAND2_X1 U14084 ( .A1(n10848), .A2(n10847), .ZN(n16060) );
  AOI22_X1 U14085 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n14618), .B1(
        n14598), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10853) );
  AOI22_X1 U14086 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n14599), .B1(
        n14579), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10852) );
  OR2_X1 U14087 ( .A1(n14601), .A2(n11242), .ZN(n10851) );
  INV_X1 U14088 ( .A(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10849) );
  OR2_X1 U14089 ( .A1(n14603), .A2(n10849), .ZN(n10850) );
  AND4_X1 U14090 ( .A1(n10853), .A2(n10852), .A3(n10851), .A4(n10850), .ZN(
        n10866) );
  AOI22_X1 U14091 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n10674), .B1(
        n14614), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10865) );
  NAND2_X1 U14092 ( .A1(n10665), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n10857) );
  NAND2_X1 U14093 ( .A1(n10496), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n10856) );
  NAND2_X1 U14094 ( .A1(n10485), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n10855) );
  NAND2_X1 U14095 ( .A1(n10673), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n10854) );
  AND4_X1 U14096 ( .A1(n10857), .A2(n10856), .A3(n10855), .A4(n10854), .ZN(
        n10864) );
  INV_X1 U14097 ( .A(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10858) );
  OR2_X1 U14098 ( .A1(n14610), .A2(n10858), .ZN(n10862) );
  INV_X1 U14099 ( .A(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n14580) );
  OR2_X1 U14100 ( .A1(n14609), .A2(n14580), .ZN(n10861) );
  NAND2_X1 U14101 ( .A1(n14613), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n10860) );
  NAND2_X1 U14102 ( .A1(n10667), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n10859) );
  AND4_X1 U14103 ( .A1(n10862), .A2(n10861), .A3(n10860), .A4(n10859), .ZN(
        n10863) );
  NAND4_X1 U14104 ( .A1(n10866), .A2(n10865), .A3(n10864), .A4(n10863), .ZN(
        n14031) );
  INV_X1 U14105 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n10868) );
  AOI22_X1 U14106 ( .A1(n12819), .A2(P2_EAX_REG_14__SCAN_IN), .B1(n10690), 
        .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n10867) );
  OAI21_X1 U14107 ( .B1(n10908), .B2(n10868), .A(n10867), .ZN(n10869) );
  AOI21_X1 U14108 ( .B1(n10870), .B2(n14031), .A(n10869), .ZN(n16050) );
  AOI22_X1 U14109 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n10674), .B1(
        n10667), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10873) );
  AOI22_X1 U14110 ( .A1(n10665), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n14618), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10872) );
  AOI22_X1 U14111 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n10485), .B1(
        n10496), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10871) );
  AND3_X1 U14112 ( .A1(n10873), .A2(n10872), .A3(n10871), .ZN(n10887) );
  AOI22_X1 U14113 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n14598), .B1(
        n14599), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10878) );
  AOI22_X1 U14114 ( .A1(n14579), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n10673), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10877) );
  OR2_X1 U14115 ( .A1(n14601), .A2(n19713), .ZN(n10876) );
  INV_X1 U14116 ( .A(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10874) );
  OR2_X1 U14117 ( .A1(n14603), .A2(n10874), .ZN(n10875) );
  NAND4_X1 U14118 ( .A1(n10878), .A2(n10877), .A3(n10876), .A4(n10875), .ZN(
        n10885) );
  INV_X1 U14119 ( .A(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n10879) );
  OR2_X1 U14120 ( .A1(n14610), .A2(n10879), .ZN(n10883) );
  INV_X1 U14121 ( .A(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n14600) );
  OR2_X1 U14122 ( .A1(n14609), .A2(n14600), .ZN(n10882) );
  NAND2_X1 U14123 ( .A1(n14614), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n10881) );
  NAND2_X1 U14124 ( .A1(n14613), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n10880) );
  NAND4_X1 U14125 ( .A1(n10883), .A2(n10882), .A3(n10881), .A4(n10880), .ZN(
        n10884) );
  NOR2_X1 U14126 ( .A1(n10885), .A2(n10884), .ZN(n10886) );
  NAND2_X1 U14127 ( .A1(n12818), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n10889) );
  AOI22_X1 U14128 ( .A1(n12819), .A2(P2_EAX_REG_15__SCAN_IN), .B1(n10690), 
        .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n10888) );
  OAI211_X1 U14129 ( .C1(n10890), .C2(n14280), .A(n10889), .B(n10888), .ZN(
        n16028) );
  NAND2_X1 U14130 ( .A1(n12818), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n10892) );
  AOI22_X1 U14131 ( .A1(n12819), .A2(P2_EAX_REG_16__SCAN_IN), .B1(n10690), 
        .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n10891) );
  NAND2_X1 U14132 ( .A1(n10892), .A2(n10891), .ZN(n14443) );
  NAND2_X1 U14133 ( .A1(n12818), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n10894) );
  AOI22_X1 U14134 ( .A1(n12819), .A2(P2_EAX_REG_17__SCAN_IN), .B1(n10690), 
        .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n10893) );
  NAND2_X1 U14135 ( .A1(n10894), .A2(n10893), .ZN(n14243) );
  NAND2_X1 U14136 ( .A1(n14445), .A2(n14243), .ZN(n14242) );
  NAND2_X1 U14137 ( .A1(n12818), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n10896) );
  AOI22_X1 U14138 ( .A1(n12819), .A2(P2_EAX_REG_18__SCAN_IN), .B1(n10690), 
        .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n10895) );
  AND2_X1 U14139 ( .A1(n10896), .A2(n10895), .ZN(n15602) );
  NAND2_X1 U14140 ( .A1(n12818), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n10900) );
  AOI22_X1 U14141 ( .A1(n12819), .A2(P2_EAX_REG_19__SCAN_IN), .B1(n10690), 
        .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n10899) );
  NAND2_X1 U14142 ( .A1(n12818), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n10902) );
  AOI22_X1 U14143 ( .A1(n12819), .A2(P2_EAX_REG_20__SCAN_IN), .B1(n10690), 
        .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n10901) );
  NAND2_X1 U14144 ( .A1(n10902), .A2(n10901), .ZN(n15590) );
  NAND2_X1 U14145 ( .A1(n12818), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n10904) );
  AOI22_X1 U14146 ( .A1(n12819), .A2(P2_EAX_REG_21__SCAN_IN), .B1(n10690), 
        .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n10903) );
  NAND2_X1 U14147 ( .A1(n10904), .A2(n10903), .ZN(n11473) );
  NAND2_X1 U14148 ( .A1(n12818), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n10906) );
  AOI22_X1 U14149 ( .A1(n12819), .A2(P2_EAX_REG_22__SCAN_IN), .B1(n10690), 
        .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n10905) );
  NAND2_X1 U14150 ( .A1(n10906), .A2(n10905), .ZN(n15570) );
  INV_X1 U14151 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n19970) );
  AOI22_X1 U14152 ( .A1(n12819), .A2(P2_EAX_REG_23__SCAN_IN), .B1(n10690), 
        .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n10907) );
  OAI21_X1 U14153 ( .B1(n10908), .B2(n19970), .A(n10907), .ZN(n15556) );
  NAND2_X1 U14154 ( .A1(n12818), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n10910) );
  AOI22_X1 U14155 ( .A1(n12819), .A2(P2_EAX_REG_24__SCAN_IN), .B1(n10690), 
        .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n10909) );
  AND2_X1 U14156 ( .A1(n10910), .A2(n10909), .ZN(n15542) );
  NAND2_X1 U14157 ( .A1(n12818), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n10912) );
  AOI22_X1 U14158 ( .A1(n12819), .A2(P2_EAX_REG_25__SCAN_IN), .B1(n10690), 
        .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n10911) );
  AND2_X1 U14159 ( .A1(n10912), .A2(n10911), .ZN(n15523) );
  NAND2_X1 U14160 ( .A1(n12818), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n10914) );
  AOI22_X1 U14161 ( .A1(n12819), .A2(P2_EAX_REG_26__SCAN_IN), .B1(n10690), 
        .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n10913) );
  NAND2_X1 U14162 ( .A1(n10914), .A2(n10913), .ZN(n15718) );
  NAND2_X1 U14163 ( .A1(n10684), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n10916) );
  AOI22_X1 U14164 ( .A1(n12819), .A2(P2_EAX_REG_27__SCAN_IN), .B1(n10690), 
        .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n10915) );
  AND2_X1 U14165 ( .A1(n10916), .A2(n10915), .ZN(n13320) );
  NAND2_X1 U14166 ( .A1(n12818), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n10918) );
  AOI22_X1 U14167 ( .A1(n12819), .A2(P2_EAX_REG_28__SCAN_IN), .B1(n10690), 
        .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n10917) );
  AND2_X1 U14168 ( .A1(n10918), .A2(n10917), .ZN(n15509) );
  NAND2_X1 U14169 ( .A1(n10684), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n10920) );
  AOI22_X1 U14170 ( .A1(n12819), .A2(P2_EAX_REG_29__SCAN_IN), .B1(n10690), 
        .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n10919) );
  NAND2_X1 U14171 ( .A1(n10920), .A2(n10919), .ZN(n12490) );
  NAND2_X1 U14172 ( .A1(n10684), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n10922) );
  AOI22_X1 U14173 ( .A1(n12819), .A2(P2_EAX_REG_30__SCAN_IN), .B1(n10690), 
        .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n10921) );
  NAND2_X1 U14174 ( .A1(n10922), .A2(n10921), .ZN(n10923) );
  INV_X1 U14175 ( .A(n12492), .ZN(n10925) );
  INV_X1 U14176 ( .A(n10923), .ZN(n10924) );
  NAND2_X1 U14177 ( .A1(n10925), .A2(n10924), .ZN(n10926) );
  INV_X1 U14178 ( .A(P2_STATE_REG_1__SCAN_IN), .ZN(n19915) );
  NOR2_X1 U14179 ( .A1(n19915), .A2(n19933), .ZN(n19924) );
  NOR2_X1 U14180 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(P2_STATE_REG_2__SCAN_IN), 
        .ZN(n19927) );
  OR3_X1 U14181 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(n19924), .A3(n19927), .ZN(
        n20063) );
  INV_X1 U14182 ( .A(n14113), .ZN(n10927) );
  NOR2_X1 U14183 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n10927), .ZN(n14128) );
  NOR2_X1 U14184 ( .A1(n16225), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n13328) );
  INV_X1 U14185 ( .A(n13328), .ZN(n13326) );
  NOR3_X1 U14186 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n10928), .A3(n20036), 
        .ZN(n16587) );
  NOR4_X4 U14187 ( .A1(n19170), .A2(n19175), .A3(n16587), .A4(n20056), .ZN(
        n19210) );
  NAND2_X1 U14188 ( .A1(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n19211), .ZN(
        n10933) );
  INV_X1 U14189 ( .A(n14128), .ZN(n10929) );
  AND2_X1 U14190 ( .A1(n13527), .A2(n10929), .ZN(n15487) );
  NOR2_X1 U14191 ( .A1(P2_EBX_REG_31__SCAN_IN), .A2(n13421), .ZN(n10930) );
  AND2_X1 U14192 ( .A1(n11127), .A2(n10930), .ZN(n10931) );
  OR2_X2 U14193 ( .A1(n15487), .A2(n10931), .ZN(n19205) );
  AOI22_X1 U14194 ( .A1(P2_REIP_REG_30__SCAN_IN), .A2(n19210), .B1(
        P2_EBX_REG_30__SCAN_IN), .B2(n19205), .ZN(n10932) );
  OAI211_X1 U14195 ( .C1(n14786), .C2(n19200), .A(n10933), .B(n10932), .ZN(
        n10934) );
  AOI21_X1 U14196 ( .B1(n12803), .B2(n19186), .A(n10934), .ZN(n11130) );
  OR2_X2 U14197 ( .A1(n10942), .A2(n19420), .ZN(n10975) );
  NAND2_X1 U14198 ( .A1(n10983), .A2(n20064), .ZN(n10947) );
  INV_X1 U14199 ( .A(n10942), .ZN(n10944) );
  OAI21_X1 U14200 ( .B1(n10968), .B2(n11487), .A(n11486), .ZN(n10943) );
  NAND2_X1 U14201 ( .A1(n10944), .A2(n10943), .ZN(n10946) );
  NOR2_X1 U14202 ( .A1(n16157), .A2(n10657), .ZN(n10945) );
  NAND2_X1 U14203 ( .A1(n10946), .A2(n10945), .ZN(n11485) );
  INV_X1 U14204 ( .A(n10966), .ZN(n10948) );
  OAI21_X1 U14205 ( .B1(n10935), .B2(n10679), .A(n10948), .ZN(n10949) );
  INV_X1 U14206 ( .A(n10949), .ZN(n11415) );
  NAND2_X1 U14207 ( .A1(n11415), .A2(n10936), .ZN(n11417) );
  NAND2_X1 U14208 ( .A1(n10968), .A2(n10938), .ZN(n11410) );
  AND2_X1 U14209 ( .A1(n11410), .A2(n19420), .ZN(n10950) );
  NAND2_X1 U14210 ( .A1(n11417), .A2(n10950), .ZN(n11483) );
  NAND2_X1 U14211 ( .A1(n11483), .A2(n19391), .ZN(n10953) );
  NAND2_X1 U14212 ( .A1(n10953), .A2(n10952), .ZN(n10982) );
  NAND2_X1 U14213 ( .A1(n19384), .A2(n20062), .ZN(n10957) );
  AND3_X2 U14214 ( .A1(n10955), .A2(n10954), .A3(n13389), .ZN(n14112) );
  INV_X1 U14215 ( .A(n11408), .ZN(n10956) );
  NAND2_X1 U14216 ( .A1(n11013), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10965) );
  INV_X1 U14217 ( .A(n10976), .ZN(n10958) );
  INV_X1 U14218 ( .A(n14104), .ZN(n10963) );
  INV_X2 U14219 ( .A(n11486), .ZN(n11481) );
  INV_X1 U14220 ( .A(n13389), .ZN(n10961) );
  NOR2_X1 U14221 ( .A1(n10961), .A2(n10960), .ZN(n10962) );
  NAND2_X1 U14222 ( .A1(n11492), .A2(n10962), .ZN(n10973) );
  NAND2_X1 U14223 ( .A1(n11469), .A2(n11481), .ZN(n13676) );
  AND2_X1 U14224 ( .A1(n10971), .A2(n10657), .ZN(n20060) );
  NAND2_X1 U14225 ( .A1(n11408), .A2(n20060), .ZN(n14073) );
  AND3_X1 U14226 ( .A1(n11481), .A2(n10072), .A3(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n10977) );
  INV_X1 U14227 ( .A(n14129), .ZN(n10987) );
  OAI22_X1 U14228 ( .A1(n13676), .A2(n14298), .B1(n10987), .B2(n20043), .ZN(
        n10978) );
  INV_X1 U14229 ( .A(n10978), .ZN(n10979) );
  NAND2_X1 U14230 ( .A1(n10980), .A2(n10979), .ZN(n11144) );
  NAND2_X1 U14231 ( .A1(n10982), .A2(n10983), .ZN(n10984) );
  NAND2_X1 U14232 ( .A1(n10981), .A2(n10984), .ZN(n10985) );
  NAND2_X1 U14233 ( .A1(n10985), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10992) );
  NAND2_X1 U14234 ( .A1(n11022), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n10990) );
  NAND2_X1 U14235 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n10986) );
  NAND2_X1 U14236 ( .A1(n11149), .A2(n11168), .ZN(n10997) );
  INV_X1 U14237 ( .A(n10993), .ZN(n10995) );
  NAND2_X1 U14238 ( .A1(n10995), .A2(n10994), .ZN(n10996) );
  NAND2_X2 U14239 ( .A1(n10997), .A2(n10996), .ZN(n11155) );
  NAND2_X1 U14240 ( .A1(n11013), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10999) );
  AOI21_X1 U14241 ( .B1(n14298), .B2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n10998) );
  INV_X1 U14242 ( .A(n11153), .ZN(n11003) );
  NAND2_X1 U14243 ( .A1(n11021), .A2(P2_EBX_REG_2__SCAN_IN), .ZN(n11001) );
  AOI22_X1 U14244 ( .A1(n11022), .A2(P2_REIP_REG_2__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11000) );
  AND2_X1 U14245 ( .A1(n11001), .A2(n11000), .ZN(n11002) );
  INV_X1 U14246 ( .A(n11137), .ZN(n11152) );
  NAND2_X1 U14247 ( .A1(n11005), .A2(n11004), .ZN(n11020) );
  INV_X1 U14248 ( .A(n11016), .ZN(n11014) );
  AND2_X1 U14249 ( .A1(n14129), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n11012) );
  INV_X1 U14250 ( .A(n11015), .ZN(n11017) );
  NAND2_X1 U14251 ( .A1(n11017), .A2(n11016), .ZN(n11018) );
  INV_X1 U14252 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n14269) );
  OR2_X1 U14253 ( .A1(n12815), .A2(n14269), .ZN(n11026) );
  NAND2_X1 U14254 ( .A1(n12812), .A2(P2_EBX_REG_4__SCAN_IN), .ZN(n11024) );
  AOI22_X1 U14255 ( .A1(n12811), .A2(P2_REIP_REG_4__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11023) );
  AND2_X1 U14256 ( .A1(n11024), .A2(n11023), .ZN(n11025) );
  NAND2_X1 U14257 ( .A1(n11026), .A2(n11025), .ZN(n13609) );
  OR2_X1 U14258 ( .A1(n12815), .A2(n14270), .ZN(n11030) );
  NAND2_X1 U14259 ( .A1(n12812), .A2(P2_EBX_REG_5__SCAN_IN), .ZN(n11028) );
  AOI22_X1 U14260 ( .A1(n12811), .A2(P2_REIP_REG_5__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11027) );
  AND2_X1 U14261 ( .A1(n11028), .A2(n11027), .ZN(n11029) );
  INV_X1 U14262 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n14488) );
  OR2_X1 U14263 ( .A1(n12815), .A2(n14488), .ZN(n11034) );
  NAND2_X1 U14264 ( .A1(n12812), .A2(P2_EBX_REG_6__SCAN_IN), .ZN(n11032) );
  INV_X2 U14265 ( .A(n11116), .ZN(n12811) );
  AOI22_X1 U14266 ( .A1(n12811), .A2(P2_REIP_REG_6__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11031) );
  AND2_X1 U14267 ( .A1(n11032), .A2(n11031), .ZN(n11033) );
  NAND2_X1 U14268 ( .A1(n11034), .A2(n11033), .ZN(n13668) );
  OR2_X1 U14269 ( .A1(n12815), .A2(n14421), .ZN(n11038) );
  NAND2_X1 U14270 ( .A1(n12812), .A2(P2_EBX_REG_7__SCAN_IN), .ZN(n11036) );
  AOI22_X1 U14271 ( .A1(n12811), .A2(P2_REIP_REG_7__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11035) );
  AND2_X1 U14272 ( .A1(n11036), .A2(n11035), .ZN(n11037) );
  AOI22_X1 U14273 ( .A1(n12811), .A2(P2_REIP_REG_8__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11040) );
  NAND2_X1 U14274 ( .A1(n12812), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n11039) );
  OAI211_X1 U14275 ( .C1(n12815), .C2(n16573), .A(n11040), .B(n11039), .ZN(
        n13819) );
  OR2_X1 U14276 ( .A1(n12815), .A2(n16072), .ZN(n11044) );
  NAND2_X1 U14277 ( .A1(n12812), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n11042) );
  AOI22_X1 U14278 ( .A1(n12811), .A2(P2_REIP_REG_9__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n11041) );
  AND2_X1 U14279 ( .A1(n11042), .A2(n11041), .ZN(n11043) );
  INV_X1 U14280 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16088) );
  OR2_X1 U14281 ( .A1(n12815), .A2(n16088), .ZN(n11048) );
  NAND2_X1 U14282 ( .A1(n12812), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n11046) );
  AOI22_X1 U14283 ( .A1(n12811), .A2(P2_REIP_REG_10__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), 
        .ZN(n11045) );
  AND2_X1 U14284 ( .A1(n11046), .A2(n11045), .ZN(n11047) );
  NAND2_X1 U14285 ( .A1(n11048), .A2(n11047), .ZN(n13707) );
  OR2_X1 U14286 ( .A1(n12815), .A2(n16080), .ZN(n11052) );
  NAND2_X1 U14287 ( .A1(n12812), .A2(P2_EBX_REG_11__SCAN_IN), .ZN(n11050) );
  AOI22_X1 U14288 ( .A1(n12811), .A2(P2_REIP_REG_11__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), 
        .ZN(n11049) );
  AND2_X1 U14289 ( .A1(n11050), .A2(n11049), .ZN(n11051) );
  OR2_X1 U14290 ( .A1(n12815), .A2(n16570), .ZN(n11057) );
  NAND2_X1 U14291 ( .A1(n12812), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n11055) );
  AOI22_X1 U14292 ( .A1(n12811), .A2(P2_REIP_REG_12__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), 
        .ZN(n11054) );
  AND2_X1 U14293 ( .A1(n11055), .A2(n11054), .ZN(n11056) );
  NAND2_X1 U14294 ( .A1(n11057), .A2(n11056), .ZN(n13827) );
  NAND2_X1 U14295 ( .A1(n13811), .A2(n13827), .ZN(n13826) );
  INV_X1 U14296 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16062) );
  OR2_X1 U14297 ( .A1(n12815), .A2(n16062), .ZN(n11060) );
  AOI22_X1 U14298 ( .A1(n12811), .A2(P2_REIP_REG_13__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), 
        .ZN(n11059) );
  NAND2_X1 U14299 ( .A1(n12812), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n11058) );
  INV_X1 U14300 ( .A(n11061), .ZN(n14027) );
  INV_X1 U14301 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n16049) );
  OR2_X1 U14302 ( .A1(n12815), .A2(n16049), .ZN(n11064) );
  AOI22_X1 U14303 ( .A1(n12811), .A2(P2_REIP_REG_14__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), 
        .ZN(n11063) );
  NAND2_X1 U14304 ( .A1(n12812), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n11062) );
  OR2_X1 U14305 ( .A1(n12815), .A2(n16034), .ZN(n11068) );
  NAND2_X1 U14306 ( .A1(n12812), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n11066) );
  AOI22_X1 U14307 ( .A1(n12811), .A2(P2_REIP_REG_15__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), 
        .ZN(n11065) );
  AND2_X1 U14308 ( .A1(n11066), .A2(n11065), .ZN(n11067) );
  NAND2_X1 U14309 ( .A1(n11068), .A2(n11067), .ZN(n14282) );
  OR2_X1 U14310 ( .A1(n12815), .A2(n16491), .ZN(n11072) );
  NAND2_X1 U14311 ( .A1(n12812), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n11070) );
  AOI22_X1 U14312 ( .A1(n12811), .A2(P2_REIP_REG_16__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), 
        .ZN(n11069) );
  AND2_X1 U14313 ( .A1(n11070), .A2(n11069), .ZN(n11071) );
  NAND2_X1 U14314 ( .A1(n11072), .A2(n11071), .ZN(n14252) );
  NAND2_X1 U14315 ( .A1(n14251), .A2(n14252), .ZN(n14250) );
  OR2_X1 U14316 ( .A1(n12815), .A2(n15990), .ZN(n11075) );
  AOI22_X1 U14317 ( .A1(n12811), .A2(P2_REIP_REG_17__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), 
        .ZN(n11074) );
  NAND2_X1 U14318 ( .A1(n12812), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n11073) );
  NAND2_X1 U14319 ( .A1(n11053), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n11079) );
  NAND2_X1 U14320 ( .A1(n12812), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n11077) );
  AOI22_X1 U14321 ( .A1(n12811), .A2(P2_REIP_REG_18__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), 
        .ZN(n11076) );
  AND2_X1 U14322 ( .A1(n11077), .A2(n11076), .ZN(n11078) );
  NAND2_X1 U14323 ( .A1(n11053), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n11082) );
  INV_X1 U14324 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n19962) );
  OAI22_X1 U14325 ( .A1(n11116), .A2(n19962), .B1(n13362), .B2(n19064), .ZN(
        n11080) );
  AOI21_X1 U14326 ( .B1(n12812), .B2(P2_EBX_REG_19__SCAN_IN), .A(n11080), .ZN(
        n11081) );
  OR2_X1 U14327 ( .A1(n12815), .A2(n15963), .ZN(n11086) );
  NAND2_X1 U14328 ( .A1(n12812), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n11084) );
  AOI22_X1 U14329 ( .A1(n12811), .A2(P2_REIP_REG_20__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), 
        .ZN(n11083) );
  AND2_X1 U14330 ( .A1(n11084), .A2(n11083), .ZN(n11085) );
  NAND2_X1 U14331 ( .A1(n11086), .A2(n11085), .ZN(n15588) );
  NAND2_X1 U14332 ( .A1(n11053), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n11089) );
  INV_X1 U14333 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n19966) );
  OAI22_X1 U14334 ( .A1(n11116), .A2(n19966), .B1(n13362), .B2(n15808), .ZN(
        n11087) );
  AOI21_X1 U14335 ( .B1(n12812), .B2(P2_EBX_REG_21__SCAN_IN), .A(n11087), .ZN(
        n11088) );
  INV_X1 U14336 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15938) );
  OR2_X1 U14337 ( .A1(n12815), .A2(n15938), .ZN(n11092) );
  AOI22_X1 U14338 ( .A1(n12811), .A2(P2_REIP_REG_22__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), 
        .ZN(n11091) );
  NAND2_X1 U14339 ( .A1(n12812), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n11090) );
  INV_X1 U14340 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n21278) );
  OR2_X1 U14341 ( .A1(n12815), .A2(n21278), .ZN(n11096) );
  NAND2_X1 U14342 ( .A1(n12812), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n11094) );
  AOI22_X1 U14343 ( .A1(n12811), .A2(P2_REIP_REG_23__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), 
        .ZN(n11093) );
  AND2_X1 U14344 ( .A1(n11094), .A2(n11093), .ZN(n11095) );
  NAND2_X1 U14345 ( .A1(n11096), .A2(n11095), .ZN(n15554) );
  OR2_X1 U14346 ( .A1(n12815), .A2(n15922), .ZN(n11100) );
  NAND2_X1 U14347 ( .A1(n12812), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n11098) );
  AOI22_X1 U14348 ( .A1(n12811), .A2(P2_REIP_REG_24__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), 
        .ZN(n11097) );
  AND2_X1 U14349 ( .A1(n11098), .A2(n11097), .ZN(n11099) );
  NAND2_X1 U14350 ( .A1(n11100), .A2(n11099), .ZN(n15538) );
  NAND2_X1 U14351 ( .A1(n11053), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n11103) );
  INV_X1 U14352 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n19973) );
  OAI22_X1 U14353 ( .A1(n11116), .A2(n19973), .B1(n13362), .B2(n15788), .ZN(
        n11101) );
  AOI21_X1 U14354 ( .B1(n12812), .B2(P2_EBX_REG_25__SCAN_IN), .A(n11101), .ZN(
        n11102) );
  NAND2_X1 U14355 ( .A1(n11053), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11107) );
  NAND2_X1 U14356 ( .A1(n12812), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n11105) );
  AOI22_X1 U14357 ( .A1(n12811), .A2(P2_REIP_REG_26__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), 
        .ZN(n11104) );
  AND2_X1 U14358 ( .A1(n11105), .A2(n11104), .ZN(n11106) );
  INV_X1 U14359 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15764) );
  OR2_X1 U14360 ( .A1(n12815), .A2(n15764), .ZN(n11111) );
  NAND2_X1 U14361 ( .A1(n12812), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n11109) );
  AOI22_X1 U14362 ( .A1(n12811), .A2(P2_REIP_REG_27__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), 
        .ZN(n11108) );
  AND2_X1 U14363 ( .A1(n11109), .A2(n11108), .ZN(n11110) );
  NAND2_X1 U14364 ( .A1(n11111), .A2(n11110), .ZN(n13318) );
  INV_X1 U14365 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n12474) );
  OR2_X1 U14366 ( .A1(n12815), .A2(n12474), .ZN(n11115) );
  NAND2_X1 U14367 ( .A1(n12812), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n11113) );
  AOI22_X1 U14368 ( .A1(n12811), .A2(P2_REIP_REG_28__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), 
        .ZN(n11112) );
  AND2_X1 U14369 ( .A1(n11113), .A2(n11112), .ZN(n11114) );
  NAND2_X1 U14370 ( .A1(n11115), .A2(n11114), .ZN(n15504) );
  NAND2_X1 U14371 ( .A1(n13316), .A2(n15504), .ZN(n12486) );
  NAND2_X1 U14372 ( .A1(n11053), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n11119) );
  INV_X1 U14373 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n19981) );
  OAI22_X1 U14374 ( .A1(n11116), .A2(n19981), .B1(n13362), .B2(n12790), .ZN(
        n11117) );
  AOI21_X1 U14375 ( .B1(n12812), .B2(P2_EBX_REG_29__SCAN_IN), .A(n11117), .ZN(
        n11118) );
  NAND2_X1 U14376 ( .A1(n11053), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11123) );
  NAND2_X1 U14377 ( .A1(n12812), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n11121) );
  AOI22_X1 U14378 ( .A1(n12811), .A2(P2_REIP_REG_30__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), 
        .ZN(n11120) );
  AND2_X1 U14379 ( .A1(n11121), .A2(n11120), .ZN(n11122) );
  AND2_X1 U14380 ( .A1(n11123), .A2(n11122), .ZN(n11124) );
  NAND2_X1 U14381 ( .A1(n12489), .A2(n11124), .ZN(n11125) );
  NAND2_X1 U14382 ( .A1(n12817), .A2(n11125), .ZN(n14789) );
  INV_X1 U14383 ( .A(n11126), .ZN(n11128) );
  NAND2_X1 U14384 ( .A1(n11132), .A2(n11131), .ZN(P2_U2825) );
  AND3_X1 U14385 ( .A1(n11133), .A2(P2_EBX_REG_21__SCAN_IN), .A3(n10543), .ZN(
        n11134) );
  OR2_X1 U14386 ( .A1(n11135), .A2(n11134), .ZN(n15583) );
  INV_X1 U14387 ( .A(n15583), .ZN(n11136) );
  NAND2_X1 U14388 ( .A1(n11136), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12435) );
  INV_X1 U14389 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n11516) );
  OAI21_X1 U14390 ( .B1(n15583), .B2(n11254), .A(n11516), .ZN(n12429) );
  OAI21_X1 U14391 ( .B1(n12435), .B2(n11254), .A(n12429), .ZN(n11362) );
  INV_X1 U14392 ( .A(n11139), .ZN(n11140) );
  NAND2_X1 U14393 ( .A1(n11155), .A2(n11142), .ZN(n11143) );
  INV_X1 U14394 ( .A(n11144), .ZN(n11147) );
  INV_X1 U14395 ( .A(n11145), .ZN(n11146) );
  NAND2_X1 U14396 ( .A1(n11147), .A2(n11146), .ZN(n11148) );
  INV_X1 U14397 ( .A(n11167), .ZN(n11150) );
  NAND2_X1 U14398 ( .A1(n14093), .A2(n11150), .ZN(n11157) );
  INV_X1 U14399 ( .A(n11157), .ZN(n11151) );
  XNOR2_X1 U14400 ( .A(n11153), .B(n11152), .ZN(n11154) );
  XNOR2_X2 U14401 ( .A(n11155), .B(n11154), .ZN(n13564) );
  NAND2_X1 U14402 ( .A1(n14093), .A2(n11167), .ZN(n11159) );
  INV_X1 U14403 ( .A(n11159), .ZN(n11156) );
  AOI22_X1 U14404 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19672), .B1(
        n19715), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11166) );
  AOI22_X1 U14405 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19433), .B1(
        n11207), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11165) );
  AND2_X2 U14406 ( .A1(n11160), .A2(n19342), .ZN(n11209) );
  AOI22_X1 U14407 ( .A1(n11208), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n11209), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11164) );
  AOI22_X1 U14408 ( .A1(n19605), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n11210), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11163) );
  AND4_X1 U14409 ( .A1(n11166), .A2(n11165), .A3(n11164), .A4(n11163), .ZN(
        n11182) );
  INV_X1 U14410 ( .A(n14093), .ZN(n19198) );
  AOI22_X1 U14411 ( .A1(n11222), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n11223), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11181) );
  INV_X1 U14412 ( .A(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11170) );
  INV_X2 U14413 ( .A(n11188), .ZN(n19373) );
  INV_X1 U14414 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11174) );
  NAND2_X1 U14415 ( .A1(n19461), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n11173) );
  OAI21_X1 U14416 ( .B1(n19373), .B2(n11174), .A(n11173), .ZN(n11175) );
  NOR2_X1 U14417 ( .A1(n11176), .A2(n11175), .ZN(n11180) );
  INV_X1 U14418 ( .A(n19572), .ZN(n11224) );
  AOI22_X1 U14419 ( .A1(n11224), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11225), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11179) );
  NAND2_X1 U14420 ( .A1(n11183), .A2(n9839), .ZN(n11184) );
  NAND2_X1 U14421 ( .A1(n11222), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n11187) );
  NAND2_X1 U14422 ( .A1(n11225), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n11186) );
  NAND2_X1 U14423 ( .A1(n11187), .A2(n11186), .ZN(n11194) );
  NAND2_X1 U14424 ( .A1(n11223), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n11192) );
  NAND2_X1 U14425 ( .A1(n11216), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n11190) );
  NAND2_X1 U14426 ( .A1(n11192), .A2(n11191), .ZN(n11193) );
  NOR2_X1 U14427 ( .A1(n11194), .A2(n11193), .ZN(n11204) );
  AOI22_X1 U14428 ( .A1(n19461), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n11207), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11198) );
  AOI22_X1 U14429 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19605), .B1(
        n11208), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11197) );
  AOI22_X1 U14430 ( .A1(n19433), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n11210), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11196) );
  AOI22_X1 U14431 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19672), .B1(
        n11209), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11195) );
  AND4_X1 U14432 ( .A1(n11198), .A2(n11197), .A3(n11196), .A4(n11195), .ZN(
        n11203) );
  AOI21_X1 U14433 ( .B1(n19715), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A(
        n9839), .ZN(n11200) );
  NAND2_X1 U14434 ( .A1(n11217), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n11199) );
  OAI211_X1 U14435 ( .C1(n19572), .C2(n19586), .A(n11200), .B(n11199), .ZN(
        n11201) );
  INV_X1 U14436 ( .A(n11201), .ZN(n11202) );
  NAND3_X1 U14437 ( .A1(n11204), .A2(n11203), .A3(n11202), .ZN(n11206) );
  OR2_X1 U14438 ( .A1(n11429), .A2(n20062), .ZN(n13344) );
  NOR2_X1 U14439 ( .A1(n13344), .A2(n11428), .ZN(n11432) );
  AOI22_X1 U14440 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19433), .B1(
        n11207), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11214) );
  AOI22_X1 U14441 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19672), .B1(
        n19715), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11213) );
  AOI22_X1 U14442 ( .A1(n11208), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n11209), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11212) );
  AOI22_X1 U14443 ( .A1(n19605), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11210), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11211) );
  INV_X1 U14444 ( .A(n19461), .ZN(n11241) );
  OR2_X1 U14445 ( .A1(n11241), .A2(n11215), .ZN(n11221) );
  OR2_X1 U14446 ( .A1(n19373), .A2(n13669), .ZN(n11220) );
  NAND2_X1 U14447 ( .A1(n11216), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n11219) );
  NAND2_X1 U14448 ( .A1(n11217), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n11218) );
  AOI22_X1 U14449 ( .A1(n11222), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11223), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11227) );
  AOI22_X1 U14450 ( .A1(n11224), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11225), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11226) );
  NAND4_X1 U14451 ( .A1(n11229), .A2(n11228), .A3(n11227), .A4(n11226), .ZN(
        n11233) );
  INV_X1 U14452 ( .A(n11230), .ZN(n11231) );
  NAND2_X1 U14453 ( .A1(n11231), .A2(n9839), .ZN(n11232) );
  AOI22_X1 U14454 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n11207), .B1(
        n11208), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11237) );
  AOI22_X1 U14455 ( .A1(n19605), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n11210), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11236) );
  AOI22_X1 U14456 ( .A1(n19433), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n19672), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11235) );
  AOI22_X1 U14457 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n11209), .B1(
        n19715), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11234) );
  AOI22_X1 U14458 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n11222), .B1(
        n11224), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11248) );
  INV_X1 U14459 ( .A(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11240) );
  INV_X1 U14460 ( .A(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11239) );
  OAI22_X1 U14461 ( .A1(n11241), .A2(n11240), .B1(n11238), .B2(n11239), .ZN(
        n11245) );
  INV_X1 U14462 ( .A(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11243) );
  OAI22_X1 U14463 ( .A1(n19373), .A2(n11243), .B1(n14295), .B2(n11242), .ZN(
        n11244) );
  NOR2_X1 U14464 ( .A1(n11245), .A2(n11244), .ZN(n11247) );
  AOI22_X1 U14465 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n11225), .B1(
        n11223), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11246) );
  NAND4_X1 U14466 ( .A1(n11249), .A2(n11248), .A3(n11247), .A4(n11246), .ZN(
        n11252) );
  NAND2_X1 U14467 ( .A1(n9839), .A2(n11250), .ZN(n11251) );
  INV_X1 U14468 ( .A(n11255), .ZN(n11300) );
  XNOR2_X1 U14469 ( .A(n11301), .B(n11300), .ZN(n19153) );
  INV_X1 U14470 ( .A(n11271), .ZN(n11257) );
  OAI21_X1 U14471 ( .B1(n11264), .B2(n11258), .A(n11257), .ZN(n14068) );
  OAI21_X1 U14472 ( .B1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n20043), .A(
        n11260), .ZN(n11391) );
  MUX2_X1 U14473 ( .A(n11391), .B(n11429), .S(n10072), .Z(n11396) );
  INV_X1 U14474 ( .A(P2_EBX_REG_0__SCAN_IN), .ZN(n11261) );
  MUX2_X1 U14475 ( .A(n11396), .B(n11261), .S(n10543), .Z(n19201) );
  NOR2_X1 U14476 ( .A1(n19201), .A2(n16105), .ZN(n13341) );
  INV_X1 U14477 ( .A(n13341), .ZN(n13333) );
  NAND3_X1 U14478 ( .A1(n10543), .A2(P2_EBX_REG_0__SCAN_IN), .A3(
        P2_EBX_REG_1__SCAN_IN), .ZN(n11262) );
  NAND2_X1 U14479 ( .A1(n11265), .A2(n11262), .ZN(n19184) );
  NOR2_X1 U14480 ( .A1(n13333), .A2(n19184), .ZN(n11263) );
  NAND2_X1 U14481 ( .A1(n13333), .A2(n19184), .ZN(n13332) );
  OAI21_X1 U14482 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n11263), .A(
        n13332), .ZN(n14802) );
  INV_X1 U14483 ( .A(n11264), .ZN(n11268) );
  NAND2_X1 U14484 ( .A1(n11266), .A2(n11265), .ZN(n11267) );
  NAND2_X1 U14485 ( .A1(n11268), .A2(n11267), .ZN(n14201) );
  XNOR2_X1 U14486 ( .A(n14201), .B(n11499), .ZN(n14801) );
  OR2_X1 U14487 ( .A1(n14802), .A2(n14801), .ZN(n14799) );
  INV_X1 U14488 ( .A(n14201), .ZN(n11269) );
  NAND2_X1 U14489 ( .A1(n11269), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11270) );
  NAND2_X1 U14490 ( .A1(n14799), .A2(n11270), .ZN(n13868) );
  XNOR2_X1 U14491 ( .A(n11272), .B(n11271), .ZN(n11273) );
  INV_X1 U14492 ( .A(n11273), .ZN(n14190) );
  NAND2_X1 U14493 ( .A1(n14190), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11274) );
  NAND2_X1 U14494 ( .A1(n11275), .A2(n11274), .ZN(n14263) );
  INV_X1 U14495 ( .A(n11301), .ZN(n11279) );
  NAND2_X1 U14496 ( .A1(n11277), .A2(n11276), .ZN(n11278) );
  NAND2_X1 U14497 ( .A1(n11279), .A2(n11278), .ZN(n19168) );
  AND2_X1 U14498 ( .A1(n19168), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11283) );
  AND2_X1 U14499 ( .A1(n11254), .A2(n14270), .ZN(n11284) );
  INV_X1 U14500 ( .A(n11284), .ZN(n11280) );
  NAND2_X1 U14501 ( .A1(n11290), .A2(n11280), .ZN(n11281) );
  NAND2_X1 U14502 ( .A1(n11282), .A2(n11281), .ZN(n11289) );
  MUX2_X1 U14503 ( .A(n11284), .B(n11283), .S(n11290), .Z(n11285) );
  NAND2_X1 U14504 ( .A1(n11285), .A2(n11291), .ZN(n11288) );
  OAI21_X1 U14505 ( .B1(n11254), .B2(n14270), .A(n19168), .ZN(n11286) );
  OAI21_X1 U14506 ( .B1(n19168), .B2(n14270), .A(n11286), .ZN(n11287) );
  OAI211_X1 U14507 ( .C1(n11291), .C2(n11289), .A(n11288), .B(n11287), .ZN(
        n14262) );
  NAND2_X1 U14508 ( .A1(n14263), .A2(n14262), .ZN(n11294) );
  OAI21_X1 U14509 ( .B1(n11446), .B2(n12808), .A(n19168), .ZN(n11292) );
  NAND2_X1 U14510 ( .A1(n11292), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11293) );
  NAND2_X1 U14511 ( .A1(n11294), .A2(n11293), .ZN(n14485) );
  NAND2_X1 U14512 ( .A1(n14484), .A2(n14485), .ZN(n11297) );
  NAND2_X1 U14513 ( .A1(n11295), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11296) );
  OAI21_X1 U14514 ( .B1(n11299), .B2(n11298), .A(n9890), .ZN(n14162) );
  OR2_X1 U14515 ( .A1(n14162), .A2(n11458), .ZN(n16530) );
  INV_X1 U14516 ( .A(n11299), .ZN(n11305) );
  NAND2_X1 U14517 ( .A1(n11301), .A2(n11300), .ZN(n11303) );
  NAND2_X1 U14518 ( .A1(n11303), .A2(n11302), .ZN(n11304) );
  NAND2_X1 U14519 ( .A1(n11305), .A2(n11304), .ZN(n19145) );
  OR2_X1 U14520 ( .A1(n19145), .A2(n14421), .ZN(n16532) );
  NAND2_X1 U14521 ( .A1(n16530), .A2(n16532), .ZN(n11306) );
  NAND3_X1 U14522 ( .A1(n11307), .A2(P2_EBX_REG_10__SCAN_IN), .A3(n10543), 
        .ZN(n11308) );
  OAI211_X1 U14523 ( .C1(n11307), .C2(P2_EBX_REG_10__SCAN_IN), .A(n11308), .B(
        n12460), .ZN(n14175) );
  OR2_X1 U14524 ( .A1(n14175), .A2(n11254), .ZN(n11309) );
  NAND2_X1 U14525 ( .A1(n11309), .A2(n16088), .ZN(n16094) );
  OR2_X1 U14526 ( .A1(n14162), .A2(n11254), .ZN(n11310) );
  NAND2_X1 U14527 ( .A1(n11310), .A2(n16573), .ZN(n16531) );
  NAND2_X1 U14528 ( .A1(n19145), .A2(n14421), .ZN(n16534) );
  AND2_X1 U14529 ( .A1(n16531), .A2(n16534), .ZN(n14539) );
  NAND2_X1 U14530 ( .A1(n10543), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n11311) );
  XNOR2_X1 U14531 ( .A(n9890), .B(n11311), .ZN(n19134) );
  NAND2_X1 U14532 ( .A1(n19134), .A2(n12808), .ZN(n11312) );
  NAND2_X1 U14533 ( .A1(n11312), .A2(n16072), .ZN(n16089) );
  AND3_X1 U14534 ( .A1(n16094), .A2(n14539), .A3(n16089), .ZN(n11313) );
  INV_X1 U14535 ( .A(n14175), .ZN(n11315) );
  NOR2_X1 U14536 ( .A1(n11254), .A2(n16088), .ZN(n11314) );
  NAND2_X1 U14537 ( .A1(n11315), .A2(n11314), .ZN(n16093) );
  NOR2_X1 U14538 ( .A1(n11254), .A2(n16072), .ZN(n11316) );
  NAND2_X1 U14539 ( .A1(n19134), .A2(n11316), .ZN(n16090) );
  AND3_X1 U14540 ( .A1(n10543), .A2(P2_EBX_REG_11__SCAN_IN), .A3(n9940), .ZN(
        n11317) );
  NOR2_X1 U14541 ( .A1(n11318), .A2(n11317), .ZN(n19120) );
  NAND2_X1 U14542 ( .A1(n19120), .A2(n12808), .ZN(n15865) );
  NAND2_X1 U14543 ( .A1(n10188), .A2(n11320), .ZN(n11321) );
  NAND2_X1 U14544 ( .A1(n11326), .A2(n11321), .ZN(n15615) );
  XNOR2_X1 U14545 ( .A(n11322), .B(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n16514) );
  NAND2_X1 U14546 ( .A1(n11322), .A2(n16570), .ZN(n11323) );
  NAND2_X1 U14547 ( .A1(n11326), .A2(n11325), .ZN(n11327) );
  AND2_X1 U14548 ( .A1(n11330), .A2(n11327), .ZN(n19110) );
  NAND2_X1 U14549 ( .A1(n19110), .A2(n12808), .ZN(n11332) );
  INV_X1 U14550 ( .A(n11332), .ZN(n11328) );
  NAND2_X1 U14551 ( .A1(n11328), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n15850) );
  NAND2_X1 U14552 ( .A1(n12442), .A2(n15850), .ZN(n16041) );
  AND2_X1 U14553 ( .A1(n11330), .A2(n11329), .ZN(n11331) );
  OR2_X1 U14554 ( .A1(n11331), .A2(n11338), .ZN(n19100) );
  OAI21_X1 U14555 ( .B1(n19100), .B2(n11254), .A(n16049), .ZN(n16039) );
  NAND2_X1 U14556 ( .A1(n11332), .A2(n16062), .ZN(n16040) );
  NAND2_X1 U14557 ( .A1(n16039), .A2(n16040), .ZN(n12427) );
  INV_X1 U14558 ( .A(n12427), .ZN(n11335) );
  INV_X1 U14559 ( .A(n19100), .ZN(n11334) );
  NOR2_X1 U14560 ( .A1(n11254), .A2(n16049), .ZN(n11333) );
  NAND2_X1 U14561 ( .A1(n11334), .A2(n11333), .ZN(n16038) );
  INV_X1 U14562 ( .A(n11336), .ZN(n11337) );
  XNOR2_X1 U14563 ( .A(n11338), .B(n11337), .ZN(n19089) );
  AOI21_X1 U14564 ( .B1(n19089), .B2(n12808), .A(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n16023) );
  NOR2_X1 U14565 ( .A1(n11254), .A2(n16034), .ZN(n11339) );
  NAND2_X1 U14566 ( .A1(n19089), .A2(n11339), .ZN(n12436) );
  NAND3_X1 U14567 ( .A1(n11341), .A2(P2_EBX_REG_16__SCAN_IN), .A3(n10543), 
        .ZN(n11340) );
  OAI211_X1 U14568 ( .C1(n11341), .C2(P2_EBX_REG_16__SCAN_IN), .A(n11340), .B(
        n12460), .ZN(n14452) );
  OR2_X1 U14569 ( .A1(n14452), .A2(n11254), .ZN(n11342) );
  XNOR2_X1 U14570 ( .A(n11342), .B(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n16015) );
  OR2_X1 U14571 ( .A1(n14452), .A2(n16491), .ZN(n12432) );
  INV_X1 U14572 ( .A(n11343), .ZN(n11344) );
  XNOR2_X1 U14573 ( .A(n9888), .B(n11344), .ZN(n19077) );
  NAND2_X1 U14574 ( .A1(n19077), .A2(n12808), .ZN(n11345) );
  NAND2_X1 U14575 ( .A1(n11345), .A2(n15990), .ZN(n15841) );
  NOR2_X1 U14576 ( .A1(n11254), .A2(n15990), .ZN(n11346) );
  NAND2_X1 U14577 ( .A1(n19077), .A2(n11346), .ZN(n15840) );
  INV_X1 U14578 ( .A(n15840), .ZN(n11347) );
  NOR2_X1 U14579 ( .A1(n11349), .A2(n11348), .ZN(n11350) );
  OR2_X1 U14580 ( .A1(n11354), .A2(n11350), .ZN(n15610) );
  INV_X1 U14581 ( .A(n15610), .ZN(n11351) );
  NAND2_X1 U14582 ( .A1(n11351), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n12433) );
  OR2_X1 U14583 ( .A1(n12433), .A2(n11254), .ZN(n15987) );
  NOR2_X1 U14584 ( .A1(n11354), .A2(n11353), .ZN(n11355) );
  OR2_X1 U14585 ( .A1(n11352), .A2(n11355), .ZN(n19065) );
  INV_X1 U14586 ( .A(n19065), .ZN(n11356) );
  NAND2_X1 U14587 ( .A1(n11356), .A2(n12808), .ZN(n11360) );
  INV_X1 U14588 ( .A(n11360), .ZN(n11357) );
  NAND2_X1 U14589 ( .A1(n11357), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15830) );
  INV_X1 U14590 ( .A(n15830), .ZN(n11358) );
  AND2_X1 U14591 ( .A1(n10543), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n11359) );
  XNOR2_X1 U14592 ( .A(n11352), .B(n11359), .ZN(n15595) );
  NAND2_X1 U14593 ( .A1(n15595), .A2(n12808), .ZN(n11361) );
  AND2_X1 U14594 ( .A1(n11361), .A2(n15963), .ZN(n15818) );
  INV_X1 U14595 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15980) );
  NAND2_X1 U14596 ( .A1(n11360), .A2(n15980), .ZN(n15829) );
  INV_X1 U14597 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n15835) );
  OAI21_X1 U14598 ( .B1(n15610), .B2(n11254), .A(n15835), .ZN(n15986) );
  NAND2_X1 U14599 ( .A1(n15829), .A2(n15986), .ZN(n15815) );
  OR2_X1 U14600 ( .A1(n15818), .A2(n15815), .ZN(n12430) );
  OR2_X1 U14601 ( .A1(n11361), .A2(n15963), .ZN(n15817) );
  NOR2_X1 U14602 ( .A1(n11363), .A2(n11379), .ZN(n11364) );
  OR2_X1 U14603 ( .A1(n11402), .A2(n11364), .ZN(n11381) );
  NAND2_X1 U14604 ( .A1(n11366), .A2(n11365), .ZN(n11399) );
  INV_X1 U14605 ( .A(n11397), .ZN(n11367) );
  OAI21_X1 U14606 ( .B1(n11391), .B2(n11367), .A(n10072), .ZN(n11371) );
  INV_X1 U14607 ( .A(n11391), .ZN(n11369) );
  OAI211_X1 U14608 ( .C1(n20062), .C2(n11369), .A(n20064), .B(n11368), .ZN(
        n11370) );
  OAI211_X1 U14609 ( .C1(n11372), .C2(n11373), .A(n11371), .B(n11370), .ZN(
        n11377) );
  NAND2_X1 U14610 ( .A1(n11384), .A2(n20062), .ZN(n11374) );
  MUX2_X1 U14611 ( .A(n11379), .B(n11374), .S(n11373), .Z(n11376) );
  AOI21_X1 U14612 ( .B1(n11377), .B2(n11376), .A(n11375), .ZN(n11378) );
  AOI21_X1 U14613 ( .B1(n11399), .B2(n11379), .A(n11378), .ZN(n11380) );
  NOR2_X1 U14614 ( .A1(n11381), .A2(n11380), .ZN(n11382) );
  MUX2_X1 U14615 ( .A(n11383), .B(n11382), .S(P2_STATE2_REG_0__SCAN_IN), .Z(
        n11387) );
  INV_X1 U14616 ( .A(n11384), .ZN(n13363) );
  NAND2_X1 U14617 ( .A1(n11402), .A2(n13363), .ZN(n11385) );
  NAND2_X1 U14618 ( .A1(n14108), .A2(n20062), .ZN(n13692) );
  OAI211_X1 U14619 ( .C1(n10657), .C2(n11387), .A(n13692), .B(n10938), .ZN(
        n11425) );
  NAND2_X1 U14620 ( .A1(n11487), .A2(n14113), .ZN(n11388) );
  OR2_X1 U14621 ( .A1(n13692), .A2(n11388), .ZN(n11424) );
  INV_X1 U14622 ( .A(n11389), .ZN(n11390) );
  INV_X1 U14623 ( .A(n14115), .ZN(n14111) );
  OAI21_X1 U14624 ( .B1(n11391), .B2(n11390), .A(n14111), .ZN(n11395) );
  NAND2_X1 U14625 ( .A1(n10436), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11392) );
  NAND2_X1 U14626 ( .A1(n11392), .A2(n11383), .ZN(n16155) );
  INV_X1 U14627 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n11393) );
  OAI21_X1 U14628 ( .B1(n10496), .B2(n16155), .A(n11393), .ZN(n11394) );
  NAND2_X1 U14629 ( .A1(n11394), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n20035) );
  OAI21_X1 U14630 ( .B1(n11395), .B2(P2_STATE2_REG_1__SCAN_IN), .A(n20035), 
        .ZN(n20047) );
  NAND3_X1 U14631 ( .A1(n20047), .A2(n14112), .A3(n20062), .ZN(n11406) );
  INV_X1 U14632 ( .A(n11396), .ZN(n11398) );
  NAND2_X1 U14633 ( .A1(n11398), .A2(n11397), .ZN(n11401) );
  AOI21_X1 U14634 ( .B1(n11401), .B2(n11400), .A(n11399), .ZN(n11403) );
  OR2_X1 U14635 ( .A1(n11403), .A2(n11402), .ZN(n20048) );
  INV_X1 U14636 ( .A(n20048), .ZN(n11404) );
  NAND2_X1 U14637 ( .A1(n11404), .A2(n20049), .ZN(n11405) );
  NAND2_X1 U14638 ( .A1(n11406), .A2(n11405), .ZN(n12786) );
  MUX2_X1 U14639 ( .A(n11408), .B(n11487), .S(n9839), .Z(n11407) );
  NAND2_X1 U14640 ( .A1(n11407), .A2(n20069), .ZN(n11421) );
  NAND2_X1 U14641 ( .A1(n11408), .A2(n14113), .ZN(n11409) );
  OR2_X1 U14642 ( .A1(n14115), .A2(n11409), .ZN(n11420) );
  AND2_X1 U14643 ( .A1(n11410), .A2(n19384), .ZN(n11414) );
  NAND2_X1 U14644 ( .A1(n10938), .A2(n9839), .ZN(n11477) );
  NAND2_X1 U14645 ( .A1(n11477), .A2(n20064), .ZN(n11411) );
  NAND2_X1 U14646 ( .A1(n11411), .A2(n19420), .ZN(n11412) );
  AOI21_X1 U14647 ( .B1(n11412), .B2(n19384), .A(n11481), .ZN(n11413) );
  OAI21_X1 U14648 ( .B1(n13686), .B2(n11414), .A(n11413), .ZN(n11480) );
  OR2_X1 U14649 ( .A1(n11415), .A2(n10937), .ZN(n11416) );
  NAND2_X1 U14650 ( .A1(n11416), .A2(n20060), .ZN(n11484) );
  NAND2_X1 U14651 ( .A1(n11484), .A2(n11417), .ZN(n11418) );
  NOR2_X1 U14652 ( .A1(n11480), .A2(n11418), .ZN(n11419) );
  AND2_X1 U14653 ( .A1(n11420), .A2(n11419), .ZN(n13688) );
  OAI21_X1 U14654 ( .B1(n14115), .B2(n11421), .A(n13688), .ZN(n11422) );
  NOR2_X1 U14655 ( .A1(n12786), .A2(n11422), .ZN(n11423) );
  NAND3_X1 U14656 ( .A1(n11425), .A2(n11424), .A3(n11423), .ZN(n11426) );
  AND2_X1 U14657 ( .A1(n14112), .A2(n10072), .ZN(n20050) );
  INV_X1 U14658 ( .A(n13344), .ZN(n11427) );
  NOR2_X1 U14659 ( .A1(n11427), .A2(n16105), .ZN(n13342) );
  XOR2_X1 U14660 ( .A(n11429), .B(n11428), .Z(n11430) );
  NAND2_X1 U14661 ( .A1(n13342), .A2(n11430), .ZN(n11431) );
  XOR2_X1 U14662 ( .A(n11430), .B(n13342), .Z(n13336) );
  NAND2_X1 U14663 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n13336), .ZN(
        n13335) );
  NAND2_X1 U14664 ( .A1(n11431), .A2(n13335), .ZN(n11434) );
  XOR2_X1 U14665 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n11434), .Z(
        n14795) );
  XOR2_X1 U14666 ( .A(n11433), .B(n11432), .Z(n14794) );
  NAND2_X1 U14667 ( .A1(n14795), .A2(n14794), .ZN(n14793) );
  NAND2_X1 U14668 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n11434), .ZN(
        n11435) );
  NAND2_X1 U14669 ( .A1(n14793), .A2(n11435), .ZN(n11436) );
  NAND2_X1 U14670 ( .A1(n11436), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11437) );
  XNOR2_X1 U14671 ( .A(n11440), .B(n11439), .ZN(n11442) );
  NAND2_X1 U14672 ( .A1(n11441), .A2(n11442), .ZN(n14049) );
  NAND2_X1 U14673 ( .A1(n14049), .A2(n14269), .ZN(n11445) );
  AND2_X2 U14674 ( .A1(n11445), .A2(n14050), .ZN(n14264) );
  NAND2_X1 U14675 ( .A1(n11446), .A2(n14270), .ZN(n14265) );
  NAND2_X1 U14676 ( .A1(n14264), .A2(n14265), .ZN(n11453) );
  INV_X1 U14677 ( .A(n11453), .ZN(n11448) );
  INV_X1 U14678 ( .A(n11447), .ZN(n11454) );
  NAND2_X1 U14679 ( .A1(n11448), .A2(n11447), .ZN(n11452) );
  INV_X1 U14680 ( .A(n11449), .ZN(n14267) );
  NAND2_X1 U14681 ( .A1(n14477), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n14478) );
  NAND2_X1 U14682 ( .A1(n11453), .A2(n14267), .ZN(n11455) );
  NAND2_X1 U14683 ( .A1(n11455), .A2(n11454), .ZN(n11456) );
  XNOR2_X1 U14684 ( .A(n11457), .B(n11254), .ZN(n14408) );
  OAI21_X1 U14686 ( .B1(n11459), .B2(n11254), .A(n16573), .ZN(n11460) );
  NAND2_X1 U14687 ( .A1(n11460), .A2(n11461), .ZN(n16538) );
  NOR2_X1 U14688 ( .A1(n16088), .A2(n16080), .ZN(n16071) );
  NAND2_X1 U14689 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n16071), .ZN(
        n16562) );
  NOR2_X1 U14690 ( .A1(n16570), .A2(n16562), .ZN(n16054) );
  AND2_X1 U14691 ( .A1(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n11462) );
  NOR2_X1 U14692 ( .A1(n11464), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n11465) );
  OR2_X1 U14693 ( .A1(n11463), .A2(n11465), .ZN(n15809) );
  AOI21_X1 U14694 ( .B1(n11467), .B2(n9863), .A(n10159), .ZN(n15812) );
  NAND2_X1 U14695 ( .A1(n14104), .A2(n20062), .ZN(n11471) );
  NAND2_X1 U14696 ( .A1(n11469), .A2(n11470), .ZN(n14106) );
  NAND2_X1 U14697 ( .A1(n11471), .A2(n14106), .ZN(n11472) );
  OR2_X1 U14698 ( .A1(n9871), .A2(n11473), .ZN(n11475) );
  INV_X1 U14699 ( .A(n15569), .ZN(n11474) );
  NAND2_X1 U14700 ( .A1(n11475), .A2(n11474), .ZN(n15745) );
  INV_X2 U14701 ( .A(n19345), .ZN(n19170) );
  NAND2_X1 U14702 ( .A1(n19170), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n15806) );
  NAND2_X1 U14703 ( .A1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n11513) );
  INV_X1 U14704 ( .A(n16004), .ZN(n11476) );
  NOR4_X1 U14705 ( .A1(n11476), .A2(n15990), .A3(n16491), .A4(n16034), .ZN(
        n15962) );
  NAND2_X1 U14706 ( .A1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n15962), .ZN(
        n11512) );
  NAND2_X1 U14707 ( .A1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16580) );
  NOR3_X1 U14708 ( .A1(n13867), .A2(n14270), .A3(n14269), .ZN(n11508) );
  INV_X1 U14709 ( .A(n11508), .ZN(n11501) );
  INV_X1 U14710 ( .A(n11477), .ZN(n11478) );
  NAND2_X1 U14711 ( .A1(n11484), .A2(n11478), .ZN(n11479) );
  NAND2_X1 U14712 ( .A1(n11505), .A2(n13379), .ZN(n19336) );
  INV_X1 U14713 ( .A(n19336), .ZN(n11500) );
  NOR2_X1 U14714 ( .A1(n16105), .A2(n19348), .ZN(n11498) );
  AND2_X1 U14715 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n11498), .ZN(
        n11504) );
  AND2_X1 U14716 ( .A1(n10983), .A2(n11481), .ZN(n11482) );
  NAND2_X1 U14717 ( .A1(n10982), .A2(n11482), .ZN(n11495) );
  NAND2_X1 U14718 ( .A1(n11483), .A2(n20062), .ZN(n14083) );
  NAND2_X1 U14719 ( .A1(n14083), .A2(n11484), .ZN(n11491) );
  INV_X1 U14720 ( .A(n13380), .ZN(n13331) );
  NAND2_X1 U14721 ( .A1(n11486), .A2(n10936), .ZN(n11488) );
  AOI22_X1 U14722 ( .A1(n13331), .A2(n11488), .B1(n10657), .B2(n11487), .ZN(
        n11489) );
  NAND2_X1 U14723 ( .A1(n11485), .A2(n11489), .ZN(n11490) );
  AOI21_X1 U14724 ( .B1(n11491), .B2(n19391), .A(n11490), .ZN(n11494) );
  AND2_X1 U14725 ( .A1(n13351), .A2(n11492), .ZN(n11493) );
  NAND2_X1 U14726 ( .A1(n10983), .A2(n11493), .ZN(n13384) );
  AND3_X1 U14727 ( .A1(n11495), .A2(n11494), .A3(n13384), .ZN(n14074) );
  INV_X1 U14728 ( .A(n11496), .ZN(n13677) );
  NAND2_X1 U14729 ( .A1(n14074), .A2(n13677), .ZN(n11497) );
  NAND2_X1 U14730 ( .A1(n11505), .A2(n11497), .ZN(n19333) );
  INV_X1 U14731 ( .A(n11498), .ZN(n19346) );
  NAND2_X1 U14732 ( .A1(n11499), .A2(n19346), .ZN(n11503) );
  OAI211_X1 U14733 ( .C1(n11500), .C2(n11504), .A(n16561), .B(n11503), .ZN(
        n14053) );
  NOR2_X1 U14734 ( .A1(n11501), .A2(n14053), .ZN(n14489) );
  NAND2_X1 U14735 ( .A1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n14489), .ZN(
        n14412) );
  INV_X1 U14736 ( .A(n16073), .ZN(n16052) );
  NOR2_X1 U14737 ( .A1(n11513), .A2(n15976), .ZN(n12483) );
  NAND2_X1 U14738 ( .A1(n12483), .A2(n11516), .ZN(n11502) );
  OAI211_X1 U14739 ( .C1(n19327), .C2(n15745), .A(n15806), .B(n11502), .ZN(
        n11518) );
  OR2_X1 U14740 ( .A1(n19336), .A2(n11503), .ZN(n19332) );
  OR2_X1 U14741 ( .A1(n19333), .A2(n11504), .ZN(n11507) );
  INV_X1 U14742 ( .A(n11505), .ZN(n11506) );
  NAND2_X1 U14743 ( .A1(n11506), .A2(n19345), .ZN(n19349) );
  AND2_X1 U14744 ( .A1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n11508), .ZN(
        n11509) );
  OR2_X1 U14745 ( .A1(n19353), .A2(n11509), .ZN(n11510) );
  NAND2_X1 U14746 ( .A1(n16561), .A2(n16580), .ZN(n11511) );
  NAND2_X1 U14747 ( .A1(n16047), .A2(n19353), .ZN(n15911) );
  NOR2_X1 U14748 ( .A1(n11513), .A2(n11512), .ZN(n11514) );
  NAND2_X1 U14749 ( .A1(n16047), .A2(n11514), .ZN(n11515) );
  NAND2_X1 U14750 ( .A1(n15911), .A2(n11515), .ZN(n12496) );
  NOR2_X1 U14751 ( .A1(n12496), .A2(n11516), .ZN(n11517) );
  AOI211_X1 U14752 ( .C1(n15812), .C2(n19341), .A(n11518), .B(n11517), .ZN(
        n11519) );
  INV_X1 U14753 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11522) );
  AND2_X2 U14754 ( .A1(n11522), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11527) );
  AOI22_X1 U14755 ( .A1(n11599), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n9826), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11525) );
  AND2_X2 U14756 ( .A1(n11528), .A2(n11527), .ZN(n12038) );
  AOI22_X1 U14757 ( .A1(n12038), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n12392), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11524) );
  AOI22_X1 U14758 ( .A1(n12043), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11612), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11523) );
  INV_X1 U14759 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11526) );
  AND2_X2 U14760 ( .A1(n11530), .A2(n11527), .ZN(n11684) );
  AOI22_X1 U14761 ( .A1(n11697), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n11622), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11533) );
  AND2_X2 U14762 ( .A1(n11530), .A2(n13958), .ZN(n11692) );
  AOI22_X1 U14763 ( .A1(n11692), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n11715), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11532) );
  AOI22_X1 U14764 ( .A1(n9849), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n11716), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11531) );
  INV_X1 U14765 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11535) );
  AND2_X2 U14766 ( .A1(n13945), .A2(n11537), .ZN(n12722) );
  AOI22_X1 U14767 ( .A1(n11766), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n12722), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11538) );
  AOI22_X1 U14768 ( .A1(n11692), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n11715), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11543) );
  AOI22_X1 U14769 ( .A1(n11697), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11622), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11542) );
  AOI22_X1 U14770 ( .A1(n11684), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n9821), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11541) );
  AOI22_X1 U14771 ( .A1(n9849), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n11716), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11540) );
  NAND4_X1 U14772 ( .A1(n11543), .A2(n11542), .A3(n11541), .A4(n11540), .ZN(
        n11549) );
  AOI22_X1 U14773 ( .A1(n11599), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n9825), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11547) );
  AOI22_X1 U14774 ( .A1(n12043), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11612), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11546) );
  AOI22_X1 U14775 ( .A1(n11766), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12722), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11544) );
  NAND4_X1 U14776 ( .A1(n11547), .A2(n11546), .A3(n11545), .A4(n11544), .ZN(
        n11548) );
  AOI22_X1 U14777 ( .A1(n12043), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11715), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11553) );
  AOI22_X1 U14778 ( .A1(n9825), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(n9821), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11552) );
  AOI22_X1 U14779 ( .A1(n12724), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n11716), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11551) );
  AOI22_X1 U14780 ( .A1(n11684), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11612), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11550) );
  AOI22_X1 U14781 ( .A1(n12392), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11599), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11555) );
  NAND2_X1 U14782 ( .A1(n11555), .A2(n11554), .ZN(n11559) );
  AOI22_X1 U14783 ( .A1(n12038), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11622), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11557) );
  AOI22_X1 U14784 ( .A1(n11697), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11692), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11556) );
  NAND2_X1 U14785 ( .A1(n11557), .A2(n11556), .ZN(n11558) );
  NAND2_X2 U14786 ( .A1(n11561), .A2(n11560), .ZN(n12766) );
  AOI22_X1 U14787 ( .A1(n11697), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11692), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11565) );
  AOI22_X1 U14788 ( .A1(n11684), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11622), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11564) );
  AOI22_X1 U14789 ( .A1(n9848), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11716), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11562) );
  AOI22_X1 U14790 ( .A1(n12392), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11599), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11569) );
  AOI22_X1 U14791 ( .A1(n12038), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11715), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11568) );
  AOI22_X1 U14792 ( .A1(n11612), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n9824), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11567) );
  AOI22_X1 U14793 ( .A1(n12043), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11612), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11576) );
  AOI22_X1 U14794 ( .A1(n11599), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n9826), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11575) );
  AOI22_X1 U14795 ( .A1(n11766), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12722), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11574) );
  NAND4_X1 U14796 ( .A1(n11577), .A2(n11576), .A3(n11575), .A4(n11574), .ZN(
        n11583) );
  AOI22_X1 U14797 ( .A1(n11697), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11622), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11580) );
  AOI22_X1 U14798 ( .A1(n11684), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12723), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11579) );
  AOI22_X1 U14799 ( .A1(n12724), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11716), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11578) );
  NAND4_X1 U14800 ( .A1(n11581), .A2(n11580), .A3(n11579), .A4(n11578), .ZN(
        n11582) );
  INV_X1 U14801 ( .A(n12766), .ZN(n11665) );
  AND2_X2 U14802 ( .A1(n11665), .A2(n11816), .ZN(n11654) );
  INV_X1 U14803 ( .A(n11584), .ZN(n11585) );
  AOI22_X1 U14804 ( .A1(n9851), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(n9826), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11589) );
  AOI22_X1 U14805 ( .A1(n9838), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11612), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11588) );
  AOI22_X1 U14806 ( .A1(n12038), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12392), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11587) );
  BUF_X4 U14807 ( .A(n12722), .Z(n12702) );
  AOI22_X1 U14808 ( .A1(n11766), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12702), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11586) );
  NAND4_X1 U14809 ( .A1(n11589), .A2(n11588), .A3(n11587), .A4(n11586), .ZN(
        n11595) );
  AOI22_X1 U14810 ( .A1(n11692), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n11715), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11593) );
  AOI22_X1 U14811 ( .A1(n11697), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11622), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11592) );
  AOI22_X1 U14812 ( .A1(n11684), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12723), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11591) );
  AOI22_X1 U14813 ( .A1(n12724), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n11716), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11590) );
  NAND4_X1 U14814 ( .A1(n11593), .A2(n11592), .A3(n11591), .A4(n11590), .ZN(
        n11594) );
  NAND2_X1 U14815 ( .A1(n11657), .A2(n20331), .ZN(n11596) );
  NAND2_X1 U14816 ( .A1(n12392), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n11603) );
  NAND2_X1 U14817 ( .A1(n12038), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n11602) );
  NAND2_X1 U14818 ( .A1(n9850), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n11601) );
  NAND2_X1 U14819 ( .A1(n9826), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n11600) );
  NAND2_X1 U14820 ( .A1(n11697), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n11607) );
  NAND2_X1 U14821 ( .A1(n11684), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n11606) );
  NAND2_X1 U14822 ( .A1(n11622), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n11605) );
  NAND2_X1 U14823 ( .A1(n11692), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n11611) );
  NAND2_X1 U14824 ( .A1(n9849), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n11610) );
  NAND2_X1 U14825 ( .A1(n11715), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n11609) );
  NAND2_X1 U14826 ( .A1(n11716), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n11608) );
  NAND2_X1 U14827 ( .A1(n11612), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n11616) );
  NAND2_X1 U14828 ( .A1(n9838), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n11615) );
  NAND2_X1 U14829 ( .A1(n11766), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n11614) );
  NAND2_X1 U14830 ( .A1(n12702), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n11613) );
  NAND4_X4 U14831 ( .A1(n11620), .A2(n11619), .A3(n11618), .A4(n11617), .ZN(
        n11644) );
  NOR2_X1 U14832 ( .A1(n11598), .A2(n11644), .ZN(n11621) );
  NAND2_X2 U14833 ( .A1(n11649), .A2(n11621), .ZN(n12757) );
  AOI22_X1 U14834 ( .A1(n11684), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n11622), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11626) );
  AOI22_X1 U14835 ( .A1(n11692), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n12723), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11625) );
  AOI22_X1 U14836 ( .A1(n12392), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n11612), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11624) );
  AOI22_X1 U14837 ( .A1(n9848), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n11716), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11623) );
  NAND4_X1 U14838 ( .A1(n11626), .A2(n11625), .A3(n11624), .A4(n11623), .ZN(
        n11632) );
  AOI22_X1 U14839 ( .A1(n12038), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n9851), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11630) );
  AOI22_X1 U14840 ( .A1(n11697), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n11715), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11629) );
  AOI22_X1 U14841 ( .A1(n12043), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n9826), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11628) );
  AOI22_X1 U14842 ( .A1(n11766), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12722), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11627) );
  NAND4_X1 U14843 ( .A1(n11630), .A2(n11629), .A3(n11628), .A4(n11627), .ZN(
        n11631) );
  NAND2_X1 U14844 ( .A1(n11634), .A2(n11633), .ZN(n13473) );
  NAND2_X1 U14845 ( .A1(n11654), .A2(n11635), .ZN(n11637) );
  NAND2_X1 U14846 ( .A1(n11641), .A2(n12766), .ZN(n11636) );
  NAND2_X1 U14847 ( .A1(n11637), .A2(n11650), .ZN(n13516) );
  INV_X1 U14848 ( .A(n13516), .ZN(n11638) );
  NAND2_X1 U14849 ( .A1(n11638), .A2(n11835), .ZN(n11919) );
  NOR2_X2 U14850 ( .A1(n11919), .A2(n11639), .ZN(n13461) );
  NAND2_X1 U14851 ( .A1(n16201), .A2(n11644), .ZN(n12857) );
  INV_X2 U14852 ( .A(n12857), .ZN(n13548) );
  XNOR2_X1 U14853 ( .A(n20928), .B(P1_STATE_REG_1__SCAN_IN), .ZN(n12941) );
  NOR2_X2 U14854 ( .A1(n16201), .A2(n11644), .ZN(n12763) );
  NAND2_X1 U14855 ( .A1(n13943), .A2(n11641), .ZN(n13543) );
  INV_X1 U14856 ( .A(n13543), .ZN(n11642) );
  INV_X1 U14857 ( .A(n20331), .ZN(n11645) );
  NAND2_X1 U14858 ( .A1(n11647), .A2(n11646), .ZN(n13511) );
  INV_X1 U14859 ( .A(n13943), .ZN(n11648) );
  NAND2_X1 U14860 ( .A1(n13775), .A2(n16201), .ZN(n13839) );
  INV_X1 U14861 ( .A(n11649), .ZN(n11664) );
  NAND2_X1 U14862 ( .A1(n11664), .A2(n13775), .ZN(n11659) );
  INV_X1 U14863 ( .A(n11650), .ZN(n11653) );
  NAND2_X1 U14864 ( .A1(n11669), .A2(n11670), .ZN(n11658) );
  NAND2_X1 U14865 ( .A1(n11670), .A2(n11644), .ZN(n11655) );
  NAND2_X1 U14866 ( .A1(n11655), .A2(n12755), .ZN(n11656) );
  NAND2_X1 U14867 ( .A1(n11658), .A2(n13521), .ZN(n11675) );
  NAND2_X1 U14868 ( .A1(n20846), .A2(n20767), .ZN(n20732) );
  AND2_X1 U14869 ( .A1(n20910), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n11736) );
  AOI21_X1 U14870 ( .B1(n12414), .B2(n20656), .A(n11736), .ZN(n11660) );
  NAND2_X1 U14871 ( .A1(n11661), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11735) );
  INV_X1 U14872 ( .A(n20910), .ZN(n16207) );
  INV_X1 U14873 ( .A(n12414), .ZN(n11745) );
  MUX2_X1 U14874 ( .A(n16207), .B(n11745), .S(n20767), .Z(n11663) );
  OAI21_X2 U14875 ( .B1(n11742), .B2(n13523), .A(n11663), .ZN(n11710) );
  NAND2_X1 U14876 ( .A1(n11664), .A2(n12763), .ZN(n13519) );
  NAND2_X1 U14877 ( .A1(n13943), .A2(n11665), .ZN(n11666) );
  NAND3_X1 U14878 ( .A1(n13839), .A2(P1_STATE2_REG_0__SCAN_IN), .A3(n20080), 
        .ZN(n11667) );
  NOR2_X1 U14879 ( .A1(n11668), .A2(n11667), .ZN(n11674) );
  INV_X1 U14880 ( .A(n11669), .ZN(n11672) );
  NAND2_X1 U14881 ( .A1(n11670), .A2(n20331), .ZN(n11671) );
  AOI22_X1 U14882 ( .A1(n21001), .A2(n11672), .B1(n13420), .B2(n11671), .ZN(
        n11673) );
  OAI211_X1 U14883 ( .C1(n11675), .C2(n11633), .A(n11674), .B(n11673), .ZN(
        n11676) );
  INV_X1 U14884 ( .A(n11676), .ZN(n11677) );
  AOI22_X1 U14885 ( .A1(n9838), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n9820), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11683) );
  AOI22_X1 U14886 ( .A1(n12038), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n11622), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11682) );
  AOI22_X1 U14887 ( .A1(n12729), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n9821), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11681) );
  AOI22_X1 U14888 ( .A1(n12250), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n12702), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11680) );
  NAND4_X1 U14889 ( .A1(n11683), .A2(n11682), .A3(n11681), .A4(n11680), .ZN(
        n11690) );
  AOI22_X1 U14890 ( .A1(n12732), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n9850), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11688) );
  AOI22_X1 U14891 ( .A1(n12374), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12731), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11687) );
  AOI22_X1 U14892 ( .A1(n12286), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n9825), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11686) );
  AOI22_X1 U14893 ( .A1(n12724), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12185), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11685) );
  NAND4_X1 U14894 ( .A1(n11688), .A2(n11687), .A3(n11686), .A4(n11685), .ZN(
        n11689) );
  NAND2_X1 U14895 ( .A1(n9933), .A2(n11834), .ZN(n11691) );
  AOI22_X1 U14896 ( .A1(n12038), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12392), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11696) );
  AOI22_X1 U14897 ( .A1(n12286), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12732), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11695) );
  AOI22_X1 U14898 ( .A1(n9838), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11612), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11694) );
  AOI22_X1 U14899 ( .A1(n11766), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n12702), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11693) );
  NAND4_X1 U14900 ( .A1(n11696), .A2(n11695), .A3(n11694), .A4(n11693), .ZN(
        n11703) );
  AOI22_X1 U14901 ( .A1(n12729), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n9852), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11700) );
  AOI22_X1 U14902 ( .A1(n12731), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n11622), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11699) );
  AOI22_X1 U14903 ( .A1(n12724), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12185), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11698) );
  NAND4_X1 U14904 ( .A1(n11701), .A2(n11700), .A3(n11699), .A4(n11698), .ZN(
        n11702) );
  INV_X1 U14905 ( .A(n11896), .ZN(n11882) );
  NAND2_X1 U14906 ( .A1(n13775), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11758) );
  INV_X1 U14907 ( .A(n11758), .ZN(n11704) );
  AOI22_X1 U14908 ( .A1(n9933), .A2(n11882), .B1(n11704), .B2(n11834), .ZN(
        n11707) );
  NAND2_X1 U14909 ( .A1(n11968), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11706) );
  XNOR2_X1 U14910 ( .A(n11710), .B(n11709), .ZN(n11993) );
  NAND2_X1 U14911 ( .A1(n11993), .A2(n20310), .ZN(n11725) );
  AOI22_X1 U14912 ( .A1(n9838), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11612), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11714) );
  AOI22_X1 U14913 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n12392), .B1(
        n11599), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11713) );
  AOI22_X1 U14914 ( .A1(n11766), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n12702), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11712) );
  AOI22_X1 U14915 ( .A1(n12038), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12356), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11711) );
  NAND4_X1 U14916 ( .A1(n11714), .A2(n11713), .A3(n11712), .A4(n11711), .ZN(
        n11722) );
  AOI22_X1 U14917 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n12729), .B1(
        n12732), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11720) );
  AOI22_X1 U14918 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n12731), .B1(
        n9825), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11719) );
  AOI22_X1 U14920 ( .A1(n9849), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12185), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11717) );
  NAND4_X1 U14921 ( .A1(n11720), .A2(n11719), .A3(n11718), .A4(n11717), .ZN(
        n11721) );
  XNOR2_X1 U14922 ( .A(n11727), .B(n11896), .ZN(n11723) );
  NAND2_X1 U14923 ( .A1(n11723), .A2(n9933), .ZN(n11724) );
  INV_X1 U14924 ( .A(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11730) );
  NAND2_X1 U14925 ( .A1(n11679), .A2(n11896), .ZN(n11726) );
  OAI211_X1 U14926 ( .C1(n11727), .C2(n11644), .A(n11726), .B(
        P1_STATE2_REG_0__SCAN_IN), .ZN(n11728) );
  INV_X1 U14927 ( .A(n11728), .ZN(n11729) );
  NAND2_X1 U14928 ( .A1(n11984), .A2(n11985), .ZN(n11734) );
  INV_X1 U14929 ( .A(n11731), .ZN(n11732) );
  INV_X1 U14930 ( .A(n11735), .ZN(n11739) );
  INV_X1 U14931 ( .A(n11736), .ZN(n11737) );
  NAND2_X1 U14932 ( .A1(n11737), .A2(n13554), .ZN(n11738) );
  NAND2_X1 U14933 ( .A1(n11739), .A2(n11738), .ZN(n11740) );
  XNOR2_X1 U14934 ( .A(n20696), .B(n20598), .ZN(n20318) );
  OR2_X1 U14935 ( .A1(n11742), .A2(n13561), .ZN(n11744) );
  NAND2_X1 U14936 ( .A1(n20910), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n11743) );
  AOI22_X1 U14937 ( .A1(n12116), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12392), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11751) );
  AOI22_X1 U14938 ( .A1(n9838), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11612), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11750) );
  AOI22_X1 U14939 ( .A1(n9851), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(n9826), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11749) );
  AOI22_X1 U14940 ( .A1(n12250), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n12702), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11748) );
  NAND4_X1 U14941 ( .A1(n11751), .A2(n11750), .A3(n11749), .A4(n11748), .ZN(
        n11757) );
  AOI22_X1 U14942 ( .A1(n12732), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12731), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11755) );
  AOI22_X1 U14943 ( .A1(n12729), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12356), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11754) );
  AOI22_X1 U14944 ( .A1(n9848), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12185), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11752) );
  NAND4_X1 U14945 ( .A1(n11755), .A2(n11754), .A3(n11753), .A4(n11752), .ZN(
        n11756) );
  INV_X1 U14946 ( .A(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11759) );
  OAI22_X1 U14947 ( .A1(n11959), .A2(n11759), .B1(n11758), .B2(n11846), .ZN(
        n11760) );
  OAI21_X1 U14948 ( .B1(n20696), .B2(n20598), .A(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n11762) );
  INV_X1 U14949 ( .A(n20696), .ZN(n20843) );
  NAND2_X1 U14950 ( .A1(n20387), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n20520) );
  INV_X1 U14951 ( .A(n20520), .ZN(n11761) );
  NAND2_X1 U14952 ( .A1(n20843), .A2(n11761), .ZN(n20562) );
  NAND2_X1 U14953 ( .A1(n11762), .A2(n20562), .ZN(n20599) );
  AOI22_X1 U14954 ( .A1(n12414), .A2(n20599), .B1(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n20910), .ZN(n11763) );
  INV_X1 U14955 ( .A(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n21089) );
  AOI22_X1 U14956 ( .A1(n12116), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12392), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11770) );
  AOI22_X1 U14957 ( .A1(n9838), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11612), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11769) );
  AOI22_X1 U14958 ( .A1(n9850), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(n9825), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11768) );
  AOI22_X1 U14959 ( .A1(n12250), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12702), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11767) );
  NAND4_X1 U14960 ( .A1(n11770), .A2(n11769), .A3(n11768), .A4(n11767), .ZN(
        n11776) );
  AOI22_X1 U14961 ( .A1(n12732), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12731), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11774) );
  AOI22_X1 U14962 ( .A1(n12729), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12356), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11773) );
  AOI22_X1 U14963 ( .A1(n9849), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12185), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11771) );
  NAND4_X1 U14964 ( .A1(n11774), .A2(n11773), .A3(n11772), .A4(n11771), .ZN(
        n11775) );
  AOI22_X1 U14965 ( .A1(n11968), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n11939), .B2(n11865), .ZN(n11777) );
  NAND2_X2 U14966 ( .A1(n11779), .A2(n13972), .ZN(n11855) );
  INV_X1 U14967 ( .A(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11791) );
  AOI22_X1 U14968 ( .A1(n9838), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12374), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11783) );
  AOI22_X1 U14969 ( .A1(n9820), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(n9851), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11782) );
  AOI22_X1 U14970 ( .A1(n12250), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n12702), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11781) );
  AOI22_X1 U14971 ( .A1(n12116), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n11622), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11780) );
  NAND4_X1 U14972 ( .A1(n11783), .A2(n11782), .A3(n11781), .A4(n11780), .ZN(
        n11789) );
  AOI22_X1 U14973 ( .A1(n12286), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n12732), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11787) );
  AOI22_X1 U14974 ( .A1(n12731), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n9826), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11786) );
  AOI22_X1 U14975 ( .A1(n9849), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n12185), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11784) );
  NAND4_X1 U14976 ( .A1(n11787), .A2(n11786), .A3(n11785), .A4(n11784), .ZN(
        n11788) );
  NAND2_X1 U14977 ( .A1(n11939), .A2(n11864), .ZN(n11790) );
  OAI21_X1 U14978 ( .B1(n11959), .B2(n11791), .A(n11790), .ZN(n11854) );
  INV_X1 U14979 ( .A(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11803) );
  AOI22_X1 U14980 ( .A1(n12116), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n9817), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11795) );
  AOI22_X1 U14981 ( .A1(n9838), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12374), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11794) );
  AOI22_X1 U14982 ( .A1(n9850), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(n9825), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11793) );
  AOI22_X1 U14983 ( .A1(n12250), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12702), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11792) );
  NAND4_X1 U14984 ( .A1(n11795), .A2(n11794), .A3(n11793), .A4(n11792), .ZN(
        n11801) );
  INV_X1 U14985 ( .A(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n21142) );
  AOI22_X1 U14986 ( .A1(n12732), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12731), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11799) );
  AOI22_X1 U14987 ( .A1(n12729), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12356), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11798) );
  AOI22_X1 U14988 ( .A1(n12724), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12185), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11796) );
  NAND4_X1 U14989 ( .A1(n11799), .A2(n11798), .A3(n11797), .A4(n11796), .ZN(
        n11800) );
  NAND2_X1 U14990 ( .A1(n11939), .A2(n11887), .ZN(n11802) );
  OAI21_X1 U14991 ( .B1(n11959), .B2(n11803), .A(n11802), .ZN(n11862) );
  INV_X1 U14992 ( .A(n11874), .ZN(n11815) );
  AOI22_X1 U14993 ( .A1(n9817), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12286), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11807) );
  AOI22_X1 U14994 ( .A1(n12116), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12732), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11806) );
  AOI22_X1 U14995 ( .A1(n9848), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12185), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11804) );
  NAND4_X1 U14996 ( .A1(n11807), .A2(n11806), .A3(n11805), .A4(n11804), .ZN(
        n11813) );
  AOI22_X1 U14997 ( .A1(n12729), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12731), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11811) );
  AOI22_X1 U14998 ( .A1(n12374), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n9826), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11810) );
  AOI22_X1 U14999 ( .A1(n9851), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n12356), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11809) );
  AOI22_X1 U15000 ( .A1(n12250), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n12702), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11808) );
  NAND4_X1 U15001 ( .A1(n11811), .A2(n11810), .A3(n11809), .A4(n11808), .ZN(
        n11812) );
  AOI22_X1 U15002 ( .A1(n11968), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n11939), .B2(n11888), .ZN(n11873) );
  INV_X1 U15003 ( .A(n11873), .ZN(n11814) );
  AND2_X1 U15004 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15347) );
  NAND2_X1 U15005 ( .A1(n15347), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15344) );
  INV_X1 U15006 ( .A(n15344), .ZN(n11912) );
  NAND2_X1 U15007 ( .A1(n11820), .A2(n11819), .ZN(n11821) );
  INV_X1 U15008 ( .A(n13971), .ZN(n11822) );
  NAND2_X1 U15009 ( .A1(n11822), .A2(n11886), .ZN(n11826) );
  NAND2_X1 U15010 ( .A1(n11834), .A2(n11833), .ZN(n11847) );
  XNOR2_X1 U15011 ( .A(n11847), .B(n11846), .ZN(n11824) );
  NAND2_X1 U15012 ( .A1(n13775), .A2(n20331), .ZN(n11828) );
  INV_X1 U15013 ( .A(n11828), .ZN(n11823) );
  AOI21_X1 U15014 ( .B1(n11824), .B2(n21001), .A(n11823), .ZN(n11825) );
  NAND2_X1 U15015 ( .A1(n11826), .A2(n11825), .ZN(n13734) );
  OAI21_X1 U15016 ( .B1(n12755), .B2(n11833), .A(n11828), .ZN(n11829) );
  INV_X1 U15017 ( .A(n11829), .ZN(n11830) );
  OAI21_X2 U15018 ( .B1(n11991), .B2(n11929), .A(n11830), .ZN(n13533) );
  INV_X1 U15019 ( .A(n11831), .ZN(n11832) );
  NAND2_X1 U15020 ( .A1(n11832), .A2(n16201), .ZN(n11839) );
  XNOR2_X1 U15021 ( .A(n11834), .B(n11833), .ZN(n11836) );
  OAI211_X1 U15022 ( .C1(n11836), .C2(n12755), .A(n11835), .B(n11816), .ZN(
        n11837) );
  INV_X1 U15023 ( .A(n11837), .ZN(n11838) );
  NAND2_X1 U15024 ( .A1(n11839), .A2(n11838), .ZN(n11841) );
  INV_X1 U15025 ( .A(n11840), .ZN(n13534) );
  NAND2_X1 U15026 ( .A1(n13534), .A2(n11841), .ZN(n11842) );
  INV_X1 U15027 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n14501) );
  NAND2_X1 U15028 ( .A1(n11843), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11844) );
  INV_X1 U15029 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n20273) );
  INV_X1 U15030 ( .A(n13972), .ZN(n13974) );
  NAND2_X2 U15031 ( .A1(n11855), .A2(n11845), .ZN(n20594) );
  OR2_X1 U15032 ( .A1(n20594), .A2(n11929), .ZN(n11851) );
  NAND2_X1 U15033 ( .A1(n11847), .A2(n11846), .ZN(n11867) );
  INV_X1 U15034 ( .A(n11865), .ZN(n11848) );
  XNOR2_X1 U15035 ( .A(n11867), .B(n11848), .ZN(n11849) );
  NAND2_X1 U15036 ( .A1(n11849), .A2(n21001), .ZN(n11850) );
  NAND2_X1 U15037 ( .A1(n11851), .A2(n11850), .ZN(n13849) );
  NAND2_X1 U15038 ( .A1(n11852), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11853) );
  XNOR2_X1 U15039 ( .A(n11855), .B(n11854), .ZN(n12017) );
  NAND2_X1 U15040 ( .A1(n12017), .A2(n11886), .ZN(n11859) );
  NAND2_X1 U15041 ( .A1(n11867), .A2(n11865), .ZN(n11856) );
  XNOR2_X1 U15042 ( .A(n11856), .B(n11864), .ZN(n11857) );
  NAND2_X1 U15043 ( .A1(n11857), .A2(n21001), .ZN(n11858) );
  NAND2_X1 U15044 ( .A1(n11859), .A2(n11858), .ZN(n11860) );
  XNOR2_X1 U15045 ( .A(n11860), .B(n20267), .ZN(n20244) );
  NAND2_X1 U15046 ( .A1(n11860), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11861) );
  XNOR2_X1 U15047 ( .A(n11863), .B(n11862), .ZN(n12018) );
  NAND2_X1 U15048 ( .A1(n12018), .A2(n11886), .ZN(n11870) );
  AND2_X1 U15049 ( .A1(n11865), .A2(n11864), .ZN(n11866) );
  NAND2_X1 U15050 ( .A1(n11867), .A2(n11866), .ZN(n11875) );
  XNOR2_X1 U15051 ( .A(n11875), .B(n11887), .ZN(n11868) );
  NAND2_X1 U15052 ( .A1(n11868), .A2(n21001), .ZN(n11869) );
  NAND2_X1 U15053 ( .A1(n11870), .A2(n11869), .ZN(n11871) );
  INV_X1 U15054 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n16430) );
  NAND2_X1 U15055 ( .A1(n11871), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11872) );
  NAND2_X1 U15056 ( .A1(n11874), .A2(n11873), .ZN(n12031) );
  INV_X1 U15057 ( .A(n11875), .ZN(n11890) );
  NAND2_X1 U15058 ( .A1(n11890), .A2(n11887), .ZN(n11876) );
  XNOR2_X1 U15059 ( .A(n11876), .B(n11888), .ZN(n11877) );
  NAND2_X1 U15060 ( .A1(n11877), .A2(n21001), .ZN(n11878) );
  NAND2_X1 U15061 ( .A1(n11879), .A2(n11878), .ZN(n16335) );
  OR2_X1 U15062 ( .A1(n16335), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11880) );
  NAND2_X1 U15063 ( .A1(n16335), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11881) );
  INV_X1 U15064 ( .A(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11883) );
  INV_X1 U15065 ( .A(n11939), .ZN(n11946) );
  OAI22_X1 U15066 ( .A1(n11959), .A2(n11883), .B1(n11946), .B2(n11882), .ZN(
        n11884) );
  NAND2_X1 U15067 ( .A1(n12037), .A2(n11886), .ZN(n11893) );
  AND2_X1 U15068 ( .A1(n11888), .A2(n11887), .ZN(n11889) );
  NAND2_X1 U15069 ( .A1(n11890), .A2(n11889), .ZN(n11895) );
  XNOR2_X1 U15070 ( .A(n11895), .B(n11896), .ZN(n11891) );
  NAND2_X1 U15071 ( .A1(n11891), .A2(n21001), .ZN(n11892) );
  NAND2_X1 U15072 ( .A1(n11893), .A2(n11892), .ZN(n11894) );
  OR2_X1 U15073 ( .A1(n11894), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16331) );
  NAND2_X1 U15074 ( .A1(n11894), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16330) );
  INV_X1 U15075 ( .A(n11895), .ZN(n11897) );
  NAND3_X1 U15076 ( .A1(n11897), .A2(n21001), .A3(n11896), .ZN(n11898) );
  NAND2_X1 U15077 ( .A1(n9844), .A2(n11898), .ZN(n14470) );
  NAND2_X1 U15078 ( .A1(n14470), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11900) );
  NAND2_X1 U15079 ( .A1(n9845), .A2(n16390), .ZN(n11901) );
  INV_X1 U15080 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15425) );
  OR2_X1 U15081 ( .A1(n11907), .A2(n15425), .ZN(n15235) );
  NAND2_X1 U15082 ( .A1(n9845), .A2(n15425), .ZN(n11902) );
  NAND2_X1 U15083 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n11903) );
  AND2_X1 U15084 ( .A1(n9845), .A2(n11903), .ZN(n15243) );
  AND2_X1 U15085 ( .A1(n9844), .A2(n15453), .ZN(n15246) );
  INV_X1 U15086 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n12892) );
  AND2_X1 U15087 ( .A1(n9844), .A2(n12892), .ZN(n15222) );
  NOR2_X1 U15088 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n11904) );
  OR2_X1 U15089 ( .A1(n9845), .A2(n11904), .ZN(n16312) );
  INV_X1 U15090 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n11905) );
  OR2_X1 U15091 ( .A1(n9844), .A2(n11905), .ZN(n16311) );
  NAND2_X1 U15092 ( .A1(n9844), .A2(n11905), .ZN(n16310) );
  INV_X1 U15093 ( .A(n16300), .ZN(n11906) );
  INV_X1 U15094 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n16359) );
  OR2_X1 U15095 ( .A1(n9844), .A2(n15453), .ZN(n15244) );
  NOR2_X1 U15096 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n11908) );
  OR2_X1 U15097 ( .A1(n9845), .A2(n11908), .ZN(n15242) );
  XNOR2_X1 U15098 ( .A(n9844), .B(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15214) );
  AND2_X1 U15099 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15287) );
  AND2_X1 U15100 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15289) );
  NAND2_X1 U15101 ( .A1(n15287), .A2(n15289), .ZN(n15276) );
  INV_X1 U15102 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15392) );
  OAI21_X2 U15103 ( .B1(n15180), .B2(n15276), .A(n11909), .ZN(n13001) );
  INV_X1 U15104 ( .A(n15213), .ZN(n15191) );
  INV_X1 U15105 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n15433) );
  INV_X1 U15106 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n21220) );
  INV_X1 U15107 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n15402) );
  INV_X1 U15108 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15410) );
  AND4_X1 U15109 ( .A1(n15433), .A2(n21220), .A3(n15402), .A4(n15410), .ZN(
        n11910) );
  INV_X1 U15110 ( .A(n11913), .ZN(n11915) );
  INV_X1 U15111 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15355) );
  INV_X1 U15112 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15362) );
  NAND2_X1 U15113 ( .A1(n15355), .A2(n15362), .ZN(n13000) );
  NOR4_X1 U15114 ( .A1(n13000), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A4(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n11914) );
  NAND2_X1 U15115 ( .A1(n11913), .A2(n11914), .ZN(n11917) );
  NAND3_X1 U15116 ( .A1(n11915), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n11916) );
  MUX2_X1 U15117 ( .A(n11917), .B(n11916), .S(n9844), .Z(n11918) );
  INV_X1 U15118 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15327) );
  AND2_X1 U15119 ( .A1(n13521), .A2(n13775), .ZN(n11920) );
  XNOR2_X1 U15120 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n11943) );
  NAND2_X1 U15121 ( .A1(n11944), .A2(n11943), .ZN(n11922) );
  NAND2_X1 U15122 ( .A1(n20846), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11921) );
  NAND2_X1 U15123 ( .A1(n11922), .A2(n11921), .ZN(n11933) );
  XNOR2_X1 U15124 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n11932) );
  NAND2_X1 U15125 ( .A1(n11933), .A2(n11932), .ZN(n11924) );
  NAND2_X1 U15126 ( .A1(n20598), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11923) );
  NAND2_X1 U15127 ( .A1(n11924), .A2(n11923), .ZN(n11931) );
  MUX2_X1 U15128 ( .A(n20387), .B(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .S(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n11930) );
  NAND2_X1 U15129 ( .A1(n11931), .A2(n11930), .ZN(n11926) );
  NAND2_X1 U15130 ( .A1(n20387), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11925) );
  NAND2_X1 U15131 ( .A1(n11926), .A2(n11925), .ZN(n11964) );
  NAND2_X1 U15132 ( .A1(n11962), .A2(n12758), .ZN(n11975) );
  XNOR2_X1 U15133 ( .A(n11931), .B(n11930), .ZN(n12761) );
  NAND2_X1 U15134 ( .A1(n11633), .A2(n11816), .ZN(n11947) );
  NAND2_X1 U15135 ( .A1(n16196), .A2(n11947), .ZN(n11937) );
  INV_X1 U15136 ( .A(n11937), .ZN(n11958) );
  XNOR2_X1 U15137 ( .A(n11933), .B(n11932), .ZN(n12760) );
  INV_X1 U15138 ( .A(n12760), .ZN(n11934) );
  AND2_X1 U15139 ( .A1(n11939), .A2(n11934), .ZN(n11935) );
  INV_X1 U15140 ( .A(n11935), .ZN(n11957) );
  AOI211_X1 U15141 ( .C1(n11968), .C2(n12760), .A(n11935), .B(n11937), .ZN(
        n11956) );
  INV_X1 U15142 ( .A(n11598), .ZN(n13790) );
  INV_X1 U15143 ( .A(n11944), .ZN(n11936) );
  OAI21_X1 U15144 ( .B1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n20767), .A(
        n11936), .ZN(n11938) );
  AOI211_X1 U15145 ( .C1(n13790), .C2(n11644), .A(n11937), .B(n11938), .ZN(
        n11942) );
  INV_X1 U15146 ( .A(n11938), .ZN(n11940) );
  AOI21_X1 U15147 ( .B1(n11940), .B2(n11939), .A(n11962), .ZN(n11941) );
  NOR2_X1 U15148 ( .A1(n11942), .A2(n11941), .ZN(n11954) );
  XNOR2_X1 U15149 ( .A(n11944), .B(n11943), .ZN(n12759) );
  NAND2_X1 U15150 ( .A1(n11641), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11945) );
  NAND2_X1 U15151 ( .A1(n11946), .A2(n11945), .ZN(n11948) );
  AOI22_X1 U15152 ( .A1(n11968), .A2(n12759), .B1(n11947), .B2(n11948), .ZN(
        n11951) );
  INV_X1 U15153 ( .A(n11951), .ZN(n11953) );
  INV_X1 U15154 ( .A(n11948), .ZN(n11949) );
  NAND2_X1 U15155 ( .A1(n11949), .A2(n16201), .ZN(n11966) );
  INV_X1 U15156 ( .A(n11954), .ZN(n11950) );
  AOI22_X1 U15157 ( .A1(n12759), .A2(n11966), .B1(n11951), .B2(n11950), .ZN(
        n11952) );
  AOI21_X1 U15158 ( .B1(n11954), .B2(n11953), .A(n11952), .ZN(n11955) );
  OAI22_X1 U15159 ( .A1(n11958), .A2(n11957), .B1(n11956), .B2(n11955), .ZN(
        n11961) );
  NAND2_X1 U15160 ( .A1(n11959), .A2(n12761), .ZN(n11960) );
  AOI22_X1 U15161 ( .A1(n11962), .A2(n12761), .B1(n11961), .B2(n11960), .ZN(
        n11971) );
  INV_X1 U15162 ( .A(n12762), .ZN(n11965) );
  NOR2_X1 U15163 ( .A1(n11968), .A2(n11965), .ZN(n11970) );
  INV_X1 U15164 ( .A(n11966), .ZN(n11967) );
  NAND3_X1 U15165 ( .A1(n11968), .A2(n11967), .A3(n12762), .ZN(n11969) );
  OAI21_X1 U15166 ( .B1(n11971), .B2(n11970), .A(n11969), .ZN(n11972) );
  AOI21_X1 U15167 ( .B1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n20310), .A(
        n11972), .ZN(n11973) );
  INV_X1 U15168 ( .A(n11973), .ZN(n11974) );
  NOR2_X1 U15169 ( .A1(n11598), .A2(n20086), .ZN(n11978) );
  NAND2_X1 U15170 ( .A1(n10042), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12013) );
  XNOR2_X1 U15171 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13936) );
  AOI21_X1 U15172 ( .B1(n12847), .B2(n13936), .A(n12747), .ZN(n11981) );
  NAND2_X1 U15173 ( .A1(n12748), .A2(P1_EAX_REG_2__SCAN_IN), .ZN(n11980) );
  OAI211_X1 U15174 ( .C1(n12013), .C2(n13561), .A(n11981), .B(n11980), .ZN(
        n11982) );
  INV_X1 U15175 ( .A(n11982), .ZN(n11983) );
  NAND2_X1 U15176 ( .A1(n12747), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11999) );
  NAND2_X1 U15177 ( .A1(n13973), .A2(n12154), .ZN(n11990) );
  AOI22_X1 U15178 ( .A1(n12748), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n20999), .ZN(n11988) );
  INV_X1 U15179 ( .A(n12013), .ZN(n11986) );
  NAND2_X1 U15180 ( .A1(n11986), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11987) );
  AND2_X1 U15181 ( .A1(n11988), .A2(n11987), .ZN(n11989) );
  NAND2_X1 U15182 ( .A1(n11991), .A2(n11665), .ZN(n11992) );
  NAND2_X1 U15183 ( .A1(n11992), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13529) );
  NAND2_X1 U15184 ( .A1(n12025), .A2(P1_EAX_REG_0__SCAN_IN), .ZN(n11995) );
  NAND2_X1 U15185 ( .A1(n20999), .A2(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n11994) );
  OAI211_X1 U15186 ( .C1(n12013), .C2(n13523), .A(n11995), .B(n11994), .ZN(
        n11996) );
  AOI21_X1 U15187 ( .B1(n20422), .B2(n12154), .A(n11996), .ZN(n11997) );
  OR2_X1 U15188 ( .A1(n13529), .A2(n11997), .ZN(n13530) );
  INV_X1 U15189 ( .A(n11997), .ZN(n13531) );
  OR2_X1 U15190 ( .A1(n13531), .A2(n12742), .ZN(n11998) );
  NAND2_X1 U15191 ( .A1(n13530), .A2(n11998), .ZN(n13541) );
  NAND2_X1 U15192 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n12001) );
  INV_X1 U15193 ( .A(n12001), .ZN(n12000) );
  INV_X1 U15194 ( .A(n12010), .ZN(n12004) );
  INV_X1 U15195 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n12002) );
  NAND2_X1 U15196 ( .A1(n12002), .A2(n12001), .ZN(n12003) );
  NAND2_X1 U15197 ( .A1(n12004), .A2(n12003), .ZN(n13890) );
  AOI22_X1 U15198 ( .A1(n13890), .A2(n12847), .B1(n12747), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n12007) );
  NAND2_X1 U15199 ( .A1(n12748), .A2(P1_EAX_REG_3__SCAN_IN), .ZN(n12006) );
  OAI211_X1 U15200 ( .C1(n12013), .C2(n11535), .A(n12007), .B(n12006), .ZN(
        n12008) );
  INV_X1 U15201 ( .A(n12008), .ZN(n12009) );
  OAI21_X2 U15202 ( .B1(n20594), .B2(n12143), .A(n12009), .ZN(n13852) );
  NAND2_X1 U15203 ( .A1(n12010), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12019) );
  OAI21_X1 U15204 ( .B1(n12010), .B2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n12019), .ZN(n20251) );
  INV_X1 U15205 ( .A(n20251), .ZN(n20155) );
  NAND2_X1 U15206 ( .A1(n20999), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12012) );
  NAND2_X1 U15207 ( .A1(n12748), .A2(P1_EAX_REG_4__SCAN_IN), .ZN(n12011) );
  OAI211_X1 U15208 ( .C1(n12013), .C2(n13478), .A(n12012), .B(n12011), .ZN(
        n12014) );
  NAND2_X1 U15209 ( .A1(n12014), .A2(n12742), .ZN(n12015) );
  OAI21_X1 U15210 ( .B1(n20155), .B2(n12742), .A(n12015), .ZN(n12016) );
  AOI21_X1 U15211 ( .B1(n12017), .B2(n12154), .A(n12016), .ZN(n14016) );
  NOR2_X2 U15212 ( .A1(n13851), .A2(n14016), .ZN(n14022) );
  NAND2_X1 U15213 ( .A1(n12018), .A2(n12154), .ZN(n12024) );
  INV_X1 U15214 ( .A(n12747), .ZN(n12086) );
  AND2_X1 U15215 ( .A1(n12019), .A2(n21092), .ZN(n12020) );
  OR2_X1 U15216 ( .A1(n12020), .A2(n12026), .ZN(n20142) );
  NAND2_X1 U15217 ( .A1(n20142), .A2(n12847), .ZN(n12021) );
  OAI21_X1 U15218 ( .B1(n21092), .B2(n12086), .A(n12021), .ZN(n12022) );
  AOI21_X1 U15219 ( .B1(n12748), .B2(P1_EAX_REG_5__SCAN_IN), .A(n12022), .ZN(
        n12023) );
  NAND2_X1 U15220 ( .A1(n12024), .A2(n12023), .ZN(n14021) );
  NAND2_X1 U15221 ( .A1(n14022), .A2(n14021), .ZN(n14020) );
  INV_X1 U15222 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n12029) );
  NOR2_X1 U15223 ( .A1(n12026), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12027) );
  OR2_X1 U15224 ( .A1(n12032), .A2(n12027), .ZN(n20127) );
  AOI22_X1 U15225 ( .A1(n20127), .A2(n12847), .B1(n12747), .B2(
        P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n12028) );
  OAI21_X1 U15226 ( .B1(n12005), .B2(n12029), .A(n12028), .ZN(n12030) );
  AOI21_X1 U15227 ( .B1(n12031), .B2(n12154), .A(n12030), .ZN(n14249) );
  INV_X1 U15228 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n12035) );
  OR2_X1 U15229 ( .A1(n12032), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12033) );
  NAND2_X1 U15230 ( .A1(n12033), .A2(n12054), .ZN(n20113) );
  AOI22_X1 U15231 ( .A1(n20113), .A2(n12847), .B1(n12747), .B2(
        P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n12034) );
  OAI21_X1 U15232 ( .B1(n12005), .B2(n12035), .A(n12034), .ZN(n12036) );
  AOI22_X1 U15233 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n12116), .B1(
        n9817), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12042) );
  AOI22_X1 U15234 ( .A1(n12374), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n9850), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12041) );
  AOI22_X1 U15235 ( .A1(n12250), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n12702), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12040) );
  AOI22_X1 U15236 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n12732), .B1(
        n11622), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12039) );
  NAND4_X1 U15237 ( .A1(n12042), .A2(n12041), .A3(n12040), .A4(n12039), .ZN(
        n12049) );
  AOI22_X1 U15238 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n9838), .B1(
        n12286), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12047) );
  AOI22_X1 U15239 ( .A1(n12729), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12731), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12046) );
  AOI22_X1 U15240 ( .A1(n9852), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n10016), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12045) );
  AOI22_X1 U15241 ( .A1(n12724), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12185), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12044) );
  NAND4_X1 U15242 ( .A1(n12047), .A2(n12046), .A3(n12045), .A4(n12044), .ZN(
        n12048) );
  OAI21_X1 U15243 ( .B1(n12049), .B2(n12048), .A(n12154), .ZN(n12053) );
  INV_X1 U15244 ( .A(n12054), .ZN(n12050) );
  XNOR2_X1 U15245 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B(n12050), .ZN(
        n14472) );
  AOI22_X1 U15246 ( .A1(n12847), .A2(n14472), .B1(n12747), .B2(
        P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n12052) );
  NAND2_X1 U15247 ( .A1(n12025), .A2(P1_EAX_REG_8__SCAN_IN), .ZN(n12051) );
  XNOR2_X1 U15248 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .B(n12079), .ZN(
        n20107) );
  INV_X1 U15249 ( .A(n20107), .ZN(n14512) );
  AOI22_X1 U15250 ( .A1(n9838), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12374), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12058) );
  AOI22_X1 U15251 ( .A1(n12729), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12731), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12057) );
  AOI22_X1 U15252 ( .A1(n12116), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n9852), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12056) );
  AOI22_X1 U15253 ( .A1(n12250), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n12702), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12055) );
  NAND4_X1 U15254 ( .A1(n12058), .A2(n12057), .A3(n12056), .A4(n12055), .ZN(
        n12064) );
  AOI22_X1 U15255 ( .A1(n9817), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n9850), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12062) );
  AOI22_X1 U15256 ( .A1(n12286), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n12356), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12060) );
  AOI22_X1 U15257 ( .A1(n9849), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11716), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12059) );
  NAND4_X1 U15258 ( .A1(n12062), .A2(n12061), .A3(n12060), .A4(n12059), .ZN(
        n12063) );
  OAI21_X1 U15259 ( .B1(n12064), .B2(n12063), .A(n12154), .ZN(n12067) );
  NAND2_X1 U15260 ( .A1(n12025), .A2(P1_EAX_REG_9__SCAN_IN), .ZN(n12066) );
  NAND2_X1 U15261 ( .A1(n12747), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n12065) );
  NAND3_X1 U15262 ( .A1(n12067), .A2(n12066), .A3(n12065), .ZN(n12068) );
  AOI21_X1 U15263 ( .B1(n14512), .B2(n12847), .A(n12068), .ZN(n14494) );
  AOI22_X1 U15264 ( .A1(n12116), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12729), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12072) );
  AOI22_X1 U15265 ( .A1(n9817), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n9851), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12071) );
  AOI22_X1 U15266 ( .A1(n9838), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n9825), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12070) );
  AOI22_X1 U15267 ( .A1(n12250), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n12702), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12069) );
  NAND4_X1 U15268 ( .A1(n12072), .A2(n12071), .A3(n12070), .A4(n12069), .ZN(
        n12078) );
  AOI22_X1 U15269 ( .A1(n12286), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12732), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12076) );
  AOI22_X1 U15270 ( .A1(n12731), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n11622), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12075) );
  AOI22_X1 U15271 ( .A1(n12374), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n10016), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12074) );
  AOI22_X1 U15272 ( .A1(n12724), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11716), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12073) );
  NAND4_X1 U15273 ( .A1(n12076), .A2(n12075), .A3(n12074), .A4(n12073), .ZN(
        n12077) );
  NOR2_X1 U15274 ( .A1(n12078), .A2(n12077), .ZN(n12082) );
  XNOR2_X1 U15275 ( .A(n12083), .B(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n15269) );
  NAND2_X1 U15276 ( .A1(n15269), .A2(n12847), .ZN(n12081) );
  AOI22_X1 U15277 ( .A1(n12748), .A2(P1_EAX_REG_10__SCAN_IN), .B1(n12747), 
        .B2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n12080) );
  OAI211_X1 U15278 ( .C1(n12082), .C2(n12143), .A(n12081), .B(n12080), .ZN(
        n14458) );
  NAND2_X1 U15279 ( .A1(n14456), .A2(n14458), .ZN(n14457) );
  INV_X1 U15280 ( .A(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n12087) );
  OAI21_X1 U15281 ( .B1(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n12084), .A(
        n12127), .ZN(n16328) );
  NAND2_X1 U15282 ( .A1(n16328), .A2(n12847), .ZN(n12085) );
  OAI21_X1 U15283 ( .B1(n12087), .B2(n12086), .A(n12085), .ZN(n12088) );
  AOI21_X1 U15284 ( .B1(n12025), .B2(P1_EAX_REG_11__SCAN_IN), .A(n12088), .ZN(
        n14977) );
  AOI22_X1 U15285 ( .A1(n9838), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12374), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12093) );
  AOI22_X1 U15286 ( .A1(n12116), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n9851), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12092) );
  AOI22_X1 U15287 ( .A1(n12250), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n12702), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12091) );
  AOI22_X1 U15288 ( .A1(n12286), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n10016), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12090) );
  NAND4_X1 U15289 ( .A1(n12093), .A2(n12092), .A3(n12091), .A4(n12090), .ZN(
        n12099) );
  AOI22_X1 U15290 ( .A1(n9817), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12731), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12097) );
  AOI22_X1 U15291 ( .A1(n12729), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n9825), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12096) );
  AOI22_X1 U15292 ( .A1(n12732), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11622), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12095) );
  AOI22_X1 U15293 ( .A1(n9848), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11716), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12094) );
  NAND4_X1 U15294 ( .A1(n12097), .A2(n12096), .A3(n12095), .A4(n12094), .ZN(
        n12098) );
  OR2_X1 U15295 ( .A1(n12099), .A2(n12098), .ZN(n12100) );
  NAND2_X1 U15296 ( .A1(n12154), .A2(n12100), .ZN(n15047) );
  INV_X1 U15297 ( .A(n15047), .ZN(n12101) );
  XNOR2_X1 U15298 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .B(n12140), .ZN(
        n15249) );
  AOI22_X1 U15299 ( .A1(n9817), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12286), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12106) );
  AOI22_X1 U15300 ( .A1(n12116), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12732), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12105) );
  AOI22_X1 U15301 ( .A1(n9838), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12731), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12104) );
  AOI22_X1 U15302 ( .A1(n9848), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12185), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12103) );
  NAND4_X1 U15303 ( .A1(n12106), .A2(n12105), .A3(n12104), .A4(n12103), .ZN(
        n12112) );
  AOI22_X1 U15304 ( .A1(n12374), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n9825), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12110) );
  AOI22_X1 U15305 ( .A1(n9850), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n12356), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12109) );
  AOI22_X1 U15306 ( .A1(n12250), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n12702), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12107) );
  NAND4_X1 U15307 ( .A1(n12110), .A2(n12109), .A3(n12108), .A4(n12107), .ZN(
        n12111) );
  OR2_X1 U15308 ( .A1(n12112), .A2(n12111), .ZN(n12113) );
  AOI22_X1 U15309 ( .A1(n12154), .A2(n12113), .B1(n12747), .B2(
        P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n12115) );
  NAND2_X1 U15310 ( .A1(n12025), .A2(P1_EAX_REG_13__SCAN_IN), .ZN(n12114) );
  OAI211_X1 U15311 ( .C1(n15249), .C2(n12742), .A(n12115), .B(n12114), .ZN(
        n14979) );
  INV_X1 U15312 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n15114) );
  AOI22_X1 U15313 ( .A1(n9838), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n9826), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12120) );
  AOI22_X1 U15314 ( .A1(n12116), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12356), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12119) );
  AOI22_X1 U15315 ( .A1(n12250), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n12702), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12117) );
  NAND4_X1 U15316 ( .A1(n12120), .A2(n12119), .A3(n12118), .A4(n12117), .ZN(
        n12126) );
  AOI22_X1 U15317 ( .A1(n9817), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12732), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12124) );
  AOI22_X1 U15318 ( .A1(n12729), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12374), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12123) );
  AOI22_X1 U15319 ( .A1(n9851), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n12731), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12122) );
  AOI22_X1 U15320 ( .A1(n12724), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n12185), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12121) );
  NAND4_X1 U15321 ( .A1(n12124), .A2(n12123), .A3(n12122), .A4(n12121), .ZN(
        n12125) );
  OAI21_X1 U15322 ( .B1(n12126), .B2(n12125), .A(n12154), .ZN(n12129) );
  XNOR2_X1 U15323 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B(n12127), .ZN(
        n16277) );
  INV_X1 U15324 ( .A(n16277), .ZN(n15260) );
  AOI22_X1 U15325 ( .A1(n12747), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        n12847), .B2(n15260), .ZN(n12128) );
  OAI211_X1 U15326 ( .C1(n12005), .C2(n15114), .A(n12129), .B(n12128), .ZN(
        n15035) );
  AOI22_X1 U15327 ( .A1(n12116), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12729), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12133) );
  AOI22_X1 U15328 ( .A1(n9817), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n9852), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12132) );
  AOI22_X1 U15329 ( .A1(n12250), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n12702), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12130) );
  NAND4_X1 U15330 ( .A1(n12133), .A2(n12132), .A3(n12131), .A4(n12130), .ZN(
        n12139) );
  AOI22_X1 U15331 ( .A1(n12732), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n9851), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12137) );
  AOI22_X1 U15332 ( .A1(n12374), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n12731), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12136) );
  AOI22_X1 U15333 ( .A1(n9838), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12356), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12135) );
  AOI22_X1 U15334 ( .A1(n9849), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12185), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12134) );
  NAND4_X1 U15335 ( .A1(n12137), .A2(n12136), .A3(n12135), .A4(n12134), .ZN(
        n12138) );
  NOR2_X1 U15336 ( .A1(n12139), .A2(n12138), .ZN(n12144) );
  XNOR2_X1 U15337 ( .A(n12145), .B(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n16267) );
  NAND2_X1 U15338 ( .A1(n16267), .A2(n12847), .ZN(n12142) );
  AOI22_X1 U15339 ( .A1(n12748), .A2(P1_EAX_REG_14__SCAN_IN), .B1(n12747), 
        .B2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n12141) );
  OAI211_X1 U15340 ( .C1(n12144), .C2(n12143), .A(n12142), .B(n12141), .ZN(
        n15028) );
  XNOR2_X1 U15341 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B(n12162), .ZN(
        n16317) );
  INV_X1 U15342 ( .A(n16317), .ZN(n12161) );
  AOI22_X1 U15343 ( .A1(n12116), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12732), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12149) );
  AOI22_X1 U15344 ( .A1(n9817), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n9851), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12148) );
  AOI22_X1 U15345 ( .A1(n9838), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n9852), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12147) );
  AOI22_X1 U15346 ( .A1(n12250), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n12702), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12146) );
  NAND4_X1 U15347 ( .A1(n12149), .A2(n12148), .A3(n12147), .A4(n12146), .ZN(
        n12156) );
  AOI22_X1 U15348 ( .A1(n12374), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n12731), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12153) );
  AOI22_X1 U15349 ( .A1(n12286), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n11622), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12152) );
  AOI22_X1 U15350 ( .A1(n9849), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12185), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12150) );
  NAND4_X1 U15351 ( .A1(n12153), .A2(n12152), .A3(n12151), .A4(n12150), .ZN(
        n12155) );
  OAI21_X1 U15352 ( .B1(n12156), .B2(n12155), .A(n12154), .ZN(n12159) );
  NAND2_X1 U15353 ( .A1(n12025), .A2(P1_EAX_REG_15__SCAN_IN), .ZN(n12158) );
  NAND2_X1 U15354 ( .A1(n12747), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n12157) );
  NAND3_X1 U15355 ( .A1(n12159), .A2(n12158), .A3(n12157), .ZN(n12160) );
  AOI21_X1 U15356 ( .B1(n12161), .B2(n12847), .A(n12160), .ZN(n15026) );
  INV_X1 U15357 ( .A(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n15227) );
  XNOR2_X1 U15358 ( .A(n12180), .B(n15227), .ZN(n15230) );
  NAND2_X1 U15359 ( .A1(n15230), .A2(n12847), .ZN(n12178) );
  AOI22_X1 U15360 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n12729), .B1(
        n12038), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12166) );
  AOI22_X1 U15361 ( .A1(n12732), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n12731), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12165) );
  AOI22_X1 U15362 ( .A1(n12374), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n12356), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12164) );
  AOI22_X1 U15363 ( .A1(n9850), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n12702), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12163) );
  NAND4_X1 U15364 ( .A1(n12166), .A2(n12165), .A3(n12164), .A4(n12163), .ZN(
        n12174) );
  AOI22_X1 U15365 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n9817), .B1(
        n12286), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12172) );
  AOI22_X1 U15366 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n9838), .B1(
        n9826), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12171) );
  NAND2_X1 U15367 ( .A1(n12250), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n12168) );
  NAND2_X1 U15368 ( .A1(n11716), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n12167) );
  AND3_X1 U15369 ( .A1(n12168), .A2(n12742), .A3(n12167), .ZN(n12169) );
  NAND4_X1 U15370 ( .A1(n12172), .A2(n12171), .A3(n12170), .A4(n12169), .ZN(
        n12173) );
  NAND2_X1 U15371 ( .A1(n12717), .A2(n12742), .ZN(n12276) );
  OAI21_X1 U15372 ( .B1(n12174), .B2(n12173), .A(n12276), .ZN(n12176) );
  AOI22_X1 U15373 ( .A1(n12748), .A2(P1_EAX_REG_16__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n20999), .ZN(n12175) );
  NAND2_X1 U15374 ( .A1(n12176), .A2(n12175), .ZN(n12177) );
  NAND2_X1 U15375 ( .A1(n12178), .A2(n12177), .ZN(n14963) );
  XNOR2_X1 U15376 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B(n12194), .ZN(
        n16306) );
  AOI22_X1 U15377 ( .A1(n12748), .A2(P1_EAX_REG_17__SCAN_IN), .B1(n12747), 
        .B2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n12193) );
  AOI22_X1 U15378 ( .A1(n9838), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12374), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12184) );
  AOI22_X1 U15379 ( .A1(n12116), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12731), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12183) );
  AOI22_X1 U15380 ( .A1(n9851), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(n9852), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12182) );
  AOI22_X1 U15381 ( .A1(n12250), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n12702), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12181) );
  NAND4_X1 U15382 ( .A1(n12184), .A2(n12183), .A3(n12182), .A4(n12181), .ZN(
        n12191) );
  AOI22_X1 U15383 ( .A1(n12729), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12732), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12189) );
  AOI22_X1 U15384 ( .A1(n12286), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12356), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12188) );
  AOI22_X1 U15385 ( .A1(n9849), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12185), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12186) );
  NAND4_X1 U15386 ( .A1(n12189), .A2(n12188), .A3(n12187), .A4(n12186), .ZN(
        n12190) );
  OAI21_X1 U15387 ( .B1(n12191), .B2(n12190), .A(n12744), .ZN(n12192) );
  OAI211_X1 U15388 ( .C1(n16306), .C2(n12742), .A(n12193), .B(n12192), .ZN(
        n14942) );
  INV_X1 U15389 ( .A(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n12195) );
  XNOR2_X1 U15390 ( .A(n12210), .B(n12195), .ZN(n16247) );
  AOI22_X1 U15391 ( .A1(n12748), .A2(P1_EAX_REG_18__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n20999), .ZN(n12209) );
  AOI22_X1 U15392 ( .A1(n9838), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11599), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12199) );
  AOI22_X1 U15393 ( .A1(n12116), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n9852), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12198) );
  AOI22_X1 U15394 ( .A1(n12374), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n12702), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12196) );
  NAND4_X1 U15395 ( .A1(n12199), .A2(n12198), .A3(n12197), .A4(n12196), .ZN(
        n12207) );
  AOI22_X1 U15396 ( .A1(n12729), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12286), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12205) );
  AOI22_X1 U15397 ( .A1(n12724), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12731), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12204) );
  AOI22_X1 U15398 ( .A1(n9817), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12356), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12203) );
  NAND2_X1 U15399 ( .A1(n12250), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(
        n12201) );
  NAND2_X1 U15400 ( .A1(n12185), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n12200) );
  AND3_X1 U15401 ( .A1(n12201), .A2(n12742), .A3(n12200), .ZN(n12202) );
  NAND4_X1 U15402 ( .A1(n12205), .A2(n12204), .A3(n12203), .A4(n12202), .ZN(
        n12206) );
  OAI21_X1 U15403 ( .B1(n12207), .B2(n12206), .A(n12276), .ZN(n12208) );
  AOI22_X1 U15404 ( .A1(n16247), .A2(n12847), .B1(n12209), .B2(n12208), .ZN(
        n15012) );
  INV_X1 U15405 ( .A(n12211), .ZN(n12213) );
  INV_X1 U15406 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n12212) );
  NAND2_X1 U15407 ( .A1(n12213), .A2(n12212), .ZN(n12214) );
  NAND2_X1 U15408 ( .A1(n12246), .A2(n12214), .ZN(n16240) );
  OR2_X1 U15409 ( .A1(n16240), .A2(n12742), .ZN(n12229) );
  AOI22_X1 U15410 ( .A1(n12116), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n9817), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12218) );
  AOI22_X1 U15411 ( .A1(n9850), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(n9825), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12217) );
  AOI22_X1 U15412 ( .A1(n12250), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n12702), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12215) );
  NAND4_X1 U15413 ( .A1(n12218), .A2(n12217), .A3(n12216), .A4(n12215), .ZN(
        n12224) );
  AOI22_X1 U15414 ( .A1(n12286), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12374), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12222) );
  AOI22_X1 U15415 ( .A1(n9838), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12731), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12221) );
  AOI22_X1 U15416 ( .A1(n12732), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12356), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12220) );
  AOI22_X1 U15417 ( .A1(n9848), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11716), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12219) );
  NAND4_X1 U15418 ( .A1(n12222), .A2(n12221), .A3(n12220), .A4(n12219), .ZN(
        n12223) );
  NOR2_X1 U15419 ( .A1(n12224), .A2(n12223), .ZN(n12227) );
  INV_X1 U15420 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n21000) );
  OAI21_X1 U15421 ( .B1(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n21000), .A(
        n20999), .ZN(n12226) );
  NAND2_X1 U15422 ( .A1(n12025), .A2(P1_EAX_REG_19__SCAN_IN), .ZN(n12225) );
  OAI211_X1 U15423 ( .C1(n12717), .C2(n12227), .A(n12226), .B(n12225), .ZN(
        n12228) );
  NAND2_X1 U15424 ( .A1(n12229), .A2(n12228), .ZN(n15005) );
  XNOR2_X1 U15425 ( .A(n12246), .B(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15204) );
  NAND2_X1 U15426 ( .A1(n15204), .A2(n12847), .ZN(n12245) );
  AOI22_X1 U15427 ( .A1(n12116), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12729), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12233) );
  AOI22_X1 U15428 ( .A1(n12374), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n12356), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12232) );
  AOI22_X1 U15429 ( .A1(n9850), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n12722), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12230) );
  NAND4_X1 U15430 ( .A1(n12233), .A2(n12232), .A3(n12231), .A4(n12230), .ZN(
        n12241) );
  AOI22_X1 U15431 ( .A1(n12732), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n9848), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12239) );
  AOI22_X1 U15432 ( .A1(n9817), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12731), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12238) );
  AOI22_X1 U15433 ( .A1(n9838), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n9825), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12237) );
  NAND2_X1 U15434 ( .A1(n12250), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n12235) );
  NAND2_X1 U15435 ( .A1(n12185), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n12234) );
  AND3_X1 U15436 ( .A1(n12235), .A2(n12742), .A3(n12234), .ZN(n12236) );
  NAND4_X1 U15437 ( .A1(n12239), .A2(n12238), .A3(n12237), .A4(n12236), .ZN(
        n12240) );
  OAI21_X1 U15438 ( .B1(n12241), .B2(n12240), .A(n12276), .ZN(n12243) );
  AOI22_X1 U15439 ( .A1(n12748), .A2(P1_EAX_REG_20__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n20999), .ZN(n12242) );
  NAND2_X1 U15440 ( .A1(n12243), .A2(n12242), .ZN(n12244) );
  NAND2_X1 U15441 ( .A1(n12245), .A2(n12244), .ZN(n14928) );
  NOR2_X2 U15442 ( .A1(n14929), .A2(n14928), .ZN(n14915) );
  INV_X1 U15443 ( .A(n12247), .ZN(n12248) );
  INV_X1 U15444 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n21259) );
  NAND2_X1 U15445 ( .A1(n12248), .A2(n21259), .ZN(n12249) );
  NAND2_X1 U15446 ( .A1(n12281), .A2(n12249), .ZN(n15195) );
  OR2_X1 U15447 ( .A1(n15195), .A2(n12742), .ZN(n12265) );
  AOI22_X1 U15448 ( .A1(n9838), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n9817), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12254) );
  AOI22_X1 U15449 ( .A1(n12286), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12732), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12253) );
  AOI22_X1 U15450 ( .A1(n12250), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n12722), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12252) );
  AOI22_X1 U15451 ( .A1(n12729), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12356), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12251) );
  NAND4_X1 U15452 ( .A1(n12254), .A2(n12253), .A3(n12252), .A4(n12251), .ZN(
        n12260) );
  AOI22_X1 U15453 ( .A1(n12116), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12374), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12258) );
  AOI22_X1 U15454 ( .A1(n9851), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n12731), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12257) );
  AOI22_X1 U15455 ( .A1(n9848), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12185), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12255) );
  NAND4_X1 U15456 ( .A1(n12258), .A2(n12257), .A3(n12256), .A4(n12255), .ZN(
        n12259) );
  NOR2_X1 U15457 ( .A1(n12260), .A2(n12259), .ZN(n12263) );
  OAI21_X1 U15458 ( .B1(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n21000), .A(
        n20999), .ZN(n12262) );
  NAND2_X1 U15459 ( .A1(n12748), .A2(P1_EAX_REG_21__SCAN_IN), .ZN(n12261) );
  OAI211_X1 U15460 ( .C1(n12717), .C2(n12263), .A(n12262), .B(n12261), .ZN(
        n12264) );
  XNOR2_X1 U15461 ( .A(n12281), .B(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15189) );
  AOI22_X1 U15462 ( .A1(n12748), .A2(P1_EAX_REG_22__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n20999), .ZN(n12280) );
  AOI22_X1 U15463 ( .A1(n12038), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12286), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12269) );
  AOI22_X1 U15464 ( .A1(n12729), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12732), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12268) );
  AOI22_X1 U15465 ( .A1(n9817), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12702), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12267) );
  AOI22_X1 U15466 ( .A1(n9851), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n11622), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12266) );
  NAND4_X1 U15467 ( .A1(n12269), .A2(n12268), .A3(n12267), .A4(n12266), .ZN(
        n12278) );
  AOI22_X1 U15468 ( .A1(n9849), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12731), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12275) );
  AOI22_X1 U15469 ( .A1(n9838), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n9826), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12274) );
  AOI22_X1 U15470 ( .A1(n12374), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n10016), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12273) );
  NAND2_X1 U15471 ( .A1(n12250), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n12271) );
  NAND2_X1 U15472 ( .A1(n11716), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n12270) );
  AND3_X1 U15473 ( .A1(n12271), .A2(n12742), .A3(n12270), .ZN(n12272) );
  NAND4_X1 U15474 ( .A1(n12275), .A2(n12274), .A3(n12273), .A4(n12272), .ZN(
        n12277) );
  OAI21_X1 U15475 ( .B1(n12278), .B2(n12277), .A(n12276), .ZN(n12279) );
  AOI22_X1 U15476 ( .A1(n15189), .A2(n12847), .B1(n12280), .B2(n12279), .ZN(
        n14901) );
  INV_X1 U15477 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n15185) );
  XNOR2_X1 U15478 ( .A(n12327), .B(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15169) );
  NAND2_X1 U15479 ( .A1(n15169), .A2(n12847), .ZN(n12318) );
  AOI22_X1 U15480 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n12116), .B1(
        n9838), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12285) );
  AOI22_X1 U15481 ( .A1(n12374), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n12702), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12284) );
  AOI22_X1 U15482 ( .A1(n9850), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10016), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12283) );
  AOI22_X1 U15483 ( .A1(n12724), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11716), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12282) );
  NAND4_X1 U15484 ( .A1(n12285), .A2(n12284), .A3(n12283), .A4(n12282), .ZN(
        n12292) );
  AOI22_X1 U15485 ( .A1(P1_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n12732), .B1(
        n12731), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12290) );
  AOI22_X1 U15486 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n12729), .B1(
        n9852), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12289) );
  AOI22_X1 U15487 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n12286), .B1(
        n12356), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12288) );
  AOI22_X1 U15488 ( .A1(n9817), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12250), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12287) );
  NAND4_X1 U15489 ( .A1(n12290), .A2(n12289), .A3(n12288), .A4(n12287), .ZN(
        n12291) );
  NOR2_X1 U15490 ( .A1(n12292), .A2(n12291), .ZN(n12322) );
  AOI22_X1 U15491 ( .A1(n9817), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n9851), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12296) );
  AOI22_X1 U15492 ( .A1(n12729), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n10016), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12295) );
  AOI22_X1 U15493 ( .A1(n12250), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n12702), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12294) );
  AOI22_X1 U15494 ( .A1(n9849), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12185), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12293) );
  NAND4_X1 U15495 ( .A1(n12296), .A2(n12295), .A3(n12294), .A4(n12293), .ZN(
        n12302) );
  AOI22_X1 U15496 ( .A1(n9838), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12374), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12300) );
  AOI22_X1 U15497 ( .A1(n12732), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12731), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12299) );
  AOI22_X1 U15498 ( .A1(n12116), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n9826), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12298) );
  AOI22_X1 U15499 ( .A1(n12286), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12356), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12297) );
  NAND4_X1 U15500 ( .A1(n12300), .A2(n12299), .A3(n12298), .A4(n12297), .ZN(
        n12301) );
  NOR2_X1 U15501 ( .A1(n12302), .A2(n12301), .ZN(n12321) );
  NOR2_X1 U15502 ( .A1(n12322), .A2(n12321), .ZN(n12343) );
  AOI22_X1 U15503 ( .A1(n12116), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n9817), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12306) );
  AOI22_X1 U15504 ( .A1(n9838), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n12374), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12305) );
  AOI22_X1 U15505 ( .A1(n9850), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(n9852), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12304) );
  AOI22_X1 U15506 ( .A1(n12250), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n12702), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12303) );
  NAND4_X1 U15507 ( .A1(n12306), .A2(n12305), .A3(n12304), .A4(n12303), .ZN(
        n12312) );
  AOI22_X1 U15508 ( .A1(n12732), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12731), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12310) );
  AOI22_X1 U15509 ( .A1(n12729), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11622), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12309) );
  AOI22_X1 U15510 ( .A1(n12286), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n10016), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12308) );
  AOI22_X1 U15511 ( .A1(n12724), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12185), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12307) );
  NAND4_X1 U15512 ( .A1(n12310), .A2(n12309), .A3(n12308), .A4(n12307), .ZN(
        n12311) );
  OR2_X1 U15513 ( .A1(n12312), .A2(n12311), .ZN(n12342) );
  XNOR2_X1 U15514 ( .A(n12343), .B(n12342), .ZN(n12316) );
  NAND2_X1 U15515 ( .A1(n20999), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n12313) );
  NAND2_X1 U15516 ( .A1(n12742), .A2(n12313), .ZN(n12314) );
  AOI21_X1 U15517 ( .B1(n12025), .B2(P1_EAX_REG_24__SCAN_IN), .A(n12314), .ZN(
        n12315) );
  OAI21_X1 U15518 ( .B1(n12316), .B2(n12717), .A(n12315), .ZN(n12317) );
  NAND2_X1 U15519 ( .A1(n12318), .A2(n12317), .ZN(n14875) );
  NAND2_X1 U15520 ( .A1(n12319), .A2(n14890), .ZN(n12320) );
  NAND2_X1 U15521 ( .A1(n12327), .A2(n12320), .ZN(n15176) );
  XNOR2_X1 U15522 ( .A(n12322), .B(n12321), .ZN(n12323) );
  NOR2_X1 U15523 ( .A1(n12323), .A2(n12717), .ZN(n12326) );
  INV_X1 U15524 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n15070) );
  NAND2_X1 U15525 ( .A1(n20999), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n12324) );
  OAI211_X1 U15526 ( .C1(n12005), .C2(n15070), .A(n12742), .B(n12324), .ZN(
        n12325) );
  OAI22_X1 U15527 ( .A1(n15176), .A2(n12742), .B1(n12326), .B2(n12325), .ZN(
        n14888) );
  INV_X1 U15528 ( .A(n12328), .ZN(n12330) );
  INV_X1 U15529 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n12329) );
  NAND2_X1 U15530 ( .A1(n12330), .A2(n12329), .ZN(n12331) );
  NAND2_X1 U15531 ( .A1(n12368), .A2(n12331), .ZN(n15160) );
  AOI22_X1 U15532 ( .A1(n12729), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12374), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12335) );
  AOI22_X1 U15533 ( .A1(n12731), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12356), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12334) );
  AOI22_X1 U15534 ( .A1(n9826), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n12722), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12333) );
  AOI22_X1 U15535 ( .A1(n9849), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12185), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12332) );
  NAND4_X1 U15536 ( .A1(n12335), .A2(n12334), .A3(n12333), .A4(n12332), .ZN(
        n12341) );
  AOI22_X1 U15537 ( .A1(n9838), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n12116), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12339) );
  AOI22_X1 U15538 ( .A1(n9817), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12286), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12338) );
  AOI22_X1 U15539 ( .A1(n9850), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12250), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12337) );
  AOI22_X1 U15540 ( .A1(n12732), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n10016), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12336) );
  NAND4_X1 U15541 ( .A1(n12339), .A2(n12338), .A3(n12337), .A4(n12336), .ZN(
        n12340) );
  NOR2_X1 U15542 ( .A1(n12341), .A2(n12340), .ZN(n12351) );
  NAND2_X1 U15543 ( .A1(n12343), .A2(n12342), .ZN(n12350) );
  XNOR2_X1 U15544 ( .A(n12351), .B(n12350), .ZN(n12347) );
  NAND2_X1 U15545 ( .A1(n20999), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n12344) );
  NAND2_X1 U15546 ( .A1(n12742), .A2(n12344), .ZN(n12345) );
  AOI21_X1 U15547 ( .B1(n12025), .B2(P1_EAX_REG_25__SCAN_IN), .A(n12345), .ZN(
        n12346) );
  OAI21_X1 U15548 ( .B1(n12347), .B2(n12717), .A(n12346), .ZN(n12348) );
  NAND2_X1 U15549 ( .A1(n12349), .A2(n12348), .ZN(n14860) );
  XNOR2_X1 U15550 ( .A(n12368), .B(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15152) );
  NOR2_X1 U15551 ( .A1(n12351), .A2(n12350), .ZN(n12386) );
  AOI22_X1 U15552 ( .A1(n12116), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n9817), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12355) );
  AOI22_X1 U15553 ( .A1(n9838), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n11612), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12354) );
  AOI22_X1 U15554 ( .A1(n9851), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(n9825), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12353) );
  AOI22_X1 U15555 ( .A1(n12250), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n12722), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12352) );
  NAND4_X1 U15556 ( .A1(n12355), .A2(n12354), .A3(n12353), .A4(n12352), .ZN(
        n12362) );
  AOI22_X1 U15557 ( .A1(n12732), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12731), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12360) );
  AOI22_X1 U15558 ( .A1(n12729), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12356), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12359) );
  AOI22_X1 U15559 ( .A1(n9848), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12185), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12357) );
  NAND4_X1 U15560 ( .A1(n12360), .A2(n12359), .A3(n12358), .A4(n12357), .ZN(
        n12361) );
  OR2_X1 U15561 ( .A1(n12362), .A2(n12361), .ZN(n12385) );
  INV_X1 U15562 ( .A(n12385), .ZN(n12363) );
  XNOR2_X1 U15563 ( .A(n12386), .B(n12363), .ZN(n12366) );
  INV_X1 U15564 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n15059) );
  NAND2_X1 U15565 ( .A1(n20999), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12364) );
  OAI211_X1 U15566 ( .C1(n12005), .C2(n15059), .A(n12742), .B(n12364), .ZN(
        n12365) );
  AOI21_X1 U15567 ( .B1(n12366), .B2(n12744), .A(n12365), .ZN(n12367) );
  AOI21_X1 U15568 ( .B1(n15152), .B2(n12847), .A(n12367), .ZN(n14854) );
  INV_X1 U15569 ( .A(n12368), .ZN(n12369) );
  INV_X1 U15570 ( .A(n12370), .ZN(n12372) );
  INV_X1 U15571 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n12371) );
  NAND2_X1 U15572 ( .A1(n12372), .A2(n12371), .ZN(n12373) );
  NAND2_X1 U15573 ( .A1(n12697), .A2(n12373), .ZN(n15140) );
  AOI22_X1 U15574 ( .A1(n9838), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n12374), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12378) );
  AOI22_X1 U15575 ( .A1(n9817), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12731), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12377) );
  AOI22_X1 U15576 ( .A1(n12250), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n12702), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12376) );
  AOI22_X1 U15577 ( .A1(n12724), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12185), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12375) );
  NAND4_X1 U15578 ( .A1(n12378), .A2(n12377), .A3(n12376), .A4(n12375), .ZN(
        n12384) );
  AOI22_X1 U15579 ( .A1(n12729), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n12286), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12382) );
  AOI22_X1 U15580 ( .A1(n11599), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n9852), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12381) );
  AOI22_X1 U15581 ( .A1(n12116), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n11622), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12380) );
  AOI22_X1 U15582 ( .A1(n12732), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n10016), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12379) );
  NAND4_X1 U15583 ( .A1(n12382), .A2(n12381), .A3(n12380), .A4(n12379), .ZN(
        n12383) );
  NOR2_X1 U15584 ( .A1(n12384), .A2(n12383), .ZN(n12404) );
  NAND2_X1 U15585 ( .A1(n12386), .A2(n12385), .ZN(n12403) );
  XNOR2_X1 U15586 ( .A(n12404), .B(n12403), .ZN(n12389) );
  AOI21_X1 U15587 ( .B1(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n20999), .A(
        n12847), .ZN(n12388) );
  NAND2_X1 U15588 ( .A1(n12748), .A2(P1_EAX_REG_27__SCAN_IN), .ZN(n12387) );
  OAI211_X1 U15589 ( .C1(n12389), .C2(n12717), .A(n12388), .B(n12387), .ZN(
        n12390) );
  OAI21_X1 U15590 ( .B1(n15140), .B2(n12742), .A(n12390), .ZN(n14834) );
  XNOR2_X1 U15591 ( .A(n12697), .B(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14523) );
  INV_X1 U15592 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n12415) );
  AOI21_X1 U15593 ( .B1(n12415), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n12391) );
  AOI21_X1 U15594 ( .B1(n12025), .B2(P1_EAX_REG_28__SCAN_IN), .A(n12391), .ZN(
        n12407) );
  AOI22_X1 U15595 ( .A1(n12038), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n9817), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12396) );
  AOI22_X1 U15596 ( .A1(n9838), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n11612), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12395) );
  AOI22_X1 U15597 ( .A1(n9850), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(n9852), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12394) );
  AOI22_X1 U15598 ( .A1(n12250), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n12722), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12393) );
  NAND4_X1 U15599 ( .A1(n12396), .A2(n12395), .A3(n12394), .A4(n12393), .ZN(
        n12402) );
  AOI22_X1 U15600 ( .A1(n12732), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12731), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12400) );
  AOI22_X1 U15601 ( .A1(n12729), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11622), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12399) );
  AOI22_X1 U15602 ( .A1(n12286), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10016), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12398) );
  AOI22_X1 U15603 ( .A1(n9848), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12185), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12397) );
  NAND4_X1 U15604 ( .A1(n12400), .A2(n12399), .A3(n12398), .A4(n12397), .ZN(
        n12401) );
  OR2_X1 U15605 ( .A1(n12402), .A2(n12401), .ZN(n12713) );
  NOR2_X1 U15606 ( .A1(n12404), .A2(n12403), .ZN(n12714) );
  XOR2_X1 U15607 ( .A(n12713), .B(n12714), .Z(n12405) );
  NAND2_X1 U15608 ( .A1(n12405), .A2(n12744), .ZN(n12406) );
  AOI22_X1 U15609 ( .A1(n14523), .A2(n12847), .B1(n12407), .B2(n12406), .ZN(
        n12409) );
  OR2_X1 U15610 ( .A1(n12408), .A2(n12409), .ZN(n12410) );
  NAND2_X1 U15611 ( .A1(P1_STATEBS16_REG_SCAN_IN), .A2(n21002), .ZN(n16437) );
  INV_X1 U15612 ( .A(n16437), .ZN(n12411) );
  NOR2_X1 U15613 ( .A1(n14516), .A2(n20306), .ZN(n12420) );
  OR2_X1 U15614 ( .A1(n12414), .A2(n20769), .ZN(n21009) );
  AND2_X1 U15615 ( .A1(n21009), .A2(n20310), .ZN(n12412) );
  NAND2_X1 U15616 ( .A1(n21000), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n12413) );
  NOR2_X1 U15617 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n20999), .ZN(n16205) );
  INV_X1 U15618 ( .A(n16205), .ZN(n21004) );
  NAND2_X1 U15619 ( .A1(n12413), .A2(n21004), .ZN(n13537) );
  NAND2_X1 U15620 ( .A1(n16316), .A2(n14523), .ZN(n12418) );
  NAND2_X1 U15621 ( .A1(n20296), .A2(P1_REIP_REG_28__SCAN_IN), .ZN(n15326) );
  OAI21_X1 U15622 ( .B1(n15228), .B2(n12415), .A(n15326), .ZN(n12416) );
  NAND2_X1 U15623 ( .A1(n12418), .A2(n12417), .ZN(n12419) );
  NOR2_X1 U15624 ( .A1(n12420), .A2(n12419), .ZN(n12421) );
  NAND2_X1 U15625 ( .A1(n15934), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15796) );
  AND2_X1 U15626 ( .A1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15895) );
  INV_X1 U15627 ( .A(n15895), .ZN(n12485) );
  INV_X1 U15628 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n12425) );
  AOI21_X1 U15629 ( .B1(n15763), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n12423) );
  NOR2_X2 U15630 ( .A1(n12968), .A2(n12423), .ZN(n12794) );
  NAND2_X1 U15631 ( .A1(n12794), .A2(n16577), .ZN(n12505) );
  XNOR2_X1 U15632 ( .A(n12469), .B(n12424), .ZN(n12426) );
  INV_X1 U15633 ( .A(n12426), .ZN(n15495) );
  NAND3_X1 U15634 ( .A1(n15495), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n12808), .ZN(n12974) );
  NAND2_X1 U15635 ( .A1(n12974), .A2(n12800), .ZN(n12482) );
  NOR2_X1 U15636 ( .A1(n16023), .A2(n12427), .ZN(n12428) );
  INV_X1 U15637 ( .A(n12430), .ZN(n12431) );
  NAND2_X1 U15638 ( .A1(n9899), .A2(n12431), .ZN(n12441) );
  NAND2_X1 U15639 ( .A1(n15595), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12434) );
  NAND4_X1 U15640 ( .A1(n12435), .A2(n12434), .A3(n12433), .A4(n12432), .ZN(
        n12439) );
  AND4_X1 U15641 ( .A1(n15840), .A2(n12436), .A3(n15850), .A4(n16038), .ZN(
        n12437) );
  NAND2_X1 U15642 ( .A1(n15830), .A2(n12437), .ZN(n12438) );
  AOI21_X1 U15643 ( .B1(n12439), .B2(n12808), .A(n12438), .ZN(n12440) );
  NAND2_X1 U15644 ( .A1(n12444), .A2(n10185), .ZN(n12445) );
  NAND2_X1 U15645 ( .A1(n12449), .A2(n12445), .ZN(n15575) );
  OR2_X1 U15646 ( .A1(n15575), .A2(n11254), .ZN(n12446) );
  NAND2_X1 U15647 ( .A1(n12446), .A2(n15938), .ZN(n15951) );
  OR2_X1 U15648 ( .A1(n11254), .A2(n15938), .ZN(n12447) );
  OR2_X1 U15649 ( .A1(n15575), .A2(n12447), .ZN(n15950) );
  NAND2_X1 U15650 ( .A1(n12449), .A2(n12448), .ZN(n12450) );
  AND2_X1 U15651 ( .A1(n15536), .A2(n12450), .ZN(n15558) );
  NAND2_X1 U15652 ( .A1(n15558), .A2(n12808), .ZN(n12451) );
  NAND2_X1 U15653 ( .A1(n15935), .A2(n15936), .ZN(n12453) );
  NAND3_X1 U15654 ( .A1(n15558), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        n12808), .ZN(n12452) );
  NAND2_X1 U15655 ( .A1(n12453), .A2(n12452), .ZN(n15794) );
  NAND2_X1 U15656 ( .A1(n12460), .A2(n12808), .ZN(n12454) );
  NAND2_X1 U15657 ( .A1(n12454), .A2(n15922), .ZN(n15792) );
  NAND2_X1 U15658 ( .A1(n15794), .A2(n15792), .ZN(n12456) );
  INV_X1 U15659 ( .A(n12454), .ZN(n12455) );
  NAND2_X1 U15660 ( .A1(n12455), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15793) );
  NOR2_X1 U15661 ( .A1(n12457), .A2(n15653), .ZN(n12458) );
  NAND2_X1 U15662 ( .A1(n10543), .A2(n12458), .ZN(n12459) );
  AND2_X1 U15663 ( .A1(n12460), .A2(n12459), .ZN(n12461) );
  NAND2_X1 U15664 ( .A1(n12462), .A2(n12461), .ZN(n15530) );
  INV_X1 U15665 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15912) );
  NAND2_X1 U15666 ( .A1(n12478), .A2(n15912), .ZN(n15780) );
  AND3_X1 U15667 ( .A1(n10543), .A2(P2_EBX_REG_26__SCAN_IN), .A3(n12462), .ZN(
        n12463) );
  NOR2_X1 U15668 ( .A1(n12804), .A2(n12463), .ZN(n16450) );
  INV_X1 U15669 ( .A(n16450), .ZN(n12464) );
  NOR2_X1 U15670 ( .A1(n12464), .A2(n11254), .ZN(n12465) );
  NAND3_X1 U15671 ( .A1(n16450), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        n12808), .ZN(n12479) );
  OAI21_X1 U15672 ( .B1(n12465), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n12479), .ZN(n15773) );
  INV_X1 U15673 ( .A(n12466), .ZN(n12467) );
  NAND2_X1 U15674 ( .A1(n12467), .A2(n9889), .ZN(n12468) );
  NAND2_X1 U15675 ( .A1(n12470), .A2(n12468), .ZN(n13315) );
  AOI21_X1 U15676 ( .B1(n12471), .B2(n12470), .A(n12469), .ZN(n15515) );
  INV_X1 U15677 ( .A(n15515), .ZN(n12472) );
  INV_X1 U15678 ( .A(n15753), .ZN(n12475) );
  NAND2_X1 U15679 ( .A1(n12475), .A2(n12474), .ZN(n12476) );
  NAND2_X1 U15680 ( .A1(n12477), .A2(n12476), .ZN(n12481) );
  NAND2_X1 U15681 ( .A1(n15781), .A2(n12479), .ZN(n15749) );
  INV_X1 U15682 ( .A(n15749), .ZN(n12480) );
  XOR2_X1 U15683 ( .A(n12482), .B(n12801), .Z(n12795) );
  NAND2_X1 U15684 ( .A1(n12483), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15955) );
  AND2_X1 U15685 ( .A1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15937) );
  NAND2_X1 U15686 ( .A1(n15937), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n12484) );
  NOR2_X1 U15687 ( .A1(n15910), .A2(n12485), .ZN(n12985) );
  NAND2_X1 U15688 ( .A1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n12985), .ZN(
        n15877) );
  XNOR2_X1 U15689 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .B(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n12501) );
  NAND2_X1 U15690 ( .A1(n12486), .A2(n12487), .ZN(n12488) );
  NAND2_X1 U15691 ( .A1(n12489), .A2(n12488), .ZN(n15630) );
  INV_X1 U15692 ( .A(n15630), .ZN(n12494) );
  NOR2_X1 U15693 ( .A1(n15510), .A2(n12490), .ZN(n12491) );
  NAND2_X1 U15694 ( .A1(n19170), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n12789) );
  OAI21_X1 U15695 ( .B1(n19327), .B2(n15697), .A(n12789), .ZN(n12493) );
  AOI21_X1 U15696 ( .B1(n12494), .B2(n19341), .A(n12493), .ZN(n12500) );
  OR2_X1 U15697 ( .A1(n19353), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12495) );
  NAND2_X1 U15698 ( .A1(n12496), .A2(n12495), .ZN(n15953) );
  OAI21_X1 U15699 ( .B1(n19353), .B2(n15937), .A(
        P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n12497) );
  INV_X1 U15700 ( .A(n15930), .ZN(n15914) );
  NAND2_X1 U15701 ( .A1(n15914), .A2(n15895), .ZN(n15886) );
  NAND2_X1 U15702 ( .A1(n15886), .A2(n15911), .ZN(n12498) );
  NAND2_X1 U15703 ( .A1(n12985), .A2(n15764), .ZN(n15883) );
  NAND2_X1 U15704 ( .A1(n12498), .A2(n15883), .ZN(n15874) );
  NAND2_X1 U15705 ( .A1(n15874), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12499) );
  OAI211_X1 U15706 ( .C1(n15877), .C2(n12501), .A(n12500), .B(n12499), .ZN(
        n12502) );
  NAND2_X1 U15707 ( .A1(n12505), .A2(n12504), .ZN(P2_U3017) );
  INV_X2 U15708 ( .A(n17340), .ZN(n17385) );
  INV_X1 U15709 ( .A(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n17277) );
  AOI22_X1 U15710 ( .A1(n17379), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n17343), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12512) );
  AOI22_X1 U15711 ( .A1(n17357), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n13120), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12511) );
  OAI211_X1 U15712 ( .C1(n13050), .C2(n17277), .A(n12512), .B(n12511), .ZN(
        n12522) );
  AOI22_X1 U15713 ( .A1(n17378), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n17245), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12520) );
  AOI22_X1 U15714 ( .A1(n12552), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n17365), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12519) );
  NAND2_X4 U15715 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n12515), .ZN(
        n17395) );
  AOI22_X1 U15716 ( .A1(n13080), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n17327), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12518) );
  NAND2_X1 U15717 ( .A1(n17344), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n12517) );
  NAND4_X1 U15718 ( .A1(n12520), .A2(n12519), .A3(n12518), .A4(n12517), .ZN(
        n12521) );
  AOI22_X1 U15719 ( .A1(n17378), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n17245), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12525) );
  OAI21_X1 U15720 ( .B1(n21308), .B2(n17283), .A(n12525), .ZN(n12535) );
  AOI22_X1 U15721 ( .A1(n13080), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n17357), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12533) );
  INV_X1 U15722 ( .A(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12526) );
  OAI22_X1 U15723 ( .A1(n17363), .A2(n17359), .B1(n9827), .B2(n12526), .ZN(
        n12531) );
  AOI22_X1 U15724 ( .A1(n17385), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n9829), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12529) );
  AOI22_X1 U15725 ( .A1(n17365), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_10__1__SCAN_IN), .B2(n17343), .ZN(n12528) );
  AOI22_X1 U15726 ( .A1(n17327), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n17361), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12527) );
  NAND3_X1 U15727 ( .A1(n12529), .A2(n12528), .A3(n12527), .ZN(n12530) );
  AOI211_X1 U15728 ( .C1(n13079), .C2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A(
        n12531), .B(n12530), .ZN(n12532) );
  OAI211_X1 U15729 ( .C1(n21090), .C2(n17252), .A(n12533), .B(n12532), .ZN(
        n12534) );
  AOI211_X4 U15730 ( .C1(n17379), .C2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A(
        n12535), .B(n12534), .ZN(n19012) );
  AOI22_X1 U15731 ( .A1(n13079), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n13089), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12536) );
  OAI21_X1 U15732 ( .B1(n13050), .B2(n17383), .A(n12536), .ZN(n12541) );
  INV_X1 U15733 ( .A(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n17394) );
  AOI22_X1 U15734 ( .A1(n17386), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n13064), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12539) );
  AOI22_X1 U15735 ( .A1(n17245), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n13120), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12538) );
  OAI211_X1 U15736 ( .C1(n17384), .C2(n17394), .A(n12539), .B(n12538), .ZN(
        n12540) );
  AOI211_X1 U15737 ( .C1(n17344), .C2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A(
        n12541), .B(n12540), .ZN(n12549) );
  INV_X1 U15738 ( .A(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n17381) );
  AOI22_X1 U15739 ( .A1(n17385), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17343), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12542) );
  OAI21_X1 U15740 ( .B1(n17283), .B2(n17381), .A(n12542), .ZN(n12547) );
  AOI22_X1 U15741 ( .A1(n17379), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17365), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12543) );
  AOI22_X1 U15742 ( .A1(n13089), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n13068), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12559) );
  INV_X1 U15743 ( .A(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12550) );
  OAI22_X1 U15744 ( .A1(n12551), .A2(n17217), .B1(n17384), .B2(n12550), .ZN(
        n12557) );
  AOI22_X1 U15745 ( .A1(n17379), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17245), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12555) );
  AOI22_X1 U15746 ( .A1(n12552), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17343), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12554) );
  AOI22_X1 U15747 ( .A1(n17344), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17361), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12553) );
  NAND3_X1 U15748 ( .A1(n12555), .A2(n12554), .A3(n12553), .ZN(n12556) );
  AOI211_X1 U15749 ( .C1(n13080), .C2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A(
        n12557), .B(n12556), .ZN(n12558) );
  OAI211_X1 U15750 ( .C1(n13051), .C2(n17308), .A(n12559), .B(n12558), .ZN(
        n12560) );
  INV_X1 U15751 ( .A(n12560), .ZN(n12566) );
  INV_X1 U15752 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17411) );
  AOI22_X1 U15753 ( .A1(n9829), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17365), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12562) );
  OAI21_X1 U15754 ( .B1(n17252), .B2(n17411), .A(n12562), .ZN(n12564) );
  AOI22_X1 U15755 ( .A1(n13080), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17327), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12572) );
  INV_X1 U15756 ( .A(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n17186) );
  AOI22_X1 U15757 ( .A1(n13120), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n17343), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12568) );
  AOI22_X1 U15758 ( .A1(n17245), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17365), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12567) );
  OAI211_X1 U15759 ( .C1(n12551), .C2(n17186), .A(n12568), .B(n12567), .ZN(
        n12571) );
  AOI22_X1 U15760 ( .A1(n17378), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n13064), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12570) );
  AOI22_X1 U15761 ( .A1(n17357), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n13068), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12569) );
  NAND2_X1 U15762 ( .A1(n18401), .A2(n17433), .ZN(n12592) );
  INV_X1 U15763 ( .A(n12592), .ZN(n18816) );
  INV_X1 U15764 ( .A(n12631), .ZN(n17340) );
  AOI22_X1 U15765 ( .A1(n9829), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17343), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12573) );
  OAI21_X1 U15766 ( .B1(n17340), .B2(n17211), .A(n12573), .ZN(n12581) );
  AOI22_X1 U15767 ( .A1(n17245), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n13080), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12580) );
  INV_X1 U15768 ( .A(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12682) );
  OAI22_X1 U15769 ( .A1(n17363), .A2(n12682), .B1(n9827), .B2(n21277), .ZN(
        n12578) );
  AOI22_X1 U15770 ( .A1(n13120), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n17365), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12576) );
  AOI22_X1 U15771 ( .A1(n12552), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17357), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12575) );
  AOI22_X1 U15772 ( .A1(n17327), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17361), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12574) );
  NAND3_X1 U15773 ( .A1(n12576), .A2(n12575), .A3(n12574), .ZN(n12577) );
  AOI211_X1 U15774 ( .C1(n13079), .C2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A(
        n12578), .B(n12577), .ZN(n12579) );
  AOI22_X1 U15775 ( .A1(n13080), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n13079), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12591) );
  INV_X1 U15776 ( .A(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n17353) );
  AOI22_X1 U15777 ( .A1(n13120), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n13064), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12583) );
  AOI22_X1 U15778 ( .A1(n17379), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17343), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12582) );
  OAI211_X1 U15779 ( .C1(n17384), .C2(n17353), .A(n12583), .B(n12582), .ZN(
        n12589) );
  AOI22_X1 U15780 ( .A1(n12552), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17378), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12587) );
  AOI22_X1 U15781 ( .A1(n17245), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n17386), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12586) );
  AOI22_X1 U15782 ( .A1(n17385), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17365), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12585) );
  NAND2_X1 U15783 ( .A1(n13089), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(
        n12584) );
  NAND4_X1 U15784 ( .A1(n12587), .A2(n12586), .A3(n12585), .A4(n12584), .ZN(
        n12588) );
  AOI211_X1 U15785 ( .C1(n17344), .C2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A(
        n12589), .B(n12588), .ZN(n12590) );
  NOR2_X1 U15786 ( .A1(n13176), .A2(n18393), .ZN(n13250) );
  NAND2_X1 U15787 ( .A1(n12592), .A2(n13198), .ZN(n13181) );
  INV_X1 U15788 ( .A(n13181), .ZN(n12593) );
  AOI22_X1 U15789 ( .A1(n13089), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n13064), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12603) );
  INV_X1 U15790 ( .A(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n17325) );
  AOI22_X1 U15791 ( .A1(n17379), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17365), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12595) );
  AOI22_X1 U15792 ( .A1(n13120), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n13068), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12594) );
  OAI211_X1 U15793 ( .C1(n17384), .C2(n17325), .A(n12595), .B(n12594), .ZN(
        n12601) );
  AOI22_X1 U15794 ( .A1(n12552), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17343), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12599) );
  AOI22_X1 U15795 ( .A1(n17378), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17386), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12598) );
  AOI22_X1 U15796 ( .A1(n13080), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n13079), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12597) );
  NAND2_X1 U15797 ( .A1(n17361), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n12596) );
  NAND4_X1 U15798 ( .A1(n12599), .A2(n12598), .A3(n12597), .A4(n12596), .ZN(
        n12600) );
  NAND2_X1 U15799 ( .A1(n18397), .A2(n18413), .ZN(n13195) );
  NOR2_X1 U15800 ( .A1(n13191), .A2(n13190), .ZN(n12604) );
  OR2_X1 U15801 ( .A1(n12609), .A2(n12610), .ZN(n12605) );
  OAI21_X1 U15802 ( .B1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n18982), .A(
        n12605), .ZN(n12606) );
  OAI22_X1 U15803 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18847), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n12606), .ZN(n12611) );
  NOR2_X1 U15804 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18847), .ZN(
        n12607) );
  NAND2_X1 U15805 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n12606), .ZN(
        n12612) );
  AOI22_X1 U15806 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n12611), .B1(
        n12607), .B2(n12612), .ZN(n12616) );
  OAI21_X1 U15807 ( .B1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n18621), .A(
        n13190), .ZN(n13189) );
  NOR2_X1 U15808 ( .A1(n13191), .A2(n13189), .ZN(n12615) );
  OAI21_X1 U15809 ( .B1(n12610), .B2(n12609), .A(n12616), .ZN(n12608) );
  AOI21_X1 U15810 ( .B1(n12612), .B2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(
        n12611), .ZN(n12613) );
  INV_X1 U15811 ( .A(n13192), .ZN(n12614) );
  INV_X1 U15812 ( .A(n18808), .ZN(n16150) );
  NOR2_X1 U15813 ( .A1(n18393), .A2(n18397), .ZN(n18815) );
  NAND2_X1 U15814 ( .A1(n12617), .A2(n18815), .ZN(n13171) );
  NAND2_X1 U15815 ( .A1(n10005), .A2(n17547), .ZN(n12618) );
  INV_X1 U15816 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n16996) );
  NAND3_X1 U15817 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .ZN(n17410) );
  NAND2_X1 U15818 ( .A1(P3_EBX_REG_5__SCAN_IN), .A2(n17413), .ZN(n17404) );
  NAND2_X1 U15819 ( .A1(n17403), .A2(P3_EBX_REG_8__SCAN_IN), .ZN(n17374) );
  NAND2_X1 U15820 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n13981), .ZN(n17257) );
  NAND2_X1 U15821 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n17271), .ZN(n17239) );
  NAND2_X1 U15822 ( .A1(P3_EBX_REG_23__SCAN_IN), .A2(n17179), .ZN(n17175) );
  INV_X1 U15823 ( .A(P3_EBX_REG_28__SCAN_IN), .ZN(n17121) );
  NOR2_X1 U15824 ( .A1(n17426), .A2(n17160), .ZN(n17161) );
  INV_X1 U15825 ( .A(n9895), .ZN(n17169) );
  NAND2_X1 U15826 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(n17169), .ZN(n12694) );
  AOI22_X1 U15827 ( .A1(n17385), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n13064), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12620) );
  OAI21_X1 U15828 ( .B1(n17306), .B2(n21208), .A(n12620), .ZN(n12629) );
  INV_X1 U15829 ( .A(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n17324) );
  AOI22_X1 U15830 ( .A1(n13080), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n17386), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12627) );
  INV_X1 U15831 ( .A(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n13058) );
  OAI22_X1 U15832 ( .A1(n12551), .A2(n21140), .B1(n9827), .B2(n13058), .ZN(
        n12625) );
  AOI22_X1 U15833 ( .A1(n12552), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n13120), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12623) );
  AOI22_X1 U15834 ( .A1(n17378), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17343), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12622) );
  AOI22_X1 U15835 ( .A1(n17344), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17327), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12621) );
  NAND3_X1 U15836 ( .A1(n12623), .A2(n12622), .A3(n12621), .ZN(n12624) );
  AOI211_X1 U15837 ( .C1(n17361), .C2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A(
        n12625), .B(n12624), .ZN(n12626) );
  OAI211_X1 U15838 ( .C1(n12537), .C2(n17324), .A(n12627), .B(n12626), .ZN(
        n12628) );
  AOI211_X1 U15839 ( .C1(n17379), .C2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A(
        n12629), .B(n12628), .ZN(n17167) );
  AOI22_X1 U15840 ( .A1(n17378), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n17245), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12630) );
  OAI21_X1 U15841 ( .B1(n17283), .B2(n21090), .A(n12630), .ZN(n12640) );
  AOI22_X1 U15842 ( .A1(n13080), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_4__1__SCAN_IN), .B2(n13120), .ZN(n12638) );
  INV_X1 U15843 ( .A(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n13091) );
  OAI22_X1 U15844 ( .A1(n13091), .A2(n17363), .B1(n17359), .B2(n9827), .ZN(
        n12636) );
  AOI22_X1 U15845 ( .A1(n17386), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_14__1__SCAN_IN), .B2(n17343), .ZN(n12634) );
  AOI22_X1 U15846 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n17365), .B1(
        n13064), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12633) );
  AOI22_X1 U15847 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n17361), .B1(
        n17327), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12632) );
  NAND3_X1 U15848 ( .A1(n12634), .A2(n12633), .A3(n12632), .ZN(n12635) );
  AOI211_X1 U15849 ( .C1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .C2(n13079), .A(
        n12636), .B(n12635), .ZN(n12637) );
  OAI211_X1 U15850 ( .C1(n21308), .C2(n17340), .A(n12638), .B(n12637), .ZN(
        n12639) );
  AOI211_X1 U15851 ( .C1(n17379), .C2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A(
        n12640), .B(n12639), .ZN(n17176) );
  INV_X1 U15852 ( .A(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n13123) );
  AOI22_X1 U15853 ( .A1(n17357), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n13089), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12650) );
  AOI22_X1 U15854 ( .A1(n13120), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17365), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12641) );
  OAI21_X1 U15855 ( .B1(n13051), .B2(n17394), .A(n12641), .ZN(n12648) );
  AOI22_X1 U15856 ( .A1(n13079), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n17361), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12646) );
  AOI22_X1 U15857 ( .A1(n12552), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n17343), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12643) );
  AOI22_X1 U15858 ( .A1(n17379), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n13068), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12642) );
  OAI211_X1 U15859 ( .C1(n17363), .C2(n13127), .A(n12643), .B(n12642), .ZN(
        n12644) );
  AOI21_X1 U15860 ( .B1(n17327), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A(
        n12644), .ZN(n12645) );
  OAI211_X1 U15861 ( .C1(n17395), .C2(n17383), .A(n12646), .B(n12645), .ZN(
        n12647) );
  AOI211_X1 U15862 ( .C1(n17245), .C2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A(
        n12648), .B(n12647), .ZN(n12649) );
  OAI211_X1 U15863 ( .C1(n12561), .C2(n13123), .A(n12650), .B(n12649), .ZN(
        n17181) );
  AOI22_X1 U15864 ( .A1(n17245), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17365), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12661) );
  AOI22_X1 U15865 ( .A1(n17379), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n17386), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12660) );
  AOI22_X1 U15866 ( .A1(n17344), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n17327), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12659) );
  INV_X1 U15867 ( .A(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n17144) );
  OAI22_X1 U15868 ( .A1(n17395), .A2(n17401), .B1(n17252), .B2(n17144), .ZN(
        n12657) );
  AOI22_X1 U15869 ( .A1(n17385), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n17343), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12655) );
  AOI22_X1 U15870 ( .A1(n12552), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n13064), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12654) );
  AOI22_X1 U15871 ( .A1(n13089), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n17361), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12653) );
  NAND2_X1 U15872 ( .A1(n13079), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n12652) );
  NAND4_X1 U15873 ( .A1(n12655), .A2(n12654), .A3(n12653), .A4(n12652), .ZN(
        n12656) );
  AOI211_X1 U15874 ( .C1(n17378), .C2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A(
        n12657), .B(n12656), .ZN(n12658) );
  NAND4_X1 U15875 ( .A1(n12661), .A2(n12660), .A3(n12659), .A4(n12658), .ZN(
        n17182) );
  NAND2_X1 U15876 ( .A1(n17181), .A2(n17182), .ZN(n17180) );
  NOR2_X1 U15877 ( .A1(n17176), .A2(n17180), .ZN(n17172) );
  AOI22_X1 U15878 ( .A1(n13079), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n17361), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12671) );
  INV_X1 U15879 ( .A(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n17341) );
  INV_X2 U15880 ( .A(n9884), .ZN(n17343) );
  AOI22_X1 U15881 ( .A1(n17357), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17343), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12663) );
  AOI22_X1 U15882 ( .A1(n17245), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n13064), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12662) );
  OAI211_X1 U15883 ( .C1(n17384), .C2(n17341), .A(n12663), .B(n12662), .ZN(
        n12669) );
  AOI22_X1 U15884 ( .A1(n12552), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n17379), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12667) );
  AOI22_X1 U15885 ( .A1(n17378), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n13068), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12666) );
  AOI22_X1 U15886 ( .A1(n13120), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n17365), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12665) );
  NAND2_X1 U15887 ( .A1(n13089), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n12664) );
  NAND4_X1 U15888 ( .A1(n12667), .A2(n12666), .A3(n12665), .A4(n12664), .ZN(
        n12668) );
  AOI211_X1 U15889 ( .C1(n17344), .C2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A(
        n12669), .B(n12668), .ZN(n12670) );
  OAI211_X1 U15890 ( .C1(n17395), .C2(n21306), .A(n12671), .B(n12670), .ZN(
        n17171) );
  NAND2_X1 U15891 ( .A1(n17172), .A2(n17171), .ZN(n17170) );
  NOR2_X1 U15892 ( .A1(n17167), .A2(n17170), .ZN(n17165) );
  AOI22_X1 U15893 ( .A1(n13120), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n13089), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12681) );
  INV_X1 U15894 ( .A(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n17305) );
  AOI22_X1 U15895 ( .A1(n17378), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n17245), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12673) );
  AOI22_X1 U15896 ( .A1(n17365), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17343), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12672) );
  OAI211_X1 U15897 ( .C1(n13050), .C2(n17305), .A(n12673), .B(n12672), .ZN(
        n12679) );
  AOI22_X1 U15898 ( .A1(n12552), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n13068), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12677) );
  AOI22_X1 U15899 ( .A1(n17357), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n13064), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12676) );
  AOI22_X1 U15900 ( .A1(n13080), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n17327), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12675) );
  NAND2_X1 U15901 ( .A1(n13079), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n12674) );
  NAND4_X1 U15902 ( .A1(n12677), .A2(n12676), .A3(n12675), .A4(n12674), .ZN(
        n12678) );
  AOI211_X1 U15903 ( .C1(n17344), .C2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A(
        n12679), .B(n12678), .ZN(n12680) );
  OAI211_X1 U15904 ( .C1(n17360), .C2(n17308), .A(n12681), .B(n12680), .ZN(
        n17164) );
  NAND2_X1 U15905 ( .A1(n17165), .A2(n17164), .ZN(n17163) );
  AOI22_X1 U15906 ( .A1(n9829), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n17365), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12692) );
  AOI22_X1 U15907 ( .A1(n17378), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n13068), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12691) );
  OAI22_X1 U15908 ( .A1(n9827), .A2(n12682), .B1(n13050), .B2(n21277), .ZN(
        n12689) );
  INV_X1 U15909 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n17407) );
  AOI22_X1 U15910 ( .A1(n13080), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n13120), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12687) );
  INV_X1 U15911 ( .A(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n17200) );
  AOI22_X1 U15912 ( .A1(n17245), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17386), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12684) );
  AOI22_X1 U15913 ( .A1(n17379), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17343), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12683) );
  OAI211_X1 U15914 ( .C1(n17363), .C2(n17200), .A(n12684), .B(n12683), .ZN(
        n12685) );
  AOI21_X1 U15915 ( .B1(n13079), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A(
        n12685), .ZN(n12686) );
  OAI211_X1 U15916 ( .C1(n17283), .C2(n17407), .A(n12687), .B(n12686), .ZN(
        n12688) );
  AOI211_X1 U15917 ( .C1(n17327), .C2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A(
        n12689), .B(n12688), .ZN(n12690) );
  NAND3_X1 U15918 ( .A1(n12692), .A2(n12691), .A3(n12690), .ZN(n17156) );
  XNOR2_X1 U15919 ( .A(n17163), .B(n17156), .ZN(n17445) );
  NAND2_X1 U15920 ( .A1(n17426), .A2(n17445), .ZN(n12693) );
  AOI21_X1 U15921 ( .B1(n17161), .B2(P3_EBX_REG_28__SCAN_IN), .A(n12695), .ZN(
        n12696) );
  INV_X1 U15922 ( .A(n12696), .ZN(P3_U2675) );
  INV_X1 U15923 ( .A(n12697), .ZN(n12698) );
  INV_X1 U15924 ( .A(n12699), .ZN(n12700) );
  INV_X1 U15925 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n14824) );
  NAND2_X1 U15926 ( .A1(n12700), .A2(n14824), .ZN(n12701) );
  NAND2_X1 U15927 ( .A1(n12845), .A2(n12701), .ZN(n15132) );
  AOI22_X1 U15928 ( .A1(n9817), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12732), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12706) );
  AOI22_X1 U15929 ( .A1(n9851), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12702), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12705) );
  AOI22_X1 U15930 ( .A1(n9838), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n11622), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12704) );
  AOI22_X1 U15931 ( .A1(n12724), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12185), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12703) );
  NAND4_X1 U15932 ( .A1(n12706), .A2(n12705), .A3(n12704), .A4(n12703), .ZN(
        n12712) );
  AOI22_X1 U15933 ( .A1(n12038), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12286), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12710) );
  AOI22_X1 U15934 ( .A1(n12729), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11612), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12709) );
  AOI22_X1 U15935 ( .A1(n9852), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n12250), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12708) );
  AOI22_X1 U15936 ( .A1(n12731), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n10016), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12707) );
  NAND4_X1 U15937 ( .A1(n12710), .A2(n12709), .A3(n12708), .A4(n12707), .ZN(
        n12711) );
  NOR2_X1 U15938 ( .A1(n12712), .A2(n12711), .ZN(n12721) );
  NAND2_X1 U15939 ( .A1(n12714), .A2(n12713), .ZN(n12720) );
  XNOR2_X1 U15940 ( .A(n12721), .B(n12720), .ZN(n12718) );
  AOI21_X1 U15941 ( .B1(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n20999), .A(
        n12847), .ZN(n12716) );
  NAND2_X1 U15942 ( .A1(n12748), .A2(P1_EAX_REG_29__SCAN_IN), .ZN(n12715) );
  OAI211_X1 U15943 ( .C1(n12718), .C2(n12717), .A(n12716), .B(n12715), .ZN(
        n12719) );
  OAI21_X1 U15944 ( .B1(n15132), .B2(n12742), .A(n12719), .ZN(n14822) );
  XNOR2_X1 U15945 ( .A(n12845), .B(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15122) );
  NOR2_X1 U15946 ( .A1(n12721), .A2(n12720), .ZN(n12740) );
  AOI22_X1 U15947 ( .A1(n9838), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n12286), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12728) );
  AOI22_X1 U15948 ( .A1(n9852), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n12722), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12727) );
  AOI22_X1 U15949 ( .A1(n12356), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n10016), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12726) );
  AOI22_X1 U15950 ( .A1(n9849), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11716), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12725) );
  NAND4_X1 U15951 ( .A1(n12728), .A2(n12727), .A3(n12726), .A4(n12725), .ZN(
        n12738) );
  AOI22_X1 U15952 ( .A1(n9817), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12729), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12736) );
  AOI22_X1 U15953 ( .A1(n12038), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11612), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12735) );
  AOI22_X1 U15954 ( .A1(n12732), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12731), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12734) );
  AOI22_X1 U15955 ( .A1(n9850), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n12250), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12733) );
  NAND4_X1 U15956 ( .A1(n12736), .A2(n12735), .A3(n12734), .A4(n12733), .ZN(
        n12737) );
  NOR2_X1 U15957 ( .A1(n12738), .A2(n12737), .ZN(n12739) );
  XNOR2_X1 U15958 ( .A(n12740), .B(n12739), .ZN(n12745) );
  INV_X1 U15959 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n13022) );
  NAND2_X1 U15960 ( .A1(n20999), .A2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12741) );
  OAI211_X1 U15961 ( .C1(n12005), .C2(n13022), .A(n12742), .B(n12741), .ZN(
        n12743) );
  AOI21_X1 U15962 ( .B1(n12745), .B2(n12744), .A(n12743), .ZN(n12746) );
  AOI22_X1 U15963 ( .A1(n12748), .A2(P1_EAX_REG_31__SCAN_IN), .B1(n12747), 
        .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n12749) );
  INV_X1 U15964 ( .A(n12749), .ZN(n12750) );
  INV_X1 U15965 ( .A(n12753), .ZN(n12754) );
  INV_X1 U15966 ( .A(n12758), .ZN(n13758) );
  OR4_X1 U15967 ( .A1(n12762), .A2(n12761), .A3(n12760), .A4(n12759), .ZN(
        n13756) );
  NAND2_X1 U15968 ( .A1(n13758), .A2(n13756), .ZN(n16192) );
  NAND2_X1 U15969 ( .A1(n12763), .A2(n21010), .ZN(n12765) );
  NAND2_X1 U15970 ( .A1(n13791), .A2(n12763), .ZN(n13792) );
  INV_X1 U15971 ( .A(n11979), .ZN(n20349) );
  NAND3_X1 U15972 ( .A1(n11679), .A2(n20349), .A3(n12766), .ZN(n13544) );
  NOR2_X1 U15973 ( .A1(n13514), .A2(n13544), .ZN(n12767) );
  AND2_X1 U15974 ( .A1(n15090), .A2(n20349), .ZN(n12769) );
  NAND2_X1 U15975 ( .A1(n13010), .A2(n12769), .ZN(n12784) );
  NOR4_X1 U15976 ( .A1(P1_ADDRESS_REG_15__SCAN_IN), .A2(
        P1_ADDRESS_REG_14__SCAN_IN), .A3(P1_ADDRESS_REG_13__SCAN_IN), .A4(
        P1_ADDRESS_REG_12__SCAN_IN), .ZN(n12773) );
  NOR4_X1 U15977 ( .A1(P1_ADDRESS_REG_19__SCAN_IN), .A2(
        P1_ADDRESS_REG_18__SCAN_IN), .A3(P1_ADDRESS_REG_17__SCAN_IN), .A4(
        P1_ADDRESS_REG_16__SCAN_IN), .ZN(n12772) );
  NOR4_X1 U15978 ( .A1(P1_ADDRESS_REG_7__SCAN_IN), .A2(
        P1_ADDRESS_REG_6__SCAN_IN), .A3(P1_ADDRESS_REG_5__SCAN_IN), .A4(
        P1_ADDRESS_REG_4__SCAN_IN), .ZN(n12771) );
  NOR4_X1 U15979 ( .A1(P1_ADDRESS_REG_11__SCAN_IN), .A2(
        P1_ADDRESS_REG_10__SCAN_IN), .A3(P1_ADDRESS_REG_9__SCAN_IN), .A4(
        P1_ADDRESS_REG_8__SCAN_IN), .ZN(n12770) );
  AND4_X1 U15980 ( .A1(n12773), .A2(n12772), .A3(n12771), .A4(n12770), .ZN(
        n12778) );
  NOR4_X1 U15981 ( .A1(P1_ADDRESS_REG_1__SCAN_IN), .A2(
        P1_ADDRESS_REG_0__SCAN_IN), .A3(P1_ADDRESS_REG_3__SCAN_IN), .A4(
        P1_ADDRESS_REG_28__SCAN_IN), .ZN(n12776) );
  NOR4_X1 U15982 ( .A1(P1_ADDRESS_REG_23__SCAN_IN), .A2(
        P1_ADDRESS_REG_22__SCAN_IN), .A3(P1_ADDRESS_REG_21__SCAN_IN), .A4(
        P1_ADDRESS_REG_20__SCAN_IN), .ZN(n12775) );
  NOR4_X1 U15983 ( .A1(P1_ADDRESS_REG_27__SCAN_IN), .A2(
        P1_ADDRESS_REG_26__SCAN_IN), .A3(P1_ADDRESS_REG_25__SCAN_IN), .A4(
        P1_ADDRESS_REG_24__SCAN_IN), .ZN(n12774) );
  AND4_X1 U15984 ( .A1(n12776), .A2(n12775), .A3(n12774), .A4(n20931), .ZN(
        n12777) );
  NAND2_X1 U15985 ( .A1(n12778), .A2(n12777), .ZN(n12779) );
  INV_X1 U15986 ( .A(n20303), .ZN(n20305) );
  INV_X1 U15987 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n20347) );
  NOR2_X1 U15988 ( .A1(n16299), .A2(n20347), .ZN(n12782) );
  AOI22_X1 U15989 ( .A1(n16295), .A2(DATAI_31_), .B1(P1_EAX_REG_31__SCAN_IN), 
        .B2(n16293), .ZN(n12780) );
  INV_X1 U15990 ( .A(n12780), .ZN(n12781) );
  NOR2_X1 U15991 ( .A1(n12782), .A2(n12781), .ZN(n12783) );
  NAND2_X1 U15992 ( .A1(n12784), .A2(n12783), .ZN(P1_U2873) );
  AND2_X1 U15993 ( .A1(n10657), .A2(n13386), .ZN(n12785) );
  NOR2_X1 U15994 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n20005) );
  INV_X1 U15995 ( .A(n20005), .ZN(n19038) );
  NAND2_X1 U15996 ( .A1(n20002), .A2(n19038), .ZN(n20039) );
  NAND2_X1 U15997 ( .A1(n20039), .A2(n14298), .ZN(n12787) );
  AND2_X1 U15998 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n20024) );
  NAND2_X1 U15999 ( .A1(n20061), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n12788) );
  NAND2_X1 U16000 ( .A1(n13350), .A2(n12788), .ZN(n13346) );
  OAI21_X1 U16001 ( .B1(n16559), .B2(n12790), .A(n12789), .ZN(n12791) );
  AOI21_X1 U16002 ( .B1(n16550), .B2(n15500), .A(n12791), .ZN(n12792) );
  OAI21_X1 U16003 ( .B1(n15630), .B2(n16545), .A(n12792), .ZN(n12793) );
  AOI21_X1 U16004 ( .B1(n12794), .B2(n16539), .A(n12793), .ZN(n12796) );
  NAND2_X1 U16005 ( .A1(n12796), .A2(n10380), .ZN(P2_U2985) );
  INV_X1 U16006 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n12797) );
  INV_X1 U16007 ( .A(n12844), .ZN(n12799) );
  NAND2_X1 U16008 ( .A1(n12799), .A2(n16577), .ZN(n12833) );
  AOI21_X1 U16009 ( .B1(n12803), .B2(n12808), .A(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n12978) );
  INV_X1 U16010 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n12983) );
  NOR2_X1 U16011 ( .A1(n11254), .A2(n12983), .ZN(n12802) );
  NAND2_X1 U16012 ( .A1(n12803), .A2(n12802), .ZN(n12976) );
  INV_X1 U16013 ( .A(n12804), .ZN(n12807) );
  NOR2_X1 U16014 ( .A1(n12805), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n12806) );
  MUX2_X1 U16015 ( .A(n12807), .B(n12806), .S(n10543), .Z(n15491) );
  NAND2_X1 U16016 ( .A1(n15491), .A2(n12808), .ZN(n12809) );
  XNOR2_X1 U16017 ( .A(n12809), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n12810) );
  NOR2_X1 U16018 ( .A1(n12839), .A2(n19363), .ZN(n12831) );
  AOI22_X1 U16019 ( .A1(n12811), .A2(P2_REIP_REG_31__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n12814) );
  NAND2_X1 U16020 ( .A1(n12812), .A2(P2_EBX_REG_31__SCAN_IN), .ZN(n12813) );
  OAI211_X1 U16021 ( .C1(n12815), .C2(n12797), .A(n12814), .B(n12813), .ZN(
        n12816) );
  NAND2_X1 U16022 ( .A1(n12818), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n12821) );
  AOI22_X1 U16023 ( .A1(n12819), .A2(P2_EAX_REG_31__SCAN_IN), .B1(n10690), 
        .B2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n12820) );
  AND2_X1 U16024 ( .A1(n12821), .A2(n12820), .ZN(n12822) );
  AND3_X1 U16025 ( .A1(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n12984) );
  NAND2_X1 U16026 ( .A1(n15895), .A2(n12984), .ZN(n12824) );
  OAI21_X1 U16027 ( .B1(n15930), .B2(n12824), .A(n15911), .ZN(n12986) );
  OAI21_X1 U16028 ( .B1(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n19353), .A(
        n12986), .ZN(n12825) );
  NAND2_X1 U16029 ( .A1(n12825), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n12826) );
  NAND2_X1 U16030 ( .A1(n19170), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n12835) );
  NAND2_X1 U16031 ( .A1(n12826), .A2(n12835), .ZN(n12827) );
  NAND2_X1 U16032 ( .A1(n12833), .A2(n12832), .ZN(P2_U3015) );
  INV_X1 U16033 ( .A(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n12837) );
  NAND2_X1 U16034 ( .A1(n16550), .A2(n12834), .ZN(n12836) );
  OAI211_X1 U16035 ( .C1(n12837), .C2(n16559), .A(n12836), .B(n12835), .ZN(
        n12838) );
  INV_X1 U16036 ( .A(n12839), .ZN(n12841) );
  OAI211_X1 U16037 ( .C1(n12844), .C2(n19319), .A(n12843), .B(n12842), .ZN(
        P2_U2983) );
  INV_X1 U16038 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n15124) );
  INV_X1 U16039 ( .A(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n12956) );
  NAND2_X1 U16040 ( .A1(n12847), .A2(n21002), .ZN(n13835) );
  NAND2_X1 U16041 ( .A1(n13010), .A2(n20131), .ZN(n12967) );
  BUF_X1 U16042 ( .A(n12848), .Z(n12934) );
  AOI22_X1 U16043 ( .A1(n13630), .A2(P1_EBX_REG_30__SCAN_IN), .B1(
        P1_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n16195), .ZN(n14808) );
  INV_X1 U16045 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n12850) );
  NAND2_X1 U16046 ( .A1(n12923), .A2(n12850), .ZN(n12854) );
  INV_X1 U16047 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n20286) );
  NAND2_X1 U16048 ( .A1(n9856), .A2(n20286), .ZN(n12852) );
  NAND2_X1 U16049 ( .A1(n13548), .A2(n12850), .ZN(n12851) );
  NAND3_X1 U16050 ( .A1(n12852), .A2(n12934), .A3(n12851), .ZN(n12853) );
  NAND2_X1 U16051 ( .A1(n9856), .A2(P1_EBX_REG_0__SCAN_IN), .ZN(n12856) );
  INV_X1 U16052 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n13633) );
  NAND2_X1 U16053 ( .A1(n12934), .A2(n13633), .ZN(n12855) );
  NAND2_X1 U16054 ( .A1(n12856), .A2(n12855), .ZN(n13631) );
  INV_X1 U16055 ( .A(n9856), .ZN(n12886) );
  INV_X1 U16056 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n13935) );
  MUX2_X1 U16057 ( .A(n12886), .B(n12923), .S(n13935), .Z(n12860) );
  NAND2_X1 U16058 ( .A1(n12886), .A2(n16195), .ZN(n12888) );
  NAND2_X1 U16059 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n16195), .ZN(
        n12858) );
  NAND2_X1 U16060 ( .A1(n12888), .A2(n12858), .ZN(n12859) );
  NOR2_X1 U16061 ( .A1(n12860), .A2(n12859), .ZN(n13753) );
  MUX2_X1 U16062 ( .A(n12927), .B(n12934), .S(P1_EBX_REG_3__SCAN_IN), .Z(
        n12861) );
  OAI21_X1 U16063 ( .B1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n13630), .A(
        n12861), .ZN(n13859) );
  INV_X1 U16064 ( .A(n12923), .ZN(n12932) );
  MUX2_X1 U16065 ( .A(n12932), .B(n9856), .S(P1_EBX_REG_4__SCAN_IN), .Z(n12864) );
  NAND2_X1 U16066 ( .A1(n16195), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12862) );
  AND2_X1 U16067 ( .A1(n12888), .A2(n12862), .ZN(n12863) );
  NAND2_X1 U16068 ( .A1(n12864), .A2(n12863), .ZN(n14044) );
  NAND2_X1 U16069 ( .A1(n12934), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12865) );
  OAI211_X1 U16070 ( .C1(n16195), .C2(P1_EBX_REG_5__SCAN_IN), .A(n9856), .B(
        n12865), .ZN(n12866) );
  OAI21_X1 U16071 ( .B1(n12927), .B2(P1_EBX_REG_5__SCAN_IN), .A(n12866), .ZN(
        n16422) );
  MUX2_X1 U16072 ( .A(n12923), .B(n12886), .S(P1_EBX_REG_6__SCAN_IN), .Z(
        n12869) );
  NAND2_X1 U16073 ( .A1(n16195), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12867) );
  NAND2_X1 U16074 ( .A1(n12888), .A2(n12867), .ZN(n12868) );
  NOR2_X1 U16075 ( .A1(n12869), .A2(n12868), .ZN(n14259) );
  NAND2_X1 U16076 ( .A1(n12934), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12870) );
  OAI211_X1 U16077 ( .C1(n16195), .C2(P1_EBX_REG_7__SCAN_IN), .A(n9856), .B(
        n12870), .ZN(n12871) );
  OAI21_X1 U16078 ( .B1(n12927), .B2(P1_EBX_REG_7__SCAN_IN), .A(n12871), .ZN(
        n16407) );
  MUX2_X1 U16079 ( .A(n12932), .B(n9856), .S(P1_EBX_REG_8__SCAN_IN), .Z(n12874) );
  NAND2_X1 U16080 ( .A1(n16195), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12872) );
  AND2_X1 U16081 ( .A1(n12888), .A2(n12872), .ZN(n12873) );
  NAND2_X1 U16082 ( .A1(n12874), .A2(n12873), .ZN(n14505) );
  INV_X1 U16083 ( .A(n12927), .ZN(n12875) );
  INV_X1 U16084 ( .A(P1_EBX_REG_9__SCAN_IN), .ZN(n20169) );
  NAND2_X1 U16085 ( .A1(n12875), .A2(n20169), .ZN(n12878) );
  NAND2_X1 U16086 ( .A1(n12934), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n12876) );
  OAI211_X1 U16087 ( .C1(n16195), .C2(P1_EBX_REG_9__SCAN_IN), .A(n9856), .B(
        n12876), .ZN(n12877) );
  AND2_X1 U16088 ( .A1(n12878), .A2(n12877), .ZN(n14504) );
  AND2_X1 U16089 ( .A1(n14505), .A2(n14504), .ZN(n12879) );
  INV_X1 U16090 ( .A(P1_EBX_REG_10__SCAN_IN), .ZN(n14463) );
  NAND2_X1 U16091 ( .A1(n12923), .A2(n14463), .ZN(n12883) );
  INV_X1 U16092 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15266) );
  NAND2_X1 U16093 ( .A1(n9856), .A2(n15266), .ZN(n12881) );
  NAND2_X1 U16094 ( .A1(n13548), .A2(n14463), .ZN(n12880) );
  NAND3_X1 U16095 ( .A1(n12881), .A2(n12934), .A3(n12880), .ZN(n12882) );
  MUX2_X1 U16096 ( .A(n12927), .B(n12934), .S(P1_EBX_REG_11__SCAN_IN), .Z(
        n12884) );
  OAI21_X1 U16097 ( .B1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n13630), .A(
        n12884), .ZN(n15041) );
  NOR2_X1 U16098 ( .A1(n15042), .A2(n15041), .ZN(n12885) );
  NAND2_X1 U16099 ( .A1(n15040), .A2(n12885), .ZN(n15044) );
  MUX2_X1 U16100 ( .A(n12923), .B(n12886), .S(P1_EBX_REG_12__SCAN_IN), .Z(
        n12890) );
  NAND2_X1 U16101 ( .A1(n16195), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n12887) );
  NAND2_X1 U16102 ( .A1(n12888), .A2(n12887), .ZN(n12889) );
  NOR2_X1 U16103 ( .A1(n12890), .A2(n12889), .ZN(n15037) );
  MUX2_X1 U16104 ( .A(n12927), .B(n12934), .S(P1_EBX_REG_13__SCAN_IN), .Z(
        n12891) );
  OAI21_X1 U16105 ( .B1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n13630), .A(
        n12891), .ZN(n14985) );
  INV_X1 U16106 ( .A(P1_EBX_REG_14__SCAN_IN), .ZN(n12893) );
  NAND2_X1 U16107 ( .A1(n12923), .A2(n12893), .ZN(n12897) );
  NAND2_X1 U16108 ( .A1(n9856), .A2(n12892), .ZN(n12895) );
  NAND2_X1 U16109 ( .A1(n13548), .A2(n12893), .ZN(n12894) );
  NAND3_X1 U16110 ( .A1(n12895), .A2(n12934), .A3(n12894), .ZN(n12896) );
  MUX2_X1 U16111 ( .A(n12927), .B(n12934), .S(P1_EBX_REG_15__SCAN_IN), .Z(
        n12898) );
  OAI21_X1 U16112 ( .B1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n13630), .A(
        n12898), .ZN(n15019) );
  NOR2_X1 U16113 ( .A1(n15029), .A2(n15019), .ZN(n12899) );
  INV_X1 U16114 ( .A(P1_EBX_REG_16__SCAN_IN), .ZN(n14970) );
  NAND2_X1 U16115 ( .A1(n12923), .A2(n14970), .ZN(n12903) );
  NAND2_X1 U16116 ( .A1(n9856), .A2(n16359), .ZN(n12901) );
  NAND2_X1 U16117 ( .A1(n13548), .A2(n14970), .ZN(n12900) );
  NAND3_X1 U16118 ( .A1(n12901), .A2(n12934), .A3(n12900), .ZN(n12902) );
  MUX2_X1 U16119 ( .A(n12927), .B(n12934), .S(P1_EBX_REG_17__SCAN_IN), .Z(
        n12904) );
  OAI21_X1 U16120 ( .B1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n13630), .A(
        n12904), .ZN(n14947) );
  NOR2_X1 U16121 ( .A1(n14965), .A2(n14947), .ZN(n12905) );
  INV_X1 U16122 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n15015) );
  NAND2_X1 U16123 ( .A1(n12923), .A2(n15015), .ZN(n12909) );
  NAND2_X1 U16124 ( .A1(n9856), .A2(n15433), .ZN(n12907) );
  NAND2_X1 U16125 ( .A1(n13548), .A2(n15015), .ZN(n12906) );
  NAND3_X1 U16126 ( .A1(n12907), .A2(n12934), .A3(n12906), .ZN(n12908) );
  AND2_X1 U16127 ( .A1(n12909), .A2(n12908), .ZN(n15013) );
  MUX2_X1 U16128 ( .A(n12927), .B(n12934), .S(P1_EBX_REG_19__SCAN_IN), .Z(
        n12910) );
  NAND2_X1 U16129 ( .A1(n10374), .A2(n12910), .ZN(n15007) );
  MUX2_X1 U16130 ( .A(n12932), .B(n9856), .S(P1_EBX_REG_20__SCAN_IN), .Z(
        n12912) );
  NAND2_X1 U16131 ( .A1(n16195), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12911) );
  NAND2_X1 U16132 ( .A1(n12912), .A2(n12911), .ZN(n14934) );
  NAND2_X1 U16133 ( .A1(n12934), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12913) );
  OAI211_X1 U16134 ( .C1(n16195), .C2(P1_EBX_REG_21__SCAN_IN), .A(n9856), .B(
        n12913), .ZN(n12914) );
  OAI21_X1 U16135 ( .B1(n12927), .B2(P1_EBX_REG_21__SCAN_IN), .A(n12914), .ZN(
        n14917) );
  INV_X1 U16136 ( .A(P1_EBX_REG_22__SCAN_IN), .ZN(n15001) );
  NAND2_X1 U16137 ( .A1(n12923), .A2(n15001), .ZN(n12917) );
  NAND2_X1 U16138 ( .A1(n9856), .A2(n15392), .ZN(n12915) );
  OAI211_X1 U16139 ( .C1(P1_EBX_REG_22__SCAN_IN), .C2(n16195), .A(n12915), .B(
        n12934), .ZN(n12916) );
  MUX2_X1 U16140 ( .A(n12927), .B(n12934), .S(P1_EBX_REG_23__SCAN_IN), .Z(
        n12918) );
  OAI21_X1 U16141 ( .B1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n13630), .A(
        n12918), .ZN(n14891) );
  NAND2_X1 U16142 ( .A1(n9856), .A2(n15362), .ZN(n12919) );
  OAI211_X1 U16143 ( .C1(P1_EBX_REG_24__SCAN_IN), .C2(n16195), .A(n12919), .B(
        n12934), .ZN(n12920) );
  OAI21_X1 U16144 ( .B1(n12932), .B2(P1_EBX_REG_24__SCAN_IN), .A(n12920), .ZN(
        n14876) );
  NAND2_X1 U16145 ( .A1(n14892), .A2(n14876), .ZN(n14878) );
  MUX2_X1 U16146 ( .A(n12927), .B(n12934), .S(P1_EBX_REG_25__SCAN_IN), .Z(
        n12921) );
  OAI21_X1 U16147 ( .B1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n13630), .A(
        n12921), .ZN(n14862) );
  INV_X1 U16148 ( .A(n12922), .ZN(n14861) );
  INV_X1 U16149 ( .A(P1_EBX_REG_26__SCAN_IN), .ZN(n14994) );
  NAND2_X1 U16150 ( .A1(n12923), .A2(n14994), .ZN(n12926) );
  INV_X1 U16151 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15348) );
  NAND2_X1 U16152 ( .A1(n9856), .A2(n15348), .ZN(n12924) );
  OAI211_X1 U16153 ( .C1(P1_EBX_REG_26__SCAN_IN), .C2(n16195), .A(n12924), .B(
        n12934), .ZN(n12925) );
  MUX2_X1 U16154 ( .A(n12927), .B(n12934), .S(P1_EBX_REG_27__SCAN_IN), .Z(
        n12928) );
  OAI21_X1 U16155 ( .B1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n13630), .A(
        n12928), .ZN(n14837) );
  NAND2_X1 U16156 ( .A1(n9856), .A2(n15327), .ZN(n12930) );
  OAI211_X1 U16157 ( .C1(P1_EBX_REG_28__SCAN_IN), .C2(n16195), .A(n12930), .B(
        n12848), .ZN(n12931) );
  OAI21_X1 U16158 ( .B1(n12932), .B2(P1_EBX_REG_28__SCAN_IN), .A(n12931), .ZN(
        n14520) );
  INV_X1 U16159 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n14992) );
  NAND2_X1 U16160 ( .A1(n13548), .A2(n14992), .ZN(n12935) );
  OR2_X1 U16161 ( .A1(n13630), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12933) );
  NAND2_X1 U16162 ( .A1(n12933), .A2(n12935), .ZN(n14806) );
  MUX2_X1 U16163 ( .A(n12935), .B(n14806), .S(n12934), .Z(n14817) );
  MUX2_X1 U16164 ( .A(n12934), .B(n14808), .S(n14819), .Z(n12937) );
  AOI22_X1 U16165 ( .A1(n13630), .A2(P1_EBX_REG_31__SCAN_IN), .B1(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n16195), .ZN(n12936) );
  NAND2_X1 U16166 ( .A1(n16194), .A2(n13768), .ZN(n13396) );
  NOR2_X1 U16167 ( .A1(n13840), .A2(n13775), .ZN(n12955) );
  NAND2_X1 U16168 ( .A1(n16201), .A2(P1_EBX_REG_31__SCAN_IN), .ZN(n12951) );
  AND2_X1 U16169 ( .A1(n21010), .A2(n21000), .ZN(n16203) );
  NOR2_X1 U16170 ( .A1(n12951), .A2(n16203), .ZN(n12939) );
  INV_X1 U16171 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n12940) );
  NAND2_X1 U16172 ( .A1(n12941), .A2(n12940), .ZN(n16223) );
  NAND2_X1 U16173 ( .A1(n11633), .A2(n16223), .ZN(n13759) );
  AND2_X1 U16174 ( .A1(n13759), .A2(n16203), .ZN(n12953) );
  NAND3_X1 U16175 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n16442), .A3(n20999), 
        .ZN(n16211) );
  OAI21_X1 U16176 ( .B1(n16211), .B2(n20310), .A(n13835), .ZN(n12942) );
  OR2_X1 U16177 ( .A1(n20296), .A2(n12942), .ZN(n12943) );
  AND2_X1 U16178 ( .A1(P1_REIP_REG_29__SCAN_IN), .A2(P1_REIP_REG_30__SCAN_IN), 
        .ZN(n12960) );
  INV_X1 U16179 ( .A(P1_REIP_REG_8__SCAN_IN), .ZN(n21260) );
  NAND4_X1 U16180 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(P1_REIP_REG_3__SCAN_IN), 
        .A3(P1_REIP_REG_1__SCAN_IN), .A4(P1_REIP_REG_2__SCAN_IN), .ZN(n20136)
         );
  NAND2_X1 U16181 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(P1_REIP_REG_5__SCAN_IN), 
        .ZN(n20112) );
  NOR2_X1 U16182 ( .A1(n20136), .A2(n20112), .ZN(n20118) );
  NAND2_X1 U16183 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(n20118), .ZN(n14393) );
  NOR2_X1 U16184 ( .A1(n21260), .A2(n14393), .ZN(n14461) );
  INV_X1 U16185 ( .A(P1_REIP_REG_12__SCAN_IN), .ZN(n20944) );
  NAND3_X1 U16186 ( .A1(P1_REIP_REG_11__SCAN_IN), .A2(P1_REIP_REG_10__SCAN_IN), 
        .A3(P1_REIP_REG_9__SCAN_IN), .ZN(n16278) );
  NOR2_X1 U16187 ( .A1(n20944), .A2(n16278), .ZN(n14955) );
  NAND2_X1 U16188 ( .A1(n14461), .A2(n14955), .ZN(n14935) );
  INV_X1 U16189 ( .A(P1_REIP_REG_17__SCAN_IN), .ZN(n20952) );
  NAND2_X1 U16190 ( .A1(P1_REIP_REG_16__SCAN_IN), .A2(P1_REIP_REG_15__SCAN_IN), 
        .ZN(n14967) );
  NOR2_X1 U16191 ( .A1(n20952), .A2(n14967), .ZN(n16238) );
  AND2_X1 U16192 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(P1_REIP_REG_13__SCAN_IN), 
        .ZN(n14956) );
  AND4_X1 U16193 ( .A1(P1_REIP_REG_19__SCAN_IN), .A2(P1_REIP_REG_20__SCAN_IN), 
        .A3(P1_REIP_REG_18__SCAN_IN), .A4(n14956), .ZN(n12944) );
  NAND2_X1 U16194 ( .A1(n16238), .A2(n12944), .ZN(n12945) );
  NOR2_X1 U16195 ( .A1(n14935), .A2(n12945), .ZN(n14906) );
  AND3_X1 U16196 ( .A1(P1_REIP_REG_23__SCAN_IN), .A2(P1_REIP_REG_21__SCAN_IN), 
        .A3(P1_REIP_REG_22__SCAN_IN), .ZN(n12946) );
  NAND2_X1 U16197 ( .A1(n14906), .A2(n12946), .ZN(n14880) );
  INV_X1 U16198 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n20965) );
  NOR2_X1 U16199 ( .A1(n14880), .A2(n20965), .ZN(n14866) );
  NAND2_X1 U16200 ( .A1(P1_REIP_REG_25__SCAN_IN), .A2(n14866), .ZN(n14848) );
  INV_X1 U16201 ( .A(n14848), .ZN(n12947) );
  AND2_X1 U16202 ( .A1(P1_REIP_REG_26__SCAN_IN), .A2(n12947), .ZN(n12957) );
  OR2_X1 U16203 ( .A1(n20151), .A2(n12957), .ZN(n12948) );
  NAND2_X1 U16204 ( .A1(n12948), .A2(n20117), .ZN(n14851) );
  INV_X1 U16205 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n20971) );
  NOR2_X1 U16206 ( .A1(n14851), .A2(n20971), .ZN(n14838) );
  NAND2_X1 U16207 ( .A1(n14838), .A2(P1_REIP_REG_28__SCAN_IN), .ZN(n12950) );
  INV_X1 U16208 ( .A(n14958), .ZN(n12949) );
  NAND2_X1 U16209 ( .A1(n12950), .A2(n12949), .ZN(n14828) );
  OAI21_X1 U16210 ( .B1(n14958), .B2(n12960), .A(n14828), .ZN(n14810) );
  INV_X1 U16211 ( .A(n12951), .ZN(n12952) );
  NOR2_X1 U16212 ( .A1(n12953), .A2(n12952), .ZN(n12954) );
  INV_X1 U16213 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n14989) );
  OAI22_X1 U16214 ( .A1(n20122), .A2(n14989), .B1(n12956), .B2(n20158), .ZN(
        n12963) );
  INV_X1 U16215 ( .A(n12957), .ZN(n12958) );
  NOR2_X1 U16216 ( .A1(n20151), .A2(n12958), .ZN(n14840) );
  AND2_X1 U16217 ( .A1(P1_REIP_REG_27__SCAN_IN), .A2(P1_REIP_REG_28__SCAN_IN), 
        .ZN(n12959) );
  NAND2_X1 U16218 ( .A1(n14840), .A2(n12959), .ZN(n14823) );
  INV_X1 U16219 ( .A(n12960), .ZN(n12961) );
  NOR3_X1 U16220 ( .A1(n14823), .A2(P1_REIP_REG_31__SCAN_IN), .A3(n12961), 
        .ZN(n12962) );
  AOI211_X1 U16221 ( .C1(n14810), .C2(P1_REIP_REG_31__SCAN_IN), .A(n12963), 
        .B(n12962), .ZN(n12964) );
  NAND2_X1 U16222 ( .A1(n12967), .A2(n12966), .ZN(P1_U2809) );
  XNOR2_X1 U16223 ( .A(n12968), .B(n12983), .ZN(n12996) );
  NAND2_X1 U16224 ( .A1(n19170), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n12987) );
  OAI21_X1 U16225 ( .B1(n16559), .B2(n12969), .A(n12987), .ZN(n12970) );
  AOI21_X1 U16226 ( .B1(n16550), .B2(n12971), .A(n12970), .ZN(n12972) );
  OAI21_X1 U16227 ( .B1(n14789), .B2(n16545), .A(n12972), .ZN(n12973) );
  AOI21_X1 U16228 ( .B1(n12996), .B2(n16539), .A(n12973), .ZN(n12982) );
  NAND2_X1 U16229 ( .A1(n12975), .A2(n12974), .ZN(n12980) );
  INV_X1 U16230 ( .A(n12976), .ZN(n12977) );
  NOR2_X1 U16231 ( .A1(n12978), .A2(n12977), .ZN(n12979) );
  XNOR2_X1 U16232 ( .A(n12980), .B(n12979), .ZN(n12997) );
  NAND2_X1 U16233 ( .A1(n12982), .A2(n12981), .ZN(P2_U2984) );
  NAND3_X1 U16234 ( .A1(n12985), .A2(n12984), .A3(n12983), .ZN(n12991) );
  INV_X1 U16235 ( .A(n12986), .ZN(n12989) );
  AOI21_X1 U16236 ( .B1(n12989), .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n12988), .ZN(n12990) );
  NAND2_X1 U16237 ( .A1(n12991), .A2(n12990), .ZN(n12992) );
  OAI21_X1 U16238 ( .B1(n14789), .B2(n19355), .A(n12994), .ZN(n12995) );
  AOI21_X1 U16239 ( .B1(n12996), .B2(n16577), .A(n12995), .ZN(n12999) );
  NAND2_X1 U16240 ( .A1(n12999), .A2(n12998), .ZN(P2_U3016) );
  NOR2_X1 U16241 ( .A1(n13001), .A2(n16302), .ZN(n15154) );
  INV_X1 U16242 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15339) );
  NAND2_X1 U16243 ( .A1(n15339), .A2(n15327), .ZN(n15331) );
  INV_X1 U16244 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15315) );
  NAND2_X1 U16245 ( .A1(n13005), .A2(n13004), .ZN(n13008) );
  AND2_X1 U16246 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15314) );
  NAND2_X1 U16247 ( .A1(n9835), .A2(n9834), .ZN(n13007) );
  NAND2_X1 U16248 ( .A1(n13010), .A2(n16325), .ZN(n13014) );
  NAND2_X1 U16249 ( .A1(n20280), .A2(P1_REIP_REG_31__SCAN_IN), .ZN(n15298) );
  NAND2_X1 U16250 ( .A1(n20242), .A2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n13011) );
  OAI211_X1 U16251 ( .C1(n13837), .C2(n20252), .A(n15298), .B(n13011), .ZN(
        n13012) );
  INV_X1 U16252 ( .A(n13012), .ZN(n13013) );
  OAI211_X1 U16253 ( .C1(n15303), .C2(n20088), .A(n13014), .B(n13013), .ZN(
        P1_U2968) );
  INV_X1 U16254 ( .A(n13015), .ZN(n13016) );
  XNOR2_X1 U16255 ( .A(n14820), .B(n13016), .ZN(n15126) );
  AND2_X1 U16256 ( .A1(n11641), .A2(n11979), .ZN(n13020) );
  INV_X1 U16257 ( .A(n13020), .ZN(n13017) );
  AND2_X1 U16258 ( .A1(n13017), .A2(n11643), .ZN(n13018) );
  NAND2_X1 U16259 ( .A1(n15126), .A2(n13019), .ZN(n13027) );
  INV_X1 U16260 ( .A(DATAI_14_), .ZN(n13021) );
  INV_X1 U16261 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n13486) );
  MUX2_X1 U16262 ( .A(n13021), .B(n13486), .S(n20303), .Z(n15111) );
  OAI22_X1 U16263 ( .A1(n15091), .A2(n15111), .B1(n13022), .B2(n15090), .ZN(
        n13023) );
  AOI21_X1 U16264 ( .B1(n16295), .B2(DATAI_30_), .A(n13023), .ZN(n13024) );
  INV_X1 U16265 ( .A(n13024), .ZN(n13025) );
  NOR2_X1 U16266 ( .A1(n13025), .A2(n10368), .ZN(n13026) );
  NAND2_X1 U16267 ( .A1(n13027), .A2(n13026), .ZN(P1_U2874) );
  AOI22_X1 U16268 ( .A1(n17365), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n17343), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n13028) );
  OAI21_X1 U16269 ( .B1(n12537), .B2(n17144), .A(n13028), .ZN(n13037) );
  AOI22_X1 U16270 ( .A1(n13080), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n17361), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n13035) );
  INV_X1 U16271 ( .A(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n17273) );
  OAI22_X1 U16272 ( .A1(n9919), .A2(n17273), .B1(n9827), .B2(n21152), .ZN(
        n13033) );
  AOI22_X1 U16273 ( .A1(n13120), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n13068), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n13031) );
  AOI22_X1 U16274 ( .A1(n12552), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n13064), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n13030) );
  AOI22_X1 U16275 ( .A1(n17344), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n13079), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n13029) );
  NAND3_X1 U16276 ( .A1(n13031), .A2(n13030), .A3(n13029), .ZN(n13032) );
  AOI211_X1 U16277 ( .C1(n17379), .C2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A(
        n13033), .B(n13032), .ZN(n13034) );
  OAI211_X1 U16278 ( .C1(n17384), .C2(n17401), .A(n13035), .B(n13034), .ZN(
        n13036) );
  AOI22_X1 U16279 ( .A1(n9829), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17343), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n13038) );
  OAI21_X1 U16280 ( .B1(n9919), .B2(n21277), .A(n13038), .ZN(n13048) );
  AOI22_X1 U16281 ( .A1(n17379), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n13080), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n13046) );
  AOI22_X1 U16282 ( .A1(n13089), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17361), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n13039) );
  OAI21_X1 U16283 ( .B1(n17384), .B2(n17407), .A(n13039), .ZN(n13044) );
  INV_X1 U16284 ( .A(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n13042) );
  AOI22_X1 U16285 ( .A1(n13120), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n17365), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13041) );
  AOI22_X1 U16286 ( .A1(n17245), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n13068), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n13040) );
  OAI211_X1 U16287 ( .C1(n17363), .C2(n13042), .A(n13041), .B(n13040), .ZN(
        n13043) );
  AOI211_X1 U16288 ( .C1(n13079), .C2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A(
        n13044), .B(n13043), .ZN(n13045) );
  OAI211_X1 U16289 ( .C1(n17283), .C2(n17200), .A(n13046), .B(n13045), .ZN(
        n13047) );
  OAI21_X1 U16290 ( .B1(n13050), .B2(n21140), .A(n13049), .ZN(n13055) );
  INV_X1 U16291 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17414) );
  INV_X1 U16292 ( .A(n13051), .ZN(n17309) );
  AOI22_X1 U16293 ( .A1(n17309), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17386), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n13053) );
  AOI22_X1 U16294 ( .A1(n17379), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17245), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n13052) );
  OAI211_X1 U16295 ( .C1(n17384), .C2(n17414), .A(n13053), .B(n13052), .ZN(
        n13054) );
  AOI211_X1 U16296 ( .C1(n13079), .C2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A(
        n13055), .B(n13054), .ZN(n13063) );
  AOI22_X1 U16297 ( .A1(n13120), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n13089), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n13062) );
  AOI22_X1 U16298 ( .A1(n17365), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17343), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n13057) );
  OAI21_X1 U16299 ( .B1(n17340), .B2(n13058), .A(n13057), .ZN(n13059) );
  INV_X1 U16300 ( .A(n13059), .ZN(n13060) );
  INV_X1 U16301 ( .A(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n21293) );
  AOI22_X1 U16302 ( .A1(n17365), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n17343), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n13066) );
  AOI22_X1 U16303 ( .A1(n12552), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n13064), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n13065) );
  OAI211_X1 U16304 ( .C1(n17363), .C2(n21293), .A(n13066), .B(n13065), .ZN(
        n13067) );
  INV_X1 U16305 ( .A(n13067), .ZN(n13072) );
  AOI22_X1 U16306 ( .A1(n13089), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n13068), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n13071) );
  NOR2_X1 U16307 ( .A1(n17252), .A2(n21306), .ZN(n13069) );
  NAND3_X1 U16308 ( .A1(n13072), .A2(n13071), .A3(n13070), .ZN(n13078) );
  AOI22_X1 U16309 ( .A1(n17379), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17245), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n13076) );
  AOI22_X1 U16310 ( .A1(n17309), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17386), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n13075) );
  AOI22_X1 U16311 ( .A1(n13080), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n13079), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n13074) );
  NAND2_X1 U16312 ( .A1(n17361), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n13073) );
  NAND4_X1 U16313 ( .A1(n13076), .A2(n13075), .A3(n13074), .A4(n13073), .ZN(
        n13077) );
  INV_X1 U16314 ( .A(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n21275) );
  AOI22_X1 U16315 ( .A1(n13080), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n13079), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n13081) );
  OAI21_X1 U16316 ( .B1(n17363), .B2(n21275), .A(n13081), .ZN(n13087) );
  AOI22_X1 U16317 ( .A1(n17379), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_7__1__SCAN_IN), .B2(n13082), .ZN(n13085) );
  AOI22_X1 U16318 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n13083), .B1(
        n13120), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n13084) );
  OAI211_X1 U16319 ( .C1(n21090), .C2(n17384), .A(n13085), .B(n13084), .ZN(
        n13086) );
  AOI211_X1 U16320 ( .C1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .C2(n17361), .A(
        n13087), .B(n13086), .ZN(n13096) );
  INV_X1 U16321 ( .A(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n17261) );
  AOI22_X1 U16322 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n12631), .B1(
        n13089), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n13090) );
  INV_X1 U16323 ( .A(n13090), .ZN(n13093) );
  NAND2_X1 U16324 ( .A1(n17568), .A2(n13214), .ZN(n13137) );
  NOR2_X1 U16325 ( .A1(n17564), .A2(n13137), .ZN(n13117) );
  AOI22_X1 U16326 ( .A1(n17344), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n17361), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n13106) );
  AOI22_X1 U16327 ( .A1(n13120), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n17385), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n13098) );
  AOI22_X1 U16328 ( .A1(n12552), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n9829), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n13097) );
  OAI211_X1 U16329 ( .C1(n17384), .C2(n17411), .A(n13098), .B(n13097), .ZN(
        n13104) );
  AOI22_X1 U16330 ( .A1(n17357), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17365), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n13102) );
  AOI22_X1 U16331 ( .A1(n17379), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17343), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n13101) );
  AOI22_X1 U16332 ( .A1(n17309), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17245), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n13100) );
  NAND2_X1 U16333 ( .A1(n13089), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n13099) );
  NAND4_X1 U16334 ( .A1(n13102), .A2(n13101), .A3(n13100), .A4(n13099), .ZN(
        n13103) );
  AOI211_X1 U16335 ( .C1(n13079), .C2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A(
        n13104), .B(n13103), .ZN(n13105) );
  OAI211_X1 U16336 ( .C1(n17395), .C2(n17217), .A(n13106), .B(n13105), .ZN(
        n13206) );
  NAND2_X1 U16337 ( .A1(n13117), .A2(n13206), .ZN(n13143) );
  AOI22_X1 U16338 ( .A1(n17309), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n13089), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n13116) );
  INV_X1 U16339 ( .A(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17290) );
  AOI22_X1 U16340 ( .A1(n17385), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n9829), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n13108) );
  AOI22_X1 U16341 ( .A1(n12552), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17343), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n13107) );
  OAI211_X1 U16342 ( .C1(n17384), .C2(n17290), .A(n13108), .B(n13107), .ZN(
        n13114) );
  AOI22_X1 U16343 ( .A1(n17245), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17365), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n13112) );
  AOI22_X1 U16344 ( .A1(n17379), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17386), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n13111) );
  AOI22_X1 U16345 ( .A1(n13080), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17361), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n13110) );
  NAND2_X1 U16346 ( .A1(n13079), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n13109) );
  NAND4_X1 U16347 ( .A1(n13112), .A2(n13111), .A3(n13110), .A4(n13109), .ZN(
        n13113) );
  AOI211_X1 U16348 ( .C1(n17344), .C2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A(
        n13114), .B(n13113), .ZN(n13115) );
  OAI211_X1 U16349 ( .C1(n17252), .C2(n21237), .A(n13116), .B(n13115), .ZN(
        n17553) );
  INV_X1 U16350 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n17744) );
  INV_X1 U16351 ( .A(n13206), .ZN(n17560) );
  XNOR2_X1 U16352 ( .A(n17560), .B(n13117), .ZN(n13141) );
  NAND2_X1 U16353 ( .A1(n17581), .A2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13134) );
  XNOR2_X1 U16354 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B(n13214), .ZN(
        n18037) );
  INV_X1 U16355 ( .A(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n17389) );
  AOI22_X1 U16356 ( .A1(n13080), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n17361), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n13119) );
  OAI21_X1 U16357 ( .B1(n17384), .B2(n17389), .A(n13119), .ZN(n13125) );
  AOI22_X1 U16358 ( .A1(n17357), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n13120), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n13122) );
  AOI22_X1 U16359 ( .A1(n17309), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n9829), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n13121) );
  OAI211_X1 U16360 ( .C1(n17363), .C2(n13123), .A(n13122), .B(n13121), .ZN(
        n13124) );
  AOI211_X1 U16361 ( .C1(n13079), .C2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A(
        n13125), .B(n13124), .ZN(n13133) );
  AOI22_X1 U16362 ( .A1(n17245), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n13089), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n13132) );
  INV_X1 U16363 ( .A(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n13982) );
  AOI22_X1 U16364 ( .A1(n12631), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17365), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n13126) );
  OAI21_X1 U16365 ( .B1(n9884), .B2(n13982), .A(n13126), .ZN(n13130) );
  INV_X1 U16366 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n18977) );
  NOR2_X1 U16367 ( .A1(n10364), .A2(n18977), .ZN(n18044) );
  NAND2_X1 U16368 ( .A1(n18037), .A2(n18044), .ZN(n18036) );
  NAND2_X1 U16369 ( .A1(n13134), .A2(n18036), .ZN(n18028) );
  NAND2_X1 U16370 ( .A1(n18029), .A2(n18028), .ZN(n18027) );
  NAND2_X1 U16371 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n13135), .ZN(
        n13136) );
  NAND2_X1 U16372 ( .A1(n18027), .A2(n13136), .ZN(n18017) );
  XOR2_X1 U16373 ( .A(n17564), .B(n13137), .Z(n13138) );
  INV_X1 U16374 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n18311) );
  XNOR2_X1 U16375 ( .A(n13138), .B(n18311), .ZN(n18018) );
  NAND2_X1 U16376 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n13138), .ZN(
        n13139) );
  XNOR2_X1 U16377 ( .A(n13141), .B(n13140), .ZN(n18009) );
  NOR2_X1 U16378 ( .A1(n13141), .A2(n13140), .ZN(n13142) );
  XOR2_X1 U16379 ( .A(n17557), .B(n13143), .Z(n17996) );
  XOR2_X1 U16380 ( .A(n17553), .B(n13144), .Z(n13145) );
  XOR2_X1 U16381 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B(n13145), .Z(
        n13742) );
  NAND2_X1 U16382 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n13145), .ZN(
        n13146) );
  NAND2_X1 U16383 ( .A1(n13741), .A2(n13146), .ZN(n13148) );
  AOI21_X1 U16384 ( .B1(n17551), .B2(n16638), .A(n17957), .ZN(n13149) );
  NAND2_X1 U16385 ( .A1(n13149), .A2(n13148), .ZN(n13150) );
  NAND2_X1 U16386 ( .A1(n17942), .A2(n18269), .ZN(n17933) );
  INV_X1 U16387 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n17920) );
  NOR3_X1 U16388 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n13151) );
  INV_X1 U16389 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n13152) );
  INV_X1 U16390 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18258) );
  NOR2_X1 U16391 ( .A1(n18269), .A2(n18258), .ZN(n18240) );
  NAND2_X1 U16392 ( .A1(n18240), .A2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n18250) );
  NAND2_X1 U16393 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n13230) );
  NOR2_X1 U16394 ( .A1(n18250), .A2(n13230), .ZN(n17869) );
  NAND2_X1 U16395 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n17869), .ZN(
        n18177) );
  NAND2_X1 U16396 ( .A1(n17896), .A2(n17853), .ZN(n13153) );
  INV_X1 U16397 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n18181) );
  INV_X1 U16398 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n17847) );
  INV_X1 U16399 ( .A(n13153), .ZN(n13154) );
  NOR2_X1 U16400 ( .A1(n13155), .A2(n13154), .ZN(n17852) );
  NAND2_X1 U16401 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n17836) );
  INV_X1 U16402 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n17801) );
  NOR2_X1 U16403 ( .A1(n18156), .A2(n18115), .ZN(n18132) );
  INV_X1 U16404 ( .A(n18132), .ZN(n17798) );
  NOR3_X1 U16405 ( .A1(n17801), .A2(n17828), .A3(n17798), .ZN(n13162) );
  NAND2_X1 U16406 ( .A1(n18161), .A2(n13162), .ZN(n18114) );
  INV_X1 U16407 ( .A(n18114), .ZN(n18120) );
  NAND2_X1 U16408 ( .A1(n18120), .A2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n18095) );
  NOR2_X1 U16409 ( .A1(n18094), .A2(n18095), .ZN(n17749) );
  INV_X1 U16410 ( .A(n17749), .ZN(n17755) );
  NAND2_X1 U16411 ( .A1(n17828), .A2(n13160), .ZN(n17827) );
  NOR2_X1 U16412 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17827), .ZN(
        n13156) );
  NAND2_X1 U16413 ( .A1(n13156), .A2(n18115), .ZN(n17796) );
  NOR2_X1 U16414 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17796), .ZN(
        n17778) );
  NAND3_X1 U16415 ( .A1(n17778), .A2(n18094), .A3(n18127), .ZN(n13157) );
  INV_X1 U16416 ( .A(n13158), .ZN(n13159) );
  INV_X1 U16417 ( .A(n17756), .ZN(n17743) );
  MUX2_X1 U16418 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B(n17743), .S(
        n13160), .Z(n13163) );
  OR2_X1 U16419 ( .A1(n17836), .A2(n17852), .ZN(n17795) );
  NAND2_X1 U16420 ( .A1(n13162), .A2(n17829), .ZN(n17779) );
  NOR2_X1 U16421 ( .A1(n18127), .A2(n17779), .ZN(n17760) );
  INV_X1 U16422 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n18054) );
  NAND2_X1 U16423 ( .A1(n17957), .A2(n13164), .ZN(n17742) );
  NAND2_X1 U16424 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n13258) );
  INV_X1 U16425 ( .A(n13258), .ZN(n17694) );
  NAND2_X1 U16426 ( .A1(n16164), .A2(n16610), .ZN(n16216) );
  INV_X1 U16427 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n16603) );
  AOI21_X1 U16428 ( .B1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n16216), .A(
        n13166), .ZN(n13170) );
  INV_X1 U16429 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n18975) );
  AOI22_X1 U16430 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n13160), .B1(
        n17957), .B2(n18975), .ZN(n13169) );
  OAI21_X1 U16431 ( .B1(n13166), .B2(n13160), .A(n16216), .ZN(n13167) );
  NAND2_X1 U16432 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n18975), .ZN(
        n13264) );
  NAND3_X1 U16433 ( .A1(n13167), .A2(n13264), .A3(n13169), .ZN(n13168) );
  OAI21_X1 U16434 ( .B1(n13170), .B2(n13169), .A(n13168), .ZN(n13256) );
  NAND2_X1 U16435 ( .A1(n16232), .A2(n18387), .ZN(n13179) );
  NAND2_X1 U16436 ( .A1(n19012), .A2(n18378), .ZN(n13182) );
  NAND2_X1 U16437 ( .A1(n13179), .A2(n13182), .ZN(n19029) );
  NOR2_X1 U16438 ( .A1(n13171), .A2(n18387), .ZN(n13174) );
  INV_X1 U16439 ( .A(n13173), .ZN(n13175) );
  NAND2_X1 U16440 ( .A1(n18393), .A2(n13184), .ZN(n16731) );
  NAND2_X1 U16441 ( .A1(n16732), .A2(n16146), .ZN(n13185) );
  NOR2_X1 U16442 ( .A1(n13175), .A2(n18397), .ZN(n13178) );
  NOR2_X1 U16443 ( .A1(n13176), .A2(n18409), .ZN(n16234) );
  INV_X1 U16444 ( .A(n16234), .ZN(n18820) );
  NOR2_X1 U16445 ( .A1(n18820), .A2(n18401), .ZN(n13177) );
  INV_X1 U16446 ( .A(n13179), .ZN(n13196) );
  OAI21_X1 U16447 ( .B1(n13196), .B2(n18393), .A(n13246), .ZN(n13180) );
  NOR2_X1 U16448 ( .A1(n17547), .A2(n16234), .ZN(n16233) );
  NOR2_X1 U16449 ( .A1(n16233), .A2(n13182), .ZN(n13243) );
  NOR2_X2 U16450 ( .A1(n18831), .A2(n18824), .ZN(n18222) );
  INV_X1 U16451 ( .A(n13185), .ZN(n13292) );
  NAND3_X1 U16452 ( .A1(n18387), .A2(n13292), .A3(n13195), .ZN(n13187) );
  NAND2_X1 U16453 ( .A1(n13187), .A2(n13186), .ZN(n18814) );
  AOI21_X4 U16454 ( .B1(n18815), .B2(n13290), .A(n18814), .ZN(n18821) );
  NOR2_X1 U16455 ( .A1(n13193), .A2(n13189), .ZN(n13252) );
  XNOR2_X1 U16456 ( .A(n13191), .B(n13190), .ZN(n13194) );
  NOR2_X1 U16457 ( .A1(n13252), .A2(n18802), .ZN(n18800) );
  NOR2_X1 U16458 ( .A1(n19012), .A2(n18393), .ZN(n13249) );
  NAND2_X1 U16459 ( .A1(n13249), .A2(n18409), .ZN(n13251) );
  AOI211_X1 U16460 ( .C1(n18401), .C2(n18820), .A(n13196), .B(n13195), .ZN(
        n13197) );
  NAND2_X1 U16461 ( .A1(n13198), .A2(n13197), .ZN(n13245) );
  NAND2_X2 U16462 ( .A1(n13232), .A2(n18387), .ZN(n18049) );
  NOR2_X2 U16463 ( .A1(n17551), .A2(n18049), .ZN(n17963) );
  NAND2_X1 U16464 ( .A1(n13256), .A2(n17963), .ZN(n13242) );
  NOR3_X1 U16465 ( .A1(n13258), .A2(n17693), .A3(n10180), .ZN(n13263) );
  NAND2_X1 U16466 ( .A1(n17749), .A2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n17729) );
  INV_X1 U16467 ( .A(n13199), .ZN(n13200) );
  NOR2_X1 U16468 ( .A1(n17896), .A2(n13200), .ZN(n18289) );
  INV_X1 U16469 ( .A(n18289), .ZN(n17960) );
  NOR2_X2 U16470 ( .A1(n17956), .A2(n18283), .ZN(n18214) );
  NAND2_X1 U16471 ( .A1(n18228), .A2(n18214), .ZN(n18217) );
  NOR2_X2 U16472 ( .A1(n13230), .A2(n18217), .ZN(n18189) );
  NAND2_X1 U16473 ( .A1(n13263), .A2(n17741), .ZN(n16625) );
  NOR2_X1 U16474 ( .A1(n16610), .A2(n16625), .ZN(n16608) );
  NAND2_X1 U16475 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16608), .ZN(
        n13201) );
  XNOR2_X1 U16476 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n13201), .ZN(
        n13271) );
  NOR2_X2 U16477 ( .A1(n16624), .A2(n18049), .ZN(n17926) );
  NOR2_X1 U16478 ( .A1(n13210), .A2(n17568), .ZN(n13208) );
  NOR2_X1 U16479 ( .A1(n13208), .A2(n17564), .ZN(n13207) );
  NAND2_X1 U16480 ( .A1(n13207), .A2(n13206), .ZN(n13204) );
  NOR2_X1 U16481 ( .A1(n17557), .A2(n13204), .ZN(n13203) );
  NAND2_X1 U16482 ( .A1(n13203), .A2(n17553), .ZN(n13202) );
  NOR2_X1 U16483 ( .A1(n17551), .A2(n13202), .ZN(n13228) );
  XNOR2_X1 U16484 ( .A(n13202), .B(n16624), .ZN(n17977) );
  XOR2_X1 U16485 ( .A(n13203), .B(n17553), .Z(n13221) );
  XOR2_X1 U16486 ( .A(n13204), .B(n17557), .Z(n13205) );
  NAND2_X1 U16487 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n13205), .ZN(
        n13220) );
  XNOR2_X1 U16488 ( .A(n18308), .B(n13205), .ZN(n17992) );
  XOR2_X1 U16489 ( .A(n13207), .B(n13206), .Z(n13218) );
  XOR2_X1 U16490 ( .A(n13208), .B(n17564), .Z(n13209) );
  NAND2_X1 U16491 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n13209), .ZN(
        n13216) );
  XNOR2_X1 U16492 ( .A(n18311), .B(n13209), .ZN(n18016) );
  NAND2_X1 U16493 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n13211), .ZN(
        n13215) );
  XOR2_X1 U16494 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n13211), .Z(
        n18026) );
  INV_X1 U16495 ( .A(n10364), .ZN(n16235) );
  AOI21_X1 U16496 ( .B1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n13214), .A(
        n16235), .ZN(n13213) );
  NOR2_X1 U16497 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n13214), .ZN(
        n13212) );
  AOI221_X1 U16498 ( .B1(n16235), .B2(n13214), .C1(n13213), .C2(n18977), .A(
        n13212), .ZN(n18025) );
  NAND2_X1 U16499 ( .A1(n18026), .A2(n18025), .ZN(n18024) );
  NAND2_X1 U16500 ( .A1(n13215), .A2(n18024), .ZN(n18015) );
  NAND2_X1 U16501 ( .A1(n18016), .A2(n18015), .ZN(n18014) );
  NAND2_X1 U16502 ( .A1(n13216), .A2(n18014), .ZN(n13217) );
  NAND2_X1 U16503 ( .A1(n13218), .A2(n13217), .ZN(n13219) );
  NAND2_X1 U16504 ( .A1(n13220), .A2(n17990), .ZN(n13222) );
  NAND2_X1 U16505 ( .A1(n13221), .A2(n13222), .ZN(n13223) );
  XOR2_X1 U16506 ( .A(n13222), .B(n13221), .Z(n13745) );
  NAND2_X1 U16507 ( .A1(n13228), .A2(n13224), .ZN(n13229) );
  INV_X1 U16508 ( .A(n13224), .ZN(n13227) );
  NAND2_X1 U16509 ( .A1(n17977), .A2(n17976), .ZN(n13226) );
  NAND2_X1 U16510 ( .A1(n13228), .A2(n13227), .ZN(n13225) );
  OAI211_X1 U16511 ( .C1(n13228), .C2(n13227), .A(n13226), .B(n13225), .ZN(
        n17959) );
  NAND2_X1 U16512 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n17959), .ZN(
        n17958) );
  NAND2_X1 U16513 ( .A1(n17734), .A2(n13263), .ZN(n16631) );
  NAND2_X1 U16514 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16609), .ZN(
        n13231) );
  XOR2_X1 U16515 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n13231), .Z(
        n13269) );
  INV_X1 U16516 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n18994) );
  NAND2_X1 U16517 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_2__SCAN_IN), .ZN(n18367) );
  NAND2_X1 U16518 ( .A1(n18967), .A2(n18367), .ZN(n19019) );
  NAND2_X1 U16519 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n18006) );
  NAND2_X1 U16520 ( .A1(n17993), .A2(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n17971) );
  NAND2_X1 U16521 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n17902) );
  NAND2_X1 U16522 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n17857) );
  NAND3_X1 U16523 ( .A1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n17805) );
  NOR2_X1 U16524 ( .A1(n17805), .A2(n17804), .ZN(n13296) );
  NAND2_X1 U16525 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n17786) );
  NAND2_X1 U16526 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n17766), .ZN(
        n17736) );
  NAND2_X1 U16527 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n17737) );
  NAND2_X1 U16528 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n17703) );
  NAND2_X1 U16529 ( .A1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n16614), .ZN(
        n13233) );
  INV_X1 U16530 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n18951) );
  NOR2_X1 U16531 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n19028) );
  NAND3_X2 U16532 ( .A1(n19028), .A2(n19017), .A3(n19027), .ZN(n18316) );
  NOR2_X1 U16533 ( .A1(n18951), .A2(n18316), .ZN(n13265) );
  NAND2_X1 U16534 ( .A1(n18994), .A2(n19027), .ZN(n19016) );
  INV_X1 U16535 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n19013) );
  OR2_X1 U16536 ( .A1(n13235), .A2(n17901), .ZN(n16599) );
  INV_X1 U16537 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n16754) );
  XOR2_X1 U16538 ( .A(n16754), .B(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .Z(
        n13237) );
  NOR2_X1 U16539 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n17776), .ZN(
        n16616) );
  NOR2_X1 U16540 ( .A1(n18040), .A2(n17702), .ZN(n16749) );
  INV_X1 U16541 ( .A(n16749), .ZN(n13234) );
  NOR2_X1 U16542 ( .A1(n13234), .A2(n17703), .ZN(n16747) );
  NAND2_X1 U16543 ( .A1(n18748), .A2(n13235), .ZN(n13236) );
  OAI211_X1 U16544 ( .C1(n16747), .C2(n18046), .A(n18045), .B(n13236), .ZN(
        n16617) );
  NOR2_X1 U16545 ( .A1(n16616), .A2(n16617), .ZN(n16598) );
  OAI22_X1 U16546 ( .A1(n16599), .A2(n13237), .B1(n16598), .B2(n16754), .ZN(
        n13238) );
  AOI211_X1 U16547 ( .C1(n17895), .C2(n17101), .A(n13265), .B(n13238), .ZN(
        n13239) );
  NAND2_X1 U16548 ( .A1(n13242), .A2(n13241), .ZN(P3_U2799) );
  AOI211_X1 U16549 ( .C1(n16731), .C2(n13245), .A(n13244), .B(n13243), .ZN(
        n16148) );
  OAI21_X1 U16550 ( .B1(n18393), .B2(n13246), .A(n10005), .ZN(n13254) );
  INV_X1 U16551 ( .A(n18802), .ZN(n16230) );
  INV_X1 U16552 ( .A(n18393), .ZN(n13247) );
  NAND2_X2 U16553 ( .A1(n18960), .A2(P3_STATE_REG_2__SCAN_IN), .ZN(n18954) );
  OAI21_X1 U16554 ( .B1(n13247), .B2(n18387), .A(n19011), .ZN(n13248) );
  OAI21_X1 U16555 ( .B1(n13249), .B2(n13248), .A(n18858), .ZN(n16729) );
  OAI22_X1 U16556 ( .A1(n13252), .A2(n13251), .B1(n13250), .B2(n16729), .ZN(
        n13253) );
  AOI22_X1 U16557 ( .A1(n18808), .A2(n13254), .B1(n16230), .B2(n13253), .ZN(
        n13255) );
  NAND2_X1 U16558 ( .A1(n13256), .A2(n18287), .ZN(n13273) );
  NAND2_X1 U16559 ( .A1(n18804), .A2(n18359), .ZN(n18358) );
  NOR2_X1 U16560 ( .A1(n16624), .A2(n18358), .ZN(n18288) );
  NAND2_X1 U16561 ( .A1(n18244), .A2(n18359), .ZN(n18326) );
  INV_X1 U16562 ( .A(n18276), .ZN(n18280) );
  NOR3_X1 U16563 ( .A1(n17693), .A2(n10180), .A3(n16610), .ZN(n16604) );
  NAND2_X1 U16564 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18315) );
  NAND3_X1 U16565 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n13748) );
  NOR2_X1 U16566 ( .A1(n18315), .A2(n13748), .ZN(n13739) );
  NAND3_X1 U16567 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A3(n13739), .ZN(n18268) );
  NOR2_X1 U16568 ( .A1(n18283), .A2(n18268), .ZN(n18239) );
  NAND2_X1 U16569 ( .A1(n17853), .A2(n18239), .ZN(n18111) );
  NOR2_X1 U16570 ( .A1(n18095), .A2(n18111), .ZN(n18056) );
  NOR3_X1 U16571 ( .A1(n18094), .A2(n18098), .A3(n13258), .ZN(n17716) );
  NAND2_X1 U16572 ( .A1(n18056), .A2(n17716), .ZN(n13260) );
  NAND2_X1 U16573 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n18239), .ZN(
        n18199) );
  NOR2_X1 U16574 ( .A1(n16637), .A2(n18199), .ZN(n18179) );
  AOI21_X1 U16575 ( .B1(n18120), .B2(n18179), .A(n18821), .ZN(n18118) );
  NAND2_X1 U16576 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n17716), .ZN(
        n17698) );
  NOR2_X1 U16577 ( .A1(n18127), .A2(n17698), .ZN(n16634) );
  AOI21_X1 U16578 ( .B1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18312) );
  NOR2_X1 U16579 ( .A1(n18312), .A2(n13748), .ZN(n13738) );
  NAND4_X1 U16580 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A4(n13738), .ZN(n18176) );
  OR2_X1 U16581 ( .A1(n16637), .A2(n18176), .ZN(n18158) );
  OAI21_X1 U16582 ( .B1(n17729), .B2(n18158), .A(n18831), .ZN(n13257) );
  INV_X1 U16583 ( .A(n13257), .ZN(n18077) );
  NOR2_X1 U16584 ( .A1(n13258), .A2(n18077), .ZN(n18055) );
  OAI22_X1 U16585 ( .A1(n18821), .A2(n16634), .B1(n18055), .B2(n18807), .ZN(
        n13259) );
  AOI211_X1 U16586 ( .C1(n18824), .C2(n13260), .A(n18118), .B(n13259), .ZN(
        n16161) );
  OAI21_X1 U16587 ( .B1(n18280), .B2(n16604), .A(n16161), .ZN(n13261) );
  AOI21_X1 U16588 ( .B1(n18359), .B2(n13261), .A(n16603), .ZN(n16221) );
  NAND2_X1 U16589 ( .A1(n18359), .A2(n18276), .ZN(n18351) );
  OAI21_X1 U16590 ( .B1(n16221), .B2(n18351), .A(n18350), .ZN(n13267) );
  INV_X1 U16591 ( .A(n18821), .ZN(n18813) );
  AOI21_X1 U16592 ( .B1(n18813), .B2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n18824), .ZN(n18337) );
  OAI22_X1 U16593 ( .A1(n18807), .A2(n18158), .B1(n18337), .B2(n18111), .ZN(
        n13262) );
  INV_X1 U16594 ( .A(n13262), .ZN(n18052) );
  NOR2_X1 U16595 ( .A1(n18052), .A2(n17729), .ZN(n18075) );
  NAND3_X1 U16596 ( .A1(n13263), .A2(n18359), .A3(n18075), .ZN(n16168) );
  NOR3_X1 U16597 ( .A1(n16610), .A2(n13264), .A3(n16168), .ZN(n13266) );
  AOI211_X1 U16598 ( .C1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .C2(n13267), .A(
        n13266), .B(n13265), .ZN(n13268) );
  NAND2_X1 U16599 ( .A1(n13273), .A2(n13272), .ZN(P3_U2831) );
  INV_X1 U16600 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n20998) );
  NOR3_X1 U16601 ( .A1(P1_BE_N_REG_2__SCAN_IN), .A2(P1_BE_N_REG_0__SCAN_IN), 
        .A3(n20998), .ZN(n13275) );
  NOR4_X1 U16602 ( .A1(P1_BE_N_REG_1__SCAN_IN), .A2(P1_BE_N_REG_3__SCAN_IN), 
        .A3(P1_D_C_N_REG_SCAN_IN), .A4(P1_ADS_N_REG_SCAN_IN), .ZN(n13274) );
  NOR4_X1 U16603 ( .A1(P2_ADDRESS_REG_15__SCAN_IN), .A2(
        P2_ADDRESS_REG_14__SCAN_IN), .A3(P2_ADDRESS_REG_13__SCAN_IN), .A4(
        P2_ADDRESS_REG_12__SCAN_IN), .ZN(n13279) );
  NOR4_X1 U16604 ( .A1(P2_ADDRESS_REG_19__SCAN_IN), .A2(
        P2_ADDRESS_REG_18__SCAN_IN), .A3(P2_ADDRESS_REG_17__SCAN_IN), .A4(
        P2_ADDRESS_REG_16__SCAN_IN), .ZN(n13278) );
  NOR4_X1 U16605 ( .A1(P2_ADDRESS_REG_6__SCAN_IN), .A2(
        P2_ADDRESS_REG_5__SCAN_IN), .A3(P2_ADDRESS_REG_4__SCAN_IN), .A4(
        P2_ADDRESS_REG_3__SCAN_IN), .ZN(n13277) );
  NOR4_X1 U16606 ( .A1(P2_ADDRESS_REG_11__SCAN_IN), .A2(
        P2_ADDRESS_REG_9__SCAN_IN), .A3(P2_ADDRESS_REG_8__SCAN_IN), .A4(
        P2_ADDRESS_REG_7__SCAN_IN), .ZN(n13276) );
  NAND4_X1 U16607 ( .A1(n13279), .A2(n13278), .A3(n13277), .A4(n13276), .ZN(
        n13284) );
  NOR4_X1 U16608 ( .A1(P2_ADDRESS_REG_1__SCAN_IN), .A2(
        P2_ADDRESS_REG_0__SCAN_IN), .A3(P2_ADDRESS_REG_10__SCAN_IN), .A4(
        P2_ADDRESS_REG_23__SCAN_IN), .ZN(n13282) );
  NOR4_X1 U16609 ( .A1(P2_ADDRESS_REG_24__SCAN_IN), .A2(
        P2_ADDRESS_REG_22__SCAN_IN), .A3(P2_ADDRESS_REG_21__SCAN_IN), .A4(
        P2_ADDRESS_REG_20__SCAN_IN), .ZN(n13281) );
  NOR4_X1 U16610 ( .A1(P2_ADDRESS_REG_28__SCAN_IN), .A2(
        P2_ADDRESS_REG_27__SCAN_IN), .A3(P2_ADDRESS_REG_26__SCAN_IN), .A4(
        P2_ADDRESS_REG_25__SCAN_IN), .ZN(n13280) );
  NAND4_X1 U16611 ( .A1(n13282), .A2(n13281), .A3(n13280), .A4(n19939), .ZN(
        n13283) );
  NOR2_X1 U16612 ( .A1(P2_BE_N_REG_0__SCAN_IN), .A2(P2_BE_N_REG_1__SCAN_IN), 
        .ZN(n13287) );
  NOR4_X1 U16613 ( .A1(P2_BE_N_REG_2__SCAN_IN), .A2(P2_BE_N_REG_3__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n13286) );
  NAND4_X1 U16614 ( .A1(P2_M_IO_N_REG_SCAN_IN), .A2(P2_W_R_N_REG_SCAN_IN), 
        .A3(n13287), .A4(n13286), .ZN(n13288) );
  NOR2_X4 U16615 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n13288), .ZN(n16717)
         );
  INV_X2 U16616 ( .A(n16717), .ZN(U215) );
  NOR3_X1 U16617 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .ZN(n17084) );
  NAND2_X1 U16618 ( .A1(n17084), .A2(n17079), .ZN(n17076) );
  NOR2_X1 U16619 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n17076), .ZN(n17053) );
  INV_X1 U16620 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n17046) );
  NAND2_X1 U16621 ( .A1(n17053), .A2(n17046), .ZN(n17045) );
  NOR2_X1 U16622 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n17045), .ZN(n17029) );
  NAND2_X1 U16623 ( .A1(n17029), .A2(n17022), .ZN(n17020) );
  NOR2_X1 U16624 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n17020), .ZN(n17005) );
  NAND2_X1 U16625 ( .A1(n17005), .A2(n16996), .ZN(n16977) );
  NOR2_X1 U16626 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n16977), .ZN(n16976) );
  NAND2_X1 U16627 ( .A1(n16976), .A2(n17322), .ZN(n16969) );
  NOR2_X1 U16628 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n16969), .ZN(n16956) );
  INV_X1 U16629 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n16950) );
  NAND2_X1 U16630 ( .A1(n16956), .A2(n16950), .ZN(n16947) );
  NOR2_X1 U16631 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n16947), .ZN(n16932) );
  NAND2_X1 U16632 ( .A1(n16932), .A2(n16923), .ZN(n16922) );
  NAND2_X1 U16633 ( .A1(n16912), .A2(n16904), .ZN(n16903) );
  NAND2_X1 U16634 ( .A1(n16887), .A2(n21148), .ZN(n16874) );
  INV_X1 U16635 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n17214) );
  NAND2_X1 U16636 ( .A1(n16862), .A2(n17214), .ZN(n16854) );
  NOR2_X1 U16637 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n16854), .ZN(n16840) );
  INV_X1 U16638 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n17119) );
  NAND2_X1 U16639 ( .A1(n16840), .A2(n17119), .ZN(n16832) );
  NOR2_X1 U16640 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n16832), .ZN(n16817) );
  INV_X1 U16641 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n16807) );
  NAND2_X1 U16642 ( .A1(n16817), .A2(n16807), .ZN(n16806) );
  NOR2_X1 U16643 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n16806), .ZN(n16800) );
  INV_X1 U16644 ( .A(n13289), .ZN(n13291) );
  NAND2_X1 U16645 ( .A1(n13291), .A2(n13290), .ZN(n16152) );
  NAND2_X1 U16646 ( .A1(n13292), .A2(n16152), .ZN(n18801) );
  INV_X1 U16647 ( .A(n13305), .ZN(n13294) );
  NAND2_X1 U16648 ( .A1(n19013), .A2(n18858), .ZN(n13293) );
  NAND4_X1 U16649 ( .A1(n13294), .A2(P3_EBX_REG_31__SCAN_IN), .A3(n18387), 
        .A4(n13293), .ZN(n17110) );
  AOI211_X1 U16650 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n16806), .A(n16800), .B(
        n17110), .ZN(n13311) );
  INV_X1 U16651 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n18941) );
  INV_X1 U16652 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n18943) );
  AOI211_X1 U16653 ( .C1(n19012), .C2(n19011), .A(n9998), .B(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n13306) );
  INV_X1 U16654 ( .A(n13306), .ZN(n18856) );
  INV_X1 U16655 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n18939) );
  INV_X1 U16656 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n18916) );
  NAND3_X1 U16657 ( .A1(P3_REIP_REG_3__SCAN_IN), .A2(P3_REIP_REG_1__SCAN_IN), 
        .A3(P3_REIP_REG_2__SCAN_IN), .ZN(n17057) );
  NOR2_X1 U16658 ( .A1(n18903), .A2(n17057), .ZN(n17039) );
  NAND2_X1 U16659 ( .A1(P3_REIP_REG_5__SCAN_IN), .A2(n17039), .ZN(n16979) );
  NAND3_X1 U16660 ( .A1(P3_REIP_REG_8__SCAN_IN), .A2(P3_REIP_REG_7__SCAN_IN), 
        .A3(P3_REIP_REG_6__SCAN_IN), .ZN(n16980) );
  NAND2_X1 U16661 ( .A1(P3_REIP_REG_10__SCAN_IN), .A2(P3_REIP_REG_9__SCAN_IN), 
        .ZN(n16967) );
  NOR4_X1 U16662 ( .A1(n18916), .A2(n16979), .A3(n16980), .A4(n16967), .ZN(
        n16959) );
  NAND2_X1 U16663 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n16959), .ZN(n16942) );
  NAND2_X1 U16664 ( .A1(P3_REIP_REG_14__SCAN_IN), .A2(P3_REIP_REG_13__SCAN_IN), 
        .ZN(n16827) );
  NOR2_X1 U16665 ( .A1(n16942), .A2(n16827), .ZN(n16808) );
  INV_X1 U16666 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n18938) );
  INV_X1 U16667 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n18931) );
  NAND3_X1 U16668 ( .A1(P3_REIP_REG_17__SCAN_IN), .A2(P3_REIP_REG_16__SCAN_IN), 
        .A3(P3_REIP_REG_15__SCAN_IN), .ZN(n16877) );
  NAND2_X1 U16669 ( .A1(P3_REIP_REG_19__SCAN_IN), .A2(P3_REIP_REG_18__SCAN_IN), 
        .ZN(n16861) );
  NOR3_X1 U16670 ( .A1(n18931), .A2(n16877), .A3(n16861), .ZN(n16839) );
  NAND3_X1 U16671 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(P3_REIP_REG_21__SCAN_IN), 
        .A3(n16839), .ZN(n16828) );
  NOR2_X1 U16672 ( .A1(n18938), .A2(n16828), .ZN(n16809) );
  NAND2_X1 U16673 ( .A1(n16808), .A2(n16809), .ZN(n16820) );
  NOR2_X1 U16674 ( .A1(n18939), .A2(n16820), .ZN(n13295) );
  NAND2_X1 U16675 ( .A1(n17083), .A2(n13295), .ZN(n16804) );
  NOR3_X1 U16676 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(P3_STATE2_REG_2__SCAN_IN), .A3(P3_STATEBS16_REG_SCAN_IN), .ZN(n18877) );
  NOR2_X1 U16677 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n18967), .ZN(n18715) );
  NAND2_X1 U16678 ( .A1(n18870), .A2(n18715), .ZN(n18862) );
  NAND3_X1 U16679 ( .A1(P3_REIP_REG_26__SCAN_IN), .A2(P3_REIP_REG_25__SCAN_IN), 
        .A3(n13295), .ZN(n16752) );
  NOR2_X1 U16680 ( .A1(n17100), .A2(n16752), .ZN(n16758) );
  NOR2_X1 U16681 ( .A1(n16909), .A2(n16758), .ZN(n16789) );
  INV_X1 U16682 ( .A(n16789), .ZN(n16803) );
  AOI221_X1 U16683 ( .B1(n18941), .B2(n18943), .C1(n16804), .C2(n18943), .A(
        n16803), .ZN(n13310) );
  NAND2_X1 U16684 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17722), .ZN(
        n17691) );
  AOI21_X1 U16685 ( .B1(n10098), .B2(n17691), .A(n16749), .ZN(n17726) );
  INV_X1 U16686 ( .A(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n17768) );
  NAND2_X1 U16687 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n9922), .ZN(
        n16908) );
  NAND2_X1 U16688 ( .A1(n13296), .A2(n16896), .ZN(n13298) );
  NOR2_X1 U16689 ( .A1(n17786), .A2(n13298), .ZN(n13297) );
  INV_X1 U16690 ( .A(n13297), .ZN(n17735) );
  NAND2_X1 U16691 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n13297), .ZN(
        n13302) );
  INV_X1 U16692 ( .A(n13302), .ZN(n13301) );
  AOI21_X1 U16693 ( .B1(n17768), .B2(n17735), .A(n13301), .ZN(n17764) );
  INV_X1 U16694 ( .A(n17764), .ZN(n16835) );
  INV_X1 U16695 ( .A(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n16841) );
  INV_X1 U16696 ( .A(n13298), .ZN(n13300) );
  NAND2_X1 U16697 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n13300), .ZN(
        n13299) );
  AOI21_X1 U16698 ( .B1(n16841), .B2(n13299), .A(n13297), .ZN(n17777) );
  INV_X1 U16699 ( .A(n17777), .ZN(n16846) );
  NOR2_X1 U16700 ( .A1(n17805), .A2(n16908), .ZN(n17774) );
  OAI21_X1 U16701 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n17774), .A(
        n13298), .ZN(n17807) );
  NAND2_X1 U16702 ( .A1(n16896), .A2(n17069), .ZN(n16897) );
  NAND2_X1 U16703 ( .A1(n17101), .A2(n16867), .ZN(n16853) );
  OAI21_X1 U16704 ( .B1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n13300), .A(
        n13299), .ZN(n17790) );
  NAND2_X1 U16705 ( .A1(n16853), .A2(n17790), .ZN(n16852) );
  NAND2_X1 U16706 ( .A1(n17101), .A2(n16852), .ZN(n16845) );
  NAND2_X1 U16707 ( .A1(n16846), .A2(n16845), .ZN(n16844) );
  NAND2_X1 U16708 ( .A1(n17101), .A2(n16844), .ZN(n16834) );
  NAND2_X1 U16709 ( .A1(n16835), .A2(n16834), .ZN(n16833) );
  NAND2_X1 U16710 ( .A1(n17101), .A2(n16833), .ZN(n16824) );
  INV_X1 U16711 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n17753) );
  AOI22_X1 U16712 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n13302), .B1(
        n13301), .B2(n17753), .ZN(n17750) );
  NAND2_X1 U16713 ( .A1(n16824), .A2(n17750), .ZN(n16823) );
  NAND2_X1 U16714 ( .A1(n17101), .A2(n16823), .ZN(n16811) );
  NOR2_X1 U16715 ( .A1(n17753), .A2(n13302), .ZN(n13303) );
  OAI21_X1 U16716 ( .B1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n13303), .A(
        n17691), .ZN(n17739) );
  NAND2_X1 U16717 ( .A1(n16811), .A2(n17739), .ZN(n16810) );
  NAND2_X1 U16718 ( .A1(n17101), .A2(n16810), .ZN(n16750) );
  INV_X1 U16719 ( .A(n16750), .ZN(n13304) );
  INV_X1 U16720 ( .A(n17726), .ZN(n16751) );
  AOI221_X1 U16721 ( .B1(n17726), .B2(n13304), .C1(n16751), .C2(n16750), .A(
        n18873), .ZN(n13309) );
  AOI211_X4 U16722 ( .C1(P3_EBX_REG_31__SCAN_IN), .C2(n18387), .A(n13306), .B(
        n13305), .ZN(n17059) );
  AOI22_X1 U16723 ( .A1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n17070), .B1(
        n17059), .B2(P3_EBX_REG_26__SCAN_IN), .ZN(n13307) );
  INV_X1 U16724 ( .A(n13307), .ZN(n13308) );
  AOI211_X1 U16725 ( .C1(n15767), .C2(n13313), .A(n13312), .B(n19214), .ZN(
        n13325) );
  INV_X1 U16726 ( .A(n19205), .ZN(n19155) );
  INV_X1 U16727 ( .A(P2_EBX_REG_27__SCAN_IN), .ZN(n13314) );
  INV_X1 U16728 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n19978) );
  OAI22_X1 U16729 ( .A1(n19155), .A2(n13314), .B1(n19978), .B2(n19181), .ZN(
        n13324) );
  OAI22_X1 U16730 ( .A1(n13315), .A2(n19202), .B1(n15765), .B2(n19180), .ZN(
        n13323) );
  NOR2_X1 U16731 ( .A1(n13317), .A2(n13318), .ZN(n13319) );
  NAND2_X1 U16732 ( .A1(n15717), .A2(n13320), .ZN(n13321) );
  NAND2_X1 U16733 ( .A1(n9886), .A2(n13321), .ZN(n15884) );
  OAI22_X1 U16734 ( .A1(n15889), .A2(n19197), .B1(n15884), .B2(n19200), .ZN(
        n13322) );
  OR4_X1 U16735 ( .A1(n13325), .A2(n13324), .A3(n13323), .A4(n13322), .ZN(
        P2_U2828) );
  INV_X1 U16736 ( .A(n19208), .ZN(n19193) );
  INV_X1 U16737 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .ZN(n13327) );
  OAI211_X1 U16738 ( .C1(n19193), .C2(n13327), .A(n13326), .B(n13421), .ZN(
        P2_U2814) );
  INV_X1 U16739 ( .A(n20056), .ZN(n13330) );
  OAI21_X1 U16740 ( .B1(n13328), .B2(P2_READREQUEST_REG_SCAN_IN), .A(n13330), 
        .ZN(n13329) );
  OAI21_X1 U16741 ( .B1(n13331), .B2(n13330), .A(n13329), .ZN(P2_U3612) );
  OAI21_X1 U16742 ( .B1(n13333), .B2(n19184), .A(n13332), .ZN(n13334) );
  XNOR2_X1 U16743 ( .A(n13334), .B(n19348), .ZN(n19362) );
  NOR2_X1 U16744 ( .A1(n16559), .A2(n19191), .ZN(n13338) );
  OAI21_X1 U16745 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n13336), .A(
        n13335), .ZN(n19357) );
  NAND2_X1 U16746 ( .A1(n19170), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n19360) );
  OAI21_X1 U16747 ( .B1(n19319), .B2(n19357), .A(n19360), .ZN(n13337) );
  AOI211_X1 U16748 ( .C1(n19191), .C2(n16550), .A(n13338), .B(n13337), .ZN(
        n13340) );
  NAND2_X1 U16749 ( .A1(n19315), .A2(n9860), .ZN(n13339) );
  OAI211_X1 U16750 ( .C1(n19362), .C2(n16553), .A(n13340), .B(n13339), .ZN(
        P2_U3013) );
  AOI21_X1 U16751 ( .B1(n19201), .B2(n16105), .A(n13341), .ZN(n13376) );
  INV_X1 U16752 ( .A(n13342), .ZN(n13343) );
  OAI21_X1 U16753 ( .B1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n13344), .A(
        n13343), .ZN(n13373) );
  NAND2_X1 U16754 ( .A1(n19170), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n13365) );
  OAI21_X1 U16755 ( .B1(n19319), .B2(n13373), .A(n13365), .ZN(n13345) );
  AOI21_X1 U16756 ( .B1(n12840), .B2(n13376), .A(n13345), .ZN(n13348) );
  OAI21_X1 U16757 ( .B1(n19313), .B2(n13346), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13347) );
  OAI211_X1 U16758 ( .C1(n16545), .C2(n19198), .A(n13348), .B(n13347), .ZN(
        P2_U3014) );
  NAND2_X1 U16759 ( .A1(n13351), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n13590) );
  NOR2_X1 U16760 ( .A1(n20002), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n13352) );
  NAND2_X1 U16761 ( .A1(n20062), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n13355) );
  AND4_X1 U16762 ( .A1(n10679), .A2(n13355), .A3(P2_STATE2_REG_0__SCAN_IN), 
        .A4(n20036), .ZN(n13356) );
  NOR2_X1 U16763 ( .A1(n15661), .A2(n19198), .ZN(n13357) );
  AOI21_X1 U16764 ( .B1(P2_EBX_REG_0__SCAN_IN), .B2(n15661), .A(n13357), .ZN(
        n13358) );
  OAI21_X1 U16765 ( .B1(n15694), .B2(n19207), .A(n13358), .ZN(P2_U2887) );
  OAI21_X1 U16766 ( .B1(n13692), .B2(n13359), .A(n13657), .ZN(n13361) );
  INV_X1 U16767 ( .A(n20063), .ZN(n13360) );
  INV_X1 U16768 ( .A(n13694), .ZN(n14296) );
  OR2_X1 U16769 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n14296), .ZN(n19309) );
  INV_X2 U16770 ( .A(n19309), .ZN(n20057) );
  INV_X1 U16771 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n21162) );
  INV_X1 U16772 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n13618) );
  INV_X1 U16773 ( .A(P2_UWORD_REG_0__SCAN_IN), .ZN(n13364) );
  OAI222_X1 U16774 ( .A1(n19312), .A2(n21162), .B1(n19276), .B2(n13618), .C1(
        n13364), .C2(n19309), .ZN(P2_U2935) );
  INV_X1 U16775 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n13616) );
  INV_X1 U16776 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n16711) );
  INV_X1 U16777 ( .A(P2_UWORD_REG_5__SCAN_IN), .ZN(n21305) );
  OAI222_X1 U16778 ( .A1(n19276), .A2(n13616), .B1(n19312), .B2(n16711), .C1(
        n21305), .C2(n19309), .ZN(P2_U2930) );
  OAI21_X1 U16779 ( .B1(n19355), .B2(n19198), .A(n13365), .ZN(n13375) );
  INV_X1 U16780 ( .A(n13366), .ZN(n13372) );
  INV_X1 U16781 ( .A(n13367), .ZN(n13370) );
  INV_X1 U16782 ( .A(n13368), .ZN(n13369) );
  NAND2_X1 U16783 ( .A1(n13370), .A2(n13369), .ZN(n13371) );
  NAND2_X1 U16784 ( .A1(n13372), .A2(n13371), .ZN(n19199) );
  OAI22_X1 U16785 ( .A1(n19356), .A2(n13373), .B1(n19327), .B2(n19199), .ZN(
        n13374) );
  AOI211_X1 U16786 ( .C1(n19331), .C2(n13376), .A(n13375), .B(n13374), .ZN(
        n13378) );
  MUX2_X1 U16787 ( .A(n19353), .B(n19349), .S(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .Z(n13377) );
  NAND2_X1 U16788 ( .A1(n13378), .A2(n13377), .ZN(P2_U3046) );
  OAI22_X1 U16789 ( .A1(n14303), .A2(BUF1_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n14302), .ZN(n13653) );
  INV_X1 U16790 ( .A(n13653), .ZN(n19220) );
  NAND2_X1 U16791 ( .A1(n14108), .A2(n13379), .ZN(n13383) );
  AND2_X1 U16792 ( .A1(n13380), .A2(n20069), .ZN(n14114) );
  NAND2_X1 U16793 ( .A1(n14104), .A2(n14114), .ZN(n13381) );
  OR2_X1 U16794 ( .A1(n14115), .A2(n13381), .ZN(n13382) );
  NAND2_X1 U16795 ( .A1(n13383), .A2(n13382), .ZN(n13687) );
  INV_X1 U16796 ( .A(n13384), .ZN(n13385) );
  AND2_X1 U16797 ( .A1(n19274), .A2(n13388), .ZN(n19221) );
  NAND2_X1 U16798 ( .A1(n19274), .A2(n13389), .ZN(n14244) );
  INV_X1 U16799 ( .A(n14244), .ZN(n13390) );
  OAI22_X1 U16800 ( .A1(n19229), .A2(n19199), .B1(n19274), .B2(n13658), .ZN(
        n13393) );
  NOR2_X1 U16801 ( .A1(n19207), .A2(n19199), .ZN(n13918) );
  AOI211_X1 U16802 ( .C1(n19207), .C2(n19199), .A(n13918), .B(n19258), .ZN(
        n13392) );
  AOI211_X1 U16803 ( .C1(n19220), .C2(n19266), .A(n13393), .B(n13392), .ZN(
        n13394) );
  INV_X1 U16804 ( .A(n13394), .ZN(P2_U2919) );
  AND2_X1 U16805 ( .A1(n20769), .A2(n16442), .ZN(n13418) );
  INV_X1 U16806 ( .A(n13637), .ZN(n13395) );
  AOI211_X1 U16807 ( .C1(P1_MEMORYFETCH_REG_SCAN_IN), .C2(n13396), .A(n13418), 
        .B(n13395), .ZN(n13397) );
  INV_X1 U16808 ( .A(n13397), .ZN(P1_U2801) );
  INV_X1 U16809 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n13481) );
  AOI22_X1 U16810 ( .A1(n20057), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n19303), 
        .B2(P2_DATAO_REG_18__SCAN_IN), .ZN(n13398) );
  OAI21_X1 U16811 ( .B1(n13481), .B2(n19276), .A(n13398), .ZN(P2_U2933) );
  INV_X1 U16812 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n13504) );
  AOI22_X1 U16813 ( .A1(n20057), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(n19303), 
        .B2(P2_DATAO_REG_26__SCAN_IN), .ZN(n13399) );
  OAI21_X1 U16814 ( .B1(n13504), .B2(n19276), .A(n13399), .ZN(P2_U2925) );
  INV_X1 U16815 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n13492) );
  AOI22_X1 U16816 ( .A1(n20057), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n19303), 
        .B2(P2_DATAO_REG_20__SCAN_IN), .ZN(n13400) );
  OAI21_X1 U16817 ( .B1(n13492), .B2(n19276), .A(n13400), .ZN(P2_U2931) );
  INV_X1 U16818 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n13402) );
  AOI22_X1 U16819 ( .A1(n20057), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n19303), 
        .B2(P2_DATAO_REG_17__SCAN_IN), .ZN(n13401) );
  OAI21_X1 U16820 ( .B1(n13402), .B2(n19276), .A(n13401), .ZN(P2_U2934) );
  INV_X1 U16821 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n13485) );
  AOI22_X1 U16822 ( .A1(n20057), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(n19303), 
        .B2(P2_DATAO_REG_24__SCAN_IN), .ZN(n13403) );
  OAI21_X1 U16823 ( .B1(n13485), .B2(n19276), .A(n13403), .ZN(P2_U2927) );
  INV_X1 U16824 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n15709) );
  AOI22_X1 U16825 ( .A1(n20057), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(n19303), 
        .B2(P2_DATAO_REG_27__SCAN_IN), .ZN(n13404) );
  OAI21_X1 U16826 ( .B1(n15709), .B2(n19276), .A(n13404), .ZN(P2_U2924) );
  INV_X1 U16827 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n13406) );
  AOI22_X1 U16828 ( .A1(n20057), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n19303), 
        .B2(P2_DATAO_REG_23__SCAN_IN), .ZN(n13405) );
  OAI21_X1 U16829 ( .B1(n13406), .B2(n19276), .A(n13405), .ZN(P2_U2928) );
  INV_X1 U16830 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n13408) );
  AOI22_X1 U16831 ( .A1(n20057), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(n19303), 
        .B2(P2_DATAO_REG_25__SCAN_IN), .ZN(n13407) );
  OAI21_X1 U16832 ( .B1(n13408), .B2(n19276), .A(n13407), .ZN(P2_U2926) );
  INV_X1 U16833 ( .A(P2_EAX_REG_30__SCAN_IN), .ZN(n13490) );
  AOI22_X1 U16834 ( .A1(n20057), .A2(P2_UWORD_REG_14__SCAN_IN), .B1(n19303), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .ZN(n13409) );
  OAI21_X1 U16835 ( .B1(n13490), .B2(n19276), .A(n13409), .ZN(P2_U2921) );
  INV_X1 U16836 ( .A(P2_EAX_REG_29__SCAN_IN), .ZN(n15698) );
  AOI22_X1 U16837 ( .A1(n20057), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(n19303), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n13410) );
  OAI21_X1 U16838 ( .B1(n15698), .B2(n19276), .A(n13410), .ZN(P2_U2922) );
  INV_X1 U16839 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n13634) );
  AOI22_X1 U16840 ( .A1(n20057), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n19303), 
        .B2(P2_DATAO_REG_19__SCAN_IN), .ZN(n13411) );
  OAI21_X1 U16841 ( .B1(n13634), .B2(n19276), .A(n13411), .ZN(P2_U2932) );
  INV_X1 U16842 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n13500) );
  AOI22_X1 U16843 ( .A1(n20057), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(n19303), 
        .B2(P2_DATAO_REG_28__SCAN_IN), .ZN(n13412) );
  OAI21_X1 U16844 ( .B1(n13500), .B2(n19276), .A(n13412), .ZN(P2_U2923) );
  NAND2_X1 U16845 ( .A1(n13582), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13413) );
  INV_X1 U16846 ( .A(n13584), .ZN(n19716) );
  NOR2_X1 U16847 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19368) );
  INV_X1 U16848 ( .A(n19368), .ZN(n19637) );
  NAND2_X1 U16849 ( .A1(n19716), .A2(n19637), .ZN(n14315) );
  NAND2_X1 U16850 ( .A1(n13413), .A2(n19579), .ZN(n13414) );
  NOR2_X1 U16851 ( .A1(n15661), .A2(n19354), .ZN(n13416) );
  AOI21_X1 U16852 ( .B1(P2_EBX_REG_1__SCAN_IN), .B2(n15661), .A(n13416), .ZN(
        n13417) );
  OAI21_X1 U16853 ( .B1(n20026), .B2(n15694), .A(n13417), .ZN(P2_U2886) );
  OAI21_X1 U16854 ( .B1(n13418), .B2(P1_READREQUEST_REG_SCAN_IN), .A(n13840), 
        .ZN(n13419) );
  OAI21_X1 U16855 ( .B1(n13420), .B2(n13840), .A(n13419), .ZN(P1_U3487) );
  AOI22_X1 U16856 ( .A1(n14302), .A2(BUF1_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n14303), .ZN(n13617) );
  INV_X1 U16857 ( .A(n13617), .ZN(n19403) );
  NOR3_X4 U16858 ( .A1(n13421), .A2(n9839), .A3(n19925), .ZN(n13615) );
  INV_X1 U16859 ( .A(n13421), .ZN(n13422) );
  AOI222_X1 U16860 ( .A1(n19403), .A2(n13615), .B1(P2_EAX_REG_5__SCAN_IN), 
        .B2(n13527), .C1(n13526), .C2(P2_LWORD_REG_5__SCAN_IN), .ZN(n13423) );
  INV_X1 U16861 ( .A(n13423), .ZN(P2_U2972) );
  AOI22_X1 U16862 ( .A1(n14302), .A2(BUF1_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n14303), .ZN(n13424) );
  INV_X1 U16863 ( .A(n13424), .ZN(n14306) );
  AOI222_X1 U16864 ( .A1(n14306), .A2(n13615), .B1(n13527), .B2(
        P2_EAX_REG_1__SCAN_IN), .C1(n13526), .C2(P2_LWORD_REG_1__SCAN_IN), 
        .ZN(n13425) );
  INV_X1 U16865 ( .A(n13425), .ZN(P2_U2968) );
  AOI22_X1 U16866 ( .A1(P2_LWORD_REG_13__SCAN_IN), .A2(n13526), .B1(n13527), 
        .B2(P2_EAX_REG_13__SCAN_IN), .ZN(n13429) );
  INV_X1 U16867 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n15049) );
  OR2_X1 U16868 ( .A1(n14303), .A2(n15049), .ZN(n13427) );
  NAND2_X1 U16869 ( .A1(n14303), .A2(BUF2_REG_13__SCAN_IN), .ZN(n13426) );
  AND2_X1 U16870 ( .A1(n13427), .A2(n13426), .ZN(n19236) );
  INV_X1 U16871 ( .A(n19236), .ZN(n13428) );
  NAND2_X1 U16872 ( .A1(n13615), .A2(n13428), .ZN(n13439) );
  NAND2_X1 U16873 ( .A1(n13429), .A2(n13439), .ZN(P2_U2980) );
  AOI22_X1 U16874 ( .A1(P2_LWORD_REG_7__SCAN_IN), .A2(n13447), .B1(n13527), 
        .B2(P2_EAX_REG_7__SCAN_IN), .ZN(n13430) );
  AOI22_X1 U16875 ( .A1(n14302), .A2(BUF1_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n14303), .ZN(n19417) );
  INV_X1 U16876 ( .A(n19417), .ZN(n15737) );
  NAND2_X1 U16877 ( .A1(n13615), .A2(n15737), .ZN(n13445) );
  NAND2_X1 U16878 ( .A1(n13430), .A2(n13445), .ZN(P2_U2974) );
  AOI22_X1 U16879 ( .A1(P2_UWORD_REG_11__SCAN_IN), .A2(n13447), .B1(n13527), 
        .B2(P2_EAX_REG_27__SCAN_IN), .ZN(n13434) );
  INV_X1 U16880 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n16673) );
  OR2_X1 U16881 ( .A1(n14303), .A2(n16673), .ZN(n13432) );
  NAND2_X1 U16882 ( .A1(n14303), .A2(BUF2_REG_11__SCAN_IN), .ZN(n13431) );
  AND2_X1 U16883 ( .A1(n13432), .A2(n13431), .ZN(n19242) );
  INV_X1 U16884 ( .A(n19242), .ZN(n13433) );
  NAND2_X1 U16885 ( .A1(n13615), .A2(n13433), .ZN(n13443) );
  NAND2_X1 U16886 ( .A1(n13434), .A2(n13443), .ZN(P2_U2963) );
  AOI22_X1 U16887 ( .A1(P2_UWORD_REG_9__SCAN_IN), .A2(n13447), .B1(n13527), 
        .B2(P2_EAX_REG_25__SCAN_IN), .ZN(n13437) );
  INV_X1 U16888 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n14495) );
  OR2_X1 U16889 ( .A1(n14303), .A2(n14495), .ZN(n13436) );
  NAND2_X1 U16890 ( .A1(n14303), .A2(BUF2_REG_9__SCAN_IN), .ZN(n13435) );
  AND2_X1 U16891 ( .A1(n13436), .A2(n13435), .ZN(n19247) );
  INV_X1 U16892 ( .A(n19247), .ZN(n15725) );
  NAND2_X1 U16893 ( .A1(n13615), .A2(n15725), .ZN(n13448) );
  NAND2_X1 U16894 ( .A1(n13437), .A2(n13448), .ZN(P2_U2961) );
  AOI22_X1 U16895 ( .A1(P2_LWORD_REG_6__SCAN_IN), .A2(n13447), .B1(n13527), 
        .B2(P2_EAX_REG_6__SCAN_IN), .ZN(n13438) );
  INV_X1 U16896 ( .A(BUF1_REG_6__SCAN_IN), .ZN(n16680) );
  INV_X1 U16897 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n18410) );
  AOI22_X1 U16898 ( .A1(n14302), .A2(n16680), .B1(n18410), .B2(n14303), .ZN(
        n19409) );
  NAND2_X1 U16899 ( .A1(n13615), .A2(n19409), .ZN(n13441) );
  NAND2_X1 U16900 ( .A1(n13438), .A2(n13441), .ZN(P2_U2973) );
  AOI22_X1 U16901 ( .A1(P2_UWORD_REG_13__SCAN_IN), .A2(n13526), .B1(n13527), 
        .B2(P2_EAX_REG_29__SCAN_IN), .ZN(n13440) );
  NAND2_X1 U16902 ( .A1(n13440), .A2(n13439), .ZN(P2_U2965) );
  AOI22_X1 U16903 ( .A1(P2_UWORD_REG_6__SCAN_IN), .A2(n13447), .B1(n13527), 
        .B2(P2_EAX_REG_22__SCAN_IN), .ZN(n13442) );
  NAND2_X1 U16904 ( .A1(n13442), .A2(n13441), .ZN(P2_U2958) );
  AOI22_X1 U16905 ( .A1(P2_LWORD_REG_11__SCAN_IN), .A2(n13447), .B1(n13527), 
        .B2(P2_EAX_REG_11__SCAN_IN), .ZN(n13444) );
  NAND2_X1 U16906 ( .A1(n13444), .A2(n13443), .ZN(P2_U2978) );
  AOI22_X1 U16907 ( .A1(P2_UWORD_REG_7__SCAN_IN), .A2(n13447), .B1(n13527), 
        .B2(P2_EAX_REG_23__SCAN_IN), .ZN(n13446) );
  NAND2_X1 U16908 ( .A1(n13446), .A2(n13445), .ZN(P2_U2959) );
  AOI22_X1 U16909 ( .A1(P2_LWORD_REG_9__SCAN_IN), .A2(n13447), .B1(n13527), 
        .B2(P2_EAX_REG_9__SCAN_IN), .ZN(n13449) );
  NAND2_X1 U16910 ( .A1(n13449), .A2(n13448), .ZN(P2_U2976) );
  AOI22_X1 U16911 ( .A1(P2_LWORD_REG_2__SCAN_IN), .A2(n13526), .B1(n13527), 
        .B2(P2_EAX_REG_2__SCAN_IN), .ZN(n13450) );
  INV_X1 U16912 ( .A(BUF1_REG_2__SCAN_IN), .ZN(n16687) );
  INV_X1 U16913 ( .A(BUF2_REG_2__SCAN_IN), .ZN(n18394) );
  AOI22_X1 U16914 ( .A1(n14302), .A2(n16687), .B1(n18394), .B2(n14303), .ZN(
        n19381) );
  NAND2_X1 U16915 ( .A1(n13615), .A2(n19381), .ZN(n13480) );
  NAND2_X1 U16916 ( .A1(n13450), .A2(n13480), .ZN(P2_U2969) );
  OAI21_X1 U16917 ( .B1(n13453), .B2(n13452), .A(n13451), .ZN(n20031) );
  XNOR2_X1 U16918 ( .A(n20029), .B(n20031), .ZN(n13919) );
  XOR2_X1 U16919 ( .A(n13918), .B(n13919), .Z(n13456) );
  AOI22_X1 U16920 ( .A1(n19265), .A2(n20031), .B1(P2_EAX_REG_1__SCAN_IN), .B2(
        n19257), .ZN(n13455) );
  NAND2_X1 U16921 ( .A1(n19266), .A2(n14306), .ZN(n13454) );
  OAI211_X1 U16922 ( .C1(n13456), .C2(n19258), .A(n13455), .B(n13454), .ZN(
        P2_U2918) );
  NAND2_X1 U16923 ( .A1(n13791), .A2(n13518), .ZN(n13457) );
  NAND2_X1 U16924 ( .A1(n13457), .A2(n12757), .ZN(n13766) );
  NOR2_X1 U16925 ( .A1(n13521), .A2(n13458), .ZN(n13770) );
  NAND2_X1 U16926 ( .A1(n16210), .A2(n13770), .ZN(n13546) );
  OAI211_X1 U16927 ( .C1(n13839), .C2(n11640), .A(n13766), .B(n13546), .ZN(
        n13459) );
  NOR2_X1 U16928 ( .A1(n13460), .A2(n13459), .ZN(n13468) );
  INV_X1 U16929 ( .A(n13462), .ZN(n13463) );
  AOI21_X1 U16930 ( .B1(n15468), .B2(n13463), .A(n16223), .ZN(n13466) );
  OAI211_X1 U16931 ( .C1(n13466), .C2(n13465), .A(n16193), .B(n21010), .ZN(
        n13467) );
  NAND2_X1 U16932 ( .A1(n13468), .A2(n13467), .ZN(n16172) );
  NAND2_X1 U16933 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n13963), .ZN(n16443) );
  INV_X1 U16934 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n20089) );
  NOR2_X1 U16935 ( .A1(n16443), .A2(n20089), .ZN(n13469) );
  AOI21_X1 U16936 ( .B1(n16172), .B2(n13768), .A(n13469), .ZN(n13476) );
  NAND2_X1 U16937 ( .A1(n20310), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n13470) );
  INV_X1 U16938 ( .A(n15484), .ZN(n15477) );
  INV_X1 U16939 ( .A(n20460), .ZN(n20729) );
  NOR2_X1 U16940 ( .A1(n13471), .A2(n20729), .ZN(n13472) );
  XNOR2_X1 U16941 ( .A(n13472), .B(n13478), .ZN(n20153) );
  INV_X1 U16942 ( .A(n13474), .ZN(n13475) );
  NAND2_X1 U16943 ( .A1(n20153), .A2(n13475), .ZN(n13962) );
  INV_X1 U16944 ( .A(n20080), .ZN(n15482) );
  OR3_X1 U16945 ( .A1(n13962), .A2(n13476), .A3(n15482), .ZN(n13477) );
  OAI21_X1 U16946 ( .B1(n13478), .B2(n15477), .A(n13477), .ZN(P1_U3468) );
  NAND2_X1 U16947 ( .A1(n13526), .A2(P2_UWORD_REG_2__SCAN_IN), .ZN(n13479) );
  OAI211_X1 U16948 ( .C1(n13481), .C2(n13657), .A(n13480), .B(n13479), .ZN(
        P2_U2954) );
  NAND2_X1 U16949 ( .A1(n14303), .A2(BUF2_REG_8__SCAN_IN), .ZN(n13483) );
  INV_X1 U16950 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n16677) );
  OR2_X1 U16951 ( .A1(n14303), .A2(n16677), .ZN(n13482) );
  NAND2_X1 U16952 ( .A1(n13483), .A2(n13482), .ZN(n19249) );
  NAND2_X1 U16953 ( .A1(n13615), .A2(n19249), .ZN(n13496) );
  NAND2_X1 U16954 ( .A1(n13526), .A2(P2_UWORD_REG_8__SCAN_IN), .ZN(n13484) );
  OAI211_X1 U16955 ( .C1(n13485), .C2(n13657), .A(n13496), .B(n13484), .ZN(
        P2_U2960) );
  NAND2_X1 U16956 ( .A1(n14303), .A2(BUF2_REG_14__SCAN_IN), .ZN(n13488) );
  OR2_X1 U16957 ( .A1(n14303), .A2(n13486), .ZN(n13487) );
  NAND2_X1 U16958 ( .A1(n13488), .A2(n13487), .ZN(n19232) );
  NAND2_X1 U16959 ( .A1(n13615), .A2(n19232), .ZN(n13506) );
  NAND2_X1 U16960 ( .A1(n13526), .A2(P2_UWORD_REG_14__SCAN_IN), .ZN(n13489) );
  OAI211_X1 U16961 ( .C1(n13490), .C2(n13657), .A(n13506), .B(n13489), .ZN(
        P2_U2966) );
  INV_X1 U16962 ( .A(BUF1_REG_4__SCAN_IN), .ZN(n16683) );
  INV_X1 U16963 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n18402) );
  AOI22_X1 U16964 ( .A1(n14302), .A2(n16683), .B1(n18402), .B2(n14303), .ZN(
        n19396) );
  NAND2_X1 U16965 ( .A1(n13615), .A2(n19396), .ZN(n13494) );
  NAND2_X1 U16966 ( .A1(n13526), .A2(P2_UWORD_REG_4__SCAN_IN), .ZN(n13491) );
  OAI211_X1 U16967 ( .C1(n13492), .C2(n13657), .A(n13494), .B(n13491), .ZN(
        P2_U2956) );
  INV_X1 U16968 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n19301) );
  NAND2_X1 U16969 ( .A1(n13526), .A2(P2_LWORD_REG_4__SCAN_IN), .ZN(n13493) );
  OAI211_X1 U16970 ( .C1(n19301), .C2(n13657), .A(n13494), .B(n13493), .ZN(
        P2_U2971) );
  INV_X1 U16971 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n19293) );
  NAND2_X1 U16972 ( .A1(n13526), .A2(P2_LWORD_REG_8__SCAN_IN), .ZN(n13495) );
  OAI211_X1 U16973 ( .C1(n19293), .C2(n13657), .A(n13496), .B(n13495), .ZN(
        P2_U2975) );
  NAND2_X1 U16974 ( .A1(n14303), .A2(BUF2_REG_12__SCAN_IN), .ZN(n13498) );
  INV_X1 U16975 ( .A(BUF1_REG_12__SCAN_IN), .ZN(n16671) );
  OR2_X1 U16976 ( .A1(n14303), .A2(n16671), .ZN(n13497) );
  NAND2_X1 U16977 ( .A1(n13498), .A2(n13497), .ZN(n19239) );
  NAND2_X1 U16978 ( .A1(n13615), .A2(n19239), .ZN(n13508) );
  NAND2_X1 U16979 ( .A1(n13526), .A2(P2_UWORD_REG_12__SCAN_IN), .ZN(n13499) );
  OAI211_X1 U16980 ( .C1(n13500), .C2(n13657), .A(n13508), .B(n13499), .ZN(
        P2_U2964) );
  NAND2_X1 U16981 ( .A1(n14303), .A2(BUF2_REG_10__SCAN_IN), .ZN(n13502) );
  INV_X1 U16982 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n14491) );
  OR2_X1 U16983 ( .A1(n14303), .A2(n14491), .ZN(n13501) );
  NAND2_X1 U16984 ( .A1(n13502), .A2(n13501), .ZN(n19244) );
  NAND2_X1 U16985 ( .A1(n13615), .A2(n19244), .ZN(n13510) );
  NAND2_X1 U16986 ( .A1(n13526), .A2(P2_UWORD_REG_10__SCAN_IN), .ZN(n13503) );
  OAI211_X1 U16987 ( .C1(n13504), .C2(n13657), .A(n13510), .B(n13503), .ZN(
        P2_U2962) );
  INV_X1 U16988 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n19282) );
  NAND2_X1 U16989 ( .A1(n13526), .A2(P2_LWORD_REG_14__SCAN_IN), .ZN(n13505) );
  OAI211_X1 U16990 ( .C1(n19282), .C2(n13657), .A(n13506), .B(n13505), .ZN(
        P2_U2981) );
  INV_X1 U16991 ( .A(P2_LWORD_REG_12__SCAN_IN), .ZN(n21221) );
  NAND2_X1 U16992 ( .A1(n13527), .A2(P2_EAX_REG_12__SCAN_IN), .ZN(n13507) );
  OAI211_X1 U16993 ( .C1(n13655), .C2(n21221), .A(n13508), .B(n13507), .ZN(
        P2_U2979) );
  INV_X1 U16994 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n19289) );
  NAND2_X1 U16995 ( .A1(n13526), .A2(P2_LWORD_REG_10__SCAN_IN), .ZN(n13509) );
  OAI211_X1 U16996 ( .C1(n19289), .C2(n13657), .A(n13510), .B(n13509), .ZN(
        P2_U2977) );
  INV_X1 U16997 ( .A(n20422), .ZN(n13967) );
  INV_X1 U16998 ( .A(n13839), .ZN(n13512) );
  AND2_X1 U16999 ( .A1(n13512), .A2(n11598), .ZN(n13776) );
  INV_X1 U17000 ( .A(n13776), .ZN(n13513) );
  NAND3_X1 U17001 ( .A1(n10040), .A2(n13514), .A3(n13513), .ZN(n13515) );
  NOR2_X1 U17002 ( .A1(n13462), .A2(n13515), .ZN(n13520) );
  OAI21_X1 U17003 ( .B1(n13516), .B2(n13943), .A(n16201), .ZN(n13517) );
  AND2_X1 U17004 ( .A1(n13518), .A2(n13517), .ZN(n13778) );
  AND4_X1 U17005 ( .A1(n13474), .A2(n13520), .A3(n13778), .A4(n13519), .ZN(
        n13944) );
  OAI22_X1 U17006 ( .A1(n13967), .A2(n13944), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n13521), .ZN(n16174) );
  OAI22_X1 U17007 ( .A1(n16442), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n15481), .ZN(n13522) );
  AOI21_X1 U17008 ( .B1(n16174), .B2(n20080), .A(n13522), .ZN(n13525) );
  AOI21_X1 U17009 ( .B1(n16175), .B2(n20080), .A(n15484), .ZN(n13524) );
  OAI22_X1 U17010 ( .A1(n13525), .A2(n15484), .B1(n13524), .B2(n13523), .ZN(
        P1_U3474) );
  AOI222_X1 U17011 ( .A1(P2_EAX_REG_17__SCAN_IN), .A2(n13527), .B1(n14306), 
        .B2(n13615), .C1(n13526), .C2(P2_UWORD_REG_1__SCAN_IN), .ZN(n13528) );
  INV_X1 U17012 ( .A(n13528), .ZN(P2_U2953) );
  INV_X1 U17013 ( .A(n13529), .ZN(n13532) );
  OAI21_X1 U17014 ( .B1(n13532), .B2(n13531), .A(n13530), .ZN(n14015) );
  INV_X1 U17015 ( .A(n13533), .ZN(n13536) );
  INV_X1 U17016 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n13535) );
  AOI21_X1 U17017 ( .B1(n13536), .B2(n13535), .A(n13534), .ZN(n20290) );
  INV_X1 U17018 ( .A(P1_REIP_REG_0__SCAN_IN), .ZN(n13863) );
  OAI21_X1 U17019 ( .B1(n20242), .B2(n13537), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13538) );
  OAI21_X1 U17020 ( .B1(n13863), .B2(n20256), .A(n13538), .ZN(n13539) );
  AOI21_X1 U17021 ( .B1(n20290), .B2(n20248), .A(n13539), .ZN(n13540) );
  OAI21_X1 U17022 ( .B1(n20306), .B2(n14015), .A(n13540), .ZN(P1_U2999) );
  OAI21_X1 U17023 ( .B1(n13542), .B2(n13541), .A(n13729), .ZN(n14010) );
  NAND2_X1 U17024 ( .A1(n13546), .A2(n13545), .ZN(n13547) );
  OR2_X1 U17025 ( .A1(n13549), .A2(n13548), .ZN(n13550) );
  AND2_X1 U17026 ( .A1(n13551), .A2(n13550), .ZN(n13841) );
  INV_X1 U17027 ( .A(n13841), .ZN(n20281) );
  AOI22_X1 U17028 ( .A1(n20171), .A2(n20281), .B1(n15032), .B2(
        P1_EBX_REG_1__SCAN_IN), .ZN(n13552) );
  OAI21_X1 U17029 ( .B1(n14010), .B2(n9828), .A(n13552), .ZN(P1_U2871) );
  XNOR2_X1 U17030 ( .A(n13554), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13556) );
  INV_X1 U17031 ( .A(n13770), .ZN(n16188) );
  NAND2_X1 U17032 ( .A1(n13792), .A2(n16188), .ZN(n13949) );
  XNOR2_X1 U17033 ( .A(n15472), .B(n13561), .ZN(n13559) );
  INV_X1 U17034 ( .A(n13559), .ZN(n13555) );
  AOI22_X1 U17035 ( .A1(n16175), .A2(n13556), .B1(n13949), .B2(n13555), .ZN(
        n13558) );
  NAND3_X1 U17036 ( .A1(n13944), .A2(n13943), .A3(n13559), .ZN(n13557) );
  OAI211_X1 U17037 ( .C1(n13553), .C2(n13944), .A(n13558), .B(n13557), .ZN(
        n13941) );
  NOR2_X1 U17038 ( .A1(n16442), .A2(n13535), .ZN(n15474) );
  INV_X1 U17039 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n21115) );
  AOI22_X1 U17040 ( .A1(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n20286), .B2(n21115), .ZN(
        n15471) );
  INV_X1 U17041 ( .A(n15481), .ZN(n13560) );
  AOI222_X1 U17042 ( .A1(n13941), .A2(n20080), .B1(n15474), .B2(n15471), .C1(
        n13560), .C2(n13559), .ZN(n13562) );
  MUX2_X1 U17043 ( .A(n13562), .B(n13561), .S(n15484), .Z(n13563) );
  INV_X1 U17044 ( .A(n13563), .ZN(P1_U3472) );
  NAND2_X1 U17045 ( .A1(n13564), .A2(n13587), .ZN(n13568) );
  NAND2_X1 U17046 ( .A1(n19716), .A2(n20023), .ZN(n13565) );
  NOR2_X1 U17047 ( .A1(n20023), .A2(n20033), .ZN(n19853) );
  NAND2_X1 U17048 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19853), .ZN(
        n19367) );
  NAND2_X1 U17049 ( .A1(n13565), .A2(n19367), .ZN(n14316) );
  NOR2_X1 U17050 ( .A1(n14316), .A2(n20002), .ZN(n13566) );
  AOI21_X1 U17051 ( .B1(n13582), .B2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n13566), .ZN(n13567) );
  INV_X1 U17052 ( .A(n13570), .ZN(n13571) );
  NOR2_X1 U17053 ( .A1(n16107), .A2(n13571), .ZN(n13572) );
  INV_X1 U17054 ( .A(n19364), .ZN(n20018) );
  INV_X1 U17055 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n14197) );
  MUX2_X1 U17056 ( .A(n14805), .B(n14197), .S(n15667), .Z(n13575) );
  OAI21_X1 U17057 ( .B1(n20018), .B2(n15694), .A(n13575), .ZN(P2_U2885) );
  INV_X1 U17058 ( .A(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13846) );
  INV_X1 U17059 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n13576) );
  OAI22_X1 U17060 ( .A1(n15228), .A2(n13846), .B1(n20256), .B2(n13576), .ZN(
        n13577) );
  AOI21_X1 U17061 ( .B1(n16316), .B2(n13846), .A(n13577), .ZN(n13581) );
  OR2_X1 U17062 ( .A1(n13578), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n20279) );
  NAND3_X1 U17063 ( .A1(n20279), .A2(n13579), .A3(n20248), .ZN(n13580) );
  OAI211_X1 U17064 ( .C1(n14010), .C2(n20306), .A(n13581), .B(n13580), .ZN(
        P1_U2998) );
  NAND2_X1 U17065 ( .A1(n13582), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13586) );
  NAND2_X1 U17066 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n20017), .ZN(
        n19539) );
  INV_X1 U17067 ( .A(n19539), .ZN(n13583) );
  AND2_X1 U17068 ( .A1(n19367), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n13585) );
  OAI21_X1 U17069 ( .B1(n19643), .B2(n13585), .A(n20006), .ZN(n14341) );
  NAND2_X1 U17070 ( .A1(n14723), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n13593) );
  NAND3_X1 U17071 ( .A1(n13619), .A2(n13624), .A3(n13588), .ZN(n13598) );
  NAND3_X1 U17072 ( .A1(n13624), .A2(n13589), .A3(n13569), .ZN(n13597) );
  INV_X1 U17073 ( .A(n13590), .ZN(n13591) );
  NAND2_X1 U17074 ( .A1(n13591), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n13596) );
  INV_X1 U17075 ( .A(n13592), .ZN(n13595) );
  INV_X1 U17076 ( .A(n13593), .ZN(n13594) );
  NAND2_X1 U17077 ( .A1(n13595), .A2(n13594), .ZN(n13623) );
  INV_X1 U17078 ( .A(n14723), .ZN(n13600) );
  INV_X1 U17079 ( .A(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13599) );
  NOR2_X1 U17080 ( .A1(n13600), .A2(n13599), .ZN(n13608) );
  NAND2_X1 U17081 ( .A1(n13702), .A2(n13608), .ZN(n13670) );
  XOR2_X1 U17082 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B(n13670), .Z(n13607)
         );
  NAND2_X1 U17083 ( .A1(n13601), .A2(n13612), .ZN(n13604) );
  INV_X1 U17084 ( .A(n13602), .ZN(n13603) );
  AND2_X1 U17085 ( .A1(n13604), .A2(n13603), .ZN(n19174) );
  NOR2_X1 U17086 ( .A1(n14287), .A2(n10544), .ZN(n13605) );
  AOI21_X1 U17087 ( .B1(n19174), .B2(n14287), .A(n13605), .ZN(n13606) );
  OAI21_X1 U17088 ( .B1(n13607), .B2(n15694), .A(n13606), .ZN(P2_U2882) );
  OAI21_X1 U17089 ( .B1(n13702), .B2(n13608), .A(n13670), .ZN(n19259) );
  NAND2_X1 U17090 ( .A1(n15667), .A2(P2_EBX_REG_4__SCAN_IN), .ZN(n13614) );
  OR2_X1 U17091 ( .A1(n13610), .A2(n13609), .ZN(n13611) );
  AND2_X1 U17092 ( .A1(n13612), .A2(n13611), .ZN(n19316) );
  NAND2_X1 U17093 ( .A1(n19316), .A2(n14287), .ZN(n13613) );
  OAI211_X1 U17094 ( .C1(n19259), .C2(n15694), .A(n13614), .B(n13613), .ZN(
        P2_U2883) );
  INV_X1 U17095 ( .A(n13615), .ZN(n13654) );
  OAI222_X1 U17096 ( .A1(n13654), .A2(n13617), .B1(n21305), .B2(n13655), .C1(
        n13657), .C2(n13616), .ZN(P2_U2957) );
  AOI22_X1 U17097 ( .A1(n14302), .A2(BUF1_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n14303), .ZN(n19230) );
  INV_X1 U17098 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n19280) );
  INV_X1 U17099 ( .A(P2_LWORD_REG_15__SCAN_IN), .ZN(n21222) );
  OAI222_X1 U17100 ( .A1(n13654), .A2(n19230), .B1(n13657), .B2(n19280), .C1(
        n21222), .C2(n13655), .ZN(P2_U2982) );
  OAI222_X1 U17101 ( .A1(n13654), .A2(n13653), .B1(n13364), .B2(n13655), .C1(
        n13657), .C2(n13618), .ZN(P2_U2952) );
  INV_X1 U17102 ( .A(n13619), .ZN(n13622) );
  CLKBUF_X1 U17103 ( .A(n13627), .Z(n14070) );
  INV_X1 U17104 ( .A(n14070), .ZN(n13893) );
  MUX2_X1 U17105 ( .A(n13893), .B(n13628), .S(n15667), .Z(n13629) );
  OAI21_X1 U17106 ( .B1(n19431), .B2(n15694), .A(n13629), .ZN(P2_U2884) );
  OR2_X1 U17107 ( .A1(n13630), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13632) );
  AND2_X1 U17108 ( .A1(n13632), .A2(n13631), .ZN(n13861) );
  INV_X1 U17109 ( .A(n13861), .ZN(n20291) );
  OAI222_X1 U17110 ( .A1(n20291), .A2(n20175), .B1(n13633), .B2(n20182), .C1(
        n14015), .C2(n9828), .ZN(P1_U2872) );
  AOI22_X1 U17111 ( .A1(n14302), .A2(BUF1_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n14303), .ZN(n14382) );
  INV_X1 U17112 ( .A(P2_UWORD_REG_3__SCAN_IN), .ZN(n13635) );
  OAI222_X1 U17113 ( .A1(n14382), .A2(n13654), .B1(n13635), .B2(n13655), .C1(
        n13657), .C2(n13634), .ZN(P2_U2955) );
  INV_X1 U17114 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n13641) );
  NAND2_X1 U17115 ( .A1(n16193), .A2(n13768), .ZN(n13636) );
  INV_X1 U17116 ( .A(n16223), .ZN(n13638) );
  INV_X1 U17117 ( .A(n13963), .ZN(n16438) );
  NOR2_X4 U17118 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n16438), .ZN(n13910) );
  NOR2_X4 U17119 ( .A1(n20187), .A2(n13910), .ZN(n20204) );
  AOI22_X1 U17120 ( .A1(P1_UWORD_REG_8__SCAN_IN), .A2(n13910), .B1(n20204), 
        .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n13640) );
  OAI21_X1 U17121 ( .B1(n13641), .B2(n13912), .A(n13640), .ZN(P1_U2912) );
  INV_X1 U17122 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n13643) );
  AOI22_X1 U17123 ( .A1(P1_UWORD_REG_12__SCAN_IN), .A2(n13910), .B1(n20204), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n13642) );
  OAI21_X1 U17124 ( .B1(n13643), .B2(n13912), .A(n13642), .ZN(P1_U2908) );
  AOI22_X1 U17125 ( .A1(P1_UWORD_REG_10__SCAN_IN), .A2(n13910), .B1(n20204), 
        .B2(P1_DATAO_REG_26__SCAN_IN), .ZN(n13644) );
  OAI21_X1 U17126 ( .B1(n15059), .B2(n13912), .A(n13644), .ZN(P1_U2910) );
  INV_X1 U17127 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n13646) );
  AOI22_X1 U17128 ( .A1(P1_UWORD_REG_9__SCAN_IN), .A2(n13910), .B1(n20204), 
        .B2(P1_DATAO_REG_25__SCAN_IN), .ZN(n13645) );
  OAI21_X1 U17129 ( .B1(n13646), .B2(n13912), .A(n13645), .ZN(P1_U2911) );
  INV_X1 U17130 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n13648) );
  AOI22_X1 U17131 ( .A1(P1_UWORD_REG_13__SCAN_IN), .A2(n13910), .B1(n20204), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n13647) );
  OAI21_X1 U17132 ( .B1(n13648), .B2(n13912), .A(n13647), .ZN(P1_U2907) );
  INV_X1 U17133 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n21309) );
  AOI22_X1 U17134 ( .A1(P1_UWORD_REG_11__SCAN_IN), .A2(n13910), .B1(n20204), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n13649) );
  OAI21_X1 U17135 ( .B1(n21309), .B2(n13912), .A(n13649), .ZN(P1_U2909) );
  AOI22_X1 U17136 ( .A1(P1_UWORD_REG_14__SCAN_IN), .A2(n13910), .B1(n20204), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .ZN(n13650) );
  OAI21_X1 U17137 ( .B1(n13022), .B2(n13912), .A(n13650), .ZN(P1_U2906) );
  INV_X1 U17138 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n13652) );
  INV_X1 U17139 ( .A(P2_LWORD_REG_3__SCAN_IN), .ZN(n13651) );
  OAI222_X1 U17140 ( .A1(n13652), .A2(n13657), .B1(n13651), .B2(n13655), .C1(
        n13654), .C2(n14382), .ZN(P2_U2970) );
  INV_X1 U17141 ( .A(P2_LWORD_REG_0__SCAN_IN), .ZN(n13656) );
  OAI222_X1 U17142 ( .A1(n13658), .A2(n13657), .B1(n13656), .B2(n13655), .C1(
        n13654), .C2(n13653), .ZN(P2_U2967) );
  AND2_X1 U17143 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13698) );
  INV_X1 U17144 ( .A(n13698), .ZN(n13659) );
  NOR2_X1 U17145 ( .A1(n13670), .A2(n13659), .ZN(n13721) );
  XNOR2_X1 U17146 ( .A(n13721), .B(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13667) );
  NAND2_X1 U17147 ( .A1(n13661), .A2(n13660), .ZN(n13664) );
  INV_X1 U17148 ( .A(n13662), .ZN(n13663) );
  NAND2_X1 U17149 ( .A1(n13664), .A2(n13663), .ZN(n19148) );
  INV_X1 U17150 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n13665) );
  MUX2_X1 U17151 ( .A(n19148), .B(n13665), .S(n15667), .Z(n13666) );
  OAI21_X1 U17152 ( .B1(n13667), .B2(n15694), .A(n13666), .ZN(P2_U2880) );
  OAI21_X1 U17153 ( .B1(n13668), .B2(n13602), .A(n13660), .ZN(n16546) );
  NOR2_X1 U17154 ( .A1(n13670), .A2(n13669), .ZN(n13672) );
  INV_X1 U17155 ( .A(n13721), .ZN(n13671) );
  OAI211_X1 U17156 ( .C1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .C2(n13672), .A(
        n13671), .B(n15685), .ZN(n13674) );
  NAND2_X1 U17157 ( .A1(n15667), .A2(P2_EBX_REG_6__SCAN_IN), .ZN(n13673) );
  OAI211_X1 U17158 ( .C1(n16546), .C2(n15661), .A(n13674), .B(n13673), .ZN(
        P2_U2881) );
  INV_X1 U17159 ( .A(n19431), .ZN(n20010) );
  INV_X1 U17160 ( .A(n14613), .ZN(n13685) );
  NAND2_X1 U17161 ( .A1(n14105), .A2(n14106), .ZN(n14076) );
  INV_X1 U17162 ( .A(n10435), .ZN(n13675) );
  NAND2_X1 U17163 ( .A1(n13675), .A2(n10144), .ZN(n14075) );
  AOI22_X1 U17164 ( .A1(n14076), .A2(n14075), .B1(n10436), .B2(n14090), .ZN(
        n13683) );
  INV_X1 U17165 ( .A(n14075), .ZN(n13680) );
  AND2_X1 U17166 ( .A1(n13677), .A2(n13676), .ZN(n14081) );
  NOR2_X1 U17167 ( .A1(n14081), .A2(n13678), .ZN(n13679) );
  AOI211_X1 U17168 ( .C1(n13681), .C2(n14090), .A(n13680), .B(n13679), .ZN(
        n13682) );
  MUX2_X1 U17169 ( .A(n13683), .B(n13682), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n13684) );
  OAI211_X1 U17170 ( .C1(n13893), .C2(n14074), .A(n13685), .B(n13684), .ZN(
        n14097) );
  AOI22_X1 U17171 ( .A1(n20010), .A2(n16589), .B1(n20005), .B2(n14097), .ZN(
        n13697) );
  NAND2_X1 U17172 ( .A1(n13686), .A2(n14113), .ZN(n13693) );
  INV_X1 U17173 ( .A(n13687), .ZN(n13691) );
  AND2_X1 U17174 ( .A1(n13689), .A2(n13688), .ZN(n13690) );
  OAI211_X1 U17175 ( .C1(n13693), .C2(n13692), .A(n13691), .B(n13690), .ZN(
        n14098) );
  INV_X1 U17176 ( .A(n14098), .ZN(n14120) );
  NAND2_X1 U17177 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n13694), .ZN(n16595) );
  INV_X1 U17178 ( .A(n16595), .ZN(n16226) );
  AOI22_X1 U17179 ( .A1(n16226), .A2(P2_FLUSH_REG_SCAN_IN), .B1(
        P2_STATE2_REG_3__SCAN_IN), .B2(n14298), .ZN(n13695) );
  OAI21_X1 U17180 ( .B1(n14120), .B2(n19040), .A(n13695), .ZN(n16160) );
  INV_X1 U17181 ( .A(n16160), .ZN(n16118) );
  NAND2_X1 U17182 ( .A1(n16118), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13696) );
  OAI21_X1 U17183 ( .B1(n13697), .B2(n16118), .A(n13696), .ZN(P2_U3596) );
  AND4_X1 U17184 ( .A1(n13722), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A3(
        P2_INSTQUEUE_REG_0__7__SCAN_IN), .A4(n13698), .ZN(n13700) );
  AND3_X1 U17185 ( .A1(n14723), .A2(n13700), .A3(n13699), .ZN(n13701) );
  INV_X1 U17186 ( .A(n13703), .ZN(n13706) );
  INV_X1 U17187 ( .A(n13704), .ZN(n13705) );
  OAI211_X1 U17188 ( .C1(n13706), .C2(n13705), .A(n15685), .B(n13813), .ZN(
        n13712) );
  INV_X1 U17189 ( .A(n13707), .ZN(n13708) );
  NAND2_X1 U17190 ( .A1(n13708), .A2(n9950), .ZN(n13710) );
  AND2_X1 U17191 ( .A1(n13710), .A2(n13709), .ZN(n16519) );
  NAND2_X1 U17192 ( .A1(n14287), .A2(n16519), .ZN(n13711) );
  OAI211_X1 U17193 ( .C1(n14287), .C2(n10175), .A(n13712), .B(n13711), .ZN(
        P2_U2877) );
  AND2_X2 U17194 ( .A1(n13808), .A2(n11633), .ZN(n20239) );
  AOI22_X1 U17195 ( .A1(n20239), .A2(P1_EAX_REG_4__SCAN_IN), .B1(n20238), .B2(
        P1_LWORD_REG_4__SCAN_IN), .ZN(n13715) );
  INV_X1 U17196 ( .A(DATAI_4_), .ZN(n13714) );
  NAND2_X1 U17197 ( .A1(n20303), .A2(BUF1_REG_4__SCAN_IN), .ZN(n13713) );
  OAI21_X1 U17198 ( .B1(n20303), .B2(n13714), .A(n13713), .ZN(n20335) );
  NAND2_X1 U17199 ( .A1(n20224), .A2(n20335), .ZN(n13719) );
  NAND2_X1 U17200 ( .A1(n13715), .A2(n13719), .ZN(P1_U2956) );
  AOI22_X1 U17201 ( .A1(n20239), .A2(P1_EAX_REG_23__SCAN_IN), .B1(n20238), 
        .B2(P1_UWORD_REG_7__SCAN_IN), .ZN(n13718) );
  NAND2_X1 U17202 ( .A1(n20305), .A2(DATAI_7_), .ZN(n13717) );
  NAND2_X1 U17203 ( .A1(n20303), .A2(BUF1_REG_7__SCAN_IN), .ZN(n13716) );
  NAND2_X1 U17204 ( .A1(n20224), .A2(n20352), .ZN(n14134) );
  NAND2_X1 U17205 ( .A1(n13718), .A2(n14134), .ZN(P1_U2944) );
  AOI22_X1 U17206 ( .A1(n20239), .A2(P1_EAX_REG_20__SCAN_IN), .B1(n20238), 
        .B2(P1_UWORD_REG_4__SCAN_IN), .ZN(n13720) );
  NAND2_X1 U17207 ( .A1(n13720), .A2(n13719), .ZN(P1_U2941) );
  INV_X1 U17208 ( .A(n15667), .ZN(n14287) );
  NAND2_X1 U17209 ( .A1(n13721), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n13821) );
  NOR2_X1 U17210 ( .A1(n13821), .A2(n13822), .ZN(n13820) );
  OAI211_X1 U17211 ( .C1(n13820), .C2(n13722), .A(n15685), .B(n13703), .ZN(
        n13726) );
  NAND2_X1 U17212 ( .A1(n13723), .A2(n13818), .ZN(n13724) );
  AND2_X1 U17213 ( .A1(n13724), .A2(n9950), .ZN(n19136) );
  NAND2_X1 U17214 ( .A1(n14287), .A2(n19136), .ZN(n13725) );
  OAI211_X1 U17215 ( .C1(n14287), .C2(n10583), .A(n13726), .B(n13725), .ZN(
        P2_U2878) );
  NAND2_X1 U17216 ( .A1(n13728), .A2(n13729), .ZN(n13730) );
  NAND2_X1 U17217 ( .A1(n13727), .A2(n13730), .ZN(n14013) );
  NAND2_X1 U17218 ( .A1(n20296), .A2(P1_REIP_REG_2__SCAN_IN), .ZN(n13773) );
  NAND2_X1 U17219 ( .A1(n20242), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13731) );
  OAI211_X1 U17220 ( .C1(n20252), .C2(n13936), .A(n13773), .B(n13731), .ZN(
        n13732) );
  INV_X1 U17221 ( .A(n13732), .ZN(n13737) );
  OR2_X1 U17222 ( .A1(n13734), .A2(n13733), .ZN(n13796) );
  NAND3_X1 U17223 ( .A1(n13796), .A2(n13735), .A3(n20248), .ZN(n13736) );
  OAI211_X1 U17224 ( .C1(n14013), .C2(n20306), .A(n13737), .B(n13736), .ZN(
        P1_U2997) );
  NAND2_X1 U17225 ( .A1(n18813), .A2(n18977), .ZN(n18313) );
  INV_X1 U17226 ( .A(n18313), .ZN(n18334) );
  NAND2_X1 U17227 ( .A1(n18837), .A2(n18821), .ZN(n18333) );
  INV_X1 U17228 ( .A(n18333), .ZN(n18164) );
  OAI22_X1 U17229 ( .A1(n18164), .A2(n13739), .B1(n13738), .B2(n18807), .ZN(
        n13740) );
  NOR2_X1 U17230 ( .A1(n18334), .A2(n13740), .ZN(n18278) );
  OAI21_X1 U17231 ( .B1(n18278), .B2(n18349), .A(n18350), .ZN(n18301) );
  INV_X1 U17232 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n18907) );
  NOR2_X1 U17233 ( .A1(n18316), .A2(n18907), .ZN(n13747) );
  OAI21_X1 U17234 ( .B1(n13743), .B2(n13742), .A(n13741), .ZN(n17982) );
  OAI21_X1 U17235 ( .B1(n13745), .B2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n13744), .ZN(n17984) );
  OAI22_X1 U17236 ( .A1(n18358), .A2(n17982), .B1(n18326), .B2(n17984), .ZN(
        n13746) );
  AOI211_X1 U17237 ( .C1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .C2(n18301), .A(
        n13747), .B(n13746), .ZN(n13752) );
  INV_X1 U17238 ( .A(n13748), .ZN(n16636) );
  INV_X1 U17239 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n13750) );
  OAI22_X1 U17240 ( .A1(n18312), .A2(n18807), .B1(n18337), .B2(n18315), .ZN(
        n18324) );
  NAND2_X1 U17241 ( .A1(n18359), .A2(n18324), .ZN(n18310) );
  INV_X1 U17242 ( .A(n18310), .ZN(n13749) );
  NAND3_X1 U17243 ( .A1(n16636), .A2(n13750), .A3(n13749), .ZN(n13751) );
  NAND2_X1 U17244 ( .A1(n13752), .A2(n13751), .ZN(P3_U2856) );
  NAND2_X1 U17245 ( .A1(n13754), .A2(n13753), .ZN(n13755) );
  NAND2_X1 U17246 ( .A1(n13858), .A2(n13755), .ZN(n13930) );
  OAI222_X1 U17247 ( .A1(n14013), .A2(n9828), .B1(n20182), .B2(n13935), .C1(
        n13930), .C2(n20175), .ZN(P1_U2870) );
  NAND2_X1 U17248 ( .A1(n16201), .A2(n16223), .ZN(n13757) );
  NAND4_X1 U17249 ( .A1(n13758), .A2(n21010), .A3(n13757), .A4(n13756), .ZN(
        n13764) );
  NAND3_X1 U17250 ( .A1(n13462), .A2(n21010), .A3(n13759), .ZN(n13760) );
  NAND3_X1 U17251 ( .A1(n13760), .A2(n11644), .A3(n11643), .ZN(n13761) );
  NAND2_X1 U17252 ( .A1(n13761), .A2(n16193), .ZN(n13763) );
  MUX2_X1 U17253 ( .A(n13764), .B(n13763), .S(n13762), .Z(n13767) );
  NAND3_X1 U17254 ( .A1(n16210), .A2(n15466), .A3(n16201), .ZN(n13765) );
  NAND3_X1 U17255 ( .A1(n13767), .A2(n13766), .A3(n13765), .ZN(n13769) );
  NAND2_X1 U17256 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n13771) );
  OAI21_X1 U17257 ( .B1(n13535), .B2(n20286), .A(n14501), .ZN(n20261) );
  OAI21_X1 U17258 ( .B1(n13771), .B2(n14501), .A(n20261), .ZN(n13789) );
  OAI22_X1 U17259 ( .A1(n12754), .A2(n16201), .B1(n11652), .B2(n10363), .ZN(
        n13772) );
  OAI21_X1 U17260 ( .B1(n20292), .B2(n13930), .A(n13773), .ZN(n13788) );
  OAI22_X1 U17261 ( .A1(n13511), .A2(n13776), .B1(n13775), .B2(n13774), .ZN(
        n13777) );
  NAND3_X1 U17262 ( .A1(n10381), .A2(n13778), .A3(n13777), .ZN(n13779) );
  INV_X1 U17263 ( .A(n20288), .ZN(n13780) );
  NAND2_X1 U17264 ( .A1(n13535), .A2(n20298), .ZN(n20275) );
  NOR2_X1 U17265 ( .A1(n20286), .A2(n20258), .ZN(n13786) );
  NAND2_X1 U17266 ( .A1(n20288), .A2(n13535), .ZN(n13783) );
  INV_X1 U17267 ( .A(n13795), .ZN(n13781) );
  NAND2_X1 U17268 ( .A1(n13781), .A2(n20256), .ZN(n13782) );
  AOI21_X1 U17269 ( .B1(n20286), .B2(n16400), .A(n20277), .ZN(n13784) );
  INV_X1 U17270 ( .A(n13784), .ZN(n13785) );
  MUX2_X1 U17271 ( .A(n13786), .B(n13785), .S(
        P1_INSTADDRPOINTER_REG_2__SCAN_IN), .Z(n13787) );
  AOI211_X1 U17272 ( .C1(n20289), .C2(n13789), .A(n13788), .B(n13787), .ZN(
        n13798) );
  NAND2_X1 U17273 ( .A1(n13791), .A2(n13790), .ZN(n16199) );
  AND2_X1 U17274 ( .A1(n13792), .A2(n16199), .ZN(n16189) );
  OAI211_X1 U17275 ( .C1(n11679), .C2(n10363), .A(n13793), .B(n16189), .ZN(
        n13794) );
  NAND3_X1 U17276 ( .A1(n13796), .A2(n13735), .A3(n20278), .ZN(n13797) );
  NAND2_X1 U17277 ( .A1(n13798), .A2(n13797), .ZN(P1_U3029) );
  INV_X1 U17278 ( .A(n20239), .ZN(n13810) );
  INV_X1 U17279 ( .A(n15111), .ZN(n13799) );
  NAND2_X1 U17280 ( .A1(n20224), .A2(n13799), .ZN(n20240) );
  NAND2_X1 U17281 ( .A1(n20238), .A2(P1_UWORD_REG_14__SCAN_IN), .ZN(n13800) );
  OAI211_X1 U17282 ( .C1(n13810), .C2(n13022), .A(n20240), .B(n13800), .ZN(
        P1_U2951) );
  INV_X1 U17283 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n21270) );
  NAND2_X1 U17284 ( .A1(n20238), .A2(P1_UWORD_REG_0__SCAN_IN), .ZN(n13803) );
  INV_X1 U17285 ( .A(DATAI_0_), .ZN(n13802) );
  NAND2_X1 U17286 ( .A1(n20303), .A2(BUF1_REG_0__SCAN_IN), .ZN(n13801) );
  OAI21_X1 U17287 ( .B1(n20303), .B2(n13802), .A(n13801), .ZN(n20316) );
  NAND2_X1 U17288 ( .A1(n20224), .A2(n20316), .ZN(n14148) );
  OAI211_X1 U17289 ( .C1(n13810), .C2(n21270), .A(n13803), .B(n14148), .ZN(
        P1_U2937) );
  INV_X1 U17290 ( .A(DATAI_11_), .ZN(n21174) );
  MUX2_X1 U17291 ( .A(n21174), .B(n16673), .S(n20303), .Z(n15117) );
  INV_X1 U17292 ( .A(n15117), .ZN(n13804) );
  NAND2_X1 U17293 ( .A1(n20224), .A2(n13804), .ZN(n20232) );
  NAND2_X1 U17294 ( .A1(n20238), .A2(P1_UWORD_REG_11__SCAN_IN), .ZN(n13805) );
  OAI211_X1 U17295 ( .C1(n13810), .C2(n21309), .A(n20232), .B(n13805), .ZN(
        P1_U2948) );
  INV_X1 U17296 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n15107) );
  INV_X1 U17297 ( .A(DATAI_15_), .ZN(n13807) );
  INV_X1 U17298 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n13806) );
  MUX2_X1 U17299 ( .A(n13807), .B(n13806), .S(n20303), .Z(n15108) );
  INV_X1 U17300 ( .A(P1_LWORD_REG_15__SCAN_IN), .ZN(n20184) );
  OAI222_X1 U17301 ( .A1(n13810), .A2(n15107), .B1(n13809), .B2(n15108), .C1(
        n20184), .C2(n13808), .ZN(P1_U2967) );
  AOI21_X1 U17302 ( .B1(n13812), .B2(n13709), .A(n13811), .ZN(n19127) );
  NOR2_X1 U17303 ( .A1(n14287), .A2(n19122), .ZN(n13816) );
  AOI211_X1 U17304 ( .C1(n13814), .C2(n13813), .A(n15694), .B(n13829), .ZN(
        n13815) );
  AOI211_X1 U17305 ( .C1(n19127), .C2(n14287), .A(n13816), .B(n13815), .ZN(
        n13817) );
  INV_X1 U17306 ( .A(n13817), .ZN(P2_U2876) );
  OAI21_X1 U17307 ( .B1(n13819), .B2(n13662), .A(n13818), .ZN(n14159) );
  NOR2_X1 U17308 ( .A1(n15661), .A2(n14159), .ZN(n13824) );
  AOI211_X1 U17309 ( .C1(n13822), .C2(n13821), .A(n15694), .B(n13820), .ZN(
        n13823) );
  AOI211_X1 U17310 ( .C1(P2_EBX_REG_8__SCAN_IN), .C2(n15661), .A(n13824), .B(
        n13823), .ZN(n13825) );
  INV_X1 U17311 ( .A(n13825), .ZN(P2_U2879) );
  OR2_X1 U17312 ( .A1(n13811), .A2(n13827), .ZN(n13828) );
  AND2_X1 U17313 ( .A1(n13826), .A2(n13828), .ZN(n16565) );
  INV_X1 U17314 ( .A(n16565), .ZN(n13834) );
  INV_X1 U17315 ( .A(n14030), .ZN(n13830) );
  OAI211_X1 U17316 ( .C1(n13829), .C2(n13831), .A(n13830), .B(n15685), .ZN(
        n13833) );
  NAND2_X1 U17317 ( .A1(n15667), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n13832) );
  OAI211_X1 U17318 ( .C1(n13834), .C2(n15661), .A(n13833), .B(n13832), .ZN(
        P2_U2875) );
  OAI21_X1 U17319 ( .B1(n16196), .B2(n13840), .A(n14988), .ZN(n20161) );
  INV_X1 U17320 ( .A(n20161), .ZN(n13940) );
  INV_X1 U17321 ( .A(n13835), .ZN(n13836) );
  NOR2_X1 U17322 ( .A1(n13840), .A2(n13839), .ZN(n20152) );
  INV_X1 U17323 ( .A(n20152), .ZN(n13884) );
  OAI22_X1 U17324 ( .A1(n20158), .A2(n13846), .B1(n13576), .B2(n20117), .ZN(
        n13843) );
  OAI22_X1 U17325 ( .A1(n13841), .A2(n20124), .B1(n20151), .B2(
        P1_REIP_REG_1__SCAN_IN), .ZN(n13842) );
  AOI211_X1 U17326 ( .C1(n20147), .C2(P1_EBX_REG_1__SCAN_IN), .A(n13843), .B(
        n13842), .ZN(n13844) );
  OAI21_X1 U17327 ( .B1(n13838), .B2(n13884), .A(n13844), .ZN(n13845) );
  AOI21_X1 U17328 ( .B1(n20154), .B2(n13846), .A(n13845), .ZN(n13847) );
  OAI21_X1 U17329 ( .B1(n13940), .B2(n14010), .A(n13847), .ZN(P1_U2839) );
  OAI21_X1 U17330 ( .B1(n13850), .B2(n13849), .A(n13848), .ZN(n20268) );
  OR2_X1 U17331 ( .A1(n13853), .A2(n13852), .ZN(n13854) );
  AND2_X1 U17332 ( .A1(n13851), .A2(n13854), .ZN(n13887) );
  AOI22_X1 U17333 ( .A1(n20242), .A2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B1(
        n20296), .B2(P1_REIP_REG_3__SCAN_IN), .ZN(n13855) );
  OAI21_X1 U17334 ( .B1(n13890), .B2(n20252), .A(n13855), .ZN(n13856) );
  AOI21_X1 U17335 ( .B1(n13887), .B2(n16325), .A(n13856), .ZN(n13857) );
  OAI21_X1 U17336 ( .B1(n20268), .B2(n20088), .A(n13857), .ZN(P1_U2996) );
  INV_X1 U17337 ( .A(n13887), .ZN(n14006) );
  INV_X1 U17338 ( .A(P1_EBX_REG_3__SCAN_IN), .ZN(n13883) );
  XOR2_X1 U17339 ( .A(n13859), .B(n13858), .Z(n20270) );
  INV_X1 U17340 ( .A(n20270), .ZN(n13860) );
  OAI222_X1 U17341 ( .A1(n14006), .A2(n9828), .B1(n20182), .B2(n13883), .C1(
        n13860), .C2(n20175), .ZN(P1_U2869) );
  AOI22_X1 U17342 ( .A1(n20149), .A2(n13861), .B1(n20147), .B2(
        P1_EBX_REG_0__SCAN_IN), .ZN(n13862) );
  OAI21_X1 U17343 ( .B1(n14958), .B2(n13863), .A(n13862), .ZN(n13864) );
  AOI21_X1 U17344 ( .B1(n20422), .B2(n20152), .A(n13864), .ZN(n13866) );
  OAI21_X1 U17345 ( .B1(n20154), .B2(n20140), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13865) );
  OAI211_X1 U17346 ( .C1(n13940), .C2(n14015), .A(n13866), .B(n13865), .ZN(
        P1_U2840) );
  XNOR2_X1 U17347 ( .A(n13868), .B(n13867), .ZN(n13869) );
  XNOR2_X1 U17348 ( .A(n13870), .B(n13869), .ZN(n13897) );
  XOR2_X1 U17349 ( .A(n9900), .B(n13871), .Z(n13895) );
  OAI21_X1 U17350 ( .B1(n13874), .B2(n13873), .A(n13872), .ZN(n20014) );
  INV_X1 U17351 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n19938) );
  OAI22_X1 U17352 ( .A1(n19327), .A2(n20014), .B1(n19938), .B2(n19345), .ZN(
        n13876) );
  NOR2_X1 U17353 ( .A1(n14054), .A2(n13867), .ZN(n13875) );
  AOI211_X1 U17354 ( .C1(n19341), .C2(n14070), .A(n13876), .B(n13875), .ZN(
        n13877) );
  OAI21_X1 U17355 ( .B1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n14053), .A(
        n13877), .ZN(n13878) );
  AOI21_X1 U17356 ( .B1(n13895), .B2(n16577), .A(n13878), .ZN(n13879) );
  OAI21_X1 U17357 ( .B1(n19363), .B2(n13897), .A(n13879), .ZN(P2_U3043) );
  INV_X1 U17358 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n20932) );
  NAND4_X1 U17359 ( .A1(n20137), .A2(n20932), .A3(P1_REIP_REG_2__SCAN_IN), 
        .A4(P1_REIP_REG_1__SCAN_IN), .ZN(n13882) );
  OAI221_X1 U17360 ( .B1(n20151), .B2(P1_REIP_REG_1__SCAN_IN), .C1(n20151), 
        .C2(P1_REIP_REG_2__SCAN_IN), .A(n20117), .ZN(n13880) );
  AOI22_X1 U17361 ( .A1(n20140), .A2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B1(
        P1_REIP_REG_3__SCAN_IN), .B2(n13880), .ZN(n13881) );
  OAI211_X1 U17362 ( .C1(n13883), .C2(n20122), .A(n13882), .B(n13881), .ZN(
        n13886) );
  INV_X1 U17363 ( .A(n20597), .ZN(n13978) );
  NOR2_X1 U17364 ( .A1(n13978), .A2(n13884), .ZN(n13885) );
  AOI211_X1 U17365 ( .C1(n20270), .C2(n20149), .A(n13886), .B(n13885), .ZN(
        n13889) );
  NAND2_X1 U17366 ( .A1(n20161), .A2(n13887), .ZN(n13888) );
  OAI211_X1 U17367 ( .C1(n20143), .C2(n13890), .A(n13889), .B(n13888), .ZN(
        P1_U2837) );
  AOI22_X1 U17368 ( .A1(n19313), .A2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .B1(
        P2_REIP_REG_3__SCAN_IN), .B2(n19170), .ZN(n13892) );
  NAND2_X1 U17369 ( .A1(n16550), .A2(n14062), .ZN(n13891) );
  OAI211_X1 U17370 ( .C1(n13893), .C2(n16545), .A(n13892), .B(n13891), .ZN(
        n13894) );
  AOI21_X1 U17371 ( .B1(n13895), .B2(n16539), .A(n13894), .ZN(n13896) );
  OAI21_X1 U17372 ( .B1(n16553), .B2(n13897), .A(n13896), .ZN(P2_U3011) );
  INV_X1 U17373 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n13899) );
  AOI22_X1 U17374 ( .A1(P1_UWORD_REG_4__SCAN_IN), .A2(n13910), .B1(n20204), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n13898) );
  OAI21_X1 U17375 ( .B1(n13899), .B2(n13912), .A(n13898), .ZN(P1_U2916) );
  INV_X1 U17376 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n13901) );
  AOI22_X1 U17377 ( .A1(P1_UWORD_REG_6__SCAN_IN), .A2(n13910), .B1(n20204), 
        .B2(P1_DATAO_REG_22__SCAN_IN), .ZN(n13900) );
  OAI21_X1 U17378 ( .B1(n13901), .B2(n13912), .A(n13900), .ZN(P1_U2914) );
  AOI22_X1 U17379 ( .A1(P1_UWORD_REG_7__SCAN_IN), .A2(n13910), .B1(n20204), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n13902) );
  OAI21_X1 U17380 ( .B1(n15070), .B2(n13912), .A(n13902), .ZN(P1_U2913) );
  INV_X1 U17381 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n13904) );
  AOI22_X1 U17382 ( .A1(P1_UWORD_REG_2__SCAN_IN), .A2(n13910), .B1(n20204), 
        .B2(P1_DATAO_REG_18__SCAN_IN), .ZN(n13903) );
  OAI21_X1 U17383 ( .B1(n13904), .B2(n13912), .A(n13903), .ZN(P1_U2918) );
  INV_X1 U17384 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n13906) );
  AOI22_X1 U17385 ( .A1(P1_UWORD_REG_1__SCAN_IN), .A2(n13910), .B1(n20204), 
        .B2(P1_DATAO_REG_17__SCAN_IN), .ZN(n13905) );
  OAI21_X1 U17386 ( .B1(n13906), .B2(n13912), .A(n13905), .ZN(P1_U2919) );
  AOI22_X1 U17387 ( .A1(P1_UWORD_REG_0__SCAN_IN), .A2(n13910), .B1(n20204), 
        .B2(P1_DATAO_REG_16__SCAN_IN), .ZN(n13907) );
  OAI21_X1 U17388 ( .B1(n21270), .B2(n13912), .A(n13907), .ZN(P1_U2920) );
  INV_X1 U17389 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n13909) );
  AOI22_X1 U17390 ( .A1(P1_UWORD_REG_3__SCAN_IN), .A2(n13910), .B1(n20204), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n13908) );
  OAI21_X1 U17391 ( .B1(n13909), .B2(n13912), .A(n13908), .ZN(P1_U2917) );
  INV_X1 U17392 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n15080) );
  AOI22_X1 U17393 ( .A1(P1_UWORD_REG_5__SCAN_IN), .A2(n13910), .B1(n20204), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n13911) );
  OAI21_X1 U17394 ( .B1(n15080), .B2(n13912), .A(n13911), .ZN(P1_U2915) );
  INV_X1 U17395 ( .A(n19266), .ZN(n19255) );
  NAND2_X1 U17396 ( .A1(n13914), .A2(n13913), .ZN(n13917) );
  INV_X1 U17397 ( .A(n13915), .ZN(n13916) );
  NAND2_X1 U17398 ( .A1(n13917), .A2(n13916), .ZN(n20021) );
  NOR2_X1 U17399 ( .A1(n19364), .A2(n20021), .ZN(n13920) );
  AOI21_X1 U17400 ( .B1(n19364), .B2(n20021), .A(n13920), .ZN(n19269) );
  OAI22_X1 U17401 ( .A1(n13919), .A2(n13918), .B1(n20029), .B2(n20031), .ZN(
        n19268) );
  NAND2_X1 U17402 ( .A1(n19269), .A2(n19268), .ZN(n19267) );
  INV_X1 U17403 ( .A(n13920), .ZN(n13921) );
  NAND2_X1 U17404 ( .A1(n19267), .A2(n13921), .ZN(n13923) );
  XOR2_X1 U17405 ( .A(n20014), .B(n19431), .Z(n13922) );
  NAND2_X1 U17406 ( .A1(n13923), .A2(n13922), .ZN(n14039) );
  OAI21_X1 U17407 ( .B1(n13923), .B2(n13922), .A(n14039), .ZN(n13924) );
  NAND2_X1 U17408 ( .A1(n13924), .A2(n19270), .ZN(n13927) );
  INV_X1 U17409 ( .A(n20014), .ZN(n13925) );
  AOI22_X1 U17410 ( .A1(n19265), .A2(n13925), .B1(P2_EAX_REG_3__SCAN_IN), .B2(
        n19257), .ZN(n13926) );
  OAI211_X1 U17411 ( .C1(n19255), .C2(n14382), .A(n13927), .B(n13926), .ZN(
        P2_U2916) );
  INV_X1 U17412 ( .A(n13553), .ZN(n20313) );
  INV_X1 U17413 ( .A(P1_REIP_REG_2__SCAN_IN), .ZN(n13929) );
  NAND2_X1 U17414 ( .A1(n13576), .A2(n13929), .ZN(n13928) );
  OAI211_X1 U17415 ( .C1(n13576), .C2(n13929), .A(n20137), .B(n13928), .ZN(
        n13934) );
  INV_X1 U17416 ( .A(n20117), .ZN(n20135) );
  INV_X1 U17417 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n13931) );
  OAI22_X1 U17418 ( .A1(n13931), .A2(n20158), .B1(n20124), .B2(n13930), .ZN(
        n13932) );
  AOI21_X1 U17419 ( .B1(n20135), .B2(P1_REIP_REG_2__SCAN_IN), .A(n13932), .ZN(
        n13933) );
  OAI211_X1 U17420 ( .C1(n20122), .C2(n13935), .A(n13934), .B(n13933), .ZN(
        n13938) );
  NOR2_X1 U17421 ( .A1(n20143), .A2(n13936), .ZN(n13937) );
  AOI211_X1 U17422 ( .C1(n20152), .C2(n20313), .A(n13938), .B(n13937), .ZN(
        n13939) );
  OAI21_X1 U17423 ( .B1(n13940), .B2(n14013), .A(n13939), .ZN(P1_U2838) );
  NOR2_X1 U17424 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(n16442), .ZN(n13955) );
  MUX2_X1 U17425 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n13941), .S(
        n16172), .Z(n16181) );
  AOI22_X1 U17426 ( .A1(n13955), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n16442), .B2(n16181), .ZN(n13957) );
  INV_X1 U17427 ( .A(n13944), .ZN(n15470) );
  AOI21_X1 U17428 ( .B1(n15472), .B2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13942) );
  NOR2_X1 U17429 ( .A1(n11716), .A2(n13942), .ZN(n15479) );
  NAND3_X1 U17430 ( .A1(n13944), .A2(n13943), .A3(n15479), .ZN(n13952) );
  XNOR2_X1 U17431 ( .A(n13945), .B(n11535), .ZN(n13950) );
  NOR2_X1 U17432 ( .A1(n13947), .A2(n13946), .ZN(n13948) );
  AOI22_X1 U17433 ( .A1(n16175), .A2(n13950), .B1(n13949), .B2(n13948), .ZN(
        n13951) );
  NAND2_X1 U17434 ( .A1(n13952), .A2(n13951), .ZN(n13953) );
  AOI21_X1 U17435 ( .B1(n20597), .B2(n15470), .A(n13953), .ZN(n15483) );
  NOR2_X1 U17436 ( .A1(n16172), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13954) );
  AOI21_X1 U17437 ( .B1(n15483), .B2(n16172), .A(n13954), .ZN(n16182) );
  AOI22_X1 U17438 ( .A1(n13955), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n16182), .B2(n16442), .ZN(n13956) );
  NOR2_X1 U17439 ( .A1(n13957), .A2(n13956), .ZN(n16185) );
  INV_X1 U17440 ( .A(n16185), .ZN(n13959) );
  NOR2_X1 U17441 ( .A1(n13959), .A2(n13958), .ZN(n13966) );
  AND2_X1 U17442 ( .A1(n16172), .A2(n16442), .ZN(n13961) );
  OAI22_X1 U17443 ( .A1(n13961), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B1(
        n16442), .B2(n20089), .ZN(n13960) );
  AOI21_X1 U17444 ( .B1(n13962), .B2(n13961), .A(n13960), .ZN(n16186) );
  NOR3_X1 U17445 ( .A1(n13966), .A2(n16186), .A3(P1_FLUSH_REG_SCAN_IN), .ZN(
        n13965) );
  NOR2_X1 U17446 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13964) );
  OR3_X1 U17447 ( .A1(n13966), .A2(n16186), .A3(n16438), .ZN(n16213) );
  INV_X1 U17448 ( .A(n16213), .ZN(n13969) );
  AND2_X1 U17449 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n20738), .ZN(n15462) );
  OAI22_X1 U17450 ( .A1(n11991), .A2(n20848), .B1(n13967), .B2(n15462), .ZN(
        n13968) );
  OAI21_X1 U17451 ( .B1(n13969), .B2(n13968), .A(n20301), .ZN(n13970) );
  OAI21_X1 U17452 ( .B1(n20301), .B2(n20767), .A(n13970), .ZN(P1_U3478) );
  NAND2_X1 U17453 ( .A1(n9853), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n20700) );
  OR2_X1 U17454 ( .A1(n20700), .A2(n20848), .ZN(n20854) );
  NOR2_X1 U17455 ( .A1(n20496), .A2(n20854), .ZN(n20567) );
  NOR3_X1 U17456 ( .A1(n20855), .A2(n20848), .A3(n20628), .ZN(n20773) );
  INV_X1 U17457 ( .A(n20773), .ZN(n13977) );
  INV_X1 U17458 ( .A(n20594), .ZN(n13975) );
  OAI211_X1 U17459 ( .C1(n20593), .C2(n21000), .A(n13975), .B(n20769), .ZN(
        n13976) );
  OAI211_X1 U17460 ( .C1(n13978), .C2(n15462), .A(n13977), .B(n13976), .ZN(
        n13979) );
  OAI21_X1 U17461 ( .B1(n20567), .B2(n13979), .A(n20301), .ZN(n13980) );
  OAI21_X1 U17462 ( .B1(n20387), .B2(n20301), .A(n13980), .ZN(P1_U3475) );
  NOR2_X1 U17463 ( .A1(n17426), .A2(n13981), .ZN(n17286) );
  AOI22_X1 U17464 ( .A1(n9829), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17343), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n13992) );
  AOI22_X1 U17465 ( .A1(n12552), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17357), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n13991) );
  OAI22_X1 U17466 ( .A1(n17395), .A2(n17389), .B1(n17340), .B2(n13982), .ZN(
        n13989) );
  AOI22_X1 U17467 ( .A1(n13089), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17361), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n13987) );
  AOI22_X1 U17468 ( .A1(n17379), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n13120), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n13984) );
  AOI22_X1 U17469 ( .A1(n17309), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n17245), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n13983) );
  OAI211_X1 U17470 ( .C1(n17363), .C2(n17381), .A(n13984), .B(n13983), .ZN(
        n13985) );
  AOI21_X1 U17471 ( .B1(n17327), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A(
        n13985), .ZN(n13986) );
  OAI211_X1 U17472 ( .C1(n12551), .C2(n17383), .A(n13987), .B(n13986), .ZN(
        n13988) );
  AOI211_X1 U17473 ( .C1(n17365), .C2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A(
        n13989), .B(n13988), .ZN(n13990) );
  NAND3_X1 U17474 ( .A1(n13992), .A2(n13991), .A3(n13990), .ZN(n17507) );
  AOI22_X1 U17475 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n17286), .B1(n17426), 
        .B2(n17507), .ZN(n13996) );
  INV_X1 U17476 ( .A(P3_EBX_REG_16__SCAN_IN), .ZN(n13994) );
  NAND3_X1 U17477 ( .A1(n17547), .A2(P3_EBX_REG_12__SCAN_IN), .A3(n9920), .ZN(
        n16137) );
  NAND2_X1 U17478 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n17301), .ZN(n17300) );
  INV_X1 U17479 ( .A(n17300), .ZN(n13993) );
  NAND3_X1 U17480 ( .A1(P3_EBX_REG_15__SCAN_IN), .A2(n13994), .A3(n13993), 
        .ZN(n13995) );
  NAND2_X1 U17481 ( .A1(n13996), .A2(n13995), .ZN(P3_U2687) );
  XNOR2_X1 U17482 ( .A(n14030), .B(n14032), .ZN(n14001) );
  NAND2_X1 U17483 ( .A1(n13826), .A2(n13997), .ZN(n13998) );
  NAND2_X1 U17484 ( .A1(n14027), .A2(n13998), .ZN(n19115) );
  INV_X1 U17485 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n13999) );
  MUX2_X1 U17486 ( .A(n19115), .B(n13999), .S(n15667), .Z(n14000) );
  OAI21_X1 U17487 ( .B1(n14001), .B2(n15694), .A(n14000), .ZN(P2_U2874) );
  INV_X1 U17488 ( .A(DATAI_3_), .ZN(n14004) );
  NAND2_X1 U17489 ( .A1(n20303), .A2(BUF1_REG_3__SCAN_IN), .ZN(n14003) );
  OAI21_X1 U17490 ( .B1(n20303), .B2(n14004), .A(n14003), .ZN(n20332) );
  INV_X1 U17491 ( .A(n20332), .ZN(n14005) );
  INV_X1 U17492 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n20201) );
  OAI222_X1 U17493 ( .A1(n14006), .A2(n15118), .B1(n15116), .B2(n14005), .C1(
        n15090), .C2(n20201), .ZN(P1_U2901) );
  INV_X1 U17494 ( .A(DATAI_1_), .ZN(n14008) );
  NAND2_X1 U17495 ( .A1(n20303), .A2(BUF1_REG_1__SCAN_IN), .ZN(n14007) );
  OAI21_X1 U17496 ( .B1(n20303), .B2(n14008), .A(n14007), .ZN(n20325) );
  INV_X1 U17497 ( .A(n20325), .ZN(n14009) );
  INV_X1 U17498 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n20206) );
  OAI222_X1 U17499 ( .A1(n14010), .A2(n15118), .B1(n14009), .B2(n15116), .C1(
        n15090), .C2(n20206), .ZN(P1_U2903) );
  NAND2_X1 U17500 ( .A1(n20305), .A2(DATAI_2_), .ZN(n14012) );
  NAND2_X1 U17501 ( .A1(n20303), .A2(BUF1_REG_2__SCAN_IN), .ZN(n14011) );
  INV_X1 U17502 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n20203) );
  OAI222_X1 U17503 ( .A1(n14013), .A2(n15118), .B1(n20328), .B2(n15116), .C1(
        n15090), .C2(n20203), .ZN(P1_U2902) );
  INV_X1 U17504 ( .A(n20316), .ZN(n14014) );
  INV_X1 U17505 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n20209) );
  OAI222_X1 U17506 ( .A1(n14015), .A2(n15118), .B1(n14014), .B2(n15116), .C1(
        n15090), .C2(n20209), .ZN(P1_U2904) );
  INV_X1 U17507 ( .A(n14016), .ZN(n14017) );
  XNOR2_X1 U17508 ( .A(n13851), .B(n14017), .ZN(n20247) );
  INV_X1 U17509 ( .A(n20247), .ZN(n14047) );
  INV_X1 U17510 ( .A(n15116), .ZN(n14018) );
  AOI22_X1 U17511 ( .A1(n14018), .A2(n20335), .B1(P1_EAX_REG_4__SCAN_IN), .B2(
        n16293), .ZN(n14019) );
  OAI21_X1 U17512 ( .B1(n14047), .B2(n15118), .A(n14019), .ZN(P1_U2900) );
  OR2_X1 U17513 ( .A1(n14022), .A2(n14021), .ZN(n14023) );
  AND2_X1 U17514 ( .A1(n14020), .A2(n14023), .ZN(n20179) );
  INV_X1 U17515 ( .A(n20179), .ZN(n14025) );
  INV_X1 U17516 ( .A(DATAI_5_), .ZN(n14024) );
  INV_X1 U17517 ( .A(BUF1_REG_5__SCAN_IN), .ZN(n16681) );
  MUX2_X1 U17518 ( .A(n14024), .B(n16681), .S(n20303), .Z(n15081) );
  INV_X1 U17519 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n20197) );
  OAI222_X1 U17520 ( .A1(n14025), .A2(n15118), .B1(n15081), .B2(n15116), .C1(
        n15090), .C2(n20197), .ZN(P1_U2899) );
  AOI21_X1 U17521 ( .B1(n14028), .B2(n14027), .A(n14026), .ZN(n19102) );
  INV_X1 U17522 ( .A(n19102), .ZN(n14036) );
  AND2_X1 U17523 ( .A1(n14031), .A2(n14032), .ZN(n14029) );
  NAND2_X1 U17524 ( .A1(n14030), .A2(n14029), .ZN(n14205) );
  AOI21_X1 U17525 ( .B1(n14030), .B2(n14032), .A(n14031), .ZN(n14033) );
  OR3_X1 U17526 ( .A1(n14281), .A2(n14033), .A3(n15694), .ZN(n14035) );
  NAND2_X1 U17527 ( .A1(n15661), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n14034) );
  OAI211_X1 U17528 ( .C1(n14036), .C2(n15661), .A(n14035), .B(n14034), .ZN(
        P2_U2873) );
  NAND2_X1 U17529 ( .A1(n19431), .A2(n20014), .ZN(n14038) );
  XNOR2_X1 U17530 ( .A(n13872), .B(n14037), .ZN(n14185) );
  INV_X1 U17531 ( .A(n14185), .ZN(n14040) );
  AOI21_X1 U17532 ( .B1(n14039), .B2(n14038), .A(n14040), .ZN(n19260) );
  XNOR2_X1 U17533 ( .A(n19260), .B(n19259), .ZN(n14043) );
  AOI22_X1 U17534 ( .A1(n19265), .A2(n14040), .B1(P2_EAX_REG_4__SCAN_IN), .B2(
        n19257), .ZN(n14042) );
  NAND2_X1 U17535 ( .A1(n19266), .A2(n19396), .ZN(n14041) );
  OAI211_X1 U17536 ( .C1(n14043), .C2(n19258), .A(n14042), .B(n14041), .ZN(
        P2_U2915) );
  OR2_X1 U17537 ( .A1(n14045), .A2(n14044), .ZN(n14046) );
  INV_X1 U17538 ( .A(P1_EBX_REG_4__SCAN_IN), .ZN(n14048) );
  OAI222_X1 U17539 ( .A1(n20257), .A2(n20175), .B1(n14048), .B2(n20182), .C1(
        n9828), .C2(n14047), .ZN(P1_U2868) );
  NAND2_X1 U17540 ( .A1(n14050), .A2(n14049), .ZN(n14051) );
  XNOR2_X1 U17541 ( .A(n14051), .B(n14269), .ZN(n19320) );
  XNOR2_X1 U17542 ( .A(n14052), .B(n9961), .ZN(n19314) );
  NOR2_X1 U17543 ( .A1(n13867), .A2(n14053), .ZN(n14268) );
  OAI21_X1 U17544 ( .B1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n19353), .A(
        n14054), .ZN(n14274) );
  INV_X1 U17545 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n21299) );
  NOR2_X1 U17546 ( .A1(n21299), .A2(n19345), .ZN(n14055) );
  AOI221_X1 U17547 ( .B1(n14268), .B2(n14269), .C1(n14274), .C2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A(n14055), .ZN(n14057) );
  NAND2_X1 U17548 ( .A1(n19316), .A2(n19341), .ZN(n14056) );
  OAI211_X1 U17549 ( .C1(n14185), .C2(n19327), .A(n14057), .B(n14056), .ZN(
        n14058) );
  AOI21_X1 U17550 ( .B1(n19331), .B2(n19314), .A(n14058), .ZN(n14059) );
  OAI21_X1 U17551 ( .B1(n19356), .B2(n19320), .A(n14059), .ZN(P2_U3042) );
  NAND2_X1 U17552 ( .A1(n10135), .A2(n14060), .ZN(n14061) );
  XNOR2_X1 U17553 ( .A(n14062), .B(n14061), .ZN(n14063) );
  NAND2_X1 U17554 ( .A1(n14063), .A2(n19175), .ZN(n14072) );
  OAI22_X1 U17555 ( .A1(n14064), .A2(n19180), .B1(n19938), .B2(n19181), .ZN(
        n14066) );
  NOR2_X1 U17556 ( .A1(n19200), .A2(n20014), .ZN(n14065) );
  AOI211_X1 U17557 ( .C1(P2_EBX_REG_3__SCAN_IN), .C2(n19205), .A(n14066), .B(
        n14065), .ZN(n14067) );
  OAI21_X1 U17558 ( .B1(n14068), .B2(n19202), .A(n14067), .ZN(n14069) );
  AOI21_X1 U17559 ( .B1(n19179), .B2(n14070), .A(n14069), .ZN(n14071) );
  OAI211_X1 U17560 ( .C1(n19431), .C2(n19208), .A(n14072), .B(n14071), .ZN(
        P2_U2852) );
  INV_X1 U17561 ( .A(n14073), .ZN(n14127) );
  INV_X1 U17562 ( .A(n14074), .ZN(n14092) );
  NAND2_X1 U17563 ( .A1(n9842), .A2(n14075), .ZN(n14080) );
  NAND2_X1 U17564 ( .A1(n14076), .A2(n14080), .ZN(n14079) );
  NAND2_X1 U17565 ( .A1(n14090), .A2(n14077), .ZN(n14078) );
  OAI211_X1 U17566 ( .C1(n14081), .C2(n14080), .A(n14079), .B(n14078), .ZN(
        n14082) );
  AOI21_X1 U17567 ( .B1(n19342), .B2(n14092), .A(n14082), .ZN(n16120) );
  NAND2_X1 U17568 ( .A1(n9860), .A2(n14092), .ZN(n14087) );
  INV_X1 U17569 ( .A(n11469), .ZN(n14084) );
  NAND2_X1 U17570 ( .A1(n14084), .A2(n14083), .ZN(n14089) );
  NOR2_X1 U17571 ( .A1(n10425), .A2(n10435), .ZN(n14085) );
  AOI22_X1 U17572 ( .A1(n14090), .A2(n10438), .B1(n14089), .B2(n14085), .ZN(
        n14086) );
  NAND2_X1 U17573 ( .A1(n14087), .A2(n14086), .ZN(n16116) );
  NAND2_X1 U17574 ( .A1(n16116), .A2(n20033), .ZN(n14094) );
  MUX2_X1 U17575 ( .A(n14090), .B(n14089), .S(n14088), .Z(n14091) );
  AOI21_X1 U17576 ( .B1(n14093), .B2(n14092), .A(n14091), .ZN(n16106) );
  NAND3_X1 U17577 ( .A1(n14094), .A2(n16106), .A3(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n14095) );
  OAI211_X1 U17578 ( .C1(n20033), .C2(n16116), .A(n14095), .B(n14098), .ZN(
        n14096) );
  AOI21_X1 U17579 ( .B1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n16120), .A(
        n14096), .ZN(n14101) );
  MUX2_X1 U17580 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n14097), .S(
        n14098), .Z(n14103) );
  MUX2_X1 U17581 ( .A(n9840), .B(n16120), .S(n14098), .Z(n14122) );
  NOR2_X1 U17582 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n14122), .ZN(
        n14099) );
  OR3_X1 U17583 ( .A1(n14101), .A2(n14103), .A3(n14099), .ZN(n14100) );
  AOI22_X1 U17584 ( .A1(n14101), .A2(n14103), .B1(n20017), .B2(n14100), .ZN(
        n14102) );
  NOR2_X1 U17585 ( .A1(n14102), .A2(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(
        n14125) );
  INV_X1 U17586 ( .A(n14103), .ZN(n14123) );
  OR2_X1 U17587 ( .A1(n14108), .A2(n14105), .ZN(n14110) );
  INV_X1 U17588 ( .A(n14106), .ZN(n14107) );
  NAND2_X1 U17589 ( .A1(n14108), .A2(n14107), .ZN(n14109) );
  OAI211_X1 U17590 ( .C1(n10963), .C2(n14111), .A(n14110), .B(n14109), .ZN(
        n20046) );
  INV_X1 U17591 ( .A(n14112), .ZN(n14118) );
  NOR4_X1 U17592 ( .A1(n14115), .A2(n10963), .A3(n14114), .A4(n14113), .ZN(
        n19041) );
  OAI21_X1 U17593 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(P2_MORE_REG_SCAN_IN), .A(
        n19041), .ZN(n14117) );
  NAND3_X1 U17594 ( .A1(n16157), .A2(n16156), .A3(n16155), .ZN(n14116) );
  OAI211_X1 U17595 ( .C1(n20064), .C2(n14118), .A(n14117), .B(n14116), .ZN(
        n14119) );
  AOI211_X1 U17596 ( .C1(n14120), .C2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(
        n20046), .B(n14119), .ZN(n14121) );
  OAI21_X1 U17597 ( .B1(n14123), .B2(n14122), .A(n14121), .ZN(n14124) );
  NOR2_X1 U17598 ( .A1(n14125), .A2(n14124), .ZN(n16593) );
  AOI21_X1 U17599 ( .B1(n16593), .B2(n13362), .A(n14298), .ZN(n14126) );
  AOI21_X1 U17600 ( .B1(n14128), .B2(n14127), .A(n14126), .ZN(n14133) );
  NOR2_X1 U17601 ( .A1(n14129), .A2(n20034), .ZN(n20059) );
  NAND2_X1 U17602 ( .A1(n14133), .A2(n20059), .ZN(n16594) );
  NAND4_X1 U17603 ( .A1(n16594), .A2(n20069), .A3(P2_STATE2_REG_0__SCAN_IN), 
        .A4(n20005), .ZN(n14132) );
  NAND2_X1 U17604 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n20034), .ZN(n19037) );
  AOI211_X1 U17605 ( .C1(n16594), .C2(n19037), .A(n20069), .B(n13362), .ZN(
        n14130) );
  NOR2_X1 U17606 ( .A1(n19175), .A2(n14130), .ZN(n14131) );
  OAI211_X1 U17607 ( .C1(n14133), .C2(n19040), .A(n14132), .B(n14131), .ZN(
        P2_U3177) );
  AOI22_X1 U17608 ( .A1(n20239), .A2(P1_EAX_REG_7__SCAN_IN), .B1(n20238), .B2(
        P1_LWORD_REG_7__SCAN_IN), .ZN(n14135) );
  NAND2_X1 U17609 ( .A1(n14135), .A2(n14134), .ZN(P1_U2959) );
  AOI22_X1 U17610 ( .A1(n20239), .A2(P1_EAX_REG_19__SCAN_IN), .B1(n20238), 
        .B2(P1_UWORD_REG_3__SCAN_IN), .ZN(n14136) );
  NAND2_X1 U17611 ( .A1(n20224), .A2(n20332), .ZN(n14144) );
  NAND2_X1 U17612 ( .A1(n14136), .A2(n14144), .ZN(P1_U2940) );
  AOI22_X1 U17613 ( .A1(n20239), .A2(P1_EAX_REG_6__SCAN_IN), .B1(n20238), .B2(
        P1_LWORD_REG_6__SCAN_IN), .ZN(n14139) );
  NAND2_X1 U17614 ( .A1(n20305), .A2(DATAI_6_), .ZN(n14138) );
  NAND2_X1 U17615 ( .A1(n20303), .A2(BUF1_REG_6__SCAN_IN), .ZN(n14137) );
  AND2_X1 U17616 ( .A1(n14138), .A2(n14137), .ZN(n15076) );
  NAND2_X1 U17617 ( .A1(n20224), .A2(n20342), .ZN(n14152) );
  NAND2_X1 U17618 ( .A1(n14139), .A2(n14152), .ZN(P1_U2958) );
  AOI22_X1 U17619 ( .A1(n20239), .A2(P1_EAX_REG_21__SCAN_IN), .B1(n20238), 
        .B2(P1_UWORD_REG_5__SCAN_IN), .ZN(n14140) );
  INV_X1 U17620 ( .A(n15081), .ZN(n20338) );
  NAND2_X1 U17621 ( .A1(n20224), .A2(n20338), .ZN(n14146) );
  NAND2_X1 U17622 ( .A1(n14140), .A2(n14146), .ZN(P1_U2942) );
  AOI22_X1 U17623 ( .A1(n20239), .A2(P1_EAX_REG_17__SCAN_IN), .B1(n20238), 
        .B2(P1_UWORD_REG_1__SCAN_IN), .ZN(n14141) );
  NAND2_X1 U17624 ( .A1(n20224), .A2(n20325), .ZN(n14154) );
  NAND2_X1 U17625 ( .A1(n14141), .A2(n14154), .ZN(P1_U2938) );
  AOI22_X1 U17626 ( .A1(n20239), .A2(P1_EAX_REG_18__SCAN_IN), .B1(n20238), 
        .B2(P1_UWORD_REG_2__SCAN_IN), .ZN(n14143) );
  INV_X1 U17627 ( .A(n20328), .ZN(n14142) );
  NAND2_X1 U17628 ( .A1(n20224), .A2(n14142), .ZN(n14150) );
  NAND2_X1 U17629 ( .A1(n14143), .A2(n14150), .ZN(P1_U2939) );
  AOI22_X1 U17630 ( .A1(n20239), .A2(P1_EAX_REG_3__SCAN_IN), .B1(n20238), .B2(
        P1_LWORD_REG_3__SCAN_IN), .ZN(n14145) );
  NAND2_X1 U17631 ( .A1(n14145), .A2(n14144), .ZN(P1_U2955) );
  AOI22_X1 U17632 ( .A1(n20239), .A2(P1_EAX_REG_5__SCAN_IN), .B1(n20238), .B2(
        P1_LWORD_REG_5__SCAN_IN), .ZN(n14147) );
  NAND2_X1 U17633 ( .A1(n14147), .A2(n14146), .ZN(P1_U2957) );
  AOI22_X1 U17634 ( .A1(n20239), .A2(P1_EAX_REG_0__SCAN_IN), .B1(n20238), .B2(
        P1_LWORD_REG_0__SCAN_IN), .ZN(n14149) );
  NAND2_X1 U17635 ( .A1(n14149), .A2(n14148), .ZN(P1_U2952) );
  AOI22_X1 U17636 ( .A1(n20239), .A2(P1_EAX_REG_2__SCAN_IN), .B1(n20238), .B2(
        P1_LWORD_REG_2__SCAN_IN), .ZN(n14151) );
  NAND2_X1 U17637 ( .A1(n14151), .A2(n14150), .ZN(P1_U2954) );
  AOI22_X1 U17638 ( .A1(n20239), .A2(P1_EAX_REG_22__SCAN_IN), .B1(n20238), 
        .B2(P1_UWORD_REG_6__SCAN_IN), .ZN(n14153) );
  NAND2_X1 U17639 ( .A1(n14153), .A2(n14152), .ZN(P1_U2943) );
  AOI22_X1 U17640 ( .A1(n20239), .A2(P1_EAX_REG_1__SCAN_IN), .B1(n20238), .B2(
        P1_LWORD_REG_1__SCAN_IN), .ZN(n14155) );
  NAND2_X1 U17641 ( .A1(n14155), .A2(n14154), .ZN(P1_U2953) );
  INV_X1 U17642 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n14167) );
  NOR2_X1 U17643 ( .A1(n19159), .A2(n14156), .ZN(n14157) );
  XNOR2_X1 U17644 ( .A(n14157), .B(n16542), .ZN(n14158) );
  NAND2_X1 U17645 ( .A1(n14158), .A2(n19175), .ZN(n14166) );
  INV_X1 U17646 ( .A(n14159), .ZN(n16578) );
  AOI21_X1 U17647 ( .B1(n14160), .B2(n14415), .A(n9877), .ZN(n19251) );
  INV_X1 U17648 ( .A(n19251), .ZN(n16572) );
  AOI22_X1 U17649 ( .A1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n19166), .B1(
        P2_EBX_REG_8__SCAN_IN), .B2(n19205), .ZN(n14161) );
  OAI211_X1 U17650 ( .C1(n19200), .C2(n16572), .A(n14161), .B(n19345), .ZN(
        n14164) );
  NOR2_X1 U17651 ( .A1(n19202), .A2(n14162), .ZN(n14163) );
  AOI211_X1 U17652 ( .C1(n16578), .C2(n19179), .A(n14164), .B(n14163), .ZN(
        n14165) );
  OAI211_X1 U17653 ( .C1(n14167), .C2(n19181), .A(n14166), .B(n14165), .ZN(
        P2_U2847) );
  INV_X1 U17654 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n14180) );
  NOR2_X1 U17655 ( .A1(n19159), .A2(n14168), .ZN(n14169) );
  XNOR2_X1 U17656 ( .A(n14169), .B(n16523), .ZN(n14170) );
  NAND2_X1 U17657 ( .A1(n14170), .A2(n19175), .ZN(n14179) );
  AOI21_X1 U17658 ( .B1(n14172), .B2(n14171), .A(n16075), .ZN(n19245) );
  INV_X1 U17659 ( .A(n19245), .ZN(n14174) );
  AOI22_X1 U17660 ( .A1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n19166), .B1(
        P2_EBX_REG_10__SCAN_IN), .B2(n19205), .ZN(n14173) );
  OAI211_X1 U17661 ( .C1(n19200), .C2(n14174), .A(n14173), .B(n19345), .ZN(
        n14177) );
  NOR2_X1 U17662 ( .A1(n14175), .A2(n19202), .ZN(n14176) );
  AOI211_X1 U17663 ( .C1(n16519), .C2(n19179), .A(n14177), .B(n14176), .ZN(
        n14178) );
  OAI211_X1 U17664 ( .C1(n19181), .C2(n14180), .A(n14179), .B(n14178), .ZN(
        P2_U2845) );
  INV_X1 U17665 ( .A(n19324), .ZN(n14184) );
  NOR2_X1 U17666 ( .A1(n19159), .A2(n14181), .ZN(n14183) );
  AOI21_X1 U17667 ( .B1(n14184), .B2(n14183), .A(n19214), .ZN(n14182) );
  OAI21_X1 U17668 ( .B1(n14184), .B2(n14183), .A(n14182), .ZN(n14194) );
  NOR2_X1 U17669 ( .A1(n19200), .A2(n14185), .ZN(n14186) );
  AOI211_X1 U17670 ( .C1(n19166), .C2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n19170), .B(n14186), .ZN(n14187) );
  OAI21_X1 U17671 ( .B1(n14188), .B2(n19155), .A(n14187), .ZN(n14189) );
  AOI21_X1 U17672 ( .B1(n14190), .B2(n19186), .A(n14189), .ZN(n14191) );
  OAI21_X1 U17673 ( .B1(n21299), .B2(n19181), .A(n14191), .ZN(n14192) );
  AOI21_X1 U17674 ( .B1(n19179), .B2(n19316), .A(n14192), .ZN(n14193) );
  OAI211_X1 U17675 ( .C1(n19208), .C2(n19259), .A(n14194), .B(n14193), .ZN(
        P2_U2851) );
  NOR2_X1 U17676 ( .A1(n19159), .A2(n14195), .ZN(n16113) );
  XNOR2_X1 U17677 ( .A(n16113), .B(n14796), .ZN(n14196) );
  NAND2_X1 U17678 ( .A1(n14196), .A2(n19175), .ZN(n14204) );
  INV_X1 U17679 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n19936) );
  OAI22_X1 U17680 ( .A1(n19155), .A2(n14197), .B1(n19936), .B2(n19181), .ZN(
        n14198) );
  AOI21_X1 U17681 ( .B1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n19166), .A(
        n14198), .ZN(n14200) );
  NAND2_X1 U17682 ( .A1(n20021), .A2(n19183), .ZN(n14199) );
  OAI211_X1 U17683 ( .C1(n19202), .C2(n14201), .A(n14200), .B(n14199), .ZN(
        n14202) );
  AOI21_X1 U17684 ( .B1(n19342), .B2(n19179), .A(n14202), .ZN(n14203) );
  OAI211_X1 U17685 ( .C1(n20018), .C2(n19208), .A(n14204), .B(n14203), .ZN(
        P2_U2853) );
  AOI22_X1 U17686 ( .A1(n14599), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n14598), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n14212) );
  AOI22_X1 U17687 ( .A1(n14579), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n10673), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n14211) );
  OR2_X1 U17688 ( .A1(n14601), .A2(n14207), .ZN(n14210) );
  INV_X1 U17689 ( .A(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n14208) );
  OR2_X1 U17690 ( .A1(n14603), .A2(n14208), .ZN(n14209) );
  AND4_X1 U17691 ( .A1(n14212), .A2(n14211), .A3(n14210), .A4(n14209), .ZN(
        n14217) );
  INV_X1 U17692 ( .A(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n14213) );
  INV_X1 U17693 ( .A(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n14344) );
  OAI22_X1 U17694 ( .A1(n14610), .A2(n14213), .B1(n14609), .B2(n14344), .ZN(
        n14214) );
  INV_X1 U17695 ( .A(n14214), .ZN(n14216) );
  AOI22_X1 U17696 ( .A1(n14614), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n14613), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n14215) );
  NAND3_X1 U17697 ( .A1(n14217), .A2(n14216), .A3(n14215), .ZN(n14222) );
  AOI22_X1 U17698 ( .A1(n10674), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n10667), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n14220) );
  AOI22_X1 U17699 ( .A1(n10665), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n14618), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n14219) );
  AOI22_X1 U17700 ( .A1(n10485), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n10496), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n14218) );
  NAND3_X1 U17701 ( .A1(n14220), .A2(n14219), .A3(n14218), .ZN(n14221) );
  NOR2_X1 U17702 ( .A1(n14222), .A2(n14221), .ZN(n14255) );
  AOI22_X1 U17703 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n14599), .B1(
        n14598), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n14228) );
  AOI22_X1 U17704 ( .A1(n14579), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n10673), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n14227) );
  OR2_X1 U17705 ( .A1(n14601), .A2(n14223), .ZN(n14226) );
  INV_X1 U17706 ( .A(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n14224) );
  OR2_X1 U17707 ( .A1(n14603), .A2(n14224), .ZN(n14225) );
  NAND4_X1 U17708 ( .A1(n14228), .A2(n14227), .A3(n14226), .A4(n14225), .ZN(
        n14236) );
  INV_X1 U17709 ( .A(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n14229) );
  OR2_X1 U17710 ( .A1(n14610), .A2(n14229), .ZN(n14234) );
  INV_X1 U17711 ( .A(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n14230) );
  OR2_X1 U17712 ( .A1(n14609), .A2(n14230), .ZN(n14233) );
  NAND2_X1 U17713 ( .A1(n14614), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n14232) );
  NAND2_X1 U17714 ( .A1(n14613), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n14231) );
  NAND4_X1 U17715 ( .A1(n14234), .A2(n14233), .A3(n14232), .A4(n14231), .ZN(
        n14235) );
  NOR2_X1 U17716 ( .A1(n14236), .A2(n14235), .ZN(n14240) );
  AOI22_X1 U17717 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n10674), .B1(
        n10667), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n14239) );
  AOI22_X1 U17718 ( .A1(n10665), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n14618), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n14238) );
  AOI22_X1 U17719 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n10496), .B1(
        n10485), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n14237) );
  NAND4_X1 U17720 ( .A1(n14240), .A2(n14239), .A3(n14238), .A4(n14237), .ZN(
        n14241) );
  INV_X1 U17721 ( .A(n14363), .ZN(n14435) );
  OAI21_X1 U17722 ( .B1(n9945), .B2(n14241), .A(n14435), .ZN(n14406) );
  OAI21_X1 U17723 ( .B1(n14445), .B2(n14243), .A(n14242), .ZN(n19080) );
  NOR2_X2 U17724 ( .A1(n14244), .A2(n14302), .ZN(n19223) );
  NOR2_X2 U17725 ( .A1(n14244), .A2(n14303), .ZN(n19222) );
  AOI22_X1 U17726 ( .A1(n19223), .A2(BUF2_REG_17__SCAN_IN), .B1(n19222), .B2(
        BUF1_REG_17__SCAN_IN), .ZN(n14246) );
  AOI22_X1 U17727 ( .A1(n19221), .A2(n14306), .B1(n19257), .B2(
        P2_EAX_REG_17__SCAN_IN), .ZN(n14245) );
  OAI211_X1 U17728 ( .C1(n19229), .C2(n19080), .A(n14246), .B(n14245), .ZN(
        n14247) );
  INV_X1 U17729 ( .A(n14247), .ZN(n14248) );
  OAI21_X1 U17730 ( .B1(n14406), .B2(n19258), .A(n14248), .ZN(P2_U2902) );
  XOR2_X1 U17731 ( .A(n14020), .B(n14249), .Z(n20132) );
  INV_X1 U17732 ( .A(n20132), .ZN(n14261) );
  OAI222_X1 U17733 ( .A1(n15118), .A2(n14261), .B1(n15090), .B2(n12029), .C1(
        n15116), .C2(n15076), .ZN(P1_U2898) );
  OR2_X1 U17734 ( .A1(n14251), .A2(n14252), .ZN(n14253) );
  NAND2_X1 U17735 ( .A1(n14250), .A2(n14253), .ZN(n16493) );
  AND2_X1 U17736 ( .A1(n14254), .A2(n14255), .ZN(n14256) );
  NOR2_X1 U17737 ( .A1(n9945), .A2(n14256), .ZN(n19225) );
  NAND2_X1 U17738 ( .A1(n19225), .A2(n15685), .ZN(n14258) );
  NAND2_X1 U17739 ( .A1(n15661), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n14257) );
  OAI211_X1 U17740 ( .C1(n16493), .C2(n15661), .A(n14258), .B(n14257), .ZN(
        P2_U2871) );
  NAND2_X1 U17741 ( .A1(n16424), .A2(n14259), .ZN(n14260) );
  AND2_X1 U17742 ( .A1(n16408), .A2(n14260), .ZN(n16417) );
  INV_X1 U17743 ( .A(n16417), .ZN(n20125) );
  INV_X1 U17744 ( .A(P1_EBX_REG_6__SCAN_IN), .ZN(n20123) );
  OAI222_X1 U17745 ( .A1(n20175), .A2(n20125), .B1(n20182), .B2(n20123), .C1(
        n9828), .C2(n14261), .ZN(P1_U2866) );
  XNOR2_X1 U17746 ( .A(n14263), .B(n14262), .ZN(n16552) );
  AOI21_X1 U17747 ( .B1(n14267), .B2(n14265), .A(n14264), .ZN(n14266) );
  AOI21_X1 U17748 ( .B1(n11448), .B2(n14267), .A(n14266), .ZN(n16551) );
  OAI221_X1 U17749 ( .B1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .C1(n14270), .C2(n14269), .A(
        n14268), .ZN(n14271) );
  INV_X1 U17750 ( .A(n14271), .ZN(n14278) );
  XNOR2_X1 U17751 ( .A(n14273), .B(n14272), .ZN(n19263) );
  NAND2_X1 U17752 ( .A1(n19341), .A2(n19174), .ZN(n14276) );
  AOI22_X1 U17753 ( .A1(n19170), .A2(P2_REIP_REG_5__SCAN_IN), .B1(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n14274), .ZN(n14275) );
  OAI211_X1 U17754 ( .C1(n19263), .C2(n19327), .A(n14276), .B(n14275), .ZN(
        n14277) );
  AOI211_X1 U17755 ( .C1(n16551), .C2(n16577), .A(n14278), .B(n14277), .ZN(
        n14279) );
  OAI21_X1 U17756 ( .B1(n19363), .B2(n16552), .A(n14279), .ZN(P2_U3041) );
  INV_X1 U17757 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n14286) );
  OAI211_X1 U17758 ( .C1(n14281), .C2(n14206), .A(n15685), .B(n14254), .ZN(
        n14285) );
  NOR2_X1 U17759 ( .A1(n14026), .A2(n14282), .ZN(n14283) );
  OR2_X1 U17760 ( .A1(n14251), .A2(n14283), .ZN(n19091) );
  INV_X1 U17761 ( .A(n19091), .ZN(n16503) );
  NAND2_X1 U17762 ( .A1(n16503), .A2(n14287), .ZN(n14284) );
  OAI211_X1 U17763 ( .C1(n14287), .C2(n14286), .A(n14285), .B(n14284), .ZN(
        P2_U2872) );
  INV_X1 U17764 ( .A(n14289), .ZN(n14291) );
  NAND2_X1 U17765 ( .A1(n14291), .A2(n14290), .ZN(n14292) );
  AND2_X1 U17766 ( .A1(n14288), .A2(n14292), .ZN(n20172) );
  INV_X1 U17767 ( .A(n20172), .ZN(n14293) );
  OAI222_X1 U17768 ( .A1(n14293), .A2(n15118), .B1(n15071), .B2(n15116), .C1(
        n15090), .C2(n12035), .ZN(P1_U2897) );
  NOR2_X1 U17769 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n20017), .ZN(
        n19720) );
  NOR3_X2 U17770 ( .A1(n20043), .A2(n19717), .A3(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19692) );
  AOI221_X1 U17771 ( .B1(P2_STATEBS16_REG_SCAN_IN), .B2(n19710), .C1(
        P2_STATEBS16_REG_SCAN_IN), .C2(n19737), .A(n19692), .ZN(n14294) );
  AOI211_X1 U17772 ( .C1(P2_STATE2_REG_2__SCAN_IN), .C2(n14295), .A(
        P2_STATE2_REG_3__SCAN_IN), .B(n14294), .ZN(n14300) );
  NOR3_X2 U17773 ( .A1(n20033), .A2(n19717), .A3(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19708) );
  AND2_X1 U17774 ( .A1(n14296), .A2(n16225), .ZN(n14297) );
  OAI21_X1 U17775 ( .B1(n14300), .B2(n19708), .A(n19861), .ZN(n14301) );
  INV_X1 U17776 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n16664) );
  INV_X1 U17777 ( .A(BUF2_REG_17__SCAN_IN), .ZN(n18389) );
  OAI22_X2 U17778 ( .A1(n16664), .A2(n19424), .B1(n18389), .B2(n19422), .ZN(
        n19869) );
  INV_X1 U17779 ( .A(BUF2_REG_25__SCAN_IN), .ZN(n18390) );
  INV_X1 U17780 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n16654) );
  OAI22_X2 U17781 ( .A1(n18390), .A2(n19422), .B1(n16654), .B2(n19424), .ZN(
        n19818) );
  AOI22_X1 U17782 ( .A1(n19737), .A2(n19869), .B1(n19710), .B2(n19818), .ZN(
        n14308) );
  OAI21_X1 U17783 ( .B1(n11217), .B2(n19708), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n14305) );
  NAND2_X1 U17784 ( .A1(n14306), .A2(n19861), .ZN(n19821) );
  AOI22_X1 U17785 ( .A1(n19709), .A2(n19868), .B1(n19708), .B2(n19867), .ZN(
        n14307) );
  OAI211_X1 U17786 ( .C1(n19714), .C2(n14309), .A(n14308), .B(n14307), .ZN(
        P2_U3129) );
  INV_X1 U17787 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n16665) );
  INV_X1 U17788 ( .A(BUF2_REG_16__SCAN_IN), .ZN(n18384) );
  OAI22_X2 U17789 ( .A1(n16665), .A2(n19424), .B1(n18384), .B2(n19422), .ZN(
        n19863) );
  INV_X1 U17790 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n16656) );
  INV_X1 U17791 ( .A(BUF2_REG_24__SCAN_IN), .ZN(n18379) );
  OAI22_X2 U17792 ( .A1(n16656), .A2(n19424), .B1(n18379), .B2(n19422), .ZN(
        n19808) );
  AOI22_X1 U17793 ( .A1(n19737), .A2(n19863), .B1(n19710), .B2(n19808), .ZN(
        n14311) );
  NAND2_X1 U17794 ( .A1(n19220), .A2(n19861), .ZN(n19817) );
  AOI22_X1 U17795 ( .A1(n19709), .A2(n19856), .B1(n19855), .B2(n19708), .ZN(
        n14310) );
  OAI211_X1 U17796 ( .C1(n19714), .C2(n14312), .A(n14311), .B(n14310), .ZN(
        P2_U3128) );
  NAND2_X1 U17797 ( .A1(n11222), .A2(n20036), .ZN(n14314) );
  NOR2_X1 U17798 ( .A1(n19539), .A2(n19637), .ZN(n19533) );
  NOR2_X1 U17799 ( .A1(n19533), .A2(n20006), .ZN(n14313) );
  NAND2_X1 U17800 ( .A1(n14314), .A2(n14313), .ZN(n14320) );
  OAI21_X1 U17801 ( .B1(n19535), .B2(n19563), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n14317) );
  INV_X1 U17802 ( .A(n14315), .ZN(n19569) );
  NOR2_X1 U17803 ( .A1(n19569), .A2(n14316), .ZN(n14338) );
  NAND2_X1 U17804 ( .A1(n14338), .A2(n20017), .ZN(n14322) );
  NAND2_X1 U17805 ( .A1(n14317), .A2(n14322), .ZN(n14318) );
  AND2_X1 U17806 ( .A1(n19861), .A2(n14318), .ZN(n14319) );
  INV_X1 U17807 ( .A(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n14327) );
  OAI21_X1 U17808 ( .B1(n11222), .B2(n19533), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n14321) );
  INV_X1 U17809 ( .A(n19867), .ZN(n14324) );
  INV_X1 U17810 ( .A(n19533), .ZN(n14329) );
  AOI22_X1 U17811 ( .A1(n19563), .A2(n19869), .B1(n19535), .B2(n19818), .ZN(
        n14323) );
  OAI21_X1 U17812 ( .B1(n14324), .B2(n14329), .A(n14323), .ZN(n14325) );
  AOI21_X1 U17813 ( .B1(n19534), .B2(n19868), .A(n14325), .ZN(n14326) );
  OAI21_X1 U17814 ( .B1(n19523), .B2(n14327), .A(n14326), .ZN(P2_U3081) );
  INV_X1 U17815 ( .A(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n14333) );
  INV_X1 U17816 ( .A(n19855), .ZN(n14330) );
  AOI22_X1 U17817 ( .A1(n19563), .A2(n19863), .B1(n19535), .B2(n19808), .ZN(
        n14328) );
  OAI21_X1 U17818 ( .B1(n14330), .B2(n14329), .A(n14328), .ZN(n14331) );
  AOI21_X1 U17819 ( .B1(n19534), .B2(n19856), .A(n14331), .ZN(n14332) );
  OAI21_X1 U17820 ( .B1(n19523), .B2(n14333), .A(n14332), .ZN(P2_U3080) );
  NAND3_X1 U17821 ( .A1(n20033), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19779) );
  NOR2_X1 U17822 ( .A1(n19779), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n19767) );
  INV_X1 U17823 ( .A(n19767), .ZN(n14337) );
  OAI21_X1 U17824 ( .B1(n11225), .B2(n20034), .A(n20036), .ZN(n14336) );
  AOI21_X1 U17825 ( .B1(n19763), .B2(n19801), .A(n20061), .ZN(n14334) );
  AOI21_X1 U17826 ( .B1(n14338), .B2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(
        n14334), .ZN(n14335) );
  AOI211_X1 U17827 ( .C1(n14337), .C2(n14336), .A(n19610), .B(n14335), .ZN(
        n19750) );
  AOI22_X1 U17828 ( .A1(n19760), .A2(n19863), .B1(n19769), .B2(n19808), .ZN(
        n14343) );
  INV_X1 U17829 ( .A(n14338), .ZN(n14340) );
  OAI21_X1 U17830 ( .B1(n11225), .B2(n19767), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n14339) );
  OAI21_X1 U17831 ( .B1(n14341), .B2(n14340), .A(n14339), .ZN(n19768) );
  AOI22_X1 U17832 ( .A1(n19768), .A2(n19856), .B1(n19855), .B2(n19767), .ZN(
        n14342) );
  OAI211_X1 U17833 ( .C1(n19750), .C2(n14344), .A(n14343), .B(n14342), .ZN(
        P2_U3144) );
  AOI22_X1 U17834 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n14599), .B1(
        n14598), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n14350) );
  AOI22_X1 U17835 ( .A1(n14579), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n10673), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n14349) );
  OR2_X1 U17836 ( .A1(n14601), .A2(n14345), .ZN(n14348) );
  INV_X1 U17837 ( .A(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n14346) );
  OR2_X1 U17838 ( .A1(n14603), .A2(n14346), .ZN(n14347) );
  NAND4_X1 U17839 ( .A1(n14350), .A2(n14349), .A3(n14348), .A4(n14347), .ZN(
        n14358) );
  INV_X1 U17840 ( .A(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n14351) );
  OR2_X1 U17841 ( .A1(n14610), .A2(n14351), .ZN(n14356) );
  INV_X1 U17842 ( .A(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n14352) );
  OR2_X1 U17843 ( .A1(n14609), .A2(n14352), .ZN(n14355) );
  NAND2_X1 U17844 ( .A1(n14614), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n14354) );
  NAND2_X1 U17845 ( .A1(n14613), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n14353) );
  NAND4_X1 U17846 ( .A1(n14356), .A2(n14355), .A3(n14354), .A4(n14353), .ZN(
        n14357) );
  NOR2_X1 U17847 ( .A1(n14358), .A2(n14357), .ZN(n14362) );
  AOI22_X1 U17848 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n10674), .B1(
        n10667), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n14361) );
  AOI22_X1 U17849 ( .A1(n10665), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n14618), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n14360) );
  AOI22_X1 U17850 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n10496), .B1(
        n10485), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n14359) );
  NAND4_X1 U17851 ( .A1(n14362), .A2(n14361), .A3(n14360), .A4(n14359), .ZN(
        n14434) );
  AOI22_X1 U17852 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n14599), .B1(
        n14598), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n14369) );
  AOI22_X1 U17853 ( .A1(n14579), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n10673), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n14368) );
  OR2_X1 U17854 ( .A1(n14601), .A2(n14364), .ZN(n14367) );
  INV_X1 U17855 ( .A(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n14365) );
  OR2_X1 U17856 ( .A1(n14603), .A2(n14365), .ZN(n14366) );
  AND4_X1 U17857 ( .A1(n14369), .A2(n14368), .A3(n14367), .A4(n14366), .ZN(
        n14375) );
  INV_X1 U17858 ( .A(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n14371) );
  INV_X1 U17859 ( .A(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n14370) );
  OAI22_X1 U17860 ( .A1(n14371), .A2(n14610), .B1(n14609), .B2(n14370), .ZN(
        n14372) );
  INV_X1 U17861 ( .A(n14372), .ZN(n14374) );
  AOI22_X1 U17862 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n14614), .B1(
        n14613), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n14373) );
  NAND3_X1 U17863 ( .A1(n14375), .A2(n14374), .A3(n14373), .ZN(n14380) );
  AOI22_X1 U17864 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n10674), .B1(
        n10667), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n14378) );
  AOI22_X1 U17865 ( .A1(n10665), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n14618), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n14377) );
  AOI22_X1 U17866 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n10496), .B1(
        n10485), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n14376) );
  NAND3_X1 U17867 ( .A1(n14378), .A2(n14377), .A3(n14376), .ZN(n14379) );
  OAI21_X1 U17868 ( .B1(n9947), .B2(n10371), .A(n14543), .ZN(n15695) );
  XNOR2_X1 U17869 ( .A(n15604), .B(n14381), .ZN(n19068) );
  AOI22_X1 U17870 ( .A1(n19223), .A2(BUF2_REG_19__SCAN_IN), .B1(n19222), .B2(
        BUF1_REG_19__SCAN_IN), .ZN(n14384) );
  INV_X1 U17871 ( .A(n14382), .ZN(n19388) );
  AOI22_X1 U17872 ( .A1(n19221), .A2(n19388), .B1(n19257), .B2(
        P2_EAX_REG_19__SCAN_IN), .ZN(n14383) );
  OAI211_X1 U17873 ( .C1(n19068), .C2(n19229), .A(n14384), .B(n14383), .ZN(
        n14385) );
  INV_X1 U17874 ( .A(n14385), .ZN(n14386) );
  OAI21_X1 U17875 ( .B1(n15695), .B2(n19258), .A(n14386), .ZN(P2_U2900) );
  NAND2_X1 U17876 ( .A1(n14288), .A2(n14388), .ZN(n14389) );
  NAND2_X1 U17877 ( .A1(n14387), .A2(n14389), .ZN(n14476) );
  INV_X1 U17878 ( .A(n14472), .ZN(n14390) );
  AOI22_X1 U17879 ( .A1(n20154), .A2(n14390), .B1(P1_EBX_REG_8__SCAN_IN), .B2(
        n20147), .ZN(n14391) );
  OAI211_X1 U17880 ( .C1(n20158), .C2(n14392), .A(n14391), .B(n20256), .ZN(
        n14397) );
  NOR3_X1 U17881 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(n20151), .A3(n14393), .ZN(
        n14396) );
  XNOR2_X1 U17882 ( .A(n16410), .B(n14505), .ZN(n16395) );
  AND2_X1 U17883 ( .A1(n20117), .A2(n14461), .ZN(n14954) );
  NOR2_X1 U17884 ( .A1(n14954), .A2(n14958), .ZN(n20108) );
  NAND2_X1 U17885 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(n20108), .ZN(n14394) );
  OAI21_X1 U17886 ( .B1(n16395), .B2(n20124), .A(n14394), .ZN(n14395) );
  NOR3_X1 U17887 ( .A1(n14397), .A2(n14396), .A3(n14395), .ZN(n14398) );
  OAI21_X1 U17888 ( .B1(n14476), .B2(n14988), .A(n14398), .ZN(P1_U2832) );
  INV_X1 U17889 ( .A(DATAI_8_), .ZN(n14399) );
  MUX2_X1 U17890 ( .A(n14399), .B(n16677), .S(n20303), .Z(n20210) );
  INV_X1 U17891 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n14400) );
  OAI222_X1 U17892 ( .A1(n14476), .A2(n15118), .B1(n20210), .B2(n15116), .C1(
        n14400), .C2(n15090), .ZN(P1_U2896) );
  INV_X1 U17893 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n14401) );
  OAI222_X1 U17894 ( .A1(n9828), .A2(n14476), .B1(n14401), .B2(n20182), .C1(
        n20175), .C2(n16395), .ZN(P1_U2864) );
  NAND2_X1 U17895 ( .A1(n15661), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n14405) );
  INV_X1 U17896 ( .A(n14432), .ZN(n14402) );
  AOI21_X1 U17897 ( .B1(n14403), .B2(n14250), .A(n14402), .ZN(n19082) );
  NAND2_X1 U17898 ( .A1(n19082), .A2(n14287), .ZN(n14404) );
  OAI211_X1 U17899 ( .C1(n14406), .C2(n15694), .A(n14405), .B(n14404), .ZN(
        P2_U2870) );
  XNOR2_X1 U17900 ( .A(n14408), .B(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n14409) );
  XNOR2_X1 U17901 ( .A(n14407), .B(n14409), .ZN(n14430) );
  NAND2_X1 U17902 ( .A1(n16532), .A2(n16534), .ZN(n14411) );
  XNOR2_X1 U17903 ( .A(n14410), .B(n14411), .ZN(n14428) );
  INV_X1 U17904 ( .A(n14412), .ZN(n16581) );
  NAND2_X1 U17905 ( .A1(n16581), .A2(n14421), .ZN(n14420) );
  INV_X1 U17906 ( .A(n19148), .ZN(n14418) );
  OR2_X1 U17907 ( .A1(n14414), .A2(n14413), .ZN(n14416) );
  NAND2_X1 U17908 ( .A1(n14416), .A2(n14415), .ZN(n19253) );
  INV_X1 U17909 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n19945) );
  OAI22_X1 U17910 ( .A1(n19327), .A2(n19253), .B1(n19945), .B2(n19345), .ZN(
        n14417) );
  AOI21_X1 U17911 ( .B1(n19341), .B2(n14418), .A(n14417), .ZN(n14419) );
  OAI211_X1 U17912 ( .C1(n16574), .C2(n14421), .A(n14420), .B(n14419), .ZN(
        n14422) );
  AOI21_X1 U17913 ( .B1(n14428), .B2(n19331), .A(n14422), .ZN(n14423) );
  OAI21_X1 U17914 ( .B1(n14430), .B2(n19356), .A(n14423), .ZN(P2_U3039) );
  OAI22_X1 U17915 ( .A1(n16559), .A2(n14424), .B1(n19945), .B2(n19345), .ZN(
        n14427) );
  INV_X1 U17916 ( .A(n19143), .ZN(n14425) );
  OAI22_X1 U17917 ( .A1(n16545), .A2(n19148), .B1(n19325), .B2(n14425), .ZN(
        n14426) );
  AOI211_X1 U17918 ( .C1(n14428), .C2(n12840), .A(n14427), .B(n14426), .ZN(
        n14429) );
  OAI21_X1 U17919 ( .B1(n14430), .B2(n19319), .A(n14429), .ZN(P2_U3007) );
  NAND2_X1 U17920 ( .A1(n14432), .A2(n14431), .ZN(n14433) );
  INV_X1 U17921 ( .A(n16486), .ZN(n14439) );
  INV_X1 U17922 ( .A(n14434), .ZN(n14436) );
  AOI21_X1 U17923 ( .B1(n14436), .B2(n14435), .A(n9947), .ZN(n16468) );
  NAND2_X1 U17924 ( .A1(n16468), .A2(n15685), .ZN(n14438) );
  NAND2_X1 U17925 ( .A1(n15661), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n14437) );
  OAI211_X1 U17926 ( .C1(n14439), .C2(n15661), .A(n14438), .B(n14437), .ZN(
        P2_U2869) );
  NOR2_X1 U17927 ( .A1(n19159), .A2(n14440), .ZN(n14441) );
  XNOR2_X1 U17928 ( .A(n14441), .B(n16499), .ZN(n14454) );
  INV_X1 U17929 ( .A(n16493), .ZN(n14449) );
  NOR2_X1 U17930 ( .A1(n14443), .A2(n14442), .ZN(n14444) );
  NOR2_X1 U17931 ( .A1(n14445), .A2(n14444), .ZN(n19224) );
  NAND2_X1 U17932 ( .A1(n19183), .A2(n19224), .ZN(n14447) );
  AOI22_X1 U17933 ( .A1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n19166), .B1(
        P2_EBX_REG_16__SCAN_IN), .B2(n19205), .ZN(n14446) );
  NAND3_X1 U17934 ( .A1(n14447), .A2(n14446), .A3(n19345), .ZN(n14448) );
  AOI21_X1 U17935 ( .B1(n14449), .B2(n19179), .A(n14448), .ZN(n14451) );
  NAND2_X1 U17936 ( .A1(n19210), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n14450) );
  OAI211_X1 U17937 ( .C1(n14452), .C2(n19202), .A(n14451), .B(n14450), .ZN(
        n14453) );
  AOI21_X1 U17938 ( .B1(n14454), .B2(n19175), .A(n14453), .ZN(n14455) );
  INV_X1 U17939 ( .A(n14455), .ZN(P2_U2839) );
  OAI21_X1 U17940 ( .B1(n14456), .B2(n14458), .A(n14457), .ZN(n15273) );
  XNOR2_X1 U17941 ( .A(n15040), .B(n15042), .ZN(n16386) );
  AOI22_X1 U17942 ( .A1(n16386), .A2(n20171), .B1(P1_EBX_REG_10__SCAN_IN), 
        .B2(n15032), .ZN(n14459) );
  OAI21_X1 U17943 ( .B1(n15273), .B2(n9828), .A(n14459), .ZN(P1_U2862) );
  INV_X1 U17944 ( .A(P1_REIP_REG_10__SCAN_IN), .ZN(n20942) );
  INV_X1 U17945 ( .A(P1_REIP_REG_9__SCAN_IN), .ZN(n20940) );
  NOR2_X1 U17946 ( .A1(n20942), .A2(n20940), .ZN(n14460) );
  AOI21_X1 U17947 ( .B1(n14460), .B2(n14954), .A(n14958), .ZN(n16289) );
  NAND2_X1 U17948 ( .A1(n20137), .A2(n14461), .ZN(n20105) );
  NOR2_X1 U17949 ( .A1(n20940), .A2(n20105), .ZN(n16285) );
  NAND2_X1 U17950 ( .A1(n16285), .A2(n20942), .ZN(n14466) );
  AOI21_X1 U17951 ( .B1(n20140), .B2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n20280), .ZN(n14462) );
  OAI21_X1 U17952 ( .B1(n20122), .B2(n14463), .A(n14462), .ZN(n14464) );
  AOI21_X1 U17953 ( .B1(n16386), .B2(n20149), .A(n14464), .ZN(n14465) );
  OAI211_X1 U17954 ( .C1(n20143), .C2(n15269), .A(n14466), .B(n14465), .ZN(
        n14467) );
  AOI21_X1 U17955 ( .B1(P1_REIP_REG_10__SCAN_IN), .B2(n16289), .A(n14467), 
        .ZN(n14468) );
  OAI21_X1 U17956 ( .B1(n15273), .B2(n14988), .A(n14468), .ZN(P1_U2830) );
  XNOR2_X1 U17957 ( .A(n14470), .B(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n14471) );
  XNOR2_X1 U17958 ( .A(n14469), .B(n14471), .ZN(n16403) );
  NAND2_X1 U17959 ( .A1(n16403), .A2(n20248), .ZN(n14475) );
  AND2_X1 U17960 ( .A1(n20296), .A2(P1_REIP_REG_8__SCAN_IN), .ZN(n16396) );
  NOR2_X1 U17961 ( .A1(n20252), .A2(n14472), .ZN(n14473) );
  AOI211_X1 U17962 ( .C1(n20242), .C2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n16396), .B(n14473), .ZN(n14474) );
  OAI211_X1 U17963 ( .C1(n20306), .C2(n14476), .A(n14475), .B(n14474), .ZN(
        P1_U2991) );
  OAI21_X1 U17964 ( .B1(n14477), .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n14479), .ZN(n16543) );
  INV_X1 U17965 ( .A(n16546), .ZN(n19162) );
  XNOR2_X1 U17966 ( .A(n14481), .B(n14480), .ZN(n19256) );
  INV_X1 U17967 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n19943) );
  OAI22_X1 U17968 ( .A1(n19327), .A2(n19256), .B1(n19943), .B2(n19345), .ZN(
        n14482) );
  AOI21_X1 U17969 ( .B1(n19341), .B2(n19162), .A(n14482), .ZN(n14483) );
  OAI21_X1 U17970 ( .B1(n16574), .B2(n14488), .A(n14483), .ZN(n14487) );
  XNOR2_X1 U17971 ( .A(n14485), .B(n14484), .ZN(n16544) );
  NOR2_X1 U17972 ( .A1(n16544), .A2(n19363), .ZN(n14486) );
  AOI211_X1 U17973 ( .C1(n14489), .C2(n14488), .A(n14487), .B(n14486), .ZN(
        n14490) );
  OAI21_X1 U17974 ( .B1(n19356), .B2(n16543), .A(n14490), .ZN(P2_U3040) );
  INV_X1 U17975 ( .A(DATAI_10_), .ZN(n14492) );
  MUX2_X1 U17976 ( .A(n14492), .B(n14491), .S(n20303), .Z(n20216) );
  INV_X1 U17977 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n14493) );
  OAI222_X1 U17978 ( .A1(n15273), .A2(n15118), .B1(n20216), .B2(n15116), .C1(
        n14493), .C2(n15090), .ZN(P1_U2894) );
  NOR2_X1 U17979 ( .A1(n14456), .A2(n10379), .ZN(n20167) );
  INV_X1 U17980 ( .A(n20167), .ZN(n14498) );
  INV_X1 U17981 ( .A(DATAI_9_), .ZN(n14496) );
  MUX2_X1 U17982 ( .A(n14496), .B(n14495), .S(n20303), .Z(n20213) );
  INV_X1 U17983 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n14497) );
  OAI222_X1 U17984 ( .A1(n14498), .A2(n15118), .B1(n20213), .B2(n15116), .C1(
        n14497), .C2(n15090), .ZN(P1_U2895) );
  XNOR2_X1 U17985 ( .A(n9845), .B(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n14500) );
  XNOR2_X1 U17986 ( .A(n14499), .B(n14500), .ZN(n14515) );
  NOR2_X1 U17987 ( .A1(n20276), .A2(n20277), .ZN(n15313) );
  NOR2_X1 U17988 ( .A1(n20267), .A2(n20273), .ZN(n20262) );
  NOR2_X1 U17989 ( .A1(n14501), .A2(n20286), .ZN(n20260) );
  NAND2_X1 U17990 ( .A1(n20262), .A2(n20260), .ZN(n16399) );
  NOR2_X1 U17991 ( .A1(n16399), .A2(n16430), .ZN(n15448) );
  INV_X1 U17992 ( .A(n15448), .ZN(n14502) );
  NAND3_X1 U17993 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n15275) );
  NAND2_X1 U17994 ( .A1(n20262), .A2(n20261), .ZN(n16425) );
  NOR2_X1 U17995 ( .A1(n16430), .A2(n16425), .ZN(n16426) );
  INV_X1 U17996 ( .A(n20289), .ZN(n20253) );
  OAI21_X1 U17997 ( .B1(n16426), .B2(n20253), .A(n15284), .ZN(n16398) );
  AOI211_X1 U17998 ( .C1(n16400), .C2(n14502), .A(n15275), .B(n16398), .ZN(
        n14503) );
  NOR2_X1 U17999 ( .A1(n15313), .A2(n14503), .ZN(n16388) );
  NAND2_X1 U18000 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16394) );
  NAND2_X1 U18001 ( .A1(n16431), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n15366) );
  NAND2_X1 U18002 ( .A1(n20289), .A2(n16426), .ZN(n15385) );
  NAND2_X1 U18003 ( .A1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n15431), .ZN(
        n16415) );
  NOR2_X1 U18004 ( .A1(n16394), .A2(n16415), .ZN(n16389) );
  AOI22_X1 U18005 ( .A1(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n16388), .B1(
        n16389), .B2(n16390), .ZN(n14508) );
  AOI21_X1 U18006 ( .B1(n16410), .B2(n14505), .A(n14504), .ZN(n14506) );
  OR2_X1 U18007 ( .A1(n15040), .A2(n14506), .ZN(n20165) );
  INV_X1 U18008 ( .A(n20165), .ZN(n20103) );
  AND2_X1 U18009 ( .A1(n20296), .A2(P1_REIP_REG_9__SCAN_IN), .ZN(n14509) );
  AOI21_X1 U18010 ( .B1(n20103), .B2(n20282), .A(n14509), .ZN(n14507) );
  OAI211_X1 U18011 ( .C1(n14515), .C2(n20293), .A(n14508), .B(n14507), .ZN(
        P1_U3022) );
  INV_X1 U18012 ( .A(n14509), .ZN(n14511) );
  NAND2_X1 U18013 ( .A1(n20242), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n14510) );
  OAI211_X1 U18014 ( .C1(n20252), .C2(n14512), .A(n14511), .B(n14510), .ZN(
        n14513) );
  AOI21_X1 U18015 ( .B1(n20167), .B2(n16325), .A(n14513), .ZN(n14514) );
  OAI21_X1 U18016 ( .B1(n14515), .B2(n20088), .A(n14514), .ZN(P1_U2990) );
  INV_X1 U18017 ( .A(DATAI_12_), .ZN(n21101) );
  MUX2_X1 U18018 ( .A(n21101), .B(n16671), .S(n20303), .Z(n20219) );
  OAI22_X1 U18019 ( .A1(n15091), .A2(n20219), .B1(n13643), .B2(n15090), .ZN(
        n14517) );
  AOI21_X1 U18020 ( .B1(n16295), .B2(DATAI_28_), .A(n14517), .ZN(n14519) );
  NAND2_X1 U18021 ( .A1(n15105), .A2(BUF1_REG_28__SCAN_IN), .ZN(n14518) );
  OAI211_X1 U18022 ( .C1(n14516), .C2(n15118), .A(n14519), .B(n14518), .ZN(
        P1_U2876) );
  INV_X1 U18023 ( .A(P1_EBX_REG_28__SCAN_IN), .ZN(n14521) );
  OAI21_X1 U18024 ( .B1(n14835), .B2(n14520), .A(n9867), .ZN(n14522) );
  OAI222_X1 U18025 ( .A1(n9828), .A2(n14516), .B1(n14521), .B2(n20182), .C1(
        n14522), .C2(n20175), .ZN(P1_U2844) );
  INV_X1 U18026 ( .A(n14522), .ZN(n15329) );
  INV_X1 U18027 ( .A(n14523), .ZN(n14527) );
  AOI22_X1 U18028 ( .A1(n20147), .A2(P1_EBX_REG_28__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n20140), .ZN(n14526) );
  INV_X1 U18029 ( .A(n14828), .ZN(n14524) );
  OAI21_X1 U18030 ( .B1(P1_REIP_REG_28__SCAN_IN), .B2(n14838), .A(n14524), 
        .ZN(n14525) );
  OAI211_X1 U18031 ( .C1(n20143), .C2(n14527), .A(n14526), .B(n14525), .ZN(
        n14528) );
  AOI21_X1 U18032 ( .B1(n15329), .B2(n20149), .A(n14528), .ZN(n14529) );
  OAI21_X1 U18033 ( .B1(n14516), .B2(n14988), .A(n14529), .ZN(P1_U2812) );
  INV_X1 U18034 ( .A(n14530), .ZN(n14531) );
  INV_X1 U18035 ( .A(n15859), .ZN(n16087) );
  OAI21_X1 U18036 ( .B1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n14530), .A(
        n16087), .ZN(n16525) );
  OAI21_X1 U18037 ( .B1(n14532), .B2(n9877), .A(n14171), .ZN(n19248) );
  INV_X1 U18038 ( .A(n19248), .ZN(n14534) );
  INV_X1 U18039 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n19948) );
  NOR2_X1 U18040 ( .A1(n19948), .A2(n19345), .ZN(n14533) );
  AOI21_X1 U18041 ( .B1(n19347), .B2(n14534), .A(n14533), .ZN(n14536) );
  NAND2_X1 U18042 ( .A1(n19341), .A2(n19136), .ZN(n14535) );
  OAI211_X1 U18043 ( .C1(n16047), .C2(n16072), .A(n14536), .B(n14535), .ZN(
        n14537) );
  AOI21_X1 U18044 ( .B1(n16073), .B2(n16072), .A(n14537), .ZN(n14542) );
  NAND2_X1 U18045 ( .A1(n14538), .A2(n14539), .ZN(n16092) );
  NAND2_X1 U18046 ( .A1(n16089), .A2(n16090), .ZN(n14540) );
  XNOR2_X1 U18047 ( .A(n16092), .B(n14540), .ZN(n16524) );
  OR2_X1 U18048 ( .A1(n16524), .A2(n19363), .ZN(n14541) );
  OAI211_X1 U18049 ( .C1(n16525), .C2(n19356), .A(n14542), .B(n14541), .ZN(
        P2_U3037) );
  AOI22_X1 U18050 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n14599), .B1(
        n14598), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n14549) );
  AOI22_X1 U18051 ( .A1(n14579), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n10673), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n14548) );
  OR2_X1 U18052 ( .A1(n14601), .A2(n14544), .ZN(n14547) );
  INV_X1 U18053 ( .A(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n14545) );
  OR2_X1 U18054 ( .A1(n14603), .A2(n14545), .ZN(n14546) );
  AND4_X1 U18055 ( .A1(n14549), .A2(n14548), .A3(n14547), .A4(n14546), .ZN(
        n14555) );
  INV_X1 U18056 ( .A(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n14551) );
  INV_X1 U18057 ( .A(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n14550) );
  OAI22_X1 U18058 ( .A1(n14551), .A2(n14610), .B1(n14609), .B2(n14550), .ZN(
        n14552) );
  INV_X1 U18059 ( .A(n14552), .ZN(n14554) );
  AOI22_X1 U18060 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n14614), .B1(
        n14613), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n14553) );
  NAND3_X1 U18061 ( .A1(n14555), .A2(n14554), .A3(n14553), .ZN(n14560) );
  AOI22_X1 U18062 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n10674), .B1(
        n10667), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n14558) );
  AOI22_X1 U18063 ( .A1(n10665), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n14618), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n14557) );
  AOI22_X1 U18064 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n10496), .B1(
        n10485), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n14556) );
  NAND3_X1 U18065 ( .A1(n14558), .A2(n14557), .A3(n14556), .ZN(n14559) );
  NOR2_X1 U18066 ( .A1(n14560), .A2(n14559), .ZN(n15684) );
  AOI22_X1 U18067 ( .A1(n14599), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n14598), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n14567) );
  AOI22_X1 U18068 ( .A1(n14579), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10673), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n14566) );
  OR2_X1 U18069 ( .A1(n14601), .A2(n14562), .ZN(n14565) );
  INV_X1 U18070 ( .A(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n14563) );
  OR2_X1 U18071 ( .A1(n14603), .A2(n14563), .ZN(n14564) );
  AND4_X1 U18072 ( .A1(n14567), .A2(n14566), .A3(n14565), .A4(n14564), .ZN(
        n14573) );
  INV_X1 U18073 ( .A(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n14569) );
  INV_X1 U18074 ( .A(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n14568) );
  OAI22_X1 U18075 ( .A1(n14610), .A2(n14569), .B1(n14609), .B2(n14568), .ZN(
        n14570) );
  INV_X1 U18076 ( .A(n14570), .ZN(n14572) );
  AOI22_X1 U18077 ( .A1(n14614), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n14613), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n14571) );
  NAND3_X1 U18078 ( .A1(n14573), .A2(n14572), .A3(n14571), .ZN(n14578) );
  AOI22_X1 U18079 ( .A1(n10674), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n10667), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n14576) );
  AOI22_X1 U18080 ( .A1(n10665), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n14618), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n14575) );
  AOI22_X1 U18081 ( .A1(n10485), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10496), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n14574) );
  NAND3_X1 U18082 ( .A1(n14576), .A2(n14575), .A3(n14574), .ZN(n14577) );
  NOR2_X1 U18083 ( .A1(n14578), .A2(n14577), .ZN(n15679) );
  AOI22_X1 U18084 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n14599), .B1(
        n14598), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n14585) );
  AOI22_X1 U18085 ( .A1(n14579), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n10673), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n14584) );
  OR2_X1 U18086 ( .A1(n14601), .A2(n14580), .ZN(n14583) );
  INV_X1 U18087 ( .A(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n14581) );
  OR2_X1 U18088 ( .A1(n14603), .A2(n14581), .ZN(n14582) );
  NAND4_X1 U18089 ( .A1(n14585), .A2(n14584), .A3(n14583), .A4(n14582), .ZN(
        n14593) );
  INV_X1 U18090 ( .A(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n14586) );
  OR2_X1 U18091 ( .A1(n14610), .A2(n14586), .ZN(n14591) );
  INV_X1 U18092 ( .A(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n14587) );
  OR2_X1 U18093 ( .A1(n14609), .A2(n14587), .ZN(n14590) );
  NAND2_X1 U18094 ( .A1(n14614), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n14589) );
  NAND2_X1 U18095 ( .A1(n14613), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n14588) );
  NAND4_X1 U18096 ( .A1(n14591), .A2(n14590), .A3(n14589), .A4(n14588), .ZN(
        n14592) );
  NOR2_X1 U18097 ( .A1(n14593), .A2(n14592), .ZN(n14597) );
  AOI22_X1 U18098 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n10674), .B1(
        n10667), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n14596) );
  AOI22_X1 U18099 ( .A1(n10665), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n14618), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n14595) );
  AOI22_X1 U18100 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n10496), .B1(
        n10485), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n14594) );
  NAND4_X1 U18101 ( .A1(n14597), .A2(n14596), .A3(n14595), .A4(n14594), .ZN(
        n15671) );
  NAND2_X1 U18102 ( .A1(n15672), .A2(n15671), .ZN(n14642) );
  AOI22_X1 U18103 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n14599), .B1(
        n14598), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n14607) );
  AOI22_X1 U18104 ( .A1(n14579), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n10673), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n14606) );
  OR2_X1 U18105 ( .A1(n14601), .A2(n14600), .ZN(n14605) );
  INV_X1 U18106 ( .A(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n14602) );
  OR2_X1 U18107 ( .A1(n14603), .A2(n14602), .ZN(n14604) );
  AND4_X1 U18108 ( .A1(n14607), .A2(n14606), .A3(n14605), .A4(n14604), .ZN(
        n14617) );
  INV_X1 U18109 ( .A(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n14611) );
  INV_X1 U18110 ( .A(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n14608) );
  OAI22_X1 U18111 ( .A1(n14611), .A2(n14610), .B1(n14609), .B2(n14608), .ZN(
        n14612) );
  INV_X1 U18112 ( .A(n14612), .ZN(n14616) );
  AOI22_X1 U18113 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n14614), .B1(
        n14613), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n14615) );
  NAND3_X1 U18114 ( .A1(n14617), .A2(n14616), .A3(n14615), .ZN(n14623) );
  AOI22_X1 U18115 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n10674), .B1(
        n10667), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n14621) );
  AOI22_X1 U18116 ( .A1(n10665), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n14618), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n14620) );
  AOI22_X1 U18117 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n10496), .B1(
        n10485), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n14619) );
  NAND3_X1 U18118 ( .A1(n14621), .A2(n14620), .A3(n14619), .ZN(n14622) );
  NOR2_X1 U18119 ( .A1(n14623), .A2(n14622), .ZN(n14659) );
  AOI22_X1 U18120 ( .A1(n9855), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n9847), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n14632) );
  AND2_X1 U18121 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n14625) );
  OR2_X1 U18122 ( .A1(n14625), .A2(n14624), .ZN(n14773) );
  INV_X1 U18123 ( .A(n14773), .ZN(n14747) );
  NAND2_X1 U18124 ( .A1(n9843), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n14628) );
  NAND2_X1 U18125 ( .A1(n9859), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n14627) );
  AND3_X1 U18126 ( .A1(n14747), .A2(n14628), .A3(n14627), .ZN(n14631) );
  AOI22_X1 U18127 ( .A1(n14770), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n9854), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n14630) );
  AOI22_X1 U18128 ( .A1(n13678), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n10644), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n14629) );
  NAND4_X1 U18129 ( .A1(n14632), .A2(n14631), .A3(n14630), .A4(n14629), .ZN(
        n14640) );
  AOI22_X1 U18130 ( .A1(n9847), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n14770), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n14638) );
  AOI22_X1 U18131 ( .A1(n9855), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(n9857), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n14637) );
  AOI22_X1 U18132 ( .A1(n9843), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n10644), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n14636) );
  NAND2_X1 U18133 ( .A1(n13678), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n14634) );
  NAND2_X1 U18134 ( .A1(n10647), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n14633) );
  AND3_X1 U18135 ( .A1(n14634), .A2(n14773), .A3(n14633), .ZN(n14635) );
  NAND4_X1 U18136 ( .A1(n14638), .A2(n14637), .A3(n14636), .A4(n14635), .ZN(
        n14639) );
  NAND2_X1 U18137 ( .A1(n14640), .A2(n14639), .ZN(n14664) );
  NOR2_X1 U18138 ( .A1(n9839), .A2(n14664), .ZN(n14641) );
  XOR2_X1 U18139 ( .A(n14659), .B(n14641), .Z(n14665) );
  INV_X1 U18140 ( .A(n14664), .ZN(n14660) );
  NAND2_X1 U18141 ( .A1(n9839), .A2(n14660), .ZN(n15664) );
  NOR2_X2 U18142 ( .A1(n15665), .A2(n15664), .ZN(n15663) );
  INV_X1 U18143 ( .A(n14642), .ZN(n15673) );
  INV_X1 U18144 ( .A(n14665), .ZN(n14643) );
  AOI22_X1 U18145 ( .A1(n9855), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n9847), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n14650) );
  NAND2_X1 U18146 ( .A1(n13678), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n14646) );
  NAND2_X1 U18147 ( .A1(n9858), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n14645) );
  AND3_X1 U18148 ( .A1(n14747), .A2(n14646), .A3(n14645), .ZN(n14649) );
  AOI22_X1 U18149 ( .A1(n14770), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n9854), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n14648) );
  AOI22_X1 U18150 ( .A1(n9843), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n10644), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n14647) );
  NAND4_X1 U18151 ( .A1(n14650), .A2(n14649), .A3(n14648), .A4(n14647), .ZN(
        n14658) );
  AOI22_X1 U18152 ( .A1(n9855), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n10646), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n14656) );
  AOI22_X1 U18153 ( .A1(n14770), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n9854), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n14655) );
  AOI22_X1 U18154 ( .A1(n10645), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n9822), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n14654) );
  NAND2_X1 U18155 ( .A1(n9841), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n14652) );
  INV_X1 U18156 ( .A(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n19586) );
  NAND2_X1 U18157 ( .A1(n9859), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n14651) );
  AND3_X1 U18158 ( .A1(n14652), .A2(n14651), .A3(n14773), .ZN(n14653) );
  NAND4_X1 U18159 ( .A1(n14656), .A2(n14655), .A3(n14654), .A4(n14653), .ZN(
        n14657) );
  INV_X1 U18160 ( .A(n14659), .ZN(n14661) );
  AND2_X1 U18161 ( .A1(n14661), .A2(n14660), .ZN(n14662) );
  NAND2_X1 U18162 ( .A1(n14662), .A2(n14663), .ZN(n14666) );
  OAI211_X1 U18163 ( .C1(n14663), .C2(n14662), .A(n14723), .B(n14666), .ZN(
        n15657) );
  NAND2_X1 U18164 ( .A1(n9839), .A2(n14663), .ZN(n15659) );
  INV_X1 U18165 ( .A(n14666), .ZN(n14681) );
  AOI22_X1 U18166 ( .A1(n9855), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n9847), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n14672) );
  NAND2_X1 U18167 ( .A1(n13678), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n14668) );
  NAND2_X1 U18168 ( .A1(n9858), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n14667) );
  AND3_X1 U18169 ( .A1(n14747), .A2(n14668), .A3(n14667), .ZN(n14671) );
  AOI22_X1 U18170 ( .A1(n14770), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n9854), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n14670) );
  AOI22_X1 U18171 ( .A1(n10645), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n10644), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n14669) );
  NAND4_X1 U18172 ( .A1(n14672), .A2(n14671), .A3(n14670), .A4(n14669), .ZN(
        n14680) );
  AOI22_X1 U18173 ( .A1(n9855), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(n9847), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n14678) );
  AOI22_X1 U18174 ( .A1(n14770), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n10647), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n14677) );
  AOI22_X1 U18175 ( .A1(n9843), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(n9823), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n14676) );
  NAND2_X1 U18176 ( .A1(n9841), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(
        n14674) );
  NAND2_X1 U18177 ( .A1(n9857), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(
        n14673) );
  AND3_X1 U18178 ( .A1(n14674), .A2(n14673), .A3(n14773), .ZN(n14675) );
  NAND4_X1 U18179 ( .A1(n14678), .A2(n14677), .A3(n14676), .A4(n14675), .ZN(
        n14679) );
  AND2_X1 U18180 ( .A1(n14680), .A2(n14679), .ZN(n14683) );
  NAND2_X1 U18181 ( .A1(n14681), .A2(n14683), .ZN(n14687) );
  OAI211_X1 U18182 ( .C1(n14681), .C2(n14683), .A(n14723), .B(n14687), .ZN(
        n14685) );
  INV_X1 U18183 ( .A(n14685), .ZN(n14682) );
  INV_X1 U18184 ( .A(n14683), .ZN(n14684) );
  NOR2_X1 U18185 ( .A1(n20062), .A2(n14684), .ZN(n15651) );
  NAND2_X1 U18186 ( .A1(n15652), .A2(n15651), .ZN(n15650) );
  INV_X1 U18187 ( .A(n14687), .ZN(n14702) );
  AOI22_X1 U18188 ( .A1(n9855), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n10646), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n14693) );
  NAND2_X1 U18189 ( .A1(n13678), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n14689) );
  NAND2_X1 U18190 ( .A1(n9857), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n14688) );
  AND3_X1 U18191 ( .A1(n14747), .A2(n14689), .A3(n14688), .ZN(n14692) );
  AOI22_X1 U18192 ( .A1(n14770), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n9854), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n14691) );
  AOI22_X1 U18193 ( .A1(n10645), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n9823), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n14690) );
  NAND4_X1 U18194 ( .A1(n14693), .A2(n14692), .A3(n14691), .A4(n14690), .ZN(
        n14701) );
  AOI22_X1 U18195 ( .A1(n9855), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(n9847), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n14699) );
  AOI22_X1 U18196 ( .A1(n14770), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n10647), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n14698) );
  AOI22_X1 U18197 ( .A1(n9843), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(n9823), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n14697) );
  NAND2_X1 U18198 ( .A1(n13678), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(
        n14695) );
  NAND2_X1 U18199 ( .A1(n9859), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n14694) );
  AND3_X1 U18200 ( .A1(n14695), .A2(n14694), .A3(n14773), .ZN(n14696) );
  NAND4_X1 U18201 ( .A1(n14699), .A2(n14698), .A3(n14697), .A4(n14696), .ZN(
        n14700) );
  AND2_X1 U18202 ( .A1(n14701), .A2(n14700), .ZN(n14704) );
  NAND2_X1 U18203 ( .A1(n14702), .A2(n14704), .ZN(n14722) );
  OAI211_X1 U18204 ( .C1(n14702), .C2(n14704), .A(n14723), .B(n14722), .ZN(
        n14705) );
  NAND2_X1 U18205 ( .A1(n9839), .A2(n14704), .ZN(n15646) );
  NOR2_X2 U18206 ( .A1(n15647), .A2(n15646), .ZN(n15645) );
  AOI22_X1 U18207 ( .A1(n9855), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(n9847), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n14713) );
  AOI22_X1 U18208 ( .A1(n14770), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n9854), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n14712) );
  AOI22_X1 U18209 ( .A1(n10645), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n9822), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n14711) );
  NAND2_X1 U18210 ( .A1(n13678), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n14709) );
  NAND2_X1 U18211 ( .A1(n9859), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n14708) );
  AND3_X1 U18212 ( .A1(n14709), .A2(n14708), .A3(n14773), .ZN(n14710) );
  NAND4_X1 U18213 ( .A1(n14713), .A2(n14712), .A3(n14711), .A4(n14710), .ZN(
        n14721) );
  AOI22_X1 U18214 ( .A1(n9855), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n9847), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n14719) );
  NAND2_X1 U18215 ( .A1(n9841), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n14715) );
  NAND2_X1 U18216 ( .A1(n9858), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n14714) );
  AND3_X1 U18217 ( .A1(n14747), .A2(n14715), .A3(n14714), .ZN(n14718) );
  AOI22_X1 U18218 ( .A1(n14770), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n10647), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n14717) );
  AOI22_X1 U18219 ( .A1(n9843), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n9823), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n14716) );
  NAND4_X1 U18220 ( .A1(n14719), .A2(n14718), .A3(n14717), .A4(n14716), .ZN(
        n14720) );
  NAND2_X1 U18221 ( .A1(n14721), .A2(n14720), .ZN(n14729) );
  INV_X1 U18222 ( .A(n14729), .ZN(n14725) );
  INV_X1 U18223 ( .A(n14722), .ZN(n14724) );
  OR2_X1 U18224 ( .A1(n14722), .A2(n14729), .ZN(n15631) );
  OAI211_X1 U18225 ( .C1(n14725), .C2(n14724), .A(n14723), .B(n15631), .ZN(
        n14726) );
  NOR2_X1 U18226 ( .A1(n20062), .A2(n14729), .ZN(n15639) );
  NAND2_X1 U18227 ( .A1(n15637), .A2(n15639), .ZN(n15638) );
  INV_X1 U18228 ( .A(n14730), .ZN(n15632) );
  AOI22_X1 U18229 ( .A1(n9855), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(n9847), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n14736) );
  AOI22_X1 U18230 ( .A1(n14770), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n9854), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n14735) );
  AOI22_X1 U18231 ( .A1(n9843), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(n9823), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n14734) );
  NAND2_X1 U18232 ( .A1(n13678), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n14732) );
  NAND2_X1 U18233 ( .A1(n9858), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n14731) );
  AND3_X1 U18234 ( .A1(n14732), .A2(n14731), .A3(n14773), .ZN(n14733) );
  NAND4_X1 U18235 ( .A1(n14736), .A2(n14735), .A3(n14734), .A4(n14733), .ZN(
        n14744) );
  AOI22_X1 U18236 ( .A1(n9855), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n10646), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n14742) );
  NAND2_X1 U18237 ( .A1(n9841), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n14738) );
  NAND2_X1 U18238 ( .A1(n9857), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n14737) );
  AND3_X1 U18239 ( .A1(n14747), .A2(n14738), .A3(n14737), .ZN(n14741) );
  AOI22_X1 U18240 ( .A1(n14770), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10647), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n14740) );
  AOI22_X1 U18241 ( .A1(n10645), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n10644), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n14739) );
  NAND4_X1 U18242 ( .A1(n14742), .A2(n14741), .A3(n14740), .A4(n14739), .ZN(
        n14743) );
  NAND2_X1 U18243 ( .A1(n14744), .A2(n14743), .ZN(n15633) );
  AOI21_X2 U18244 ( .B1(n15638), .B2(n15632), .A(n15633), .ZN(n15626) );
  AOI22_X1 U18245 ( .A1(n9847), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n14770), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n14751) );
  NAND2_X1 U18246 ( .A1(n10644), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n14746) );
  NAND2_X1 U18247 ( .A1(n9857), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n14745) );
  AND3_X1 U18248 ( .A1(n14747), .A2(n14746), .A3(n14745), .ZN(n14750) );
  AOI22_X1 U18249 ( .A1(n9855), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n9854), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n14749) );
  AOI22_X1 U18250 ( .A1(n9843), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n13678), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n14748) );
  NAND4_X1 U18251 ( .A1(n14751), .A2(n14750), .A3(n14749), .A4(n14748), .ZN(
        n14759) );
  AOI22_X1 U18252 ( .A1(n10646), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n14770), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n14757) );
  AOI22_X1 U18253 ( .A1(n9855), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n10647), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n14756) );
  AOI22_X1 U18254 ( .A1(n10645), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n9822), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n14755) );
  NAND2_X1 U18255 ( .A1(n9841), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(
        n14753) );
  NAND2_X1 U18256 ( .A1(n9859), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n14752) );
  AND3_X1 U18257 ( .A1(n14753), .A2(n14752), .A3(n14773), .ZN(n14754) );
  NAND4_X1 U18258 ( .A1(n14757), .A2(n14756), .A3(n14755), .A4(n14754), .ZN(
        n14758) );
  NAND2_X1 U18259 ( .A1(n14759), .A2(n14758), .ZN(n14763) );
  INV_X1 U18260 ( .A(n15633), .ZN(n14760) );
  NAND2_X1 U18261 ( .A1(n20062), .A2(n14760), .ZN(n14761) );
  OR2_X1 U18262 ( .A1(n15631), .A2(n14761), .ZN(n14762) );
  NOR2_X1 U18263 ( .A1(n14762), .A2(n14763), .ZN(n14764) );
  AOI21_X1 U18264 ( .B1(n14763), .B2(n14762), .A(n14764), .ZN(n15625) );
  NAND2_X1 U18265 ( .A1(n15626), .A2(n15625), .ZN(n15627) );
  INV_X1 U18266 ( .A(n14764), .ZN(n14765) );
  NAND2_X1 U18267 ( .A1(n15627), .A2(n14765), .ZN(n14783) );
  AOI22_X1 U18268 ( .A1(n9855), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n10646), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n14767) );
  AOI22_X1 U18269 ( .A1(n14770), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n9854), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n14766) );
  NAND2_X1 U18270 ( .A1(n14767), .A2(n14766), .ZN(n14780) );
  AOI21_X1 U18271 ( .B1(n9858), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A(
        n14773), .ZN(n14769) );
  AOI22_X1 U18272 ( .A1(n13678), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n9822), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n14768) );
  OAI211_X1 U18273 ( .C1(n14626), .C2(n19713), .A(n14769), .B(n14768), .ZN(
        n14779) );
  AOI22_X1 U18274 ( .A1(n9847), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n14770), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n14772) );
  AOI22_X1 U18275 ( .A1(n9855), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n10647), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n14771) );
  NAND2_X1 U18276 ( .A1(n14772), .A2(n14771), .ZN(n14778) );
  AOI22_X1 U18277 ( .A1(n10645), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n13678), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n14776) );
  NAND2_X1 U18278 ( .A1(n9859), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n14775) );
  NAND2_X1 U18279 ( .A1(n9823), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n14774) );
  NAND4_X1 U18280 ( .A1(n14776), .A2(n14775), .A3(n14774), .A4(n14773), .ZN(
        n14777) );
  OAI22_X1 U18281 ( .A1(n14780), .A2(n14779), .B1(n14778), .B2(n14777), .ZN(
        n14781) );
  INV_X1 U18282 ( .A(n14781), .ZN(n14782) );
  XNOR2_X1 U18283 ( .A(n14783), .B(n14782), .ZN(n14792) );
  AOI22_X1 U18284 ( .A1(n19223), .A2(BUF2_REG_30__SCAN_IN), .B1(n19222), .B2(
        BUF1_REG_30__SCAN_IN), .ZN(n14785) );
  AOI22_X1 U18285 ( .A1(n19221), .A2(n19232), .B1(n19257), .B2(
        P2_EAX_REG_30__SCAN_IN), .ZN(n14784) );
  OAI211_X1 U18286 ( .C1(n14786), .C2(n19229), .A(n14785), .B(n14784), .ZN(
        n14787) );
  INV_X1 U18287 ( .A(n14787), .ZN(n14788) );
  OAI21_X1 U18288 ( .B1(n14792), .B2(n19258), .A(n14788), .ZN(P2_U2889) );
  NOR2_X1 U18289 ( .A1(n14789), .A2(n15661), .ZN(n14790) );
  AOI21_X1 U18290 ( .B1(P2_EBX_REG_30__SCAN_IN), .B2(n15661), .A(n14790), .ZN(
        n14791) );
  OAI21_X1 U18291 ( .B1(n14792), .B2(n15694), .A(n14791), .ZN(P2_U2857) );
  OAI21_X1 U18292 ( .B1(n14795), .B2(n14794), .A(n14793), .ZN(n19326) );
  OAI22_X1 U18293 ( .A1(n19319), .A2(n19326), .B1(n19936), .B2(n19345), .ZN(
        n14798) );
  NOR2_X1 U18294 ( .A1(n19325), .A2(n14796), .ZN(n14797) );
  AOI211_X1 U18295 ( .C1(n19313), .C2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A(
        n14798), .B(n14797), .ZN(n14804) );
  INV_X1 U18296 ( .A(n14799), .ZN(n14800) );
  AOI21_X1 U18297 ( .B1(n14802), .B2(n14801), .A(n14800), .ZN(n19330) );
  NAND2_X1 U18298 ( .A1(n19330), .A2(n12840), .ZN(n14803) );
  OAI211_X1 U18299 ( .C1(n16545), .C2(n14805), .A(n14804), .B(n14803), .ZN(
        P2_U3012) );
  INV_X1 U18300 ( .A(n15126), .ZN(n14991) );
  OAI22_X1 U18301 ( .A1(n14819), .A2(n12848), .B1(n14806), .B2(n9867), .ZN(
        n14809) );
  XNOR2_X1 U18302 ( .A(n14809), .B(n14808), .ZN(n15310) );
  INV_X1 U18303 ( .A(n15122), .ZN(n14814) );
  AOI22_X1 U18304 ( .A1(n20147), .A2(P1_EBX_REG_30__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n20140), .ZN(n14813) );
  INV_X1 U18305 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n20974) );
  NOR2_X1 U18306 ( .A1(n14823), .A2(n20974), .ZN(n14811) );
  OAI21_X1 U18307 ( .B1(P1_REIP_REG_30__SCAN_IN), .B2(n14811), .A(n14810), 
        .ZN(n14812) );
  OAI211_X1 U18308 ( .C1(n20143), .C2(n14814), .A(n14813), .B(n14812), .ZN(
        n14815) );
  AOI21_X1 U18309 ( .B1(n15310), .B2(n20149), .A(n14815), .ZN(n14816) );
  OAI21_X1 U18310 ( .B1(n14991), .B2(n14988), .A(n14816), .ZN(P1_U2810) );
  AND2_X1 U18311 ( .A1(n9867), .A2(n14817), .ZN(n14818) );
  NAND2_X1 U18312 ( .A1(n15134), .A2(n20131), .ZN(n14832) );
  INV_X1 U18313 ( .A(n15132), .ZN(n14830) );
  INV_X1 U18314 ( .A(n14823), .ZN(n14826) );
  OAI22_X1 U18315 ( .A1(n20122), .A2(n14992), .B1(n14824), .B2(n20158), .ZN(
        n14825) );
  AOI21_X1 U18316 ( .B1(n14826), .B2(n20974), .A(n14825), .ZN(n14827) );
  OAI21_X1 U18317 ( .B1(n14828), .B2(n20974), .A(n14827), .ZN(n14829) );
  AOI21_X1 U18318 ( .B1(n20154), .B2(n14830), .A(n14829), .ZN(n14831) );
  OAI211_X1 U18319 ( .C1(n20124), .C2(n15322), .A(n14832), .B(n14831), .ZN(
        P1_U2811) );
  AOI21_X1 U18320 ( .B1(n14834), .B2(n14833), .A(n12408), .ZN(n15142) );
  INV_X1 U18321 ( .A(n15142), .ZN(n15058) );
  INV_X1 U18322 ( .A(n14846), .ZN(n14836) );
  AOI21_X1 U18323 ( .B1(n14837), .B2(n14836), .A(n14835), .ZN(n15338) );
  AOI22_X1 U18324 ( .A1(n20147), .A2(P1_EBX_REG_27__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n20140), .ZN(n14842) );
  INV_X1 U18325 ( .A(n14838), .ZN(n14839) );
  OAI21_X1 U18326 ( .B1(P1_REIP_REG_27__SCAN_IN), .B2(n14840), .A(n14839), 
        .ZN(n14841) );
  OAI211_X1 U18327 ( .C1(n20143), .C2(n15140), .A(n14842), .B(n14841), .ZN(
        n14843) );
  AOI21_X1 U18328 ( .B1(n15338), .B2(n20149), .A(n14843), .ZN(n14844) );
  OAI21_X1 U18329 ( .B1(n15058), .B2(n14988), .A(n14844), .ZN(P1_U2813) );
  AND2_X1 U18330 ( .A1(n14861), .A2(n14845), .ZN(n14847) );
  OR2_X1 U18331 ( .A1(n14847), .A2(n14846), .ZN(n15346) );
  INV_X1 U18332 ( .A(P1_REIP_REG_26__SCAN_IN), .ZN(n20968) );
  OAI21_X1 U18333 ( .B1(n20151), .B2(n14848), .A(n20968), .ZN(n14850) );
  INV_X1 U18334 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n15148) );
  OAI22_X1 U18335 ( .A1(n20122), .A2(n14994), .B1(n15148), .B2(n20158), .ZN(
        n14849) );
  AOI21_X1 U18336 ( .B1(n14851), .B2(n14850), .A(n14849), .ZN(n14852) );
  OAI21_X1 U18337 ( .B1(n15346), .B2(n20124), .A(n14852), .ZN(n14856) );
  OAI21_X1 U18338 ( .B1(n14853), .B2(n14854), .A(n14833), .ZN(n15149) );
  NOR2_X1 U18339 ( .A1(n15149), .A2(n14988), .ZN(n14855) );
  AOI211_X1 U18340 ( .C1(n20154), .C2(n15152), .A(n14856), .B(n14855), .ZN(
        n14857) );
  INV_X1 U18341 ( .A(n14857), .ZN(P1_U2814) );
  AOI21_X1 U18342 ( .B1(n14860), .B2(n14859), .A(n14853), .ZN(n15162) );
  INV_X1 U18343 ( .A(n15162), .ZN(n14996) );
  AOI21_X1 U18344 ( .B1(n14862), .B2(n14878), .A(n12922), .ZN(n15358) );
  NOR2_X1 U18345 ( .A1(n20143), .A2(n15160), .ZN(n14871) );
  INV_X1 U18346 ( .A(n14880), .ZN(n14863) );
  AND2_X1 U18347 ( .A1(n20117), .A2(n14863), .ZN(n14864) );
  OR2_X1 U18348 ( .A1(n14958), .A2(n14864), .ZN(n14879) );
  INV_X1 U18349 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n14869) );
  AOI22_X1 U18350 ( .A1(n20147), .A2(P1_EBX_REG_25__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n20140), .ZN(n14868) );
  NAND2_X1 U18351 ( .A1(P1_REIP_REG_25__SCAN_IN), .A2(P1_REIP_REG_24__SCAN_IN), 
        .ZN(n14865) );
  OAI211_X1 U18352 ( .C1(P1_REIP_REG_25__SCAN_IN), .C2(n14866), .A(n20137), 
        .B(n14865), .ZN(n14867) );
  OAI211_X1 U18353 ( .C1(n14879), .C2(n14869), .A(n14868), .B(n14867), .ZN(
        n14870) );
  AOI211_X1 U18354 ( .C1(n15358), .C2(n20149), .A(n14871), .B(n14870), .ZN(
        n14872) );
  OAI21_X1 U18355 ( .B1(n14996), .B2(n14988), .A(n14872), .ZN(P1_U2815) );
  OR2_X1 U18356 ( .A1(n14873), .A2(n14888), .ZN(n14886) );
  INV_X1 U18357 ( .A(n14859), .ZN(n14874) );
  AOI21_X1 U18358 ( .B1(n14875), .B2(n14886), .A(n14874), .ZN(n15170) );
  INV_X1 U18359 ( .A(n15170), .ZN(n15069) );
  OR2_X1 U18360 ( .A1(n14892), .A2(n14876), .ZN(n14877) );
  AND2_X1 U18361 ( .A1(n14878), .A2(n14877), .ZN(n15365) );
  INV_X1 U18362 ( .A(n15365), .ZN(n14997) );
  INV_X1 U18363 ( .A(n14879), .ZN(n14897) );
  INV_X1 U18364 ( .A(P1_EBX_REG_24__SCAN_IN), .ZN(n14998) );
  OAI22_X1 U18365 ( .A1(n20122), .A2(n14998), .B1(n15167), .B2(n20158), .ZN(
        n14882) );
  NOR3_X1 U18366 ( .A1(n20151), .A2(P1_REIP_REG_24__SCAN_IN), .A3(n14880), 
        .ZN(n14881) );
  AOI211_X1 U18367 ( .C1(n14897), .C2(P1_REIP_REG_24__SCAN_IN), .A(n14882), 
        .B(n14881), .ZN(n14883) );
  OAI21_X1 U18368 ( .B1(n14997), .B2(n20124), .A(n14883), .ZN(n14884) );
  AOI21_X1 U18369 ( .B1(n15169), .B2(n20154), .A(n14884), .ZN(n14885) );
  OAI21_X1 U18370 ( .B1(n15069), .B2(n14988), .A(n14885), .ZN(P1_U2816) );
  INV_X1 U18371 ( .A(n14886), .ZN(n14887) );
  AOI21_X1 U18372 ( .B1(n14888), .B2(n14873), .A(n14887), .ZN(n15178) );
  NAND2_X1 U18373 ( .A1(n15178), .A2(n20131), .ZN(n14899) );
  NAND3_X1 U18374 ( .A1(n20137), .A2(P1_REIP_REG_21__SCAN_IN), .A3(n14906), 
        .ZN(n14907) );
  INV_X1 U18375 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n20962) );
  INV_X1 U18376 ( .A(P1_REIP_REG_23__SCAN_IN), .ZN(n14889) );
  OAI21_X1 U18377 ( .B1(n14907), .B2(n20962), .A(n14889), .ZN(n14896) );
  INV_X1 U18378 ( .A(P1_EBX_REG_23__SCAN_IN), .ZN(n14999) );
  OAI22_X1 U18379 ( .A1(n20122), .A2(n14999), .B1(n14890), .B2(n20158), .ZN(
        n14895) );
  AND2_X1 U18380 ( .A1(n14903), .A2(n14891), .ZN(n14893) );
  OR2_X1 U18381 ( .A1(n14893), .A2(n14892), .ZN(n15375) );
  NOR2_X1 U18382 ( .A1(n15375), .A2(n20124), .ZN(n14894) );
  AOI211_X1 U18383 ( .C1(n14897), .C2(n14896), .A(n14895), .B(n14894), .ZN(
        n14898) );
  OAI211_X1 U18384 ( .C1(n20143), .C2(n15176), .A(n14899), .B(n14898), .ZN(
        P1_U2817) );
  OR2_X1 U18385 ( .A1(n14900), .A2(n14901), .ZN(n14902) );
  NAND2_X1 U18386 ( .A1(n14873), .A2(n14902), .ZN(n15186) );
  INV_X1 U18387 ( .A(n14903), .ZN(n14904) );
  AOI21_X1 U18388 ( .B1(n14905), .B2(n14919), .A(n14904), .ZN(n15394) );
  INV_X1 U18389 ( .A(n15394), .ZN(n15000) );
  INV_X1 U18390 ( .A(n14906), .ZN(n14921) );
  AOI21_X1 U18391 ( .B1(n20137), .B2(n14921), .A(n20135), .ZN(n14920) );
  OAI21_X1 U18392 ( .B1(P1_REIP_REG_21__SCAN_IN), .B2(n20151), .A(n14920), 
        .ZN(n14910) );
  OAI22_X1 U18393 ( .A1(n20122), .A2(n15001), .B1(n15185), .B2(n20158), .ZN(
        n14909) );
  NOR2_X1 U18394 ( .A1(n14907), .A2(P1_REIP_REG_22__SCAN_IN), .ZN(n14908) );
  AOI211_X1 U18395 ( .C1(P1_REIP_REG_22__SCAN_IN), .C2(n14910), .A(n14909), 
        .B(n14908), .ZN(n14911) );
  OAI21_X1 U18396 ( .B1(n15000), .B2(n20124), .A(n14911), .ZN(n14912) );
  AOI21_X1 U18397 ( .B1(n15189), .B2(n20154), .A(n14912), .ZN(n14913) );
  OAI21_X1 U18398 ( .B1(n15186), .B2(n14988), .A(n14913), .ZN(P1_U2818) );
  INV_X1 U18399 ( .A(n14914), .ZN(n14916) );
  INV_X1 U18400 ( .A(n14915), .ZN(n14930) );
  AOI21_X1 U18401 ( .B1(n14916), .B2(n14930), .A(n14900), .ZN(n15197) );
  INV_X1 U18402 ( .A(n15197), .ZN(n15085) );
  INV_X1 U18403 ( .A(n15195), .ZN(n14926) );
  NAND2_X1 U18404 ( .A1(n14933), .A2(n14917), .ZN(n14918) );
  NAND2_X1 U18405 ( .A1(n14919), .A2(n14918), .ZN(n15399) );
  INV_X1 U18406 ( .A(n14920), .ZN(n14936) );
  INV_X1 U18407 ( .A(P1_EBX_REG_21__SCAN_IN), .ZN(n15002) );
  OAI22_X1 U18408 ( .A1(n20122), .A2(n15002), .B1(n21259), .B2(n20158), .ZN(
        n14923) );
  NOR3_X1 U18409 ( .A1(n20151), .A2(P1_REIP_REG_21__SCAN_IN), .A3(n14921), 
        .ZN(n14922) );
  AOI211_X1 U18410 ( .C1(n14936), .C2(P1_REIP_REG_21__SCAN_IN), .A(n14923), 
        .B(n14922), .ZN(n14924) );
  OAI21_X1 U18411 ( .B1(n15399), .B2(n20124), .A(n14924), .ZN(n14925) );
  AOI21_X1 U18412 ( .B1(n20154), .B2(n14926), .A(n14925), .ZN(n14927) );
  OAI21_X1 U18413 ( .B1(n15085), .B2(n14988), .A(n14927), .ZN(P1_U2819) );
  INV_X1 U18414 ( .A(n14928), .ZN(n14932) );
  INV_X1 U18415 ( .A(n14929), .ZN(n14931) );
  OAI21_X1 U18416 ( .B1(n15009), .B2(n14934), .A(n14933), .ZN(n15416) );
  AOI22_X1 U18417 ( .A1(n20147), .A2(P1_EBX_REG_20__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n20140), .ZN(n14939) );
  NOR2_X1 U18418 ( .A1(n20151), .A2(n14935), .ZN(n16264) );
  AND4_X1 U18419 ( .A1(n16237), .A2(P1_REIP_REG_19__SCAN_IN), .A3(
        P1_REIP_REG_18__SCAN_IN), .A4(n16238), .ZN(n14937) );
  OAI21_X1 U18420 ( .B1(n14937), .B2(P1_REIP_REG_20__SCAN_IN), .A(n14936), 
        .ZN(n14938) );
  OAI211_X1 U18421 ( .C1(n15416), .C2(n20124), .A(n14939), .B(n14938), .ZN(
        n14940) );
  AOI21_X1 U18422 ( .B1(n20154), .B2(n15204), .A(n14940), .ZN(n14941) );
  OAI21_X1 U18423 ( .B1(n15207), .B2(n14988), .A(n14941), .ZN(P1_U2820) );
  INV_X1 U18424 ( .A(n14942), .ZN(n14946) );
  INV_X1 U18425 ( .A(n14943), .ZN(n14945) );
  AOI21_X1 U18426 ( .B1(n14946), .B2(n14945), .A(n14944), .ZN(n16307) );
  INV_X1 U18427 ( .A(n16307), .ZN(n15100) );
  INV_X1 U18428 ( .A(n14966), .ZN(n15021) );
  OAI21_X1 U18429 ( .B1(n15021), .B2(n14965), .A(n14947), .ZN(n14948) );
  NAND2_X1 U18430 ( .A1(n14948), .A2(n9927), .ZN(n16346) );
  NOR2_X1 U18431 ( .A1(n16346), .A2(n20124), .ZN(n14953) );
  INV_X1 U18432 ( .A(P1_EBX_REG_17__SCAN_IN), .ZN(n14949) );
  OR2_X1 U18433 ( .A1(n20122), .A2(n14949), .ZN(n14950) );
  OAI211_X1 U18434 ( .C1(n14951), .C2(n20158), .A(n14950), .B(n20256), .ZN(
        n14952) );
  AOI211_X1 U18435 ( .C1(n20154), .C2(n16306), .A(n14953), .B(n14952), .ZN(
        n14961) );
  AOI21_X1 U18436 ( .B1(n14955), .B2(n14954), .A(n14958), .ZN(n16280) );
  NOR2_X1 U18437 ( .A1(n14958), .A2(n14956), .ZN(n14957) );
  INV_X1 U18438 ( .A(n16260), .ZN(n16273) );
  OAI21_X1 U18439 ( .B1(n14958), .B2(n16238), .A(n16273), .ZN(n16251) );
  INV_X1 U18440 ( .A(n16237), .ZN(n16263) );
  OAI21_X1 U18441 ( .B1(n14967), .B2(n16263), .A(n20952), .ZN(n14959) );
  NAND2_X1 U18442 ( .A1(n16251), .A2(n14959), .ZN(n14960) );
  OAI211_X1 U18443 ( .C1(n15100), .C2(n14988), .A(n14961), .B(n14960), .ZN(
        P1_U2823) );
  INV_X1 U18444 ( .A(n14962), .ZN(n15025) );
  AOI21_X1 U18445 ( .B1(n14963), .B2(n15025), .A(n14943), .ZN(n14964) );
  INV_X1 U18446 ( .A(n14964), .ZN(n15233) );
  INV_X1 U18447 ( .A(n15230), .ZN(n14973) );
  XNOR2_X1 U18448 ( .A(n14966), .B(n14965), .ZN(n16356) );
  OAI211_X1 U18449 ( .C1(P1_REIP_REG_16__SCAN_IN), .C2(P1_REIP_REG_15__SCAN_IN), .A(n16237), .B(n14967), .ZN(n14969) );
  AOI21_X1 U18450 ( .B1(n20140), .B2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n20280), .ZN(n14968) );
  OAI211_X1 U18451 ( .C1(n14970), .C2(n20122), .A(n14969), .B(n14968), .ZN(
        n14971) );
  AOI21_X1 U18452 ( .B1(n16356), .B2(n20149), .A(n14971), .ZN(n14972) );
  OAI21_X1 U18453 ( .B1(n20143), .B2(n14973), .A(n14972), .ZN(n14974) );
  AOI21_X1 U18454 ( .B1(n16260), .B2(P1_REIP_REG_16__SCAN_IN), .A(n14974), 
        .ZN(n14975) );
  OAI21_X1 U18455 ( .B1(n15233), .B2(n14988), .A(n14975), .ZN(P1_U2824) );
  NAND2_X1 U18456 ( .A1(n14457), .A2(n14977), .ZN(n14978) );
  NAND2_X1 U18457 ( .A1(n14976), .A2(n14978), .ZN(n15046) );
  OAI21_X1 U18458 ( .B1(n15046), .B2(n15047), .A(n14976), .ZN(n15036) );
  NAND2_X1 U18459 ( .A1(n15036), .A2(n15035), .ZN(n15034) );
  INV_X1 U18460 ( .A(n14979), .ZN(n14981) );
  AOI21_X1 U18461 ( .B1(n15034), .B2(n14981), .A(n14980), .ZN(n15253) );
  INV_X1 U18462 ( .A(n15253), .ZN(n15113) );
  INV_X1 U18463 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n20947) );
  AOI21_X1 U18464 ( .B1(n20154), .B2(n15249), .A(n20280), .ZN(n14982) );
  OAI21_X1 U18465 ( .B1(n14983), .B2(n20158), .A(n14982), .ZN(n14984) );
  AOI221_X1 U18466 ( .B1(n16280), .B2(P1_REIP_REG_13__SCAN_IN), .C1(n16264), 
        .C2(n20947), .A(n14984), .ZN(n14987) );
  AOI21_X1 U18467 ( .B1(n14985), .B2(n15039), .A(n15030), .ZN(n15443) );
  AOI22_X1 U18468 ( .A1(n15443), .A2(n20149), .B1(n20147), .B2(
        P1_EBX_REG_13__SCAN_IN), .ZN(n14986) );
  OAI211_X1 U18469 ( .C1(n15113), .C2(n14988), .A(n14987), .B(n14986), .ZN(
        P1_U2827) );
  OAI22_X1 U18470 ( .A1(n15274), .A2(n20175), .B1(n20182), .B2(n14989), .ZN(
        P1_U2841) );
  AOI22_X1 U18471 ( .A1(n15310), .A2(n20171), .B1(P1_EBX_REG_30__SCAN_IN), 
        .B2(n15032), .ZN(n14990) );
  OAI21_X1 U18472 ( .B1(n14991), .B2(n9828), .A(n14990), .ZN(P1_U2842) );
  INV_X1 U18473 ( .A(n15134), .ZN(n15054) );
  OAI222_X1 U18474 ( .A1(n9828), .A2(n15054), .B1(n14992), .B2(n20182), .C1(
        n15322), .C2(n20175), .ZN(P1_U2843) );
  AOI22_X1 U18475 ( .A1(n15338), .A2(n20171), .B1(P1_EBX_REG_27__SCAN_IN), 
        .B2(n15032), .ZN(n14993) );
  OAI21_X1 U18476 ( .B1(n15058), .B2(n9828), .A(n14993), .ZN(P1_U2845) );
  OAI222_X1 U18477 ( .A1(n9828), .A2(n15149), .B1(n14994), .B2(n20182), .C1(
        n15346), .C2(n20175), .ZN(P1_U2846) );
  AOI22_X1 U18478 ( .A1(n15358), .A2(n20171), .B1(P1_EBX_REG_25__SCAN_IN), 
        .B2(n15032), .ZN(n14995) );
  OAI21_X1 U18479 ( .B1(n14996), .B2(n9828), .A(n14995), .ZN(P1_U2847) );
  OAI222_X1 U18480 ( .A1(n9828), .A2(n15069), .B1(n14998), .B2(n20182), .C1(
        n14997), .C2(n20175), .ZN(P1_U2848) );
  INV_X1 U18481 ( .A(n15178), .ZN(n15075) );
  OAI222_X1 U18482 ( .A1(n9828), .A2(n15075), .B1(n14999), .B2(n20182), .C1(
        n15375), .C2(n20175), .ZN(P1_U2849) );
  OAI222_X1 U18483 ( .A1(n9828), .A2(n15186), .B1(n15001), .B2(n20182), .C1(
        n15000), .C2(n20175), .ZN(P1_U2850) );
  OAI222_X1 U18484 ( .A1(n9828), .A2(n15085), .B1(n15002), .B2(n20182), .C1(
        n15399), .C2(n20175), .ZN(P1_U2851) );
  INV_X1 U18485 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n15003) );
  OAI222_X1 U18486 ( .A1(n9828), .A2(n15207), .B1(n20182), .B2(n15003), .C1(
        n15416), .C2(n20175), .ZN(P1_U2852) );
  NAND2_X1 U18487 ( .A1(n15004), .A2(n15005), .ZN(n15006) );
  INV_X1 U18488 ( .A(n16296), .ZN(n15011) );
  INV_X1 U18489 ( .A(P1_EBX_REG_19__SCAN_IN), .ZN(n15010) );
  AND2_X1 U18490 ( .A1(n9887), .A2(n15007), .ZN(n15008) );
  OR2_X1 U18491 ( .A1(n15009), .A2(n15008), .ZN(n16246) );
  OAI222_X1 U18492 ( .A1(n9828), .A2(n15011), .B1(n15010), .B2(n20182), .C1(
        n16246), .C2(n20175), .ZN(P1_U2853) );
  XOR2_X1 U18493 ( .A(n15012), .B(n14944), .Z(n16252) );
  NAND2_X1 U18494 ( .A1(n9927), .A2(n15013), .ZN(n15014) );
  NAND2_X1 U18495 ( .A1(n9887), .A2(n15014), .ZN(n16255) );
  OAI22_X1 U18496 ( .A1(n16255), .A2(n20175), .B1(n15015), .B2(n20182), .ZN(
        n15016) );
  AOI21_X1 U18497 ( .B1(n16252), .B2(n20178), .A(n15016), .ZN(n15017) );
  INV_X1 U18498 ( .A(n15017), .ZN(P1_U2854) );
  OAI222_X1 U18499 ( .A1(n15100), .A2(n9828), .B1(n14949), .B2(n20182), .C1(
        n20175), .C2(n16346), .ZN(P1_U2855) );
  AOI22_X1 U18500 ( .A1(n16356), .A2(n20171), .B1(P1_EBX_REG_16__SCAN_IN), 
        .B2(n15032), .ZN(n15018) );
  OAI21_X1 U18501 ( .B1(n15233), .B2(n9828), .A(n15018), .ZN(P1_U2856) );
  INV_X1 U18502 ( .A(n15030), .ZN(n15020) );
  OAI21_X1 U18503 ( .B1(n15020), .B2(n15029), .A(n15019), .ZN(n15022) );
  NAND2_X1 U18504 ( .A1(n15022), .A2(n15021), .ZN(n16256) );
  INV_X1 U18505 ( .A(P1_EBX_REG_15__SCAN_IN), .ZN(n15027) );
  AOI21_X1 U18506 ( .B1(n15026), .B2(n15024), .A(n14962), .ZN(n16318) );
  INV_X1 U18507 ( .A(n16318), .ZN(n15109) );
  OAI222_X1 U18508 ( .A1(n16256), .A2(n20175), .B1(n15027), .B2(n20182), .C1(
        n15109), .C2(n9828), .ZN(P1_U2857) );
  OAI21_X1 U18509 ( .B1(n14980), .B2(n15028), .A(n15024), .ZN(n16265) );
  XNOR2_X1 U18510 ( .A(n15030), .B(n15029), .ZN(n16371) );
  AOI22_X1 U18511 ( .A1(n16371), .A2(n20171), .B1(P1_EBX_REG_14__SCAN_IN), 
        .B2(n15032), .ZN(n15031) );
  OAI21_X1 U18512 ( .B1(n16265), .B2(n9828), .A(n15031), .ZN(P1_U2858) );
  AOI22_X1 U18513 ( .A1(n15443), .A2(n20171), .B1(P1_EBX_REG_13__SCAN_IN), 
        .B2(n15032), .ZN(n15033) );
  OAI21_X1 U18514 ( .B1(n15113), .B2(n9828), .A(n15033), .ZN(P1_U2859) );
  OAI21_X1 U18515 ( .B1(n15036), .B2(n15035), .A(n15034), .ZN(n15258) );
  INV_X1 U18516 ( .A(P1_EBX_REG_12__SCAN_IN), .ZN(n16274) );
  NAND2_X1 U18517 ( .A1(n15044), .A2(n15037), .ZN(n15038) );
  NAND2_X1 U18518 ( .A1(n15039), .A2(n15038), .ZN(n16275) );
  OAI222_X1 U18519 ( .A1(n15258), .A2(n9828), .B1(n16274), .B2(n20182), .C1(
        n16275), .C2(n20175), .ZN(P1_U2860) );
  INV_X1 U18520 ( .A(n15040), .ZN(n15043) );
  OAI21_X1 U18521 ( .B1(n15043), .B2(n15042), .A(n15041), .ZN(n15045) );
  NAND2_X1 U18522 ( .A1(n15045), .A2(n15044), .ZN(n16286) );
  INV_X1 U18523 ( .A(P1_EBX_REG_11__SCAN_IN), .ZN(n15048) );
  XOR2_X1 U18524 ( .A(n15047), .B(n15046), .Z(n16324) );
  INV_X1 U18525 ( .A(n16324), .ZN(n15119) );
  OAI222_X1 U18526 ( .A1(n16286), .A2(n20175), .B1(n15048), .B2(n20182), .C1(
        n15119), .C2(n9828), .ZN(P1_U2861) );
  INV_X1 U18527 ( .A(DATAI_13_), .ZN(n15050) );
  MUX2_X1 U18528 ( .A(n15050), .B(n15049), .S(n20303), .Z(n20222) );
  OAI22_X1 U18529 ( .A1(n15091), .A2(n20222), .B1(n13648), .B2(n15090), .ZN(
        n15051) );
  AOI21_X1 U18530 ( .B1(n16295), .B2(DATAI_29_), .A(n15051), .ZN(n15053) );
  NAND2_X1 U18531 ( .A1(n15105), .A2(BUF1_REG_29__SCAN_IN), .ZN(n15052) );
  OAI211_X1 U18532 ( .C1(n15054), .C2(n15118), .A(n15053), .B(n15052), .ZN(
        P1_U2875) );
  OAI22_X1 U18533 ( .A1(n15091), .A2(n15117), .B1(n21309), .B2(n15090), .ZN(
        n15055) );
  AOI21_X1 U18534 ( .B1(n16295), .B2(DATAI_27_), .A(n15055), .ZN(n15057) );
  NAND2_X1 U18535 ( .A1(n15105), .A2(BUF1_REG_27__SCAN_IN), .ZN(n15056) );
  OAI211_X1 U18536 ( .C1(n15058), .C2(n15118), .A(n15057), .B(n15056), .ZN(
        P1_U2877) );
  OAI22_X1 U18537 ( .A1(n15091), .A2(n20216), .B1(n15059), .B2(n15090), .ZN(
        n15060) );
  AOI21_X1 U18538 ( .B1(n16295), .B2(DATAI_26_), .A(n15060), .ZN(n15062) );
  NAND2_X1 U18539 ( .A1(n15105), .A2(BUF1_REG_26__SCAN_IN), .ZN(n15061) );
  OAI211_X1 U18540 ( .C1(n15149), .C2(n15118), .A(n15062), .B(n15061), .ZN(
        P1_U2878) );
  NAND2_X1 U18541 ( .A1(n15162), .A2(n13019), .ZN(n15065) );
  OAI22_X1 U18542 ( .A1(n15091), .A2(n20213), .B1(n13646), .B2(n15090), .ZN(
        n15063) );
  AOI21_X1 U18543 ( .B1(n16295), .B2(DATAI_25_), .A(n15063), .ZN(n15064) );
  OAI211_X1 U18544 ( .C1(n16654), .C2(n16299), .A(n15065), .B(n15064), .ZN(
        P1_U2879) );
  OAI22_X1 U18545 ( .A1(n15091), .A2(n20210), .B1(n13641), .B2(n15090), .ZN(
        n15066) );
  AOI21_X1 U18546 ( .B1(n16295), .B2(DATAI_24_), .A(n15066), .ZN(n15068) );
  NAND2_X1 U18547 ( .A1(n15105), .A2(BUF1_REG_24__SCAN_IN), .ZN(n15067) );
  OAI211_X1 U18548 ( .C1(n15069), .C2(n15118), .A(n15068), .B(n15067), .ZN(
        P1_U2880) );
  OAI22_X1 U18549 ( .A1(n15091), .A2(n15071), .B1(n15070), .B2(n15090), .ZN(
        n15072) );
  AOI21_X1 U18550 ( .B1(n16295), .B2(DATAI_23_), .A(n15072), .ZN(n15074) );
  NAND2_X1 U18551 ( .A1(n15105), .A2(BUF1_REG_23__SCAN_IN), .ZN(n15073) );
  OAI211_X1 U18552 ( .C1(n15075), .C2(n15118), .A(n15074), .B(n15073), .ZN(
        P1_U2881) );
  OAI22_X1 U18553 ( .A1(n15091), .A2(n15076), .B1(n13901), .B2(n15090), .ZN(
        n15077) );
  AOI21_X1 U18554 ( .B1(n16295), .B2(DATAI_22_), .A(n15077), .ZN(n15079) );
  NAND2_X1 U18555 ( .A1(n15105), .A2(BUF1_REG_22__SCAN_IN), .ZN(n15078) );
  OAI211_X1 U18556 ( .C1(n15186), .C2(n15118), .A(n15079), .B(n15078), .ZN(
        P1_U2882) );
  OAI22_X1 U18557 ( .A1(n15091), .A2(n15081), .B1(n15080), .B2(n15090), .ZN(
        n15082) );
  AOI21_X1 U18558 ( .B1(n16295), .B2(DATAI_21_), .A(n15082), .ZN(n15084) );
  NAND2_X1 U18559 ( .A1(n15105), .A2(BUF1_REG_21__SCAN_IN), .ZN(n15083) );
  OAI211_X1 U18560 ( .C1(n15085), .C2(n15118), .A(n15084), .B(n15083), .ZN(
        P1_U2883) );
  INV_X1 U18561 ( .A(DATAI_20_), .ZN(n15087) );
  INV_X1 U18562 ( .A(n15091), .ZN(n16294) );
  AOI22_X1 U18563 ( .A1(n16294), .A2(n20335), .B1(P1_EAX_REG_20__SCAN_IN), 
        .B2(n16293), .ZN(n15086) );
  OAI21_X1 U18564 ( .B1(n15103), .B2(n15087), .A(n15086), .ZN(n15088) );
  AOI21_X1 U18565 ( .B1(n15105), .B2(BUF1_REG_20__SCAN_IN), .A(n15088), .ZN(
        n15089) );
  OAI21_X1 U18566 ( .B1(n15207), .B2(n15118), .A(n15089), .ZN(P1_U2884) );
  INV_X1 U18567 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n15095) );
  NAND2_X1 U18568 ( .A1(n16252), .A2(n13019), .ZN(n15094) );
  OAI22_X1 U18569 ( .A1(n15091), .A2(n20328), .B1(n13904), .B2(n15090), .ZN(
        n15092) );
  AOI21_X1 U18570 ( .B1(n16295), .B2(DATAI_18_), .A(n15092), .ZN(n15093) );
  OAI211_X1 U18571 ( .C1(n16299), .C2(n15095), .A(n15094), .B(n15093), .ZN(
        P1_U2886) );
  INV_X1 U18572 ( .A(DATAI_17_), .ZN(n15097) );
  AOI22_X1 U18573 ( .A1(n16294), .A2(n20325), .B1(P1_EAX_REG_17__SCAN_IN), 
        .B2(n16293), .ZN(n15096) );
  OAI21_X1 U18574 ( .B1(n15103), .B2(n15097), .A(n15096), .ZN(n15098) );
  AOI21_X1 U18575 ( .B1(n15105), .B2(BUF1_REG_17__SCAN_IN), .A(n15098), .ZN(
        n15099) );
  OAI21_X1 U18576 ( .B1(n15100), .B2(n15118), .A(n15099), .ZN(P1_U2887) );
  INV_X1 U18577 ( .A(DATAI_16_), .ZN(n15102) );
  AOI22_X1 U18578 ( .A1(n16294), .A2(n20316), .B1(P1_EAX_REG_16__SCAN_IN), 
        .B2(n16293), .ZN(n15101) );
  OAI21_X1 U18579 ( .B1(n15103), .B2(n15102), .A(n15101), .ZN(n15104) );
  AOI21_X1 U18580 ( .B1(n15105), .B2(BUF1_REG_16__SCAN_IN), .A(n15104), .ZN(
        n15106) );
  OAI21_X1 U18581 ( .B1(n15233), .B2(n15118), .A(n15106), .ZN(P1_U2888) );
  OAI222_X1 U18582 ( .A1(n15109), .A2(n15118), .B1(n15116), .B2(n15108), .C1(
        n15090), .C2(n15107), .ZN(P1_U2889) );
  INV_X1 U18583 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n15110) );
  OAI222_X1 U18584 ( .A1(n16265), .A2(n15118), .B1(n15111), .B2(n15116), .C1(
        n15110), .C2(n15090), .ZN(P1_U2890) );
  INV_X1 U18585 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n15112) );
  OAI222_X1 U18586 ( .A1(n15113), .A2(n15118), .B1(n20222), .B2(n15116), .C1(
        n15112), .C2(n15090), .ZN(P1_U2891) );
  OAI222_X1 U18587 ( .A1(n15258), .A2(n15118), .B1(n20219), .B2(n15116), .C1(
        n15114), .C2(n15090), .ZN(P1_U2892) );
  INV_X1 U18588 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n15115) );
  OAI222_X1 U18589 ( .A1(n15119), .A2(n15118), .B1(n15117), .B2(n15116), .C1(
        n15115), .C2(n15090), .ZN(P1_U2893) );
  NAND2_X1 U18590 ( .A1(n9836), .A2(n15120), .ZN(n15121) );
  XNOR2_X1 U18591 ( .A(n15121), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15312) );
  NAND2_X1 U18592 ( .A1(n15122), .A2(n16316), .ZN(n15123) );
  NAND2_X1 U18593 ( .A1(n20296), .A2(P1_REIP_REG_30__SCAN_IN), .ZN(n15304) );
  OAI211_X1 U18594 ( .C1(n15124), .C2(n15228), .A(n15123), .B(n15304), .ZN(
        n15125) );
  AOI21_X1 U18595 ( .B1(n15126), .B2(n16325), .A(n15125), .ZN(n15127) );
  OAI21_X1 U18596 ( .B1(n15312), .B2(n20088), .A(n15127), .ZN(P1_U2969) );
  MUX2_X1 U18597 ( .A(n9844), .B(n15129), .S(n15128), .Z(n15130) );
  XNOR2_X1 U18598 ( .A(n15130), .B(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15325) );
  NAND2_X1 U18599 ( .A1(n20280), .A2(P1_REIP_REG_29__SCAN_IN), .ZN(n15320) );
  NAND2_X1 U18600 ( .A1(n20242), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15131) );
  OAI211_X1 U18601 ( .C1(n15132), .C2(n20252), .A(n15320), .B(n15131), .ZN(
        n15133) );
  AOI21_X1 U18602 ( .B1(n15134), .B2(n16325), .A(n15133), .ZN(n15135) );
  OAI21_X1 U18603 ( .B1(n15325), .B2(n20088), .A(n15135), .ZN(P1_U2970) );
  NAND2_X1 U18604 ( .A1(n9909), .A2(n13001), .ZN(n15136) );
  MUX2_X1 U18605 ( .A(n15137), .B(n15136), .S(n9845), .Z(n15138) );
  XNOR2_X1 U18606 ( .A(n15138), .B(n15339), .ZN(n15343) );
  NOR2_X1 U18607 ( .A1(n20256), .A2(n20971), .ZN(n15337) );
  AOI21_X1 U18608 ( .B1(n20242), .B2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n15337), .ZN(n15139) );
  OAI21_X1 U18609 ( .B1(n15140), .B2(n20252), .A(n15139), .ZN(n15141) );
  AOI21_X1 U18610 ( .B1(n15142), .B2(n16325), .A(n15141), .ZN(n15143) );
  OAI21_X1 U18611 ( .B1(n20088), .B2(n15343), .A(n15143), .ZN(P1_U2972) );
  INV_X1 U18612 ( .A(n15174), .ZN(n15144) );
  OAI21_X1 U18613 ( .B1(n15144), .B2(n15344), .A(n9844), .ZN(n15145) );
  NAND2_X1 U18614 ( .A1(n15146), .A2(n15145), .ZN(n15147) );
  XNOR2_X1 U18615 ( .A(n15147), .B(n15348), .ZN(n15353) );
  NAND2_X1 U18616 ( .A1(n20296), .A2(P1_REIP_REG_26__SCAN_IN), .ZN(n15345) );
  OAI21_X1 U18617 ( .B1(n15228), .B2(n15148), .A(n15345), .ZN(n15151) );
  NOR2_X1 U18618 ( .A1(n15149), .A2(n20306), .ZN(n15150) );
  AOI211_X1 U18619 ( .C1(n16316), .C2(n15152), .A(n15151), .B(n15150), .ZN(
        n15153) );
  OAI21_X1 U18620 ( .B1(n20088), .B2(n15353), .A(n15153), .ZN(P1_U2973) );
  INV_X1 U18621 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15377) );
  NOR2_X1 U18622 ( .A1(n15154), .A2(n15377), .ZN(n15165) );
  INV_X1 U18623 ( .A(n15165), .ZN(n15157) );
  MUX2_X1 U18624 ( .A(n15155), .B(n15362), .S(n9845), .Z(n15156) );
  AOI21_X1 U18625 ( .B1(n15157), .B2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n15156), .ZN(n15158) );
  XNOR2_X1 U18626 ( .A(n15158), .B(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15361) );
  NAND2_X1 U18627 ( .A1(n20280), .A2(P1_REIP_REG_25__SCAN_IN), .ZN(n15354) );
  NAND2_X1 U18628 ( .A1(n20242), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15159) );
  OAI211_X1 U18629 ( .C1(n15160), .C2(n20252), .A(n15354), .B(n15159), .ZN(
        n15161) );
  AOI21_X1 U18630 ( .B1(n15162), .B2(n16325), .A(n15161), .ZN(n15163) );
  OAI21_X1 U18631 ( .B1(n20088), .B2(n15361), .A(n15163), .ZN(P1_U2974) );
  NOR2_X1 U18632 ( .A1(n15165), .A2(n15174), .ZN(n15164) );
  MUX2_X1 U18633 ( .A(n15165), .B(n15164), .S(n16302), .Z(n15166) );
  XNOR2_X1 U18634 ( .A(n15166), .B(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15371) );
  NOR2_X1 U18635 ( .A1(n20256), .A2(n20965), .ZN(n15364) );
  NOR2_X1 U18636 ( .A1(n15228), .A2(n15167), .ZN(n15168) );
  AOI211_X1 U18637 ( .C1(n15169), .C2(n16316), .A(n15364), .B(n15168), .ZN(
        n15172) );
  NAND2_X1 U18638 ( .A1(n15170), .A2(n16325), .ZN(n15171) );
  OAI211_X1 U18639 ( .C1(n15371), .C2(n20088), .A(n15172), .B(n15171), .ZN(
        P1_U2975) );
  XNOR2_X1 U18640 ( .A(n9844), .B(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15173) );
  XNOR2_X1 U18641 ( .A(n15174), .B(n15173), .ZN(n15380) );
  NAND2_X1 U18642 ( .A1(n20280), .A2(P1_REIP_REG_23__SCAN_IN), .ZN(n15374) );
  NAND2_X1 U18643 ( .A1(n20242), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15175) );
  OAI211_X1 U18644 ( .C1(n15176), .C2(n20252), .A(n15374), .B(n15175), .ZN(
        n15177) );
  AOI21_X1 U18645 ( .B1(n15178), .B2(n16325), .A(n15177), .ZN(n15179) );
  OAI21_X1 U18646 ( .B1(n15380), .B2(n20088), .A(n15179), .ZN(P1_U2976) );
  INV_X1 U18647 ( .A(n15181), .ZN(n15192) );
  NAND3_X1 U18648 ( .A1(n15192), .A2(n15287), .A3(
        P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n15183) );
  AOI21_X1 U18649 ( .B1(n15183), .B2(n9845), .A(n15182), .ZN(n15184) );
  XNOR2_X1 U18650 ( .A(n15184), .B(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15396) );
  NAND2_X1 U18651 ( .A1(n20296), .A2(P1_REIP_REG_22__SCAN_IN), .ZN(n15390) );
  OAI21_X1 U18652 ( .B1(n15228), .B2(n15185), .A(n15390), .ZN(n15188) );
  NOR2_X1 U18653 ( .A1(n15186), .A2(n20306), .ZN(n15187) );
  AOI211_X1 U18654 ( .C1(n16316), .C2(n15189), .A(n15188), .B(n15187), .ZN(
        n15190) );
  OAI21_X1 U18655 ( .B1(n20088), .B2(n15396), .A(n15190), .ZN(P1_U2977) );
  NAND4_X1 U18656 ( .A1(n15191), .A2(n16302), .A3(n15410), .A4(n15433), .ZN(
        n15199) );
  NAND3_X1 U18657 ( .A1(n15192), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        n9844), .ZN(n15200) );
  MUX2_X1 U18658 ( .A(n15199), .B(n15200), .S(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .Z(n15193) );
  XNOR2_X1 U18659 ( .A(n15193), .B(n15402), .ZN(n15405) );
  NAND2_X1 U18660 ( .A1(n20296), .A2(P1_REIP_REG_21__SCAN_IN), .ZN(n15397) );
  NAND2_X1 U18661 ( .A1(n20242), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15194) );
  OAI211_X1 U18662 ( .C1(n15195), .C2(n20252), .A(n15397), .B(n15194), .ZN(
        n15196) );
  AOI21_X1 U18663 ( .B1(n15197), .B2(n16325), .A(n15196), .ZN(n15198) );
  OAI21_X1 U18664 ( .B1(n15405), .B2(n20088), .A(n15198), .ZN(P1_U2978) );
  NAND2_X1 U18665 ( .A1(n15200), .A2(n15199), .ZN(n15201) );
  XNOR2_X1 U18666 ( .A(n15201), .B(n21220), .ZN(n15406) );
  NAND2_X1 U18667 ( .A1(n15406), .A2(n20248), .ZN(n15206) );
  INV_X1 U18668 ( .A(P1_REIP_REG_20__SCAN_IN), .ZN(n20959) );
  NOR2_X1 U18669 ( .A1(n20256), .A2(n20959), .ZN(n15412) );
  NOR2_X1 U18670 ( .A1(n15228), .A2(n15202), .ZN(n15203) );
  AOI211_X1 U18671 ( .C1(n15204), .C2(n16316), .A(n15412), .B(n15203), .ZN(
        n15205) );
  OAI211_X1 U18672 ( .C1(n20306), .C2(n15207), .A(n15206), .B(n15205), .ZN(
        P1_U2979) );
  OAI21_X1 U18673 ( .B1(n15433), .B2(n9844), .A(n15181), .ZN(n15209) );
  XNOR2_X1 U18674 ( .A(n9845), .B(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15208) );
  XNOR2_X1 U18675 ( .A(n15209), .B(n15208), .ZN(n15424) );
  AND2_X1 U18676 ( .A1(n20296), .A2(P1_REIP_REG_19__SCAN_IN), .ZN(n15417) );
  AOI21_X1 U18677 ( .B1(n20242), .B2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n15417), .ZN(n15210) );
  OAI21_X1 U18678 ( .B1(n16240), .B2(n20252), .A(n15210), .ZN(n15211) );
  AOI21_X1 U18679 ( .B1(n16296), .B2(n16325), .A(n15211), .ZN(n15212) );
  OAI21_X1 U18680 ( .B1(n15424), .B2(n20088), .A(n15212), .ZN(P1_U2980) );
  OAI21_X1 U18681 ( .B1(n15213), .B2(n15214), .A(n15181), .ZN(n15437) );
  INV_X1 U18682 ( .A(n16247), .ZN(n15216) );
  AOI22_X1 U18683 ( .A1(n20242), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B1(
        n20296), .B2(P1_REIP_REG_18__SCAN_IN), .ZN(n15215) );
  OAI21_X1 U18684 ( .B1(n15216), .B2(n20252), .A(n15215), .ZN(n15217) );
  AOI21_X1 U18685 ( .B1(n16252), .B2(n16325), .A(n15217), .ZN(n15218) );
  OAI21_X1 U18686 ( .B1(n20088), .B2(n15437), .A(n15218), .ZN(P1_U2981) );
  AOI21_X1 U18687 ( .B1(n15219), .B2(n15221), .A(n15220), .ZN(n15234) );
  INV_X1 U18688 ( .A(n15222), .ZN(n15223) );
  NAND2_X1 U18689 ( .A1(n15234), .A2(n15223), .ZN(n16313) );
  AOI21_X1 U18690 ( .B1(n16313), .B2(n15224), .A(n10047), .ZN(n15225) );
  XOR2_X1 U18691 ( .A(n15226), .B(n15225), .Z(n16358) );
  NAND2_X1 U18692 ( .A1(n16358), .A2(n20248), .ZN(n15232) );
  NAND2_X1 U18693 ( .A1(n20280), .A2(P1_REIP_REG_16__SCAN_IN), .ZN(n16354) );
  OAI21_X1 U18694 ( .B1(n15228), .B2(n15227), .A(n16354), .ZN(n15229) );
  AOI21_X1 U18695 ( .B1(n15230), .B2(n16316), .A(n15229), .ZN(n15231) );
  OAI211_X1 U18696 ( .C1(n20306), .C2(n15233), .A(n15232), .B(n15231), .ZN(
        P1_U2983) );
  INV_X1 U18697 ( .A(n15234), .ZN(n15236) );
  NAND2_X1 U18698 ( .A1(n15236), .A2(n15235), .ZN(n15238) );
  MUX2_X1 U18699 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B(n12892), .S(
        n9844), .Z(n15237) );
  XNOR2_X1 U18700 ( .A(n15238), .B(n15237), .ZN(n16372) );
  NAND2_X1 U18701 ( .A1(n16372), .A2(n20248), .ZN(n15241) );
  AND2_X1 U18702 ( .A1(n20296), .A2(P1_REIP_REG_14__SCAN_IN), .ZN(n16370) );
  NOR2_X1 U18703 ( .A1(n16267), .A2(n20252), .ZN(n15239) );
  AOI211_X1 U18704 ( .C1(n20242), .C2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n16370), .B(n15239), .ZN(n15240) );
  OAI211_X1 U18705 ( .C1(n20306), .C2(n16265), .A(n15241), .B(n15240), .ZN(
        P1_U2985) );
  OAI21_X1 U18706 ( .B1(n15219), .B2(n15243), .A(n15242), .ZN(n15257) );
  INV_X1 U18707 ( .A(n15246), .ZN(n15245) );
  NAND2_X1 U18708 ( .A1(n15245), .A2(n15244), .ZN(n15256) );
  NOR2_X1 U18709 ( .A1(n15257), .A2(n15256), .ZN(n15255) );
  NOR2_X1 U18710 ( .A1(n15255), .A2(n15246), .ZN(n15247) );
  XOR2_X1 U18711 ( .A(n15248), .B(n15247), .Z(n15447) );
  INV_X1 U18712 ( .A(n15249), .ZN(n15251) );
  NAND2_X1 U18713 ( .A1(n20280), .A2(P1_REIP_REG_13__SCAN_IN), .ZN(n15439) );
  NAND2_X1 U18714 ( .A1(n20242), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n15250) );
  OAI211_X1 U18715 ( .C1(n15251), .C2(n20252), .A(n15439), .B(n15250), .ZN(
        n15252) );
  AOI21_X1 U18716 ( .B1(n15253), .B2(n16325), .A(n15252), .ZN(n15254) );
  OAI21_X1 U18717 ( .B1(n15447), .B2(n20088), .A(n15254), .ZN(P1_U2986) );
  AOI21_X1 U18718 ( .B1(n15257), .B2(n15256), .A(n15255), .ZN(n15457) );
  INV_X1 U18719 ( .A(n15258), .ZN(n16281) );
  AOI22_X1 U18720 ( .A1(n20242), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        n20296), .B2(P1_REIP_REG_12__SCAN_IN), .ZN(n15259) );
  OAI21_X1 U18721 ( .B1(n15260), .B2(n20252), .A(n15259), .ZN(n15261) );
  AOI21_X1 U18722 ( .B1(n16281), .B2(n16325), .A(n15261), .ZN(n15262) );
  OAI21_X1 U18723 ( .B1(n15457), .B2(n20088), .A(n15262), .ZN(P1_U2987) );
  NAND2_X1 U18724 ( .A1(n15263), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n15265) );
  XNOR2_X1 U18725 ( .A(n15219), .B(n15266), .ZN(n15264) );
  MUX2_X1 U18726 ( .A(n15265), .B(n15264), .S(n9845), .Z(n15268) );
  INV_X1 U18727 ( .A(n15263), .ZN(n15267) );
  NAND3_X1 U18728 ( .A1(n15267), .A2(n16302), .A3(n15266), .ZN(n16321) );
  NAND2_X1 U18729 ( .A1(n15268), .A2(n16321), .ZN(n16387) );
  NAND2_X1 U18730 ( .A1(n16387), .A2(n20248), .ZN(n15272) );
  AND2_X1 U18731 ( .A1(n20296), .A2(P1_REIP_REG_10__SCAN_IN), .ZN(n16385) );
  NOR2_X1 U18732 ( .A1(n20252), .A2(n15269), .ZN(n15270) );
  AOI211_X1 U18733 ( .C1(n20242), .C2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n16385), .B(n15270), .ZN(n15271) );
  OAI211_X1 U18734 ( .C1(n20306), .C2(n15273), .A(n15272), .B(n15271), .ZN(
        P1_U2989) );
  INV_X1 U18735 ( .A(n15274), .ZN(n15301) );
  NOR3_X1 U18736 ( .A1(n15266), .A2(n16390), .A3(n15275), .ZN(n16380) );
  NAND2_X1 U18737 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n16380), .ZN(
        n15452) );
  NOR2_X1 U18738 ( .A1(n15452), .A2(n15453), .ZN(n15381) );
  NAND2_X1 U18739 ( .A1(n15381), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n16369) );
  INV_X1 U18740 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15432) );
  NAND3_X1 U18741 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n16348) );
  NOR2_X1 U18742 ( .A1(n15432), .A2(n16348), .ZN(n15429) );
  NAND2_X1 U18743 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n15429), .ZN(
        n15281) );
  NOR2_X1 U18744 ( .A1(n16369), .A2(n15281), .ZN(n15280) );
  INV_X1 U18745 ( .A(n15276), .ZN(n15277) );
  AND2_X1 U18746 ( .A1(n15280), .A2(n15277), .ZN(n15278) );
  NOR2_X1 U18747 ( .A1(n15344), .A2(n15348), .ZN(n15279) );
  NAND3_X1 U18748 ( .A1(n15340), .A2(n15314), .A3(
        P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15307) );
  NAND2_X1 U18749 ( .A1(n21115), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15299) );
  AND2_X1 U18750 ( .A1(n15280), .A2(n16426), .ZN(n15286) );
  NAND2_X1 U18751 ( .A1(n15381), .A2(n15448), .ZN(n15426) );
  NOR2_X1 U18752 ( .A1(n15425), .A2(n15281), .ZN(n15386) );
  INV_X1 U18753 ( .A(n15386), .ZN(n15282) );
  OR2_X1 U18754 ( .A1(n15426), .A2(n15282), .ZN(n15283) );
  NAND2_X1 U18755 ( .A1(n16400), .A2(n15283), .ZN(n15285) );
  OAI211_X1 U18756 ( .C1(n15286), .C2(n20253), .A(n15285), .B(n15284), .ZN(
        n15418) );
  INV_X1 U18757 ( .A(n15287), .ZN(n15388) );
  NOR2_X1 U18758 ( .A1(n15418), .A2(n15388), .ZN(n15288) );
  OR2_X1 U18759 ( .A1(n15313), .A2(n15288), .ZN(n15398) );
  INV_X1 U18760 ( .A(n15289), .ZN(n15389) );
  NAND2_X1 U18761 ( .A1(n20276), .A2(n15389), .ZN(n15290) );
  INV_X1 U18762 ( .A(n15347), .ZN(n15291) );
  NAND2_X1 U18763 ( .A1(n20276), .A2(n15291), .ZN(n15292) );
  AND2_X1 U18764 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15293) );
  NAND2_X1 U18765 ( .A1(n15356), .A2(n15293), .ZN(n15294) );
  INV_X1 U18766 ( .A(n15313), .ZN(n15296) );
  NAND2_X1 U18767 ( .A1(n15294), .A2(n15296), .ZN(n15335) );
  NAND2_X1 U18768 ( .A1(n15335), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15318) );
  INV_X1 U18769 ( .A(n15314), .ZN(n15330) );
  NOR2_X1 U18770 ( .A1(n15318), .A2(n15330), .ZN(n15295) );
  OAI21_X1 U18771 ( .B1(n15295), .B2(n15313), .A(
        P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15305) );
  NAND3_X1 U18772 ( .A1(n15305), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n15296), .ZN(n15297) );
  OAI211_X1 U18773 ( .C1(n15307), .C2(n15299), .A(n15298), .B(n15297), .ZN(
        n15300) );
  AOI21_X1 U18774 ( .B1(n15301), .B2(n20282), .A(n15300), .ZN(n15302) );
  OAI21_X1 U18775 ( .B1(n15303), .B2(n20293), .A(n15302), .ZN(P1_U3000) );
  INV_X1 U18776 ( .A(n15304), .ZN(n15309) );
  INV_X1 U18777 ( .A(n15305), .ZN(n15306) );
  AOI21_X1 U18778 ( .B1(n15307), .B2(n13004), .A(n15306), .ZN(n15308) );
  AOI211_X1 U18779 ( .C1(n15310), .C2(n20282), .A(n15309), .B(n15308), .ZN(
        n15311) );
  OAI21_X1 U18780 ( .B1(n15312), .B2(n20293), .A(n15311), .ZN(P1_U3001) );
  NOR2_X1 U18781 ( .A1(n15313), .A2(n15314), .ZN(n15319) );
  NAND2_X1 U18782 ( .A1(n15340), .A2(n15314), .ZN(n15316) );
  NAND2_X1 U18783 ( .A1(n15316), .A2(n15315), .ZN(n15317) );
  OAI21_X1 U18784 ( .B1(n15319), .B2(n15318), .A(n15317), .ZN(n15321) );
  OAI211_X1 U18785 ( .C1(n15322), .C2(n20292), .A(n15321), .B(n15320), .ZN(
        n15323) );
  INV_X1 U18786 ( .A(n15323), .ZN(n15324) );
  OAI21_X1 U18787 ( .B1(n15325), .B2(n20293), .A(n15324), .ZN(P1_U3002) );
  OAI21_X1 U18788 ( .B1(n15335), .B2(n15327), .A(n15326), .ZN(n15328) );
  AOI21_X1 U18789 ( .B1(n15329), .B2(n20282), .A(n15328), .ZN(n15333) );
  NAND3_X1 U18790 ( .A1(n15340), .A2(n15331), .A3(n15330), .ZN(n15332) );
  OAI211_X1 U18791 ( .C1(n15334), .C2(n20293), .A(n15333), .B(n15332), .ZN(
        P1_U3003) );
  NOR2_X1 U18792 ( .A1(n15335), .A2(n15339), .ZN(n15336) );
  AOI211_X1 U18793 ( .C1(n15338), .C2(n20282), .A(n15337), .B(n15336), .ZN(
        n15342) );
  NAND2_X1 U18794 ( .A1(n15340), .A2(n15339), .ZN(n15341) );
  OAI211_X1 U18795 ( .C1(n15343), .C2(n20293), .A(n15342), .B(n15341), .ZN(
        P1_U3004) );
  NOR2_X1 U18796 ( .A1(n15344), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15351) );
  OAI21_X1 U18797 ( .B1(n15346), .B2(n20292), .A(n15345), .ZN(n15350) );
  NAND3_X1 U18798 ( .A1(n15378), .A2(n15347), .A3(n15355), .ZN(n15359) );
  AOI21_X1 U18799 ( .B1(n15359), .B2(n15356), .A(n15348), .ZN(n15349) );
  AOI211_X1 U18800 ( .C1(n15378), .C2(n15351), .A(n15350), .B(n15349), .ZN(
        n15352) );
  OAI21_X1 U18801 ( .B1(n15353), .B2(n20293), .A(n15352), .ZN(P1_U3005) );
  OAI21_X1 U18802 ( .B1(n15356), .B2(n15355), .A(n15354), .ZN(n15357) );
  AOI21_X1 U18803 ( .B1(n15358), .B2(n20282), .A(n15357), .ZN(n15360) );
  OAI211_X1 U18804 ( .C1(n15361), .C2(n20293), .A(n15360), .B(n15359), .ZN(
        P1_U3006) );
  AND3_X1 U18805 ( .A1(n15378), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        n15362), .ZN(n15363) );
  AOI211_X1 U18806 ( .C1(n20282), .C2(n15365), .A(n15364), .B(n15363), .ZN(
        n15370) );
  AOI21_X1 U18807 ( .B1(n15366), .B2(n20253), .A(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15368) );
  INV_X1 U18808 ( .A(n15367), .ZN(n15372) );
  OAI21_X1 U18809 ( .B1(n15368), .B2(n15372), .A(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15369) );
  OAI211_X1 U18810 ( .C1(n15371), .C2(n20293), .A(n15370), .B(n15369), .ZN(
        P1_U3007) );
  NAND2_X1 U18811 ( .A1(n15372), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15373) );
  OAI211_X1 U18812 ( .C1(n15375), .C2(n20292), .A(n15374), .B(n15373), .ZN(
        n15376) );
  AOI21_X1 U18813 ( .B1(n15378), .B2(n15377), .A(n15376), .ZN(n15379) );
  OAI21_X1 U18814 ( .B1(n15380), .B2(n20293), .A(n15379), .ZN(P1_U3008) );
  INV_X1 U18815 ( .A(n15381), .ZN(n15384) );
  INV_X1 U18816 ( .A(n15426), .ZN(n15382) );
  NAND3_X1 U18817 ( .A1(n20288), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A3(
        n15382), .ZN(n15383) );
  OAI21_X1 U18818 ( .B1(n15385), .B2(n15384), .A(n15383), .ZN(n15444) );
  NOR2_X1 U18819 ( .A1(n20298), .A2(n15426), .ZN(n15438) );
  OR2_X1 U18820 ( .A1(n15444), .A2(n15438), .ZN(n15387) );
  NAND2_X1 U18821 ( .A1(n15387), .A2(n15386), .ZN(n15420) );
  NOR2_X1 U18822 ( .A1(n15420), .A2(n15388), .ZN(n15403) );
  OAI211_X1 U18823 ( .C1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A(n15403), .B(n15389), .ZN(
        n15391) );
  OAI211_X1 U18824 ( .C1(n15398), .C2(n15392), .A(n15391), .B(n15390), .ZN(
        n15393) );
  AOI21_X1 U18825 ( .B1(n15394), .B2(n20282), .A(n15393), .ZN(n15395) );
  OAI21_X1 U18826 ( .B1(n15396), .B2(n20293), .A(n15395), .ZN(P1_U3009) );
  OAI21_X1 U18827 ( .B1(n15398), .B2(n15402), .A(n15397), .ZN(n15401) );
  NOR2_X1 U18828 ( .A1(n15399), .A2(n20292), .ZN(n15400) );
  AOI211_X1 U18829 ( .C1(n15403), .C2(n15402), .A(n15401), .B(n15400), .ZN(
        n15404) );
  OAI21_X1 U18830 ( .B1(n15405), .B2(n20293), .A(n15404), .ZN(P1_U3010) );
  NAND2_X1 U18831 ( .A1(n15406), .A2(n20278), .ZN(n15415) );
  INV_X1 U18832 ( .A(n20298), .ZN(n15407) );
  NOR2_X1 U18833 ( .A1(n15444), .A2(n15407), .ZN(n15409) );
  INV_X1 U18834 ( .A(n15418), .ZN(n15408) );
  OAI21_X1 U18835 ( .B1(n15409), .B2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n15408), .ZN(n15413) );
  NOR3_X1 U18836 ( .A1(n15420), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A3(
        n15410), .ZN(n15411) );
  AOI211_X1 U18837 ( .C1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .C2(n15413), .A(
        n15412), .B(n15411), .ZN(n15414) );
  OAI211_X1 U18838 ( .C1(n20292), .C2(n15416), .A(n15415), .B(n15414), .ZN(
        P1_U3011) );
  INV_X1 U18839 ( .A(n16246), .ZN(n15422) );
  AOI21_X1 U18840 ( .B1(n15418), .B2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n15417), .ZN(n15419) );
  OAI21_X1 U18841 ( .B1(n15420), .B2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n15419), .ZN(n15421) );
  AOI21_X1 U18842 ( .B1(n15422), .B2(n20282), .A(n15421), .ZN(n15423) );
  OAI21_X1 U18843 ( .B1(n15424), .B2(n20293), .A(n15423), .ZN(P1_U3012) );
  INV_X1 U18844 ( .A(n20276), .ZN(n16402) );
  INV_X1 U18845 ( .A(n16400), .ZN(n20254) );
  NOR2_X1 U18846 ( .A1(n15426), .A2(n15425), .ZN(n15440) );
  INV_X1 U18847 ( .A(n16398), .ZN(n15427) );
  OAI21_X1 U18848 ( .B1(n20254), .B2(n15440), .A(n15427), .ZN(n15428) );
  AOI21_X1 U18849 ( .B1(n20289), .B2(n16369), .A(n15428), .ZN(n16357) );
  OAI21_X1 U18850 ( .B1(n16402), .B2(n15429), .A(n16357), .ZN(n16349) );
  INV_X1 U18851 ( .A(P1_REIP_REG_18__SCAN_IN), .ZN(n20955) );
  OAI22_X1 U18852 ( .A1(n16255), .A2(n20292), .B1(n20955), .B2(n20256), .ZN(
        n15430) );
  AOI21_X1 U18853 ( .B1(n16349), .B2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n15430), .ZN(n15436) );
  NOR4_X1 U18854 ( .A1(n16421), .A2(n16369), .A3(n15432), .A4(n16348), .ZN(
        n15434) );
  NAND2_X1 U18855 ( .A1(n15434), .A2(n15433), .ZN(n15435) );
  OAI211_X1 U18856 ( .C1(n15437), .C2(n20293), .A(n15436), .B(n15435), .ZN(
        P1_U3013) );
  INV_X1 U18857 ( .A(n15438), .ZN(n15441) );
  OAI21_X1 U18858 ( .B1(n15441), .B2(n15440), .A(n15439), .ZN(n15442) );
  AOI21_X1 U18859 ( .B1(n15443), .B2(n20282), .A(n15442), .ZN(n15446) );
  INV_X1 U18860 ( .A(n16357), .ZN(n16373) );
  OAI21_X1 U18861 ( .B1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n15444), .A(
        n16373), .ZN(n15445) );
  OAI211_X1 U18862 ( .C1(n15447), .C2(n20293), .A(n15446), .B(n15445), .ZN(
        P1_U3018) );
  AOI21_X1 U18863 ( .B1(n16380), .B2(n15448), .A(n20254), .ZN(n15449) );
  AOI211_X1 U18864 ( .C1(n20289), .C2(n15452), .A(n15449), .B(n16398), .ZN(
        n16384) );
  OAI21_X1 U18865 ( .B1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n20258), .A(
        n16384), .ZN(n15451) );
  OAI22_X1 U18866 ( .A1(n16275), .A2(n20292), .B1(n20944), .B2(n20256), .ZN(
        n15450) );
  AOI21_X1 U18867 ( .B1(n15451), .B2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n15450), .ZN(n15456) );
  NOR2_X1 U18868 ( .A1(n16421), .A2(n15452), .ZN(n15454) );
  NAND2_X1 U18869 ( .A1(n15454), .A2(n15453), .ZN(n15455) );
  OAI211_X1 U18870 ( .C1(n15457), .C2(n20293), .A(n15456), .B(n15455), .ZN(
        P1_U3019) );
  NAND2_X1 U18871 ( .A1(n20700), .A2(n20769), .ZN(n15460) );
  NOR2_X1 U18872 ( .A1(n9853), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n15458) );
  OAI22_X1 U18873 ( .A1(n15460), .A2(n15458), .B1(n13838), .B2(n15462), .ZN(
        n15459) );
  MUX2_X1 U18874 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n15459), .S(
        n20301), .Z(P1_U3477) );
  MUX2_X1 U18875 ( .A(n15460), .B(n20854), .S(n20593), .Z(n15461) );
  OAI21_X1 U18876 ( .B1(n15462), .B2(n13553), .A(n15461), .ZN(n15463) );
  MUX2_X1 U18877 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n15463), .S(
        n20301), .Z(P1_U3476) );
  INV_X1 U18878 ( .A(n15472), .ZN(n15465) );
  INV_X1 U18879 ( .A(n13958), .ZN(n15464) );
  NAND3_X1 U18880 ( .A1(n15466), .A2(n15465), .A3(n15464), .ZN(n15467) );
  OAI21_X1 U18881 ( .B1(n15468), .B2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n15467), .ZN(n15469) );
  AOI21_X1 U18882 ( .B1(n20799), .B2(n15470), .A(n15469), .ZN(n16171) );
  INV_X1 U18883 ( .A(n15471), .ZN(n15475) );
  NOR3_X1 U18884 ( .A1(n13958), .A2(n15472), .A3(n15481), .ZN(n15473) );
  AOI21_X1 U18885 ( .B1(n15475), .B2(n15474), .A(n15473), .ZN(n15476) );
  OAI21_X1 U18886 ( .B1(n16171), .B2(n15482), .A(n15476), .ZN(n15478) );
  MUX2_X1 U18887 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n15478), .S(
        n15477), .Z(P1_U3473) );
  INV_X1 U18888 ( .A(n15479), .ZN(n15480) );
  OAI22_X1 U18889 ( .A1(n15483), .A2(n15482), .B1(n15481), .B2(n15480), .ZN(
        n15485) );
  MUX2_X1 U18890 ( .A(n15485), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n15484), .Z(P1_U3469) );
  NOR2_X1 U18891 ( .A1(n19159), .A2(n19214), .ZN(n15586) );
  NAND2_X1 U18892 ( .A1(n15486), .A2(n15586), .ZN(n15493) );
  NAND2_X1 U18893 ( .A1(n19210), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n15489) );
  AOI22_X1 U18894 ( .A1(n15487), .A2(P2_EBX_REG_31__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n19166), .ZN(n15488) );
  OAI211_X1 U18895 ( .C1(n19216), .C2(n19200), .A(n15489), .B(n15488), .ZN(
        n15490) );
  AOI21_X1 U18896 ( .B1(n15491), .B2(n19186), .A(n15490), .ZN(n15492) );
  OAI211_X1 U18897 ( .C1(n15494), .C2(n19197), .A(n15493), .B(n15492), .ZN(
        P2_U2824) );
  AOI22_X1 U18898 ( .A1(P2_REIP_REG_29__SCAN_IN), .A2(n19210), .B1(
        P2_EBX_REG_29__SCAN_IN), .B2(n19205), .ZN(n15497) );
  AOI22_X1 U18899 ( .A1(n15495), .A2(n19186), .B1(
        P2_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n19166), .ZN(n15496) );
  OAI211_X1 U18900 ( .C1(n15697), .C2(n19200), .A(n15497), .B(n15496), .ZN(
        n15502) );
  AOI211_X1 U18901 ( .C1(n15500), .C2(n15499), .A(n15498), .B(n19214), .ZN(
        n15501) );
  NOR2_X1 U18902 ( .A1(n15502), .A2(n15501), .ZN(n15503) );
  OAI21_X1 U18903 ( .B1(n15630), .B2(n19197), .A(n15503), .ZN(P2_U2826) );
  OR2_X1 U18904 ( .A1(n13316), .A2(n15504), .ZN(n15505) );
  NAND2_X1 U18905 ( .A1(n12486), .A2(n15505), .ZN(n15869) );
  AOI211_X1 U18906 ( .C1(n15758), .C2(n15507), .A(n15506), .B(n19214), .ZN(
        n15508) );
  INV_X1 U18907 ( .A(n15508), .ZN(n15517) );
  AND2_X1 U18908 ( .A1(n9886), .A2(n15509), .ZN(n15511) );
  OR2_X1 U18909 ( .A1(n15511), .A2(n15510), .ZN(n15871) );
  NAND2_X1 U18910 ( .A1(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n19211), .ZN(
        n15513) );
  AOI22_X1 U18911 ( .A1(P2_REIP_REG_28__SCAN_IN), .A2(n19210), .B1(
        P2_EBX_REG_28__SCAN_IN), .B2(n19205), .ZN(n15512) );
  OAI211_X1 U18912 ( .C1(n19200), .C2(n15871), .A(n15513), .B(n15512), .ZN(
        n15514) );
  AOI21_X1 U18913 ( .B1(n15515), .B2(n19186), .A(n15514), .ZN(n15516) );
  OAI211_X1 U18914 ( .C1(n19197), .C2(n15869), .A(n15517), .B(n15516), .ZN(
        P2_U2827) );
  AOI211_X1 U18915 ( .C1(n15519), .C2(n15786), .A(n19214), .B(n15518), .ZN(
        n15520) );
  INV_X1 U18916 ( .A(n15520), .ZN(n15529) );
  INV_X1 U18917 ( .A(n15643), .ZN(n15521) );
  AOI21_X1 U18918 ( .B1(n15522), .B2(n15540), .A(n15521), .ZN(n15917) );
  AND2_X1 U18919 ( .A1(n15544), .A2(n15523), .ZN(n15524) );
  NOR2_X1 U18920 ( .A1(n15719), .A2(n15524), .ZN(n15907) );
  NAND2_X1 U18921 ( .A1(n19183), .A2(n15907), .ZN(n15526) );
  AOI22_X1 U18922 ( .A1(P2_REIP_REG_25__SCAN_IN), .A2(n19210), .B1(
        P2_EBX_REG_25__SCAN_IN), .B2(n19205), .ZN(n15525) );
  OAI211_X1 U18923 ( .C1(n19180), .C2(n15788), .A(n15526), .B(n15525), .ZN(
        n15527) );
  AOI21_X1 U18924 ( .B1(n15917), .B2(n19179), .A(n15527), .ZN(n15528) );
  OAI211_X1 U18925 ( .C1(n19202), .C2(n15530), .A(n15529), .B(n15528), .ZN(
        P2_U2830) );
  AOI211_X1 U18926 ( .C1(n15533), .C2(n15532), .A(n15531), .B(n19214), .ZN(
        n15535) );
  INV_X1 U18927 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n19972) );
  OAI22_X1 U18928 ( .A1(n19155), .A2(n10183), .B1(n19972), .B2(n19181), .ZN(
        n15534) );
  AOI211_X1 U18929 ( .C1(n19211), .C2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n15535), .B(n15534), .ZN(n15548) );
  XNOR2_X1 U18930 ( .A(n15536), .B(n10183), .ZN(n15546) );
  OR2_X1 U18931 ( .A1(n15537), .A2(n15538), .ZN(n15539) );
  NAND2_X1 U18932 ( .A1(n15540), .A2(n15539), .ZN(n15926) );
  NAND2_X1 U18933 ( .A1(n15541), .A2(n15542), .ZN(n15543) );
  NAND2_X1 U18934 ( .A1(n15544), .A2(n15543), .ZN(n15925) );
  OAI22_X1 U18935 ( .A1(n15926), .A2(n19197), .B1(n19200), .B2(n15925), .ZN(
        n15545) );
  AOI21_X1 U18936 ( .B1(n15546), .B2(n19186), .A(n15545), .ZN(n15547) );
  NAND2_X1 U18937 ( .A1(n15548), .A2(n15547), .ZN(P2_U2831) );
  AOI211_X1 U18938 ( .C1(n16472), .C2(n15550), .A(n15549), .B(n19214), .ZN(
        n15552) );
  INV_X1 U18939 ( .A(P2_EBX_REG_23__SCAN_IN), .ZN(n15670) );
  OAI22_X1 U18940 ( .A1(n19155), .A2(n15670), .B1(n19970), .B2(n19181), .ZN(
        n15551) );
  AOI211_X1 U18941 ( .C1(n19211), .C2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n15552), .B(n15551), .ZN(n15560) );
  NOR2_X1 U18942 ( .A1(n15553), .A2(n15554), .ZN(n15555) );
  OR2_X1 U18943 ( .A1(n15537), .A2(n15555), .ZN(n15666) );
  OAI21_X1 U18944 ( .B1(n15572), .B2(n15556), .A(n15541), .ZN(n15942) );
  OAI22_X1 U18945 ( .A1(n15666), .A2(n19197), .B1(n19200), .B2(n15942), .ZN(
        n15557) );
  AOI21_X1 U18946 ( .B1(n15558), .B2(n19186), .A(n15557), .ZN(n15559) );
  NAND2_X1 U18947 ( .A1(n15560), .A2(n15559), .ZN(P2_U2832) );
  OAI21_X1 U18948 ( .B1(n16484), .B2(n15561), .A(n19175), .ZN(n15563) );
  AOI22_X1 U18949 ( .A1(P2_REIP_REG_22__SCAN_IN), .A2(n19210), .B1(
        P2_EBX_REG_22__SCAN_IN), .B2(n19205), .ZN(n15562) );
  OAI21_X1 U18950 ( .B1(n15564), .B2(n15563), .A(n15562), .ZN(n15565) );
  AOI21_X1 U18951 ( .B1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n19211), .A(
        n15565), .ZN(n15574) );
  INV_X1 U18952 ( .A(n15566), .ZN(n15568) );
  INV_X1 U18953 ( .A(n15553), .ZN(n15567) );
  OAI21_X1 U18954 ( .B1(n10159), .B2(n15568), .A(n15567), .ZN(n15959) );
  INV_X1 U18955 ( .A(n15959), .ZN(n16481) );
  NOR2_X1 U18956 ( .A1(n15570), .A2(n15569), .ZN(n15571) );
  NOR2_X1 U18957 ( .A1(n15572), .A2(n15571), .ZN(n16457) );
  AOI22_X1 U18958 ( .A1(n16481), .A2(n19179), .B1(n19183), .B2(n16457), .ZN(
        n15573) );
  OAI211_X1 U18959 ( .C1(n15575), .C2(n19202), .A(n15574), .B(n15573), .ZN(
        P2_U2833) );
  AND2_X1 U18960 ( .A1(n10135), .A2(n15585), .ZN(n15577) );
  OAI21_X1 U18961 ( .B1(n15805), .B2(n15577), .A(n19175), .ZN(n15576) );
  AOI21_X1 U18962 ( .B1(n15805), .B2(n15577), .A(n15576), .ZN(n15579) );
  OAI22_X1 U18963 ( .A1(n15808), .A2(n19180), .B1(n19966), .B2(n19181), .ZN(
        n15578) );
  AOI211_X1 U18964 ( .C1(P2_EBX_REG_21__SCAN_IN), .C2(n19205), .A(n15579), .B(
        n15578), .ZN(n15582) );
  INV_X1 U18965 ( .A(n15745), .ZN(n15580) );
  AOI22_X1 U18966 ( .A1(n15812), .A2(n19179), .B1(n15580), .B2(n19183), .ZN(
        n15581) );
  OAI211_X1 U18967 ( .C1(n15583), .C2(n19202), .A(n15582), .B(n15581), .ZN(
        P2_U2834) );
  INV_X1 U18968 ( .A(n15823), .ZN(n15584) );
  NOR2_X1 U18969 ( .A1(n10135), .A2(n19214), .ZN(n19192) );
  AOI22_X1 U18970 ( .A1(P2_EBX_REG_20__SCAN_IN), .A2(n19205), .B1(n15584), 
        .B2(n19192), .ZN(n15598) );
  OAI211_X1 U18971 ( .C1(n15587), .C2(n15823), .A(n15586), .B(n15585), .ZN(
        n15597) );
  OR2_X1 U18972 ( .A1(n15691), .A2(n15588), .ZN(n15589) );
  NAND2_X1 U18973 ( .A1(n9863), .A2(n15589), .ZN(n15968) );
  AOI22_X1 U18974 ( .A1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n19166), .B1(
        P2_REIP_REG_20__SCAN_IN), .B2(n19210), .ZN(n15593) );
  NOR2_X1 U18975 ( .A1(n9941), .A2(n15590), .ZN(n15591) );
  NAND2_X1 U18976 ( .A1(n19183), .A2(n9921), .ZN(n15592) );
  OAI211_X1 U18977 ( .C1(n15968), .C2(n19197), .A(n15593), .B(n15592), .ZN(
        n15594) );
  AOI21_X1 U18978 ( .B1(n15595), .B2(n19186), .A(n15594), .ZN(n15596) );
  NAND3_X1 U18979 ( .A1(n15598), .A2(n15597), .A3(n15596), .ZN(P2_U2835) );
  NOR2_X1 U18980 ( .A1(n19159), .A2(n15599), .ZN(n15600) );
  XNOR2_X1 U18981 ( .A(n15600), .B(n16490), .ZN(n15601) );
  NAND2_X1 U18982 ( .A1(n15601), .A2(n19175), .ZN(n15609) );
  NAND2_X1 U18983 ( .A1(n14242), .A2(n15602), .ZN(n15603) );
  NAND2_X1 U18984 ( .A1(n15604), .A2(n15603), .ZN(n16466) );
  AOI22_X1 U18985 ( .A1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n19166), .B1(
        P2_EBX_REG_18__SCAN_IN), .B2(n19205), .ZN(n15605) );
  OAI211_X1 U18986 ( .C1(n19200), .C2(n16466), .A(n15605), .B(n19345), .ZN(
        n15607) );
  INV_X1 U18987 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n15994) );
  NOR2_X1 U18988 ( .A1(n19181), .A2(n15994), .ZN(n15606) );
  AOI211_X1 U18989 ( .C1(n16486), .C2(n19179), .A(n15607), .B(n15606), .ZN(
        n15608) );
  OAI211_X1 U18990 ( .C1(n19202), .C2(n15610), .A(n15609), .B(n15608), .ZN(
        P2_U2837) );
  NOR2_X1 U18991 ( .A1(n19159), .A2(n15611), .ZN(n15612) );
  XNOR2_X1 U18992 ( .A(n15612), .B(n16517), .ZN(n15613) );
  NAND2_X1 U18993 ( .A1(n15613), .A2(n19175), .ZN(n15623) );
  INV_X1 U18994 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n19952) );
  INV_X1 U18995 ( .A(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n15614) );
  OAI22_X1 U18996 ( .A1(n15615), .A2(n19202), .B1(n15614), .B2(n19180), .ZN(
        n15616) );
  INV_X1 U18997 ( .A(n15616), .ZN(n15617) );
  OAI211_X1 U18998 ( .C1(n19952), .C2(n19181), .A(n15617), .B(n19345), .ZN(
        n15618) );
  AOI21_X1 U18999 ( .B1(P2_EBX_REG_12__SCAN_IN), .B2(n19205), .A(n15618), .ZN(
        n15622) );
  AOI21_X1 U19000 ( .B1(n15620), .B2(n16074), .A(n15619), .ZN(n19238) );
  AOI22_X1 U19001 ( .A1(n19179), .A2(n16565), .B1(n19183), .B2(n19238), .ZN(
        n15621) );
  NAND3_X1 U19002 ( .A1(n15623), .A2(n15622), .A3(n15621), .ZN(P2_U2843) );
  MUX2_X1 U19003 ( .A(n15624), .B(P2_EBX_REG_31__SCAN_IN), .S(n15667), .Z(
        P2_U2856) );
  OR2_X1 U19004 ( .A1(n15626), .A2(n15625), .ZN(n15696) );
  NAND3_X1 U19005 ( .A1(n15696), .A2(n15627), .A3(n15685), .ZN(n15629) );
  NAND2_X1 U19006 ( .A1(n15667), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n15628) );
  OAI211_X1 U19007 ( .C1(n15667), .C2(n15630), .A(n15629), .B(n15628), .ZN(
        P2_U2858) );
  NAND2_X1 U19008 ( .A1(n15632), .A2(n15631), .ZN(n15634) );
  XNOR2_X1 U19009 ( .A(n15634), .B(n15633), .ZN(n15707) );
  NAND2_X1 U19010 ( .A1(n15707), .A2(n15685), .ZN(n15636) );
  NAND2_X1 U19011 ( .A1(n15667), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n15635) );
  OAI211_X1 U19012 ( .C1(n15869), .C2(n15661), .A(n15636), .B(n15635), .ZN(
        P2_U2859) );
  OAI21_X1 U19013 ( .B1(n9832), .B2(n15639), .A(n15638), .ZN(n15715) );
  NOR2_X1 U19014 ( .A1(n15889), .A2(n15661), .ZN(n15640) );
  AOI21_X1 U19015 ( .B1(P2_EBX_REG_27__SCAN_IN), .B2(n15661), .A(n15640), .ZN(
        n15641) );
  OAI21_X1 U19016 ( .B1(n15715), .B2(n15694), .A(n15641), .ZN(P2_U2860) );
  AND2_X1 U19017 ( .A1(n15643), .A2(n15642), .ZN(n15644) );
  AOI21_X1 U19018 ( .B1(n15647), .B2(n15646), .A(n15645), .ZN(n15716) );
  NAND2_X1 U19019 ( .A1(n15716), .A2(n15685), .ZN(n15649) );
  NAND2_X1 U19020 ( .A1(n15667), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n15648) );
  OAI211_X1 U19021 ( .C1(n16452), .C2(n15667), .A(n15649), .B(n15648), .ZN(
        P2_U2861) );
  OAI21_X1 U19022 ( .B1(n15652), .B2(n15651), .A(n15650), .ZN(n15731) );
  NOR2_X1 U19023 ( .A1(n14287), .A2(n15653), .ZN(n15654) );
  AOI21_X1 U19024 ( .B1(n15917), .B2(n14287), .A(n15654), .ZN(n15655) );
  OAI21_X1 U19025 ( .B1(n15731), .B2(n15694), .A(n15655), .ZN(P2_U2862) );
  AOI21_X1 U19026 ( .B1(n15656), .B2(n15657), .A(n9928), .ZN(n15658) );
  XOR2_X1 U19027 ( .A(n15659), .B(n15658), .Z(n15736) );
  NOR2_X1 U19028 ( .A1(n15926), .A2(n15661), .ZN(n15660) );
  AOI21_X1 U19029 ( .B1(P2_EBX_REG_24__SCAN_IN), .B2(n15661), .A(n15660), .ZN(
        n15662) );
  OAI21_X1 U19030 ( .B1(n15736), .B2(n15694), .A(n15662), .ZN(P2_U2863) );
  AOI21_X1 U19031 ( .B1(n15665), .B2(n15664), .A(n15663), .ZN(n15741) );
  NAND2_X1 U19032 ( .A1(n15741), .A2(n15685), .ZN(n15669) );
  NAND2_X1 U19033 ( .A1(n16476), .A2(n14287), .ZN(n15668) );
  OAI211_X1 U19034 ( .C1(n14287), .C2(n15670), .A(n15669), .B(n15668), .ZN(
        P2_U2864) );
  INV_X1 U19035 ( .A(n15671), .ZN(n15675) );
  INV_X1 U19036 ( .A(n15672), .ZN(n15674) );
  AOI21_X1 U19037 ( .B1(n15675), .B2(n15674), .A(n15673), .ZN(n16458) );
  NAND2_X1 U19038 ( .A1(n16458), .A2(n15685), .ZN(n15677) );
  NAND2_X1 U19039 ( .A1(n15661), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n15676) );
  OAI211_X1 U19040 ( .C1(n15959), .C2(n15667), .A(n15677), .B(n15676), .ZN(
        P2_U2865) );
  AOI21_X1 U19041 ( .B1(n15679), .B2(n15682), .A(n15672), .ZN(n15747) );
  NAND2_X1 U19042 ( .A1(n15747), .A2(n15685), .ZN(n15681) );
  NAND2_X1 U19043 ( .A1(n15812), .A2(n14287), .ZN(n15680) );
  OAI211_X1 U19044 ( .C1(n14287), .C2(n10189), .A(n15681), .B(n15680), .ZN(
        P2_U2866) );
  INV_X1 U19045 ( .A(n15682), .ZN(n15683) );
  AOI21_X1 U19046 ( .B1(n15684), .B2(n14543), .A(n15683), .ZN(n16462) );
  NAND2_X1 U19047 ( .A1(n16462), .A2(n15685), .ZN(n15687) );
  NAND2_X1 U19048 ( .A1(n15661), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n15686) );
  OAI211_X1 U19049 ( .C1(n15968), .C2(n15667), .A(n15687), .B(n15686), .ZN(
        P2_U2867) );
  NAND2_X1 U19050 ( .A1(n15661), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n15693) );
  AND2_X1 U19051 ( .A1(n15689), .A2(n15688), .ZN(n15690) );
  NOR2_X1 U19052 ( .A1(n15691), .A2(n15690), .ZN(n19070) );
  NAND2_X1 U19053 ( .A1(n19070), .A2(n14287), .ZN(n15692) );
  OAI211_X1 U19054 ( .C1(n15695), .C2(n15694), .A(n15693), .B(n15692), .ZN(
        P2_U2868) );
  NAND3_X1 U19055 ( .A1(n15696), .A2(n15627), .A3(n19270), .ZN(n15703) );
  INV_X1 U19056 ( .A(n15697), .ZN(n15700) );
  INV_X1 U19057 ( .A(n19221), .ZN(n15710) );
  OAI22_X1 U19058 ( .A1(n15710), .A2(n19236), .B1(n19274), .B2(n15698), .ZN(
        n15699) );
  AOI21_X1 U19059 ( .B1(n19265), .B2(n15700), .A(n15699), .ZN(n15702) );
  AOI22_X1 U19060 ( .A1(n19223), .A2(BUF2_REG_29__SCAN_IN), .B1(n19222), .B2(
        BUF1_REG_29__SCAN_IN), .ZN(n15701) );
  NAND3_X1 U19061 ( .A1(n15703), .A2(n15702), .A3(n15701), .ZN(P2_U2890) );
  AOI22_X1 U19062 ( .A1(n19223), .A2(BUF2_REG_28__SCAN_IN), .B1(n19222), .B2(
        BUF1_REG_28__SCAN_IN), .ZN(n15705) );
  AOI22_X1 U19063 ( .A1(n19221), .A2(n19239), .B1(n19257), .B2(
        P2_EAX_REG_28__SCAN_IN), .ZN(n15704) );
  OAI211_X1 U19064 ( .C1(n19229), .C2(n15871), .A(n15705), .B(n15704), .ZN(
        n15706) );
  AOI21_X1 U19065 ( .B1(n15707), .B2(n19270), .A(n15706), .ZN(n15708) );
  INV_X1 U19066 ( .A(n15708), .ZN(P2_U2891) );
  INV_X1 U19067 ( .A(n15884), .ZN(n15712) );
  OAI22_X1 U19068 ( .A1(n15710), .A2(n19242), .B1(n19274), .B2(n15709), .ZN(
        n15711) );
  AOI21_X1 U19069 ( .B1(n19265), .B2(n15712), .A(n15711), .ZN(n15714) );
  AOI22_X1 U19070 ( .A1(n19223), .A2(BUF2_REG_27__SCAN_IN), .B1(n19222), .B2(
        BUF1_REG_27__SCAN_IN), .ZN(n15713) );
  OAI211_X1 U19071 ( .C1(n15715), .C2(n19258), .A(n15714), .B(n15713), .ZN(
        P2_U2892) );
  NAND2_X1 U19072 ( .A1(n15716), .A2(n19270), .ZN(n15724) );
  OAI21_X1 U19073 ( .B1(n15719), .B2(n15718), .A(n15717), .ZN(n15720) );
  INV_X1 U19074 ( .A(n15720), .ZN(n16455) );
  AOI22_X1 U19075 ( .A1(n19265), .A2(n16455), .B1(P2_EAX_REG_26__SCAN_IN), 
        .B2(n19257), .ZN(n15723) );
  AOI22_X1 U19076 ( .A1(n19223), .A2(BUF2_REG_26__SCAN_IN), .B1(n19222), .B2(
        BUF1_REG_26__SCAN_IN), .ZN(n15722) );
  NAND2_X1 U19077 ( .A1(n19221), .A2(n19244), .ZN(n15721) );
  NAND4_X1 U19078 ( .A1(n15724), .A2(n15723), .A3(n15722), .A4(n15721), .ZN(
        P2_U2893) );
  INV_X1 U19079 ( .A(n15907), .ZN(n15728) );
  AOI22_X1 U19080 ( .A1(n19223), .A2(BUF2_REG_25__SCAN_IN), .B1(n19222), .B2(
        BUF1_REG_25__SCAN_IN), .ZN(n15727) );
  AOI22_X1 U19081 ( .A1(n19221), .A2(n15725), .B1(n19257), .B2(
        P2_EAX_REG_25__SCAN_IN), .ZN(n15726) );
  OAI211_X1 U19082 ( .C1(n19229), .C2(n15728), .A(n15727), .B(n15726), .ZN(
        n15729) );
  INV_X1 U19083 ( .A(n15729), .ZN(n15730) );
  OAI21_X1 U19084 ( .B1(n15731), .B2(n19258), .A(n15730), .ZN(P2_U2894) );
  AOI22_X1 U19085 ( .A1(n19223), .A2(BUF2_REG_24__SCAN_IN), .B1(n19222), .B2(
        BUF1_REG_24__SCAN_IN), .ZN(n15733) );
  AOI22_X1 U19086 ( .A1(n19221), .A2(n19249), .B1(n19257), .B2(
        P2_EAX_REG_24__SCAN_IN), .ZN(n15732) );
  OAI211_X1 U19087 ( .C1(n19229), .C2(n15925), .A(n15733), .B(n15732), .ZN(
        n15734) );
  INV_X1 U19088 ( .A(n15734), .ZN(n15735) );
  OAI21_X1 U19089 ( .B1(n15736), .B2(n19258), .A(n15735), .ZN(P2_U2895) );
  AOI22_X1 U19090 ( .A1(n19223), .A2(BUF2_REG_23__SCAN_IN), .B1(n19222), .B2(
        BUF1_REG_23__SCAN_IN), .ZN(n15739) );
  AOI22_X1 U19091 ( .A1(n19221), .A2(n15737), .B1(n19257), .B2(
        P2_EAX_REG_23__SCAN_IN), .ZN(n15738) );
  OAI211_X1 U19092 ( .C1(n19229), .C2(n15942), .A(n15739), .B(n15738), .ZN(
        n15740) );
  AOI21_X1 U19093 ( .B1(n15741), .B2(n19270), .A(n15740), .ZN(n15742) );
  INV_X1 U19094 ( .A(n15742), .ZN(P2_U2896) );
  AOI22_X1 U19095 ( .A1(n19223), .A2(BUF2_REG_21__SCAN_IN), .B1(n19222), .B2(
        BUF1_REG_21__SCAN_IN), .ZN(n15744) );
  AOI22_X1 U19096 ( .A1(n19221), .A2(n19403), .B1(n19257), .B2(
        P2_EAX_REG_21__SCAN_IN), .ZN(n15743) );
  OAI211_X1 U19097 ( .C1(n19229), .C2(n15745), .A(n15744), .B(n15743), .ZN(
        n15746) );
  AOI21_X1 U19098 ( .B1(n15747), .B2(n19270), .A(n15746), .ZN(n15748) );
  INV_X1 U19099 ( .A(n15748), .ZN(P2_U2898) );
  XNOR2_X1 U19100 ( .A(n15750), .B(n15752), .ZN(n15762) );
  INV_X1 U19101 ( .A(n15750), .ZN(n15751) );
  AOI22_X1 U19102 ( .A1(n15762), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B1(
        n15752), .B2(n15751), .ZN(n15755) );
  XNOR2_X1 U19103 ( .A(n15753), .B(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n15754) );
  XNOR2_X1 U19104 ( .A(n15755), .B(n15754), .ZN(n15881) );
  XNOR2_X1 U19105 ( .A(n12422), .B(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n15879) );
  NAND2_X1 U19106 ( .A1(n19170), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n15870) );
  OAI21_X1 U19107 ( .B1(n16559), .B2(n15756), .A(n15870), .ZN(n15757) );
  AOI21_X1 U19108 ( .B1(n16550), .B2(n15758), .A(n15757), .ZN(n15759) );
  OAI21_X1 U19109 ( .B1(n15869), .B2(n16545), .A(n15759), .ZN(n15760) );
  AOI21_X1 U19110 ( .B1(n15879), .B2(n16539), .A(n15760), .ZN(n15761) );
  OAI21_X1 U19111 ( .B1(n15881), .B2(n16553), .A(n15761), .ZN(P2_U2986) );
  XNOR2_X1 U19112 ( .A(n15762), .B(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15893) );
  AOI21_X1 U19113 ( .B1(n15764), .B2(n9864), .A(n15763), .ZN(n15891) );
  NAND2_X1 U19114 ( .A1(n19170), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n15882) );
  OAI21_X1 U19115 ( .B1(n16559), .B2(n15765), .A(n15882), .ZN(n15766) );
  AOI21_X1 U19116 ( .B1(n16550), .B2(n15767), .A(n15766), .ZN(n15768) );
  OAI21_X1 U19117 ( .B1(n15889), .B2(n16545), .A(n15768), .ZN(n15769) );
  AOI21_X1 U19118 ( .B1(n15891), .B2(n16539), .A(n15769), .ZN(n15770) );
  OAI21_X1 U19119 ( .B1(n15893), .B2(n16553), .A(n15770), .ZN(P2_U2987) );
  NOR2_X1 U19120 ( .A1(n15798), .A2(n15912), .ZN(n15785) );
  OAI21_X1 U19121 ( .B1(n15785), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n9864), .ZN(n15904) );
  NAND2_X1 U19122 ( .A1(n15772), .A2(n15781), .ZN(n15774) );
  XNOR2_X1 U19123 ( .A(n15774), .B(n15773), .ZN(n15902) );
  NOR2_X1 U19124 ( .A1(n16452), .A2(n16545), .ZN(n15778) );
  NAND2_X1 U19125 ( .A1(n19170), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n15894) );
  NAND2_X1 U19126 ( .A1(n19313), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15775) );
  OAI211_X1 U19127 ( .C1(n19325), .C2(n15776), .A(n15894), .B(n15775), .ZN(
        n15777) );
  AOI211_X1 U19128 ( .C1(n15902), .C2(n12840), .A(n15778), .B(n15777), .ZN(
        n15779) );
  OAI21_X1 U19129 ( .B1(n15904), .B2(n19319), .A(n15779), .ZN(P2_U2988) );
  INV_X1 U19130 ( .A(n15781), .ZN(n15784) );
  AND2_X1 U19131 ( .A1(n15781), .A2(n15780), .ZN(n15783) );
  OAI22_X1 U19132 ( .A1(n15772), .A2(n15784), .B1(n15783), .B2(n15782), .ZN(
        n15920) );
  INV_X1 U19133 ( .A(n15785), .ZN(n15906) );
  NAND2_X1 U19134 ( .A1(n15798), .A2(n15912), .ZN(n15905) );
  NAND3_X1 U19135 ( .A1(n15906), .A2(n16539), .A3(n15905), .ZN(n15791) );
  NAND2_X1 U19136 ( .A1(n16550), .A2(n15786), .ZN(n15787) );
  NAND2_X1 U19137 ( .A1(n19170), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n15908) );
  OAI211_X1 U19138 ( .C1(n16559), .C2(n15788), .A(n15787), .B(n15908), .ZN(
        n15789) );
  AOI21_X1 U19139 ( .B1(n15917), .B2(n19315), .A(n15789), .ZN(n15790) );
  OAI211_X1 U19140 ( .C1(n16553), .C2(n15920), .A(n15791), .B(n15790), .ZN(
        P2_U2989) );
  NAND2_X1 U19141 ( .A1(n15793), .A2(n15792), .ZN(n15795) );
  XOR2_X1 U19142 ( .A(n15795), .B(n15794), .Z(n15933) );
  BUF_X1 U19143 ( .A(n15796), .Z(n15797) );
  AOI21_X1 U19144 ( .B1(n15922), .B2(n15797), .A(n15771), .ZN(n15921) );
  NAND2_X1 U19145 ( .A1(n15921), .A2(n16539), .ZN(n15804) );
  INV_X1 U19146 ( .A(n15926), .ZN(n15802) );
  NAND2_X1 U19147 ( .A1(n19170), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n15924) );
  NAND2_X1 U19148 ( .A1(n19313), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15799) );
  OAI211_X1 U19149 ( .C1(n19325), .C2(n15800), .A(n15924), .B(n15799), .ZN(
        n15801) );
  AOI21_X1 U19150 ( .B1(n15802), .B2(n19315), .A(n15801), .ZN(n15803) );
  OAI211_X1 U19151 ( .C1(n15933), .C2(n16553), .A(n15804), .B(n15803), .ZN(
        P2_U2990) );
  NAND2_X1 U19152 ( .A1(n16550), .A2(n15805), .ZN(n15807) );
  OAI211_X1 U19153 ( .C1(n16559), .C2(n15808), .A(n15807), .B(n15806), .ZN(
        n15811) );
  NOR2_X1 U19154 ( .A1(n15809), .A2(n19319), .ZN(n15810) );
  AOI211_X1 U19155 ( .C1(n19315), .C2(n15812), .A(n15811), .B(n15810), .ZN(
        n15813) );
  OAI21_X1 U19156 ( .B1(n15814), .B2(n16553), .A(n15813), .ZN(P2_U2993) );
  NOR2_X1 U19157 ( .A1(n15816), .A2(n15815), .ZN(n15821) );
  INV_X1 U19158 ( .A(n15817), .ZN(n15819) );
  NOR2_X1 U19159 ( .A1(n15819), .A2(n15818), .ZN(n15820) );
  XNOR2_X1 U19160 ( .A(n15821), .B(n15820), .ZN(n15973) );
  AOI21_X1 U19161 ( .B1(n15963), .B2(n15822), .A(n11464), .ZN(n15971) );
  INV_X1 U19162 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n19964) );
  NOR2_X1 U19163 ( .A1(n19345), .A2(n19964), .ZN(n15966) );
  NOR2_X1 U19164 ( .A1(n19325), .A2(n15823), .ZN(n15824) );
  AOI211_X1 U19165 ( .C1(n19313), .C2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n15966), .B(n15824), .ZN(n15825) );
  OAI21_X1 U19166 ( .B1(n15968), .B2(n16545), .A(n15825), .ZN(n15826) );
  AOI21_X1 U19167 ( .B1(n15971), .B2(n16539), .A(n15826), .ZN(n15827) );
  OAI21_X1 U19168 ( .B1(n15973), .B2(n16553), .A(n15827), .ZN(P2_U2994) );
  NAND2_X1 U19169 ( .A1(n15828), .A2(n15986), .ZN(n15832) );
  NAND2_X1 U19170 ( .A1(n15830), .A2(n15829), .ZN(n15831) );
  XNOR2_X1 U19171 ( .A(n15832), .B(n15831), .ZN(n15985) );
  NAND2_X1 U19172 ( .A1(n16550), .A2(n19063), .ZN(n15833) );
  NAND2_X1 U19173 ( .A1(n19170), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n15975) );
  OAI211_X1 U19174 ( .C1(n16559), .C2(n19064), .A(n15833), .B(n15975), .ZN(
        n15838) );
  OAI21_X1 U19175 ( .B1(n15834), .B2(n15835), .A(n15980), .ZN(n15836) );
  NAND2_X1 U19176 ( .A1(n15836), .A2(n15822), .ZN(n15974) );
  NOR2_X1 U19177 ( .A1(n15974), .A2(n19319), .ZN(n15837) );
  AOI211_X1 U19178 ( .C1(n19315), .C2(n19070), .A(n15838), .B(n15837), .ZN(
        n15839) );
  OAI21_X1 U19179 ( .B1(n15985), .B2(n16553), .A(n15839), .ZN(P2_U2995) );
  NAND2_X1 U19180 ( .A1(n15841), .A2(n15840), .ZN(n15843) );
  XOR2_X1 U19181 ( .A(n15843), .B(n15842), .Z(n16010) );
  INV_X1 U19182 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n19959) );
  NOR2_X1 U19183 ( .A1(n19959), .A2(n19345), .ZN(n15847) );
  INV_X1 U19184 ( .A(n19076), .ZN(n15844) );
  OAI22_X1 U19185 ( .A1(n16559), .A2(n15845), .B1(n19325), .B2(n15844), .ZN(
        n15846) );
  AOI211_X1 U19186 ( .C1(n19082), .C2(n19315), .A(n15847), .B(n15846), .ZN(
        n15849) );
  OAI211_X1 U19187 ( .C1(n9861), .C2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n16539), .B(n15834), .ZN(n15848) );
  OAI211_X1 U19188 ( .C1(n16010), .C2(n16553), .A(n15849), .B(n15848), .ZN(
        P2_U2997) );
  NAND2_X1 U19189 ( .A1(n15850), .A2(n16040), .ZN(n15851) );
  XNOR2_X1 U19190 ( .A(n12442), .B(n15851), .ZN(n16070) );
  AND2_X1 U19191 ( .A1(n14530), .A2(n16054), .ZN(n16511) );
  INV_X1 U19192 ( .A(n16511), .ZN(n15853) );
  NAND2_X1 U19193 ( .A1(n16511), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n16045) );
  INV_X1 U19194 ( .A(n16045), .ZN(n15852) );
  AOI21_X1 U19195 ( .B1(n16062), .B2(n15853), .A(n15852), .ZN(n16066) );
  INV_X1 U19196 ( .A(n15854), .ZN(n19109) );
  OAI22_X1 U19197 ( .A1(n16559), .A2(n19111), .B1(n19325), .B2(n19109), .ZN(
        n15857) );
  INV_X1 U19198 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n15855) );
  OAI22_X1 U19199 ( .A1(n16545), .A2(n19115), .B1(n15855), .B2(n19345), .ZN(
        n15856) );
  AOI211_X1 U19200 ( .C1(n16066), .C2(n16539), .A(n15857), .B(n15856), .ZN(
        n15858) );
  OAI21_X1 U19201 ( .B1(n16553), .B2(n16070), .A(n15858), .ZN(P2_U3001) );
  NOR2_X1 U19202 ( .A1(n16087), .A2(n16088), .ZN(n16086) );
  NAND2_X1 U19203 ( .A1(n15859), .A2(n16071), .ZN(n16512) );
  OAI21_X1 U19204 ( .B1(n16086), .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n16512), .ZN(n16085) );
  INV_X1 U19205 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n15860) );
  NOR2_X1 U19206 ( .A1(n19345), .A2(n15860), .ZN(n16078) );
  INV_X1 U19207 ( .A(n19126), .ZN(n15861) );
  OAI22_X1 U19208 ( .A1(n16559), .A2(n15862), .B1(n19325), .B2(n15861), .ZN(
        n15863) );
  AOI211_X1 U19209 ( .C1(n19315), .C2(n19127), .A(n16078), .B(n15863), .ZN(
        n15868) );
  XNOR2_X1 U19210 ( .A(n15865), .B(n16080), .ZN(n15866) );
  XNOR2_X1 U19211 ( .A(n15864), .B(n15866), .ZN(n16083) );
  NAND2_X1 U19212 ( .A1(n16083), .A2(n12840), .ZN(n15867) );
  OAI211_X1 U19213 ( .C1(n16085), .C2(n19319), .A(n15868), .B(n15867), .ZN(
        P2_U3003) );
  INV_X1 U19214 ( .A(n15869), .ZN(n15873) );
  OAI21_X1 U19215 ( .B1(n19327), .B2(n15871), .A(n15870), .ZN(n15872) );
  NAND2_X1 U19216 ( .A1(n15874), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n15875) );
  OAI211_X1 U19217 ( .C1(n15877), .C2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n15876), .B(n15875), .ZN(n15878) );
  AOI21_X1 U19218 ( .B1(n15879), .B2(n16577), .A(n15878), .ZN(n15880) );
  OAI21_X1 U19219 ( .B1(n15881), .B2(n19363), .A(n15880), .ZN(P2_U3018) );
  OAI211_X1 U19220 ( .C1(n19327), .C2(n15884), .A(n15883), .B(n15882), .ZN(
        n15885) );
  INV_X1 U19221 ( .A(n15885), .ZN(n15888) );
  NAND3_X1 U19222 ( .A1(n15886), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A3(
        n15911), .ZN(n15887) );
  OAI211_X1 U19223 ( .C1(n15889), .C2(n19355), .A(n15888), .B(n15887), .ZN(
        n15890) );
  AOI21_X1 U19224 ( .B1(n15891), .B2(n16577), .A(n15890), .ZN(n15892) );
  OAI21_X1 U19225 ( .B1(n15893), .B2(n19363), .A(n15892), .ZN(P2_U3019) );
  INV_X1 U19226 ( .A(n15894), .ZN(n15898) );
  INV_X1 U19227 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15896) );
  AOI211_X1 U19228 ( .C1(n15896), .C2(n15912), .A(n15895), .B(n15910), .ZN(
        n15897) );
  AOI211_X1 U19229 ( .C1(n19347), .C2(n16455), .A(n15898), .B(n15897), .ZN(
        n15900) );
  NAND3_X1 U19230 ( .A1(n15930), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        n15911), .ZN(n15899) );
  OAI211_X1 U19231 ( .C1(n16452), .C2(n19355), .A(n15900), .B(n15899), .ZN(
        n15901) );
  AOI21_X1 U19232 ( .B1(n15902), .B2(n19331), .A(n15901), .ZN(n15903) );
  OAI21_X1 U19233 ( .B1(n15904), .B2(n19356), .A(n15903), .ZN(P2_U3020) );
  NAND3_X1 U19234 ( .A1(n15906), .A2(n16577), .A3(n15905), .ZN(n15919) );
  NAND2_X1 U19235 ( .A1(n19347), .A2(n15907), .ZN(n15909) );
  OAI211_X1 U19236 ( .C1(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .C2(n15910), .A(
        n15909), .B(n15908), .ZN(n15916) );
  INV_X1 U19237 ( .A(n15911), .ZN(n15913) );
  NOR3_X1 U19238 ( .A1(n15914), .A2(n15913), .A3(n15912), .ZN(n15915) );
  AOI211_X1 U19239 ( .C1(n15917), .C2(n19341), .A(n15916), .B(n15915), .ZN(
        n15918) );
  OAI211_X1 U19240 ( .C1(n15920), .C2(n19363), .A(n15919), .B(n15918), .ZN(
        P2_U3021) );
  NAND2_X1 U19241 ( .A1(n15921), .A2(n16577), .ZN(n15932) );
  INV_X1 U19242 ( .A(n15937), .ZN(n15923) );
  OAI21_X1 U19243 ( .B1(n15955), .B2(n15923), .A(n15922), .ZN(n15929) );
  OAI21_X1 U19244 ( .B1(n19327), .B2(n15925), .A(n15924), .ZN(n15928) );
  NOR2_X1 U19245 ( .A1(n15926), .A2(n19355), .ZN(n15927) );
  AOI211_X1 U19246 ( .C1(n15930), .C2(n15929), .A(n15928), .B(n15927), .ZN(
        n15931) );
  OAI211_X1 U19247 ( .C1(n15933), .C2(n19363), .A(n15932), .B(n15931), .ZN(
        P2_U3022) );
  OAI21_X1 U19248 ( .B1(n15934), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n15797), .ZN(n16474) );
  XNOR2_X1 U19249 ( .A(n15935), .B(n15936), .ZN(n16473) );
  NOR2_X1 U19250 ( .A1(n19970), .A2(n19345), .ZN(n15940) );
  AOI211_X1 U19251 ( .C1(n21278), .C2(n15938), .A(n15937), .B(n15955), .ZN(
        n15939) );
  NOR2_X1 U19252 ( .A1(n15940), .A2(n15939), .ZN(n15941) );
  OAI21_X1 U19253 ( .B1(n19327), .B2(n15942), .A(n15941), .ZN(n15943) );
  AOI21_X1 U19254 ( .B1(n16476), .B2(n19341), .A(n15943), .ZN(n15945) );
  NAND2_X1 U19255 ( .A1(n15953), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15944) );
  OAI211_X1 U19256 ( .C1(n16473), .C2(n19363), .A(n15945), .B(n15944), .ZN(
        n15946) );
  INV_X1 U19257 ( .A(n15946), .ZN(n15947) );
  OAI21_X1 U19258 ( .B1(n16474), .B2(n19356), .A(n15947), .ZN(P2_U3023) );
  INV_X1 U19259 ( .A(n15934), .ZN(n15948) );
  NAND2_X1 U19260 ( .A1(n15951), .A2(n15950), .ZN(n15952) );
  XNOR2_X1 U19261 ( .A(n15949), .B(n15952), .ZN(n16482) );
  NAND2_X1 U19262 ( .A1(n15953), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15958) );
  NAND2_X1 U19263 ( .A1(P2_REIP_REG_22__SCAN_IN), .A2(n19170), .ZN(n15954) );
  OAI21_X1 U19264 ( .B1(n15955), .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n15954), .ZN(n15956) );
  AOI21_X1 U19265 ( .B1(n19347), .B2(n16457), .A(n15956), .ZN(n15957) );
  OAI211_X1 U19266 ( .C1(n15959), .C2(n19355), .A(n15958), .B(n15957), .ZN(
        n15960) );
  AOI21_X1 U19267 ( .B1(n16482), .B2(n19331), .A(n15960), .ZN(n15961) );
  OAI21_X1 U19268 ( .B1(n16480), .B2(n19356), .A(n15961), .ZN(P2_U3024) );
  NAND2_X1 U19269 ( .A1(n16073), .A2(n16004), .ZN(n16001) );
  NOR2_X1 U19270 ( .A1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n16001), .ZN(
        n15991) );
  OAI21_X1 U19271 ( .B1(n15962), .B2(n19353), .A(n16047), .ZN(n15993) );
  NOR2_X1 U19272 ( .A1(n15991), .A2(n15993), .ZN(n15981) );
  NOR2_X1 U19273 ( .A1(n15981), .A2(n15963), .ZN(n15970) );
  XNOR2_X1 U19274 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .B(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15964) );
  NOR2_X1 U19275 ( .A1(n15964), .A2(n15976), .ZN(n15965) );
  AOI211_X1 U19276 ( .C1(n19347), .C2(n9921), .A(n15966), .B(n15965), .ZN(
        n15967) );
  OAI21_X1 U19277 ( .B1(n15968), .B2(n19355), .A(n15967), .ZN(n15969) );
  AOI211_X1 U19278 ( .C1(n15971), .C2(n16577), .A(n15970), .B(n15969), .ZN(
        n15972) );
  OAI21_X1 U19279 ( .B1(n15973), .B2(n19363), .A(n15972), .ZN(P2_U3026) );
  INV_X1 U19280 ( .A(n15974), .ZN(n15983) );
  NOR2_X1 U19281 ( .A1(n19327), .A2(n19068), .ZN(n15978) );
  OAI21_X1 U19282 ( .B1(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n15976), .A(
        n15975), .ZN(n15977) );
  AOI211_X1 U19283 ( .C1(n19070), .C2(n19341), .A(n15978), .B(n15977), .ZN(
        n15979) );
  OAI21_X1 U19284 ( .B1(n15981), .B2(n15980), .A(n15979), .ZN(n15982) );
  AOI21_X1 U19285 ( .B1(n15983), .B2(n16577), .A(n15982), .ZN(n15984) );
  OAI21_X1 U19286 ( .B1(n15985), .B2(n19363), .A(n15984), .ZN(P2_U3027) );
  NAND2_X1 U19287 ( .A1(n15987), .A2(n15986), .ZN(n15989) );
  XOR2_X1 U19288 ( .A(n15989), .B(n15988), .Z(n16487) );
  NAND2_X1 U19289 ( .A1(n16487), .A2(n19331), .ZN(n15999) );
  NOR3_X1 U19290 ( .A1(n16034), .A2(n16491), .A3(n15990), .ZN(n15992) );
  AOI22_X1 U19291 ( .A1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n15993), .B1(
        n15992), .B2(n15991), .ZN(n15998) );
  OAI22_X1 U19292 ( .A1(n19327), .A2(n16466), .B1(n15994), .B2(n19345), .ZN(
        n15995) );
  AOI21_X1 U19293 ( .B1(n16486), .B2(n19341), .A(n15995), .ZN(n15997) );
  XNOR2_X1 U19294 ( .A(n15834), .B(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n16485) );
  NAND2_X1 U19295 ( .A1(n16485), .A2(n16577), .ZN(n15996) );
  NAND4_X1 U19296 ( .A1(n15999), .A2(n15998), .A3(n15997), .A4(n15996), .ZN(
        P2_U3028) );
  OAI22_X1 U19297 ( .A1(n19327), .A2(n19080), .B1(n19959), .B2(n19345), .ZN(
        n16003) );
  INV_X1 U19298 ( .A(n16001), .ZN(n16035) );
  AOI22_X1 U19299 ( .A1(n16020), .A2(n16577), .B1(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n16035), .ZN(n16012) );
  NOR3_X1 U19300 ( .A1(n16012), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A3(
        n16491), .ZN(n16002) );
  AOI211_X1 U19301 ( .C1(n19082), .C2(n19341), .A(n16003), .B(n16002), .ZN(
        n16009) );
  INV_X1 U19302 ( .A(n19333), .ZN(n19334) );
  OR2_X1 U19303 ( .A1(n19353), .A2(n16004), .ZN(n16005) );
  NAND2_X1 U19304 ( .A1(n16047), .A2(n16005), .ZN(n16026) );
  AOI21_X1 U19305 ( .B1(n19356), .B2(n19336), .A(n9861), .ZN(n16006) );
  AOI211_X1 U19306 ( .C1(n19334), .C2(n16034), .A(n16026), .B(n16006), .ZN(
        n16018) );
  OAI21_X1 U19307 ( .B1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n19353), .A(
        n16018), .ZN(n16007) );
  NAND2_X1 U19308 ( .A1(n16007), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n16008) );
  OAI211_X1 U19309 ( .C1(n16010), .C2(n19363), .A(n16009), .B(n16008), .ZN(
        P2_U3029) );
  INV_X1 U19310 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n16011) );
  OAI22_X1 U19311 ( .A1(n19355), .A2(n16493), .B1(n16011), .B2(n19345), .ZN(
        n16014) );
  NOR2_X1 U19312 ( .A1(n16012), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n16013) );
  AOI211_X1 U19313 ( .C1(n19347), .C2(n19224), .A(n16014), .B(n16013), .ZN(
        n16017) );
  XNOR2_X1 U19314 ( .A(n9898), .B(n16015), .ZN(n16496) );
  NAND2_X1 U19315 ( .A1(n16496), .A2(n19331), .ZN(n16016) );
  OAI211_X1 U19316 ( .C1(n16018), .C2(n16491), .A(n16017), .B(n16016), .ZN(
        P2_U3030) );
  AND2_X1 U19317 ( .A1(n16019), .A2(n16034), .ZN(n16021) );
  OR2_X1 U19318 ( .A1(n16021), .A2(n16020), .ZN(n16500) );
  OAI21_X1 U19319 ( .B1(n16023), .B2(n16025), .A(n16022), .ZN(n16024) );
  OAI21_X1 U19320 ( .B1(n9906), .B2(n16025), .A(n16024), .ZN(n16501) );
  OR2_X1 U19321 ( .A1(n16501), .A2(n19363), .ZN(n16037) );
  NAND2_X1 U19322 ( .A1(n16026), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n16032) );
  INV_X1 U19323 ( .A(n14442), .ZN(n16027) );
  OAI21_X1 U19324 ( .B1(n16028), .B2(n9865), .A(n16027), .ZN(n19231) );
  INV_X1 U19325 ( .A(n19231), .ZN(n16030) );
  INV_X1 U19326 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n19956) );
  NOR2_X1 U19327 ( .A1(n19956), .A2(n19345), .ZN(n16029) );
  AOI21_X1 U19328 ( .B1(n19347), .B2(n16030), .A(n16029), .ZN(n16031) );
  OAI211_X1 U19329 ( .C1(n19355), .C2(n19091), .A(n16032), .B(n16031), .ZN(
        n16033) );
  AOI21_X1 U19330 ( .B1(n16035), .B2(n16034), .A(n16033), .ZN(n16036) );
  OAI211_X1 U19331 ( .C1(n16500), .C2(n19356), .A(n16037), .B(n16036), .ZN(
        P2_U3031) );
  NAND2_X1 U19332 ( .A1(n16039), .A2(n16038), .ZN(n16043) );
  NAND2_X1 U19333 ( .A1(n16041), .A2(n16040), .ZN(n16042) );
  XOR2_X1 U19334 ( .A(n16043), .B(n16042), .Z(n16508) );
  INV_X1 U19335 ( .A(n16508), .ZN(n16059) );
  INV_X1 U19336 ( .A(n16019), .ZN(n16044) );
  AOI21_X1 U19337 ( .B1(n16045), .B2(n16049), .A(n16044), .ZN(n16507) );
  NAND3_X1 U19338 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n16071), .A3(
        n16073), .ZN(n16046) );
  NOR2_X1 U19339 ( .A1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n16046), .ZN(
        n16563) );
  INV_X1 U19340 ( .A(n16047), .ZN(n16560) );
  AOI211_X1 U19341 ( .C1(n16562), .C2(n16561), .A(n16563), .B(n16560), .ZN(
        n16063) );
  NAND4_X1 U19342 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n16071), .A3(
        n16073), .A4(n16062), .ZN(n16061) );
  NAND2_X1 U19343 ( .A1(P2_REIP_REG_14__SCAN_IN), .A2(n19170), .ZN(n16048) );
  OAI221_X1 U19344 ( .B1(n16049), .B2(n16063), .C1(n16049), .C2(n16061), .A(
        n16048), .ZN(n16057) );
  AOI21_X1 U19345 ( .B1(n16051), .B2(n16050), .A(n9865), .ZN(n19103) );
  INV_X1 U19346 ( .A(n19103), .ZN(n19234) );
  NOR3_X1 U19347 ( .A1(n16062), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A3(
        n16052), .ZN(n16053) );
  AOI22_X1 U19348 ( .A1(n19341), .A2(n19102), .B1(n16054), .B2(n16053), .ZN(
        n16055) );
  OAI21_X1 U19349 ( .B1(n19234), .B2(n19327), .A(n16055), .ZN(n16056) );
  AOI211_X1 U19350 ( .C1(n16507), .C2(n16577), .A(n16057), .B(n16056), .ZN(
        n16058) );
  OAI21_X1 U19351 ( .B1(n16059), .B2(n19363), .A(n16058), .ZN(P2_U3032) );
  XOR2_X1 U19352 ( .A(n15619), .B(n16060), .Z(n19235) );
  OAI22_X1 U19353 ( .A1(n16063), .A2(n16062), .B1(n16570), .B2(n16061), .ZN(
        n16065) );
  OAI22_X1 U19354 ( .A1(n19355), .A2(n19115), .B1(n15855), .B2(n19345), .ZN(
        n16064) );
  OR2_X1 U19355 ( .A1(n16065), .A2(n16064), .ZN(n16068) );
  AND2_X1 U19356 ( .A1(n16066), .A2(n16577), .ZN(n16067) );
  AOI211_X1 U19357 ( .C1(n19347), .C2(n19235), .A(n16068), .B(n16067), .ZN(
        n16069) );
  OAI21_X1 U19358 ( .B1(n19363), .B2(n16070), .A(n16069), .ZN(P2_U3033) );
  NAND2_X1 U19359 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n16073), .ZN(
        n16099) );
  AOI211_X1 U19360 ( .C1(n16088), .C2(n16080), .A(n16071), .B(n16099), .ZN(
        n16082) );
  AOI21_X1 U19361 ( .B1(n16073), .B2(n16072), .A(n16560), .ZN(n16098) );
  OAI21_X1 U19362 ( .B1(n16076), .B2(n16075), .A(n16074), .ZN(n19243) );
  NOR2_X1 U19363 ( .A1(n19327), .A2(n19243), .ZN(n16077) );
  AOI211_X1 U19364 ( .C1(n19341), .C2(n19127), .A(n16078), .B(n16077), .ZN(
        n16079) );
  OAI21_X1 U19365 ( .B1(n16098), .B2(n16080), .A(n16079), .ZN(n16081) );
  AOI211_X1 U19366 ( .C1(n16083), .C2(n19331), .A(n16082), .B(n16081), .ZN(
        n16084) );
  OAI21_X1 U19367 ( .B1(n16085), .B2(n19356), .A(n16084), .ZN(P2_U3035) );
  AOI21_X1 U19368 ( .B1(n16088), .B2(n16087), .A(n16086), .ZN(n16518) );
  NAND2_X1 U19369 ( .A1(n16518), .A2(n16577), .ZN(n16104) );
  AOI22_X1 U19370 ( .A1(n19341), .A2(n16519), .B1(n19347), .B2(n19245), .ZN(
        n16103) );
  INV_X1 U19371 ( .A(n16089), .ZN(n16091) );
  OAI21_X1 U19372 ( .B1(n16092), .B2(n16091), .A(n16090), .ZN(n16096) );
  NAND2_X1 U19373 ( .A1(n16094), .A2(n16093), .ZN(n16095) );
  XNOR2_X1 U19374 ( .A(n16096), .B(n16095), .ZN(n16520) );
  NAND2_X1 U19375 ( .A1(n16520), .A2(n19331), .ZN(n16102) );
  NAND2_X1 U19376 ( .A1(P2_REIP_REG_10__SCAN_IN), .A2(n19170), .ZN(n16097) );
  OAI221_X1 U19377 ( .B1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n16099), 
        .C1(n16088), .C2(n16098), .A(n16097), .ZN(n16100) );
  INV_X1 U19378 ( .A(n16100), .ZN(n16101) );
  NAND4_X1 U19379 ( .A1(n16104), .A2(n16103), .A3(n16102), .A4(n16101), .ZN(
        P2_U3036) );
  AOI221_X1 U19380 ( .B1(n19215), .B2(n10135), .C1(n16105), .C2(n19159), .A(
        n13362), .ZN(n16121) );
  INV_X1 U19381 ( .A(n16121), .ZN(n16110) );
  OAI21_X1 U19382 ( .B1(n16106), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n13362), 
        .ZN(n16109) );
  INV_X1 U19383 ( .A(n16107), .ZN(n16108) );
  AOI22_X1 U19384 ( .A1(n16110), .A2(n16109), .B1(n16108), .B2(n16589), .ZN(
        n16112) );
  NAND2_X1 U19385 ( .A1(n16118), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n16111) );
  OAI21_X1 U19386 ( .B1(n16112), .B2(n16118), .A(n16111), .ZN(P2_U3601) );
  OAI21_X1 U19387 ( .B1(n19215), .B2(n16114), .A(n16113), .ZN(n19196) );
  OAI21_X1 U19388 ( .B1(n10135), .B2(n19348), .A(n19196), .ZN(n16122) );
  INV_X1 U19389 ( .A(n16122), .ZN(n16115) );
  AOI222_X1 U19390 ( .A1(n16116), .A2(n20005), .B1(n16589), .B2(n20029), .C1(
        n16115), .C2(n16121), .ZN(n16119) );
  NAND2_X1 U19391 ( .A1(n16118), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n16117) );
  OAI21_X1 U19392 ( .B1(n16119), .B2(n16118), .A(n16117), .ZN(P2_U3600) );
  INV_X1 U19393 ( .A(n16120), .ZN(n16123) );
  AOI222_X1 U19394 ( .A1(n16123), .A2(n20005), .B1(n16122), .B2(n16121), .C1(
        n16589), .C2(n19364), .ZN(n16124) );
  MUX2_X1 U19395 ( .A(n10144), .B(n16124), .S(n16160), .Z(n16126) );
  INV_X1 U19396 ( .A(n16126), .ZN(P2_U3599) );
  AOI22_X1 U19397 ( .A1(n13120), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17343), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n16127) );
  OAI21_X1 U19398 ( .B1(n13051), .B2(n17200), .A(n16127), .ZN(n16136) );
  AOI22_X1 U19399 ( .A1(n12552), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n13089), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n16134) );
  AOI22_X1 U19400 ( .A1(n13080), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17361), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n16128) );
  OAI21_X1 U19401 ( .B1(n17363), .B2(n17201), .A(n16128), .ZN(n16132) );
  AOI22_X1 U19402 ( .A1(n17379), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17245), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n16130) );
  AOI22_X1 U19403 ( .A1(n17385), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n17365), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n16129) );
  OAI211_X1 U19404 ( .C1(n12551), .C2(n17407), .A(n16130), .B(n16129), .ZN(
        n16131) );
  AOI211_X1 U19405 ( .C1(n17327), .C2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A(
        n16132), .B(n16131), .ZN(n16133) );
  OAI211_X1 U19406 ( .C1(n12561), .C2(n17211), .A(n16134), .B(n16133), .ZN(
        n16135) );
  AOI211_X1 U19407 ( .C1(n17357), .C2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A(
        n16136), .B(n16135), .ZN(n17525) );
  INV_X1 U19408 ( .A(n16137), .ZN(n17321) );
  AOI21_X1 U19409 ( .B1(P3_EBX_REG_13__SCAN_IN), .B2(n17418), .A(n17321), .ZN(
        n16138) );
  OAI22_X1 U19410 ( .A1(n17525), .A2(n17418), .B1(n17301), .B2(n16138), .ZN(
        P3_U2690) );
  NOR2_X1 U19411 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18967), .ZN(
        n18423) );
  NAND3_X1 U19412 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_0__SCAN_IN), .A3(P3_STATE2_REG_2__SCAN_IN), .ZN(n18965)
         );
  INV_X1 U19413 ( .A(n18965), .ZN(n18875) );
  INV_X1 U19414 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n18812) );
  NAND3_X1 U19415 ( .A1(n17395), .A2(n16153), .A3(n18812), .ZN(n18368) );
  INV_X1 U19416 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n18369) );
  NOR2_X1 U19417 ( .A1(n18369), .A2(n18965), .ZN(n16151) );
  AOI211_X1 U19418 ( .C1(n18875), .C2(n18368), .A(n18720), .B(n16151), .ZN(
        n16139) );
  NOR2_X1 U19419 ( .A1(n18423), .A2(n16139), .ZN(n16141) );
  INV_X1 U19420 ( .A(n16145), .ZN(n18717) );
  INV_X1 U19421 ( .A(n16139), .ZN(n18374) );
  INV_X1 U19422 ( .A(n18006), .ZN(n17890) );
  OAI22_X1 U19423 ( .A1(n17890), .A2(n19019), .B1(n18621), .B2(n18967), .ZN(
        n16144) );
  NAND3_X1 U19424 ( .A1(n18620), .A2(n18374), .A3(n16144), .ZN(n16140) );
  OAI221_X1 U19425 ( .B1(n18620), .B2(n16141), .C1(n18620), .C2(n18717), .A(
        n16140), .ZN(P3_U2864) );
  NAND2_X1 U19426 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18531) );
  NOR2_X1 U19427 ( .A1(n17890), .A2(n19019), .ZN(n16143) );
  INV_X1 U19428 ( .A(n16141), .ZN(n16142) );
  AOI221_X1 U19429 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n18531), .C1(n16143), 
        .C2(n18531), .A(n16142), .ZN(n18373) );
  OAI221_X1 U19430 ( .B1(n16145), .B2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .C1(n16145), .C2(n16144), .A(n18374), .ZN(n18371) );
  AOI22_X1 U19431 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18373), .B1(
        n18371), .B2(n18845), .ZN(P3_U2865) );
  NAND2_X1 U19432 ( .A1(n19012), .A2(n17632), .ZN(n18857) );
  OAI211_X1 U19433 ( .C1(n17582), .C2(n16229), .A(n16230), .B(n18858), .ZN(
        n16147) );
  OAI211_X1 U19434 ( .C1(n16150), .C2(n16149), .A(n16148), .B(n16147), .ZN(
        n18842) );
  NOR2_X1 U19435 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18967), .ZN(n18375) );
  INV_X1 U19436 ( .A(n18998), .ZN(n18996) );
  AOI21_X1 U19437 ( .B1(n16153), .B2(n18812), .A(n16152), .ZN(n18854) );
  NAND3_X1 U19438 ( .A1(n18996), .A2(n19028), .A3(n18854), .ZN(n16154) );
  OAI21_X1 U19439 ( .B1(n18996), .B2(n18812), .A(n16154), .ZN(P3_U3284) );
  AND4_X1 U19440 ( .A1(n16157), .A2(n16156), .A3(n20005), .A4(n16155), .ZN(
        n16158) );
  NAND2_X1 U19441 ( .A1(n16160), .A2(n16158), .ZN(n16159) );
  OAI21_X1 U19442 ( .B1(n16160), .B2(n11383), .A(n16159), .ZN(P2_U3595) );
  OAI21_X1 U19443 ( .B1(n18222), .B2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n16161), .ZN(n16630) );
  INV_X1 U19444 ( .A(n18288), .ZN(n18089) );
  OAI22_X1 U19445 ( .A1(n16608), .A2(n18089), .B1(n16609), .B2(n18326), .ZN(
        n16162) );
  NOR2_X1 U19446 ( .A1(n18344), .A2(n16162), .ZN(n16220) );
  OAI21_X1 U19447 ( .B1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n18351), .A(
        n16220), .ZN(n16163) );
  AOI21_X1 U19448 ( .B1(n18359), .B2(n16630), .A(n16163), .ZN(n16170) );
  NOR2_X1 U19449 ( .A1(n16165), .A2(n16164), .ZN(n16166) );
  XNOR2_X1 U19450 ( .A(n16166), .B(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16613) );
  OR2_X1 U19451 ( .A1(n16625), .A2(n18089), .ZN(n16167) );
  OAI211_X1 U19452 ( .C1(n18326), .C2(n16631), .A(n16168), .B(n16167), .ZN(
        n16215) );
  AOI22_X1 U19453 ( .A1(n18287), .A2(n16613), .B1(n16610), .B2(n16215), .ZN(
        n16169) );
  NAND2_X1 U19454 ( .A1(n18096), .A2(P3_REIP_REG_29__SCAN_IN), .ZN(n16620) );
  OAI211_X1 U19455 ( .C1(n16170), .C2(n16610), .A(n16169), .B(n16620), .ZN(
        P3_U2833) );
  INV_X1 U19456 ( .A(n16171), .ZN(n16173) );
  NAND2_X1 U19457 ( .A1(n16173), .A2(n16172), .ZN(n16179) );
  AOI21_X1 U19458 ( .B1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n16175), .A(
        n16174), .ZN(n16176) );
  AOI22_X1 U19459 ( .A1(n16179), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B1(
        n16176), .B2(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n16177) );
  INV_X1 U19460 ( .A(n16177), .ZN(n16178) );
  OAI21_X1 U19461 ( .B1(n16179), .B2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(
        n16178), .ZN(n16180) );
  AOI222_X1 U19462 ( .A1(n20598), .A2(n16181), .B1(n20598), .B2(n16180), .C1(
        n16181), .C2(n16180), .ZN(n16184) );
  INV_X1 U19463 ( .A(n16182), .ZN(n16183) );
  AOI222_X1 U19464 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n16184), 
        .B1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n16183), .C1(n16184), 
        .C2(n16183), .ZN(n16187) );
  AOI211_X1 U19465 ( .C1(n16187), .C2(n20302), .A(n16186), .B(n16185), .ZN(
        n16200) );
  NOR2_X1 U19466 ( .A1(n16188), .A2(n16210), .ZN(n16191) );
  AOI21_X1 U19467 ( .B1(n16189), .B2(n12754), .A(n16193), .ZN(n16190) );
  AOI211_X1 U19468 ( .C1(n11634), .C2(n16192), .A(n16191), .B(n16190), .ZN(
        n21397) );
  OAI22_X1 U19469 ( .A1(n16194), .A2(n12753), .B1(n12763), .B2(n16193), .ZN(
        n20081) );
  NAND3_X1 U19470 ( .A1(n16196), .A2(n16223), .A3(n16195), .ZN(n16197) );
  AND2_X1 U19471 ( .A1(n16197), .A2(n21010), .ZN(n21007) );
  NOR2_X1 U19472 ( .A1(n20081), .A2(n21007), .ZN(n20087) );
  OAI21_X1 U19473 ( .B1(P1_FLUSH_REG_SCAN_IN), .B2(P1_MORE_REG_SCAN_IN), .A(
        n20087), .ZN(n16198) );
  NAND4_X1 U19474 ( .A1(n16200), .A2(n21397), .A3(n16199), .A4(n16198), .ZN(
        n16206) );
  NOR3_X1 U19475 ( .A1(n12754), .A2(n16201), .A3(n16223), .ZN(n16202) );
  NAND2_X1 U19476 ( .A1(n16203), .A2(n16202), .ZN(n16204) );
  OAI221_X1 U19477 ( .B1(n16207), .B2(n16205), .C1(n16207), .C2(n20919), .A(
        n16204), .ZN(n16440) );
  AOI221_X1 U19478 ( .B1(n20310), .B2(n16442), .C1(n16206), .C2(n16442), .A(
        n16440), .ZN(n16208) );
  NOR2_X1 U19479 ( .A1(n16208), .A2(n20310), .ZN(n20912) );
  OAI211_X1 U19480 ( .C1(P1_STATE2_REG_2__SCAN_IN), .C2(n21010), .A(n20912), 
        .B(n16211), .ZN(n16441) );
  AOI21_X1 U19481 ( .B1(n16207), .B2(n16206), .A(n16441), .ZN(n16214) );
  INV_X1 U19482 ( .A(n16208), .ZN(n16209) );
  OAI21_X1 U19483 ( .B1(n16211), .B2(n16210), .A(n16209), .ZN(n16212) );
  AOI22_X1 U19484 ( .A1(n16214), .A2(n16213), .B1(n20310), .B2(n16212), .ZN(
        P1_U3161) );
  AOI21_X1 U19485 ( .B1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n16215), .A(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n16222) );
  NAND2_X1 U19486 ( .A1(n16217), .A2(n16216), .ZN(n16218) );
  XNOR2_X1 U19487 ( .A(n16218), .B(n16603), .ZN(n16601) );
  AOI22_X1 U19488 ( .A1(n18096), .A2(P3_REIP_REG_30__SCAN_IN), .B1(n18287), 
        .B2(n16601), .ZN(n16219) );
  OAI221_X1 U19489 ( .B1(n16222), .B2(n16221), .C1(n16222), .C2(n16220), .A(
        n16219), .ZN(P3_U2832) );
  INV_X1 U19490 ( .A(HOLD), .ZN(n20920) );
  NOR2_X1 U19491 ( .A1(n20928), .A2(n20920), .ZN(n20915) );
  AOI22_X1 U19492 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(HOLD), .B1(
        P1_STATE_REG_0__SCAN_IN), .B2(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n16224) );
  INV_X1 U19493 ( .A(P1_STATE_REG_1__SCAN_IN), .ZN(n20077) );
  NOR2_X1 U19494 ( .A1(n20077), .A2(n21010), .ZN(n20921) );
  INV_X1 U19495 ( .A(n20921), .ZN(n20913) );
  OAI211_X1 U19496 ( .C1(n20915), .C2(n16224), .A(n16223), .B(n20913), .ZN(
        P1_U3195) );
  AND2_X1 U19497 ( .A1(n20204), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(P1_U2905)
         );
  INV_X1 U19498 ( .A(n16225), .ZN(n20067) );
  NOR3_X1 U19499 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(P2_STATEBS16_REG_SCAN_IN), .ZN(n16227) );
  NOR2_X1 U19500 ( .A1(n20069), .A2(n19037), .ZN(n16586) );
  NOR4_X1 U19501 ( .A1(n20067), .A2(n16227), .A3(n16586), .A4(n16226), .ZN(
        P2_U3178) );
  OAI221_X1 U19502 ( .B1(n11393), .B2(n16595), .C1(n20047), .C2(n16595), .A(
        n19610), .ZN(n20041) );
  NOR2_X1 U19503 ( .A1(n16228), .A2(n20041), .ZN(P2_U3047) );
  NAND2_X1 U19504 ( .A1(n17547), .A2(n17432), .ZN(n17473) );
  INV_X1 U19505 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n17630) );
  NAND2_X1 U19506 ( .A1(n16233), .A2(n17432), .ZN(n17567) );
  AOI22_X1 U19507 ( .A1(n17578), .A2(BUF2_REG_0__SCAN_IN), .B1(n17569), .B2(
        n16235), .ZN(n16236) );
  OAI221_X1 U19508 ( .B1(P3_EAX_REG_0__SCAN_IN), .B2(n17473), .C1(n17630), 
        .C2(n17432), .A(n16236), .ZN(P3_U2735) );
  INV_X1 U19509 ( .A(P1_REIP_REG_19__SCAN_IN), .ZN(n20957) );
  NAND2_X1 U19510 ( .A1(n16238), .A2(n16237), .ZN(n16249) );
  AOI221_X1 U19511 ( .B1(P1_REIP_REG_19__SCAN_IN), .B2(P1_REIP_REG_18__SCAN_IN), .C1(n20957), .C2(n20955), .A(n16249), .ZN(n16239) );
  AOI211_X1 U19512 ( .C1(n20140), .C2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n16239), .B(n20280), .ZN(n16243) );
  INV_X1 U19513 ( .A(n16240), .ZN(n16241) );
  AOI22_X1 U19514 ( .A1(n20154), .A2(n16241), .B1(n20147), .B2(
        P1_EBX_REG_19__SCAN_IN), .ZN(n16242) );
  AND2_X1 U19515 ( .A1(n16243), .A2(n16242), .ZN(n16245) );
  AOI22_X1 U19516 ( .A1(n16296), .A2(n20131), .B1(P1_REIP_REG_19__SCAN_IN), 
        .B2(n16251), .ZN(n16244) );
  OAI211_X1 U19517 ( .C1(n20124), .C2(n16246), .A(n16245), .B(n16244), .ZN(
        P1_U2821) );
  AOI22_X1 U19518 ( .A1(n20154), .A2(n16247), .B1(n20147), .B2(
        P1_EBX_REG_18__SCAN_IN), .ZN(n16248) );
  OAI21_X1 U19519 ( .B1(P1_REIP_REG_18__SCAN_IN), .B2(n16249), .A(n16248), 
        .ZN(n16250) );
  AOI211_X1 U19520 ( .C1(n20140), .C2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n20280), .B(n16250), .ZN(n16254) );
  AOI22_X1 U19521 ( .A1(n16252), .A2(n20131), .B1(P1_REIP_REG_18__SCAN_IN), 
        .B2(n16251), .ZN(n16253) );
  OAI211_X1 U19522 ( .C1(n20124), .C2(n16255), .A(n16254), .B(n16253), .ZN(
        P1_U2822) );
  INV_X1 U19523 ( .A(n16256), .ZN(n16363) );
  AOI22_X1 U19524 ( .A1(n16363), .A2(n20149), .B1(n20147), .B2(
        P1_EBX_REG_15__SCAN_IN), .ZN(n16257) );
  OAI211_X1 U19525 ( .C1(n20158), .C2(n16258), .A(n16257), .B(n20256), .ZN(
        n16259) );
  AOI21_X1 U19526 ( .B1(n16317), .B2(n20154), .A(n16259), .ZN(n16262) );
  AOI22_X1 U19527 ( .A1(n16318), .A2(n20131), .B1(P1_REIP_REG_15__SCAN_IN), 
        .B2(n16260), .ZN(n16261) );
  OAI211_X1 U19528 ( .C1(P1_REIP_REG_15__SCAN_IN), .C2(n16263), .A(n16262), 
        .B(n16261), .ZN(P1_U2825) );
  AOI21_X1 U19529 ( .B1(P1_REIP_REG_13__SCAN_IN), .B2(n16264), .A(
        P1_REIP_REG_14__SCAN_IN), .ZN(n16272) );
  AOI22_X1 U19530 ( .A1(n16371), .A2(n20149), .B1(n20147), .B2(
        P1_EBX_REG_14__SCAN_IN), .ZN(n16271) );
  INV_X1 U19531 ( .A(n16265), .ZN(n16269) );
  AOI21_X1 U19532 ( .B1(n20140), .B2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n20280), .ZN(n16266) );
  OAI21_X1 U19533 ( .B1(n20143), .B2(n16267), .A(n16266), .ZN(n16268) );
  AOI21_X1 U19534 ( .B1(n16269), .B2(n20131), .A(n16268), .ZN(n16270) );
  OAI211_X1 U19535 ( .C1(n16273), .C2(n16272), .A(n16271), .B(n16270), .ZN(
        P1_U2826) );
  OAI22_X1 U19536 ( .A1(n16275), .A2(n20124), .B1(n20122), .B2(n16274), .ZN(
        n16276) );
  INV_X1 U19537 ( .A(n16276), .ZN(n16284) );
  AOI22_X1 U19538 ( .A1(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n20140), .B1(
        n16277), .B2(n20154), .ZN(n16283) );
  OAI21_X1 U19539 ( .B1(n16278), .B2(n20105), .A(n20944), .ZN(n16279) );
  AOI22_X1 U19540 ( .A1(n20131), .A2(n16281), .B1(n16280), .B2(n16279), .ZN(
        n16282) );
  NAND4_X1 U19541 ( .A1(n16284), .A2(n16283), .A3(n16282), .A4(n20256), .ZN(
        P1_U2828) );
  NAND2_X1 U19542 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(n16285), .ZN(n16292) );
  INV_X1 U19543 ( .A(n16286), .ZN(n16377) );
  AOI22_X1 U19544 ( .A1(n16377), .A2(n20149), .B1(n20147), .B2(
        P1_EBX_REG_11__SCAN_IN), .ZN(n16287) );
  OAI21_X1 U19545 ( .B1(n16328), .B2(n20143), .A(n16287), .ZN(n16288) );
  AOI211_X1 U19546 ( .C1(n20140), .C2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .A(
        n20280), .B(n16288), .ZN(n16291) );
  AOI22_X1 U19547 ( .A1(P1_REIP_REG_11__SCAN_IN), .A2(n16289), .B1(n20131), 
        .B2(n16324), .ZN(n16290) );
  OAI211_X1 U19548 ( .C1(P1_REIP_REG_11__SCAN_IN), .C2(n16292), .A(n16291), 
        .B(n16290), .ZN(P1_U2829) );
  INV_X1 U19549 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n19393) );
  AOI22_X1 U19550 ( .A1(n16294), .A2(n20332), .B1(P1_EAX_REG_19__SCAN_IN), 
        .B2(n16293), .ZN(n16298) );
  AOI22_X1 U19551 ( .A1(n16296), .A2(n13019), .B1(n16295), .B2(DATAI_19_), 
        .ZN(n16297) );
  OAI211_X1 U19552 ( .C1(n16299), .C2(n19393), .A(n16298), .B(n16297), .ZN(
        P1_U2885) );
  AOI21_X1 U19553 ( .B1(n15219), .B2(n16301), .A(n16300), .ZN(n16304) );
  NOR2_X1 U19554 ( .A1(n16304), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n16303) );
  MUX2_X1 U19555 ( .A(n16304), .B(n16303), .S(n16302), .Z(n16305) );
  XNOR2_X1 U19556 ( .A(n16305), .B(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n16353) );
  AOI22_X1 U19557 ( .A1(n20242), .A2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B1(
        n20296), .B2(P1_REIP_REG_17__SCAN_IN), .ZN(n16309) );
  AOI22_X1 U19558 ( .A1(n16307), .A2(n16325), .B1(n16316), .B2(n16306), .ZN(
        n16308) );
  OAI211_X1 U19559 ( .C1(n16353), .C2(n20088), .A(n16309), .B(n16308), .ZN(
        P1_U2982) );
  NAND2_X1 U19560 ( .A1(n16311), .A2(n16310), .ZN(n16315) );
  NAND2_X1 U19561 ( .A1(n16313), .A2(n16312), .ZN(n16314) );
  XOR2_X1 U19562 ( .A(n16315), .B(n16314), .Z(n16368) );
  AOI22_X1 U19563 ( .A1(n20242), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B1(
        n20296), .B2(P1_REIP_REG_15__SCAN_IN), .ZN(n16320) );
  AOI22_X1 U19564 ( .A1(n16318), .A2(n16325), .B1(n16317), .B2(n16316), .ZN(
        n16319) );
  OAI211_X1 U19565 ( .C1(n16368), .C2(n20088), .A(n16320), .B(n16319), .ZN(
        P1_U2984) );
  AOI22_X1 U19566 ( .A1(n20242), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B1(
        n20296), .B2(P1_REIP_REG_11__SCAN_IN), .ZN(n16327) );
  NAND2_X1 U19567 ( .A1(n9845), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n16322) );
  OAI21_X1 U19568 ( .B1(n15219), .B2(n16322), .A(n16321), .ZN(n16323) );
  INV_X1 U19569 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16383) );
  XNOR2_X1 U19570 ( .A(n16323), .B(n16383), .ZN(n16378) );
  AOI22_X1 U19571 ( .A1(n20248), .A2(n16378), .B1(n16325), .B2(n16324), .ZN(
        n16326) );
  OAI211_X1 U19572 ( .C1(n20252), .C2(n16328), .A(n16327), .B(n16326), .ZN(
        P1_U2988) );
  AOI22_X1 U19573 ( .A1(n20242), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B1(
        n20296), .B2(P1_REIP_REG_7__SCAN_IN), .ZN(n16334) );
  NAND2_X1 U19574 ( .A1(n16331), .A2(n16330), .ZN(n16332) );
  XNOR2_X1 U19575 ( .A(n16329), .B(n16332), .ZN(n16412) );
  AOI22_X1 U19576 ( .A1(n16412), .A2(n20248), .B1(n16325), .B2(n20172), .ZN(
        n16333) );
  OAI211_X1 U19577 ( .C1(n20252), .C2(n20113), .A(n16334), .B(n16333), .ZN(
        P1_U2992) );
  AOI22_X1 U19578 ( .A1(n20242), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B1(
        n20296), .B2(P1_REIP_REG_6__SCAN_IN), .ZN(n16339) );
  XNOR2_X1 U19579 ( .A(n16335), .B(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n16336) );
  XNOR2_X1 U19580 ( .A(n16337), .B(n16336), .ZN(n16416) );
  AOI22_X1 U19581 ( .A1(n16416), .A2(n20248), .B1(n16325), .B2(n20132), .ZN(
        n16338) );
  OAI211_X1 U19582 ( .C1(n20252), .C2(n20127), .A(n16339), .B(n16338), .ZN(
        P1_U2993) );
  AOI22_X1 U19583 ( .A1(n20242), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .B1(
        n20296), .B2(P1_REIP_REG_5__SCAN_IN), .ZN(n16345) );
  OAI21_X1 U19584 ( .B1(n16342), .B2(n16341), .A(n16340), .ZN(n16343) );
  INV_X1 U19585 ( .A(n16343), .ZN(n16429) );
  AOI22_X1 U19586 ( .A1(n16429), .A2(n20248), .B1(n16325), .B2(n20179), .ZN(
        n16344) );
  OAI211_X1 U19587 ( .C1(n20252), .C2(n20142), .A(n16345), .B(n16344), .ZN(
        P1_U2994) );
  INV_X1 U19588 ( .A(n16346), .ZN(n16347) );
  AOI22_X1 U19589 ( .A1(n16347), .A2(n20282), .B1(n20280), .B2(
        P1_REIP_REG_17__SCAN_IN), .ZN(n16352) );
  NOR3_X1 U19590 ( .A1(n16421), .A2(n16348), .A3(n16369), .ZN(n16350) );
  OAI21_X1 U19591 ( .B1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n16350), .A(
        n16349), .ZN(n16351) );
  OAI211_X1 U19592 ( .C1(n16353), .C2(n20293), .A(n16352), .B(n16351), .ZN(
        P1_U3014) );
  INV_X1 U19593 ( .A(n16354), .ZN(n16355) );
  AOI21_X1 U19594 ( .B1(n16356), .B2(n20282), .A(n16355), .ZN(n16362) );
  OAI21_X1 U19595 ( .B1(n16402), .B2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n16357), .ZN(n16365) );
  AOI22_X1 U19596 ( .A1(n16358), .A2(n20278), .B1(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n16365), .ZN(n16361) );
  NOR3_X1 U19597 ( .A1(n16421), .A2(n16369), .A3(n12892), .ZN(n16364) );
  OAI221_X1 U19598 ( .B1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .C1(n11905), .C2(n16359), .A(
        n16364), .ZN(n16360) );
  NAND3_X1 U19599 ( .A1(n16362), .A2(n16361), .A3(n16360), .ZN(P1_U3015) );
  AOI22_X1 U19600 ( .A1(n16363), .A2(n20282), .B1(n20280), .B2(
        P1_REIP_REG_15__SCAN_IN), .ZN(n16367) );
  AOI22_X1 U19601 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n16365), .B1(
        n16364), .B2(n11905), .ZN(n16366) );
  OAI211_X1 U19602 ( .C1(n16368), .C2(n20293), .A(n16367), .B(n16366), .ZN(
        P1_U3016) );
  OR2_X1 U19603 ( .A1(n16369), .A2(n16421), .ZN(n16376) );
  AOI21_X1 U19604 ( .B1(n16371), .B2(n20282), .A(n16370), .ZN(n16375) );
  AOI22_X1 U19605 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n16373), .B1(
        n20278), .B2(n16372), .ZN(n16374) );
  OAI211_X1 U19606 ( .C1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n16376), .A(
        n16375), .B(n16374), .ZN(P1_U3017) );
  AOI22_X1 U19607 ( .A1(n16377), .A2(n20282), .B1(n20280), .B2(
        P1_REIP_REG_11__SCAN_IN), .ZN(n16382) );
  NOR2_X1 U19608 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n16421), .ZN(
        n16379) );
  AOI22_X1 U19609 ( .A1(n16380), .A2(n16379), .B1(n20278), .B2(n16378), .ZN(
        n16381) );
  OAI211_X1 U19610 ( .C1(n16384), .C2(n16383), .A(n16382), .B(n16381), .ZN(
        P1_U3020) );
  AOI21_X1 U19611 ( .B1(n16386), .B2(n20282), .A(n16385), .ZN(n16393) );
  AOI22_X1 U19612 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n16388), .B1(
        n20278), .B2(n16387), .ZN(n16392) );
  OAI221_X1 U19613 ( .B1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .C1(n15266), .C2(n16390), .A(
        n16389), .ZN(n16391) );
  NAND3_X1 U19614 ( .A1(n16393), .A2(n16392), .A3(n16391), .ZN(P1_U3021) );
  OAI21_X1 U19615 ( .B1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A(n16394), .ZN(n16406) );
  INV_X1 U19616 ( .A(n16395), .ZN(n16397) );
  AOI21_X1 U19617 ( .B1(n16397), .B2(n20282), .A(n16396), .ZN(n16405) );
  AOI21_X1 U19618 ( .B1(n16400), .B2(n16399), .A(n16398), .ZN(n16401) );
  INV_X1 U19619 ( .A(n16401), .ZN(n16428) );
  AOI21_X1 U19620 ( .B1(n16431), .B2(n16430), .A(n16428), .ZN(n16419) );
  OAI21_X1 U19621 ( .B1(n16402), .B2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n16419), .ZN(n16411) );
  AOI22_X1 U19622 ( .A1(n16403), .A2(n20278), .B1(
        P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n16411), .ZN(n16404) );
  OAI211_X1 U19623 ( .C1(n16415), .C2(n16406), .A(n16405), .B(n16404), .ZN(
        P1_U3023) );
  AND2_X1 U19624 ( .A1(n16408), .A2(n16407), .ZN(n16409) );
  NOR2_X1 U19625 ( .A1(n16410), .A2(n16409), .ZN(n20170) );
  AOI22_X1 U19626 ( .A1(n20170), .A2(n20282), .B1(n20280), .B2(
        P1_REIP_REG_7__SCAN_IN), .ZN(n16414) );
  AOI22_X1 U19627 ( .A1(n16412), .A2(n20278), .B1(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n16411), .ZN(n16413) );
  OAI211_X1 U19628 ( .C1(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .C2(n16415), .A(
        n16414), .B(n16413), .ZN(P1_U3024) );
  INV_X1 U19629 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n16420) );
  AOI222_X1 U19630 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(n20296), .B1(n20282), 
        .B2(n16417), .C1(n20278), .C2(n16416), .ZN(n16418) );
  OAI221_X1 U19631 ( .B1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n16421), .C1(
        n16420), .C2(n16419), .A(n16418), .ZN(P1_U3025) );
  NAND2_X1 U19632 ( .A1(n16424), .A2(n16423), .ZN(n20176) );
  INV_X1 U19633 ( .A(n20176), .ZN(n20138) );
  NOR2_X1 U19634 ( .A1(n16426), .A2(n16425), .ZN(n16427) );
  AOI22_X1 U19635 ( .A1(n20138), .A2(n20282), .B1(n20289), .B2(n16427), .ZN(
        n16435) );
  AOI22_X1 U19636 ( .A1(n16429), .A2(n20278), .B1(
        P1_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n16428), .ZN(n16434) );
  NAND2_X1 U19637 ( .A1(n16431), .A2(n16430), .ZN(n16433) );
  NAND2_X1 U19638 ( .A1(n20296), .A2(P1_REIP_REG_5__SCAN_IN), .ZN(n16432) );
  NAND4_X1 U19639 ( .A1(n16435), .A2(n16434), .A3(n16433), .A4(n16432), .ZN(
        P1_U3026) );
  NAND4_X1 U19640 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(
        P1_STATE2_REG_0__SCAN_IN), .A3(n20999), .A4(n21010), .ZN(n16436) );
  AND2_X1 U19641 ( .A1(n16437), .A2(n16436), .ZN(n20911) );
  NAND2_X1 U19642 ( .A1(n20911), .A2(n16438), .ZN(n16439) );
  AOI22_X1 U19643 ( .A1(n16442), .A2(n16441), .B1(n16440), .B2(n16439), .ZN(
        P1_U3162) );
  OAI21_X1 U19644 ( .B1(n20912), .B2(n20738), .A(n16443), .ZN(P1_U3466) );
  AOI211_X1 U19645 ( .C1(n16446), .C2(n16445), .A(n16444), .B(n19214), .ZN(
        n16454) );
  NAND2_X1 U19646 ( .A1(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n19166), .ZN(
        n16448) );
  AOI22_X1 U19647 ( .A1(P2_REIP_REG_26__SCAN_IN), .A2(n19210), .B1(
        P2_EBX_REG_26__SCAN_IN), .B2(n19205), .ZN(n16447) );
  NAND2_X1 U19648 ( .A1(n16448), .A2(n16447), .ZN(n16449) );
  AOI21_X1 U19649 ( .B1(n16450), .B2(n19186), .A(n16449), .ZN(n16451) );
  OAI21_X1 U19650 ( .B1(n16452), .B2(n19197), .A(n16451), .ZN(n16453) );
  AOI211_X1 U19651 ( .C1(n19183), .C2(n16455), .A(n16454), .B(n16453), .ZN(
        n16456) );
  INV_X1 U19652 ( .A(n16456), .ZN(P2_U2829) );
  AOI22_X1 U19653 ( .A1(n19221), .A2(n19409), .B1(n19257), .B2(
        P2_EAX_REG_22__SCAN_IN), .ZN(n16461) );
  AOI22_X1 U19654 ( .A1(n19223), .A2(BUF2_REG_22__SCAN_IN), .B1(n19222), .B2(
        BUF1_REG_22__SCAN_IN), .ZN(n16460) );
  AOI22_X1 U19655 ( .A1(n16458), .A2(n19270), .B1(n19265), .B2(n16457), .ZN(
        n16459) );
  NAND3_X1 U19656 ( .A1(n16461), .A2(n16460), .A3(n16459), .ZN(P2_U2897) );
  AOI22_X1 U19657 ( .A1(n19221), .A2(n19396), .B1(n19257), .B2(
        P2_EAX_REG_20__SCAN_IN), .ZN(n16465) );
  AOI22_X1 U19658 ( .A1(n19223), .A2(BUF2_REG_20__SCAN_IN), .B1(n19222), .B2(
        BUF1_REG_20__SCAN_IN), .ZN(n16464) );
  AOI22_X1 U19659 ( .A1(n16462), .A2(n19270), .B1(n19265), .B2(n9921), .ZN(
        n16463) );
  NAND3_X1 U19660 ( .A1(n16465), .A2(n16464), .A3(n16463), .ZN(P2_U2899) );
  AOI22_X1 U19661 ( .A1(n19221), .A2(n19381), .B1(n19257), .B2(
        P2_EAX_REG_18__SCAN_IN), .ZN(n16471) );
  AOI22_X1 U19662 ( .A1(n19223), .A2(BUF2_REG_18__SCAN_IN), .B1(n19222), .B2(
        BUF1_REG_18__SCAN_IN), .ZN(n16470) );
  INV_X1 U19663 ( .A(n16466), .ZN(n16467) );
  AOI22_X1 U19664 ( .A1(n16468), .A2(n19270), .B1(n19265), .B2(n16467), .ZN(
        n16469) );
  NAND3_X1 U19665 ( .A1(n16471), .A2(n16470), .A3(n16469), .ZN(P2_U2901) );
  AOI22_X1 U19666 ( .A1(P2_REIP_REG_23__SCAN_IN), .A2(n19170), .B1(n16550), 
        .B2(n16472), .ZN(n16478) );
  OAI22_X1 U19667 ( .A1(n16474), .A2(n19319), .B1(n16473), .B2(n16553), .ZN(
        n16475) );
  AOI21_X1 U19668 ( .B1(n19315), .B2(n16476), .A(n16475), .ZN(n16477) );
  OAI211_X1 U19669 ( .C1(n16559), .C2(n16479), .A(n16478), .B(n16477), .ZN(
        P2_U2991) );
  AOI22_X1 U19670 ( .A1(n19313), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B1(
        P2_REIP_REG_22__SCAN_IN), .B2(n19170), .ZN(n16483) );
  AOI22_X1 U19671 ( .A1(n19313), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .B1(
        P2_REIP_REG_18__SCAN_IN), .B2(n19170), .ZN(n16489) );
  AOI222_X1 U19672 ( .A1(n16487), .A2(n12840), .B1(n19315), .B2(n16486), .C1(
        n16539), .C2(n16485), .ZN(n16488) );
  OAI211_X1 U19673 ( .C1(n19325), .C2(n16490), .A(n16489), .B(n16488), .ZN(
        P2_U2996) );
  AOI22_X1 U19674 ( .A1(n19313), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B1(
        P2_REIP_REG_16__SCAN_IN), .B2(n19170), .ZN(n16498) );
  NAND2_X1 U19675 ( .A1(n16019), .A2(n16491), .ZN(n16492) );
  OAI211_X1 U19676 ( .C1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(n16492), .B(n16539), .ZN(
        n16494) );
  OAI22_X1 U19677 ( .A1(n9861), .A2(n16494), .B1(n16493), .B2(n16545), .ZN(
        n16495) );
  AOI21_X1 U19678 ( .B1(n16496), .B2(n12840), .A(n16495), .ZN(n16497) );
  OAI211_X1 U19679 ( .C1(n19325), .C2(n16499), .A(n16498), .B(n16497), .ZN(
        P2_U2998) );
  AOI22_X1 U19680 ( .A1(P2_REIP_REG_15__SCAN_IN), .A2(n19170), .B1(n16550), 
        .B2(n19087), .ZN(n16505) );
  OAI22_X1 U19681 ( .A1(n16501), .A2(n16553), .B1(n19319), .B2(n16500), .ZN(
        n16502) );
  AOI21_X1 U19682 ( .B1(n19315), .B2(n16503), .A(n16502), .ZN(n16504) );
  OAI211_X1 U19683 ( .C1(n16559), .C2(n16506), .A(n16505), .B(n16504), .ZN(
        P2_U2999) );
  AOI22_X1 U19684 ( .A1(n19313), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(
        P2_REIP_REG_14__SCAN_IN), .B2(n19170), .ZN(n16510) );
  AOI222_X1 U19685 ( .A1(n16508), .A2(n12840), .B1(n16507), .B2(n16539), .C1(
        n19315), .C2(n19102), .ZN(n16509) );
  OAI211_X1 U19686 ( .C1(n19325), .C2(n19097), .A(n16510), .B(n16509), .ZN(
        P2_U3000) );
  AOI22_X1 U19687 ( .A1(n19313), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        P2_REIP_REG_12__SCAN_IN), .B2(n19170), .ZN(n16516) );
  AOI21_X1 U19688 ( .B1(n16512), .B2(n16570), .A(n16511), .ZN(n16567) );
  XNOR2_X1 U19689 ( .A(n16513), .B(n16514), .ZN(n16566) );
  AOI222_X1 U19690 ( .A1(n16567), .A2(n16539), .B1(n12840), .B2(n16566), .C1(
        n19315), .C2(n16565), .ZN(n16515) );
  OAI211_X1 U19691 ( .C1(n19325), .C2(n16517), .A(n16516), .B(n16515), .ZN(
        P2_U3002) );
  AOI22_X1 U19692 ( .A1(n19313), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B1(
        P2_REIP_REG_10__SCAN_IN), .B2(n19170), .ZN(n16522) );
  AOI222_X1 U19693 ( .A1(n16520), .A2(n12840), .B1(n19315), .B2(n16519), .C1(
        n16539), .C2(n16518), .ZN(n16521) );
  OAI211_X1 U19694 ( .C1(n19325), .C2(n16523), .A(n16522), .B(n16521), .ZN(
        P2_U3004) );
  AOI22_X1 U19695 ( .A1(P2_REIP_REG_9__SCAN_IN), .A2(n19170), .B1(n16550), 
        .B2(n19132), .ZN(n16528) );
  OAI22_X1 U19696 ( .A1(n16525), .A2(n19319), .B1(n16553), .B2(n16524), .ZN(
        n16526) );
  AOI21_X1 U19697 ( .B1(n19315), .B2(n19136), .A(n16526), .ZN(n16527) );
  OAI211_X1 U19698 ( .C1(n16559), .C2(n16529), .A(n16528), .B(n16527), .ZN(
        P2_U3005) );
  AOI22_X1 U19699 ( .A1(n19313), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B1(
        P2_REIP_REG_8__SCAN_IN), .B2(n19170), .ZN(n16541) );
  NAND2_X1 U19700 ( .A1(n16531), .A2(n16530), .ZN(n16536) );
  INV_X1 U19701 ( .A(n16532), .ZN(n16533) );
  AOI21_X1 U19702 ( .B1(n14410), .B2(n16534), .A(n16533), .ZN(n16535) );
  XOR2_X1 U19703 ( .A(n16536), .B(n16535), .Z(n16579) );
  XOR2_X1 U19704 ( .A(n16537), .B(n16538), .Z(n16576) );
  AOI222_X1 U19705 ( .A1(n16579), .A2(n12840), .B1(n19315), .B2(n16578), .C1(
        n16539), .C2(n16576), .ZN(n16540) );
  OAI211_X1 U19706 ( .C1(n19325), .C2(n16542), .A(n16541), .B(n16540), .ZN(
        P2_U3006) );
  AOI22_X1 U19707 ( .A1(n19313), .A2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B1(
        P2_REIP_REG_6__SCAN_IN), .B2(n19170), .ZN(n16549) );
  OAI222_X1 U19708 ( .A1(n16546), .A2(n16545), .B1(n16544), .B2(n16553), .C1(
        n19319), .C2(n16543), .ZN(n16547) );
  INV_X1 U19709 ( .A(n16547), .ZN(n16548) );
  OAI211_X1 U19710 ( .C1(n19325), .C2(n19160), .A(n16549), .B(n16548), .ZN(
        P2_U3008) );
  AOI22_X1 U19711 ( .A1(P2_REIP_REG_5__SCAN_IN), .A2(n19170), .B1(n16550), 
        .B2(n19173), .ZN(n16557) );
  INV_X1 U19712 ( .A(n16551), .ZN(n16554) );
  OAI22_X1 U19713 ( .A1(n16554), .A2(n19319), .B1(n16553), .B2(n16552), .ZN(
        n16555) );
  AOI21_X1 U19714 ( .B1(n19315), .B2(n19174), .A(n16555), .ZN(n16556) );
  OAI211_X1 U19715 ( .C1(n16559), .C2(n16558), .A(n16557), .B(n16556), .ZN(
        P2_U3009) );
  AOI21_X1 U19716 ( .B1(n16562), .B2(n16561), .A(n16560), .ZN(n16571) );
  NOR2_X1 U19717 ( .A1(n19345), .A2(n19952), .ZN(n16564) );
  AOI211_X1 U19718 ( .C1(n19238), .C2(n19347), .A(n16564), .B(n16563), .ZN(
        n16569) );
  AOI222_X1 U19719 ( .A1(n16567), .A2(n16577), .B1(n19331), .B2(n16566), .C1(
        n19341), .C2(n16565), .ZN(n16568) );
  OAI211_X1 U19720 ( .C1(n16571), .C2(n16570), .A(n16569), .B(n16568), .ZN(
        P2_U3034) );
  OAI22_X1 U19721 ( .A1(n16574), .A2(n16573), .B1(n19327), .B2(n16572), .ZN(
        n16575) );
  INV_X1 U19722 ( .A(n16575), .ZN(n16585) );
  AOI222_X1 U19723 ( .A1(n16579), .A2(n19331), .B1(n19341), .B2(n16578), .C1(
        n16577), .C2(n16576), .ZN(n16584) );
  NAND2_X1 U19724 ( .A1(P2_REIP_REG_8__SCAN_IN), .A2(n19170), .ZN(n16583) );
  OAI211_X1 U19725 ( .C1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(n16581), .B(n16580), .ZN(n16582) );
  NAND4_X1 U19726 ( .A1(n16585), .A2(n16584), .A3(n16583), .A4(n16582), .ZN(
        P2_U3038) );
  OAI21_X1 U19727 ( .B1(n20035), .B2(n20034), .A(n16594), .ZN(n16588) );
  AOI211_X1 U19728 ( .C1(P2_STATE2_REG_0__SCAN_IN), .C2(n16588), .A(n16587), 
        .B(n16586), .ZN(n16592) );
  AOI21_X1 U19729 ( .B1(n20067), .B2(n16589), .A(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n16590) );
  OAI21_X1 U19730 ( .B1(n16594), .B2(n20069), .A(n16590), .ZN(n16591) );
  OAI211_X1 U19731 ( .C1(n16593), .C2(n19040), .A(n16592), .B(n16591), .ZN(
        P2_U3176) );
  AND2_X1 U19732 ( .A1(n16594), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n16596) );
  OAI21_X1 U19733 ( .B1(n16596), .B2(n20036), .A(n16595), .ZN(P2_U3593) );
  XOR2_X1 U19734 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B(n16614), .Z(
        n16765) );
  INV_X1 U19735 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n16769) );
  INV_X2 U19736 ( .A(n18316), .ZN(n18096) );
  NAND2_X1 U19737 ( .A1(n18096), .A2(P3_REIP_REG_30__SCAN_IN), .ZN(n16597) );
  OAI221_X1 U19738 ( .B1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n16599), .C1(
        n16769), .C2(n16598), .A(n16597), .ZN(n16600) );
  AOI21_X1 U19739 ( .B1(n17895), .B2(n16765), .A(n16600), .ZN(n16607) );
  INV_X1 U19740 ( .A(n17926), .ZN(n17961) );
  OAI22_X1 U19741 ( .A1(n16609), .A2(n18050), .B1(n16608), .B2(n17961), .ZN(
        n16602) );
  AOI22_X1 U19742 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16602), .B1(
        n17963), .B2(n16601), .ZN(n16606) );
  AOI22_X2 U19743 ( .A1(n18039), .A2(n18215), .B1(n17926), .B2(n18214), .ZN(
        n17953) );
  NOR2_X2 U19744 ( .A1(n17953), .A2(n16637), .ZN(n17849) );
  NOR2_X1 U19745 ( .A1(n18095), .A2(n17864), .ZN(n17772) );
  NAND4_X1 U19746 ( .A1(n17716), .A2(n16604), .A3(n17772), .A4(n16603), .ZN(
        n16605) );
  NAND3_X1 U19747 ( .A1(n16607), .A2(n16606), .A3(n16605), .ZN(P3_U2800) );
  AOI211_X1 U19748 ( .C1(n16610), .C2(n16625), .A(n16608), .B(n17961), .ZN(
        n16612) );
  AOI211_X1 U19749 ( .C1(n16631), .C2(n16610), .A(n16609), .B(n18050), .ZN(
        n16611) );
  AOI211_X1 U19750 ( .C1(n17963), .C2(n16613), .A(n16612), .B(n16611), .ZN(
        n16621) );
  INV_X1 U19751 ( .A(n16747), .ZN(n16615) );
  AOI21_X1 U19752 ( .B1(n10099), .B2(n16615), .A(n16614), .ZN(n16776) );
  OAI21_X1 U19753 ( .B1(n16616), .B2(n17895), .A(n16776), .ZN(n16619) );
  OAI221_X1 U19754 ( .B1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n18748), .C1(
        P3_PHYADDRPOINTER_REG_29__SCAN_IN), .C2(n9962), .A(n16617), .ZN(n16618) );
  NAND4_X1 U19755 ( .A1(n16621), .A2(n16620), .A3(n16619), .A4(n16618), .ZN(
        P3_U2801) );
  INV_X1 U19756 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n18948) );
  INV_X1 U19757 ( .A(n16638), .ZN(n16622) );
  AOI22_X1 U19758 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n13160), .B1(
        n17957), .B2(n17693), .ZN(n17696) );
  AOI21_X1 U19759 ( .B1(n16623), .B2(n16622), .A(n17695), .ZN(n16629) );
  NOR2_X1 U19760 ( .A1(n16625), .A2(n16624), .ZN(n16627) );
  AOI211_X1 U19761 ( .C1(n18244), .C2(n16631), .A(n18349), .B(n16630), .ZN(
        n16632) );
  AOI21_X1 U19762 ( .B1(n16633), .B2(n16632), .A(n18096), .ZN(n16643) );
  INV_X1 U19763 ( .A(n16634), .ZN(n16639) );
  INV_X1 U19764 ( .A(n18244), .ZN(n18806) );
  NAND2_X1 U19765 ( .A1(n18804), .A2(n17551), .ZN(n18113) );
  OAI22_X1 U19766 ( .A1(n18806), .A2(n18194), .B1(n18188), .B2(n18113), .ZN(
        n16635) );
  INV_X1 U19767 ( .A(n16635), .ZN(n18051) );
  NAND3_X1 U19768 ( .A1(n16636), .A2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A3(
        n18324), .ZN(n18294) );
  NOR2_X1 U19769 ( .A1(n18295), .A2(n18294), .ZN(n18213) );
  NAND2_X1 U19770 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n18213), .ZN(
        n18186) );
  AOI211_X1 U19771 ( .C1(n18051), .C2(n18186), .A(n16637), .B(n18349), .ZN(
        n18182) );
  INV_X1 U19772 ( .A(n18182), .ZN(n18148) );
  OAI33_X1 U19773 ( .A1(n16639), .A2(n18114), .A3(n18148), .B1(n18211), .B2(
        n16638), .B3(n17695), .ZN(n16642) );
  INV_X1 U19774 ( .A(n17696), .ZN(n16640) );
  NOR3_X1 U19775 ( .A1(n16640), .A2(n18211), .A3(n17709), .ZN(n16641) );
  OAI21_X1 U19776 ( .B1(n18316), .B2(n18948), .A(n16644), .ZN(P3_U2834) );
  NOR3_X1 U19777 ( .A1(P3_W_R_N_REG_SCAN_IN), .A2(P3_BE_N_REG_0__SCAN_IN), 
        .A3(P3_BE_N_REG_1__SCAN_IN), .ZN(n16646) );
  NOR4_X1 U19778 ( .A1(P3_BE_N_REG_2__SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(P3_D_C_N_REG_SCAN_IN), .A4(P3_ADS_N_REG_SCAN_IN), .ZN(n16645) );
  NAND4_X1 U19779 ( .A1(P3_M_IO_N_REG_SCAN_IN), .A2(n16646), .A3(n16645), .A4(
        U215), .ZN(U213) );
  INV_X1 U19780 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n19275) );
  INV_X2 U19781 ( .A(U214), .ZN(n16691) );
  NOR2_X1 U19782 ( .A1(n16691), .A2(n16647), .ZN(n16690) );
  INV_X1 U19783 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n16721) );
  OAI222_X1 U19784 ( .A1(U212), .A2(n19275), .B1(n16686), .B2(n20347), .C1(
        U214), .C2(n16721), .ZN(U216) );
  INV_X1 U19785 ( .A(BUF1_REG_30__SCAN_IN), .ZN(n19410) );
  INV_X1 U19786 ( .A(U212), .ZN(n16689) );
  AOI22_X1 U19787 ( .A1(P1_DATAO_REG_30__SCAN_IN), .A2(n16691), .B1(
        P2_DATAO_REG_30__SCAN_IN), .B2(n16689), .ZN(n16648) );
  OAI21_X1 U19788 ( .B1(n19410), .B2(n16686), .A(n16648), .ZN(U217) );
  INV_X1 U19789 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n19404) );
  AOI22_X1 U19790 ( .A1(P1_DATAO_REG_29__SCAN_IN), .A2(n16691), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n16689), .ZN(n16649) );
  OAI21_X1 U19791 ( .B1(n19404), .B2(n16686), .A(n16649), .ZN(U218) );
  INV_X1 U19792 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n19398) );
  AOI22_X1 U19793 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(n16691), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(n16689), .ZN(n16650) );
  OAI21_X1 U19794 ( .B1(n19398), .B2(n16686), .A(n16650), .ZN(U219) );
  INV_X1 U19795 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n19390) );
  AOI22_X1 U19796 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(n16691), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(n16689), .ZN(n16651) );
  OAI21_X1 U19797 ( .B1(n19390), .B2(n16686), .A(n16651), .ZN(U220) );
  INV_X1 U19798 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n19383) );
  AOI22_X1 U19799 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(n16691), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(n16689), .ZN(n16652) );
  OAI21_X1 U19800 ( .B1(n19383), .B2(n16686), .A(n16652), .ZN(U221) );
  AOI22_X1 U19801 ( .A1(P1_DATAO_REG_25__SCAN_IN), .A2(n16691), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(n16689), .ZN(n16653) );
  OAI21_X1 U19802 ( .B1(n16654), .B2(n16686), .A(n16653), .ZN(U222) );
  AOI22_X1 U19803 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n16691), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(n16689), .ZN(n16655) );
  OAI21_X1 U19804 ( .B1(n16656), .B2(n16686), .A(n16655), .ZN(U223) );
  INV_X1 U19805 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n19425) );
  AOI22_X1 U19806 ( .A1(P1_DATAO_REG_23__SCAN_IN), .A2(n16691), .B1(
        P2_DATAO_REG_23__SCAN_IN), .B2(n16689), .ZN(n16657) );
  OAI21_X1 U19807 ( .B1(n19425), .B2(n16686), .A(n16657), .ZN(U224) );
  INV_X1 U19808 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n16658) );
  INV_X1 U19809 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n19414) );
  INV_X1 U19810 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n21269) );
  OAI222_X1 U19811 ( .A1(U214), .A2(n16658), .B1(n16686), .B2(n19414), .C1(
        U212), .C2(n21269), .ZN(U225) );
  INV_X1 U19812 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n19406) );
  INV_X1 U19813 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n16659) );
  OAI222_X1 U19814 ( .A1(U212), .A2(n16711), .B1(n16686), .B2(n19406), .C1(
        U214), .C2(n16659), .ZN(U226) );
  INV_X1 U19815 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n19400) );
  AOI22_X1 U19816 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n16691), .B1(
        P2_DATAO_REG_20__SCAN_IN), .B2(n16689), .ZN(n16660) );
  OAI21_X1 U19817 ( .B1(n19400), .B2(n16686), .A(n16660), .ZN(U227) );
  AOI22_X1 U19818 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(n16691), .B1(
        P2_DATAO_REG_19__SCAN_IN), .B2(n16689), .ZN(n16661) );
  OAI21_X1 U19819 ( .B1(n19393), .B2(n16686), .A(n16661), .ZN(U228) );
  AOI22_X1 U19820 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(n16691), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n16689), .ZN(n16662) );
  OAI21_X1 U19821 ( .B1(n15095), .B2(n16686), .A(n16662), .ZN(U229) );
  AOI22_X1 U19822 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(n16691), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n16689), .ZN(n16663) );
  OAI21_X1 U19823 ( .B1(n16664), .B2(n16686), .A(n16663), .ZN(U230) );
  INV_X1 U19824 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n16666) );
  OAI222_X1 U19825 ( .A1(U214), .A2(n16666), .B1(n16686), .B2(n16665), .C1(
        U212), .C2(n21162), .ZN(U231) );
  INV_X1 U19826 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n19279) );
  AOI22_X1 U19827 ( .A1(BUF1_REG_15__SCAN_IN), .A2(n16690), .B1(
        P1_DATAO_REG_15__SCAN_IN), .B2(n16691), .ZN(n16667) );
  OAI21_X1 U19828 ( .B1(n19279), .B2(U212), .A(n16667), .ZN(U232) );
  INV_X1 U19829 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n16705) );
  AOI22_X1 U19830 ( .A1(BUF1_REG_14__SCAN_IN), .A2(n16690), .B1(
        P1_DATAO_REG_14__SCAN_IN), .B2(n16691), .ZN(n16668) );
  OAI21_X1 U19831 ( .B1(n16705), .B2(U212), .A(n16668), .ZN(U233) );
  INV_X1 U19832 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n16703) );
  AOI22_X1 U19833 ( .A1(BUF1_REG_13__SCAN_IN), .A2(n16690), .B1(
        P1_DATAO_REG_13__SCAN_IN), .B2(n16691), .ZN(n16669) );
  OAI21_X1 U19834 ( .B1(n16703), .B2(U212), .A(n16669), .ZN(U234) );
  AOI22_X1 U19835 ( .A1(P1_DATAO_REG_12__SCAN_IN), .A2(n16691), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n16689), .ZN(n16670) );
  OAI21_X1 U19836 ( .B1(n16671), .B2(n16686), .A(n16670), .ZN(U235) );
  AOI22_X1 U19837 ( .A1(P1_DATAO_REG_11__SCAN_IN), .A2(n16691), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n16689), .ZN(n16672) );
  OAI21_X1 U19838 ( .B1(n16673), .B2(n16686), .A(n16672), .ZN(U236) );
  AOI222_X1 U19839 ( .A1(n16689), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n16690), 
        .B2(BUF1_REG_10__SCAN_IN), .C1(n16691), .C2(P1_DATAO_REG_10__SCAN_IN), 
        .ZN(n16674) );
  INV_X1 U19840 ( .A(n16674), .ZN(U237) );
  INV_X1 U19841 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n16700) );
  AOI22_X1 U19842 ( .A1(BUF1_REG_9__SCAN_IN), .A2(n16690), .B1(
        P1_DATAO_REG_9__SCAN_IN), .B2(n16691), .ZN(n16675) );
  OAI21_X1 U19843 ( .B1(n16700), .B2(U212), .A(n16675), .ZN(U238) );
  AOI22_X1 U19844 ( .A1(P1_DATAO_REG_8__SCAN_IN), .A2(n16691), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n16689), .ZN(n16676) );
  OAI21_X1 U19845 ( .B1(n16677), .B2(n16686), .A(n16676), .ZN(U239) );
  INV_X1 U19846 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n16698) );
  AOI22_X1 U19847 ( .A1(BUF1_REG_7__SCAN_IN), .A2(n16690), .B1(
        P1_DATAO_REG_7__SCAN_IN), .B2(n16691), .ZN(n16678) );
  OAI21_X1 U19848 ( .B1(n16698), .B2(U212), .A(n16678), .ZN(U240) );
  AOI22_X1 U19849 ( .A1(P1_DATAO_REG_6__SCAN_IN), .A2(n16691), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n16689), .ZN(n16679) );
  OAI21_X1 U19850 ( .B1(n16680), .B2(n16686), .A(n16679), .ZN(U241) );
  INV_X1 U19851 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n16696) );
  INV_X1 U19852 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n21289) );
  OAI222_X1 U19853 ( .A1(U212), .A2(n16696), .B1(n16686), .B2(n16681), .C1(
        U214), .C2(n21289), .ZN(U242) );
  AOI22_X1 U19854 ( .A1(P1_DATAO_REG_4__SCAN_IN), .A2(n16691), .B1(
        P2_DATAO_REG_4__SCAN_IN), .B2(n16689), .ZN(n16682) );
  OAI21_X1 U19855 ( .B1(n16683), .B2(n16686), .A(n16682), .ZN(U243) );
  INV_X1 U19856 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n16694) );
  AOI22_X1 U19857 ( .A1(BUF1_REG_3__SCAN_IN), .A2(n16690), .B1(
        P1_DATAO_REG_3__SCAN_IN), .B2(n16691), .ZN(n16684) );
  OAI21_X1 U19858 ( .B1(n16694), .B2(U212), .A(n16684), .ZN(U244) );
  AOI22_X1 U19859 ( .A1(P1_DATAO_REG_2__SCAN_IN), .A2(n16691), .B1(
        P2_DATAO_REG_2__SCAN_IN), .B2(n16689), .ZN(n16685) );
  OAI21_X1 U19860 ( .B1(n16687), .B2(n16686), .A(n16685), .ZN(U245) );
  AOI222_X1 U19861 ( .A1(n16689), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(n16690), 
        .B2(BUF1_REG_1__SCAN_IN), .C1(n16691), .C2(P1_DATAO_REG_1__SCAN_IN), 
        .ZN(n16688) );
  INV_X1 U19862 ( .A(n16688), .ZN(U246) );
  AOI222_X1 U19863 ( .A1(n16691), .A2(P1_DATAO_REG_0__SCAN_IN), .B1(n16690), 
        .B2(BUF1_REG_0__SCAN_IN), .C1(n16689), .C2(P2_DATAO_REG_0__SCAN_IN), 
        .ZN(n16692) );
  INV_X1 U19864 ( .A(n16692), .ZN(U247) );
  INV_X1 U19865 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n21122) );
  INV_X1 U19866 ( .A(BUF2_REG_0__SCAN_IN), .ZN(n18380) );
  AOI22_X1 U19867 ( .A1(n16717), .A2(n21122), .B1(n18380), .B2(U215), .ZN(U251) );
  INV_X1 U19868 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n19306) );
  INV_X1 U19869 ( .A(BUF2_REG_1__SCAN_IN), .ZN(n18388) );
  AOI22_X1 U19870 ( .A1(n16717), .A2(n19306), .B1(n18388), .B2(U215), .ZN(U252) );
  INV_X1 U19871 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n16693) );
  AOI22_X1 U19872 ( .A1(n16717), .A2(n16693), .B1(n18394), .B2(U215), .ZN(U253) );
  INV_X1 U19873 ( .A(BUF2_REG_3__SCAN_IN), .ZN(n18398) );
  AOI22_X1 U19874 ( .A1(n16717), .A2(n16694), .B1(n18398), .B2(U215), .ZN(U254) );
  INV_X1 U19875 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n16695) );
  AOI22_X1 U19876 ( .A1(n16717), .A2(n16695), .B1(n18402), .B2(U215), .ZN(U255) );
  INV_X1 U19877 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n18406) );
  AOI22_X1 U19878 ( .A1(n16717), .A2(n16696), .B1(n18406), .B2(U215), .ZN(U256) );
  INV_X1 U19879 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n16697) );
  AOI22_X1 U19880 ( .A1(n16717), .A2(n16697), .B1(n18410), .B2(U215), .ZN(U257) );
  INV_X1 U19881 ( .A(BUF2_REG_7__SCAN_IN), .ZN(n18416) );
  AOI22_X1 U19882 ( .A1(n16717), .A2(n16698), .B1(n18416), .B2(U215), .ZN(U258) );
  INV_X1 U19883 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n16699) );
  INV_X1 U19884 ( .A(BUF2_REG_8__SCAN_IN), .ZN(n17668) );
  AOI22_X1 U19885 ( .A1(n16717), .A2(n16699), .B1(n17668), .B2(U215), .ZN(U259) );
  INV_X1 U19886 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n17670) );
  AOI22_X1 U19887 ( .A1(n16717), .A2(n16700), .B1(n17670), .B2(U215), .ZN(U260) );
  INV_X1 U19888 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n19288) );
  INV_X1 U19889 ( .A(BUF2_REG_10__SCAN_IN), .ZN(n17672) );
  AOI22_X1 U19890 ( .A1(n16717), .A2(n19288), .B1(n17672), .B2(U215), .ZN(U261) );
  OAI22_X1 U19891 ( .A1(U215), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(
        BUF2_REG_11__SCAN_IN), .B2(n16717), .ZN(n16701) );
  INV_X1 U19892 ( .A(n16701), .ZN(U262) );
  INV_X1 U19893 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n16702) );
  INV_X1 U19894 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n17676) );
  AOI22_X1 U19895 ( .A1(n16717), .A2(n16702), .B1(n17676), .B2(U215), .ZN(U263) );
  INV_X1 U19896 ( .A(BUF2_REG_13__SCAN_IN), .ZN(n17681) );
  AOI22_X1 U19897 ( .A1(n16717), .A2(n16703), .B1(n17681), .B2(U215), .ZN(U264) );
  INV_X1 U19898 ( .A(BUF2_REG_14__SCAN_IN), .ZN(n16704) );
  AOI22_X1 U19899 ( .A1(n16717), .A2(n16705), .B1(n16704), .B2(U215), .ZN(U265) );
  INV_X1 U19900 ( .A(BUF2_REG_15__SCAN_IN), .ZN(n16706) );
  AOI22_X1 U19901 ( .A1(n16717), .A2(n19279), .B1(n16706), .B2(U215), .ZN(U266) );
  AOI22_X1 U19902 ( .A1(n16717), .A2(n21162), .B1(n18384), .B2(U215), .ZN(U267) );
  INV_X1 U19903 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n16707) );
  AOI22_X1 U19904 ( .A1(n16717), .A2(n16707), .B1(n18389), .B2(U215), .ZN(U268) );
  INV_X1 U19905 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n16708) );
  INV_X1 U19906 ( .A(BUF2_REG_18__SCAN_IN), .ZN(n19385) );
  AOI22_X1 U19907 ( .A1(n16717), .A2(n16708), .B1(n19385), .B2(U215), .ZN(U269) );
  INV_X1 U19908 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n16709) );
  AOI22_X1 U19909 ( .A1(n16717), .A2(n16709), .B1(n19392), .B2(U215), .ZN(U270) );
  INV_X1 U19910 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n16710) );
  INV_X1 U19911 ( .A(BUF2_REG_20__SCAN_IN), .ZN(n19399) );
  AOI22_X1 U19912 ( .A1(n16717), .A2(n16710), .B1(n19399), .B2(U215), .ZN(U271) );
  INV_X1 U19913 ( .A(BUF2_REG_21__SCAN_IN), .ZN(n21192) );
  AOI22_X1 U19914 ( .A1(n16717), .A2(n16711), .B1(n21192), .B2(U215), .ZN(U272) );
  INV_X1 U19915 ( .A(BUF2_REG_22__SCAN_IN), .ZN(n19413) );
  AOI22_X1 U19916 ( .A1(n16717), .A2(n21269), .B1(n19413), .B2(U215), .ZN(U273) );
  INV_X1 U19917 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n16712) );
  INV_X1 U19918 ( .A(BUF2_REG_23__SCAN_IN), .ZN(n19423) );
  AOI22_X1 U19919 ( .A1(n16717), .A2(n16712), .B1(n19423), .B2(U215), .ZN(U274) );
  INV_X1 U19920 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n16713) );
  AOI22_X1 U19921 ( .A1(n16717), .A2(n16713), .B1(n18379), .B2(U215), .ZN(U275) );
  INV_X1 U19922 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n16714) );
  AOI22_X1 U19923 ( .A1(n16717), .A2(n16714), .B1(n18390), .B2(U215), .ZN(U276) );
  INV_X1 U19924 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n16715) );
  INV_X1 U19925 ( .A(BUF2_REG_26__SCAN_IN), .ZN(n19382) );
  AOI22_X1 U19926 ( .A1(n16717), .A2(n16715), .B1(n19382), .B2(U215), .ZN(U277) );
  INV_X1 U19927 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n16716) );
  AOI22_X1 U19928 ( .A1(n16717), .A2(n16716), .B1(n19389), .B2(U215), .ZN(U278) );
  INV_X1 U19929 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n16718) );
  INV_X1 U19930 ( .A(BUF2_REG_28__SCAN_IN), .ZN(n19397) );
  AOI22_X1 U19931 ( .A1(n16717), .A2(n16718), .B1(n19397), .B2(U215), .ZN(U279) );
  INV_X1 U19932 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n16719) );
  INV_X1 U19933 ( .A(BUF2_REG_29__SCAN_IN), .ZN(n19405) );
  AOI22_X1 U19934 ( .A1(n16717), .A2(n16719), .B1(n19405), .B2(U215), .ZN(U280) );
  INV_X1 U19935 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n16720) );
  INV_X1 U19936 ( .A(BUF2_REG_30__SCAN_IN), .ZN(n19411) );
  AOI22_X1 U19937 ( .A1(n16717), .A2(n16720), .B1(n19411), .B2(U215), .ZN(U281) );
  INV_X1 U19938 ( .A(BUF2_REG_31__SCAN_IN), .ZN(n19418) );
  AOI22_X1 U19939 ( .A1(n16717), .A2(n19275), .B1(n19418), .B2(U215), .ZN(U282) );
  AOI222_X1 U19940 ( .A1(n16721), .A2(P1_DATAO_REG_30__SCAN_IN), .B1(n19275), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .C1(n17583), .C2(
        P3_DATAO_REG_30__SCAN_IN), .ZN(n16722) );
  INV_X2 U19941 ( .A(n16724), .ZN(n16723) );
  INV_X1 U19942 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n18915) );
  INV_X1 U19943 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n19950) );
  AOI22_X1 U19944 ( .A1(n16723), .A2(n18915), .B1(n19950), .B2(n16724), .ZN(
        U347) );
  INV_X1 U19945 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n18913) );
  INV_X1 U19946 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n19949) );
  AOI22_X1 U19947 ( .A1(n16723), .A2(n18913), .B1(n19949), .B2(n16724), .ZN(
        U348) );
  INV_X1 U19948 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n18911) );
  INV_X1 U19949 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n19947) );
  AOI22_X1 U19950 ( .A1(n16723), .A2(n18911), .B1(n19947), .B2(n16724), .ZN(
        U349) );
  INV_X1 U19951 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n18910) );
  INV_X1 U19952 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n19946) );
  AOI22_X1 U19953 ( .A1(n16723), .A2(n18910), .B1(n19946), .B2(n16724), .ZN(
        U350) );
  INV_X1 U19954 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n18908) );
  INV_X1 U19955 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n19944) );
  AOI22_X1 U19956 ( .A1(n16723), .A2(n18908), .B1(n19944), .B2(n16724), .ZN(
        U351) );
  INV_X1 U19957 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n18905) );
  INV_X1 U19958 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n19942) );
  AOI22_X1 U19959 ( .A1(n16723), .A2(n18905), .B1(n19942), .B2(n16724), .ZN(
        U352) );
  INV_X1 U19960 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n18904) );
  INV_X1 U19961 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n19940) );
  AOI22_X1 U19962 ( .A1(n16723), .A2(n18904), .B1(n19940), .B2(n16724), .ZN(
        U353) );
  INV_X1 U19963 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n18902) );
  AOI22_X1 U19964 ( .A1(n16723), .A2(n18902), .B1(n19939), .B2(n16724), .ZN(
        U354) );
  INV_X1 U19965 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n18952) );
  INV_X1 U19966 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n19985) );
  AOI22_X1 U19967 ( .A1(n16723), .A2(n18952), .B1(n19985), .B2(n16724), .ZN(
        U355) );
  INV_X1 U19968 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n18950) );
  INV_X1 U19969 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n19982) );
  AOI22_X1 U19970 ( .A1(n16723), .A2(n18950), .B1(n19982), .B2(n16724), .ZN(
        U356) );
  INV_X1 U19971 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n18947) );
  INV_X1 U19972 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n19980) );
  AOI22_X1 U19973 ( .A1(n16723), .A2(n18947), .B1(n19980), .B2(n16724), .ZN(
        U357) );
  INV_X1 U19974 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n21093) );
  INV_X1 U19975 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n19977) );
  AOI22_X1 U19976 ( .A1(n16723), .A2(n21093), .B1(n19977), .B2(n16724), .ZN(
        U358) );
  INV_X1 U19977 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n18944) );
  INV_X1 U19978 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n19976) );
  AOI22_X1 U19979 ( .A1(n16723), .A2(n18944), .B1(n19976), .B2(n16724), .ZN(
        U359) );
  INV_X1 U19980 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n18942) );
  INV_X1 U19981 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n19974) );
  AOI22_X1 U19982 ( .A1(n16723), .A2(n18942), .B1(n19974), .B2(n16724), .ZN(
        U360) );
  INV_X1 U19983 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n18940) );
  INV_X1 U19984 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n21195) );
  AOI22_X1 U19985 ( .A1(n16723), .A2(n18940), .B1(n21195), .B2(n16724), .ZN(
        U361) );
  INV_X1 U19986 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n18937) );
  INV_X1 U19987 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n19971) );
  AOI22_X1 U19988 ( .A1(n16723), .A2(n18937), .B1(n19971), .B2(n16724), .ZN(
        U362) );
  INV_X1 U19989 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n18936) );
  INV_X1 U19990 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n19969) );
  AOI22_X1 U19991 ( .A1(n16723), .A2(n18936), .B1(n19969), .B2(n16724), .ZN(
        U363) );
  INV_X1 U19992 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n18934) );
  INV_X1 U19993 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n19967) );
  AOI22_X1 U19994 ( .A1(n16723), .A2(n18934), .B1(n19967), .B2(n16724), .ZN(
        U364) );
  INV_X1 U19995 ( .A(P3_ADDRESS_REG_1__SCAN_IN), .ZN(n18900) );
  INV_X1 U19996 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n19937) );
  AOI22_X1 U19997 ( .A1(n16723), .A2(n18900), .B1(n19937), .B2(n16724), .ZN(
        U365) );
  INV_X1 U19998 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n18932) );
  INV_X1 U19999 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n19965) );
  AOI22_X1 U20000 ( .A1(n16723), .A2(n18932), .B1(n19965), .B2(n16724), .ZN(
        U366) );
  INV_X1 U20001 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n18930) );
  INV_X1 U20002 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n19963) );
  AOI22_X1 U20003 ( .A1(n16723), .A2(n18930), .B1(n19963), .B2(n16724), .ZN(
        U367) );
  INV_X1 U20004 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n18928) );
  INV_X1 U20005 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n19961) );
  AOI22_X1 U20006 ( .A1(n16723), .A2(n18928), .B1(n19961), .B2(n16724), .ZN(
        U368) );
  INV_X1 U20007 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n18925) );
  INV_X1 U20008 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n19960) );
  AOI22_X1 U20009 ( .A1(n16723), .A2(n18925), .B1(n19960), .B2(n16724), .ZN(
        U369) );
  INV_X1 U20010 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n18924) );
  INV_X1 U20011 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n19958) );
  AOI22_X1 U20012 ( .A1(n16723), .A2(n18924), .B1(n19958), .B2(n16724), .ZN(
        U370) );
  INV_X1 U20013 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n18922) );
  INV_X1 U20014 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n19957) );
  AOI22_X1 U20015 ( .A1(n16722), .A2(n18922), .B1(n19957), .B2(n16724), .ZN(
        U371) );
  INV_X1 U20016 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n21129) );
  INV_X1 U20017 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n19955) );
  AOI22_X1 U20018 ( .A1(n16723), .A2(n21129), .B1(n19955), .B2(n16724), .ZN(
        U372) );
  INV_X1 U20019 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n18920) );
  INV_X1 U20020 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n19954) );
  AOI22_X1 U20021 ( .A1(n16722), .A2(n18920), .B1(n19954), .B2(n16724), .ZN(
        U373) );
  INV_X1 U20022 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n21302) );
  INV_X1 U20023 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n19953) );
  AOI22_X1 U20024 ( .A1(n16722), .A2(n21302), .B1(n19953), .B2(n16724), .ZN(
        U374) );
  INV_X1 U20025 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n18917) );
  INV_X1 U20026 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n19951) );
  AOI22_X1 U20027 ( .A1(n16722), .A2(n18917), .B1(n19951), .B2(n16724), .ZN(
        U375) );
  INV_X1 U20028 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n18898) );
  INV_X1 U20029 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n19935) );
  AOI22_X1 U20030 ( .A1(n16723), .A2(n18898), .B1(n19935), .B2(n16724), .ZN(
        U376) );
  INV_X1 U20031 ( .A(P3_ADS_N_REG_SCAN_IN), .ZN(n16725) );
  NAND2_X1 U20032 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(n18897), .ZN(n18888) );
  OR2_X1 U20033 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(P3_STATE_REG_1__SCAN_IN), 
        .ZN(n18881) );
  OAI21_X1 U20034 ( .B1(n18894), .B2(n18888), .A(n18881), .ZN(n18964) );
  OAI21_X1 U20035 ( .B1(n18894), .B2(n16725), .A(n18879), .ZN(P3_U2633) );
  INV_X1 U20036 ( .A(P3_CODEFETCH_REG_SCAN_IN), .ZN(n21272) );
  NAND2_X1 U20037 ( .A1(n16732), .A2(n16731), .ZN(n16727) );
  NAND3_X1 U20038 ( .A1(n18870), .A2(n19027), .A3(n18967), .ZN(n16726) );
  OAI221_X1 U20039 ( .B1(n21272), .B2(n17631), .C1(n21272), .C2(n16727), .A(
        n16726), .ZN(P3_U2634) );
  AOI22_X1 U20040 ( .A1(n18960), .A2(n21272), .B1(P3_D_C_N_REG_SCAN_IN), .B2(
        n19025), .ZN(n16728) );
  OAI21_X1 U20041 ( .B1(P3_STATE_REG_2__SCAN_IN), .B2(n18881), .A(n16728), 
        .ZN(P3_U2635) );
  NOR2_X1 U20042 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(P3_STATE_REG_2__SCAN_IN), 
        .ZN(n18880) );
  OAI21_X1 U20043 ( .B1(n18880), .B2(BS16), .A(n18964), .ZN(n18963) );
  OAI21_X1 U20044 ( .B1(n18964), .B2(n19013), .A(n18963), .ZN(P3_U2636) );
  INV_X1 U20045 ( .A(n16729), .ZN(n16730) );
  AOI211_X1 U20046 ( .C1(n16732), .C2(n16731), .A(n16730), .B(n18802), .ZN(
        n18809) );
  NOR2_X1 U20047 ( .A1(n18809), .A2(n18864), .ZN(n19009) );
  OAI21_X1 U20048 ( .B1(n19009), .B2(n18369), .A(n16733), .ZN(P3_U2637) );
  NOR4_X1 U20049 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_21__SCAN_IN), .A3(P3_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_23__SCAN_IN), .ZN(n16737) );
  NOR4_X1 U20050 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_16__SCAN_IN), .A3(P3_DATAWIDTH_REG_17__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_18__SCAN_IN), .ZN(n16736) );
  NOR4_X1 U20051 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_29__SCAN_IN), .A3(P3_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_31__SCAN_IN), .ZN(n16735) );
  NOR4_X1 U20052 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_25__SCAN_IN), .A3(P3_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_27__SCAN_IN), .ZN(n16734) );
  NAND4_X1 U20053 ( .A1(n16737), .A2(n16736), .A3(n16735), .A4(n16734), .ZN(
        n16743) );
  NOR4_X1 U20054 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_3__SCAN_IN), .A3(P3_DATAWIDTH_REG_4__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_5__SCAN_IN), .ZN(n16741) );
  AOI211_X1 U20055 ( .C1(P3_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_6__SCAN_IN), .B(
        P3_DATAWIDTH_REG_20__SCAN_IN), .ZN(n16740) );
  NOR4_X1 U20056 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_12__SCAN_IN), .A3(P3_DATAWIDTH_REG_13__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_14__SCAN_IN), .ZN(n16739) );
  NOR4_X1 U20057 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_8__SCAN_IN), .A3(P3_DATAWIDTH_REG_9__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_10__SCAN_IN), .ZN(n16738) );
  NAND4_X1 U20058 ( .A1(n16741), .A2(n16740), .A3(n16739), .A4(n16738), .ZN(
        n16742) );
  NOR2_X1 U20059 ( .A1(n16743), .A2(n16742), .ZN(n19003) );
  INV_X1 U20060 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n18959) );
  NOR3_X1 U20061 ( .A1(P3_DATAWIDTH_REG_1__SCAN_IN), .A2(
        P3_REIP_REG_0__SCAN_IN), .A3(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(n16745)
         );
  OAI21_X1 U20062 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(n16745), .A(n19003), .ZN(
        n16744) );
  OAI21_X1 U20063 ( .B1(n19003), .B2(n18959), .A(n16744), .ZN(P3_U2638) );
  INV_X1 U20064 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n18999) );
  INV_X1 U20065 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n21109) );
  AOI21_X1 U20066 ( .B1(n18999), .B2(n21109), .A(n16745), .ZN(n16746) );
  INV_X1 U20067 ( .A(P3_BYTEENABLE_REG_3__SCAN_IN), .ZN(n18956) );
  INV_X1 U20068 ( .A(n19003), .ZN(n19006) );
  AOI22_X1 U20069 ( .A1(n19003), .A2(n16746), .B1(n18956), .B2(n19006), .ZN(
        P3_U2639) );
  NAND2_X1 U20070 ( .A1(n16800), .A2(n17120), .ZN(n16799) );
  NOR2_X1 U20071 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n16799), .ZN(n16784) );
  INV_X1 U20072 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n17159) );
  NAND2_X1 U20073 ( .A1(n16784), .A2(n17159), .ZN(n16763) );
  NOR2_X1 U20074 ( .A1(n17110), .A2(n16763), .ZN(n16766) );
  INV_X1 U20075 ( .A(n16766), .ZN(n16762) );
  INV_X1 U20076 ( .A(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n16792) );
  NAND2_X1 U20077 ( .A1(n16749), .A2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n16748) );
  AOI21_X1 U20078 ( .B1(n16792), .B2(n16748), .A(n16747), .ZN(n17692) );
  OAI21_X1 U20079 ( .B1(n16749), .B2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n16748), .ZN(n17711) );
  INV_X1 U20080 ( .A(n17711), .ZN(n16795) );
  OAI21_X1 U20081 ( .B1(n16751), .B2(n17068), .A(n16750), .ZN(n16794) );
  NOR2_X1 U20082 ( .A1(n16793), .A2(n17068), .ZN(n16786) );
  NOR2_X1 U20083 ( .A1(n17692), .A2(n16786), .ZN(n16785) );
  NOR2_X1 U20084 ( .A1(n16785), .A2(n17068), .ZN(n16775) );
  NOR2_X1 U20085 ( .A1(n16774), .A2(n17068), .ZN(n16764) );
  NOR4_X1 U20086 ( .A1(n16765), .A2(n16764), .A3(n17068), .A4(n18873), .ZN(
        n16756) );
  NAND2_X1 U20087 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .ZN(n16770) );
  INV_X1 U20088 ( .A(n16770), .ZN(n16782) );
  NAND3_X1 U20089 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(n16782), .A3(n16798), 
        .ZN(n16759) );
  NAND2_X1 U20090 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n18951), .ZN(n16753) );
  OAI22_X1 U20091 ( .A1(n16754), .A2(n17102), .B1(n16759), .B2(n16753), .ZN(
        n16755) );
  AOI211_X1 U20092 ( .C1(n17059), .C2(P3_EBX_REG_31__SCAN_IN), .A(n16756), .B(
        n16755), .ZN(n16761) );
  INV_X1 U20093 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n18949) );
  NOR2_X1 U20094 ( .A1(n18949), .A2(n16770), .ZN(n16757) );
  AOI21_X1 U20095 ( .B1(n16758), .B2(n16757), .A(n16909), .ZN(n16779) );
  NOR2_X1 U20096 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n16759), .ZN(n16767) );
  OAI21_X1 U20097 ( .B1(n16779), .B2(n16767), .A(P3_REIP_REG_31__SCAN_IN), 
        .ZN(n16760) );
  OAI211_X1 U20098 ( .C1(P3_EBX_REG_30__SCAN_IN), .C2(n16762), .A(n16761), .B(
        n16760), .ZN(P3_U2640) );
  NAND2_X1 U20099 ( .A1(n17086), .A2(n16763), .ZN(n16772) );
  AOI21_X1 U20100 ( .B1(P3_REIP_REG_30__SCAN_IN), .B2(n16779), .A(n16767), 
        .ZN(n16768) );
  NOR2_X1 U20101 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(n16770), .ZN(n16771) );
  AOI22_X1 U20102 ( .A1(n17059), .A2(P3_EBX_REG_29__SCAN_IN), .B1(n16798), 
        .B2(n16771), .ZN(n16781) );
  INV_X1 U20103 ( .A(n16784), .ZN(n16773) );
  AOI21_X1 U20104 ( .B1(P3_EBX_REG_29__SCAN_IN), .B2(n16773), .A(n16772), .ZN(
        n16778) );
  AOI211_X1 U20105 ( .C1(n16776), .C2(n16775), .A(n16774), .B(n18873), .ZN(
        n16777) );
  AOI211_X1 U20106 ( .C1(n16779), .C2(P3_REIP_REG_29__SCAN_IN), .A(n16778), 
        .B(n16777), .ZN(n16780) );
  OAI211_X1 U20107 ( .C1(n10099), .C2(n17102), .A(n16781), .B(n16780), .ZN(
        P3_U2642) );
  INV_X1 U20108 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n18945) );
  AOI21_X1 U20109 ( .B1(n18948), .B2(n18945), .A(n16782), .ZN(n16783) );
  AOI22_X1 U20110 ( .A1(n17059), .A2(P3_EBX_REG_28__SCAN_IN), .B1(n16798), 
        .B2(n16783), .ZN(n16791) );
  AOI211_X1 U20111 ( .C1(P3_EBX_REG_28__SCAN_IN), .C2(n16799), .A(n16784), .B(
        n17110), .ZN(n16788) );
  AOI211_X1 U20112 ( .C1(n17692), .C2(n16786), .A(n16785), .B(n18873), .ZN(
        n16787) );
  AOI211_X1 U20113 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(n16789), .A(n16788), 
        .B(n16787), .ZN(n16790) );
  OAI211_X1 U20114 ( .C1(n16792), .C2(n17102), .A(n16791), .B(n16790), .ZN(
        P3_U2643) );
  AOI211_X1 U20115 ( .C1(n16795), .C2(n16794), .A(n16793), .B(n18873), .ZN(
        n16797) );
  INV_X1 U20116 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n17714) );
  OAI22_X1 U20117 ( .A1(n17714), .A2(n17102), .B1(n17111), .B2(n17120), .ZN(
        n16796) );
  AOI211_X1 U20118 ( .C1(n16798), .C2(n18945), .A(n16797), .B(n16796), .ZN(
        n16802) );
  OAI211_X1 U20119 ( .C1(n16800), .C2(n17120), .A(n17086), .B(n16799), .ZN(
        n16801) );
  OAI211_X1 U20120 ( .C1(n16803), .C2(n18945), .A(n16802), .B(n16801), .ZN(
        P3_U2644) );
  OAI22_X1 U20121 ( .A1(P3_REIP_REG_25__SCAN_IN), .A2(n16804), .B1(n16807), 
        .B2(n17111), .ZN(n16805) );
  AOI21_X1 U20122 ( .B1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n17070), .A(
        n16805), .ZN(n16815) );
  OAI211_X1 U20123 ( .C1(n16817), .C2(n16807), .A(n17086), .B(n16806), .ZN(
        n16814) );
  NAND2_X1 U20124 ( .A1(n16808), .A2(n17114), .ZN(n16876) );
  AOI21_X1 U20125 ( .B1(n16809), .B2(n16934), .A(n16909), .ZN(n16816) );
  NOR2_X1 U20126 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n17104), .ZN(n16818) );
  OAI21_X1 U20127 ( .B1(n16816), .B2(n16818), .A(P3_REIP_REG_25__SCAN_IN), 
        .ZN(n16813) );
  INV_X1 U20128 ( .A(n18873), .ZN(n17094) );
  OAI211_X1 U20129 ( .C1(n17739), .C2(n16811), .A(n17094), .B(n16810), .ZN(
        n16812) );
  NAND4_X1 U20130 ( .A1(n16815), .A2(n16814), .A3(n16813), .A4(n16812), .ZN(
        P3_U2646) );
  INV_X1 U20131 ( .A(n16816), .ZN(n16829) );
  AOI211_X1 U20132 ( .C1(P3_EBX_REG_24__SCAN_IN), .C2(n16832), .A(n16817), .B(
        n17110), .ZN(n16822) );
  INV_X1 U20133 ( .A(n16818), .ZN(n16819) );
  OAI22_X1 U20134 ( .A1(n17111), .A2(n21285), .B1(n16820), .B2(n16819), .ZN(
        n16821) );
  AOI211_X1 U20135 ( .C1(n17070), .C2(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n16822), .B(n16821), .ZN(n16826) );
  OAI211_X1 U20136 ( .C1(n17750), .C2(n16824), .A(n17094), .B(n16823), .ZN(
        n16825) );
  OAI211_X1 U20137 ( .C1(n16829), .C2(n18939), .A(n16826), .B(n16825), .ZN(
        P3_U2647) );
  INV_X1 U20138 ( .A(n16927), .ZN(n16860) );
  NOR3_X1 U20139 ( .A1(P3_REIP_REG_23__SCAN_IN), .A2(n16828), .A3(n16860), 
        .ZN(n16831) );
  OAI22_X1 U20140 ( .A1(n18938), .A2(n16829), .B1(n17111), .B2(n17119), .ZN(
        n16830) );
  AOI211_X1 U20141 ( .C1(n17070), .C2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n16831), .B(n16830), .ZN(n16838) );
  OAI211_X1 U20142 ( .C1(n16840), .C2(n17119), .A(n17086), .B(n16832), .ZN(
        n16837) );
  OAI211_X1 U20143 ( .C1(n16835), .C2(n16834), .A(n17094), .B(n16833), .ZN(
        n16836) );
  NAND3_X1 U20144 ( .A1(n16838), .A2(n16837), .A3(n16836), .ZN(P3_U2648) );
  INV_X1 U20145 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n18933) );
  INV_X1 U20146 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n18935) );
  AOI22_X1 U20147 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(n18933), .B1(
        P3_REIP_REG_21__SCAN_IN), .B2(n18935), .ZN(n16849) );
  NAND2_X1 U20148 ( .A1(n16839), .A2(n16927), .ZN(n16850) );
  AOI21_X1 U20149 ( .B1(n16839), .B2(n16934), .A(n16909), .ZN(n16859) );
  AOI211_X1 U20150 ( .C1(P3_EBX_REG_22__SCAN_IN), .C2(n16854), .A(n16840), .B(
        n17110), .ZN(n16843) );
  OAI22_X1 U20151 ( .A1(n16841), .A2(n17102), .B1(n17111), .B2(n17118), .ZN(
        n16842) );
  AOI211_X1 U20152 ( .C1(n16859), .C2(P3_REIP_REG_22__SCAN_IN), .A(n16843), 
        .B(n16842), .ZN(n16848) );
  OAI211_X1 U20153 ( .C1(n16846), .C2(n16845), .A(n17094), .B(n16844), .ZN(
        n16847) );
  OAI211_X1 U20154 ( .C1(n16849), .C2(n16850), .A(n16848), .B(n16847), .ZN(
        P3_U2649) );
  AOI22_X1 U20155 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n17070), .B1(
        n17059), .B2(P3_EBX_REG_21__SCAN_IN), .ZN(n16858) );
  INV_X1 U20156 ( .A(n16850), .ZN(n16851) );
  AOI22_X1 U20157 ( .A1(P3_REIP_REG_21__SCAN_IN), .A2(n16859), .B1(n16851), 
        .B2(n18933), .ZN(n16857) );
  OAI211_X1 U20158 ( .C1(n17790), .C2(n16853), .A(n17094), .B(n16852), .ZN(
        n16856) );
  OAI211_X1 U20159 ( .C1(n16862), .C2(n17214), .A(n17086), .B(n16854), .ZN(
        n16855) );
  NAND4_X1 U20160 ( .A1(n16858), .A2(n16857), .A3(n16856), .A4(n16855), .ZN(
        P3_U2650) );
  INV_X1 U20161 ( .A(n16859), .ZN(n16871) );
  NAND2_X1 U20162 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(P3_REIP_REG_15__SCAN_IN), 
        .ZN(n16914) );
  NOR2_X1 U20163 ( .A1(n16914), .A2(n16860), .ZN(n16901) );
  NAND2_X1 U20164 ( .A1(P3_REIP_REG_17__SCAN_IN), .A2(n16901), .ZN(n16893) );
  NOR3_X1 U20165 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(n16861), .A3(n16893), 
        .ZN(n16866) );
  AOI211_X1 U20166 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n16874), .A(n16862), .B(
        n17110), .ZN(n16865) );
  INV_X1 U20167 ( .A(P3_EBX_REG_20__SCAN_IN), .ZN(n16863) );
  OAI22_X1 U20168 ( .A1(n17804), .A2(n17102), .B1(n17111), .B2(n16863), .ZN(
        n16864) );
  NOR3_X1 U20169 ( .A1(n16866), .A2(n16865), .A3(n16864), .ZN(n16870) );
  OAI211_X1 U20170 ( .C1(n17807), .C2(n16868), .A(n17094), .B(n16867), .ZN(
        n16869) );
  OAI211_X1 U20171 ( .C1(n16871), .C2(n18931), .A(n16870), .B(n16869), .ZN(
        P3_U2651) );
  INV_X1 U20172 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n17834) );
  NAND2_X1 U20173 ( .A1(n9922), .A2(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n17818) );
  NOR2_X1 U20174 ( .A1(n18040), .A2(n17818), .ZN(n17817) );
  INV_X1 U20175 ( .A(n17817), .ZN(n16895) );
  NOR2_X1 U20176 ( .A1(n17834), .A2(n16895), .ZN(n16883) );
  INV_X1 U20177 ( .A(n17774), .ZN(n16872) );
  OAI21_X1 U20178 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n16883), .A(
        n16872), .ZN(n17821) );
  AOI21_X1 U20179 ( .B1(n16883), .B2(n17069), .A(n17068), .ZN(n16873) );
  XOR2_X1 U20180 ( .A(n17821), .B(n16873), .Z(n16882) );
  OAI211_X1 U20181 ( .C1(n16887), .C2(n21148), .A(n17086), .B(n16874), .ZN(
        n16875) );
  OAI211_X1 U20182 ( .C1(n17111), .C2(n21148), .A(n18316), .B(n16875), .ZN(
        n16880) );
  INV_X1 U20183 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n18929) );
  XOR2_X1 U20184 ( .A(n18929), .B(P3_REIP_REG_18__SCAN_IN), .Z(n16878) );
  INV_X1 U20185 ( .A(n16909), .ZN(n17112) );
  OAI21_X1 U20186 ( .B1(n16877), .B2(n16876), .A(n17112), .ZN(n16894) );
  OAI22_X1 U20187 ( .A1(n16893), .A2(n16878), .B1(n16894), .B2(n18929), .ZN(
        n16879) );
  AOI211_X1 U20188 ( .C1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .C2(n17070), .A(
        n16880), .B(n16879), .ZN(n16881) );
  OAI21_X1 U20189 ( .B1(n18873), .B2(n16882), .A(n16881), .ZN(P3_U2652) );
  INV_X1 U20190 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n18927) );
  AOI21_X1 U20191 ( .B1(n17834), .B2(n16895), .A(n16883), .ZN(n16884) );
  INV_X1 U20192 ( .A(n16884), .ZN(n17831) );
  OAI21_X1 U20193 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16895), .A(
        n17101), .ZN(n16886) );
  OAI21_X1 U20194 ( .B1(n17831), .B2(n16886), .A(n17094), .ZN(n16885) );
  AOI21_X1 U20195 ( .B1(n17831), .B2(n16886), .A(n16885), .ZN(n16891) );
  AOI211_X1 U20196 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n16903), .A(n16887), .B(
        n17110), .ZN(n16890) );
  INV_X1 U20197 ( .A(P3_EBX_REG_18__SCAN_IN), .ZN(n16888) );
  OAI22_X1 U20198 ( .A1(n17834), .A2(n17102), .B1(n17111), .B2(n16888), .ZN(
        n16889) );
  NOR4_X1 U20199 ( .A1(n18096), .A2(n16891), .A3(n16890), .A4(n16889), .ZN(
        n16892) );
  OAI221_X1 U20200 ( .B1(P3_REIP_REG_18__SCAN_IN), .B2(n16893), .C1(n18927), 
        .C2(n16894), .A(n16892), .ZN(P3_U2653) );
  AOI22_X1 U20201 ( .A1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n17070), .B1(
        n17059), .B2(P3_EBX_REG_17__SCAN_IN), .ZN(n16907) );
  INV_X1 U20202 ( .A(n16894), .ZN(n16902) );
  INV_X1 U20203 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n18926) );
  OAI21_X1 U20204 ( .B1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n16896), .A(
        n16895), .ZN(n17842) );
  NAND2_X1 U20205 ( .A1(n17101), .A2(n16897), .ZN(n16899) );
  OAI21_X1 U20206 ( .B1(n17842), .B2(n16899), .A(n17094), .ZN(n16898) );
  AOI21_X1 U20207 ( .B1(n17842), .B2(n16899), .A(n16898), .ZN(n16900) );
  AOI221_X1 U20208 ( .B1(n16902), .B2(P3_REIP_REG_17__SCAN_IN), .C1(n16901), 
        .C2(n18926), .A(n16900), .ZN(n16906) );
  OAI211_X1 U20209 ( .C1(n16912), .C2(n16904), .A(n17086), .B(n16903), .ZN(
        n16905) );
  NAND4_X1 U20210 ( .A1(n16907), .A2(n16906), .A3(n18316), .A4(n16905), .ZN(
        P3_U2654) );
  INV_X1 U20211 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n17866) );
  NOR2_X1 U20212 ( .A1(n18040), .A2(n17856), .ZN(n17855) );
  INV_X1 U20213 ( .A(n17855), .ZN(n16936) );
  NOR2_X1 U20214 ( .A1(n17866), .A2(n16936), .ZN(n16910) );
  OAI21_X1 U20215 ( .B1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n16910), .A(
        n16908), .ZN(n17860) );
  INV_X1 U20216 ( .A(n17860), .ZN(n16920) );
  INV_X1 U20217 ( .A(n16910), .ZN(n16921) );
  NOR2_X1 U20218 ( .A1(n17068), .A2(n18873), .ZN(n16993) );
  OAI21_X1 U20219 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16921), .A(
        n16993), .ZN(n16930) );
  NOR2_X1 U20220 ( .A1(n16909), .A2(n16934), .ZN(n16937) );
  NAND2_X1 U20221 ( .A1(n16910), .A2(n17069), .ZN(n16911) );
  AOI211_X1 U20222 ( .C1(n17101), .C2(n16911), .A(n18873), .B(n17860), .ZN(
        n16918) );
  AOI211_X1 U20223 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n16922), .A(n16912), .B(
        n17110), .ZN(n16913) );
  AOI211_X1 U20224 ( .C1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .C2(n17070), .A(
        n18096), .B(n16913), .ZN(n16916) );
  OAI211_X1 U20225 ( .C1(P3_REIP_REG_16__SCAN_IN), .C2(P3_REIP_REG_15__SCAN_IN), .A(n16927), .B(n16914), .ZN(n16915) );
  OAI211_X1 U20226 ( .C1(n13994), .C2(n17111), .A(n16916), .B(n16915), .ZN(
        n16917) );
  AOI211_X1 U20227 ( .C1(P3_REIP_REG_16__SCAN_IN), .C2(n16937), .A(n16918), 
        .B(n16917), .ZN(n16919) );
  OAI21_X1 U20228 ( .B1(n16920), .B2(n16930), .A(n16919), .ZN(P3_U2655) );
  OAI21_X1 U20229 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n17855), .A(
        n16921), .ZN(n17879) );
  INV_X1 U20230 ( .A(n17879), .ZN(n16931) );
  AOI21_X1 U20231 ( .B1(n17101), .B2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A(
        n18873), .ZN(n17107) );
  OAI21_X1 U20232 ( .B1(n17855), .B2(n17068), .A(n17107), .ZN(n16929) );
  INV_X1 U20233 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n18921) );
  AOI22_X1 U20234 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n17070), .B1(
        n17059), .B2(P3_EBX_REG_15__SCAN_IN), .ZN(n16925) );
  OAI211_X1 U20235 ( .C1(n16932), .C2(n16923), .A(n17086), .B(n16922), .ZN(
        n16924) );
  NAND3_X1 U20236 ( .A1(n16925), .A2(n18316), .A3(n16924), .ZN(n16926) );
  AOI221_X1 U20237 ( .B1(n16937), .B2(P3_REIP_REG_15__SCAN_IN), .C1(n16927), 
        .C2(n18921), .A(n16926), .ZN(n16928) );
  OAI221_X1 U20238 ( .B1(n16931), .B2(n16930), .C1(n17879), .C2(n16929), .A(
        n16928), .ZN(P3_U2656) );
  AOI211_X1 U20239 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n16947), .A(n16932), .B(
        n17110), .ZN(n16933) );
  AOI21_X1 U20240 ( .B1(P3_EBX_REG_14__SCAN_IN), .B2(n17059), .A(n16933), .ZN(
        n16941) );
  NOR3_X1 U20241 ( .A1(n16934), .A2(n16942), .A3(n17104), .ZN(n16935) );
  AOI22_X1 U20242 ( .A1(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n17070), .B1(
        P3_REIP_REG_13__SCAN_IN), .B2(n16935), .ZN(n16940) );
  NAND2_X1 U20243 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17069), .ZN(
        n16991) );
  INV_X1 U20244 ( .A(n16991), .ZN(n17095) );
  AOI21_X1 U20245 ( .B1(n17882), .B2(n17095), .A(n17068), .ZN(n16946) );
  NOR3_X1 U20246 ( .A1(n18040), .A2(n17921), .A3(n17924), .ZN(n16961) );
  INV_X1 U20247 ( .A(n16961), .ZN(n17891) );
  NOR2_X1 U20248 ( .A1(n17902), .A2(n17891), .ZN(n16944) );
  OAI21_X1 U20249 ( .B1(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n16944), .A(
        n16936), .ZN(n17885) );
  XNOR2_X1 U20250 ( .A(n16946), .B(n17885), .ZN(n16938) );
  AOI22_X1 U20251 ( .A1(n17094), .A2(n16938), .B1(P3_REIP_REG_14__SCAN_IN), 
        .B2(n16937), .ZN(n16939) );
  NAND4_X1 U20252 ( .A1(n16941), .A2(n16940), .A3(n16939), .A4(n18316), .ZN(
        P3_U2657) );
  NOR2_X1 U20253 ( .A1(n17104), .A2(n16942), .ZN(n16943) );
  INV_X1 U20254 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n18919) );
  AOI22_X1 U20255 ( .A1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n17070), .B1(
        n16943), .B2(n18919), .ZN(n16955) );
  NOR2_X1 U20256 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n17104), .ZN(n16958) );
  OAI21_X1 U20257 ( .B1(n16959), .B2(n17104), .A(n17114), .ZN(n16973) );
  INV_X1 U20258 ( .A(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n16952) );
  NAND2_X1 U20259 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n16961), .ZN(
        n16960) );
  AOI21_X1 U20260 ( .B1(n16952), .B2(n16960), .A(n16944), .ZN(n17894) );
  INV_X1 U20261 ( .A(n17894), .ZN(n16945) );
  NAND3_X1 U20262 ( .A1(n17094), .A2(n16946), .A3(n16945), .ZN(n16949) );
  OAI211_X1 U20263 ( .C1(n16956), .C2(n16950), .A(n17086), .B(n16947), .ZN(
        n16948) );
  OAI211_X1 U20264 ( .C1(n16950), .C2(n17111), .A(n16949), .B(n16948), .ZN(
        n16951) );
  AOI221_X1 U20265 ( .B1(n16958), .B2(P3_REIP_REG_13__SCAN_IN), .C1(n16973), 
        .C2(P3_REIP_REG_13__SCAN_IN), .A(n16951), .ZN(n16954) );
  OAI211_X1 U20266 ( .C1(n16952), .C2(n17068), .A(n17894), .B(n17107), .ZN(
        n16953) );
  NAND4_X1 U20267 ( .A1(n16955), .A2(n16954), .A3(n18316), .A4(n16953), .ZN(
        P3_U2658) );
  AOI211_X1 U20268 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n16969), .A(n16956), .B(
        n17110), .ZN(n16957) );
  AOI21_X1 U20269 ( .B1(n17070), .B2(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n16957), .ZN(n16966) );
  AOI22_X1 U20270 ( .A1(n17059), .A2(P3_EBX_REG_12__SCAN_IN), .B1(n16959), 
        .B2(n16958), .ZN(n16965) );
  OAI21_X1 U20271 ( .B1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n16961), .A(
        n16960), .ZN(n17918) );
  OAI21_X1 U20272 ( .B1(n17900), .B2(n16991), .A(n17101), .ZN(n16962) );
  XOR2_X1 U20273 ( .A(n17918), .B(n16962), .Z(n16963) );
  AOI22_X1 U20274 ( .A1(n17094), .A2(n16963), .B1(P3_REIP_REG_12__SCAN_IN), 
        .B2(n16973), .ZN(n16964) );
  NAND4_X1 U20275 ( .A1(n16966), .A2(n16965), .A3(n16964), .A4(n18316), .ZN(
        P3_U2659) );
  INV_X1 U20276 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n18909) );
  NAND4_X1 U20277 ( .A1(n17083), .A2(P3_REIP_REG_5__SCAN_IN), .A3(n17039), 
        .A4(P3_REIP_REG_6__SCAN_IN), .ZN(n17027) );
  NOR2_X1 U20278 ( .A1(n18909), .A2(n17027), .ZN(n17006) );
  NAND2_X1 U20279 ( .A1(P3_REIP_REG_8__SCAN_IN), .A2(n17006), .ZN(n17000) );
  OAI21_X1 U20280 ( .B1(n16967), .B2(n17000), .A(n18916), .ZN(n16974) );
  NOR2_X1 U20281 ( .A1(n18040), .A2(n17921), .ZN(n16981) );
  OAI21_X1 U20282 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n16981), .A(
        n17891), .ZN(n17922) );
  OAI21_X1 U20283 ( .B1(n17921), .B2(n16991), .A(n17101), .ZN(n16983) );
  AOI21_X1 U20284 ( .B1(n17922), .B2(n16983), .A(n18873), .ZN(n16968) );
  OAI21_X1 U20285 ( .B1(n17922), .B2(n16983), .A(n16968), .ZN(n16971) );
  OAI211_X1 U20286 ( .C1(n16976), .C2(n17322), .A(n17086), .B(n16969), .ZN(
        n16970) );
  OAI211_X1 U20287 ( .C1(n17102), .C2(n17924), .A(n16971), .B(n16970), .ZN(
        n16972) );
  AOI21_X1 U20288 ( .B1(n16974), .B2(n16973), .A(n16972), .ZN(n16975) );
  OAI211_X1 U20289 ( .C1(n17111), .C2(n17322), .A(n16975), .B(n18316), .ZN(
        P3_U2660) );
  INV_X1 U20290 ( .A(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n16990) );
  AOI211_X1 U20291 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n16977), .A(n16976), .B(
        n17110), .ZN(n16978) );
  AOI211_X1 U20292 ( .C1(n17059), .C2(P3_EBX_REG_10__SCAN_IN), .A(n18096), .B(
        n16978), .ZN(n16989) );
  INV_X1 U20293 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n18912) );
  NOR2_X1 U20294 ( .A1(n18912), .A2(n17000), .ZN(n16987) );
  INV_X1 U20295 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n18914) );
  AOI21_X1 U20296 ( .B1(n16979), .B2(n17083), .A(n17100), .ZN(n17042) );
  INV_X1 U20297 ( .A(n17042), .ZN(n17035) );
  AOI21_X1 U20298 ( .B1(n17112), .B2(n16980), .A(n17035), .ZN(n17012) );
  OAI21_X1 U20299 ( .B1(P3_REIP_REG_9__SCAN_IN), .B2(n17000), .A(n17012), .ZN(
        n16986) );
  NOR2_X1 U20300 ( .A1(n18040), .A2(n17945), .ZN(n17007) );
  NAND2_X1 U20301 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n17007), .ZN(
        n16992) );
  AOI21_X1 U20302 ( .B1(n16990), .B2(n16992), .A(n16981), .ZN(n17932) );
  INV_X1 U20303 ( .A(n17932), .ZN(n16984) );
  NAND2_X1 U20304 ( .A1(n17094), .A2(n17068), .ZN(n17098) );
  NOR2_X1 U20305 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n16992), .ZN(
        n17004) );
  OAI21_X1 U20306 ( .B1(n17004), .B2(n16984), .A(n17094), .ZN(n16982) );
  AOI22_X1 U20307 ( .A1(n16984), .A2(n16983), .B1(n17098), .B2(n16982), .ZN(
        n16985) );
  AOI221_X1 U20308 ( .B1(n16987), .B2(n18914), .C1(n16986), .C2(
        P3_REIP_REG_10__SCAN_IN), .A(n16985), .ZN(n16988) );
  OAI211_X1 U20309 ( .C1(n16990), .C2(n17102), .A(n16989), .B(n16988), .ZN(
        P3_U2661) );
  NOR2_X1 U20310 ( .A1(n18873), .A2(n16991), .ZN(n17055) );
  OAI21_X1 U20311 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n17007), .A(
        n16992), .ZN(n17947) );
  AOI22_X1 U20312 ( .A1(n16994), .A2(n17055), .B1(n16993), .B2(n17947), .ZN(
        n17003) );
  NOR3_X1 U20313 ( .A1(P3_EBX_REG_9__SCAN_IN), .A2(n17005), .A3(n17110), .ZN(
        n16999) );
  AOI21_X1 U20314 ( .B1(n17086), .B2(n17005), .A(n17059), .ZN(n16995) );
  OAI22_X1 U20315 ( .A1(n16996), .A2(n16995), .B1(n17947), .B2(n17098), .ZN(
        n16998) );
  INV_X1 U20316 ( .A(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n17931) );
  OAI22_X1 U20317 ( .A1(n17012), .A2(n18912), .B1(n17931), .B2(n17102), .ZN(
        n16997) );
  NOR4_X1 U20318 ( .A1(n18096), .A2(n16999), .A3(n16998), .A4(n16997), .ZN(
        n17002) );
  OR2_X1 U20319 ( .A1(n17000), .A2(P3_REIP_REG_9__SCAN_IN), .ZN(n17001) );
  OAI211_X1 U20320 ( .C1(n17004), .C2(n17003), .A(n17002), .B(n17001), .ZN(
        P3_U2662) );
  INV_X1 U20321 ( .A(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n17964) );
  AOI211_X1 U20322 ( .C1(P3_EBX_REG_8__SCAN_IN), .C2(n17020), .A(n17005), .B(
        n17110), .ZN(n17014) );
  NOR2_X1 U20323 ( .A1(P3_REIP_REG_8__SCAN_IN), .A2(n17006), .ZN(n17011) );
  INV_X1 U20324 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n17973) );
  NAND2_X1 U20325 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17954), .ZN(
        n17028) );
  NOR2_X1 U20326 ( .A1(n17973), .A2(n17028), .ZN(n17017) );
  INV_X1 U20327 ( .A(n17017), .ZN(n17008) );
  AOI21_X1 U20328 ( .B1(n17964), .B2(n17008), .A(n17007), .ZN(n17955) );
  AOI21_X1 U20329 ( .B1(n17017), .B2(n17069), .A(n17068), .ZN(n17009) );
  XNOR2_X1 U20330 ( .A(n17955), .B(n17009), .ZN(n17010) );
  OAI22_X1 U20331 ( .A1(n17012), .A2(n17011), .B1(n18873), .B2(n17010), .ZN(
        n17013) );
  AOI211_X1 U20332 ( .C1(P3_EBX_REG_8__SCAN_IN), .C2(n17059), .A(n17014), .B(
        n17013), .ZN(n17015) );
  OAI211_X1 U20333 ( .C1(n17964), .C2(n17102), .A(n17015), .B(n18316), .ZN(
        P3_U2663) );
  NAND3_X1 U20334 ( .A1(n17083), .A2(P3_REIP_REG_5__SCAN_IN), .A3(n17039), 
        .ZN(n17016) );
  NOR2_X1 U20335 ( .A1(P3_REIP_REG_6__SCAN_IN), .A2(n17016), .ZN(n17034) );
  NOR2_X1 U20336 ( .A1(n17035), .A2(n17034), .ZN(n17026) );
  AOI21_X1 U20337 ( .B1(n17973), .B2(n17028), .A(n17017), .ZN(n17979) );
  INV_X1 U20338 ( .A(n17028), .ZN(n17018) );
  AOI21_X1 U20339 ( .B1(n17018), .B2(n17069), .A(n17068), .ZN(n17032) );
  OAI21_X1 U20340 ( .B1(n17979), .B2(n17032), .A(n17094), .ZN(n17019) );
  AOI21_X1 U20341 ( .B1(n17979), .B2(n17032), .A(n17019), .ZN(n17024) );
  OAI211_X1 U20342 ( .C1(n17029), .C2(n17022), .A(n17086), .B(n17020), .ZN(
        n17021) );
  OAI211_X1 U20343 ( .C1(n17111), .C2(n17022), .A(n18316), .B(n17021), .ZN(
        n17023) );
  AOI211_X1 U20344 ( .C1(n17070), .C2(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A(
        n17024), .B(n17023), .ZN(n17025) );
  OAI221_X1 U20345 ( .B1(P3_REIP_REG_7__SCAN_IN), .B2(n17027), .C1(n18909), 
        .C2(n17026), .A(n17025), .ZN(P3_U2664) );
  NOR2_X1 U20346 ( .A1(n18040), .A2(n17971), .ZN(n17040) );
  OAI21_X1 U20347 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n17040), .A(
        n17028), .ZN(n17985) );
  OAI21_X1 U20348 ( .B1(n17989), .B2(n17068), .A(n17107), .ZN(n17038) );
  AOI211_X1 U20349 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n17045), .A(n17029), .B(
        n17110), .ZN(n17031) );
  OAI22_X1 U20350 ( .A1(n17989), .A2(n17102), .B1(n17111), .B2(n21274), .ZN(
        n17030) );
  NOR3_X1 U20351 ( .A1(n18096), .A2(n17031), .A3(n17030), .ZN(n17037) );
  AND3_X1 U20352 ( .A1(n17094), .A2(n17032), .A3(n17985), .ZN(n17033) );
  AOI211_X1 U20353 ( .C1(n17035), .C2(P3_REIP_REG_6__SCAN_IN), .A(n17034), .B(
        n17033), .ZN(n17036) );
  OAI211_X1 U20354 ( .C1(n17985), .C2(n17038), .A(n17037), .B(n17036), .ZN(
        P3_U2665) );
  INV_X1 U20355 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n17049) );
  AOI21_X1 U20356 ( .B1(n17083), .B2(n17039), .A(P3_REIP_REG_5__SCAN_IN), .ZN(
        n17043) );
  NAND2_X1 U20357 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17993), .ZN(
        n17050) );
  AOI21_X1 U20358 ( .B1(n17049), .B2(n17050), .A(n17040), .ZN(n18001) );
  AOI21_X1 U20359 ( .B1(n17993), .B2(n17095), .A(n17068), .ZN(n17060) );
  XNOR2_X1 U20360 ( .A(n18001), .B(n17060), .ZN(n17041) );
  OAI22_X1 U20361 ( .A1(n17043), .A2(n17042), .B1(n18873), .B2(n17041), .ZN(
        n17044) );
  AOI211_X1 U20362 ( .C1(n17059), .C2(P3_EBX_REG_5__SCAN_IN), .A(n18096), .B(
        n17044), .ZN(n17048) );
  OAI211_X1 U20363 ( .C1(n17053), .C2(n17046), .A(n17086), .B(n17045), .ZN(
        n17047) );
  OAI211_X1 U20364 ( .C1(n17102), .C2(n17049), .A(n17048), .B(n17047), .ZN(
        P3_U2666) );
  NOR2_X1 U20365 ( .A1(n18040), .A2(n17052), .ZN(n17066) );
  OAI21_X1 U20366 ( .B1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n17066), .A(
        n17050), .ZN(n18010) );
  NOR2_X1 U20367 ( .A1(n18378), .A2(n17051), .ZN(n19032) );
  INV_X1 U20368 ( .A(n19032), .ZN(n17117) );
  NOR2_X1 U20369 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n17052), .ZN(
        n18005) );
  AOI211_X1 U20370 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n17076), .A(n17053), .B(
        n17110), .ZN(n17054) );
  AOI211_X1 U20371 ( .C1(n18005), .C2(n17055), .A(n18096), .B(n17054), .ZN(
        n17056) );
  OAI221_X1 U20372 ( .B1(n17117), .B2(n17384), .C1(n17117), .C2(n18812), .A(
        n17056), .ZN(n17064) );
  AOI21_X1 U20373 ( .B1(n17083), .B2(n17057), .A(n17100), .ZN(n17072) );
  NOR3_X1 U20374 ( .A1(P3_REIP_REG_4__SCAN_IN), .A2(n17104), .A3(n17057), .ZN(
        n17058) );
  AOI21_X1 U20375 ( .B1(P3_EBX_REG_4__SCAN_IN), .B2(n17059), .A(n17058), .ZN(
        n17062) );
  NAND3_X1 U20376 ( .A1(n17094), .A2(n17060), .A3(n18010), .ZN(n17061) );
  OAI211_X1 U20377 ( .C1(n17072), .C2(n18903), .A(n17062), .B(n17061), .ZN(
        n17063) );
  AOI211_X1 U20378 ( .C1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .C2(n17070), .A(
        n17064), .B(n17063), .ZN(n17065) );
  OAI21_X1 U20379 ( .B1(n17098), .B2(n18010), .A(n17065), .ZN(P3_U2667) );
  INV_X1 U20380 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n18033) );
  NOR2_X1 U20381 ( .A1(n18040), .A2(n18033), .ZN(n17080) );
  INV_X1 U20382 ( .A(n17066), .ZN(n17067) );
  OAI21_X1 U20383 ( .B1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n17080), .A(
        n17067), .ZN(n18019) );
  AOI21_X1 U20384 ( .B1(n17080), .B2(n17069), .A(n17068), .ZN(n17093) );
  XNOR2_X1 U20385 ( .A(n18019), .B(n17093), .ZN(n17075) );
  NAND3_X1 U20386 ( .A1(n17083), .A2(P3_REIP_REG_1__SCAN_IN), .A3(
        P3_REIP_REG_2__SCAN_IN), .ZN(n17073) );
  INV_X1 U20387 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n18901) );
  NAND2_X1 U20388 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18838), .ZN(
        n18834) );
  AOI21_X1 U20389 ( .B1(n18972), .B2(n18834), .A(n17327), .ZN(n18968) );
  AOI22_X1 U20390 ( .A1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n17070), .B1(
        n19032), .B2(n18968), .ZN(n17071) );
  OAI221_X1 U20391 ( .B1(P3_REIP_REG_3__SCAN_IN), .B2(n17073), .C1(n18901), 
        .C2(n17072), .A(n17071), .ZN(n17074) );
  AOI21_X1 U20392 ( .B1(n17075), .B2(n17094), .A(n17074), .ZN(n17078) );
  OAI211_X1 U20393 ( .C1(n17084), .C2(n17079), .A(n17086), .B(n17076), .ZN(
        n17077) );
  OAI211_X1 U20394 ( .C1(n17079), .C2(n17111), .A(n17078), .B(n17077), .ZN(
        P3_U2668) );
  AOI21_X1 U20395 ( .B1(n18040), .B2(n18033), .A(n17080), .ZN(n17081) );
  INV_X1 U20396 ( .A(n17081), .ZN(n18030) );
  INV_X1 U20397 ( .A(P3_EBX_REG_2__SCAN_IN), .ZN(n17087) );
  OAI22_X1 U20398 ( .A1(n18033), .A2(n17102), .B1(n17111), .B2(n17087), .ZN(
        n17092) );
  NAND2_X1 U20399 ( .A1(n18982), .A2(n18840), .ZN(n18830) );
  NAND2_X1 U20400 ( .A1(n18834), .A2(n18830), .ZN(n18978) );
  NAND2_X1 U20401 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_2__SCAN_IN), 
        .ZN(n17082) );
  OAI211_X1 U20402 ( .C1(P3_REIP_REG_1__SCAN_IN), .C2(P3_REIP_REG_2__SCAN_IN), 
        .A(n17083), .B(n17082), .ZN(n17090) );
  NOR2_X1 U20403 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n17088) );
  INV_X1 U20404 ( .A(n17084), .ZN(n17085) );
  OAI211_X1 U20405 ( .C1(n17088), .C2(n17087), .A(n17086), .B(n17085), .ZN(
        n17089) );
  OAI211_X1 U20406 ( .C1(n17117), .C2(n18978), .A(n17090), .B(n17089), .ZN(
        n17091) );
  AOI211_X1 U20407 ( .C1(n17100), .C2(P3_REIP_REG_2__SCAN_IN), .A(n17092), .B(
        n17091), .ZN(n17097) );
  OAI211_X1 U20408 ( .C1(n17095), .C2(n18030), .A(n17094), .B(n17093), .ZN(
        n17096) );
  OAI211_X1 U20409 ( .C1(n18030), .C2(n17098), .A(n17097), .B(n17096), .ZN(
        P3_U2669) );
  NAND2_X1 U20410 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n17417) );
  OAI21_X1 U20411 ( .B1(P3_EBX_REG_0__SCAN_IN), .B2(P3_EBX_REG_1__SCAN_IN), 
        .A(n17417), .ZN(n17424) );
  INV_X1 U20412 ( .A(n18840), .ZN(n18817) );
  NOR2_X1 U20413 ( .A1(n17099), .A2(n18817), .ZN(n18987) );
  AOI22_X1 U20414 ( .A1(n17100), .A2(P3_REIP_REG_1__SCAN_IN), .B1(n18987), 
        .B2(n19032), .ZN(n17109) );
  NAND2_X1 U20415 ( .A1(n17101), .A2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n17103) );
  OAI21_X1 U20416 ( .B1(n18873), .B2(n17103), .A(n17102), .ZN(n17106) );
  INV_X1 U20417 ( .A(P3_EBX_REG_1__SCAN_IN), .ZN(n17423) );
  OAI22_X1 U20418 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n17104), .B1(n17111), 
        .B2(n17423), .ZN(n17105) );
  AOI221_X1 U20419 ( .B1(n17107), .B2(n18040), .C1(n17106), .C2(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A(n17105), .ZN(n17108) );
  OAI211_X1 U20420 ( .C1(n17110), .C2(n17424), .A(n17109), .B(n17108), .ZN(
        P3_U2670) );
  NAND2_X1 U20421 ( .A1(n17111), .A2(n17110), .ZN(n17113) );
  AOI22_X1 U20422 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(n17113), .B1(
        P3_REIP_REG_0__SCAN_IN), .B2(n17112), .ZN(n17116) );
  INV_X1 U20423 ( .A(n19028), .ZN(n18993) );
  NAND3_X1 U20424 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n18993), .A3(
        n17114), .ZN(n17115) );
  OAI211_X1 U20425 ( .C1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .C2(n17117), .A(
        n17116), .B(n17115), .ZN(P3_U2671) );
  INV_X1 U20426 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n17127) );
  NOR4_X1 U20427 ( .A1(n21285), .A2(n17119), .A3(n17118), .A4(n17214), .ZN(
        n17123) );
  NOR4_X1 U20428 ( .A1(n17159), .A2(n17121), .A3(n17120), .A4(n17198), .ZN(
        n17122) );
  NAND4_X1 U20429 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(P3_EBX_REG_25__SCAN_IN), 
        .A3(n17123), .A4(n17122), .ZN(n17126) );
  NAND2_X1 U20430 ( .A1(n17418), .A2(P3_EBX_REG_31__SCAN_IN), .ZN(n17125) );
  NAND2_X1 U20431 ( .A1(n17154), .A2(n17547), .ZN(n17124) );
  OAI22_X1 U20432 ( .A1(n17154), .A2(n17125), .B1(P3_EBX_REG_31__SCAN_IN), 
        .B2(n17124), .ZN(P3_U2672) );
  NAND2_X1 U20433 ( .A1(n17127), .A2(n17126), .ZN(n17128) );
  NAND2_X1 U20434 ( .A1(n17128), .A2(n17418), .ZN(n17153) );
  INV_X1 U20435 ( .A(n17163), .ZN(n17155) );
  AOI22_X1 U20436 ( .A1(n17245), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n9829), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n17139) );
  INV_X1 U20437 ( .A(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n17131) );
  AOI22_X1 U20438 ( .A1(n17357), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17343), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n17130) );
  AOI22_X1 U20439 ( .A1(n17309), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n17385), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n17129) );
  OAI211_X1 U20440 ( .C1(n13050), .C2(n17131), .A(n17130), .B(n17129), .ZN(
        n17137) );
  AOI22_X1 U20441 ( .A1(n12552), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n17379), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n17135) );
  AOI22_X1 U20442 ( .A1(n13120), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17365), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n17134) );
  AOI22_X1 U20443 ( .A1(n13079), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n13089), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n17133) );
  NAND2_X1 U20444 ( .A1(n17344), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n17132) );
  NAND4_X1 U20445 ( .A1(n17135), .A2(n17134), .A3(n17133), .A4(n17132), .ZN(
        n17136) );
  AOI211_X1 U20446 ( .C1(n17327), .C2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A(
        n17137), .B(n17136), .ZN(n17138) );
  OAI211_X1 U20447 ( .C1(n17395), .C2(n21237), .A(n17139), .B(n17138), .ZN(
        n17158) );
  NAND3_X1 U20448 ( .A1(n17156), .A2(n17155), .A3(n17158), .ZN(n17152) );
  AOI22_X1 U20449 ( .A1(n17357), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n17365), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n17140) );
  OAI21_X1 U20450 ( .B1(n12537), .B2(n21152), .A(n17140), .ZN(n17150) );
  AOI22_X1 U20451 ( .A1(n17379), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n9829), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n17148) );
  AOI22_X1 U20452 ( .A1(n17344), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n13089), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n17141) );
  OAI21_X1 U20453 ( .B1(n13050), .B2(n17273), .A(n17141), .ZN(n17146) );
  AOI22_X1 U20454 ( .A1(n17385), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n17343), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n17143) );
  AOI22_X1 U20455 ( .A1(n12552), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n13120), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n17142) );
  OAI211_X1 U20456 ( .C1(n17384), .C2(n17144), .A(n17143), .B(n17142), .ZN(
        n17145) );
  AOI211_X1 U20457 ( .C1(n13079), .C2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A(
        n17146), .B(n17145), .ZN(n17147) );
  OAI211_X1 U20458 ( .C1(n17395), .C2(n17277), .A(n17148), .B(n17147), .ZN(
        n17149) );
  AOI211_X1 U20459 ( .C1(n17378), .C2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A(
        n17150), .B(n17149), .ZN(n17151) );
  XNOR2_X1 U20460 ( .A(n17152), .B(n17151), .ZN(n17439) );
  OAI22_X1 U20461 ( .A1(n17154), .A2(n17153), .B1(n17439), .B2(n17418), .ZN(
        P3_U2673) );
  NAND2_X1 U20462 ( .A1(n17156), .A2(n17155), .ZN(n17157) );
  XOR2_X1 U20463 ( .A(n17158), .B(n17157), .Z(n17444) );
  AOI22_X1 U20464 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n17161), .B1(n17160), 
        .B2(n17159), .ZN(n17162) );
  OAI21_X1 U20465 ( .B1(n17418), .B2(n17444), .A(n17162), .ZN(P3_U2674) );
  OAI21_X1 U20466 ( .B1(n17165), .B2(n17164), .A(n17163), .ZN(n17453) );
  NAND3_X1 U20467 ( .A1(n9895), .A2(P3_EBX_REG_27__SCAN_IN), .A3(n17418), .ZN(
        n17166) );
  OAI221_X1 U20468 ( .B1(n9895), .B2(P3_EBX_REG_27__SCAN_IN), .C1(n17418), 
        .C2(n17453), .A(n17166), .ZN(P3_U2676) );
  AOI21_X1 U20469 ( .B1(P3_EBX_REG_26__SCAN_IN), .B2(n17418), .A(n17174), .ZN(
        n17168) );
  XNOR2_X1 U20470 ( .A(n17167), .B(n17170), .ZN(n17458) );
  OAI22_X1 U20471 ( .A1(n17169), .A2(n17168), .B1(n17418), .B2(n17458), .ZN(
        P3_U2677) );
  AOI21_X1 U20472 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n17418), .A(n17178), .ZN(
        n17173) );
  OAI21_X1 U20473 ( .B1(n17172), .B2(n17171), .A(n17170), .ZN(n17462) );
  OAI22_X1 U20474 ( .A1(n17174), .A2(n17173), .B1(n17418), .B2(n17462), .ZN(
        P3_U2678) );
  INV_X1 U20475 ( .A(n17175), .ZN(n17184) );
  AOI21_X1 U20476 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n17418), .A(n17184), .ZN(
        n17177) );
  XNOR2_X1 U20477 ( .A(n17176), .B(n17180), .ZN(n17467) );
  OAI22_X1 U20478 ( .A1(n17178), .A2(n17177), .B1(n17418), .B2(n17467), .ZN(
        P3_U2679) );
  AOI21_X1 U20479 ( .B1(P3_EBX_REG_23__SCAN_IN), .B2(n17418), .A(n17179), .ZN(
        n17183) );
  OAI21_X1 U20480 ( .B1(n17182), .B2(n17181), .A(n17180), .ZN(n17472) );
  OAI22_X1 U20481 ( .A1(n17184), .A2(n17183), .B1(n17418), .B2(n17472), .ZN(
        P3_U2680) );
  INV_X1 U20482 ( .A(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n17299) );
  AOI22_X1 U20483 ( .A1(n17385), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17343), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n17185) );
  OAI21_X1 U20484 ( .B1(n9919), .B2(n17299), .A(n17185), .ZN(n17195) );
  AOI22_X1 U20485 ( .A1(n17344), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n13089), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n17193) );
  OAI22_X1 U20486 ( .A1(n13051), .A2(n17186), .B1(n17395), .B2(n17290), .ZN(
        n17191) );
  AOI22_X1 U20487 ( .A1(n13120), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n9829), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n17189) );
  AOI22_X1 U20488 ( .A1(n17245), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17365), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n17188) );
  AOI22_X1 U20489 ( .A1(n17327), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17361), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n17187) );
  NAND3_X1 U20490 ( .A1(n17189), .A2(n17188), .A3(n17187), .ZN(n17190) );
  AOI211_X1 U20491 ( .C1(n17379), .C2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A(
        n17191), .B(n17190), .ZN(n17192) );
  OAI211_X1 U20492 ( .C1(n12551), .C2(n21237), .A(n17193), .B(n17192), .ZN(
        n17194) );
  AOI211_X1 U20493 ( .C1(n12552), .C2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A(
        n17195), .B(n17194), .ZN(n17476) );
  NAND3_X1 U20494 ( .A1(n17197), .A2(P3_EBX_REG_22__SCAN_IN), .A3(n17418), 
        .ZN(n17196) );
  OAI221_X1 U20495 ( .B1(n17197), .B2(P3_EBX_REG_22__SCAN_IN), .C1(n17418), 
        .C2(n17476), .A(n17196), .ZN(P3_U2681) );
  NAND2_X1 U20496 ( .A1(n17418), .A2(n17198), .ZN(n17227) );
  AOI22_X1 U20497 ( .A1(n13079), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n17361), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n17210) );
  AOI22_X1 U20498 ( .A1(n13120), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n17365), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n17199) );
  OAI21_X1 U20499 ( .B1(n9884), .B2(n17200), .A(n17199), .ZN(n17208) );
  OAI22_X1 U20500 ( .A1(n17395), .A2(n17407), .B1(n17340), .B2(n17201), .ZN(
        n17202) );
  AOI21_X1 U20501 ( .B1(n12552), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A(
        n17202), .ZN(n17206) );
  AOI22_X1 U20502 ( .A1(n17309), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17357), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n17205) );
  AOI22_X1 U20503 ( .A1(n17245), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n9829), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n17204) );
  AOI22_X1 U20504 ( .A1(n17344), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17327), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n17203) );
  NAND4_X1 U20505 ( .A1(n17206), .A2(n17205), .A3(n17204), .A4(n17203), .ZN(
        n17207) );
  AOI211_X1 U20506 ( .C1(n17379), .C2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A(
        n17208), .B(n17207), .ZN(n17209) );
  OAI211_X1 U20507 ( .C1(n9827), .C2(n17211), .A(n17210), .B(n17209), .ZN(
        n17481) );
  AOI22_X1 U20508 ( .A1(n17426), .A2(n17481), .B1(n17212), .B2(n17214), .ZN(
        n17213) );
  OAI21_X1 U20509 ( .B1(n17214), .B2(n17227), .A(n17213), .ZN(P3_U2682) );
  NOR2_X1 U20510 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n17215), .ZN(n17228) );
  AOI22_X1 U20511 ( .A1(n17245), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17365), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n17216) );
  OAI21_X1 U20512 ( .B1(n13051), .B2(n17217), .A(n17216), .ZN(n17226) );
  INV_X1 U20513 ( .A(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n17317) );
  AOI22_X1 U20514 ( .A1(n13120), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n13089), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n17224) );
  INV_X1 U20515 ( .A(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n17307) );
  OAI22_X1 U20516 ( .A1(n17395), .A2(n17411), .B1(n12551), .B2(n17307), .ZN(
        n17222) );
  AOI22_X1 U20517 ( .A1(n9829), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17343), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n17220) );
  AOI22_X1 U20518 ( .A1(n17379), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n17385), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n17219) );
  AOI22_X1 U20519 ( .A1(n17327), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17361), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n17218) );
  NAND3_X1 U20520 ( .A1(n17220), .A2(n17219), .A3(n17218), .ZN(n17221) );
  AOI211_X1 U20521 ( .C1(n17344), .C2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A(
        n17222), .B(n17221), .ZN(n17223) );
  OAI211_X1 U20522 ( .C1(n9919), .C2(n17317), .A(n17224), .B(n17223), .ZN(
        n17225) );
  AOI211_X1 U20523 ( .C1(n12552), .C2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A(
        n17226), .B(n17225), .ZN(n17489) );
  OAI22_X1 U20524 ( .A1(n17228), .A2(n17227), .B1(n17489), .B2(n17418), .ZN(
        P3_U2683) );
  NAND2_X1 U20525 ( .A1(n17418), .A2(n17239), .ZN(n17255) );
  AOI22_X1 U20526 ( .A1(n17245), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17357), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n17238) );
  AOI22_X1 U20527 ( .A1(n17309), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n17343), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n17230) );
  AOI22_X1 U20528 ( .A1(n9829), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17365), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n17229) );
  OAI211_X1 U20529 ( .C1(n17384), .C2(n21140), .A(n17230), .B(n17229), .ZN(
        n17236) );
  AOI22_X1 U20530 ( .A1(n17379), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n17385), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n17234) );
  AOI22_X1 U20531 ( .A1(n12552), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n13120), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n17233) );
  AOI22_X1 U20532 ( .A1(n13079), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n13089), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n17232) );
  NAND2_X1 U20533 ( .A1(n17344), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(
        n17231) );
  NAND4_X1 U20534 ( .A1(n17234), .A2(n17233), .A3(n17232), .A4(n17231), .ZN(
        n17235) );
  AOI211_X1 U20535 ( .C1(n17361), .C2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A(
        n17236), .B(n17235), .ZN(n17237) );
  OAI211_X1 U20536 ( .C1(n17395), .C2(n17414), .A(n17238), .B(n17237), .ZN(
        n17490) );
  NOR3_X1 U20537 ( .A1(P3_EBX_REG_19__SCAN_IN), .A2(n18413), .A3(n17239), .ZN(
        n17240) );
  AOI21_X1 U20538 ( .B1(n17426), .B2(n17490), .A(n17240), .ZN(n17241) );
  OAI21_X1 U20539 ( .B1(n21148), .B2(n17255), .A(n17241), .ZN(P3_U2684) );
  AOI22_X1 U20540 ( .A1(n9829), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n17343), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n17242) );
  OAI21_X1 U20541 ( .B1(n17360), .B2(n21293), .A(n17242), .ZN(n17254) );
  AOI22_X1 U20542 ( .A1(n13080), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n17357), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n17251) );
  INV_X1 U20543 ( .A(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n17244) );
  AOI22_X1 U20544 ( .A1(n17344), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n13089), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n17243) );
  OAI21_X1 U20545 ( .B1(n17384), .B2(n17244), .A(n17243), .ZN(n17249) );
  AOI22_X1 U20546 ( .A1(n12552), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n17245), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n17247) );
  AOI22_X1 U20547 ( .A1(n17385), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17365), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n17246) );
  OAI211_X1 U20548 ( .C1(n12551), .C2(n21306), .A(n17247), .B(n17246), .ZN(
        n17248) );
  AOI211_X1 U20549 ( .C1(n17361), .C2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A(
        n17249), .B(n17248), .ZN(n17250) );
  OAI211_X1 U20550 ( .C1(n17252), .C2(n17341), .A(n17251), .B(n17250), .ZN(
        n17253) );
  AOI211_X1 U20551 ( .C1(n17378), .C2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A(
        n17254), .B(n17253), .ZN(n17499) );
  NOR2_X1 U20552 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n17271), .ZN(n17256) );
  OAI22_X1 U20553 ( .A1(n17499), .A2(n17418), .B1(n17256), .B2(n17255), .ZN(
        P3_U2685) );
  INV_X1 U20554 ( .A(n17257), .ZN(n17258) );
  OAI21_X1 U20555 ( .B1(P3_EBX_REG_17__SCAN_IN), .B2(n17258), .A(n17418), .ZN(
        n17270) );
  AOI22_X1 U20556 ( .A1(n17378), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_11__1__SCAN_IN), .B2(n17385), .ZN(n17259) );
  OAI21_X1 U20557 ( .B1(n17359), .B2(n12561), .A(n17259), .ZN(n17269) );
  AOI22_X1 U20558 ( .A1(n17245), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n13080), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n17267) );
  AOI22_X1 U20559 ( .A1(n13079), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n13089), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n17260) );
  OAI21_X1 U20560 ( .B1(n17261), .B2(n13050), .A(n17260), .ZN(n17265) );
  AOI22_X1 U20561 ( .A1(n12552), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_6__1__SCAN_IN), .B2(n17365), .ZN(n17263) );
  AOI22_X1 U20562 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n17343), .B1(
        n13120), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n17262) );
  OAI211_X1 U20563 ( .C1(n21308), .C2(n17363), .A(n17263), .B(n17262), .ZN(
        n17264) );
  AOI211_X1 U20564 ( .C1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .C2(n17327), .A(
        n17265), .B(n17264), .ZN(n17266) );
  OAI211_X1 U20565 ( .C1(n17360), .C2(n21275), .A(n17267), .B(n17266), .ZN(
        n17268) );
  AOI211_X1 U20566 ( .C1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .C2(n17386), .A(
        n17269), .B(n17268), .ZN(n17506) );
  OAI22_X1 U20567 ( .A1(n17271), .A2(n17270), .B1(n17506), .B2(n17418), .ZN(
        P3_U2686) );
  AOI22_X1 U20568 ( .A1(n17357), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n9829), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n17272) );
  OAI21_X1 U20569 ( .B1(n17306), .B2(n17273), .A(n17272), .ZN(n17285) );
  INV_X1 U20570 ( .A(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n17282) );
  AOI22_X1 U20571 ( .A1(n13080), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n17343), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n17281) );
  AOI22_X1 U20572 ( .A1(n13089), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n17361), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n17274) );
  OAI21_X1 U20573 ( .B1(n12551), .B2(n17401), .A(n17274), .ZN(n17279) );
  AOI22_X1 U20574 ( .A1(n17309), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n13120), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n17276) );
  AOI22_X1 U20575 ( .A1(n17245), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n17385), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n17275) );
  OAI211_X1 U20576 ( .C1(n17384), .C2(n17277), .A(n17276), .B(n17275), .ZN(
        n17278) );
  AOI211_X1 U20577 ( .C1(n17344), .C2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A(
        n17279), .B(n17278), .ZN(n17280) );
  OAI211_X1 U20578 ( .C1(n17283), .C2(n17282), .A(n17281), .B(n17280), .ZN(
        n17284) );
  AOI211_X1 U20579 ( .C1(n17379), .C2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A(
        n17285), .B(n17284), .ZN(n17519) );
  OAI21_X1 U20580 ( .B1(P3_EBX_REG_15__SCAN_IN), .B2(n9954), .A(n17286), .ZN(
        n17287) );
  OAI21_X1 U20581 ( .B1(n17519), .B2(n17418), .A(n17287), .ZN(P3_U2688) );
  AOI22_X1 U20582 ( .A1(n17344), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17327), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n17298) );
  AOI22_X1 U20583 ( .A1(n12552), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17385), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n17289) );
  AOI22_X1 U20584 ( .A1(n17365), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17343), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n17288) );
  OAI211_X1 U20585 ( .C1(n12551), .C2(n17290), .A(n17289), .B(n17288), .ZN(
        n17296) );
  AOI22_X1 U20586 ( .A1(n17379), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n9829), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n17294) );
  AOI22_X1 U20587 ( .A1(n17245), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17357), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n17293) );
  AOI22_X1 U20588 ( .A1(n17309), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n13120), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n17292) );
  NAND2_X1 U20589 ( .A1(n13080), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n17291) );
  NAND4_X1 U20590 ( .A1(n17294), .A2(n17293), .A3(n17292), .A4(n17291), .ZN(
        n17295) );
  AOI211_X1 U20591 ( .C1(n17361), .C2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A(
        n17296), .B(n17295), .ZN(n17297) );
  OAI211_X1 U20592 ( .C1(n9827), .C2(n17299), .A(n17298), .B(n17297), .ZN(
        n17521) );
  INV_X1 U20593 ( .A(n17521), .ZN(n17303) );
  OAI211_X1 U20594 ( .C1(n17301), .C2(P3_EBX_REG_14__SCAN_IN), .A(n17418), .B(
        n17300), .ZN(n17302) );
  OAI21_X1 U20595 ( .B1(n17303), .B2(n17418), .A(n17302), .ZN(P3_U2689) );
  AOI22_X1 U20596 ( .A1(n17245), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17357), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n17304) );
  OAI21_X1 U20597 ( .B1(n17306), .B2(n17305), .A(n17304), .ZN(n17319) );
  AOI22_X1 U20598 ( .A1(n9829), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17343), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n17316) );
  OAI22_X1 U20599 ( .A1(n17363), .A2(n17308), .B1(n17384), .B2(n17307), .ZN(
        n17314) );
  AOI22_X1 U20600 ( .A1(n17379), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n13120), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n17312) );
  AOI22_X1 U20601 ( .A1(n17309), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17385), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n17311) );
  AOI22_X1 U20602 ( .A1(n13079), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n17361), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n17310) );
  NAND3_X1 U20603 ( .A1(n17312), .A2(n17311), .A3(n17310), .ZN(n17313) );
  AOI211_X1 U20604 ( .C1(n13080), .C2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A(
        n17314), .B(n17313), .ZN(n17315) );
  OAI211_X1 U20605 ( .C1(n9827), .C2(n17317), .A(n17316), .B(n17315), .ZN(
        n17318) );
  AOI211_X1 U20606 ( .C1(n12552), .C2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A(
        n17319), .B(n17318), .ZN(n17529) );
  AOI22_X1 U20607 ( .A1(n17547), .A2(n9920), .B1(P3_EBX_REG_12__SCAN_IN), .B2(
        n17418), .ZN(n17320) );
  OAI22_X1 U20608 ( .A1(n17529), .A2(n17418), .B1(n17321), .B2(n17320), .ZN(
        P3_U2691) );
  AOI21_X1 U20609 ( .B1(n17322), .B2(n17354), .A(n17426), .ZN(n17323) );
  INV_X1 U20610 ( .A(n17323), .ZN(n17338) );
  AOI22_X1 U20611 ( .A1(n17245), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17343), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n17336) );
  AOI22_X1 U20612 ( .A1(n9829), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17365), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n17335) );
  OAI22_X1 U20613 ( .A1(n9919), .A2(n17324), .B1(n9827), .B2(n21208), .ZN(
        n17333) );
  OAI22_X1 U20614 ( .A1(n17395), .A2(n17325), .B1(n12551), .B2(n17414), .ZN(
        n17326) );
  AOI21_X1 U20615 ( .B1(n17344), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A(
        n17326), .ZN(n17331) );
  AOI22_X1 U20616 ( .A1(n17378), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17385), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n17330) );
  AOI22_X1 U20617 ( .A1(n12552), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n13120), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n17329) );
  AOI22_X1 U20618 ( .A1(n17327), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n17361), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n17328) );
  NAND4_X1 U20619 ( .A1(n17331), .A2(n17330), .A3(n17329), .A4(n17328), .ZN(
        n17332) );
  AOI211_X1 U20620 ( .C1(n17379), .C2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A(
        n17333), .B(n17332), .ZN(n17334) );
  NAND3_X1 U20621 ( .A1(n17336), .A2(n17335), .A3(n17334), .ZN(n17532) );
  INV_X1 U20622 ( .A(n17532), .ZN(n17337) );
  OAI22_X1 U20623 ( .A1(n9920), .A2(n17338), .B1(n17337), .B2(n17418), .ZN(
        P3_U2692) );
  AOI22_X1 U20624 ( .A1(n17378), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17365), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n17352) );
  AOI22_X1 U20625 ( .A1(n17245), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n9829), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n17339) );
  OAI21_X1 U20626 ( .B1(n17340), .B2(n21293), .A(n17339), .ZN(n17350) );
  OAI22_X1 U20627 ( .A1(n17384), .A2(n21306), .B1(n13050), .B2(n17341), .ZN(
        n17342) );
  AOI21_X1 U20628 ( .B1(n13089), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A(
        n17342), .ZN(n17348) );
  AOI22_X1 U20629 ( .A1(n17357), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n13120), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n17347) );
  AOI22_X1 U20630 ( .A1(n12552), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n17343), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n17346) );
  AOI22_X1 U20631 ( .A1(n17344), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n13079), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17345) );
  NAND4_X1 U20632 ( .A1(n17348), .A2(n17347), .A3(n17346), .A4(n17345), .ZN(
        n17349) );
  AOI211_X1 U20633 ( .C1(n17379), .C2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A(
        n17350), .B(n17349), .ZN(n17351) );
  OAI211_X1 U20634 ( .C1(n17395), .C2(n17353), .A(n17352), .B(n17351), .ZN(
        n17535) );
  INV_X1 U20635 ( .A(n17535), .ZN(n17356) );
  OAI21_X1 U20636 ( .B1(P3_EBX_REG_10__SCAN_IN), .B2(n17375), .A(n17354), .ZN(
        n17355) );
  AOI22_X1 U20637 ( .A1(n17426), .A2(n17356), .B1(n17355), .B2(n17418), .ZN(
        P3_U2693) );
  AOI22_X1 U20638 ( .A1(n17357), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_8__1__SCAN_IN), .B2(n9829), .ZN(n17358) );
  OAI21_X1 U20639 ( .B1(n17360), .B2(n17359), .A(n17358), .ZN(n17373) );
  AOI22_X1 U20640 ( .A1(n12552), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_7__1__SCAN_IN), .B2(n13089), .ZN(n17371) );
  INV_X1 U20641 ( .A(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n17364) );
  AOI22_X1 U20642 ( .A1(n13080), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n17361), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n17362) );
  OAI21_X1 U20643 ( .B1(n17364), .B2(n17363), .A(n17362), .ZN(n17369) );
  AOI22_X1 U20644 ( .A1(n17378), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_5__1__SCAN_IN), .B2(n17365), .ZN(n17367) );
  AOI22_X1 U20645 ( .A1(n17245), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n17385), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n17366) );
  OAI211_X1 U20646 ( .C1(n21090), .C2(n12551), .A(n17367), .B(n17366), .ZN(
        n17368) );
  AOI211_X1 U20647 ( .C1(n17327), .C2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A(
        n17369), .B(n17368), .ZN(n17370) );
  OAI211_X1 U20648 ( .C1(n21308), .C2(n9884), .A(n17371), .B(n17370), .ZN(
        n17372) );
  AOI211_X1 U20649 ( .C1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .C2(n13120), .A(
        n17373), .B(n17372), .ZN(n17539) );
  NAND2_X1 U20650 ( .A1(n17418), .A2(n17374), .ZN(n17398) );
  NAND2_X1 U20651 ( .A1(n17547), .A2(n17375), .ZN(n17376) );
  OAI21_X1 U20652 ( .B1(P3_EBX_REG_9__SCAN_IN), .B2(n17398), .A(n17376), .ZN(
        n17377) );
  AOI21_X1 U20653 ( .B1(n17426), .B2(n17539), .A(n17377), .ZN(P3_U2694) );
  AOI22_X1 U20654 ( .A1(n17379), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17378), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n17380) );
  OAI21_X1 U20655 ( .B1(n9884), .B2(n17381), .A(n17380), .ZN(n17397) );
  AOI22_X1 U20656 ( .A1(n17245), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17365), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n17393) );
  AOI22_X1 U20657 ( .A1(n13089), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17361), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n17382) );
  OAI21_X1 U20658 ( .B1(n17384), .B2(n17383), .A(n17382), .ZN(n17391) );
  AOI22_X1 U20659 ( .A1(n13120), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n17385), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n17388) );
  AOI22_X1 U20660 ( .A1(n17386), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n9829), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n17387) );
  OAI211_X1 U20661 ( .C1(n12551), .C2(n17389), .A(n17388), .B(n17387), .ZN(
        n17390) );
  AOI211_X1 U20662 ( .C1(n17344), .C2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A(
        n17391), .B(n17390), .ZN(n17392) );
  OAI211_X1 U20663 ( .C1(n17395), .C2(n17394), .A(n17393), .B(n17392), .ZN(
        n17396) );
  AOI211_X1 U20664 ( .C1(n12552), .C2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A(
        n17397), .B(n17396), .ZN(n17546) );
  NAND3_X1 U20665 ( .A1(n17547), .A2(P3_EBX_REG_5__SCAN_IN), .A3(n17413), .ZN(
        n17406) );
  NOR2_X1 U20666 ( .A1(n21274), .A2(n17406), .ZN(n17400) );
  AOI21_X1 U20667 ( .B1(P3_EBX_REG_7__SCAN_IN), .B2(n17400), .A(
        P3_EBX_REG_8__SCAN_IN), .ZN(n17399) );
  OAI22_X1 U20668 ( .A1(n17546), .A2(n17418), .B1(n17399), .B2(n17398), .ZN(
        P3_U2695) );
  AOI21_X1 U20669 ( .B1(P3_EBX_REG_7__SCAN_IN), .B2(n17418), .A(n17400), .ZN(
        n17402) );
  OAI22_X1 U20670 ( .A1(n17403), .A2(n17402), .B1(n17401), .B2(n17418), .ZN(
        P3_U2696) );
  NAND2_X1 U20671 ( .A1(n17418), .A2(n17404), .ZN(n17408) );
  NAND2_X1 U20672 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n17426), .ZN(
        n17405) );
  OAI221_X1 U20673 ( .B1(P3_EBX_REG_6__SCAN_IN), .B2(n17406), .C1(n21274), 
        .C2(n17408), .A(n17405), .ZN(P3_U2697) );
  NOR2_X1 U20674 ( .A1(P3_EBX_REG_5__SCAN_IN), .A2(n17413), .ZN(n17409) );
  OAI22_X1 U20675 ( .A1(n17409), .A2(n17408), .B1(n17407), .B2(n17418), .ZN(
        P3_U2698) );
  NOR3_X1 U20676 ( .A1(n18413), .A2(n17425), .A3(n17410), .ZN(n17421) );
  AND2_X1 U20677 ( .A1(P3_EBX_REG_3__SCAN_IN), .A2(n17421), .ZN(n17416) );
  AOI21_X1 U20678 ( .B1(P3_EBX_REG_4__SCAN_IN), .B2(n17418), .A(n17416), .ZN(
        n17412) );
  OAI22_X1 U20679 ( .A1(n17413), .A2(n17412), .B1(n17411), .B2(n17418), .ZN(
        P3_U2699) );
  AOI21_X1 U20680 ( .B1(P3_EBX_REG_3__SCAN_IN), .B2(n17418), .A(n17421), .ZN(
        n17415) );
  OAI22_X1 U20681 ( .A1(n17416), .A2(n17415), .B1(n17414), .B2(n17418), .ZN(
        P3_U2700) );
  AOI21_X1 U20682 ( .B1(n17547), .B2(n17417), .A(n17425), .ZN(n17419) );
  OAI22_X1 U20683 ( .A1(P3_EBX_REG_2__SCAN_IN), .A2(n17419), .B1(
        P3_INSTQUEUE_REG_0__2__SCAN_IN), .B2(n17418), .ZN(n17420) );
  NOR2_X1 U20684 ( .A1(n17421), .A2(n17420), .ZN(P3_U2701) );
  INV_X1 U20685 ( .A(n17425), .ZN(n17422) );
  NAND2_X1 U20686 ( .A1(n17547), .A2(n17422), .ZN(n17428) );
  OAI222_X1 U20687 ( .A1(n17428), .A2(n17424), .B1(n17423), .B2(n17422), .C1(
        n21090), .C2(n17418), .ZN(P3_U2702) );
  AOI22_X1 U20688 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n17426), .B1(
        P3_EBX_REG_0__SCAN_IN), .B2(n17425), .ZN(n17427) );
  OAI21_X1 U20689 ( .B1(P3_EBX_REG_0__SCAN_IN), .B2(n17428), .A(n17427), .ZN(
        P3_U2703) );
  INV_X1 U20690 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n17587) );
  INV_X1 U20691 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n21227) );
  NOR2_X2 U20692 ( .A1(n17659), .A2(n17576), .ZN(n17574) );
  INV_X1 U20693 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n17666) );
  NAND4_X1 U20694 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(P3_EAX_REG_2__SCAN_IN), 
        .A3(P3_EAX_REG_6__SCAN_IN), .A4(P3_EAX_REG_5__SCAN_IN), .ZN(n17429) );
  NOR3_X1 U20695 ( .A1(n21127), .A2(n17666), .A3(n17429), .ZN(n17520) );
  NAND4_X1 U20696 ( .A1(P3_EAX_REG_14__SCAN_IN), .A2(P3_EAX_REG_11__SCAN_IN), 
        .A3(P3_EAX_REG_10__SCAN_IN), .A4(P3_EAX_REG_9__SCAN_IN), .ZN(n17430)
         );
  NAND2_X1 U20697 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(P3_EAX_REG_20__SCAN_IN), 
        .ZN(n17475) );
  NAND4_X1 U20698 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(P3_EAX_REG_19__SCAN_IN), 
        .A3(P3_EAX_REG_18__SCAN_IN), .A4(P3_EAX_REG_17__SCAN_IN), .ZN(n17431)
         );
  NAND2_X1 U20699 ( .A1(P3_EAX_REG_23__SCAN_IN), .A2(n17469), .ZN(n17468) );
  NAND2_X1 U20700 ( .A1(n17440), .A2(P3_EAX_REG_30__SCAN_IN), .ZN(n17436) );
  OAI22_X1 U20701 ( .A1(P3_EAX_REG_30__SCAN_IN), .A2(n17473), .B1(n17575), 
        .B2(n17440), .ZN(n17434) );
  AOI22_X1 U20702 ( .A1(BUF2_REG_31__SCAN_IN), .A2(n17508), .B1(
        P3_EAX_REG_31__SCAN_IN), .B2(n17434), .ZN(n17435) );
  OAI21_X1 U20703 ( .B1(P3_EAX_REG_31__SCAN_IN), .B2(n17436), .A(n17435), .ZN(
        P3_U2704) );
  AOI22_X1 U20704 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17500), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n17508), .ZN(n17438) );
  OAI211_X1 U20705 ( .C1(n17440), .C2(P3_EAX_REG_30__SCAN_IN), .A(n17571), .B(
        n17436), .ZN(n17437) );
  OAI211_X1 U20706 ( .C1(n17439), .C2(n17580), .A(n17438), .B(n17437), .ZN(
        P3_U2705) );
  AOI22_X1 U20707 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17500), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n17508), .ZN(n17443) );
  AOI211_X1 U20708 ( .C1(n17587), .C2(n17446), .A(n17440), .B(n17575), .ZN(
        n17441) );
  INV_X1 U20709 ( .A(n17441), .ZN(n17442) );
  OAI211_X1 U20710 ( .C1(n17580), .C2(n17444), .A(n17443), .B(n17442), .ZN(
        P3_U2706) );
  INV_X1 U20711 ( .A(n17508), .ZN(n17495) );
  AOI22_X1 U20712 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17500), .B1(n17445), .B2(
        n17569), .ZN(n17449) );
  OAI211_X1 U20713 ( .C1(n17447), .C2(P3_EAX_REG_28__SCAN_IN), .A(n17571), .B(
        n17446), .ZN(n17448) );
  OAI211_X1 U20714 ( .C1(n17495), .C2(n19397), .A(n17449), .B(n17448), .ZN(
        P3_U2707) );
  AOI22_X1 U20715 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17500), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n17508), .ZN(n17452) );
  OAI211_X1 U20716 ( .C1(n17454), .C2(P3_EAX_REG_27__SCAN_IN), .A(n17571), .B(
        n17450), .ZN(n17451) );
  OAI211_X1 U20717 ( .C1(n17580), .C2(n17453), .A(n17452), .B(n17451), .ZN(
        P3_U2708) );
  AOI22_X1 U20718 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17500), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n17508), .ZN(n17457) );
  AOI211_X1 U20719 ( .C1(n21227), .C2(n9885), .A(n17454), .B(n17575), .ZN(
        n17455) );
  INV_X1 U20720 ( .A(n17455), .ZN(n17456) );
  OAI211_X1 U20721 ( .C1(n17580), .C2(n17458), .A(n17457), .B(n17456), .ZN(
        P3_U2709) );
  AOI22_X1 U20722 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17500), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n17508), .ZN(n17461) );
  OAI211_X1 U20723 ( .C1(n17459), .C2(P3_EAX_REG_25__SCAN_IN), .A(n17571), .B(
        n9885), .ZN(n17460) );
  OAI211_X1 U20724 ( .C1(n17580), .C2(n17462), .A(n17461), .B(n17460), .ZN(
        P3_U2710) );
  AOI22_X1 U20725 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17500), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n17508), .ZN(n17466) );
  OAI211_X1 U20726 ( .C1(n17464), .C2(P3_EAX_REG_24__SCAN_IN), .A(n17571), .B(
        n17463), .ZN(n17465) );
  OAI211_X1 U20727 ( .C1(n17467), .C2(n17580), .A(n17466), .B(n17465), .ZN(
        P3_U2711) );
  AOI22_X1 U20728 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17500), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n17508), .ZN(n17471) );
  OAI211_X1 U20729 ( .C1(P3_EAX_REG_23__SCAN_IN), .C2(n17469), .A(n17571), .B(
        n17468), .ZN(n17470) );
  OAI211_X1 U20730 ( .C1(n17472), .C2(n17580), .A(n17471), .B(n17470), .ZN(
        P3_U2712) );
  INV_X1 U20731 ( .A(n17500), .ZN(n17513) );
  INV_X1 U20732 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n17640) );
  INV_X1 U20733 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n17636) );
  NAND2_X1 U20734 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n17501), .ZN(n17496) );
  NAND2_X1 U20735 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n17491), .ZN(n17486) );
  NAND2_X1 U20736 ( .A1(n17571), .A2(n17486), .ZN(n17482) );
  OAI21_X1 U20737 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n17473), .A(n17482), .ZN(
        n17479) );
  INV_X1 U20738 ( .A(n17491), .ZN(n17474) );
  NOR3_X1 U20739 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(n17475), .A3(n17474), .ZN(
        n17478) );
  OAI22_X1 U20740 ( .A1(n17476), .A2(n17580), .B1(n19413), .B2(n17495), .ZN(
        n17477) );
  AOI211_X1 U20741 ( .C1(P3_EAX_REG_22__SCAN_IN), .C2(n17479), .A(n17478), .B(
        n17477), .ZN(n17480) );
  OAI21_X1 U20742 ( .B1(n18410), .B2(n17513), .A(n17480), .ZN(P3_U2713) );
  AOI22_X1 U20743 ( .A1(BUF2_REG_21__SCAN_IN), .A2(n17508), .B1(n17569), .B2(
        n17481), .ZN(n17485) );
  INV_X1 U20744 ( .A(n17482), .ZN(n17483) );
  AOI22_X1 U20745 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17500), .B1(
        P3_EAX_REG_21__SCAN_IN), .B2(n17483), .ZN(n17484) );
  OAI211_X1 U20746 ( .C1(P3_EAX_REG_21__SCAN_IN), .C2(n17486), .A(n17485), .B(
        n17484), .ZN(P3_U2714) );
  AOI22_X1 U20747 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17500), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n17508), .ZN(n17488) );
  OAI211_X1 U20748 ( .C1(n17491), .C2(P3_EAX_REG_20__SCAN_IN), .A(n17571), .B(
        n17486), .ZN(n17487) );
  OAI211_X1 U20749 ( .C1(n17489), .C2(n17580), .A(n17488), .B(n17487), .ZN(
        P3_U2715) );
  AOI22_X1 U20750 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17500), .B1(n17569), .B2(
        n17490), .ZN(n17494) );
  AOI211_X1 U20751 ( .C1(n17640), .C2(n17496), .A(n17491), .B(n17575), .ZN(
        n17492) );
  INV_X1 U20752 ( .A(n17492), .ZN(n17493) );
  OAI211_X1 U20753 ( .C1(n17495), .C2(n19392), .A(n17494), .B(n17493), .ZN(
        P3_U2716) );
  AOI22_X1 U20754 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17500), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n17508), .ZN(n17498) );
  OAI211_X1 U20755 ( .C1(n17501), .C2(P3_EAX_REG_18__SCAN_IN), .A(n17571), .B(
        n17496), .ZN(n17497) );
  OAI211_X1 U20756 ( .C1(n17499), .C2(n17580), .A(n17498), .B(n17497), .ZN(
        P3_U2717) );
  AOI22_X1 U20757 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17500), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n17508), .ZN(n17505) );
  INV_X1 U20758 ( .A(n17509), .ZN(n17503) );
  INV_X1 U20759 ( .A(n17501), .ZN(n17502) );
  OAI211_X1 U20760 ( .C1(n17503), .C2(P3_EAX_REG_17__SCAN_IN), .A(n17571), .B(
        n17502), .ZN(n17504) );
  OAI211_X1 U20761 ( .C1(n17506), .C2(n17580), .A(n17505), .B(n17504), .ZN(
        P3_U2718) );
  AOI22_X1 U20762 ( .A1(BUF2_REG_16__SCAN_IN), .A2(n17508), .B1(n17569), .B2(
        n17507), .ZN(n17512) );
  OAI211_X1 U20763 ( .C1(P3_EAX_REG_16__SCAN_IN), .C2(n17510), .A(n17571), .B(
        n17509), .ZN(n17511) );
  OAI211_X1 U20764 ( .C1(n17513), .C2(n18380), .A(n17512), .B(n17511), .ZN(
        P3_U2719) );
  NOR2_X1 U20765 ( .A1(n18413), .A2(n17514), .ZN(n17516) );
  NAND2_X1 U20766 ( .A1(n17571), .A2(n17514), .ZN(n17523) );
  INV_X1 U20767 ( .A(n17523), .ZN(n17515) );
  MUX2_X1 U20768 ( .A(n17516), .B(n17515), .S(P3_EAX_REG_15__SCAN_IN), .Z(
        n17517) );
  AOI21_X1 U20769 ( .B1(BUF2_REG_15__SCAN_IN), .B2(n17578), .A(n17517), .ZN(
        n17518) );
  OAI21_X1 U20770 ( .B1(n17519), .B2(n17580), .A(n17518), .ZN(P3_U2720) );
  INV_X1 U20771 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n17674) );
  INV_X1 U20772 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n17616) );
  NAND3_X1 U20773 ( .A1(n17547), .A2(n17574), .A3(n17520), .ZN(n17549) );
  NAND2_X1 U20774 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(n17542), .ZN(n17537) );
  NAND2_X1 U20775 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n17541), .ZN(n17534) );
  NOR2_X1 U20776 ( .A1(n17674), .A2(n17534), .ZN(n17528) );
  NAND2_X1 U20777 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(n17531), .ZN(n17524) );
  INV_X1 U20778 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n17683) );
  AOI22_X1 U20779 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17578), .B1(n17569), .B2(
        n17521), .ZN(n17522) );
  OAI221_X1 U20780 ( .B1(P3_EAX_REG_14__SCAN_IN), .B2(n17524), .C1(n17683), 
        .C2(n17523), .A(n17522), .ZN(P3_U2721) );
  INV_X1 U20781 ( .A(n17524), .ZN(n17527) );
  AOI21_X1 U20782 ( .B1(P3_EAX_REG_13__SCAN_IN), .B2(n17571), .A(n17531), .ZN(
        n17526) );
  OAI222_X1 U20783 ( .A1(n17567), .A2(n17681), .B1(n17527), .B2(n17526), .C1(
        n17580), .C2(n17525), .ZN(P3_U2722) );
  AOI21_X1 U20784 ( .B1(P3_EAX_REG_12__SCAN_IN), .B2(n17571), .A(n17528), .ZN(
        n17530) );
  OAI222_X1 U20785 ( .A1(n17567), .A2(n17676), .B1(n17531), .B2(n17530), .C1(
        n17580), .C2(n17529), .ZN(P3_U2723) );
  NAND2_X1 U20786 ( .A1(n17571), .A2(n17534), .ZN(n17538) );
  AOI22_X1 U20787 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17578), .B1(n17569), .B2(
        n17532), .ZN(n17533) );
  OAI221_X1 U20788 ( .B1(P3_EAX_REG_11__SCAN_IN), .B2(n17534), .C1(n17674), 
        .C2(n17538), .A(n17533), .ZN(P3_U2724) );
  INV_X1 U20789 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n17612) );
  AOI22_X1 U20790 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17578), .B1(n17569), .B2(
        n17535), .ZN(n17536) );
  OAI221_X1 U20791 ( .B1(n17538), .B2(n17612), .C1(n17538), .C2(n17537), .A(
        n17536), .ZN(P3_U2725) );
  AOI21_X1 U20792 ( .B1(P3_EAX_REG_9__SCAN_IN), .B2(n17571), .A(n17542), .ZN(
        n17540) );
  OAI222_X1 U20793 ( .A1(n17567), .A2(n17670), .B1(n17541), .B2(n17540), .C1(
        n17580), .C2(n17539), .ZN(P3_U2726) );
  AOI211_X1 U20794 ( .C1(n17543), .C2(n17616), .A(n17575), .B(n17542), .ZN(
        n17544) );
  AOI21_X1 U20795 ( .B1(n17578), .B2(BUF2_REG_8__SCAN_IN), .A(n17544), .ZN(
        n17545) );
  OAI21_X1 U20796 ( .B1(n17546), .B2(n17580), .A(n17545), .ZN(P3_U2727) );
  INV_X1 U20797 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n17624) );
  NAND3_X1 U20798 ( .A1(n17547), .A2(n17574), .A3(P3_EAX_REG_2__SCAN_IN), .ZN(
        n17570) );
  NOR2_X1 U20799 ( .A1(n17624), .A2(n17570), .ZN(n17566) );
  NAND2_X1 U20800 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n17562), .ZN(n17552) );
  INV_X1 U20801 ( .A(n17552), .ZN(n17559) );
  NAND2_X1 U20802 ( .A1(P3_EAX_REG_6__SCAN_IN), .A2(n17559), .ZN(n17555) );
  OAI21_X1 U20803 ( .B1(n17575), .B2(n17666), .A(n17555), .ZN(n17548) );
  AOI22_X1 U20804 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17578), .B1(n17549), .B2(
        n17548), .ZN(n17550) );
  OAI21_X1 U20805 ( .B1(n17551), .B2(n17580), .A(n17550), .ZN(P3_U2728) );
  INV_X1 U20806 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n17619) );
  OAI21_X1 U20807 ( .B1(n17619), .B2(n17575), .A(n17552), .ZN(n17554) );
  AOI222_X1 U20808 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17578), .B1(n17555), .B2(
        n17554), .C1(n17569), .C2(n17553), .ZN(n17556) );
  INV_X1 U20809 ( .A(n17556), .ZN(P3_U2729) );
  AOI21_X1 U20810 ( .B1(P3_EAX_REG_5__SCAN_IN), .B2(n17571), .A(n17562), .ZN(
        n17558) );
  OAI222_X1 U20811 ( .A1(n18406), .A2(n17567), .B1(n17559), .B2(n17558), .C1(
        n17580), .C2(n17557), .ZN(P3_U2730) );
  AOI21_X1 U20812 ( .B1(P3_EAX_REG_4__SCAN_IN), .B2(n17571), .A(n17566), .ZN(
        n17561) );
  OAI222_X1 U20813 ( .A1(n18402), .A2(n17567), .B1(n17562), .B2(n17561), .C1(
        n17580), .C2(n17560), .ZN(P3_U2731) );
  INV_X1 U20814 ( .A(n17570), .ZN(n17563) );
  AOI21_X1 U20815 ( .B1(P3_EAX_REG_3__SCAN_IN), .B2(n17571), .A(n17563), .ZN(
        n17565) );
  OAI222_X1 U20816 ( .A1(n18398), .A2(n17567), .B1(n17566), .B2(n17565), .C1(
        n17580), .C2(n17564), .ZN(P3_U2732) );
  AOI22_X1 U20817 ( .A1(n17578), .A2(BUF2_REG_2__SCAN_IN), .B1(n17569), .B2(
        n17568), .ZN(n17573) );
  OAI211_X1 U20818 ( .C1(n17574), .C2(P3_EAX_REG_2__SCAN_IN), .A(n17571), .B(
        n17570), .ZN(n17572) );
  NAND2_X1 U20819 ( .A1(n17573), .A2(n17572), .ZN(P3_U2733) );
  AOI211_X1 U20820 ( .C1(n17659), .C2(n17576), .A(n17575), .B(n17574), .ZN(
        n17577) );
  AOI21_X1 U20821 ( .B1(n17578), .B2(BUF2_REG_1__SCAN_IN), .A(n17577), .ZN(
        n17579) );
  OAI21_X1 U20822 ( .B1(n17581), .B2(n17580), .A(n17579), .ZN(P3_U2734) );
  INV_X2 U20823 ( .A(n19021), .ZN(n18866) );
  NOR2_X4 U20824 ( .A1(n18866), .A2(n17584), .ZN(n17602) );
  NOR2_X1 U20825 ( .A1(n17609), .A2(n17583), .ZN(P3_U2736) );
  INV_X1 U20826 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n17656) );
  AOI22_X1 U20827 ( .A1(n18866), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(n17602), 
        .B2(P3_DATAO_REG_30__SCAN_IN), .ZN(n17585) );
  OAI21_X1 U20828 ( .B1(n17656), .B2(n17604), .A(n17585), .ZN(P3_U2737) );
  AOI22_X1 U20829 ( .A1(n18866), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n17602), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n17586) );
  OAI21_X1 U20830 ( .B1(n17587), .B2(n17604), .A(n17586), .ZN(P3_U2738) );
  INV_X1 U20831 ( .A(P3_UWORD_REG_12__SCAN_IN), .ZN(n21160) );
  INV_X1 U20832 ( .A(n17604), .ZN(n17595) );
  AOI22_X1 U20833 ( .A1(P3_EAX_REG_28__SCAN_IN), .A2(n17595), .B1(n17602), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n17588) );
  OAI21_X1 U20834 ( .B1(n19021), .B2(n21160), .A(n17588), .ZN(P3_U2739) );
  INV_X1 U20835 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n17652) );
  AOI22_X1 U20836 ( .A1(n18866), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n17602), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n17589) );
  OAI21_X1 U20837 ( .B1(n17652), .B2(n17604), .A(n17589), .ZN(P3_U2740) );
  AOI22_X1 U20838 ( .A1(n18866), .A2(P3_UWORD_REG_10__SCAN_IN), .B1(
        P3_DATAO_REG_26__SCAN_IN), .B2(n17602), .ZN(n17590) );
  OAI21_X1 U20839 ( .B1(n21227), .B2(n17604), .A(n17590), .ZN(P3_U2741) );
  INV_X1 U20840 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n17592) );
  AOI22_X1 U20841 ( .A1(n18866), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n17602), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n17591) );
  OAI21_X1 U20842 ( .B1(n17592), .B2(n17604), .A(n17591), .ZN(P3_U2742) );
  AOI22_X1 U20843 ( .A1(n18866), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n17602), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n17593) );
  OAI21_X1 U20844 ( .B1(n10007), .B2(n17604), .A(n17593), .ZN(P3_U2743) );
  INV_X1 U20845 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n17647) );
  AOI22_X1 U20846 ( .A1(n18866), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n17602), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n17594) );
  OAI21_X1 U20847 ( .B1(n17647), .B2(n17604), .A(n17594), .ZN(P3_U2744) );
  INV_X1 U20848 ( .A(P3_DATAO_REG_22__SCAN_IN), .ZN(n21336) );
  AOI22_X1 U20849 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(n17595), .B1(n18866), 
        .B2(P3_UWORD_REG_6__SCAN_IN), .ZN(n17596) );
  OAI21_X1 U20850 ( .B1(n21336), .B2(n17609), .A(n17596), .ZN(P3_U2745) );
  INV_X1 U20851 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n17644) );
  AOI22_X1 U20852 ( .A1(n18866), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n17602), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n17597) );
  OAI21_X1 U20853 ( .B1(n17644), .B2(n17604), .A(n17597), .ZN(P3_U2746) );
  INV_X1 U20854 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n17642) );
  AOI22_X1 U20855 ( .A1(n18866), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n17602), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n17598) );
  OAI21_X1 U20856 ( .B1(n17642), .B2(n17604), .A(n17598), .ZN(P3_U2747) );
  AOI22_X1 U20857 ( .A1(n18866), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n17602), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n17599) );
  OAI21_X1 U20858 ( .B1(n17640), .B2(n17604), .A(n17599), .ZN(P3_U2748) );
  INV_X1 U20859 ( .A(P3_EAX_REG_18__SCAN_IN), .ZN(n17638) );
  AOI22_X1 U20860 ( .A1(n18866), .A2(P3_UWORD_REG_2__SCAN_IN), .B1(n17602), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n17600) );
  OAI21_X1 U20861 ( .B1(n17638), .B2(n17604), .A(n17600), .ZN(P3_U2749) );
  AOI22_X1 U20862 ( .A1(n18866), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n17602), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n17601) );
  OAI21_X1 U20863 ( .B1(n17636), .B2(n17604), .A(n17601), .ZN(P3_U2750) );
  INV_X1 U20864 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n17634) );
  AOI22_X1 U20865 ( .A1(n18866), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n17602), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n17603) );
  OAI21_X1 U20866 ( .B1(n17634), .B2(n17604), .A(n17603), .ZN(P3_U2751) );
  AOI22_X1 U20867 ( .A1(n18866), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n17602), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n17605) );
  OAI21_X1 U20868 ( .B1(n17688), .B2(n17629), .A(n17605), .ZN(P3_U2752) );
  INV_X1 U20869 ( .A(P3_DATAO_REG_14__SCAN_IN), .ZN(n21196) );
  INV_X1 U20870 ( .A(P3_LWORD_REG_14__SCAN_IN), .ZN(n17606) );
  OAI222_X1 U20871 ( .A1(n17609), .A2(n21196), .B1(n17629), .B2(n17683), .C1(
        n19021), .C2(n17606), .ZN(P3_U2753) );
  INV_X1 U20872 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n21210) );
  AOI22_X1 U20873 ( .A1(n18866), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n17602), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n17607) );
  OAI21_X1 U20874 ( .B1(n21210), .B2(n17629), .A(n17607), .ZN(P3_U2754) );
  INV_X1 U20875 ( .A(P3_DATAO_REG_12__SCAN_IN), .ZN(n21242) );
  INV_X1 U20876 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n21292) );
  INV_X1 U20877 ( .A(P3_LWORD_REG_12__SCAN_IN), .ZN(n17608) );
  OAI222_X1 U20878 ( .A1(n17609), .A2(n21242), .B1(n17629), .B2(n21292), .C1(
        n19021), .C2(n17608), .ZN(P3_U2755) );
  AOI22_X1 U20879 ( .A1(n18866), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n17602), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n17610) );
  OAI21_X1 U20880 ( .B1(n17674), .B2(n17629), .A(n17610), .ZN(P3_U2756) );
  AOI22_X1 U20881 ( .A1(n18866), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n17602), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n17611) );
  OAI21_X1 U20882 ( .B1(n17612), .B2(n17629), .A(n17611), .ZN(P3_U2757) );
  INV_X1 U20883 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n17614) );
  AOI22_X1 U20884 ( .A1(n18866), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n17602), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n17613) );
  OAI21_X1 U20885 ( .B1(n17614), .B2(n17629), .A(n17613), .ZN(P3_U2758) );
  AOI22_X1 U20886 ( .A1(n18866), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n17602), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n17615) );
  OAI21_X1 U20887 ( .B1(n17616), .B2(n17629), .A(n17615), .ZN(P3_U2759) );
  AOI22_X1 U20888 ( .A1(n18866), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n17602), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n17617) );
  OAI21_X1 U20889 ( .B1(n17666), .B2(n17629), .A(n17617), .ZN(P3_U2760) );
  AOI22_X1 U20890 ( .A1(n18866), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n17602), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n17618) );
  OAI21_X1 U20891 ( .B1(n17619), .B2(n17629), .A(n17618), .ZN(P3_U2761) );
  INV_X1 U20892 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n17621) );
  AOI22_X1 U20893 ( .A1(n18866), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n17602), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n17620) );
  OAI21_X1 U20894 ( .B1(n17621), .B2(n17629), .A(n17620), .ZN(P3_U2762) );
  AOI22_X1 U20895 ( .A1(n18866), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n17602), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n17622) );
  OAI21_X1 U20896 ( .B1(n21127), .B2(n17629), .A(n17622), .ZN(P3_U2763) );
  AOI22_X1 U20897 ( .A1(n18866), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n17602), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n17623) );
  OAI21_X1 U20898 ( .B1(n17624), .B2(n17629), .A(n17623), .ZN(P3_U2764) );
  INV_X1 U20899 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n17626) );
  AOI22_X1 U20900 ( .A1(n18866), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n17602), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n17625) );
  OAI21_X1 U20901 ( .B1(n17626), .B2(n17629), .A(n17625), .ZN(P3_U2765) );
  AOI22_X1 U20902 ( .A1(n18866), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n17602), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n17627) );
  OAI21_X1 U20903 ( .B1(n17659), .B2(n17629), .A(n17627), .ZN(P3_U2766) );
  AOI22_X1 U20904 ( .A1(n18866), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n17602), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n17628) );
  OAI21_X1 U20905 ( .B1(n17630), .B2(n17629), .A(n17628), .ZN(P3_U2767) );
  AOI22_X1 U20906 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17685), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n17684), .ZN(n17633) );
  OAI21_X1 U20907 ( .B1(n17634), .B2(n17687), .A(n17633), .ZN(P3_U2768) );
  AOI22_X1 U20908 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17685), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n17684), .ZN(n17635) );
  OAI21_X1 U20909 ( .B1(n17636), .B2(n17687), .A(n17635), .ZN(P3_U2769) );
  AOI22_X1 U20910 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17685), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n17684), .ZN(n17637) );
  OAI21_X1 U20911 ( .B1(n17638), .B2(n17687), .A(n17637), .ZN(P3_U2770) );
  AOI22_X1 U20912 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17685), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n17684), .ZN(n17639) );
  OAI21_X1 U20913 ( .B1(n17640), .B2(n17687), .A(n17639), .ZN(P3_U2771) );
  AOI22_X1 U20914 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17685), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n17684), .ZN(n17641) );
  OAI21_X1 U20915 ( .B1(n17642), .B2(n17687), .A(n17641), .ZN(P3_U2772) );
  AOI22_X1 U20916 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17685), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n17684), .ZN(n17643) );
  OAI21_X1 U20917 ( .B1(n17644), .B2(n17687), .A(n17643), .ZN(P3_U2773) );
  AOI22_X1 U20918 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(n17678), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n17684), .ZN(n17645) );
  OAI21_X1 U20919 ( .B1(n18410), .B2(n17680), .A(n17645), .ZN(P3_U2774) );
  AOI22_X1 U20920 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17685), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n17684), .ZN(n17646) );
  OAI21_X1 U20921 ( .B1(n17647), .B2(n17687), .A(n17646), .ZN(P3_U2775) );
  AOI22_X1 U20922 ( .A1(P3_EAX_REG_24__SCAN_IN), .A2(n17678), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n17684), .ZN(n17648) );
  OAI21_X1 U20923 ( .B1(n17668), .B2(n17680), .A(n17648), .ZN(P3_U2776) );
  AOI22_X1 U20924 ( .A1(P3_EAX_REG_25__SCAN_IN), .A2(n17678), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n17684), .ZN(n17649) );
  OAI21_X1 U20925 ( .B1(n17670), .B2(n17680), .A(n17649), .ZN(P3_U2777) );
  AOI22_X1 U20926 ( .A1(P3_EAX_REG_26__SCAN_IN), .A2(n17678), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n17684), .ZN(n17650) );
  OAI21_X1 U20927 ( .B1(n17672), .B2(n17680), .A(n17650), .ZN(P3_U2778) );
  AOI22_X1 U20928 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17685), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n17684), .ZN(n17651) );
  OAI21_X1 U20929 ( .B1(n17652), .B2(n17687), .A(n17651), .ZN(P3_U2779) );
  AOI22_X1 U20930 ( .A1(P3_EAX_REG_28__SCAN_IN), .A2(n17678), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n17684), .ZN(n17653) );
  OAI21_X1 U20931 ( .B1(n17676), .B2(n17680), .A(n17653), .ZN(P3_U2780) );
  AOI22_X1 U20932 ( .A1(P3_EAX_REG_29__SCAN_IN), .A2(n17678), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n17684), .ZN(n17654) );
  OAI21_X1 U20933 ( .B1(n17681), .B2(n17680), .A(n17654), .ZN(P3_U2781) );
  AOI22_X1 U20934 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17685), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n17684), .ZN(n17655) );
  OAI21_X1 U20935 ( .B1(n17656), .B2(n17687), .A(n17655), .ZN(P3_U2782) );
  AOI22_X1 U20936 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(n17678), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n17684), .ZN(n17657) );
  OAI21_X1 U20937 ( .B1(n18380), .B2(n17680), .A(n17657), .ZN(P3_U2783) );
  AOI22_X1 U20938 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17685), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n17684), .ZN(n17658) );
  OAI21_X1 U20939 ( .B1(n17659), .B2(n17687), .A(n17658), .ZN(P3_U2784) );
  AOI22_X1 U20940 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(n17678), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n17684), .ZN(n17660) );
  OAI21_X1 U20941 ( .B1(n18394), .B2(n17680), .A(n17660), .ZN(P3_U2785) );
  AOI22_X1 U20942 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n17678), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n17684), .ZN(n17661) );
  OAI21_X1 U20943 ( .B1(n18398), .B2(n17680), .A(n17661), .ZN(P3_U2786) );
  AOI22_X1 U20944 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(n17678), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n17677), .ZN(n17662) );
  OAI21_X1 U20945 ( .B1(n18402), .B2(n17680), .A(n17662), .ZN(P3_U2787) );
  AOI22_X1 U20946 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n17678), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n17677), .ZN(n17663) );
  OAI21_X1 U20947 ( .B1(n18406), .B2(n17680), .A(n17663), .ZN(P3_U2788) );
  AOI22_X1 U20948 ( .A1(P3_EAX_REG_6__SCAN_IN), .A2(n17678), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n17677), .ZN(n17664) );
  OAI21_X1 U20949 ( .B1(n18410), .B2(n17680), .A(n17664), .ZN(P3_U2789) );
  AOI22_X1 U20950 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17685), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n17677), .ZN(n17665) );
  OAI21_X1 U20951 ( .B1(n17666), .B2(n17687), .A(n17665), .ZN(P3_U2790) );
  AOI22_X1 U20952 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n17678), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n17677), .ZN(n17667) );
  OAI21_X1 U20953 ( .B1(n17668), .B2(n17680), .A(n17667), .ZN(P3_U2791) );
  AOI22_X1 U20954 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(n17678), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n17677), .ZN(n17669) );
  OAI21_X1 U20955 ( .B1(n17670), .B2(n17680), .A(n17669), .ZN(P3_U2792) );
  AOI22_X1 U20956 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n17678), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n17677), .ZN(n17671) );
  OAI21_X1 U20957 ( .B1(n17672), .B2(n17680), .A(n17671), .ZN(P3_U2793) );
  AOI22_X1 U20958 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17685), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n17677), .ZN(n17673) );
  OAI21_X1 U20959 ( .B1(n17674), .B2(n17687), .A(n17673), .ZN(P3_U2794) );
  AOI22_X1 U20960 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n17678), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n17677), .ZN(n17675) );
  OAI21_X1 U20961 ( .B1(n17676), .B2(n17680), .A(n17675), .ZN(P3_U2795) );
  AOI22_X1 U20962 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(n17678), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n17677), .ZN(n17679) );
  OAI21_X1 U20963 ( .B1(n17681), .B2(n17680), .A(n17679), .ZN(P3_U2796) );
  AOI22_X1 U20964 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17685), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n17684), .ZN(n17682) );
  OAI21_X1 U20965 ( .B1(n17683), .B2(n17687), .A(n17682), .ZN(P3_U2797) );
  AOI22_X1 U20966 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n17685), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n17684), .ZN(n17686) );
  OAI21_X1 U20967 ( .B1(n17688), .B2(n17687), .A(n17686), .ZN(P3_U2798) );
  INV_X1 U20968 ( .A(n18045), .ZN(n18034) );
  AOI21_X1 U20969 ( .B1(n17702), .B2(n17890), .A(n18034), .ZN(n17689) );
  INV_X1 U20970 ( .A(n17689), .ZN(n17690) );
  AOI21_X1 U20971 ( .B1(n17892), .B2(n17691), .A(n17690), .ZN(n17724) );
  OAI21_X1 U20972 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n17776), .A(
        n17724), .ZN(n17713) );
  AOI22_X1 U20973 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n17713), .B1(
        n17895), .B2(n17692), .ZN(n17707) );
  NOR2_X1 U20974 ( .A1(n18039), .A2(n17926), .ZN(n17810) );
  NOR2_X1 U20975 ( .A1(n17810), .A2(n17693), .ZN(n17701) );
  NAND2_X1 U20976 ( .A1(n17734), .A2(n17694), .ZN(n18059) );
  NAND3_X1 U20977 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(n17741), .ZN(n18058) );
  AOI22_X1 U20978 ( .A1(n18039), .A2(n18059), .B1(n17926), .B2(n18058), .ZN(
        n17732) );
  NAND2_X1 U20979 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n17732), .ZN(
        n17718) );
  AOI211_X1 U20980 ( .C1(n17697), .C2(n17696), .A(n17695), .B(n17889), .ZN(
        n17700) );
  INV_X1 U20981 ( .A(n17772), .ZN(n17717) );
  NOR3_X1 U20982 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17698), .A3(
        n17717), .ZN(n17699) );
  AOI211_X1 U20983 ( .C1(n17701), .C2(n17718), .A(n17700), .B(n17699), .ZN(
        n17706) );
  NAND2_X1 U20984 ( .A1(n18096), .A2(P3_REIP_REG_28__SCAN_IN), .ZN(n17705) );
  NOR2_X1 U20985 ( .A1(n17901), .A2(n17702), .ZN(n17715) );
  OAI211_X1 U20986 ( .C1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A(n17715), .B(n17703), .ZN(n17704) );
  NAND4_X1 U20987 ( .A1(n17707), .A2(n17706), .A3(n17705), .A4(n17704), .ZN(
        P3_U2802) );
  NAND2_X1 U20988 ( .A1(n17709), .A2(n17708), .ZN(n17710) );
  XNOR2_X1 U20989 ( .A(n17957), .B(n17710), .ZN(n18068) );
  OAI22_X1 U20990 ( .A1(n18316), .A2(n18945), .B1(n17919), .B2(n17711), .ZN(
        n17712) );
  AOI221_X1 U20991 ( .B1(n17715), .B2(n17714), .C1(n17713), .C2(
        P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A(n17712), .ZN(n17721) );
  INV_X1 U20992 ( .A(n17716), .ZN(n18053) );
  NOR2_X1 U20993 ( .A1(n18053), .A2(n17717), .ZN(n17719) );
  OAI21_X1 U20994 ( .B1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n17719), .A(
        n17718), .ZN(n17720) );
  OAI211_X1 U20995 ( .C1(n18068), .C2(n17889), .A(n17721), .B(n17720), .ZN(
        P3_U2803) );
  AOI21_X1 U20996 ( .B1(n17722), .B2(n18748), .A(
        P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n17723) );
  OAI22_X1 U20997 ( .A1(n17724), .A2(n17723), .B1(n18316), .B2(n18943), .ZN(
        n17725) );
  AOI221_X1 U20998 ( .B1(n17895), .B2(n17726), .C1(n17806), .C2(n17726), .A(
        n17725), .ZN(n17731) );
  OAI21_X1 U20999 ( .B1(n17728), .B2(n18054), .A(n17727), .ZN(n18070) );
  NOR3_X1 U21000 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n17744), .A3(
        n17729), .ZN(n18069) );
  AOI22_X1 U21001 ( .A1(n17963), .A2(n18070), .B1(n17849), .B2(n18069), .ZN(
        n17730) );
  OAI211_X1 U21002 ( .C1(n17732), .C2(n18054), .A(n17731), .B(n17730), .ZN(
        P3_U2804) );
  INV_X1 U21003 ( .A(n17734), .ZN(n17733) );
  AOI22_X1 U21004 ( .A1(n17734), .A2(n17744), .B1(
        P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n17733), .ZN(n18084) );
  AND2_X1 U21005 ( .A1(n17736), .A2(n18748), .ZN(n17765) );
  AOI211_X1 U21006 ( .C1(n17892), .C2(n17735), .A(n18034), .B(n17765), .ZN(
        n17769) );
  OAI21_X1 U21007 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n17776), .A(
        n17769), .ZN(n17752) );
  NOR2_X1 U21008 ( .A1(n17901), .A2(n17736), .ZN(n17754) );
  OAI211_X1 U21009 ( .C1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A(n17754), .B(n17737), .ZN(n17738) );
  NAND2_X1 U21010 ( .A1(n18096), .A2(P3_REIP_REG_25__SCAN_IN), .ZN(n18081) );
  OAI211_X1 U21011 ( .C1(n17919), .C2(n17739), .A(n17738), .B(n18081), .ZN(
        n17747) );
  NAND2_X1 U21012 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n17741), .ZN(
        n17740) );
  OAI21_X1 U21013 ( .B1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n17741), .A(
        n17740), .ZN(n18088) );
  OAI21_X1 U21014 ( .B1(n17957), .B2(n17743), .A(n17742), .ZN(n17745) );
  XNOR2_X1 U21015 ( .A(n17745), .B(n17744), .ZN(n18083) );
  OAI22_X1 U21016 ( .A1(n17961), .A2(n18088), .B1(n17889), .B2(n18083), .ZN(
        n17746) );
  AOI211_X1 U21017 ( .C1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .C2(n17752), .A(
        n17747), .B(n17746), .ZN(n17748) );
  OAI21_X1 U21018 ( .B1(n18050), .B2(n18084), .A(n17748), .ZN(P3_U2805) );
  NAND2_X1 U21019 ( .A1(n17749), .A2(n18098), .ZN(n18104) );
  OAI22_X1 U21020 ( .A1(n18316), .A2(n18939), .B1(n17919), .B2(n17750), .ZN(
        n17751) );
  AOI221_X1 U21021 ( .B1(n17754), .B2(n17753), .C1(n17752), .C2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A(n17751), .ZN(n17759) );
  NOR2_X1 U21022 ( .A1(n17755), .A2(n18188), .ZN(n18091) );
  NOR2_X1 U21023 ( .A1(n18194), .A2(n17755), .ZN(n18090) );
  OAI22_X1 U21024 ( .A1(n18091), .A2(n17961), .B1(n18090), .B2(n18050), .ZN(
        n17771) );
  OAI21_X1 U21025 ( .B1(n17757), .B2(n18098), .A(n17756), .ZN(n18101) );
  AOI22_X1 U21026 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17771), .B1(
        n17963), .B2(n18101), .ZN(n17758) );
  OAI211_X1 U21027 ( .C1(n17864), .C2(n18104), .A(n17759), .B(n17758), .ZN(
        P3_U2806) );
  OAI22_X1 U21028 ( .A1(n17957), .A2(n18127), .B1(n17760), .B2(n17778), .ZN(
        n17761) );
  NOR2_X1 U21029 ( .A1(n17761), .A2(n17811), .ZN(n17762) );
  XNOR2_X1 U21030 ( .A(n17762), .B(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n18110) );
  AOI22_X1 U21031 ( .A1(n17766), .A2(n17765), .B1(n17764), .B2(n17763), .ZN(
        n17767) );
  NAND2_X1 U21032 ( .A1(n18096), .A2(P3_REIP_REG_23__SCAN_IN), .ZN(n18109) );
  OAI211_X1 U21033 ( .C1(n17769), .C2(n17768), .A(n17767), .B(n18109), .ZN(
        n17770) );
  AOI221_X1 U21034 ( .B1(n17772), .B2(n18094), .C1(n17771), .C2(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A(n17770), .ZN(n17773) );
  OAI21_X1 U21035 ( .B1(n17889), .B2(n18110), .A(n17773), .ZN(P3_U2807) );
  OAI21_X1 U21036 ( .B1(n17774), .B2(n18046), .A(n18045), .ZN(n17775) );
  AOI21_X1 U21037 ( .B1(n17890), .B2(n17785), .A(n17775), .ZN(n17803) );
  OAI21_X1 U21038 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n17776), .A(
        n17803), .ZN(n17792) );
  AOI22_X1 U21039 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n17792), .B1(
        n17895), .B2(n17777), .ZN(n17789) );
  INV_X1 U21040 ( .A(n17778), .ZN(n17780) );
  AOI21_X1 U21041 ( .B1(n17780), .B2(n17779), .A(n17811), .ZN(n17781) );
  XNOR2_X1 U21042 ( .A(n17781), .B(n18127), .ZN(n18123) );
  NOR2_X1 U21043 ( .A1(n18114), .A2(n17864), .ZN(n17783) );
  AOI22_X1 U21044 ( .A1(n18194), .A2(n18039), .B1(n18188), .B2(n17926), .ZN(
        n17863) );
  OAI21_X1 U21045 ( .B1(n18120), .B2(n17810), .A(n17863), .ZN(n17782) );
  INV_X1 U21046 ( .A(n17782), .ZN(n17802) );
  MUX2_X1 U21047 ( .A(n17783), .B(n17782), .S(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .Z(n17784) );
  AOI21_X1 U21048 ( .B1(n17963), .B2(n18123), .A(n17784), .ZN(n17788) );
  NAND2_X1 U21049 ( .A1(n18096), .A2(P3_REIP_REG_22__SCAN_IN), .ZN(n18125) );
  NOR2_X1 U21050 ( .A1(n17901), .A2(n17785), .ZN(n17794) );
  OAI211_X1 U21051 ( .C1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A(n17794), .B(n17786), .ZN(n17787) );
  NAND4_X1 U21052 ( .A1(n17789), .A2(n17788), .A3(n18125), .A4(n17787), .ZN(
        P3_U2808) );
  INV_X1 U21053 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n17793) );
  OAI22_X1 U21054 ( .A1(n18316), .A2(n18933), .B1(n17919), .B2(n17790), .ZN(
        n17791) );
  AOI221_X1 U21055 ( .B1(n17794), .B2(n17793), .C1(n17792), .C2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A(n17791), .ZN(n17800) );
  OR3_X1 U21056 ( .A1(n17828), .A2(n13160), .A3(n17795), .ZN(n17815) );
  OAI22_X1 U21057 ( .A1(n17798), .A2(n17815), .B1(n17829), .B2(n17796), .ZN(
        n17797) );
  XOR2_X1 U21058 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .B(n17797), .Z(
        n18136) );
  NOR4_X1 U21059 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17836), .A3(
        n17828), .A4(n17798), .ZN(n18135) );
  AOI22_X1 U21060 ( .A1(n17963), .A2(n18136), .B1(n17849), .B2(n18135), .ZN(
        n17799) );
  OAI211_X1 U21061 ( .C1(n17802), .C2(n17801), .A(n17800), .B(n17799), .ZN(
        P3_U2809) );
  NAND2_X1 U21062 ( .A1(n18161), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n18128) );
  NOR2_X1 U21063 ( .A1(n18156), .A2(n18128), .ZN(n18141) );
  NAND2_X1 U21064 ( .A1(n18141), .A2(n18115), .ZN(n18149) );
  NAND2_X1 U21065 ( .A1(n9922), .A2(n18748), .ZN(n17840) );
  AOI221_X1 U21066 ( .B1(n17805), .B2(n17804), .C1(n17840), .C2(n17804), .A(
        n17803), .ZN(n17809) );
  AOI21_X1 U21067 ( .B1(n17919), .B2(n17776), .A(n17807), .ZN(n17808) );
  AOI211_X1 U21068 ( .C1(P3_REIP_REG_20__SCAN_IN), .C2(n18096), .A(n17809), 
        .B(n17808), .ZN(n17814) );
  OAI21_X1 U21069 ( .B1(n17810), .B2(n18141), .A(n17863), .ZN(n17823) );
  AOI221_X1 U21070 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n17815), 
        .C1(n18156), .C2(n17827), .A(n17811), .ZN(n17812) );
  XNOR2_X1 U21071 ( .A(n17812), .B(n18115), .ZN(n18144) );
  AOI22_X1 U21072 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n17823), .B1(
        n17963), .B2(n18144), .ZN(n17813) );
  OAI211_X1 U21073 ( .C1(n17864), .C2(n18149), .A(n17814), .B(n17813), .ZN(
        P3_U2810) );
  OAI21_X1 U21074 ( .B1(n17827), .B2(n17829), .A(n17815), .ZN(n17816) );
  XOR2_X1 U21075 ( .A(n17816), .B(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .Z(
        n18152) );
  INV_X1 U21076 ( .A(n18152), .ZN(n17826) );
  AOI21_X1 U21077 ( .B1(n17890), .B2(n17818), .A(n18034), .ZN(n17839) );
  OAI21_X1 U21078 ( .B1(n17817), .B2(n18046), .A(n17839), .ZN(n17833) );
  NOR2_X1 U21079 ( .A1(n17901), .A2(n17818), .ZN(n17835) );
  NAND2_X1 U21080 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n17819) );
  OAI211_X1 U21081 ( .C1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(n17835), .B(n17819), .ZN(n17820) );
  NAND2_X1 U21082 ( .A1(n18096), .A2(P3_REIP_REG_19__SCAN_IN), .ZN(n18153) );
  OAI211_X1 U21083 ( .C1(n17919), .C2(n17821), .A(n17820), .B(n18153), .ZN(
        n17822) );
  AOI21_X1 U21084 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n17833), .A(
        n17822), .ZN(n17825) );
  NOR2_X1 U21085 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18128), .ZN(
        n18150) );
  AOI22_X1 U21086 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17823), .B1(
        n17849), .B2(n18150), .ZN(n17824) );
  OAI211_X1 U21087 ( .C1(n17826), .C2(n17889), .A(n17825), .B(n17824), .ZN(
        P3_U2811) );
  OAI21_X1 U21088 ( .B1(n13160), .B2(n17828), .A(n17827), .ZN(n17830) );
  XNOR2_X1 U21089 ( .A(n17830), .B(n17829), .ZN(n18169) );
  NAND2_X1 U21090 ( .A1(n18096), .A2(P3_REIP_REG_18__SCAN_IN), .ZN(n18167) );
  OAI21_X1 U21091 ( .B1(n17919), .B2(n17831), .A(n18167), .ZN(n17832) );
  AOI221_X1 U21092 ( .B1(n17835), .B2(n17834), .C1(n17833), .C2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(n17832), .ZN(n17838) );
  OAI21_X1 U21093 ( .B1(n18161), .B2(n17864), .A(n17863), .ZN(n17845) );
  NOR2_X1 U21094 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17836), .ZN(
        n18165) );
  AOI22_X1 U21095 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17845), .B1(
        n17849), .B2(n18165), .ZN(n17837) );
  OAI211_X1 U21096 ( .C1(n17889), .C2(n18169), .A(n17838), .B(n17837), .ZN(
        P3_U2812) );
  INV_X1 U21097 ( .A(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n17841) );
  AOI21_X1 U21098 ( .B1(n17841), .B2(n17840), .A(n17839), .ZN(n17844) );
  NAND2_X1 U21099 ( .A1(n18096), .A2(P3_REIP_REG_17__SCAN_IN), .ZN(n18172) );
  OAI21_X1 U21100 ( .B1(n18031), .B2(n17842), .A(n18172), .ZN(n17843) );
  AOI211_X1 U21101 ( .C1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .C2(n17845), .A(
        n17844), .B(n17843), .ZN(n17851) );
  OAI21_X1 U21102 ( .B1(n17848), .B2(n17847), .A(n17846), .ZN(n18171) );
  NOR2_X1 U21103 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n18181), .ZN(
        n18170) );
  AOI22_X1 U21104 ( .A1(n17963), .A2(n18171), .B1(n17849), .B2(n18170), .ZN(
        n17850) );
  NAND2_X1 U21105 ( .A1(n17851), .A2(n17850), .ZN(P3_U2813) );
  NAND2_X1 U21106 ( .A1(n17957), .A2(n17896), .ZN(n17934) );
  INV_X1 U21107 ( .A(n17934), .ZN(n17943) );
  AOI22_X1 U21108 ( .A1(n17943), .A2(n17853), .B1(n17852), .B2(n13160), .ZN(
        n17854) );
  XNOR2_X1 U21109 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B(n17854), .ZN(
        n18183) );
  AOI21_X1 U21110 ( .B1(n17890), .B2(n17856), .A(n18034), .ZN(n17884) );
  OAI21_X1 U21111 ( .B1(n17855), .B2(n18046), .A(n17884), .ZN(n17865) );
  AOI22_X1 U21112 ( .A1(n18096), .A2(P3_REIP_REG_16__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n17865), .ZN(n17859) );
  NOR2_X1 U21113 ( .A1(n17901), .A2(n17856), .ZN(n17867) );
  OAI211_X1 U21114 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(n17867), .B(n17857), .ZN(n17858) );
  OAI211_X1 U21115 ( .C1(n17919), .C2(n17860), .A(n17859), .B(n17858), .ZN(
        n17861) );
  AOI21_X1 U21116 ( .B1(n17963), .B2(n18183), .A(n17861), .ZN(n17862) );
  OAI221_X1 U21117 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n17864), 
        .C1(n18181), .C2(n17863), .A(n17862), .ZN(P3_U2814) );
  NOR2_X1 U21118 ( .A1(n18316), .A2(n18921), .ZN(n18192) );
  AOI221_X1 U21119 ( .B1(n17867), .B2(n17866), .C1(n17865), .C2(
        P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A(n18192), .ZN(n17878) );
  AND2_X1 U21120 ( .A1(n18194), .A2(n18039), .ZN(n17876) );
  OR2_X1 U21121 ( .A1(n18195), .A2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n17875) );
  NOR2_X1 U21122 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n18189), .ZN(
        n17873) );
  NAND2_X1 U21123 ( .A1(n17926), .A2(n18188), .ZN(n17872) );
  AOI21_X1 U21124 ( .B1(n17896), .B2(n17869), .A(n17868), .ZN(n17870) );
  AOI221_X1 U21125 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n18237), 
        .C1(n13160), .C2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A(n17870), .ZN(
        n17871) );
  XNOR2_X1 U21126 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B(n17871), .ZN(
        n18198) );
  OAI22_X1 U21127 ( .A1(n17873), .A2(n17872), .B1(n17889), .B2(n18198), .ZN(
        n17874) );
  AOI21_X1 U21128 ( .B1(n17876), .B2(n17875), .A(n17874), .ZN(n17877) );
  OAI211_X1 U21129 ( .C1(n17919), .C2(n17879), .A(n17878), .B(n17877), .ZN(
        P3_U2815) );
  NAND2_X1 U21130 ( .A1(n18228), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n18200) );
  INV_X1 U21131 ( .A(n18200), .ZN(n17880) );
  AOI22_X1 U21132 ( .A1(n17880), .A2(n17943), .B1(n17868), .B2(n18237), .ZN(
        n17881) );
  XOR2_X1 U21133 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B(n17881), .Z(
        n18212) );
  AOI21_X1 U21134 ( .B1(n17882), .B2(n18748), .A(
        P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n17883) );
  OAI22_X1 U21135 ( .A1(n18031), .A2(n17885), .B1(n17884), .B2(n17883), .ZN(
        n17886) );
  AOI21_X1 U21136 ( .B1(n18096), .B2(P3_REIP_REG_14__SCAN_IN), .A(n17886), 
        .ZN(n17888) );
  INV_X1 U21137 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n18202) );
  AOI221_X1 U21138 ( .B1(n10166), .B2(n18202), .C1(n18221), .C2(n18202), .A(
        n18195), .ZN(n18207) );
  AOI221_X1 U21139 ( .B1(n10166), .B2(n18202), .C1(n18217), .C2(n18202), .A(
        n18189), .ZN(n18208) );
  AOI22_X1 U21140 ( .A1(n18039), .A2(n18207), .B1(n17926), .B2(n18208), .ZN(
        n17887) );
  OAI211_X1 U21141 ( .C1(n18212), .C2(n17889), .A(n17888), .B(n17887), .ZN(
        P3_U2816) );
  AOI22_X1 U21142 ( .A1(n17892), .A2(n17891), .B1(n17890), .B2(n17900), .ZN(
        n17893) );
  NAND2_X1 U21143 ( .A1(n17893), .A2(n18045), .ZN(n17907) );
  AOI22_X1 U21144 ( .A1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n17907), .B1(
        n17895), .B2(n17894), .ZN(n17906) );
  AOI22_X1 U21145 ( .A1(n17896), .A2(n18228), .B1(n18237), .B2(n13160), .ZN(
        n17897) );
  AOI21_X1 U21146 ( .B1(n17910), .B2(n13160), .A(n17897), .ZN(n17898) );
  XNOR2_X1 U21147 ( .A(n17898), .B(n10166), .ZN(n18216) );
  NAND2_X1 U21148 ( .A1(n18228), .A2(n10166), .ZN(n18227) );
  AOI22_X1 U21149 ( .A1(n18039), .A2(n18221), .B1(n17926), .B2(n18217), .ZN(
        n17912) );
  OAI22_X1 U21150 ( .A1(n17953), .A2(n18227), .B1(n17912), .B2(n10166), .ZN(
        n17899) );
  AOI21_X1 U21151 ( .B1(n17963), .B2(n18216), .A(n17899), .ZN(n17905) );
  NAND2_X1 U21152 ( .A1(n18096), .A2(P3_REIP_REG_13__SCAN_IN), .ZN(n17904) );
  NOR2_X1 U21153 ( .A1(n17901), .A2(n17900), .ZN(n17909) );
  OAI211_X1 U21154 ( .C1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A(n17909), .B(n17902), .ZN(n17903) );
  NAND4_X1 U21155 ( .A1(n17906), .A2(n17905), .A3(n17904), .A4(n17903), .ZN(
        P3_U2817) );
  INV_X1 U21156 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n17908) );
  INV_X1 U21157 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n18918) );
  NOR2_X1 U21158 ( .A1(n18316), .A2(n18918), .ZN(n18234) );
  AOI221_X1 U21159 ( .B1(n17909), .B2(n17908), .C1(n17907), .C2(
        P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A(n18234), .ZN(n17917) );
  OAI21_X1 U21160 ( .B1(n18250), .B2(n17934), .A(n17910), .ZN(n17911) );
  XNOR2_X1 U21161 ( .A(n17911), .B(n18237), .ZN(n18233) );
  NOR2_X1 U21162 ( .A1(n17953), .A2(n18250), .ZN(n17914) );
  INV_X1 U21163 ( .A(n17912), .ZN(n17913) );
  MUX2_X1 U21164 ( .A(n17914), .B(n17913), .S(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .Z(n17915) );
  AOI21_X1 U21165 ( .B1(n17963), .B2(n18233), .A(n17915), .ZN(n17916) );
  OAI211_X1 U21166 ( .C1(n17919), .C2(n17918), .A(n17917), .B(n17916), .ZN(
        P3_U2818) );
  NAND2_X1 U21167 ( .A1(n18240), .A2(n17920), .ZN(n18255) );
  NOR2_X1 U21168 ( .A1(n17921), .A2(n18418), .ZN(n17941) );
  NOR2_X1 U21169 ( .A1(n17924), .A2(n17941), .ZN(n17925) );
  OAI22_X1 U21170 ( .A1(n18031), .A2(n17922), .B1(n18316), .B2(n18916), .ZN(
        n17923) );
  AOI221_X1 U21171 ( .B1(n18041), .B2(n17925), .C1(n17924), .C2(n17941), .A(
        n17923), .ZN(n17930) );
  INV_X1 U21172 ( .A(n18215), .ZN(n18243) );
  INV_X1 U21173 ( .A(n18214), .ZN(n18241) );
  AOI22_X1 U21174 ( .A1(n18039), .A2(n18243), .B1(n17926), .B2(n18241), .ZN(
        n17952) );
  OAI21_X1 U21175 ( .B1(n18240), .B2(n17953), .A(n17952), .ZN(n17937) );
  AOI21_X1 U21176 ( .B1(n18240), .B2(n17943), .A(n17927), .ZN(n17928) );
  XNOR2_X1 U21177 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n17928), .ZN(
        n18238) );
  AOI22_X1 U21178 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n17937), .B1(
        n17963), .B2(n18238), .ZN(n17929) );
  OAI211_X1 U21179 ( .C1(n17953), .C2(n18255), .A(n17930), .B(n17929), .ZN(
        P3_U2819) );
  NOR3_X1 U21180 ( .A1(n17945), .A2(n17931), .A3(n18418), .ZN(n17949) );
  AOI21_X1 U21181 ( .B1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n18041), .A(
        n17949), .ZN(n17940) );
  AOI22_X1 U21182 ( .A1(n18096), .A2(P3_REIP_REG_10__SCAN_IN), .B1(n17932), 
        .B2(n17763), .ZN(n17939) );
  OAI21_X1 U21183 ( .B1(n18269), .B2(n17934), .A(n17933), .ZN(n17935) );
  XNOR2_X1 U21184 ( .A(n17935), .B(n18258), .ZN(n18263) );
  OAI21_X1 U21185 ( .B1(n17953), .B2(n18269), .A(n18258), .ZN(n17936) );
  AOI22_X1 U21186 ( .A1(n17963), .A2(n18263), .B1(n17937), .B2(n17936), .ZN(
        n17938) );
  OAI211_X1 U21187 ( .C1(n17941), .C2(n17940), .A(n17939), .B(n17938), .ZN(
        P3_U2820) );
  NOR2_X1 U21188 ( .A1(n17943), .A2(n17942), .ZN(n17944) );
  XNOR2_X1 U21189 ( .A(n17944), .B(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n18273) );
  NOR2_X1 U21190 ( .A1(n18316), .A2(n18912), .ZN(n18272) );
  NOR2_X1 U21191 ( .A1(n17945), .A2(n18418), .ZN(n17946) );
  AOI21_X1 U21192 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n18041), .A(
        n17946), .ZN(n17948) );
  OAI22_X1 U21193 ( .A1(n17949), .A2(n17948), .B1(n18031), .B2(n17947), .ZN(
        n17950) );
  AOI211_X1 U21194 ( .C1(n17963), .C2(n18273), .A(n18272), .B(n17950), .ZN(
        n17951) );
  OAI221_X1 U21195 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n17953), .C1(
        n18269), .C2(n17952), .A(n17951), .ZN(P3_U2821) );
  OAI21_X1 U21196 ( .B1(n17954), .B2(n18006), .A(n18045), .ZN(n17972) );
  AOI22_X1 U21197 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n17972), .B1(
        n17955), .B2(n17763), .ZN(n17968) );
  AOI21_X1 U21198 ( .B1(n17957), .B2(n17960), .A(n17956), .ZN(n18286) );
  OAI21_X1 U21199 ( .B1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n17959), .A(
        n17958), .ZN(n18292) );
  OAI22_X1 U21200 ( .A1(n18050), .A2(n18292), .B1(n17961), .B2(n17960), .ZN(
        n17962) );
  AOI21_X1 U21201 ( .B1(n17963), .B2(n18286), .A(n17962), .ZN(n17967) );
  NAND2_X1 U21202 ( .A1(n18096), .A2(P3_REIP_REG_8__SCAN_IN), .ZN(n18281) );
  OAI221_X1 U21203 ( .B1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n17965), .C1(
        n17964), .C2(n17973), .A(n18748), .ZN(n17966) );
  NAND4_X1 U21204 ( .A1(n17968), .A2(n17967), .A3(n18281), .A4(n17966), .ZN(
        P3_U2822) );
  OAI21_X1 U21205 ( .B1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n17970), .A(
        n17969), .ZN(n18300) );
  OR2_X1 U21206 ( .A1(n17971), .A2(n18418), .ZN(n17983) );
  NOR2_X1 U21207 ( .A1(n17989), .A2(n17983), .ZN(n17974) );
  NOR2_X1 U21208 ( .A1(n18316), .A2(n18909), .ZN(n18297) );
  AOI221_X1 U21209 ( .B1(n17974), .B2(n17973), .C1(n17972), .C2(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A(n18297), .ZN(n17981) );
  AOI21_X1 U21210 ( .B1(n17977), .B2(n17976), .A(n17975), .ZN(n17978) );
  XNOR2_X1 U21211 ( .A(n17978), .B(n18295), .ZN(n18298) );
  AOI22_X1 U21212 ( .A1(n18039), .A2(n18298), .B1(n17979), .B2(n17763), .ZN(
        n17980) );
  OAI211_X1 U21213 ( .C1(n18049), .C2(n18300), .A(n17981), .B(n17980), .ZN(
        P3_U2823) );
  NAND2_X1 U21214 ( .A1(n18041), .A2(n17983), .ZN(n17998) );
  OAI22_X1 U21215 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n17983), .B1(
        n18049), .B2(n17982), .ZN(n17987) );
  OAI22_X1 U21216 ( .A1(n18031), .A2(n17985), .B1(n18050), .B2(n17984), .ZN(
        n17986) );
  AOI211_X1 U21217 ( .C1(n18096), .C2(P3_REIP_REG_6__SCAN_IN), .A(n17987), .B(
        n17986), .ZN(n17988) );
  OAI21_X1 U21218 ( .B1(n17989), .B2(n17998), .A(n17988), .ZN(P3_U2824) );
  OAI21_X1 U21219 ( .B1(n17992), .B2(n17991), .A(n17990), .ZN(n18302) );
  AOI21_X1 U21220 ( .B1(n17993), .B2(n18045), .A(
        P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n17999) );
  OAI21_X1 U21221 ( .B1(n17996), .B2(n17995), .A(n17994), .ZN(n17997) );
  XNOR2_X1 U21222 ( .A(n17997), .B(n18308), .ZN(n18303) );
  OAI22_X1 U21223 ( .A1(n17999), .A2(n17998), .B1(n18049), .B2(n18303), .ZN(
        n18000) );
  AOI21_X1 U21224 ( .B1(n18001), .B2(n17763), .A(n18000), .ZN(n18002) );
  NAND2_X1 U21225 ( .A1(n18096), .A2(P3_REIP_REG_5__SCAN_IN), .ZN(n18306) );
  OAI211_X1 U21226 ( .C1(n18050), .C2(n18302), .A(n18002), .B(n18306), .ZN(
        P3_U2825) );
  OAI21_X1 U21227 ( .B1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n18004), .A(
        n18003), .ZN(n18323) );
  AOI22_X1 U21228 ( .A1(n18096), .A2(P3_REIP_REG_4__SCAN_IN), .B1(n18748), 
        .B2(n18005), .ZN(n18013) );
  OAI21_X1 U21229 ( .B1(n18007), .B2(n18006), .A(n18045), .ZN(n18022) );
  AOI21_X1 U21230 ( .B1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n18009), .A(
        n18008), .ZN(n18317) );
  OAI22_X1 U21231 ( .A1(n18031), .A2(n18010), .B1(n18317), .B2(n18049), .ZN(
        n18011) );
  AOI21_X1 U21232 ( .B1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n18022), .A(
        n18011), .ZN(n18012) );
  OAI211_X1 U21233 ( .C1(n18050), .C2(n18323), .A(n18013), .B(n18012), .ZN(
        P3_U2826) );
  OAI21_X1 U21234 ( .B1(n18016), .B2(n18015), .A(n18014), .ZN(n18325) );
  NOR2_X1 U21235 ( .A1(n18034), .A2(n18033), .ZN(n18021) );
  OAI22_X1 U21236 ( .A1(n18031), .A2(n18019), .B1(n18049), .B2(n18332), .ZN(
        n18020) );
  AOI221_X1 U21237 ( .B1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n18022), .C1(
        n18021), .C2(n18022), .A(n18020), .ZN(n18023) );
  NAND2_X1 U21238 ( .A1(n18096), .A2(P3_REIP_REG_3__SCAN_IN), .ZN(n18330) );
  OAI211_X1 U21239 ( .C1(n18050), .C2(n18325), .A(n18023), .B(n18330), .ZN(
        P3_U2827) );
  OAI21_X1 U21240 ( .B1(n18026), .B2(n18025), .A(n18024), .ZN(n18342) );
  OAI21_X1 U21241 ( .B1(n18029), .B2(n18028), .A(n18027), .ZN(n18347) );
  OAI22_X1 U21242 ( .A1(n18031), .A2(n18030), .B1(n18049), .B2(n18347), .ZN(
        n18032) );
  AOI221_X1 U21243 ( .B1(n18034), .B2(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .C1(
        n18748), .C2(n18033), .A(n18032), .ZN(n18035) );
  NAND2_X1 U21244 ( .A1(n18096), .A2(P3_REIP_REG_2__SCAN_IN), .ZN(n18345) );
  OAI211_X1 U21245 ( .C1(n18050), .C2(n18342), .A(n18035), .B(n18345), .ZN(
        P3_U2828) );
  OAI21_X1 U21246 ( .B1(n18037), .B2(n18044), .A(n18036), .ZN(n18357) );
  NAND2_X1 U21247 ( .A1(n18977), .A2(n10364), .ZN(n18038) );
  XNOR2_X1 U21248 ( .A(n18038), .B(n18037), .ZN(n18354) );
  AOI22_X1 U21249 ( .A1(n18039), .A2(n18354), .B1(n18096), .B2(
        P3_REIP_REG_1__SCAN_IN), .ZN(n18043) );
  AOI22_X1 U21250 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18041), .B1(
        n17763), .B2(n18040), .ZN(n18042) );
  OAI211_X1 U21251 ( .C1(n18049), .C2(n18357), .A(n18043), .B(n18042), .ZN(
        P3_U2829) );
  AOI21_X1 U21252 ( .B1(n10364), .B2(n18977), .A(n18044), .ZN(n18361) );
  INV_X1 U21253 ( .A(n18361), .ZN(n18363) );
  NAND3_X1 U21254 ( .A1(n18994), .A2(n18046), .A3(n18045), .ZN(n18047) );
  AOI22_X1 U21255 ( .A1(n18096), .A2(P3_REIP_REG_0__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n18047), .ZN(n18048) );
  OAI221_X1 U21256 ( .B1(n18361), .B2(n18050), .C1(n18363), .C2(n18049), .A(
        n18048), .ZN(P3_U2830) );
  NAND2_X1 U21257 ( .A1(n18052), .A2(n18051), .ZN(n18119) );
  NAND3_X1 U21258 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n18120), .A3(
        n18119), .ZN(n18105) );
  OAI21_X1 U21259 ( .B1(n18053), .B2(n18105), .A(n10180), .ZN(n18065) );
  AOI21_X1 U21260 ( .B1(n18824), .B2(n18054), .A(n10180), .ZN(n18063) );
  NOR2_X1 U21261 ( .A1(n18831), .A2(n18813), .ZN(n18348) );
  OAI22_X1 U21262 ( .A1(n18837), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B1(
        n18055), .B2(n18348), .ZN(n18062) );
  NAND2_X1 U21263 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n18057) );
  OAI21_X1 U21264 ( .B1(n18164), .B2(n18056), .A(n18313), .ZN(n18093) );
  AOI21_X1 U21265 ( .B1(n18333), .B2(n18057), .A(n18093), .ZN(n18076) );
  INV_X1 U21266 ( .A(n18113), .ZN(n18242) );
  AOI22_X1 U21267 ( .A1(n18244), .A2(n18059), .B1(n18242), .B2(n18058), .ZN(
        n18060) );
  NAND2_X1 U21268 ( .A1(n18076), .A2(n18060), .ZN(n18061) );
  OAI21_X1 U21269 ( .B1(n18062), .B2(n18061), .A(n18359), .ZN(n18071) );
  OAI21_X1 U21270 ( .B1(n18063), .B2(n18349), .A(n18071), .ZN(n18064) );
  AOI22_X1 U21271 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n18344), .B1(
        n18065), .B2(n18064), .ZN(n18067) );
  NAND2_X1 U21272 ( .A1(n18096), .A2(P3_REIP_REG_27__SCAN_IN), .ZN(n18066) );
  OAI211_X1 U21273 ( .C1(n18068), .C2(n18211), .A(n18067), .B(n18066), .ZN(
        P3_U2835) );
  INV_X1 U21274 ( .A(n18148), .ZN(n18151) );
  AOI22_X1 U21275 ( .A1(n18287), .A2(n18070), .B1(n18151), .B2(n18069), .ZN(
        n18074) );
  INV_X1 U21276 ( .A(n18071), .ZN(n18072) );
  OAI21_X1 U21277 ( .B1(n18344), .B2(n18072), .A(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n18073) );
  OAI211_X1 U21278 ( .C1(n18943), .C2(n18316), .A(n18074), .B(n18073), .ZN(
        P3_U2836) );
  INV_X1 U21279 ( .A(n18075), .ZN(n18080) );
  INV_X1 U21280 ( .A(n18076), .ZN(n18078) );
  NOR2_X1 U21281 ( .A1(n18078), .A2(n18077), .ZN(n18079) );
  MUX2_X1 U21282 ( .A(n18080), .B(n18079), .S(
        P3_INSTADDRPOINTER_REG_25__SCAN_IN), .Z(n18082) );
  OAI21_X1 U21283 ( .B1(n18349), .B2(n18082), .A(n18081), .ZN(n18086) );
  OAI22_X1 U21284 ( .A1(n18326), .A2(n18084), .B1(n18211), .B2(n18083), .ZN(
        n18085) );
  AOI211_X1 U21285 ( .C1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .C2(n18344), .A(
        n18086), .B(n18085), .ZN(n18087) );
  OAI21_X1 U21286 ( .B1(n18089), .B2(n18088), .A(n18087), .ZN(P3_U2837) );
  OAI22_X1 U21287 ( .A1(n18091), .A2(n18113), .B1(n18090), .B2(n18806), .ZN(
        n18092) );
  NOR3_X1 U21288 ( .A1(n18344), .A2(n18093), .A3(n18092), .ZN(n18099) );
  AOI221_X1 U21289 ( .B1(n18095), .B2(n18831), .C1(n18158), .C2(n18831), .A(
        n18094), .ZN(n18097) );
  AOI21_X1 U21290 ( .B1(n18099), .B2(n18097), .A(n18096), .ZN(n18106) );
  AOI21_X1 U21291 ( .B1(n18280), .B2(n18099), .A(n18098), .ZN(n18100) );
  AOI22_X1 U21292 ( .A1(n18287), .A2(n18101), .B1(n18106), .B2(n18100), .ZN(
        n18103) );
  NAND2_X1 U21293 ( .A1(n18096), .A2(P3_REIP_REG_24__SCAN_IN), .ZN(n18102) );
  OAI211_X1 U21294 ( .C1(n18104), .C2(n18148), .A(n18103), .B(n18102), .ZN(
        P3_U2838) );
  NOR2_X1 U21295 ( .A1(n18344), .A2(n18105), .ZN(n18107) );
  OAI21_X1 U21296 ( .B1(n18107), .B2(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n18106), .ZN(n18108) );
  OAI211_X1 U21297 ( .C1(n18110), .C2(n18211), .A(n18109), .B(n18108), .ZN(
        P3_U2839) );
  INV_X1 U21298 ( .A(n18111), .ZN(n18157) );
  AOI21_X1 U21299 ( .B1(n18157), .B2(n18141), .A(n18837), .ZN(n18112) );
  AOI221_X1 U21300 ( .B1(n18158), .B2(n18831), .C1(n18128), .C2(n18831), .A(
        n18112), .ZN(n18140) );
  NAND2_X1 U21301 ( .A1(n18806), .A2(n18113), .ZN(n18248) );
  AOI22_X1 U21302 ( .A1(n18824), .A2(n18115), .B1(n18114), .B2(n18248), .ZN(
        n18116) );
  NAND2_X1 U21303 ( .A1(n18140), .A2(n18116), .ZN(n18134) );
  OAI22_X1 U21304 ( .A1(n18222), .A2(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .B1(
        n18132), .B2(n18807), .ZN(n18117) );
  NOR4_X1 U21305 ( .A1(n18118), .A2(n18127), .A3(n18134), .A4(n18117), .ZN(
        n18122) );
  AOI22_X1 U21306 ( .A1(n18244), .A2(n18194), .B1(n18242), .B2(n18188), .ZN(
        n18130) );
  NAND2_X1 U21307 ( .A1(n18120), .A2(n18119), .ZN(n18121) );
  AOI22_X1 U21308 ( .A1(n18122), .A2(n18130), .B1(n18127), .B2(n18121), .ZN(
        n18124) );
  AOI22_X1 U21309 ( .A1(n18359), .A2(n18124), .B1(n18287), .B2(n18123), .ZN(
        n18126) );
  OAI211_X1 U21310 ( .C1(n18350), .C2(n18127), .A(n18126), .B(n18125), .ZN(
        P3_U2840) );
  INV_X1 U21311 ( .A(n18128), .ZN(n18129) );
  AOI21_X1 U21312 ( .B1(n18179), .B2(n18129), .A(n18821), .ZN(n18131) );
  NAND2_X1 U21313 ( .A1(n18359), .A2(n18130), .ZN(n18180) );
  NOR2_X1 U21314 ( .A1(n18131), .A2(n18180), .ZN(n18139) );
  OAI21_X1 U21315 ( .B1(n18132), .B2(n18348), .A(n18139), .ZN(n18133) );
  OAI21_X1 U21316 ( .B1(n18134), .B2(n18133), .A(
        P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n18138) );
  AOI22_X1 U21317 ( .A1(n18287), .A2(n18136), .B1(n18151), .B2(n18135), .ZN(
        n18137) );
  OAI221_X1 U21318 ( .B1(n18096), .B2(n18138), .C1(n18316), .C2(n18933), .A(
        n18137), .ZN(P3_U2841) );
  NAND2_X1 U21319 ( .A1(n18156), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n18143) );
  INV_X1 U21320 ( .A(n18248), .ZN(n18159) );
  OAI211_X1 U21321 ( .C1(n18141), .C2(n18159), .A(n18140), .B(n18139), .ZN(
        n18142) );
  NAND2_X1 U21322 ( .A1(n18316), .A2(n18142), .ZN(n18155) );
  OAI21_X1 U21323 ( .B1(n18348), .B2(n18143), .A(n18155), .ZN(n18145) );
  AOI22_X1 U21324 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n18145), .B1(
        n18287), .B2(n18144), .ZN(n18147) );
  NAND2_X1 U21325 ( .A1(n18096), .A2(P3_REIP_REG_20__SCAN_IN), .ZN(n18146) );
  OAI211_X1 U21326 ( .C1(n18149), .C2(n18148), .A(n18147), .B(n18146), .ZN(
        P3_U2842) );
  AOI22_X1 U21327 ( .A1(n18287), .A2(n18152), .B1(n18151), .B2(n18150), .ZN(
        n18154) );
  OAI211_X1 U21328 ( .C1(n18156), .C2(n18155), .A(n18154), .B(n18153), .ZN(
        P3_U2843) );
  NAND3_X1 U21329 ( .A1(n18157), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        n18313), .ZN(n18163) );
  NAND2_X1 U21330 ( .A1(n18831), .A2(n18158), .ZN(n18160) );
  AOI22_X1 U21331 ( .A1(n18161), .A2(n18160), .B1(n18159), .B2(n18807), .ZN(
        n18162) );
  AOI211_X1 U21332 ( .C1(n18333), .C2(n18163), .A(n18162), .B(n18180), .ZN(
        n18175) );
  AOI221_X1 U21333 ( .B1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n18175), 
        .C1(n18164), .C2(n18175), .A(n18096), .ZN(n18166) );
  AOI22_X1 U21334 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n18166), .B1(
        n18182), .B2(n18165), .ZN(n18168) );
  OAI211_X1 U21335 ( .C1(n18211), .C2(n18169), .A(n18168), .B(n18167), .ZN(
        P3_U2844) );
  NAND2_X1 U21336 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n18316), .ZN(
        n18174) );
  AOI22_X1 U21337 ( .A1(n18287), .A2(n18171), .B1(n18182), .B2(n18170), .ZN(
        n18173) );
  OAI211_X1 U21338 ( .C1(n18175), .C2(n18174), .A(n18173), .B(n18172), .ZN(
        P3_U2845) );
  INV_X1 U21339 ( .A(n18222), .ZN(n18256) );
  NAND2_X1 U21340 ( .A1(n18831), .A2(n18176), .ZN(n18245) );
  OAI21_X1 U21341 ( .B1(n18837), .B2(n18239), .A(n18245), .ZN(n18220) );
  AOI21_X1 U21342 ( .B1(n18256), .B2(n18177), .A(n18220), .ZN(n18178) );
  OAI211_X1 U21343 ( .C1(n18179), .C2(n18821), .A(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B(n18178), .ZN(n18187) );
  OAI221_X1 U21344 ( .B1(n18180), .B2(n18276), .C1(n18180), .C2(n18187), .A(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n18185) );
  INV_X1 U21345 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n18923) );
  AOI22_X1 U21346 ( .A1(n18287), .A2(n18183), .B1(n18182), .B2(n18181), .ZN(
        n18184) );
  OAI221_X1 U21347 ( .B1(n18096), .B2(n18185), .C1(n18316), .C2(n18923), .A(
        n18184), .ZN(P3_U2846) );
  NOR2_X1 U21348 ( .A1(n18186), .A2(n18200), .ZN(n18201) );
  OAI221_X1 U21349 ( .B1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .C1(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n18201), .A(n18187), .ZN(
        n18191) );
  OAI211_X1 U21350 ( .C1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n18189), .A(
        n18242), .B(n18188), .ZN(n18190) );
  AOI21_X1 U21351 ( .B1(n18191), .B2(n18190), .A(n18349), .ZN(n18193) );
  AOI211_X1 U21352 ( .C1(n18344), .C2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n18193), .B(n18192), .ZN(n18197) );
  OAI211_X1 U21353 ( .C1(n18195), .C2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n18364), .B(n18194), .ZN(n18196) );
  OAI211_X1 U21354 ( .C1(n18198), .C2(n18211), .A(n18197), .B(n18196), .ZN(
        P3_U2847) );
  INV_X1 U21355 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n21228) );
  NOR2_X1 U21356 ( .A1(n18316), .A2(n21228), .ZN(n18206) );
  INV_X1 U21357 ( .A(n18199), .ZN(n18265) );
  AOI21_X1 U21358 ( .B1(n18228), .B2(n18265), .A(n18821), .ZN(n18224) );
  AOI211_X1 U21359 ( .C1(n18276), .C2(n18200), .A(n18224), .B(n18220), .ZN(
        n18204) );
  INV_X1 U21360 ( .A(n18201), .ZN(n18203) );
  AOI221_X1 U21361 ( .B1(n18204), .B2(P3_INSTADDRPOINTER_REG_14__SCAN_IN), 
        .C1(n18203), .C2(n18202), .A(n18349), .ZN(n18205) );
  AOI211_X1 U21362 ( .C1(n18344), .C2(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n18206), .B(n18205), .ZN(n18210) );
  AOI22_X1 U21363 ( .A1(n18288), .A2(n18208), .B1(n18364), .B2(n18207), .ZN(
        n18209) );
  OAI211_X1 U21364 ( .C1(n18212), .C2(n18211), .A(n18210), .B(n18209), .ZN(
        P3_U2848) );
  AND2_X1 U21365 ( .A1(n18359), .A2(n18213), .ZN(n18284) );
  AOI222_X1 U21366 ( .A1(n18215), .A2(n18364), .B1(n18288), .B2(n18214), .C1(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .C2(n18284), .ZN(n18275) );
  AOI22_X1 U21367 ( .A1(n18096), .A2(P3_REIP_REG_13__SCAN_IN), .B1(n18287), 
        .B2(n18216), .ZN(n18226) );
  AOI22_X1 U21368 ( .A1(n18217), .A2(n18242), .B1(n18256), .B2(n18250), .ZN(
        n18218) );
  INV_X1 U21369 ( .A(n18218), .ZN(n18219) );
  AOI211_X1 U21370 ( .C1(n18244), .C2(n18221), .A(n18220), .B(n18219), .ZN(
        n18229) );
  OAI211_X1 U21371 ( .C1(n18222), .C2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n18359), .B(n18229), .ZN(n18223) );
  OAI211_X1 U21372 ( .C1(n18224), .C2(n18223), .A(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B(n18316), .ZN(n18225) );
  OAI211_X1 U21373 ( .C1(n18275), .C2(n18227), .A(n18226), .B(n18225), .ZN(
        P3_U2849) );
  AND2_X1 U21374 ( .A1(n18228), .A2(n18265), .ZN(n18230) );
  OAI211_X1 U21375 ( .C1(n18230), .C2(n18821), .A(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B(n18229), .ZN(n18232) );
  OAI22_X1 U21376 ( .A1(n18275), .A2(n18250), .B1(n18237), .B2(n18349), .ZN(
        n18231) );
  AOI22_X1 U21377 ( .A1(n18287), .A2(n18233), .B1(n18232), .B2(n18231), .ZN(
        n18236) );
  INV_X1 U21378 ( .A(n18234), .ZN(n18235) );
  OAI211_X1 U21379 ( .C1(n18350), .C2(n18237), .A(n18236), .B(n18235), .ZN(
        P3_U2850) );
  AOI22_X1 U21380 ( .A1(n18096), .A2(P3_REIP_REG_11__SCAN_IN), .B1(n18287), 
        .B2(n18238), .ZN(n18254) );
  NOR2_X1 U21381 ( .A1(n18837), .A2(n18239), .ZN(n18257) );
  INV_X1 U21382 ( .A(n18240), .ZN(n18249) );
  AOI21_X1 U21383 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18265), .A(
        n18821), .ZN(n18247) );
  AOI22_X1 U21384 ( .A1(n18244), .A2(n18243), .B1(n18242), .B2(n18241), .ZN(
        n18246) );
  NAND3_X1 U21385 ( .A1(n18359), .A2(n18246), .A3(n18245), .ZN(n18266) );
  AOI211_X1 U21386 ( .C1(n18249), .C2(n18248), .A(n18247), .B(n18266), .ZN(
        n18260) );
  NAND2_X1 U21387 ( .A1(n18256), .A2(n18250), .ZN(n18251) );
  OAI211_X1 U21388 ( .C1(n18821), .C2(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n18260), .B(n18251), .ZN(n18252) );
  OAI211_X1 U21389 ( .C1(n18257), .C2(n18252), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n18316), .ZN(n18253) );
  OAI211_X1 U21390 ( .C1(n18275), .C2(n18255), .A(n18254), .B(n18253), .ZN(
        P3_U2851) );
  OAI21_X1 U21391 ( .B1(n18257), .B2(n18269), .A(n18256), .ZN(n18259) );
  AOI211_X1 U21392 ( .C1(n18260), .C2(n18259), .A(n18096), .B(n18258), .ZN(
        n18262) );
  NOR3_X1 U21393 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n18275), .A3(
        n18269), .ZN(n18261) );
  AOI211_X1 U21394 ( .C1(n18287), .C2(n18263), .A(n18262), .B(n18261), .ZN(
        n18264) );
  OAI21_X1 U21395 ( .B1(n18316), .B2(n18914), .A(n18264), .ZN(P3_U2852) );
  AOI221_X1 U21396 ( .B1(n18837), .B2(n18821), .C1(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .C2(n18821), .A(n18265), .ZN(
        n18267) );
  AOI211_X1 U21397 ( .C1(n18824), .C2(n18268), .A(n18267), .B(n18266), .ZN(
        n18270) );
  NOR3_X1 U21398 ( .A1(n18096), .A2(n18270), .A3(n18269), .ZN(n18271) );
  AOI211_X1 U21399 ( .C1(n18287), .C2(n18273), .A(n18272), .B(n18271), .ZN(
        n18274) );
  OAI21_X1 U21400 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18275), .A(
        n18274), .ZN(P3_U2853) );
  AOI21_X1 U21401 ( .B1(n18276), .B2(n13750), .A(n18295), .ZN(n18277) );
  AOI21_X1 U21402 ( .B1(n18278), .B2(n18277), .A(n18349), .ZN(n18279) );
  NOR2_X1 U21403 ( .A1(n18344), .A2(n18279), .ZN(n18293) );
  AOI21_X1 U21404 ( .B1(n18280), .B2(n18350), .A(n18293), .ZN(n18285) );
  INV_X1 U21405 ( .A(n18281), .ZN(n18282) );
  AOI221_X1 U21406 ( .B1(n18285), .B2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .C1(
        n18284), .C2(n18283), .A(n18282), .ZN(n18291) );
  AOI22_X1 U21407 ( .A1(n18289), .A2(n18288), .B1(n18287), .B2(n18286), .ZN(
        n18290) );
  OAI211_X1 U21408 ( .C1(n18326), .C2(n18292), .A(n18291), .B(n18290), .ZN(
        P3_U2854) );
  AOI221_X1 U21409 ( .B1(n18349), .B2(n18295), .C1(n18294), .C2(n18295), .A(
        n18293), .ZN(n18296) );
  AOI211_X1 U21410 ( .C1(n18298), .C2(n18364), .A(n18297), .B(n18296), .ZN(
        n18299) );
  OAI21_X1 U21411 ( .B1(n18358), .B2(n18300), .A(n18299), .ZN(P3_U2855) );
  INV_X1 U21412 ( .A(n18301), .ZN(n18309) );
  NOR3_X1 U21413 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n18311), .A3(
        n18310), .ZN(n18305) );
  OAI22_X1 U21414 ( .A1(n18358), .A2(n18303), .B1(n18326), .B2(n18302), .ZN(
        n18304) );
  AOI21_X1 U21415 ( .B1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n18305), .A(
        n18304), .ZN(n18307) );
  OAI211_X1 U21416 ( .C1(n18309), .C2(n18308), .A(n18307), .B(n18306), .ZN(
        P3_U2857) );
  NOR2_X1 U21417 ( .A1(n18311), .A2(n18310), .ZN(n18321) );
  INV_X1 U21418 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n18320) );
  NAND2_X1 U21419 ( .A1(n18831), .A2(n18312), .ZN(n18340) );
  NAND3_X1 U21420 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n18313), .A3(
        n18340), .ZN(n18314) );
  AOI21_X1 U21421 ( .B1(n18333), .B2(n18315), .A(n18314), .ZN(n18328) );
  OAI21_X1 U21422 ( .B1(n18328), .B2(n18351), .A(n18350), .ZN(n18319) );
  OAI22_X1 U21423 ( .A1(n18317), .A2(n18358), .B1(n18316), .B2(n18903), .ZN(
        n18318) );
  AOI221_X1 U21424 ( .B1(n18321), .B2(n18320), .C1(n18319), .C2(
        P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A(n18318), .ZN(n18322) );
  OAI21_X1 U21425 ( .B1(n18326), .B2(n18323), .A(n18322), .ZN(P3_U2858) );
  OAI21_X1 U21426 ( .B1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n18324), .A(
        n18359), .ZN(n18327) );
  OAI22_X1 U21427 ( .A1(n18328), .A2(n18327), .B1(n18326), .B2(n18325), .ZN(
        n18329) );
  AOI21_X1 U21428 ( .B1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n18344), .A(
        n18329), .ZN(n18331) );
  OAI211_X1 U21429 ( .C1(n18332), .C2(n18358), .A(n18331), .B(n18330), .ZN(
        P3_U2859) );
  NAND2_X1 U21430 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18336) );
  INV_X1 U21431 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18976) );
  OAI21_X1 U21432 ( .B1(n18334), .B2(n18976), .A(n18333), .ZN(n18335) );
  OAI21_X1 U21433 ( .B1(n18336), .B2(n18807), .A(n18335), .ZN(n18339) );
  NOR2_X1 U21434 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n18337), .ZN(
        n18338) );
  AOI22_X1 U21435 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n18339), .B1(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n18338), .ZN(n18341) );
  OAI211_X1 U21436 ( .C1(n18342), .C2(n18806), .A(n18341), .B(n18340), .ZN(
        n18343) );
  AOI22_X1 U21437 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n18344), .B1(
        n18359), .B2(n18343), .ZN(n18346) );
  OAI211_X1 U21438 ( .C1(n18347), .C2(n18358), .A(n18346), .B(n18345), .ZN(
        P3_U2860) );
  OR3_X1 U21439 ( .A1(n18349), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A3(
        n18348), .ZN(n18365) );
  AOI21_X1 U21440 ( .B1(n18350), .B2(n18365), .A(n18976), .ZN(n18353) );
  AOI211_X1 U21441 ( .C1(n18837), .C2(n18977), .A(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B(n18351), .ZN(n18352) );
  AOI211_X1 U21442 ( .C1(n18364), .C2(n18354), .A(n18353), .B(n18352), .ZN(
        n18356) );
  NAND2_X1 U21443 ( .A1(n18096), .A2(P3_REIP_REG_1__SCAN_IN), .ZN(n18355) );
  OAI211_X1 U21444 ( .C1(n18357), .C2(n18358), .A(n18356), .B(n18355), .ZN(
        P3_U2861) );
  INV_X1 U21445 ( .A(P3_REIP_REG_0__SCAN_IN), .ZN(n19005) );
  INV_X1 U21446 ( .A(n18358), .ZN(n18362) );
  AOI211_X1 U21447 ( .C1(n18837), .C2(n18359), .A(n18096), .B(n18977), .ZN(
        n18360) );
  AOI221_X1 U21448 ( .B1(n18364), .B2(n18363), .C1(n18362), .C2(n18361), .A(
        n18360), .ZN(n18366) );
  OAI211_X1 U21449 ( .C1(n19005), .C2(n18316), .A(n18366), .B(n18365), .ZN(
        P3_U2862) );
  AOI21_X1 U21450 ( .B1(n18369), .B2(n18368), .A(n18367), .ZN(n18859) );
  OAI21_X1 U21451 ( .B1(n18859), .B2(n18423), .A(n18374), .ZN(n18370) );
  OAI221_X1 U21452 ( .B1(n18621), .B2(n19019), .C1(n18621), .C2(n18374), .A(
        n18370), .ZN(P3_U2863) );
  NOR2_X1 U21453 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18845), .ZN(
        n18556) );
  NOR2_X1 U21454 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18846), .ZN(
        n18645) );
  NOR2_X1 U21455 ( .A1(n18556), .A2(n18645), .ZN(n18372) );
  OAI22_X1 U21456 ( .A1(n18373), .A2(n18846), .B1(n18372), .B2(n18371), .ZN(
        P3_U2866) );
  NOR2_X1 U21457 ( .A1(n18847), .A2(n18374), .ZN(P3_U2867) );
  INV_X1 U21458 ( .A(n18375), .ZN(n18376) );
  NOR2_X1 U21459 ( .A1(n18377), .A2(n18376), .ZN(n18414) );
  NOR2_X1 U21460 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18826) );
  NAND2_X1 U21461 ( .A1(n18845), .A2(n18846), .ZN(n18444) );
  INV_X1 U21462 ( .A(n18444), .ZN(n18466) );
  NAND2_X1 U21463 ( .A1(n18826), .A2(n18466), .ZN(n18422) );
  NOR2_X2 U21464 ( .A1(n18379), .A2(n18418), .ZN(n18744) );
  NAND2_X1 U21465 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18620), .ZN(
        n18508) );
  NAND2_X1 U21466 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18691) );
  NOR2_X2 U21467 ( .A1(n18508), .A2(n18691), .ZN(n18793) );
  NOR2_X2 U21468 ( .A1(n18415), .A2(n18380), .ZN(n18743) );
  NOR2_X1 U21469 ( .A1(n18620), .A2(n18621), .ZN(n18825) );
  INV_X1 U21470 ( .A(n18825), .ZN(n18381) );
  NOR2_X2 U21471 ( .A1(n18381), .A2(n18691), .ZN(n18742) );
  NOR2_X1 U21472 ( .A1(n18742), .A2(n18482), .ZN(n18445) );
  NOR2_X1 U21473 ( .A1(n18715), .A2(n18445), .ZN(n18417) );
  AOI22_X1 U21474 ( .A1(n18744), .A2(n18793), .B1(n18743), .B2(n18417), .ZN(
        n18386) );
  NOR2_X1 U21475 ( .A1(n18846), .A2(n18531), .ZN(n18746) );
  NAND2_X1 U21476 ( .A1(n18746), .A2(n18621), .ZN(n18741) );
  NAND2_X1 U21477 ( .A1(n18741), .A2(n18713), .ZN(n18714) );
  AOI21_X1 U21478 ( .B1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(
        P3_STATE2_REG_3__SCAN_IN), .A(n18415), .ZN(n18383) );
  INV_X1 U21479 ( .A(n18445), .ZN(n18382) );
  AOI22_X1 U21480 ( .A1(n18748), .A2(n18714), .B1(n18383), .B2(n18382), .ZN(
        n18419) );
  NOR2_X2 U21481 ( .A1(n18418), .A2(n18384), .ZN(n18749) );
  AOI22_X1 U21482 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n18419), .B1(
        n18749), .B2(n18721), .ZN(n18385) );
  OAI211_X1 U21483 ( .C1(n18752), .C2(n18422), .A(n18386), .B(n18385), .ZN(
        P3_U2868) );
  NOR2_X2 U21484 ( .A1(n18415), .A2(n18388), .ZN(n18753) );
  NOR2_X2 U21485 ( .A1(n18418), .A2(n18389), .ZN(n18755) );
  AOI22_X1 U21486 ( .A1(n18753), .A2(n18417), .B1(n18755), .B2(n18721), .ZN(
        n18392) );
  NOR2_X2 U21487 ( .A1(n18390), .A2(n18418), .ZN(n18754) );
  AOI22_X1 U21488 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n18419), .B1(
        n18754), .B2(n18793), .ZN(n18391) );
  OAI211_X1 U21489 ( .C1(n18758), .C2(n18422), .A(n18392), .B(n18391), .ZN(
        P3_U2869) );
  NAND2_X1 U21490 ( .A1(n18414), .A2(n18393), .ZN(n18764) );
  NOR2_X2 U21491 ( .A1(n18418), .A2(n19385), .ZN(n18761) );
  NOR2_X2 U21492 ( .A1(n18415), .A2(n18394), .ZN(n18759) );
  AOI22_X1 U21493 ( .A1(n18761), .A2(n18721), .B1(n18759), .B2(n18417), .ZN(
        n18396) );
  NOR2_X2 U21494 ( .A1(n19382), .A2(n18418), .ZN(n18760) );
  AOI22_X1 U21495 ( .A1(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n18419), .B1(
        n18760), .B2(n18793), .ZN(n18395) );
  OAI211_X1 U21496 ( .C1(n18764), .C2(n18422), .A(n18396), .B(n18395), .ZN(
        P3_U2870) );
  NAND2_X1 U21497 ( .A1(n18414), .A2(n18397), .ZN(n18770) );
  NOR2_X2 U21498 ( .A1(n18415), .A2(n18398), .ZN(n18765) );
  NOR2_X2 U21499 ( .A1(n19389), .A2(n18418), .ZN(n18767) );
  AOI22_X1 U21500 ( .A1(n18765), .A2(n18417), .B1(n18767), .B2(n18793), .ZN(
        n18400) );
  NOR2_X2 U21501 ( .A1(n18418), .A2(n19392), .ZN(n18766) );
  AOI22_X1 U21502 ( .A1(P3_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n18419), .B1(
        n18766), .B2(n18721), .ZN(n18399) );
  OAI211_X1 U21503 ( .C1(n18770), .C2(n18422), .A(n18400), .B(n18399), .ZN(
        P3_U2871) );
  NOR2_X2 U21504 ( .A1(n19397), .A2(n18418), .ZN(n18772) );
  NOR2_X2 U21505 ( .A1(n18415), .A2(n18402), .ZN(n18771) );
  AOI22_X1 U21506 ( .A1(n18772), .A2(n18793), .B1(n18771), .B2(n18417), .ZN(
        n18404) );
  NOR2_X2 U21507 ( .A1(n18418), .A2(n19399), .ZN(n18773) );
  AOI22_X1 U21508 ( .A1(P3_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n18419), .B1(
        n18773), .B2(n18721), .ZN(n18403) );
  OAI211_X1 U21509 ( .C1(n18776), .C2(n18422), .A(n18404), .B(n18403), .ZN(
        P3_U2872) );
  NOR2_X2 U21510 ( .A1(n18418), .A2(n21192), .ZN(n18778) );
  NOR2_X2 U21511 ( .A1(n18415), .A2(n18406), .ZN(n18777) );
  AOI22_X1 U21512 ( .A1(n18778), .A2(n18721), .B1(n18777), .B2(n18417), .ZN(
        n18408) );
  NOR2_X2 U21513 ( .A1(n19405), .A2(n18418), .ZN(n18779) );
  AOI22_X1 U21514 ( .A1(P3_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n18419), .B1(
        n18779), .B2(n18793), .ZN(n18407) );
  OAI211_X1 U21515 ( .C1(n18782), .C2(n18422), .A(n18408), .B(n18407), .ZN(
        P3_U2873) );
  NAND2_X1 U21516 ( .A1(n18414), .A2(n18409), .ZN(n18788) );
  NOR2_X2 U21517 ( .A1(n18418), .A2(n19413), .ZN(n18785) );
  NOR2_X2 U21518 ( .A1(n18415), .A2(n18410), .ZN(n18784) );
  AOI22_X1 U21519 ( .A1(n18785), .A2(n18721), .B1(n18784), .B2(n18417), .ZN(
        n18412) );
  NOR2_X2 U21520 ( .A1(n19411), .A2(n18418), .ZN(n18783) );
  AOI22_X1 U21521 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n18419), .B1(
        n18783), .B2(n18793), .ZN(n18411) );
  OAI211_X1 U21522 ( .C1(n18788), .C2(n18422), .A(n18412), .B(n18411), .ZN(
        P3_U2874) );
  NOR2_X2 U21523 ( .A1(n18416), .A2(n18415), .ZN(n18790) );
  NOR2_X2 U21524 ( .A1(n19423), .A2(n18418), .ZN(n18794) );
  AOI22_X1 U21525 ( .A1(n18790), .A2(n18417), .B1(n18794), .B2(n18721), .ZN(
        n18421) );
  NOR2_X2 U21526 ( .A1(n18418), .A2(n19418), .ZN(n18792) );
  AOI22_X1 U21527 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n18419), .B1(
        n18792), .B2(n18793), .ZN(n18420) );
  OAI211_X1 U21528 ( .C1(n18799), .C2(n18422), .A(n18421), .B(n18420), .ZN(
        P3_U2875) );
  NOR2_X2 U21529 ( .A1(n18444), .A2(n18508), .ZN(n18503) );
  INV_X1 U21530 ( .A(n18715), .ZN(n18868) );
  NAND2_X1 U21531 ( .A1(n18620), .A2(n18868), .ZN(n18690) );
  NOR2_X1 U21532 ( .A1(n18444), .A2(n18690), .ZN(n18439) );
  AOI22_X1 U21533 ( .A1(n18744), .A2(n18721), .B1(n18743), .B2(n18439), .ZN(
        n18426) );
  INV_X1 U21534 ( .A(n18423), .ZN(n18424) );
  NAND2_X1 U21535 ( .A1(n18720), .A2(n18424), .ZN(n18646) );
  NOR2_X1 U21536 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18646), .ZN(
        n18692) );
  AOI22_X1 U21537 ( .A1(n18748), .A2(n18746), .B1(n18466), .B2(n18692), .ZN(
        n18440) );
  AOI22_X1 U21538 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n18440), .B1(
        n18749), .B2(n18742), .ZN(n18425) );
  OAI211_X1 U21539 ( .C1(n18443), .C2(n18752), .A(n18426), .B(n18425), .ZN(
        P3_U2876) );
  AOI22_X1 U21540 ( .A1(n18754), .A2(n18721), .B1(n18753), .B2(n18439), .ZN(
        n18428) );
  AOI22_X1 U21541 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n18440), .B1(
        n18755), .B2(n18742), .ZN(n18427) );
  OAI211_X1 U21542 ( .C1(n18443), .C2(n18758), .A(n18428), .B(n18427), .ZN(
        P3_U2877) );
  AOI22_X1 U21543 ( .A1(n18761), .A2(n18742), .B1(n18759), .B2(n18439), .ZN(
        n18430) );
  AOI22_X1 U21544 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n18440), .B1(
        n18760), .B2(n18721), .ZN(n18429) );
  OAI211_X1 U21545 ( .C1(n18443), .C2(n18764), .A(n18430), .B(n18429), .ZN(
        P3_U2878) );
  AOI22_X1 U21546 ( .A1(n18765), .A2(n18439), .B1(n18767), .B2(n18721), .ZN(
        n18432) );
  AOI22_X1 U21547 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n18440), .B1(
        n18766), .B2(n18742), .ZN(n18431) );
  OAI211_X1 U21548 ( .C1(n18443), .C2(n18770), .A(n18432), .B(n18431), .ZN(
        P3_U2879) );
  AOI22_X1 U21549 ( .A1(n18772), .A2(n18721), .B1(n18771), .B2(n18439), .ZN(
        n18434) );
  AOI22_X1 U21550 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n18440), .B1(
        n18773), .B2(n18742), .ZN(n18433) );
  OAI211_X1 U21551 ( .C1(n18443), .C2(n18776), .A(n18434), .B(n18433), .ZN(
        P3_U2880) );
  AOI22_X1 U21552 ( .A1(n18778), .A2(n18742), .B1(n18777), .B2(n18439), .ZN(
        n18436) );
  AOI22_X1 U21553 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n18440), .B1(
        n18779), .B2(n18721), .ZN(n18435) );
  OAI211_X1 U21554 ( .C1(n18443), .C2(n18782), .A(n18436), .B(n18435), .ZN(
        P3_U2881) );
  AOI22_X1 U21555 ( .A1(n18785), .A2(n18742), .B1(n18784), .B2(n18439), .ZN(
        n18438) );
  AOI22_X1 U21556 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n18440), .B1(
        n18783), .B2(n18721), .ZN(n18437) );
  OAI211_X1 U21557 ( .C1(n18443), .C2(n18788), .A(n18438), .B(n18437), .ZN(
        P3_U2882) );
  AOI22_X1 U21558 ( .A1(n18792), .A2(n18721), .B1(n18790), .B2(n18439), .ZN(
        n18442) );
  AOI22_X1 U21559 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n18440), .B1(
        n18794), .B2(n18742), .ZN(n18441) );
  OAI211_X1 U21560 ( .C1(n18443), .C2(n18799), .A(n18442), .B(n18441), .ZN(
        P3_U2883) );
  NOR2_X1 U21561 ( .A1(n18620), .A2(n18444), .ZN(n18511) );
  NAND2_X1 U21562 ( .A1(n18621), .A2(n18511), .ZN(n18465) );
  INV_X1 U21563 ( .A(n18465), .ZN(n18527) );
  NOR2_X1 U21564 ( .A1(n18527), .A2(n18503), .ZN(n18486) );
  NOR2_X1 U21565 ( .A1(n18715), .A2(n18486), .ZN(n18461) );
  AOI22_X1 U21566 ( .A1(n18744), .A2(n18742), .B1(n18743), .B2(n18461), .ZN(
        n18448) );
  OAI21_X1 U21567 ( .B1(n18445), .B2(n18717), .A(n18486), .ZN(n18446) );
  OAI211_X1 U21568 ( .C1(n18527), .C2(n18967), .A(n18720), .B(n18446), .ZN(
        n18462) );
  AOI22_X1 U21569 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n18462), .B1(
        n18749), .B2(n18482), .ZN(n18447) );
  OAI211_X1 U21570 ( .C1(n18465), .C2(n18752), .A(n18448), .B(n18447), .ZN(
        P3_U2884) );
  AOI22_X1 U21571 ( .A1(n18753), .A2(n18461), .B1(n18755), .B2(n18482), .ZN(
        n18450) );
  AOI22_X1 U21572 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n18462), .B1(
        n18754), .B2(n18742), .ZN(n18449) );
  OAI211_X1 U21573 ( .C1(n18465), .C2(n18758), .A(n18450), .B(n18449), .ZN(
        P3_U2885) );
  AOI22_X1 U21574 ( .A1(n18760), .A2(n18742), .B1(n18759), .B2(n18461), .ZN(
        n18452) );
  AOI22_X1 U21575 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n18462), .B1(
        n18761), .B2(n18482), .ZN(n18451) );
  OAI211_X1 U21576 ( .C1(n18465), .C2(n18764), .A(n18452), .B(n18451), .ZN(
        P3_U2886) );
  AOI22_X1 U21577 ( .A1(n18765), .A2(n18461), .B1(n18767), .B2(n18742), .ZN(
        n18454) );
  AOI22_X1 U21578 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n18462), .B1(
        n18766), .B2(n18482), .ZN(n18453) );
  OAI211_X1 U21579 ( .C1(n18465), .C2(n18770), .A(n18454), .B(n18453), .ZN(
        P3_U2887) );
  AOI22_X1 U21580 ( .A1(n18773), .A2(n18482), .B1(n18771), .B2(n18461), .ZN(
        n18456) );
  AOI22_X1 U21581 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n18462), .B1(
        n18772), .B2(n18742), .ZN(n18455) );
  OAI211_X1 U21582 ( .C1(n18465), .C2(n18776), .A(n18456), .B(n18455), .ZN(
        P3_U2888) );
  AOI22_X1 U21583 ( .A1(n18779), .A2(n18742), .B1(n18777), .B2(n18461), .ZN(
        n18458) );
  AOI22_X1 U21584 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n18462), .B1(
        n18778), .B2(n18482), .ZN(n18457) );
  OAI211_X1 U21585 ( .C1(n18465), .C2(n18782), .A(n18458), .B(n18457), .ZN(
        P3_U2889) );
  AOI22_X1 U21586 ( .A1(n18785), .A2(n18482), .B1(n18784), .B2(n18461), .ZN(
        n18460) );
  AOI22_X1 U21587 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n18462), .B1(
        n18783), .B2(n18742), .ZN(n18459) );
  OAI211_X1 U21588 ( .C1(n18465), .C2(n18788), .A(n18460), .B(n18459), .ZN(
        P3_U2890) );
  AOI22_X1 U21589 ( .A1(n18792), .A2(n18742), .B1(n18790), .B2(n18461), .ZN(
        n18464) );
  AOI22_X1 U21590 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n18462), .B1(
        n18794), .B2(n18482), .ZN(n18463) );
  OAI211_X1 U21591 ( .C1(n18465), .C2(n18799), .A(n18464), .B(n18463), .ZN(
        P3_U2891) );
  NAND2_X1 U21592 ( .A1(n18825), .A2(n18466), .ZN(n18509) );
  AND2_X1 U21593 ( .A1(n18868), .A2(n18511), .ZN(n18481) );
  AOI22_X1 U21594 ( .A1(n18503), .A2(n18749), .B1(n18743), .B2(n18481), .ZN(
        n18468) );
  AOI21_X1 U21595 ( .B1(n18620), .B2(n18717), .A(n18646), .ZN(n18555) );
  NAND2_X1 U21596 ( .A1(n18466), .A2(n18555), .ZN(n18483) );
  AOI22_X1 U21597 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n18483), .B1(
        n18744), .B2(n18482), .ZN(n18467) );
  OAI211_X1 U21598 ( .C1(n18509), .C2(n18752), .A(n18468), .B(n18467), .ZN(
        P3_U2892) );
  AOI22_X1 U21599 ( .A1(n18754), .A2(n18482), .B1(n18753), .B2(n18481), .ZN(
        n18470) );
  AOI22_X1 U21600 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n18483), .B1(
        n18503), .B2(n18755), .ZN(n18469) );
  OAI211_X1 U21601 ( .C1(n18509), .C2(n18758), .A(n18470), .B(n18469), .ZN(
        P3_U2893) );
  AOI22_X1 U21602 ( .A1(n18760), .A2(n18482), .B1(n18759), .B2(n18481), .ZN(
        n18472) );
  AOI22_X1 U21603 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n18483), .B1(
        n18503), .B2(n18761), .ZN(n18471) );
  OAI211_X1 U21604 ( .C1(n18509), .C2(n18764), .A(n18472), .B(n18471), .ZN(
        P3_U2894) );
  AOI22_X1 U21605 ( .A1(n18503), .A2(n18766), .B1(n18765), .B2(n18481), .ZN(
        n18474) );
  AOI22_X1 U21606 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n18483), .B1(
        n18767), .B2(n18482), .ZN(n18473) );
  OAI211_X1 U21607 ( .C1(n18509), .C2(n18770), .A(n18474), .B(n18473), .ZN(
        P3_U2895) );
  AOI22_X1 U21608 ( .A1(n18772), .A2(n18482), .B1(n18771), .B2(n18481), .ZN(
        n18476) );
  AOI22_X1 U21609 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n18483), .B1(
        n18503), .B2(n18773), .ZN(n18475) );
  OAI211_X1 U21610 ( .C1(n18509), .C2(n18776), .A(n18476), .B(n18475), .ZN(
        P3_U2896) );
  AOI22_X1 U21611 ( .A1(n18779), .A2(n18482), .B1(n18777), .B2(n18481), .ZN(
        n18478) );
  AOI22_X1 U21612 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n18483), .B1(
        n18503), .B2(n18778), .ZN(n18477) );
  OAI211_X1 U21613 ( .C1(n18509), .C2(n18782), .A(n18478), .B(n18477), .ZN(
        P3_U2897) );
  AOI22_X1 U21614 ( .A1(n18503), .A2(n18785), .B1(n18784), .B2(n18481), .ZN(
        n18480) );
  AOI22_X1 U21615 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n18483), .B1(
        n18783), .B2(n18482), .ZN(n18479) );
  OAI211_X1 U21616 ( .C1(n18509), .C2(n18788), .A(n18480), .B(n18479), .ZN(
        P3_U2898) );
  AOI22_X1 U21617 ( .A1(n18503), .A2(n18794), .B1(n18790), .B2(n18481), .ZN(
        n18485) );
  AOI22_X1 U21618 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n18483), .B1(
        n18792), .B2(n18482), .ZN(n18484) );
  OAI211_X1 U21619 ( .C1(n18509), .C2(n18799), .A(n18485), .B(n18484), .ZN(
        P3_U2899) );
  NAND2_X1 U21620 ( .A1(n18826), .A2(n18556), .ZN(n18507) );
  AOI21_X1 U21621 ( .B1(n18507), .B2(n18509), .A(n18715), .ZN(n18502) );
  AOI22_X1 U21622 ( .A1(n18503), .A2(n18744), .B1(n18743), .B2(n18502), .ZN(
        n18489) );
  AOI221_X1 U21623 ( .B1(n18486), .B2(n18509), .C1(n18717), .C2(n18509), .A(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n18487) );
  OAI21_X1 U21624 ( .B1(n18572), .B2(n18487), .A(n18720), .ZN(n18504) );
  AOI22_X1 U21625 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n18504), .B1(
        n18527), .B2(n18749), .ZN(n18488) );
  OAI211_X1 U21626 ( .C1(n18507), .C2(n18752), .A(n18489), .B(n18488), .ZN(
        P3_U2900) );
  AOI22_X1 U21627 ( .A1(n18527), .A2(n18755), .B1(n18502), .B2(n18753), .ZN(
        n18491) );
  AOI22_X1 U21628 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n18504), .B1(
        n18503), .B2(n18754), .ZN(n18490) );
  OAI211_X1 U21629 ( .C1(n18507), .C2(n18758), .A(n18491), .B(n18490), .ZN(
        P3_U2901) );
  AOI22_X1 U21630 ( .A1(n18527), .A2(n18761), .B1(n18502), .B2(n18759), .ZN(
        n18493) );
  AOI22_X1 U21631 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n18504), .B1(
        n18503), .B2(n18760), .ZN(n18492) );
  OAI211_X1 U21632 ( .C1(n18507), .C2(n18764), .A(n18493), .B(n18492), .ZN(
        P3_U2902) );
  AOI22_X1 U21633 ( .A1(n18503), .A2(n18767), .B1(n18502), .B2(n18765), .ZN(
        n18495) );
  AOI22_X1 U21634 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n18504), .B1(
        n18527), .B2(n18766), .ZN(n18494) );
  OAI211_X1 U21635 ( .C1(n18507), .C2(n18770), .A(n18495), .B(n18494), .ZN(
        P3_U2903) );
  AOI22_X1 U21636 ( .A1(n18527), .A2(n18773), .B1(n18502), .B2(n18771), .ZN(
        n18497) );
  AOI22_X1 U21637 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n18504), .B1(
        n18503), .B2(n18772), .ZN(n18496) );
  OAI211_X1 U21638 ( .C1(n18507), .C2(n18776), .A(n18497), .B(n18496), .ZN(
        P3_U2904) );
  AOI22_X1 U21639 ( .A1(n18503), .A2(n18779), .B1(n18502), .B2(n18777), .ZN(
        n18499) );
  AOI22_X1 U21640 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n18504), .B1(
        n18527), .B2(n18778), .ZN(n18498) );
  OAI211_X1 U21641 ( .C1(n18507), .C2(n18782), .A(n18499), .B(n18498), .ZN(
        P3_U2905) );
  AOI22_X1 U21642 ( .A1(n18503), .A2(n18783), .B1(n18502), .B2(n18784), .ZN(
        n18501) );
  AOI22_X1 U21643 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n18504), .B1(
        n18527), .B2(n18785), .ZN(n18500) );
  OAI211_X1 U21644 ( .C1(n18507), .C2(n18788), .A(n18501), .B(n18500), .ZN(
        P3_U2906) );
  AOI22_X1 U21645 ( .A1(n18527), .A2(n18794), .B1(n18502), .B2(n18790), .ZN(
        n18506) );
  AOI22_X1 U21646 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n18504), .B1(
        n18503), .B2(n18792), .ZN(n18505) );
  OAI211_X1 U21647 ( .C1(n18507), .C2(n18799), .A(n18506), .B(n18505), .ZN(
        P3_U2907) );
  INV_X1 U21648 ( .A(n18508), .ZN(n18599) );
  NAND2_X1 U21649 ( .A1(n18556), .A2(n18599), .ZN(n18532) );
  INV_X1 U21650 ( .A(n18556), .ZN(n18510) );
  NOR2_X1 U21651 ( .A1(n18510), .A2(n18690), .ZN(n18526) );
  AOI22_X1 U21652 ( .A1(n18550), .A2(n18749), .B1(n18743), .B2(n18526), .ZN(
        n18513) );
  AOI22_X1 U21653 ( .A1(n18748), .A2(n18511), .B1(n18556), .B2(n18692), .ZN(
        n18528) );
  AOI22_X1 U21654 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n18528), .B1(
        n18527), .B2(n18744), .ZN(n18512) );
  OAI211_X1 U21655 ( .C1(n18752), .C2(n18532), .A(n18513), .B(n18512), .ZN(
        P3_U2908) );
  AOI22_X1 U21656 ( .A1(n18527), .A2(n18754), .B1(n18753), .B2(n18526), .ZN(
        n18515) );
  AOI22_X1 U21657 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n18528), .B1(
        n18550), .B2(n18755), .ZN(n18514) );
  OAI211_X1 U21658 ( .C1(n18758), .C2(n18532), .A(n18515), .B(n18514), .ZN(
        P3_U2909) );
  AOI22_X1 U21659 ( .A1(n18527), .A2(n18760), .B1(n18759), .B2(n18526), .ZN(
        n18517) );
  AOI22_X1 U21660 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n18528), .B1(
        n18550), .B2(n18761), .ZN(n18516) );
  OAI211_X1 U21661 ( .C1(n18764), .C2(n18532), .A(n18517), .B(n18516), .ZN(
        P3_U2910) );
  AOI22_X1 U21662 ( .A1(n18527), .A2(n18767), .B1(n18765), .B2(n18526), .ZN(
        n18519) );
  AOI22_X1 U21663 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n18528), .B1(
        n18550), .B2(n18766), .ZN(n18518) );
  OAI211_X1 U21664 ( .C1(n18770), .C2(n18532), .A(n18519), .B(n18518), .ZN(
        P3_U2911) );
  AOI22_X1 U21665 ( .A1(n18527), .A2(n18772), .B1(n18771), .B2(n18526), .ZN(
        n18521) );
  AOI22_X1 U21666 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n18528), .B1(
        n18550), .B2(n18773), .ZN(n18520) );
  OAI211_X1 U21667 ( .C1(n18776), .C2(n18532), .A(n18521), .B(n18520), .ZN(
        P3_U2912) );
  AOI22_X1 U21668 ( .A1(n18550), .A2(n18778), .B1(n18777), .B2(n18526), .ZN(
        n18523) );
  AOI22_X1 U21669 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n18528), .B1(
        n18527), .B2(n18779), .ZN(n18522) );
  OAI211_X1 U21670 ( .C1(n18782), .C2(n18532), .A(n18523), .B(n18522), .ZN(
        P3_U2913) );
  AOI22_X1 U21671 ( .A1(n18550), .A2(n18785), .B1(n18784), .B2(n18526), .ZN(
        n18525) );
  AOI22_X1 U21672 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n18528), .B1(
        n18527), .B2(n18783), .ZN(n18524) );
  OAI211_X1 U21673 ( .C1(n18788), .C2(n18532), .A(n18525), .B(n18524), .ZN(
        P3_U2914) );
  AOI22_X1 U21674 ( .A1(n18550), .A2(n18794), .B1(n18790), .B2(n18526), .ZN(
        n18530) );
  AOI22_X1 U21675 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n18528), .B1(
        n18527), .B2(n18792), .ZN(n18529) );
  OAI211_X1 U21676 ( .C1(n18799), .C2(n18532), .A(n18530), .B(n18529), .ZN(
        P3_U2915) );
  NOR2_X1 U21677 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18531), .ZN(
        n18600) );
  NAND2_X1 U21678 ( .A1(n18600), .A2(n18621), .ZN(n18554) );
  NOR2_X1 U21679 ( .A1(n18594), .A2(n18615), .ZN(n18577) );
  NOR2_X1 U21680 ( .A1(n18715), .A2(n18577), .ZN(n18549) );
  AOI22_X1 U21681 ( .A1(n18550), .A2(n18744), .B1(n18743), .B2(n18549), .ZN(
        n18536) );
  NOR2_X1 U21682 ( .A1(n18572), .A2(n18550), .ZN(n18533) );
  OAI21_X1 U21683 ( .B1(n18533), .B2(n18717), .A(n18577), .ZN(n18534) );
  OAI211_X1 U21684 ( .C1(n18615), .C2(n18967), .A(n18720), .B(n18534), .ZN(
        n18551) );
  AOI22_X1 U21685 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n18551), .B1(
        n18572), .B2(n18749), .ZN(n18535) );
  OAI211_X1 U21686 ( .C1(n18752), .C2(n18554), .A(n18536), .B(n18535), .ZN(
        P3_U2916) );
  AOI22_X1 U21687 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n18551), .B1(
        n18753), .B2(n18549), .ZN(n18538) );
  AOI22_X1 U21688 ( .A1(n18572), .A2(n18755), .B1(n18550), .B2(n18754), .ZN(
        n18537) );
  OAI211_X1 U21689 ( .C1(n18758), .C2(n18554), .A(n18538), .B(n18537), .ZN(
        P3_U2917) );
  AOI22_X1 U21690 ( .A1(n18550), .A2(n18760), .B1(n18759), .B2(n18549), .ZN(
        n18540) );
  AOI22_X1 U21691 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n18551), .B1(
        n18572), .B2(n18761), .ZN(n18539) );
  OAI211_X1 U21692 ( .C1(n18764), .C2(n18554), .A(n18540), .B(n18539), .ZN(
        P3_U2918) );
  AOI22_X1 U21693 ( .A1(n18572), .A2(n18766), .B1(n18765), .B2(n18549), .ZN(
        n18542) );
  AOI22_X1 U21694 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n18551), .B1(
        n18550), .B2(n18767), .ZN(n18541) );
  OAI211_X1 U21695 ( .C1(n18770), .C2(n18554), .A(n18542), .B(n18541), .ZN(
        P3_U2919) );
  AOI22_X1 U21696 ( .A1(n18550), .A2(n18772), .B1(n18771), .B2(n18549), .ZN(
        n18544) );
  AOI22_X1 U21697 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n18551), .B1(
        n18572), .B2(n18773), .ZN(n18543) );
  OAI211_X1 U21698 ( .C1(n18776), .C2(n18554), .A(n18544), .B(n18543), .ZN(
        P3_U2920) );
  AOI22_X1 U21699 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n18551), .B1(
        n18777), .B2(n18549), .ZN(n18546) );
  AOI22_X1 U21700 ( .A1(n18572), .A2(n18778), .B1(n18550), .B2(n18779), .ZN(
        n18545) );
  OAI211_X1 U21701 ( .C1(n18782), .C2(n18554), .A(n18546), .B(n18545), .ZN(
        P3_U2921) );
  AOI22_X1 U21702 ( .A1(n18550), .A2(n18783), .B1(n18784), .B2(n18549), .ZN(
        n18548) );
  AOI22_X1 U21703 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n18551), .B1(
        n18572), .B2(n18785), .ZN(n18547) );
  OAI211_X1 U21704 ( .C1(n18788), .C2(n18554), .A(n18548), .B(n18547), .ZN(
        P3_U2922) );
  AOI22_X1 U21705 ( .A1(n18572), .A2(n18794), .B1(n18790), .B2(n18549), .ZN(
        n18553) );
  AOI22_X1 U21706 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n18551), .B1(
        n18550), .B2(n18792), .ZN(n18552) );
  OAI211_X1 U21707 ( .C1(n18799), .C2(n18554), .A(n18553), .B(n18552), .ZN(
        P3_U2923) );
  NAND2_X1 U21708 ( .A1(n18825), .A2(n18556), .ZN(n18576) );
  AND2_X1 U21709 ( .A1(n18868), .A2(n18600), .ZN(n18571) );
  AOI22_X1 U21710 ( .A1(n18572), .A2(n18744), .B1(n18743), .B2(n18571), .ZN(
        n18558) );
  NAND2_X1 U21711 ( .A1(n18556), .A2(n18555), .ZN(n18573) );
  AOI22_X1 U21712 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n18573), .B1(
        n18749), .B2(n18594), .ZN(n18557) );
  OAI211_X1 U21713 ( .C1(n18752), .C2(n18576), .A(n18558), .B(n18557), .ZN(
        P3_U2924) );
  AOI22_X1 U21714 ( .A1(n18753), .A2(n18571), .B1(n18755), .B2(n18594), .ZN(
        n18560) );
  AOI22_X1 U21715 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n18573), .B1(
        n18572), .B2(n18754), .ZN(n18559) );
  OAI211_X1 U21716 ( .C1(n18758), .C2(n18576), .A(n18560), .B(n18559), .ZN(
        P3_U2925) );
  AOI22_X1 U21717 ( .A1(n18761), .A2(n18594), .B1(n18759), .B2(n18571), .ZN(
        n18562) );
  AOI22_X1 U21718 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n18573), .B1(
        n18572), .B2(n18760), .ZN(n18561) );
  OAI211_X1 U21719 ( .C1(n18764), .C2(n18576), .A(n18562), .B(n18561), .ZN(
        P3_U2926) );
  AOI22_X1 U21720 ( .A1(n18572), .A2(n18767), .B1(n18765), .B2(n18571), .ZN(
        n18564) );
  AOI22_X1 U21721 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n18573), .B1(
        n18766), .B2(n18594), .ZN(n18563) );
  OAI211_X1 U21722 ( .C1(n18770), .C2(n18576), .A(n18564), .B(n18563), .ZN(
        P3_U2927) );
  AOI22_X1 U21723 ( .A1(n18773), .A2(n18594), .B1(n18771), .B2(n18571), .ZN(
        n18566) );
  AOI22_X1 U21724 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n18573), .B1(
        n18572), .B2(n18772), .ZN(n18565) );
  OAI211_X1 U21725 ( .C1(n18776), .C2(n18576), .A(n18566), .B(n18565), .ZN(
        P3_U2928) );
  AOI22_X1 U21726 ( .A1(n18572), .A2(n18779), .B1(n18777), .B2(n18571), .ZN(
        n18568) );
  AOI22_X1 U21727 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n18573), .B1(
        n18778), .B2(n18594), .ZN(n18567) );
  OAI211_X1 U21728 ( .C1(n18782), .C2(n18576), .A(n18568), .B(n18567), .ZN(
        P3_U2929) );
  AOI22_X1 U21729 ( .A1(n18785), .A2(n18594), .B1(n18784), .B2(n18571), .ZN(
        n18570) );
  AOI22_X1 U21730 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n18573), .B1(
        n18572), .B2(n18783), .ZN(n18569) );
  OAI211_X1 U21731 ( .C1(n18788), .C2(n18576), .A(n18570), .B(n18569), .ZN(
        P3_U2930) );
  AOI22_X1 U21732 ( .A1(n18572), .A2(n18792), .B1(n18790), .B2(n18571), .ZN(
        n18575) );
  AOI22_X1 U21733 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n18573), .B1(
        n18794), .B2(n18594), .ZN(n18574) );
  OAI211_X1 U21734 ( .C1(n18799), .C2(n18576), .A(n18575), .B(n18574), .ZN(
        P3_U2931) );
  NAND2_X1 U21735 ( .A1(n18826), .A2(n18645), .ZN(n18598) );
  INV_X1 U21736 ( .A(n18576), .ZN(n18640) );
  NOR2_X1 U21737 ( .A1(n18640), .A2(n18663), .ZN(n18623) );
  NOR2_X1 U21738 ( .A1(n18715), .A2(n18623), .ZN(n18593) );
  AOI22_X1 U21739 ( .A1(n18744), .A2(n18594), .B1(n18743), .B2(n18593), .ZN(
        n18580) );
  OAI21_X1 U21740 ( .B1(n18577), .B2(n18717), .A(n18623), .ZN(n18578) );
  OAI211_X1 U21741 ( .C1(n18663), .C2(n18967), .A(n18720), .B(n18578), .ZN(
        n18595) );
  AOI22_X1 U21742 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n18595), .B1(
        n18749), .B2(n18615), .ZN(n18579) );
  OAI211_X1 U21743 ( .C1(n18752), .C2(n18598), .A(n18580), .B(n18579), .ZN(
        P3_U2932) );
  AOI22_X1 U21744 ( .A1(n18754), .A2(n18594), .B1(n18753), .B2(n18593), .ZN(
        n18582) );
  AOI22_X1 U21745 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n18595), .B1(
        n18755), .B2(n18615), .ZN(n18581) );
  OAI211_X1 U21746 ( .C1(n18758), .C2(n18598), .A(n18582), .B(n18581), .ZN(
        P3_U2933) );
  AOI22_X1 U21747 ( .A1(n18761), .A2(n18615), .B1(n18759), .B2(n18593), .ZN(
        n18584) );
  AOI22_X1 U21748 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n18595), .B1(
        n18760), .B2(n18594), .ZN(n18583) );
  OAI211_X1 U21749 ( .C1(n18764), .C2(n18598), .A(n18584), .B(n18583), .ZN(
        P3_U2934) );
  AOI22_X1 U21750 ( .A1(n18766), .A2(n18615), .B1(n18765), .B2(n18593), .ZN(
        n18586) );
  AOI22_X1 U21751 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n18595), .B1(
        n18767), .B2(n18594), .ZN(n18585) );
  OAI211_X1 U21752 ( .C1(n18770), .C2(n18598), .A(n18586), .B(n18585), .ZN(
        P3_U2935) );
  AOI22_X1 U21753 ( .A1(n18773), .A2(n18615), .B1(n18771), .B2(n18593), .ZN(
        n18588) );
  AOI22_X1 U21754 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n18595), .B1(
        n18772), .B2(n18594), .ZN(n18587) );
  OAI211_X1 U21755 ( .C1(n18776), .C2(n18598), .A(n18588), .B(n18587), .ZN(
        P3_U2936) );
  AOI22_X1 U21756 ( .A1(n18778), .A2(n18615), .B1(n18777), .B2(n18593), .ZN(
        n18590) );
  AOI22_X1 U21757 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n18595), .B1(
        n18779), .B2(n18594), .ZN(n18589) );
  OAI211_X1 U21758 ( .C1(n18782), .C2(n18598), .A(n18590), .B(n18589), .ZN(
        P3_U2937) );
  AOI22_X1 U21759 ( .A1(n18785), .A2(n18615), .B1(n18784), .B2(n18593), .ZN(
        n18592) );
  AOI22_X1 U21760 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n18595), .B1(
        n18783), .B2(n18594), .ZN(n18591) );
  OAI211_X1 U21761 ( .C1(n18788), .C2(n18598), .A(n18592), .B(n18591), .ZN(
        P3_U2938) );
  AOI22_X1 U21762 ( .A1(n18790), .A2(n18593), .B1(n18794), .B2(n18615), .ZN(
        n18597) );
  AOI22_X1 U21763 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n18595), .B1(
        n18792), .B2(n18594), .ZN(n18596) );
  OAI211_X1 U21764 ( .C1(n18799), .C2(n18598), .A(n18597), .B(n18596), .ZN(
        P3_U2939) );
  NAND2_X1 U21765 ( .A1(n18599), .A2(n18645), .ZN(n18622) );
  INV_X1 U21766 ( .A(n18645), .ZN(n18619) );
  NOR2_X1 U21767 ( .A1(n18619), .A2(n18690), .ZN(n18647) );
  AOI22_X1 U21768 ( .A1(n18749), .A2(n18640), .B1(n18743), .B2(n18647), .ZN(
        n18602) );
  AOI22_X1 U21769 ( .A1(n18748), .A2(n18600), .B1(n18645), .B2(n18692), .ZN(
        n18616) );
  AOI22_X1 U21770 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n18616), .B1(
        n18744), .B2(n18615), .ZN(n18601) );
  OAI211_X1 U21771 ( .C1(n18752), .C2(n18622), .A(n18602), .B(n18601), .ZN(
        P3_U2940) );
  AOI22_X1 U21772 ( .A1(n18753), .A2(n18647), .B1(n18755), .B2(n18640), .ZN(
        n18604) );
  AOI22_X1 U21773 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n18616), .B1(
        n18754), .B2(n18615), .ZN(n18603) );
  OAI211_X1 U21774 ( .C1(n18758), .C2(n18622), .A(n18604), .B(n18603), .ZN(
        P3_U2941) );
  AOI22_X1 U21775 ( .A1(n18760), .A2(n18615), .B1(n18759), .B2(n18647), .ZN(
        n18606) );
  AOI22_X1 U21776 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n18616), .B1(
        n18761), .B2(n18640), .ZN(n18605) );
  OAI211_X1 U21777 ( .C1(n18764), .C2(n18622), .A(n18606), .B(n18605), .ZN(
        P3_U2942) );
  AOI22_X1 U21778 ( .A1(n18765), .A2(n18647), .B1(n18767), .B2(n18615), .ZN(
        n18608) );
  AOI22_X1 U21779 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n18616), .B1(
        n18766), .B2(n18640), .ZN(n18607) );
  OAI211_X1 U21780 ( .C1(n18770), .C2(n18622), .A(n18608), .B(n18607), .ZN(
        P3_U2943) );
  AOI22_X1 U21781 ( .A1(n18772), .A2(n18615), .B1(n18771), .B2(n18647), .ZN(
        n18610) );
  AOI22_X1 U21782 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n18616), .B1(
        n18773), .B2(n18640), .ZN(n18609) );
  OAI211_X1 U21783 ( .C1(n18776), .C2(n18622), .A(n18610), .B(n18609), .ZN(
        P3_U2944) );
  AOI22_X1 U21784 ( .A1(n18779), .A2(n18615), .B1(n18777), .B2(n18647), .ZN(
        n18612) );
  AOI22_X1 U21785 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n18616), .B1(
        n18778), .B2(n18640), .ZN(n18611) );
  OAI211_X1 U21786 ( .C1(n18782), .C2(n18622), .A(n18612), .B(n18611), .ZN(
        P3_U2945) );
  AOI22_X1 U21787 ( .A1(n18784), .A2(n18647), .B1(n18783), .B2(n18615), .ZN(
        n18614) );
  AOI22_X1 U21788 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n18616), .B1(
        n18785), .B2(n18640), .ZN(n18613) );
  OAI211_X1 U21789 ( .C1(n18788), .C2(n18622), .A(n18614), .B(n18613), .ZN(
        P3_U2946) );
  AOI22_X1 U21790 ( .A1(n18790), .A2(n18647), .B1(n18794), .B2(n18640), .ZN(
        n18618) );
  AOI22_X1 U21791 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n18616), .B1(
        n18792), .B2(n18615), .ZN(n18617) );
  OAI211_X1 U21792 ( .C1(n18799), .C2(n18622), .A(n18618), .B(n18617), .ZN(
        P3_U2947) );
  NOR2_X1 U21793 ( .A1(n18620), .A2(n18619), .ZN(n18694) );
  NAND2_X1 U21794 ( .A1(n18694), .A2(n18621), .ZN(n18644) );
  NOR2_X1 U21795 ( .A1(n18685), .A2(n18709), .ZN(n18668) );
  NOR2_X1 U21796 ( .A1(n18715), .A2(n18668), .ZN(n18639) );
  AOI22_X1 U21797 ( .A1(n18744), .A2(n18640), .B1(n18743), .B2(n18639), .ZN(
        n18626) );
  OAI21_X1 U21798 ( .B1(n18623), .B2(n18717), .A(n18668), .ZN(n18624) );
  OAI211_X1 U21799 ( .C1(n18709), .C2(n18967), .A(n18720), .B(n18624), .ZN(
        n18641) );
  AOI22_X1 U21800 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n18641), .B1(
        n18749), .B2(n18663), .ZN(n18625) );
  OAI211_X1 U21801 ( .C1(n18752), .C2(n18644), .A(n18626), .B(n18625), .ZN(
        P3_U2948) );
  AOI22_X1 U21802 ( .A1(n18754), .A2(n18640), .B1(n18753), .B2(n18639), .ZN(
        n18628) );
  AOI22_X1 U21803 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n18641), .B1(
        n18755), .B2(n18663), .ZN(n18627) );
  OAI211_X1 U21804 ( .C1(n18758), .C2(n18644), .A(n18628), .B(n18627), .ZN(
        P3_U2949) );
  AOI22_X1 U21805 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n18641), .B1(
        n18759), .B2(n18639), .ZN(n18630) );
  AOI22_X1 U21806 ( .A1(n18760), .A2(n18640), .B1(n18761), .B2(n18663), .ZN(
        n18629) );
  OAI211_X1 U21807 ( .C1(n18764), .C2(n18644), .A(n18630), .B(n18629), .ZN(
        P3_U2950) );
  AOI22_X1 U21808 ( .A1(n18765), .A2(n18639), .B1(n18767), .B2(n18640), .ZN(
        n18632) );
  AOI22_X1 U21809 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n18641), .B1(
        n18766), .B2(n18663), .ZN(n18631) );
  OAI211_X1 U21810 ( .C1(n18770), .C2(n18644), .A(n18632), .B(n18631), .ZN(
        P3_U2951) );
  AOI22_X1 U21811 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n18641), .B1(
        n18771), .B2(n18639), .ZN(n18634) );
  AOI22_X1 U21812 ( .A1(n18772), .A2(n18640), .B1(n18773), .B2(n18663), .ZN(
        n18633) );
  OAI211_X1 U21813 ( .C1(n18776), .C2(n18644), .A(n18634), .B(n18633), .ZN(
        P3_U2952) );
  AOI22_X1 U21814 ( .A1(n18778), .A2(n18663), .B1(n18777), .B2(n18639), .ZN(
        n18636) );
  AOI22_X1 U21815 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n18641), .B1(
        n18779), .B2(n18640), .ZN(n18635) );
  OAI211_X1 U21816 ( .C1(n18782), .C2(n18644), .A(n18636), .B(n18635), .ZN(
        P3_U2953) );
  AOI22_X1 U21817 ( .A1(n18785), .A2(n18663), .B1(n18784), .B2(n18639), .ZN(
        n18638) );
  AOI22_X1 U21818 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n18641), .B1(
        n18783), .B2(n18640), .ZN(n18637) );
  OAI211_X1 U21819 ( .C1(n18788), .C2(n18644), .A(n18638), .B(n18637), .ZN(
        P3_U2954) );
  AOI22_X1 U21820 ( .A1(n18790), .A2(n18639), .B1(n18794), .B2(n18663), .ZN(
        n18643) );
  AOI22_X1 U21821 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n18641), .B1(
        n18792), .B2(n18640), .ZN(n18642) );
  OAI211_X1 U21822 ( .C1(n18799), .C2(n18644), .A(n18643), .B(n18642), .ZN(
        P3_U2955) );
  NAND2_X1 U21823 ( .A1(n18825), .A2(n18645), .ZN(n18667) );
  AND2_X1 U21824 ( .A1(n18868), .A2(n18694), .ZN(n18662) );
  AOI22_X1 U21825 ( .A1(n18744), .A2(n18663), .B1(n18743), .B2(n18662), .ZN(
        n18649) );
  INV_X1 U21826 ( .A(n18646), .ZN(n18745) );
  AOI22_X1 U21827 ( .A1(n18748), .A2(n18647), .B1(n18745), .B2(n18694), .ZN(
        n18664) );
  AOI22_X1 U21828 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n18664), .B1(
        n18749), .B2(n18685), .ZN(n18648) );
  OAI211_X1 U21829 ( .C1(n18752), .C2(n18667), .A(n18649), .B(n18648), .ZN(
        P3_U2956) );
  AOI22_X1 U21830 ( .A1(n18754), .A2(n18663), .B1(n18753), .B2(n18662), .ZN(
        n18651) );
  AOI22_X1 U21831 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n18664), .B1(
        n18755), .B2(n18685), .ZN(n18650) );
  OAI211_X1 U21832 ( .C1(n18758), .C2(n18667), .A(n18651), .B(n18650), .ZN(
        P3_U2957) );
  AOI22_X1 U21833 ( .A1(n18760), .A2(n18663), .B1(n18759), .B2(n18662), .ZN(
        n18653) );
  AOI22_X1 U21834 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n18664), .B1(
        n18761), .B2(n18685), .ZN(n18652) );
  OAI211_X1 U21835 ( .C1(n18764), .C2(n18667), .A(n18653), .B(n18652), .ZN(
        P3_U2958) );
  AOI22_X1 U21836 ( .A1(n18765), .A2(n18662), .B1(n18767), .B2(n18663), .ZN(
        n18655) );
  AOI22_X1 U21837 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n18664), .B1(
        n18766), .B2(n18685), .ZN(n18654) );
  OAI211_X1 U21838 ( .C1(n18770), .C2(n18667), .A(n18655), .B(n18654), .ZN(
        P3_U2959) );
  AOI22_X1 U21839 ( .A1(n18772), .A2(n18663), .B1(n18771), .B2(n18662), .ZN(
        n18657) );
  AOI22_X1 U21840 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n18664), .B1(
        n18773), .B2(n18685), .ZN(n18656) );
  OAI211_X1 U21841 ( .C1(n18776), .C2(n18667), .A(n18657), .B(n18656), .ZN(
        P3_U2960) );
  AOI22_X1 U21842 ( .A1(n18779), .A2(n18663), .B1(n18777), .B2(n18662), .ZN(
        n18659) );
  AOI22_X1 U21843 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n18664), .B1(
        n18778), .B2(n18685), .ZN(n18658) );
  OAI211_X1 U21844 ( .C1(n18782), .C2(n18667), .A(n18659), .B(n18658), .ZN(
        P3_U2961) );
  AOI22_X1 U21845 ( .A1(n18784), .A2(n18662), .B1(n18783), .B2(n18663), .ZN(
        n18661) );
  AOI22_X1 U21846 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n18664), .B1(
        n18785), .B2(n18685), .ZN(n18660) );
  OAI211_X1 U21847 ( .C1(n18788), .C2(n18667), .A(n18661), .B(n18660), .ZN(
        P3_U2962) );
  AOI22_X1 U21848 ( .A1(n18790), .A2(n18662), .B1(n18794), .B2(n18685), .ZN(
        n18666) );
  AOI22_X1 U21849 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n18664), .B1(
        n18792), .B2(n18663), .ZN(n18665) );
  OAI211_X1 U21850 ( .C1(n18799), .C2(n18667), .A(n18666), .B(n18665), .ZN(
        P3_U2963) );
  INV_X1 U21851 ( .A(n18691), .ZN(n18693) );
  NAND2_X1 U21852 ( .A1(n18826), .A2(n18693), .ZN(n18689) );
  INV_X1 U21853 ( .A(n18689), .ZN(n18791) );
  NOR2_X1 U21854 ( .A1(n18737), .A2(n18791), .ZN(n18718) );
  NOR2_X1 U21855 ( .A1(n18715), .A2(n18718), .ZN(n18684) );
  AOI22_X1 U21856 ( .A1(n18749), .A2(n18709), .B1(n18743), .B2(n18684), .ZN(
        n18671) );
  OAI21_X1 U21857 ( .B1(n18668), .B2(n18717), .A(n18718), .ZN(n18669) );
  OAI211_X1 U21858 ( .C1(n18791), .C2(n18967), .A(n18720), .B(n18669), .ZN(
        n18686) );
  AOI22_X1 U21859 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n18686), .B1(
        n18744), .B2(n18685), .ZN(n18670) );
  OAI211_X1 U21860 ( .C1(n18752), .C2(n18689), .A(n18671), .B(n18670), .ZN(
        P3_U2964) );
  AOI22_X1 U21861 ( .A1(n18754), .A2(n18685), .B1(n18753), .B2(n18684), .ZN(
        n18673) );
  AOI22_X1 U21862 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n18686), .B1(
        n18755), .B2(n18709), .ZN(n18672) );
  OAI211_X1 U21863 ( .C1(n18758), .C2(n18689), .A(n18673), .B(n18672), .ZN(
        P3_U2965) );
  AOI22_X1 U21864 ( .A1(n18760), .A2(n18685), .B1(n18759), .B2(n18684), .ZN(
        n18675) );
  AOI22_X1 U21865 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n18686), .B1(
        n18761), .B2(n18709), .ZN(n18674) );
  OAI211_X1 U21866 ( .C1(n18764), .C2(n18689), .A(n18675), .B(n18674), .ZN(
        P3_U2966) );
  AOI22_X1 U21867 ( .A1(n18766), .A2(n18709), .B1(n18765), .B2(n18684), .ZN(
        n18677) );
  AOI22_X1 U21868 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n18686), .B1(
        n18767), .B2(n18685), .ZN(n18676) );
  OAI211_X1 U21869 ( .C1(n18770), .C2(n18689), .A(n18677), .B(n18676), .ZN(
        P3_U2967) );
  AOI22_X1 U21870 ( .A1(n18773), .A2(n18709), .B1(n18771), .B2(n18684), .ZN(
        n18679) );
  AOI22_X1 U21871 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n18686), .B1(
        n18772), .B2(n18685), .ZN(n18678) );
  OAI211_X1 U21872 ( .C1(n18776), .C2(n18689), .A(n18679), .B(n18678), .ZN(
        P3_U2968) );
  AOI22_X1 U21873 ( .A1(n18778), .A2(n18709), .B1(n18777), .B2(n18684), .ZN(
        n18681) );
  AOI22_X1 U21874 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n18686), .B1(
        n18779), .B2(n18685), .ZN(n18680) );
  OAI211_X1 U21875 ( .C1(n18782), .C2(n18689), .A(n18681), .B(n18680), .ZN(
        P3_U2969) );
  AOI22_X1 U21876 ( .A1(n18784), .A2(n18684), .B1(n18783), .B2(n18685), .ZN(
        n18683) );
  AOI22_X1 U21877 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n18686), .B1(
        n18785), .B2(n18709), .ZN(n18682) );
  OAI211_X1 U21878 ( .C1(n18788), .C2(n18689), .A(n18683), .B(n18682), .ZN(
        P3_U2970) );
  AOI22_X1 U21879 ( .A1(n18792), .A2(n18685), .B1(n18790), .B2(n18684), .ZN(
        n18688) );
  AOI22_X1 U21880 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n18686), .B1(
        n18794), .B2(n18709), .ZN(n18687) );
  OAI211_X1 U21881 ( .C1(n18799), .C2(n18689), .A(n18688), .B(n18687), .ZN(
        P3_U2971) );
  NOR2_X1 U21882 ( .A1(n18691), .A2(n18690), .ZN(n18747) );
  AOI22_X1 U21883 ( .A1(n18744), .A2(n18709), .B1(n18743), .B2(n18747), .ZN(
        n18696) );
  AOI22_X1 U21884 ( .A1(n18748), .A2(n18694), .B1(n18693), .B2(n18692), .ZN(
        n18710) );
  AOI22_X1 U21885 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n18710), .B1(
        n18749), .B2(n18737), .ZN(n18695) );
  OAI211_X1 U21886 ( .C1(n18752), .C2(n18713), .A(n18696), .B(n18695), .ZN(
        P3_U2972) );
  AOI22_X1 U21887 ( .A1(n18753), .A2(n18747), .B1(n18755), .B2(n18737), .ZN(
        n18698) );
  AOI22_X1 U21888 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n18710), .B1(
        n18754), .B2(n18709), .ZN(n18697) );
  OAI211_X1 U21889 ( .C1(n18758), .C2(n18713), .A(n18698), .B(n18697), .ZN(
        P3_U2973) );
  AOI22_X1 U21890 ( .A1(n18761), .A2(n18737), .B1(n18759), .B2(n18747), .ZN(
        n18700) );
  AOI22_X1 U21891 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n18710), .B1(
        n18760), .B2(n18709), .ZN(n18699) );
  OAI211_X1 U21892 ( .C1(n18764), .C2(n18713), .A(n18700), .B(n18699), .ZN(
        P3_U2974) );
  AOI22_X1 U21893 ( .A1(n18765), .A2(n18747), .B1(n18767), .B2(n18709), .ZN(
        n18702) );
  AOI22_X1 U21894 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n18710), .B1(
        n18766), .B2(n18737), .ZN(n18701) );
  OAI211_X1 U21895 ( .C1(n18770), .C2(n18713), .A(n18702), .B(n18701), .ZN(
        P3_U2975) );
  AOI22_X1 U21896 ( .A1(n18772), .A2(n18709), .B1(n18771), .B2(n18747), .ZN(
        n18704) );
  AOI22_X1 U21897 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n18710), .B1(
        n18773), .B2(n18737), .ZN(n18703) );
  OAI211_X1 U21898 ( .C1(n18776), .C2(n18713), .A(n18704), .B(n18703), .ZN(
        P3_U2976) );
  AOI22_X1 U21899 ( .A1(n18778), .A2(n18737), .B1(n18777), .B2(n18747), .ZN(
        n18706) );
  AOI22_X1 U21900 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n18710), .B1(
        n18779), .B2(n18709), .ZN(n18705) );
  OAI211_X1 U21901 ( .C1(n18782), .C2(n18713), .A(n18706), .B(n18705), .ZN(
        P3_U2977) );
  AOI22_X1 U21902 ( .A1(n18784), .A2(n18747), .B1(n18783), .B2(n18709), .ZN(
        n18708) );
  AOI22_X1 U21903 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n18710), .B1(
        n18785), .B2(n18737), .ZN(n18707) );
  OAI211_X1 U21904 ( .C1(n18788), .C2(n18713), .A(n18708), .B(n18707), .ZN(
        P3_U2978) );
  AOI22_X1 U21905 ( .A1(n18792), .A2(n18709), .B1(n18790), .B2(n18747), .ZN(
        n18712) );
  AOI22_X1 U21906 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n18710), .B1(
        n18794), .B2(n18737), .ZN(n18711) );
  OAI211_X1 U21907 ( .C1(n18799), .C2(n18713), .A(n18712), .B(n18711), .ZN(
        P3_U2979) );
  INV_X1 U21908 ( .A(n18714), .ZN(n18716) );
  NOR2_X1 U21909 ( .A1(n18715), .A2(n18716), .ZN(n18736) );
  AOI22_X1 U21910 ( .A1(n18749), .A2(n18791), .B1(n18743), .B2(n18736), .ZN(
        n18723) );
  OAI21_X1 U21911 ( .B1(n18718), .B2(n18717), .A(n18716), .ZN(n18719) );
  OAI211_X1 U21912 ( .C1(n18721), .C2(n18967), .A(n18720), .B(n18719), .ZN(
        n18738) );
  AOI22_X1 U21913 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n18738), .B1(
        n18744), .B2(n18737), .ZN(n18722) );
  OAI211_X1 U21914 ( .C1(n18752), .C2(n18741), .A(n18723), .B(n18722), .ZN(
        P3_U2980) );
  AOI22_X1 U21915 ( .A1(n18753), .A2(n18736), .B1(n18755), .B2(n18791), .ZN(
        n18725) );
  AOI22_X1 U21916 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n18738), .B1(
        n18754), .B2(n18737), .ZN(n18724) );
  OAI211_X1 U21917 ( .C1(n18758), .C2(n18741), .A(n18725), .B(n18724), .ZN(
        P3_U2981) );
  AOI22_X1 U21918 ( .A1(n18761), .A2(n18791), .B1(n18759), .B2(n18736), .ZN(
        n18727) );
  AOI22_X1 U21919 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n18738), .B1(
        n18760), .B2(n18737), .ZN(n18726) );
  OAI211_X1 U21920 ( .C1(n18764), .C2(n18741), .A(n18727), .B(n18726), .ZN(
        P3_U2982) );
  AOI22_X1 U21921 ( .A1(n18765), .A2(n18736), .B1(n18767), .B2(n18737), .ZN(
        n18729) );
  AOI22_X1 U21922 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n18738), .B1(
        n18766), .B2(n18791), .ZN(n18728) );
  OAI211_X1 U21923 ( .C1(n18770), .C2(n18741), .A(n18729), .B(n18728), .ZN(
        P3_U2983) );
  AOI22_X1 U21924 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n18738), .B1(
        n18771), .B2(n18736), .ZN(n18731) );
  AOI22_X1 U21925 ( .A1(n18772), .A2(n18737), .B1(n18773), .B2(n18791), .ZN(
        n18730) );
  OAI211_X1 U21926 ( .C1(n18776), .C2(n18741), .A(n18731), .B(n18730), .ZN(
        P3_U2984) );
  AOI22_X1 U21927 ( .A1(n18779), .A2(n18737), .B1(n18777), .B2(n18736), .ZN(
        n18733) );
  AOI22_X1 U21928 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n18738), .B1(
        n18778), .B2(n18791), .ZN(n18732) );
  OAI211_X1 U21929 ( .C1(n18782), .C2(n18741), .A(n18733), .B(n18732), .ZN(
        P3_U2985) );
  AOI22_X1 U21930 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n18738), .B1(
        n18784), .B2(n18736), .ZN(n18735) );
  AOI22_X1 U21931 ( .A1(n18785), .A2(n18791), .B1(n18783), .B2(n18737), .ZN(
        n18734) );
  OAI211_X1 U21932 ( .C1(n18788), .C2(n18741), .A(n18735), .B(n18734), .ZN(
        P3_U2986) );
  AOI22_X1 U21933 ( .A1(n18790), .A2(n18736), .B1(n18794), .B2(n18791), .ZN(
        n18740) );
  AOI22_X1 U21934 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n18738), .B1(
        n18792), .B2(n18737), .ZN(n18739) );
  OAI211_X1 U21935 ( .C1(n18799), .C2(n18741), .A(n18740), .B(n18739), .ZN(
        P3_U2987) );
  INV_X1 U21936 ( .A(n18742), .ZN(n18798) );
  AND2_X1 U21937 ( .A1(n18868), .A2(n18746), .ZN(n18789) );
  AOI22_X1 U21938 ( .A1(n18744), .A2(n18791), .B1(n18743), .B2(n18789), .ZN(
        n18751) );
  AOI22_X1 U21939 ( .A1(n18748), .A2(n18747), .B1(n18746), .B2(n18745), .ZN(
        n18795) );
  AOI22_X1 U21940 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n18795), .B1(
        n18749), .B2(n18793), .ZN(n18750) );
  OAI211_X1 U21941 ( .C1(n18752), .C2(n18798), .A(n18751), .B(n18750), .ZN(
        P3_U2988) );
  AOI22_X1 U21942 ( .A1(n18754), .A2(n18791), .B1(n18753), .B2(n18789), .ZN(
        n18757) );
  AOI22_X1 U21943 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n18795), .B1(
        n18755), .B2(n18793), .ZN(n18756) );
  OAI211_X1 U21944 ( .C1(n18758), .C2(n18798), .A(n18757), .B(n18756), .ZN(
        P3_U2989) );
  AOI22_X1 U21945 ( .A1(n18760), .A2(n18791), .B1(n18759), .B2(n18789), .ZN(
        n18763) );
  AOI22_X1 U21946 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n18795), .B1(
        n18761), .B2(n18793), .ZN(n18762) );
  OAI211_X1 U21947 ( .C1(n18764), .C2(n18798), .A(n18763), .B(n18762), .ZN(
        P3_U2990) );
  AOI22_X1 U21948 ( .A1(n18766), .A2(n18793), .B1(n18765), .B2(n18789), .ZN(
        n18769) );
  AOI22_X1 U21949 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n18795), .B1(
        n18767), .B2(n18791), .ZN(n18768) );
  OAI211_X1 U21950 ( .C1(n18770), .C2(n18798), .A(n18769), .B(n18768), .ZN(
        P3_U2991) );
  AOI22_X1 U21951 ( .A1(n18772), .A2(n18791), .B1(n18771), .B2(n18789), .ZN(
        n18775) );
  AOI22_X1 U21952 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n18795), .B1(
        n18773), .B2(n18793), .ZN(n18774) );
  OAI211_X1 U21953 ( .C1(n18776), .C2(n18798), .A(n18775), .B(n18774), .ZN(
        P3_U2992) );
  AOI22_X1 U21954 ( .A1(n18778), .A2(n18793), .B1(n18777), .B2(n18789), .ZN(
        n18781) );
  AOI22_X1 U21955 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n18795), .B1(
        n18779), .B2(n18791), .ZN(n18780) );
  OAI211_X1 U21956 ( .C1(n18782), .C2(n18798), .A(n18781), .B(n18780), .ZN(
        P3_U2993) );
  AOI22_X1 U21957 ( .A1(n18784), .A2(n18789), .B1(n18783), .B2(n18791), .ZN(
        n18787) );
  AOI22_X1 U21958 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n18795), .B1(
        n18785), .B2(n18793), .ZN(n18786) );
  OAI211_X1 U21959 ( .C1(n18788), .C2(n18798), .A(n18787), .B(n18786), .ZN(
        P3_U2994) );
  AOI22_X1 U21960 ( .A1(n18792), .A2(n18791), .B1(n18790), .B2(n18789), .ZN(
        n18797) );
  AOI22_X1 U21961 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n18795), .B1(
        n18794), .B2(n18793), .ZN(n18796) );
  OAI211_X1 U21962 ( .C1(n18799), .C2(n18798), .A(n18797), .B(n18796), .ZN(
        P3_U2995) );
  INV_X1 U21963 ( .A(n18800), .ZN(n18803) );
  AOI22_X1 U21964 ( .A1(n18804), .A2(n18803), .B1(n18802), .B2(n18801), .ZN(
        n18805) );
  OAI221_X1 U21965 ( .B1(n18808), .B2(n18807), .C1(n18808), .C2(n18806), .A(
        n18805), .ZN(n19010) );
  OAI21_X1 U21966 ( .B1(P3_MORE_REG_SCAN_IN), .B2(P3_FLUSH_REG_SCAN_IN), .A(
        n18809), .ZN(n18810) );
  OAI211_X1 U21967 ( .C1(n18812), .C2(n18842), .A(n18811), .B(n18810), .ZN(
        n18853) );
  AOI21_X1 U21968 ( .B1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n18813), .A(
        n18824), .ZN(n18822) );
  AOI211_X1 U21969 ( .C1(n18982), .C2(n12506), .A(n18822), .B(n18838), .ZN(
        n18819) );
  AOI21_X1 U21970 ( .B1(n18816), .B2(n18815), .A(n18814), .ZN(n18835) );
  NOR3_X1 U21971 ( .A1(n18817), .A2(n18835), .A3(n18982), .ZN(n18818) );
  AOI211_X1 U21972 ( .C1(n18831), .C2(n18978), .A(n18819), .B(n18818), .ZN(
        n18979) );
  MUX2_X1 U21973 ( .A(n18982), .B(n18979), .S(n18842), .Z(n18829) );
  NAND2_X1 U21974 ( .A1(n18821), .A2(n18820), .ZN(n18823) );
  INV_X1 U21975 ( .A(n18822), .ZN(n18832) );
  AOI22_X1 U21976 ( .A1(n18987), .A2(n18823), .B1(n12506), .B2(n18832), .ZN(
        n18983) );
  AOI222_X1 U21977 ( .A1(n18983), .A2(n18992), .B1(n18983), .B2(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .C1(n18992), .C2(n18825), .ZN(
        n18827) );
  AOI21_X1 U21978 ( .B1(n18827), .B2(n18842), .A(n18826), .ZN(n18828) );
  AOI21_X1 U21979 ( .B1(n18829), .B2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        n18828), .ZN(n18843) );
  INV_X1 U21980 ( .A(n18829), .ZN(n18844) );
  AOI221_X1 U21981 ( .B1(n18843), .B2(n18847), .C1(n18846), .C2(n18847), .A(
        n18844), .ZN(n18851) );
  AOI22_X1 U21982 ( .A1(n18838), .A2(n18832), .B1(n18831), .B2(n18830), .ZN(
        n18833) );
  NOR2_X1 U21983 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n18833), .ZN(
        n18969) );
  INV_X1 U21984 ( .A(n18834), .ZN(n18836) );
  OAI22_X1 U21985 ( .A1(n18838), .A2(n18837), .B1(n18836), .B2(n18835), .ZN(
        n18839) );
  AOI21_X1 U21986 ( .B1(n18982), .B2(n18840), .A(n18839), .ZN(n18970) );
  NAND2_X1 U21987 ( .A1(n18842), .A2(n18970), .ZN(n18841) );
  AOI22_X1 U21988 ( .A1(n18842), .A2(n18969), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n18841), .ZN(n18850) );
  AOI21_X1 U21989 ( .B1(n18845), .B2(n18844), .A(n18843), .ZN(n18849) );
  NAND2_X1 U21990 ( .A1(n18847), .A2(n18846), .ZN(n18848) );
  OAI22_X1 U21991 ( .A1(n18851), .A2(n18850), .B1(n18849), .B2(n18848), .ZN(
        n18852) );
  NOR4_X1 U21992 ( .A1(n18854), .A2(n19010), .A3(n18853), .A4(n18852), .ZN(
        n18865) );
  INV_X1 U21993 ( .A(n19016), .ZN(n18878) );
  AOI22_X1 U21994 ( .A1(n18988), .A2(n18878), .B1(n9998), .B2(n18866), .ZN(
        n18855) );
  INV_X1 U21995 ( .A(n18855), .ZN(n18861) );
  OAI211_X1 U21996 ( .C1(n18857), .C2(n18856), .A(n19020), .B(n18865), .ZN(
        n18966) );
  OAI21_X1 U21997 ( .B1(P3_STATE2_REG_2__SCAN_IN), .B2(n18858), .A(n18966), 
        .ZN(n18867) );
  NOR2_X1 U21998 ( .A1(n18859), .A2(n18867), .ZN(n18860) );
  MUX2_X1 U21999 ( .A(n18861), .B(n18860), .S(P3_STATE2_REG_0__SCAN_IN), .Z(
        n18863) );
  OAI211_X1 U22000 ( .C1(n18865), .C2(n18864), .A(n18863), .B(n18862), .ZN(
        P3_U2996) );
  NAND2_X1 U22001 ( .A1(n9998), .A2(n18866), .ZN(n18872) );
  NAND4_X1 U22002 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(
        P3_STATE2_REG_1__SCAN_IN), .A3(n9998), .A4(n19027), .ZN(n18874) );
  INV_X1 U22003 ( .A(n18867), .ZN(n18869) );
  NAND3_X1 U22004 ( .A1(n18870), .A2(n18869), .A3(n18868), .ZN(n18871) );
  NAND4_X1 U22005 ( .A1(n18873), .A2(n18872), .A3(n18874), .A4(n18871), .ZN(
        P3_U2997) );
  INV_X1 U22006 ( .A(n18874), .ZN(n18876) );
  NOR4_X1 U22007 ( .A1(n18878), .A2(n18877), .A3(n18876), .A4(n18875), .ZN(
        P3_U2998) );
  AND2_X1 U22008 ( .A1(P3_DATAWIDTH_REG_31__SCAN_IN), .A2(n18879), .ZN(
        P3_U2999) );
  AND2_X1 U22009 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n18879), .ZN(
        P3_U3000) );
  AND2_X1 U22010 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n18879), .ZN(
        P3_U3001) );
  AND2_X1 U22011 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n18879), .ZN(
        P3_U3002) );
  AND2_X1 U22012 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n18879), .ZN(
        P3_U3003) );
  AND2_X1 U22013 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n18879), .ZN(
        P3_U3004) );
  AND2_X1 U22014 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n18879), .ZN(
        P3_U3005) );
  AND2_X1 U22015 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n18879), .ZN(
        P3_U3006) );
  AND2_X1 U22016 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n18879), .ZN(
        P3_U3007) );
  AND2_X1 U22017 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n18879), .ZN(
        P3_U3008) );
  AND2_X1 U22018 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n18879), .ZN(
        P3_U3009) );
  INV_X1 U22019 ( .A(P3_DATAWIDTH_REG_20__SCAN_IN), .ZN(n21150) );
  NOR2_X1 U22020 ( .A1(n21150), .A2(n18964), .ZN(P3_U3010) );
  AND2_X1 U22021 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n18879), .ZN(
        P3_U3011) );
  AND2_X1 U22022 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n18879), .ZN(
        P3_U3012) );
  AND2_X1 U22023 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n18879), .ZN(
        P3_U3013) );
  AND2_X1 U22024 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n18879), .ZN(
        P3_U3014) );
  AND2_X1 U22025 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n18879), .ZN(
        P3_U3015) );
  AND2_X1 U22026 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n18879), .ZN(
        P3_U3016) );
  AND2_X1 U22027 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n18879), .ZN(
        P3_U3017) );
  AND2_X1 U22028 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n18879), .ZN(
        P3_U3018) );
  AND2_X1 U22029 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n18879), .ZN(
        P3_U3019) );
  AND2_X1 U22030 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n18879), .ZN(
        P3_U3020) );
  AND2_X1 U22031 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n18879), .ZN(P3_U3021) );
  AND2_X1 U22032 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n18879), .ZN(P3_U3022) );
  AND2_X1 U22033 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n18879), .ZN(P3_U3023) );
  AND2_X1 U22034 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n18879), .ZN(P3_U3024) );
  AND2_X1 U22035 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n18879), .ZN(P3_U3025) );
  AND2_X1 U22036 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n18879), .ZN(P3_U3026) );
  AND2_X1 U22037 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n18879), .ZN(P3_U3027) );
  AND2_X1 U22038 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n18879), .ZN(P3_U3028) );
  OAI21_X1 U22039 ( .B1(n20920), .B2(n18880), .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n18882) );
  NAND2_X1 U22040 ( .A1(n9998), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n18890) );
  NAND2_X1 U22041 ( .A1(n18890), .A2(P3_STATE_REG_0__SCAN_IN), .ZN(n18889) );
  INV_X1 U22042 ( .A(NA), .ZN(n20924) );
  OAI21_X1 U22043 ( .B1(n20924), .B2(n18881), .A(P3_STATE_REG_2__SCAN_IN), 
        .ZN(n18895) );
  AOI22_X1 U22044 ( .A1(n19025), .A2(n18882), .B1(n18889), .B2(n18895), .ZN(
        n18883) );
  INV_X1 U22045 ( .A(n18883), .ZN(P3_U3029) );
  NOR2_X1 U22046 ( .A1(n18897), .A2(n20920), .ZN(n18892) );
  INV_X1 U22047 ( .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n18884) );
  NOR3_X1 U22048 ( .A1(n18892), .A2(n18884), .A3(n18894), .ZN(n18886) );
  INV_X1 U22049 ( .A(n18890), .ZN(n18885) );
  NOR2_X1 U22050 ( .A1(n18886), .A2(n18885), .ZN(n18887) );
  OAI211_X1 U22051 ( .C1(n20920), .C2(n18888), .A(n18887), .B(n19011), .ZN(
        P3_U3030) );
  INV_X1 U22052 ( .A(n18889), .ZN(n18896) );
  OAI22_X1 U22053 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(
        P3_REQUESTPENDING_REG_SCAN_IN), .B1(NA), .B2(n18890), .ZN(n18891) );
  OAI22_X1 U22054 ( .A1(n18892), .A2(n18891), .B1(
        P3_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .ZN(n18893) );
  OAI22_X1 U22055 ( .A1(n18896), .A2(n18895), .B1(n18894), .B2(n18893), .ZN(
        P3_U3031) );
  INV_X1 U22056 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n18899) );
  OAI222_X1 U22057 ( .A1(n18999), .A2(n18954), .B1(n18898), .B2(n18960), .C1(
        n18899), .C2(n18946), .ZN(P3_U3032) );
  OAI222_X1 U22058 ( .A1(n18946), .A2(n18901), .B1(n18900), .B2(n18960), .C1(
        n18899), .C2(n18954), .ZN(P3_U3033) );
  OAI222_X1 U22059 ( .A1(n18946), .A2(n18903), .B1(n18902), .B2(n18960), .C1(
        n18901), .C2(n18954), .ZN(P3_U3034) );
  INV_X1 U22060 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n18906) );
  OAI222_X1 U22061 ( .A1(n18946), .A2(n18906), .B1(n18904), .B2(n18960), .C1(
        n18903), .C2(n18954), .ZN(P3_U3035) );
  OAI222_X1 U22062 ( .A1(n18906), .A2(n18954), .B1(n18905), .B2(n18960), .C1(
        n18907), .C2(n18946), .ZN(P3_U3036) );
  OAI222_X1 U22063 ( .A1(n18946), .A2(n18909), .B1(n18908), .B2(n18960), .C1(
        n18907), .C2(n18954), .ZN(P3_U3037) );
  INV_X1 U22064 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n21239) );
  OAI222_X1 U22065 ( .A1(n18946), .A2(n21239), .B1(n18910), .B2(n18960), .C1(
        n18909), .C2(n18954), .ZN(P3_U3038) );
  OAI222_X1 U22066 ( .A1(n21239), .A2(n18954), .B1(n18911), .B2(n18960), .C1(
        n18912), .C2(n18946), .ZN(P3_U3039) );
  OAI222_X1 U22067 ( .A1(n18946), .A2(n18914), .B1(n18913), .B2(n18960), .C1(
        n18912), .C2(n18954), .ZN(P3_U3040) );
  OAI222_X1 U22068 ( .A1(n18946), .A2(n18916), .B1(n18915), .B2(n18960), .C1(
        n18914), .C2(n18954), .ZN(P3_U3041) );
  OAI222_X1 U22069 ( .A1(n18946), .A2(n18918), .B1(n18917), .B2(n18960), .C1(
        n18916), .C2(n18954), .ZN(P3_U3042) );
  OAI222_X1 U22070 ( .A1(n18918), .A2(n18954), .B1(n21302), .B2(n18960), .C1(
        n18919), .C2(n18946), .ZN(P3_U3043) );
  OAI222_X1 U22071 ( .A1(n18946), .A2(n21228), .B1(n18920), .B2(n18960), .C1(
        n18919), .C2(n18954), .ZN(P3_U3044) );
  OAI222_X1 U22072 ( .A1(n21228), .A2(n18954), .B1(n21129), .B2(n18960), .C1(
        n18921), .C2(n18946), .ZN(P3_U3045) );
  OAI222_X1 U22073 ( .A1(n18946), .A2(n18923), .B1(n18922), .B2(n18960), .C1(
        n18921), .C2(n18954), .ZN(P3_U3046) );
  OAI222_X1 U22074 ( .A1(n18946), .A2(n18926), .B1(n18924), .B2(n18960), .C1(
        n18923), .C2(n18954), .ZN(P3_U3047) );
  OAI222_X1 U22075 ( .A1(n18926), .A2(n18954), .B1(n18925), .B2(n18960), .C1(
        n18927), .C2(n18946), .ZN(P3_U3048) );
  OAI222_X1 U22076 ( .A1(n18946), .A2(n18929), .B1(n18928), .B2(n18960), .C1(
        n18927), .C2(n18954), .ZN(P3_U3049) );
  OAI222_X1 U22077 ( .A1(n18946), .A2(n18931), .B1(n18930), .B2(n18960), .C1(
        n18929), .C2(n18954), .ZN(P3_U3050) );
  OAI222_X1 U22078 ( .A1(n18946), .A2(n18933), .B1(n18932), .B2(n18960), .C1(
        n18931), .C2(n18954), .ZN(P3_U3051) );
  OAI222_X1 U22079 ( .A1(n18946), .A2(n18935), .B1(n18934), .B2(n18960), .C1(
        n18933), .C2(n18954), .ZN(P3_U3052) );
  OAI222_X1 U22080 ( .A1(n18946), .A2(n18938), .B1(n18936), .B2(n18960), .C1(
        n18935), .C2(n18954), .ZN(P3_U3053) );
  OAI222_X1 U22081 ( .A1(n18938), .A2(n18954), .B1(n18937), .B2(n18960), .C1(
        n18939), .C2(n18946), .ZN(P3_U3054) );
  OAI222_X1 U22082 ( .A1(n18946), .A2(n18941), .B1(n18940), .B2(n18960), .C1(
        n18939), .C2(n18954), .ZN(P3_U3055) );
  OAI222_X1 U22083 ( .A1(n18946), .A2(n18943), .B1(n18942), .B2(n18960), .C1(
        n18941), .C2(n18954), .ZN(P3_U3056) );
  OAI222_X1 U22084 ( .A1(n18946), .A2(n18945), .B1(n18944), .B2(n18960), .C1(
        n18943), .C2(n18954), .ZN(P3_U3057) );
  OAI222_X1 U22085 ( .A1(n18946), .A2(n18948), .B1(n21093), .B2(n18960), .C1(
        n18945), .C2(n18954), .ZN(P3_U3058) );
  OAI222_X1 U22086 ( .A1(n18948), .A2(n18954), .B1(n18947), .B2(n18960), .C1(
        n18949), .C2(n18946), .ZN(P3_U3059) );
  INV_X1 U22087 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n18953) );
  OAI222_X1 U22088 ( .A1(n18946), .A2(n18953), .B1(n18950), .B2(n18960), .C1(
        n18949), .C2(n18954), .ZN(P3_U3060) );
  OAI222_X1 U22089 ( .A1(n18954), .A2(n18953), .B1(n18952), .B2(n18960), .C1(
        n18951), .C2(n18946), .ZN(P3_U3061) );
  INV_X1 U22090 ( .A(P3_BE_N_REG_3__SCAN_IN), .ZN(n18955) );
  AOI22_X1 U22091 ( .A1(n18960), .A2(n18956), .B1(n18955), .B2(n19025), .ZN(
        P3_U3274) );
  INV_X1 U22092 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n19001) );
  INV_X1 U22093 ( .A(P3_BE_N_REG_2__SCAN_IN), .ZN(n18957) );
  AOI22_X1 U22094 ( .A1(n18960), .A2(n19001), .B1(n18957), .B2(n19025), .ZN(
        P3_U3275) );
  INV_X1 U22095 ( .A(P3_BE_N_REG_1__SCAN_IN), .ZN(n18958) );
  AOI22_X1 U22096 ( .A1(n18960), .A2(n18959), .B1(n18958), .B2(n19025), .ZN(
        P3_U3276) );
  INV_X1 U22097 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n19007) );
  INV_X1 U22098 ( .A(P3_BE_N_REG_0__SCAN_IN), .ZN(n18961) );
  AOI22_X1 U22099 ( .A1(n18960), .A2(n19007), .B1(n18961), .B2(n19025), .ZN(
        P3_U3277) );
  OAI21_X1 U22100 ( .B1(n18964), .B2(P3_DATAWIDTH_REG_0__SCAN_IN), .A(n18963), 
        .ZN(n18962) );
  INV_X1 U22101 ( .A(n18962), .ZN(P3_U3280) );
  OAI21_X1 U22102 ( .B1(n18964), .B2(n21109), .A(n18963), .ZN(P3_U3281) );
  OAI221_X1 U22103 ( .B1(n18967), .B2(P3_STATE2_REG_0__SCAN_IN), .C1(n18967), 
        .C2(n18966), .A(n18965), .ZN(P3_U3282) );
  AOI22_X1 U22104 ( .A1(n19028), .A2(n18969), .B1(n18988), .B2(n18968), .ZN(
        n18974) );
  INV_X1 U22105 ( .A(n18970), .ZN(n18971) );
  AOI21_X1 U22106 ( .B1(n19028), .B2(n18971), .A(n18998), .ZN(n18973) );
  OAI22_X1 U22107 ( .A1(n18998), .A2(n18974), .B1(n18973), .B2(n18972), .ZN(
        P3_U3285) );
  AOI22_X1 U22108 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n18976), .B2(n18975), .ZN(
        n18984) );
  NOR2_X1 U22109 ( .A1(n18994), .A2(n18977), .ZN(n18985) );
  INV_X1 U22110 ( .A(n18988), .ZN(n18991) );
  OAI22_X1 U22111 ( .A1(n18979), .A2(n18993), .B1(n18991), .B2(n18978), .ZN(
        n18980) );
  AOI21_X1 U22112 ( .B1(n18984), .B2(n18985), .A(n18980), .ZN(n18981) );
  AOI22_X1 U22113 ( .A1(n18998), .A2(n18982), .B1(n18981), .B2(n18996), .ZN(
        P3_U3288) );
  INV_X1 U22114 ( .A(n18983), .ZN(n18989) );
  INV_X1 U22115 ( .A(n18984), .ZN(n18986) );
  AOI222_X1 U22116 ( .A1(n18989), .A2(n19028), .B1(n18988), .B2(n18987), .C1(
        n18986), .C2(n18985), .ZN(n18990) );
  AOI22_X1 U22117 ( .A1(n18998), .A2(n12506), .B1(n18990), .B2(n18996), .ZN(
        P3_U3289) );
  OAI222_X1 U22118 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n18994), .B1(
        n18993), .B2(n18992), .C1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .C2(
        n18991), .ZN(n18995) );
  INV_X1 U22119 ( .A(n18995), .ZN(n18997) );
  AOI21_X1 U22120 ( .B1(P3_REIP_REG_0__SCAN_IN), .B2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n19000) );
  AOI22_X1 U22121 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_0__SCAN_IN), 
        .B1(n19000), .B2(n18999), .ZN(n19002) );
  AOI22_X1 U22122 ( .A1(n19003), .A2(n19002), .B1(n19001), .B2(n19006), .ZN(
        P3_U3292) );
  NOR2_X1 U22123 ( .A1(n19006), .A2(P3_REIP_REG_1__SCAN_IN), .ZN(n19004) );
  AOI22_X1 U22124 ( .A1(n19007), .A2(n19006), .B1(n19005), .B2(n19004), .ZN(
        P3_U3293) );
  INV_X1 U22125 ( .A(P3_W_R_N_REG_SCAN_IN), .ZN(n19008) );
  AOI22_X1 U22126 ( .A1(n18960), .A2(P3_READREQUEST_REG_SCAN_IN), .B1(n19008), 
        .B2(n19025), .ZN(P3_U3294) );
  MUX2_X1 U22127 ( .A(P3_MORE_REG_SCAN_IN), .B(n19010), .S(n19009), .Z(
        P3_U3295) );
  AOI21_X1 U22128 ( .B1(n19013), .B2(n19012), .A(n19011), .ZN(n19014) );
  INV_X1 U22129 ( .A(n19014), .ZN(n19015) );
  AOI211_X1 U22130 ( .C1(n19029), .C2(n19015), .A(n9998), .B(n19027), .ZN(
        n19018) );
  OAI21_X1 U22131 ( .B1(n19018), .B2(n19017), .A(n19016), .ZN(n19024) );
  OAI22_X1 U22132 ( .A1(n9998), .A2(n19021), .B1(n19020), .B2(n19019), .ZN(
        n19022) );
  NOR2_X1 U22133 ( .A1(n19030), .A2(n19022), .ZN(n19023) );
  MUX2_X1 U22134 ( .A(n19024), .B(P3_REQUESTPENDING_REG_SCAN_IN), .S(n19023), 
        .Z(P3_U3296) );
  INV_X1 U22135 ( .A(P3_MEMORYFETCH_REG_SCAN_IN), .ZN(n19033) );
  INV_X1 U22136 ( .A(P3_M_IO_N_REG_SCAN_IN), .ZN(n19026) );
  AOI22_X1 U22137 ( .A1(n18960), .A2(n19033), .B1(n19026), .B2(n19025), .ZN(
        P3_U3297) );
  AOI21_X1 U22138 ( .B1(n19028), .B2(n19027), .A(n19030), .ZN(n19034) );
  INV_X1 U22139 ( .A(P3_READREQUEST_REG_SCAN_IN), .ZN(n19031) );
  AOI22_X1 U22140 ( .A1(n19034), .A2(n19031), .B1(n19030), .B2(n19029), .ZN(
        P3_U3298) );
  AOI21_X1 U22141 ( .B1(n19034), .B2(n19033), .A(n19032), .ZN(P3_U3299) );
  INV_X1 U22142 ( .A(P2_ADS_N_REG_SCAN_IN), .ZN(n19035) );
  NAND2_X1 U22143 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n19933), .ZN(n19922) );
  NAND2_X1 U22144 ( .A1(n21257), .A2(n19915), .ZN(n19919) );
  OAI21_X1 U22145 ( .B1(n21257), .B2(n19035), .A(n19914), .ZN(P2_U2815) );
  INV_X1 U22146 ( .A(P2_CODEFETCH_REG_SCAN_IN), .ZN(n19036) );
  OAI22_X1 U22147 ( .A1(n19038), .A2(n19037), .B1(n20056), .B2(n19036), .ZN(
        P2_U2816) );
  NAND2_X1 U22148 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n21257), .ZN(n20075) );
  AOI21_X1 U22149 ( .B1(n21257), .B2(n19933), .A(P2_D_C_N_REG_SCAN_IN), .ZN(
        n19039) );
  AOI22_X1 U22150 ( .A1(n19994), .A2(P2_CODEFETCH_REG_SCAN_IN), .B1(n19039), 
        .B2(n20075), .ZN(P2_U2817) );
  OAI21_X1 U22151 ( .B1(n19927), .B2(BS16), .A(n20000), .ZN(n19998) );
  OAI21_X1 U22152 ( .B1(n20000), .B2(n20061), .A(n19998), .ZN(P2_U2818) );
  NOR2_X1 U22153 ( .A1(n19041), .A2(n19040), .ZN(n20054) );
  OAI21_X1 U22154 ( .B1(n20054), .B2(n11393), .A(n19042), .ZN(P2_U2819) );
  NOR4_X1 U22155 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_21__SCAN_IN), .A3(P2_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_23__SCAN_IN), .ZN(n19046) );
  NOR4_X1 U22156 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_17__SCAN_IN), .A3(P2_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_19__SCAN_IN), .ZN(n19045) );
  NOR4_X1 U22157 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_29__SCAN_IN), .A3(P2_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_31__SCAN_IN), .ZN(n19044) );
  NOR4_X1 U22158 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_25__SCAN_IN), .A3(P2_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_27__SCAN_IN), .ZN(n19043) );
  NAND4_X1 U22159 ( .A1(n19046), .A2(n19045), .A3(n19044), .A4(n19043), .ZN(
        n19052) );
  NOR4_X1 U22160 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_4__SCAN_IN), .A3(P2_DATAWIDTH_REG_5__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_6__SCAN_IN), .ZN(n19050) );
  AOI211_X1 U22161 ( .C1(P2_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_0__SCAN_IN), .A(P2_DATAWIDTH_REG_8__SCAN_IN), .B(
        P2_DATAWIDTH_REG_2__SCAN_IN), .ZN(n19049) );
  NOR4_X1 U22162 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_13__SCAN_IN), .A3(P2_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_15__SCAN_IN), .ZN(n19048) );
  NOR4_X1 U22163 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_9__SCAN_IN), .A3(P2_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_11__SCAN_IN), .ZN(n19047) );
  NAND4_X1 U22164 ( .A1(n19050), .A2(n19049), .A3(n19048), .A4(n19047), .ZN(
        n19051) );
  NOR2_X1 U22165 ( .A1(n19052), .A2(n19051), .ZN(n19060) );
  INV_X1 U22166 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n19996) );
  OAI21_X1 U22167 ( .B1(P2_REIP_REG_0__SCAN_IN), .B2(P2_REIP_REG_1__SCAN_IN), 
        .A(n19060), .ZN(n19053) );
  OAI21_X1 U22168 ( .B1(n19060), .B2(n19996), .A(n19053), .ZN(P2_U2820) );
  INV_X1 U22169 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n19993) );
  NOR3_X1 U22170 ( .A1(P2_REIP_REG_0__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_1__SCAN_IN), .A3(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n19057) );
  OAI21_X1 U22171 ( .B1(P2_REIP_REG_1__SCAN_IN), .B2(n19057), .A(n19060), .ZN(
        n19054) );
  OAI21_X1 U22172 ( .B1(n19060), .B2(n19993), .A(n19054), .ZN(P2_U2821) );
  AOI21_X1 U22173 ( .B1(P2_REIP_REG_0__SCAN_IN), .B2(
        P2_DATAWIDTH_REG_0__SCAN_IN), .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n19055) );
  OAI22_X1 U22174 ( .A1(P2_REIP_REG_0__SCAN_IN), .A2(n19934), .B1(
        P2_REIP_REG_1__SCAN_IN), .B2(n19055), .ZN(n19056) );
  INV_X1 U22175 ( .A(P2_BYTEENABLE_REG_2__SCAN_IN), .ZN(n19991) );
  INV_X1 U22176 ( .A(n19060), .ZN(n19058) );
  AOI22_X1 U22177 ( .A1(n19060), .A2(n19056), .B1(n19991), .B2(n19058), .ZN(
        P2_U2822) );
  INV_X1 U22178 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n19999) );
  AOI21_X1 U22179 ( .B1(n19934), .B2(n19999), .A(n19057), .ZN(n19059) );
  INV_X1 U22180 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n19989) );
  AOI22_X1 U22181 ( .A1(n19060), .A2(n19059), .B1(n19989), .B2(n19058), .ZN(
        P2_U2823) );
  NAND2_X1 U22182 ( .A1(n10135), .A2(n19061), .ZN(n19062) );
  XOR2_X1 U22183 ( .A(n19063), .B(n19062), .Z(n19073) );
  OAI21_X1 U22184 ( .B1(n19962), .B2(n19181), .A(n19345), .ZN(n19067) );
  OAI22_X1 U22185 ( .A1(n19065), .A2(n19202), .B1(n19064), .B2(n19180), .ZN(
        n19066) );
  AOI211_X1 U22186 ( .C1(P2_EBX_REG_19__SCAN_IN), .C2(n19205), .A(n19067), .B(
        n19066), .ZN(n19072) );
  INV_X1 U22187 ( .A(n19068), .ZN(n19069) );
  AOI22_X1 U22188 ( .A1(n19070), .A2(n19179), .B1(n19183), .B2(n19069), .ZN(
        n19071) );
  OAI211_X1 U22189 ( .C1(n19214), .C2(n19073), .A(n19072), .B(n19071), .ZN(
        P2_U2836) );
  NAND2_X1 U22190 ( .A1(n10135), .A2(n19074), .ZN(n19075) );
  XOR2_X1 U22191 ( .A(n19076), .B(n19075), .Z(n19085) );
  AOI22_X1 U22192 ( .A1(n19077), .A2(n19186), .B1(
        P2_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n19166), .ZN(n19078) );
  OAI211_X1 U22193 ( .C1(n19959), .C2(n19181), .A(n19078), .B(n19345), .ZN(
        n19079) );
  AOI21_X1 U22194 ( .B1(P2_EBX_REG_17__SCAN_IN), .B2(n19205), .A(n19079), .ZN(
        n19084) );
  INV_X1 U22195 ( .A(n19080), .ZN(n19081) );
  AOI22_X1 U22196 ( .A1(n19082), .A2(n19179), .B1(n19183), .B2(n19081), .ZN(
        n19083) );
  OAI211_X1 U22197 ( .C1(n19214), .C2(n19085), .A(n19084), .B(n19083), .ZN(
        P2_U2838) );
  NAND2_X1 U22198 ( .A1(n10135), .A2(n19086), .ZN(n19088) );
  XOR2_X1 U22199 ( .A(n19088), .B(n19087), .Z(n19095) );
  AOI22_X1 U22200 ( .A1(n19089), .A2(n19186), .B1(P2_EBX_REG_15__SCAN_IN), 
        .B2(n19205), .ZN(n19090) );
  OAI211_X1 U22201 ( .C1(n19956), .C2(n19181), .A(n19090), .B(n19345), .ZN(
        n19093) );
  OAI22_X1 U22202 ( .A1(n19091), .A2(n19197), .B1(n19200), .B2(n19231), .ZN(
        n19092) );
  AOI211_X1 U22203 ( .C1(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(n19211), .A(
        n19093), .B(n19092), .ZN(n19094) );
  OAI21_X1 U22204 ( .B1(n19095), .B2(n19214), .A(n19094), .ZN(P2_U2840) );
  NOR2_X1 U22205 ( .A1(n19159), .A2(n19096), .ZN(n19098) );
  XOR2_X1 U22206 ( .A(n19098), .B(n19097), .Z(n19106) );
  AOI22_X1 U22207 ( .A1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n19166), .B1(
        P2_EBX_REG_14__SCAN_IN), .B2(n19205), .ZN(n19099) );
  OAI21_X1 U22208 ( .B1(n19100), .B2(n19202), .A(n19099), .ZN(n19101) );
  AOI211_X1 U22209 ( .C1(P2_REIP_REG_14__SCAN_IN), .C2(n19210), .A(n19170), 
        .B(n19101), .ZN(n19105) );
  AOI22_X1 U22210 ( .A1(n19103), .A2(n19183), .B1(n19179), .B2(n19102), .ZN(
        n19104) );
  OAI211_X1 U22211 ( .C1(n19214), .C2(n19106), .A(n19105), .B(n19104), .ZN(
        P2_U2841) );
  NAND2_X1 U22212 ( .A1(n10135), .A2(n19107), .ZN(n19108) );
  XNOR2_X1 U22213 ( .A(n19109), .B(n19108), .ZN(n19119) );
  OAI21_X1 U22214 ( .B1(n15855), .B2(n19181), .A(n19345), .ZN(n19114) );
  INV_X1 U22215 ( .A(n19110), .ZN(n19112) );
  OAI22_X1 U22216 ( .A1(n19112), .A2(n19202), .B1(n19111), .B2(n19180), .ZN(
        n19113) );
  AOI211_X1 U22217 ( .C1(P2_EBX_REG_13__SCAN_IN), .C2(n19205), .A(n19114), .B(
        n19113), .ZN(n19118) );
  INV_X1 U22218 ( .A(n19115), .ZN(n19116) );
  AOI22_X1 U22219 ( .A1(n19235), .A2(n19183), .B1(n19179), .B2(n19116), .ZN(
        n19117) );
  OAI211_X1 U22220 ( .C1(n19214), .C2(n19119), .A(n19118), .B(n19117), .ZN(
        P2_U2842) );
  AOI22_X1 U22221 ( .A1(n19120), .A2(n19186), .B1(
        P2_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n19166), .ZN(n19121) );
  OAI21_X1 U22222 ( .B1(n19155), .B2(n19122), .A(n19121), .ZN(n19123) );
  AOI211_X1 U22223 ( .C1(P2_REIP_REG_11__SCAN_IN), .C2(n19210), .A(n19170), 
        .B(n19123), .ZN(n19130) );
  NAND2_X1 U22224 ( .A1(n10135), .A2(n19124), .ZN(n19125) );
  XNOR2_X1 U22225 ( .A(n19126), .B(n19125), .ZN(n19128) );
  AOI22_X1 U22226 ( .A1(n19128), .A2(n19175), .B1(n19179), .B2(n19127), .ZN(
        n19129) );
  OAI211_X1 U22227 ( .C1(n19243), .C2(n19200), .A(n19130), .B(n19129), .ZN(
        P2_U2844) );
  NAND2_X1 U22228 ( .A1(n10135), .A2(n19131), .ZN(n19133) );
  XOR2_X1 U22229 ( .A(n19133), .B(n19132), .Z(n19141) );
  AOI22_X1 U22230 ( .A1(n19134), .A2(n19186), .B1(P2_EBX_REG_9__SCAN_IN), .B2(
        n19205), .ZN(n19135) );
  OAI211_X1 U22231 ( .C1(n19948), .C2(n19181), .A(n19135), .B(n19345), .ZN(
        n19139) );
  INV_X1 U22232 ( .A(n19136), .ZN(n19137) );
  OAI22_X1 U22233 ( .A1(n19200), .A2(n19248), .B1(n19197), .B2(n19137), .ZN(
        n19138) );
  AOI211_X1 U22234 ( .C1(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .C2(n19211), .A(
        n19139), .B(n19138), .ZN(n19140) );
  OAI21_X1 U22235 ( .B1(n19141), .B2(n19214), .A(n19140), .ZN(P2_U2846) );
  NAND2_X1 U22236 ( .A1(n10135), .A2(n19142), .ZN(n19144) );
  XOR2_X1 U22237 ( .A(n19144), .B(n19143), .Z(n19152) );
  INV_X1 U22238 ( .A(n19145), .ZN(n19146) );
  AOI22_X1 U22239 ( .A1(n19146), .A2(n19186), .B1(n19205), .B2(
        P2_EBX_REG_7__SCAN_IN), .ZN(n19147) );
  OAI211_X1 U22240 ( .C1(n19945), .C2(n19181), .A(n19147), .B(n19345), .ZN(
        n19150) );
  OAI22_X1 U22241 ( .A1(n19200), .A2(n19253), .B1(n19197), .B2(n19148), .ZN(
        n19149) );
  AOI211_X1 U22242 ( .C1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .C2(n19211), .A(
        n19150), .B(n19149), .ZN(n19151) );
  OAI21_X1 U22243 ( .B1(n19152), .B2(n19214), .A(n19151), .ZN(P2_U2848) );
  OAI21_X1 U22244 ( .B1(n19943), .B2(n19181), .A(n19345), .ZN(n19157) );
  INV_X1 U22245 ( .A(P2_EBX_REG_6__SCAN_IN), .ZN(n19154) );
  OAI22_X1 U22246 ( .A1(n19155), .A2(n19154), .B1(n19202), .B2(n19153), .ZN(
        n19156) );
  AOI211_X1 U22247 ( .C1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .C2(n19211), .A(
        n19157), .B(n19156), .ZN(n19165) );
  NOR2_X1 U22248 ( .A1(n19159), .A2(n19158), .ZN(n19161) );
  XNOR2_X1 U22249 ( .A(n19161), .B(n19160), .ZN(n19163) );
  AOI22_X1 U22250 ( .A1(n19163), .A2(n19175), .B1(n19179), .B2(n19162), .ZN(
        n19164) );
  OAI211_X1 U22251 ( .C1(n19200), .C2(n19256), .A(n19165), .B(n19164), .ZN(
        P2_U2849) );
  AOI22_X1 U22252 ( .A1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n19166), .B1(
        P2_EBX_REG_5__SCAN_IN), .B2(n19205), .ZN(n19167) );
  OAI21_X1 U22253 ( .B1(n19202), .B2(n19168), .A(n19167), .ZN(n19169) );
  AOI211_X1 U22254 ( .C1(P2_REIP_REG_5__SCAN_IN), .C2(n19210), .A(n19170), .B(
        n19169), .ZN(n19178) );
  NAND2_X1 U22255 ( .A1(n10135), .A2(n19171), .ZN(n19172) );
  XNOR2_X1 U22256 ( .A(n19173), .B(n19172), .ZN(n19176) );
  AOI22_X1 U22257 ( .A1(n19176), .A2(n19175), .B1(n19179), .B2(n19174), .ZN(
        n19177) );
  OAI211_X1 U22258 ( .C1(n19200), .C2(n19263), .A(n19178), .B(n19177), .ZN(
        P2_U2850) );
  NAND2_X1 U22259 ( .A1(n9860), .A2(n19179), .ZN(n19190) );
  OAI22_X1 U22260 ( .A1(n19934), .A2(n19181), .B1(n19191), .B2(n19180), .ZN(
        n19182) );
  AOI21_X1 U22261 ( .B1(n19183), .B2(n20031), .A(n19182), .ZN(n19189) );
  NAND2_X1 U22262 ( .A1(n19205), .A2(P2_EBX_REG_1__SCAN_IN), .ZN(n19188) );
  INV_X1 U22263 ( .A(n19184), .ZN(n19185) );
  NAND2_X1 U22264 ( .A1(n19186), .A2(n19185), .ZN(n19187) );
  AND4_X1 U22265 ( .A1(n19190), .A2(n19189), .A3(n19188), .A4(n19187), .ZN(
        n19195) );
  AOI22_X1 U22266 ( .A1(n20029), .A2(n19193), .B1(n19192), .B2(n19191), .ZN(
        n19194) );
  OAI211_X1 U22267 ( .C1(n19214), .C2(n19196), .A(n19195), .B(n19194), .ZN(
        P2_U2854) );
  NOR2_X1 U22268 ( .A1(n19198), .A2(n19197), .ZN(n19204) );
  OAI22_X1 U22269 ( .A1(n19202), .A2(n19201), .B1(n19200), .B2(n19199), .ZN(
        n19203) );
  AOI211_X1 U22270 ( .C1(P2_EBX_REG_0__SCAN_IN), .C2(n19205), .A(n19204), .B(
        n19203), .ZN(n19206) );
  OAI21_X1 U22271 ( .B1(n19208), .B2(n19207), .A(n19206), .ZN(n19209) );
  AOI21_X1 U22272 ( .B1(P2_REIP_REG_0__SCAN_IN), .B2(n19210), .A(n19209), .ZN(
        n19213) );
  NAND2_X1 U22273 ( .A1(P2_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n19211), .ZN(
        n19212) );
  OAI211_X1 U22274 ( .C1(n19215), .C2(n19214), .A(n19213), .B(n19212), .ZN(
        P2_U2855) );
  INV_X1 U22275 ( .A(n19216), .ZN(n19217) );
  AOI22_X1 U22276 ( .A1(n19222), .A2(BUF1_REG_31__SCAN_IN), .B1(n19265), .B2(
        n19217), .ZN(n19219) );
  AOI22_X1 U22277 ( .A1(P2_EAX_REG_31__SCAN_IN), .A2(n19257), .B1(n19223), 
        .B2(BUF2_REG_31__SCAN_IN), .ZN(n19218) );
  NAND2_X1 U22278 ( .A1(n19219), .A2(n19218), .ZN(P2_U2888) );
  AOI22_X1 U22279 ( .A1(n19221), .A2(n19220), .B1(n19257), .B2(
        P2_EAX_REG_16__SCAN_IN), .ZN(n19228) );
  AOI22_X1 U22280 ( .A1(n19223), .A2(BUF2_REG_16__SCAN_IN), .B1(n19222), .B2(
        BUF1_REG_16__SCAN_IN), .ZN(n19227) );
  AOI22_X1 U22281 ( .A1(n19225), .A2(n19270), .B1(n19265), .B2(n19224), .ZN(
        n19226) );
  NAND3_X1 U22282 ( .A1(n19228), .A2(n19227), .A3(n19226), .ZN(P2_U2903) );
  OAI222_X1 U22283 ( .A1(n19231), .A2(n19264), .B1(n19280), .B2(n19274), .C1(
        n19230), .C2(n19255), .ZN(P2_U2904) );
  AOI22_X1 U22284 ( .A1(P2_EAX_REG_14__SCAN_IN), .A2(n19257), .B1(n19232), 
        .B2(n19266), .ZN(n19233) );
  OAI21_X1 U22285 ( .B1(n19264), .B2(n19234), .A(n19233), .ZN(P2_U2905) );
  INV_X1 U22286 ( .A(n19235), .ZN(n19237) );
  INV_X1 U22287 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n19284) );
  OAI222_X1 U22288 ( .A1(n19237), .A2(n19264), .B1(n19284), .B2(n19274), .C1(
        n19255), .C2(n19236), .ZN(P2_U2906) );
  INV_X1 U22289 ( .A(n19238), .ZN(n19241) );
  AOI22_X1 U22290 ( .A1(P2_EAX_REG_12__SCAN_IN), .A2(n19257), .B1(n19239), 
        .B2(n19266), .ZN(n19240) );
  OAI21_X1 U22291 ( .B1(n19264), .B2(n19241), .A(n19240), .ZN(P2_U2907) );
  INV_X1 U22292 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n19287) );
  OAI222_X1 U22293 ( .A1(n19243), .A2(n19264), .B1(n19287), .B2(n19274), .C1(
        n19255), .C2(n19242), .ZN(P2_U2908) );
  INV_X1 U22294 ( .A(n19264), .ZN(n19250) );
  AOI22_X1 U22295 ( .A1(n19245), .A2(n19250), .B1(n19244), .B2(n19266), .ZN(
        n19246) );
  OAI21_X1 U22296 ( .B1(n19274), .B2(n19289), .A(n19246), .ZN(P2_U2909) );
  INV_X1 U22297 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n19291) );
  OAI222_X1 U22298 ( .A1(n19248), .A2(n19264), .B1(n19291), .B2(n19274), .C1(
        n19255), .C2(n19247), .ZN(P2_U2910) );
  AOI22_X1 U22299 ( .A1(n19251), .A2(n19250), .B1(n19249), .B2(n19266), .ZN(
        n19252) );
  OAI21_X1 U22300 ( .B1(n19274), .B2(n19293), .A(n19252), .ZN(P2_U2911) );
  INV_X1 U22301 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n19295) );
  OAI222_X1 U22302 ( .A1(n19253), .A2(n19264), .B1(n19295), .B2(n19274), .C1(
        n19255), .C2(n19417), .ZN(P2_U2912) );
  INV_X1 U22303 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n19297) );
  INV_X1 U22304 ( .A(n19409), .ZN(n19254) );
  OAI222_X1 U22305 ( .A1(n19256), .A2(n19264), .B1(n19297), .B2(n19274), .C1(
        n19255), .C2(n19254), .ZN(P2_U2913) );
  AOI22_X1 U22306 ( .A1(P2_EAX_REG_5__SCAN_IN), .A2(n19257), .B1(n19403), .B2(
        n19266), .ZN(n19262) );
  OR3_X1 U22307 ( .A1(n19260), .A2(n19259), .A3(n19258), .ZN(n19261) );
  OAI211_X1 U22308 ( .C1(n19264), .C2(n19263), .A(n19262), .B(n19261), .ZN(
        P2_U2914) );
  INV_X1 U22309 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n19305) );
  AOI22_X1 U22310 ( .A1(n19266), .A2(n19381), .B1(n19265), .B2(n20021), .ZN(
        n19273) );
  OAI21_X1 U22311 ( .B1(n19269), .B2(n19268), .A(n19267), .ZN(n19271) );
  NAND2_X1 U22312 ( .A1(n19271), .A2(n19270), .ZN(n19272) );
  OAI211_X1 U22313 ( .C1(n19274), .C2(n19305), .A(n19273), .B(n19272), .ZN(
        P2_U2917) );
  NOR2_X1 U22314 ( .A1(n19312), .A2(n19275), .ZN(P2_U2920) );
  INV_X1 U22315 ( .A(n19276), .ZN(n19277) );
  AOI22_X1 U22316 ( .A1(n19277), .A2(P2_EAX_REG_22__SCAN_IN), .B1(n20057), 
        .B2(P2_UWORD_REG_6__SCAN_IN), .ZN(n19278) );
  OAI21_X1 U22317 ( .B1(n21269), .B2(n19312), .A(n19278), .ZN(P2_U2929) );
  OAI222_X1 U22318 ( .A1(n19309), .A2(n21222), .B1(n19308), .B2(n19280), .C1(
        n19312), .C2(n19279), .ZN(P2_U2936) );
  AOI22_X1 U22319 ( .A1(n20057), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n19303), 
        .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n19281) );
  OAI21_X1 U22320 ( .B1(n19282), .B2(n19308), .A(n19281), .ZN(P2_U2937) );
  AOI22_X1 U22321 ( .A1(n20057), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n19303), 
        .B2(P2_DATAO_REG_13__SCAN_IN), .ZN(n19283) );
  OAI21_X1 U22322 ( .B1(n19284), .B2(n19308), .A(n19283), .ZN(P2_U2938) );
  AOI22_X1 U22323 ( .A1(P2_EAX_REG_12__SCAN_IN), .A2(n19310), .B1(n19303), 
        .B2(P2_DATAO_REG_12__SCAN_IN), .ZN(n19285) );
  OAI21_X1 U22324 ( .B1(n21221), .B2(n19309), .A(n19285), .ZN(P2_U2939) );
  AOI22_X1 U22325 ( .A1(n20057), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n19303), 
        .B2(P2_DATAO_REG_11__SCAN_IN), .ZN(n19286) );
  OAI21_X1 U22326 ( .B1(n19287), .B2(n19308), .A(n19286), .ZN(P2_U2940) );
  INV_X1 U22327 ( .A(P2_LWORD_REG_10__SCAN_IN), .ZN(n21284) );
  OAI222_X1 U22328 ( .A1(n19309), .A2(n21284), .B1(n19308), .B2(n19289), .C1(
        n19312), .C2(n19288), .ZN(P2_U2941) );
  AOI22_X1 U22329 ( .A1(n20057), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n19303), 
        .B2(P2_DATAO_REG_9__SCAN_IN), .ZN(n19290) );
  OAI21_X1 U22330 ( .B1(n19291), .B2(n19308), .A(n19290), .ZN(P2_U2942) );
  AOI22_X1 U22331 ( .A1(n20057), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n19303), 
        .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n19292) );
  OAI21_X1 U22332 ( .B1(n19293), .B2(n19308), .A(n19292), .ZN(P2_U2943) );
  AOI22_X1 U22333 ( .A1(n20057), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n19303), 
        .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n19294) );
  OAI21_X1 U22334 ( .B1(n19295), .B2(n19308), .A(n19294), .ZN(P2_U2944) );
  AOI22_X1 U22335 ( .A1(n20057), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n19303), 
        .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n19296) );
  OAI21_X1 U22336 ( .B1(n19297), .B2(n19308), .A(n19296), .ZN(P2_U2945) );
  INV_X1 U22337 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n19299) );
  AOI22_X1 U22338 ( .A1(n20057), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n19303), 
        .B2(P2_DATAO_REG_5__SCAN_IN), .ZN(n19298) );
  OAI21_X1 U22339 ( .B1(n19299), .B2(n19308), .A(n19298), .ZN(P2_U2946) );
  AOI22_X1 U22340 ( .A1(n20057), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n19303), 
        .B2(P2_DATAO_REG_4__SCAN_IN), .ZN(n19300) );
  OAI21_X1 U22341 ( .B1(n19301), .B2(n19308), .A(n19300), .ZN(P2_U2947) );
  AOI22_X1 U22342 ( .A1(n20057), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n19303), 
        .B2(P2_DATAO_REG_3__SCAN_IN), .ZN(n19302) );
  OAI21_X1 U22343 ( .B1(n13652), .B2(n19308), .A(n19302), .ZN(P2_U2948) );
  AOI22_X1 U22344 ( .A1(n20057), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n19303), 
        .B2(P2_DATAO_REG_2__SCAN_IN), .ZN(n19304) );
  OAI21_X1 U22345 ( .B1(n19305), .B2(n19308), .A(n19304), .ZN(P2_U2949) );
  INV_X1 U22346 ( .A(P2_LWORD_REG_1__SCAN_IN), .ZN(n21236) );
  INV_X1 U22347 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n19307) );
  OAI222_X1 U22348 ( .A1(n19309), .A2(n21236), .B1(n19308), .B2(n19307), .C1(
        n19312), .C2(n19306), .ZN(P2_U2950) );
  AOI22_X1 U22349 ( .A1(P2_EAX_REG_0__SCAN_IN), .A2(n19310), .B1(n20057), .B2(
        P2_LWORD_REG_0__SCAN_IN), .ZN(n19311) );
  OAI21_X1 U22350 ( .B1(n21122), .B2(n19312), .A(n19311), .ZN(P2_U2951) );
  AOI22_X1 U22351 ( .A1(n19313), .A2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B1(
        P2_REIP_REG_4__SCAN_IN), .B2(n19170), .ZN(n19323) );
  NAND2_X1 U22352 ( .A1(n19314), .A2(n12840), .ZN(n19318) );
  NAND2_X1 U22353 ( .A1(n19316), .A2(n19315), .ZN(n19317) );
  OAI211_X1 U22354 ( .C1(n19320), .C2(n19319), .A(n19318), .B(n19317), .ZN(
        n19321) );
  INV_X1 U22355 ( .A(n19321), .ZN(n19322) );
  OAI211_X1 U22356 ( .C1(n19325), .C2(n19324), .A(n19323), .B(n19322), .ZN(
        P2_U3010) );
  INV_X1 U22357 ( .A(n20021), .ZN(n19328) );
  OAI22_X1 U22358 ( .A1(n19328), .A2(n19327), .B1(n19356), .B2(n19326), .ZN(
        n19329) );
  AOI21_X1 U22359 ( .B1(n19331), .B2(n19330), .A(n19329), .ZN(n19344) );
  INV_X1 U22360 ( .A(n19332), .ZN(n19340) );
  NOR2_X1 U22361 ( .A1(n19333), .A2(n19346), .ZN(n19338) );
  NAND2_X1 U22362 ( .A1(n19334), .A2(n19346), .ZN(n19335) );
  OAI211_X1 U22363 ( .C1(n19346), .C2(n19336), .A(n19335), .B(n19349), .ZN(
        n19337) );
  MUX2_X1 U22364 ( .A(n19338), .B(n19337), .S(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .Z(n19339) );
  AOI211_X1 U22365 ( .C1(n19342), .C2(n19341), .A(n19340), .B(n19339), .ZN(
        n19343) );
  OAI211_X1 U22366 ( .C1(n19936), .C2(n19345), .A(n19344), .B(n19343), .ZN(
        P2_U3044) );
  OAI21_X1 U22367 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(n19346), .ZN(n19352) );
  NAND2_X1 U22368 ( .A1(n19347), .A2(n20031), .ZN(n19351) );
  OR2_X1 U22369 ( .A1(n19349), .A2(n19348), .ZN(n19350) );
  OAI211_X1 U22370 ( .C1(n19353), .C2(n19352), .A(n19351), .B(n19350), .ZN(
        n19359) );
  OAI22_X1 U22371 ( .A1(n19357), .A2(n19356), .B1(n19355), .B2(n19354), .ZN(
        n19358) );
  NOR2_X1 U22372 ( .A1(n19359), .A2(n19358), .ZN(n19361) );
  OAI211_X1 U22373 ( .C1(n19363), .C2(n19362), .A(n19361), .B(n19360), .ZN(
        P2_U3045) );
  INV_X1 U22374 ( .A(n19454), .ZN(n19365) );
  NAND3_X1 U22375 ( .A1(n19370), .A2(n20006), .A3(n19365), .ZN(n19366) );
  NOR2_X1 U22376 ( .A1(n20002), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19635) );
  INV_X1 U22377 ( .A(n19635), .ZN(n19804) );
  NAND2_X1 U22378 ( .A1(n19366), .A2(n19804), .ZN(n19371) );
  NOR2_X1 U22379 ( .A1(n19367), .A2(n20017), .ZN(n19903) );
  NOR2_X1 U22380 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19458) );
  NAND2_X1 U22381 ( .A1(n19368), .A2(n19458), .ZN(n19372) );
  OR2_X1 U22382 ( .A1(n19903), .A2(n19421), .ZN(n19375) );
  AOI21_X1 U22383 ( .B1(n19373), .B2(n19372), .A(n20034), .ZN(n19369) );
  AOI22_X1 U22384 ( .A1(n19908), .A2(n19808), .B1(n19855), .B2(n19421), .ZN(
        n19378) );
  INV_X1 U22385 ( .A(n19371), .ZN(n19376) );
  OAI211_X1 U22386 ( .C1(n19373), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19372), 
        .B(n20002), .ZN(n19374) );
  OAI211_X1 U22387 ( .C1(n19376), .C2(n19375), .A(n19861), .B(n19374), .ZN(
        n19426) );
  AOI22_X1 U22388 ( .A1(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n19426), .B1(
        n19454), .B2(n19863), .ZN(n19377) );
  OAI211_X1 U22389 ( .C1(n19429), .C2(n19817), .A(n19378), .B(n19377), .ZN(
        P2_U3048) );
  AOI22_X1 U22390 ( .A1(n19908), .A2(n19818), .B1(n19867), .B2(n19421), .ZN(
        n19380) );
  AOI22_X1 U22391 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n19426), .B1(
        n19454), .B2(n19869), .ZN(n19379) );
  OAI211_X1 U22392 ( .C1(n19429), .C2(n19821), .A(n19380), .B(n19379), .ZN(
        P2_U3049) );
  NAND2_X1 U22393 ( .A1(n19381), .A2(n19861), .ZN(n19825) );
  OAI22_X2 U22394 ( .A1(n19383), .A2(n19424), .B1(n19382), .B2(n19422), .ZN(
        n19822) );
  AOI22_X1 U22395 ( .A1(n19908), .A2(n19822), .B1(n9966), .B2(n19421), .ZN(
        n19387) );
  OAI22_X2 U22396 ( .A1(n15095), .A2(n19424), .B1(n19385), .B2(n19422), .ZN(
        n19875) );
  AOI22_X1 U22397 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n19426), .B1(
        n19454), .B2(n19875), .ZN(n19386) );
  OAI211_X1 U22398 ( .C1(n19429), .C2(n19825), .A(n19387), .B(n19386), .ZN(
        P2_U3050) );
  NAND2_X1 U22399 ( .A1(n19388), .A2(n19861), .ZN(n19829) );
  AOI22_X1 U22400 ( .A1(n19908), .A2(n19826), .B1(n19879), .B2(n19421), .ZN(
        n19395) );
  OAI22_X2 U22401 ( .A1(n19393), .A2(n19424), .B1(n19392), .B2(n19422), .ZN(
        n19881) );
  AOI22_X1 U22402 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n19426), .B1(
        n19454), .B2(n19881), .ZN(n19394) );
  OAI211_X1 U22403 ( .C1(n19429), .C2(n19829), .A(n19395), .B(n19394), .ZN(
        P2_U3051) );
  NAND2_X1 U22404 ( .A1(n19396), .A2(n19861), .ZN(n19833) );
  NOR2_X2 U22405 ( .A1(n10936), .A2(n19412), .ZN(n19885) );
  AOI22_X1 U22406 ( .A1(n19908), .A2(n19830), .B1(n19885), .B2(n19421), .ZN(
        n19402) );
  OAI22_X2 U22407 ( .A1(n19400), .A2(n19424), .B1(n19399), .B2(n19422), .ZN(
        n19887) );
  AOI22_X1 U22408 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n19426), .B1(
        n19454), .B2(n19887), .ZN(n19401) );
  OAI211_X1 U22409 ( .C1(n19429), .C2(n19833), .A(n19402), .B(n19401), .ZN(
        P2_U3052) );
  NAND2_X1 U22410 ( .A1(n19403), .A2(n19861), .ZN(n19837) );
  NOR2_X2 U22411 ( .A1(n10543), .A2(n19412), .ZN(n19891) );
  AOI22_X1 U22412 ( .A1(n19908), .A2(n19834), .B1(n19891), .B2(n19421), .ZN(
        n19408) );
  OAI22_X2 U22413 ( .A1(n19406), .A2(n19424), .B1(n21192), .B2(n19422), .ZN(
        n19893) );
  AOI22_X1 U22414 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n19426), .B1(
        n19454), .B2(n19893), .ZN(n19407) );
  OAI211_X1 U22415 ( .C1(n19429), .C2(n19837), .A(n19408), .B(n19407), .ZN(
        P2_U3053) );
  NAND2_X1 U22416 ( .A1(n19409), .A2(n19861), .ZN(n19841) );
  NOR2_X2 U22417 ( .A1(n10679), .A2(n19412), .ZN(n19897) );
  AOI22_X1 U22418 ( .A1(n19908), .A2(n19838), .B1(n19897), .B2(n19421), .ZN(
        n19416) );
  OAI22_X2 U22419 ( .A1(n19414), .A2(n19424), .B1(n19413), .B2(n19422), .ZN(
        n19899) );
  AOI22_X1 U22420 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n19426), .B1(
        n19454), .B2(n19899), .ZN(n19415) );
  OAI211_X1 U22421 ( .C1(n19429), .C2(n19841), .A(n19416), .B(n19415), .ZN(
        P2_U3054) );
  NOR2_X2 U22422 ( .A1(n19417), .A2(n19610), .ZN(n19905) );
  INV_X1 U22423 ( .A(n19905), .ZN(n19849) );
  AOI22_X1 U22424 ( .A1(n19908), .A2(n19843), .B1(n19904), .B2(n19421), .ZN(
        n19428) );
  OAI22_X2 U22425 ( .A1(n19425), .A2(n19424), .B1(n19423), .B2(n19422), .ZN(
        n19907) );
  AOI22_X1 U22426 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n19426), .B1(
        n19454), .B2(n19907), .ZN(n19427) );
  OAI211_X1 U22427 ( .C1(n19429), .C2(n19849), .A(n19428), .B(n19427), .ZN(
        P2_U3055) );
  INV_X1 U22428 ( .A(n19863), .ZN(n19728) );
  NAND2_X1 U22429 ( .A1(n19458), .A2(n20033), .ZN(n19432) );
  NOR2_X1 U22430 ( .A1(n20043), .A2(n19432), .ZN(n19452) );
  OAI21_X1 U22431 ( .B1(n19433), .B2(n19452), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19430) );
  OAI21_X1 U22432 ( .B1(n19432), .B2(n20002), .A(n19430), .ZN(n19453) );
  AOI22_X1 U22433 ( .A1(n19453), .A2(n19856), .B1(n19855), .B2(n19452), .ZN(
        n19439) );
  NAND2_X1 U22434 ( .A1(n19431), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n20003) );
  OAI21_X1 U22435 ( .B1(n20003), .B2(n19667), .A(n19432), .ZN(n19437) );
  INV_X1 U22436 ( .A(n19433), .ZN(n19435) );
  INV_X1 U22437 ( .A(n19452), .ZN(n19434) );
  OAI211_X1 U22438 ( .C1(n19435), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n20002), 
        .B(n19434), .ZN(n19436) );
  NAND3_X1 U22439 ( .A1(n19437), .A2(n19861), .A3(n19436), .ZN(n19455) );
  AOI22_X1 U22440 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19455), .B1(
        n19454), .B2(n19808), .ZN(n19438) );
  OAI211_X1 U22441 ( .C1(n19728), .C2(n19462), .A(n19439), .B(n19438), .ZN(
        P2_U3056) );
  INV_X1 U22442 ( .A(n19869), .ZN(n19731) );
  AOI22_X1 U22443 ( .A1(n19453), .A2(n19868), .B1(n19867), .B2(n19452), .ZN(
        n19441) );
  AOI22_X1 U22444 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19455), .B1(
        n19454), .B2(n19818), .ZN(n19440) );
  OAI211_X1 U22445 ( .C1(n19731), .C2(n19462), .A(n19441), .B(n19440), .ZN(
        P2_U3057) );
  AOI22_X1 U22446 ( .A1(n19453), .A2(n19874), .B1(n9966), .B2(n19452), .ZN(
        n19443) );
  AOI22_X1 U22447 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19455), .B1(
        n19454), .B2(n19822), .ZN(n19442) );
  OAI211_X1 U22448 ( .C1(n19755), .C2(n19462), .A(n19443), .B(n19442), .ZN(
        P2_U3058) );
  INV_X1 U22449 ( .A(n19881), .ZN(n19736) );
  AOI22_X1 U22450 ( .A1(n19453), .A2(n19880), .B1(n19879), .B2(n19452), .ZN(
        n19445) );
  AOI22_X1 U22451 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19455), .B1(
        n19454), .B2(n19826), .ZN(n19444) );
  OAI211_X1 U22452 ( .C1(n19736), .C2(n19462), .A(n19445), .B(n19444), .ZN(
        P2_U3059) );
  INV_X1 U22453 ( .A(n19887), .ZN(n19479) );
  AOI22_X1 U22454 ( .A1(n19453), .A2(n19886), .B1(n19885), .B2(n19452), .ZN(
        n19447) );
  AOI22_X1 U22455 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19455), .B1(
        n19454), .B2(n19830), .ZN(n19446) );
  OAI211_X1 U22456 ( .C1(n19479), .C2(n19462), .A(n19447), .B(n19446), .ZN(
        P2_U3060) );
  INV_X1 U22457 ( .A(n19893), .ZN(n19482) );
  AOI22_X1 U22458 ( .A1(n19453), .A2(n19892), .B1(n19891), .B2(n19452), .ZN(
        n19449) );
  AOI22_X1 U22459 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19455), .B1(
        n19454), .B2(n19834), .ZN(n19448) );
  OAI211_X1 U22460 ( .C1(n19482), .C2(n19462), .A(n19449), .B(n19448), .ZN(
        P2_U3061) );
  AOI22_X1 U22461 ( .A1(n19453), .A2(n19898), .B1(n19897), .B2(n19452), .ZN(
        n19451) );
  AOI22_X1 U22462 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19455), .B1(
        n19454), .B2(n19838), .ZN(n19450) );
  OAI211_X1 U22463 ( .C1(n19766), .C2(n19462), .A(n19451), .B(n19450), .ZN(
        P2_U3062) );
  INV_X1 U22464 ( .A(n19907), .ZN(n19773) );
  AOI22_X1 U22465 ( .A1(n19453), .A2(n19905), .B1(n19904), .B2(n19452), .ZN(
        n19457) );
  AOI22_X1 U22466 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19455), .B1(
        n19454), .B2(n19843), .ZN(n19456) );
  OAI211_X1 U22467 ( .C1(n19773), .C2(n19462), .A(n19457), .B(n19456), .ZN(
        P2_U3063) );
  INV_X1 U22468 ( .A(n19458), .ZN(n19491) );
  NOR2_X1 U22469 ( .A1(n20033), .A2(n19491), .ZN(n19495) );
  INV_X1 U22470 ( .A(n19495), .ZN(n19497) );
  NOR2_X1 U22471 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19497), .ZN(
        n19485) );
  OAI21_X1 U22472 ( .B1(n19461), .B2(n19485), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19460) );
  NOR2_X1 U22473 ( .A1(n19491), .A2(n19579), .ZN(n19463) );
  INV_X1 U22474 ( .A(n19463), .ZN(n19459) );
  NAND2_X1 U22475 ( .A1(n19460), .A2(n19459), .ZN(n19486) );
  AOI22_X1 U22476 ( .A1(n19486), .A2(n19856), .B1(n19855), .B2(n19485), .ZN(
        n19470) );
  INV_X1 U22477 ( .A(n19485), .ZN(n19467) );
  OAI21_X1 U22478 ( .B1(n19461), .B2(n20034), .A(n20013), .ZN(n19466) );
  AOI21_X1 U22479 ( .B1(n19519), .B2(n19462), .A(n20061), .ZN(n19464) );
  NOR3_X1 U22480 ( .A1(n19464), .A2(n19463), .A3(n20002), .ZN(n19465) );
  AOI211_X1 U22481 ( .C1(n19467), .C2(n19466), .A(n19610), .B(n19465), .ZN(
        n19468) );
  AOI22_X1 U22482 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19488), .B1(
        n19487), .B2(n19808), .ZN(n19469) );
  OAI211_X1 U22483 ( .C1(n19728), .C2(n19519), .A(n19470), .B(n19469), .ZN(
        P2_U3064) );
  AOI22_X1 U22484 ( .A1(n19486), .A2(n19868), .B1(n19867), .B2(n19485), .ZN(
        n19472) );
  AOI22_X1 U22485 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19488), .B1(
        n19487), .B2(n19818), .ZN(n19471) );
  OAI211_X1 U22486 ( .C1(n19731), .C2(n19519), .A(n19472), .B(n19471), .ZN(
        P2_U3065) );
  AOI22_X1 U22487 ( .A1(n19486), .A2(n19874), .B1(n9966), .B2(n19485), .ZN(
        n19474) );
  AOI22_X1 U22488 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19488), .B1(
        n19487), .B2(n19822), .ZN(n19473) );
  OAI211_X1 U22489 ( .C1(n19755), .C2(n19519), .A(n19474), .B(n19473), .ZN(
        P2_U3066) );
  AOI22_X1 U22490 ( .A1(n19486), .A2(n19880), .B1(n19879), .B2(n19485), .ZN(
        n19476) );
  AOI22_X1 U22491 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19488), .B1(
        n19487), .B2(n19826), .ZN(n19475) );
  OAI211_X1 U22492 ( .C1(n19736), .C2(n19519), .A(n19476), .B(n19475), .ZN(
        P2_U3067) );
  AOI22_X1 U22493 ( .A1(n19486), .A2(n19886), .B1(n19885), .B2(n19485), .ZN(
        n19478) );
  AOI22_X1 U22494 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19488), .B1(
        n19487), .B2(n19830), .ZN(n19477) );
  OAI211_X1 U22495 ( .C1(n19479), .C2(n19519), .A(n19478), .B(n19477), .ZN(
        P2_U3068) );
  AOI22_X1 U22496 ( .A1(n19486), .A2(n19892), .B1(n19891), .B2(n19485), .ZN(
        n19481) );
  AOI22_X1 U22497 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19488), .B1(
        n19487), .B2(n19834), .ZN(n19480) );
  OAI211_X1 U22498 ( .C1(n19482), .C2(n19519), .A(n19481), .B(n19480), .ZN(
        P2_U3069) );
  AOI22_X1 U22499 ( .A1(n19486), .A2(n19898), .B1(n19897), .B2(n19485), .ZN(
        n19484) );
  AOI22_X1 U22500 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19488), .B1(
        n19487), .B2(n19838), .ZN(n19483) );
  OAI211_X1 U22501 ( .C1(n19766), .C2(n19519), .A(n19484), .B(n19483), .ZN(
        P2_U3070) );
  AOI22_X1 U22502 ( .A1(n19486), .A2(n19905), .B1(n19904), .B2(n19485), .ZN(
        n19490) );
  AOI22_X1 U22503 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19488), .B1(
        n19487), .B2(n19843), .ZN(n19489) );
  OAI211_X1 U22504 ( .C1(n19773), .C2(n19519), .A(n19490), .B(n19489), .ZN(
        P2_U3071) );
  INV_X1 U22505 ( .A(n19808), .ZN(n19866) );
  NOR2_X1 U22506 ( .A1(n19491), .A2(n19716), .ZN(n19514) );
  AOI22_X1 U22507 ( .A1(n19535), .A2(n19863), .B1(n19855), .B2(n19514), .ZN(
        n19500) );
  OAI21_X1 U22508 ( .B1(n20003), .B2(n20004), .A(n20006), .ZN(n19498) );
  INV_X1 U22509 ( .A(n11208), .ZN(n19493) );
  INV_X1 U22510 ( .A(n19514), .ZN(n19492) );
  OAI211_X1 U22511 ( .C1(n19493), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n20002), 
        .B(n19492), .ZN(n19494) );
  OAI211_X1 U22512 ( .C1(n19498), .C2(n19495), .A(n19861), .B(n19494), .ZN(
        n19516) );
  OAI21_X1 U22513 ( .B1(n11208), .B2(n19514), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19496) );
  AOI22_X1 U22514 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19516), .B1(
        n19856), .B2(n19515), .ZN(n19499) );
  OAI211_X1 U22515 ( .C1(n19866), .C2(n19519), .A(n19500), .B(n19499), .ZN(
        P2_U3072) );
  INV_X1 U22516 ( .A(n19818), .ZN(n19872) );
  AOI22_X1 U22517 ( .A1(n19535), .A2(n19869), .B1(n19867), .B2(n19514), .ZN(
        n19502) );
  AOI22_X1 U22518 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19516), .B1(
        n19868), .B2(n19515), .ZN(n19501) );
  OAI211_X1 U22519 ( .C1(n19872), .C2(n19519), .A(n19502), .B(n19501), .ZN(
        P2_U3073) );
  INV_X1 U22520 ( .A(n19822), .ZN(n19878) );
  AOI22_X1 U22521 ( .A1(n19535), .A2(n19875), .B1(n19514), .B2(n9966), .ZN(
        n19504) );
  AOI22_X1 U22522 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19516), .B1(
        n19874), .B2(n19515), .ZN(n19503) );
  OAI211_X1 U22523 ( .C1(n19878), .C2(n19519), .A(n19504), .B(n19503), .ZN(
        P2_U3074) );
  AOI22_X1 U22524 ( .A1(n19535), .A2(n19881), .B1(n19514), .B2(n19879), .ZN(
        n19506) );
  AOI22_X1 U22525 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19516), .B1(
        n19880), .B2(n19515), .ZN(n19505) );
  OAI211_X1 U22526 ( .C1(n19884), .C2(n19519), .A(n19506), .B(n19505), .ZN(
        P2_U3075) );
  AOI22_X1 U22527 ( .A1(n19535), .A2(n19887), .B1(n19514), .B2(n19885), .ZN(
        n19508) );
  AOI22_X1 U22528 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19516), .B1(
        n19886), .B2(n19515), .ZN(n19507) );
  OAI211_X1 U22529 ( .C1(n19890), .C2(n19519), .A(n19508), .B(n19507), .ZN(
        P2_U3076) );
  AOI22_X1 U22530 ( .A1(n19535), .A2(n19893), .B1(n19514), .B2(n19891), .ZN(
        n19510) );
  AOI22_X1 U22531 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19516), .B1(
        n19892), .B2(n19515), .ZN(n19509) );
  OAI211_X1 U22532 ( .C1(n19896), .C2(n19519), .A(n19510), .B(n19509), .ZN(
        P2_U3077) );
  INV_X1 U22533 ( .A(n19519), .ZN(n19511) );
  AOI22_X1 U22534 ( .A1(n19511), .A2(n19838), .B1(n19514), .B2(n19897), .ZN(
        n19513) );
  AOI22_X1 U22535 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19516), .B1(
        n19898), .B2(n19515), .ZN(n19512) );
  OAI211_X1 U22536 ( .C1(n19766), .C2(n19530), .A(n19513), .B(n19512), .ZN(
        P2_U3078) );
  INV_X1 U22537 ( .A(n19843), .ZN(n19913) );
  AOI22_X1 U22538 ( .A1(n19535), .A2(n19907), .B1(n19514), .B2(n19904), .ZN(
        n19518) );
  AOI22_X1 U22539 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19516), .B1(
        n19905), .B2(n19515), .ZN(n19517) );
  OAI211_X1 U22540 ( .C1(n19913), .C2(n19519), .A(n19518), .B(n19517), .ZN(
        P2_U3079) );
  INV_X1 U22541 ( .A(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n19522) );
  AOI22_X1 U22542 ( .A1(n19534), .A2(n19874), .B1(n9966), .B2(n19533), .ZN(
        n19521) );
  AOI22_X1 U22543 ( .A1(n19535), .A2(n19822), .B1(n19563), .B2(n19875), .ZN(
        n19520) );
  OAI211_X1 U22544 ( .C1(n19523), .C2(n19522), .A(n19521), .B(n19520), .ZN(
        P2_U3082) );
  AOI22_X1 U22545 ( .A1(n19534), .A2(n19880), .B1(n19879), .B2(n19533), .ZN(
        n19525) );
  AOI22_X1 U22546 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19536), .B1(
        n19563), .B2(n19881), .ZN(n19524) );
  OAI211_X1 U22547 ( .C1(n19884), .C2(n19530), .A(n19525), .B(n19524), .ZN(
        P2_U3083) );
  AOI22_X1 U22548 ( .A1(n19534), .A2(n19886), .B1(n19885), .B2(n19533), .ZN(
        n19527) );
  AOI22_X1 U22549 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19536), .B1(
        n19563), .B2(n19887), .ZN(n19526) );
  OAI211_X1 U22550 ( .C1(n19890), .C2(n19530), .A(n19527), .B(n19526), .ZN(
        P2_U3084) );
  AOI22_X1 U22551 ( .A1(n19534), .A2(n19892), .B1(n19891), .B2(n19533), .ZN(
        n19529) );
  AOI22_X1 U22552 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19536), .B1(
        n19563), .B2(n19893), .ZN(n19528) );
  OAI211_X1 U22553 ( .C1(n19896), .C2(n19530), .A(n19529), .B(n19528), .ZN(
        P2_U3085) );
  AOI22_X1 U22554 ( .A1(n19534), .A2(n19898), .B1(n19897), .B2(n19533), .ZN(
        n19532) );
  AOI22_X1 U22555 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19536), .B1(
        n19535), .B2(n19838), .ZN(n19531) );
  OAI211_X1 U22556 ( .C1(n19766), .C2(n19561), .A(n19532), .B(n19531), .ZN(
        P2_U3086) );
  AOI22_X1 U22557 ( .A1(n19534), .A2(n19905), .B1(n19904), .B2(n19533), .ZN(
        n19538) );
  AOI22_X1 U22558 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19536), .B1(
        n19535), .B2(n19843), .ZN(n19537) );
  OAI211_X1 U22559 ( .C1(n19773), .C2(n19561), .A(n19538), .B(n19537), .ZN(
        P2_U3087) );
  NOR3_X2 U22560 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20043), .A3(
        n19539), .ZN(n19562) );
  AOI22_X1 U22561 ( .A1(n19563), .A2(n19808), .B1(n19855), .B2(n19562), .ZN(
        n19548) );
  OAI21_X1 U22562 ( .B1(n20003), .B2(n19781), .A(n20006), .ZN(n19546) );
  NAND2_X1 U22563 ( .A1(n20033), .A2(n13583), .ZN(n19545) );
  INV_X1 U22564 ( .A(n19545), .ZN(n19543) );
  OAI21_X1 U22565 ( .B1(n11207), .B2(n20034), .A(n20036), .ZN(n19541) );
  INV_X1 U22566 ( .A(n19562), .ZN(n19540) );
  AOI21_X1 U22567 ( .B1(n19541), .B2(n19540), .A(n19610), .ZN(n19542) );
  OAI21_X1 U22568 ( .B1(n11207), .B2(n19562), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19544) );
  AOI22_X1 U22569 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n19565), .B1(
        n19856), .B2(n19564), .ZN(n19547) );
  OAI211_X1 U22570 ( .C1(n19728), .C2(n19603), .A(n19548), .B(n19547), .ZN(
        P2_U3088) );
  AOI22_X1 U22571 ( .A1(n19563), .A2(n19818), .B1(n19867), .B2(n19562), .ZN(
        n19550) );
  AOI22_X1 U22572 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19565), .B1(
        n19868), .B2(n19564), .ZN(n19549) );
  OAI211_X1 U22573 ( .C1(n19731), .C2(n19603), .A(n19550), .B(n19549), .ZN(
        P2_U3089) );
  AOI22_X1 U22574 ( .A1(n19563), .A2(n19822), .B1(n19562), .B2(n9966), .ZN(
        n19552) );
  AOI22_X1 U22575 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19565), .B1(
        n19874), .B2(n19564), .ZN(n19551) );
  OAI211_X1 U22576 ( .C1(n19755), .C2(n19603), .A(n19552), .B(n19551), .ZN(
        P2_U3090) );
  AOI22_X1 U22577 ( .A1(n19583), .A2(n19881), .B1(n19879), .B2(n19562), .ZN(
        n19554) );
  AOI22_X1 U22578 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19565), .B1(
        n19880), .B2(n19564), .ZN(n19553) );
  OAI211_X1 U22579 ( .C1(n19884), .C2(n19561), .A(n19554), .B(n19553), .ZN(
        P2_U3091) );
  AOI22_X1 U22580 ( .A1(n19583), .A2(n19887), .B1(n19562), .B2(n19885), .ZN(
        n19556) );
  AOI22_X1 U22581 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19565), .B1(
        n19886), .B2(n19564), .ZN(n19555) );
  OAI211_X1 U22582 ( .C1(n19890), .C2(n19561), .A(n19556), .B(n19555), .ZN(
        P2_U3092) );
  AOI22_X1 U22583 ( .A1(n19583), .A2(n19893), .B1(n19562), .B2(n19891), .ZN(
        n19558) );
  AOI22_X1 U22584 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19565), .B1(
        n19892), .B2(n19564), .ZN(n19557) );
  OAI211_X1 U22585 ( .C1(n19896), .C2(n19561), .A(n19558), .B(n19557), .ZN(
        P2_U3093) );
  INV_X1 U22586 ( .A(n19838), .ZN(n19902) );
  AOI22_X1 U22587 ( .A1(n19583), .A2(n19899), .B1(n19562), .B2(n19897), .ZN(
        n19560) );
  AOI22_X1 U22588 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19565), .B1(
        n19898), .B2(n19564), .ZN(n19559) );
  OAI211_X1 U22589 ( .C1(n19902), .C2(n19561), .A(n19560), .B(n19559), .ZN(
        P2_U3094) );
  AOI22_X1 U22590 ( .A1(n19563), .A2(n19843), .B1(n19562), .B2(n19904), .ZN(
        n19567) );
  AOI22_X1 U22591 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19565), .B1(
        n19905), .B2(n19564), .ZN(n19566) );
  OAI211_X1 U22592 ( .C1(n19773), .C2(n19603), .A(n19567), .B(n19566), .ZN(
        P2_U3095) );
  OAI21_X1 U22593 ( .B1(n19583), .B2(n19604), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19571) );
  NAND2_X1 U22594 ( .A1(n19569), .A2(n13583), .ZN(n19570) );
  NAND2_X1 U22595 ( .A1(n19571), .A2(n19570), .ZN(n19577) );
  NAND2_X1 U22596 ( .A1(n19572), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n19573) );
  NAND2_X1 U22597 ( .A1(n19573), .A2(n20036), .ZN(n19575) );
  NAND2_X1 U22598 ( .A1(n19853), .A2(n20017), .ZN(n19612) );
  NOR2_X1 U22599 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19612), .ZN(
        n19598) );
  INV_X1 U22600 ( .A(n19598), .ZN(n19574) );
  AOI21_X1 U22601 ( .B1(n19575), .B2(n19574), .A(n19610), .ZN(n19576) );
  OAI21_X1 U22602 ( .B1(n11224), .B2(n19598), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19578) );
  AOI22_X1 U22603 ( .A1(n19599), .A2(n19856), .B1(n19855), .B2(n19598), .ZN(
        n19581) );
  AOI22_X1 U22604 ( .A1(n19604), .A2(n19863), .B1(n19583), .B2(n19808), .ZN(
        n19580) );
  OAI211_X1 U22605 ( .C1(n19587), .C2(n19582), .A(n19581), .B(n19580), .ZN(
        P2_U3096) );
  AOI22_X1 U22606 ( .A1(n19599), .A2(n19868), .B1(n19867), .B2(n19598), .ZN(
        n19585) );
  AOI22_X1 U22607 ( .A1(n19604), .A2(n19869), .B1(n19583), .B2(n19818), .ZN(
        n19584) );
  OAI211_X1 U22608 ( .C1(n19587), .C2(n19586), .A(n19585), .B(n19584), .ZN(
        P2_U3097) );
  AOI22_X1 U22609 ( .A1(n19599), .A2(n19874), .B1(n9966), .B2(n19598), .ZN(
        n19589) );
  AOI22_X1 U22610 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19600), .B1(
        n19604), .B2(n19875), .ZN(n19588) );
  OAI211_X1 U22611 ( .C1(n19878), .C2(n19603), .A(n19589), .B(n19588), .ZN(
        P2_U3098) );
  AOI22_X1 U22612 ( .A1(n19599), .A2(n19880), .B1(n19879), .B2(n19598), .ZN(
        n19591) );
  AOI22_X1 U22613 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19600), .B1(
        n19604), .B2(n19881), .ZN(n19590) );
  OAI211_X1 U22614 ( .C1(n19884), .C2(n19603), .A(n19591), .B(n19590), .ZN(
        P2_U3099) );
  AOI22_X1 U22615 ( .A1(n19599), .A2(n19886), .B1(n19885), .B2(n19598), .ZN(
        n19593) );
  AOI22_X1 U22616 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19600), .B1(
        n19604), .B2(n19887), .ZN(n19592) );
  OAI211_X1 U22617 ( .C1(n19890), .C2(n19603), .A(n19593), .B(n19592), .ZN(
        P2_U3100) );
  AOI22_X1 U22618 ( .A1(n19599), .A2(n19892), .B1(n19891), .B2(n19598), .ZN(
        n19595) );
  AOI22_X1 U22619 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19600), .B1(
        n19604), .B2(n19893), .ZN(n19594) );
  OAI211_X1 U22620 ( .C1(n19896), .C2(n19603), .A(n19595), .B(n19594), .ZN(
        P2_U3101) );
  AOI22_X1 U22621 ( .A1(n19599), .A2(n19898), .B1(n19897), .B2(n19598), .ZN(
        n19597) );
  AOI22_X1 U22622 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19600), .B1(
        n19604), .B2(n19899), .ZN(n19596) );
  OAI211_X1 U22623 ( .C1(n19902), .C2(n19603), .A(n19597), .B(n19596), .ZN(
        P2_U3102) );
  AOI22_X1 U22624 ( .A1(n19599), .A2(n19905), .B1(n19904), .B2(n19598), .ZN(
        n19602) );
  AOI22_X1 U22625 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19600), .B1(
        n19604), .B2(n19907), .ZN(n19601) );
  OAI211_X1 U22626 ( .C1(n19913), .C2(n19603), .A(n19602), .B(n19601), .ZN(
        P2_U3103) );
  NOR3_X1 U22627 ( .A1(n19605), .A2(n19643), .A3(n20034), .ZN(n19611) );
  INV_X1 U22628 ( .A(n19612), .ZN(n19606) );
  AOI21_X1 U22629 ( .B1(n20013), .B2(n19606), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19607) );
  NOR2_X1 U22630 ( .A1(n19611), .A2(n19607), .ZN(n19630) );
  AOI22_X1 U22631 ( .A1(n19630), .A2(n19856), .B1(n19643), .B2(n19855), .ZN(
        n19617) );
  INV_X1 U22632 ( .A(n20003), .ZN(n19609) );
  INV_X1 U22633 ( .A(n20001), .ZN(n19608) );
  NAND2_X1 U22634 ( .A1(n19609), .A2(n19608), .ZN(n19613) );
  AOI211_X1 U22635 ( .C1(n19613), .C2(n19612), .A(n19611), .B(n19610), .ZN(
        n19614) );
  AOI22_X1 U22636 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n19631), .B1(
        n19662), .B2(n19863), .ZN(n19616) );
  OAI211_X1 U22637 ( .C1(n19866), .C2(n19634), .A(n19617), .B(n19616), .ZN(
        P2_U3104) );
  AOI22_X1 U22638 ( .A1(n19630), .A2(n19868), .B1(n19643), .B2(n19867), .ZN(
        n19619) );
  AOI22_X1 U22639 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19631), .B1(
        n19662), .B2(n19869), .ZN(n19618) );
  OAI211_X1 U22640 ( .C1(n19872), .C2(n19634), .A(n19619), .B(n19618), .ZN(
        P2_U3105) );
  AOI22_X1 U22641 ( .A1(n19630), .A2(n19874), .B1(n19643), .B2(n9966), .ZN(
        n19621) );
  AOI22_X1 U22642 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19631), .B1(
        n19662), .B2(n19875), .ZN(n19620) );
  OAI211_X1 U22643 ( .C1(n19878), .C2(n19634), .A(n19621), .B(n19620), .ZN(
        P2_U3106) );
  AOI22_X1 U22644 ( .A1(n19630), .A2(n19880), .B1(n19643), .B2(n19879), .ZN(
        n19623) );
  AOI22_X1 U22645 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19631), .B1(
        n19662), .B2(n19881), .ZN(n19622) );
  OAI211_X1 U22646 ( .C1(n19884), .C2(n19634), .A(n19623), .B(n19622), .ZN(
        P2_U3107) );
  AOI22_X1 U22647 ( .A1(n19630), .A2(n19886), .B1(n19643), .B2(n19885), .ZN(
        n19625) );
  AOI22_X1 U22648 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19631), .B1(
        n19662), .B2(n19887), .ZN(n19624) );
  OAI211_X1 U22649 ( .C1(n19890), .C2(n19634), .A(n19625), .B(n19624), .ZN(
        P2_U3108) );
  AOI22_X1 U22650 ( .A1(n19630), .A2(n19892), .B1(n19643), .B2(n19891), .ZN(
        n19627) );
  AOI22_X1 U22651 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19631), .B1(
        n19662), .B2(n19893), .ZN(n19626) );
  OAI211_X1 U22652 ( .C1(n19896), .C2(n19634), .A(n19627), .B(n19626), .ZN(
        P2_U3109) );
  AOI22_X1 U22653 ( .A1(n19630), .A2(n19898), .B1(n19643), .B2(n19897), .ZN(
        n19629) );
  AOI22_X1 U22654 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19631), .B1(
        n19662), .B2(n19899), .ZN(n19628) );
  OAI211_X1 U22655 ( .C1(n19902), .C2(n19634), .A(n19629), .B(n19628), .ZN(
        P2_U3110) );
  AOI22_X1 U22656 ( .A1(n19630), .A2(n19905), .B1(n19643), .B2(n19904), .ZN(
        n19633) );
  AOI22_X1 U22657 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19631), .B1(
        n19662), .B2(n19907), .ZN(n19632) );
  OAI211_X1 U22658 ( .C1(n19913), .C2(n19634), .A(n19633), .B(n19632), .ZN(
        P2_U3111) );
  NOR3_X1 U22659 ( .A1(n19680), .A2(n19662), .A3(n20002), .ZN(n19636) );
  NOR2_X1 U22660 ( .A1(n19636), .A2(n19635), .ZN(n19644) );
  INV_X1 U22661 ( .A(n19644), .ZN(n19642) );
  INV_X1 U22662 ( .A(n19643), .ZN(n19640) );
  NOR2_X1 U22663 ( .A1(n19637), .A2(n19717), .ZN(n19661) );
  INV_X1 U22664 ( .A(n19661), .ZN(n19639) );
  NAND2_X1 U22665 ( .A1(n11216), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n19638) );
  OAI211_X1 U22666 ( .C1(n19644), .C2(n19640), .A(n19639), .B(n19638), .ZN(
        n19641) );
  AOI22_X1 U22667 ( .A1(n19680), .A2(n19863), .B1(n19855), .B2(n19661), .ZN(
        n19648) );
  NOR2_X1 U22668 ( .A1(n19644), .A2(n19643), .ZN(n19645) );
  AOI211_X1 U22669 ( .C1(P2_STATE2_REG_2__SCAN_IN), .C2(n11238), .A(
        P2_STATE2_REG_3__SCAN_IN), .B(n19645), .ZN(n19646) );
  AOI22_X1 U22670 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19663), .B1(
        n19662), .B2(n19808), .ZN(n19647) );
  OAI211_X1 U22671 ( .C1(n19817), .C2(n19666), .A(n19648), .B(n19647), .ZN(
        P2_U3112) );
  AOI22_X1 U22672 ( .A1(n19680), .A2(n19869), .B1(n19867), .B2(n19661), .ZN(
        n19650) );
  AOI22_X1 U22673 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19663), .B1(
        n19662), .B2(n19818), .ZN(n19649) );
  OAI211_X1 U22674 ( .C1(n19666), .C2(n19821), .A(n19650), .B(n19649), .ZN(
        P2_U3113) );
  AOI22_X1 U22675 ( .A1(n19662), .A2(n19822), .B1(n9966), .B2(n19661), .ZN(
        n19652) );
  AOI22_X1 U22676 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19663), .B1(
        n19680), .B2(n19875), .ZN(n19651) );
  OAI211_X1 U22677 ( .C1(n19666), .C2(n19825), .A(n19652), .B(n19651), .ZN(
        P2_U3114) );
  AOI22_X1 U22678 ( .A1(n19680), .A2(n19881), .B1(n19879), .B2(n19661), .ZN(
        n19654) );
  AOI22_X1 U22679 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19663), .B1(
        n19662), .B2(n19826), .ZN(n19653) );
  OAI211_X1 U22680 ( .C1(n19666), .C2(n19829), .A(n19654), .B(n19653), .ZN(
        P2_U3115) );
  AOI22_X1 U22681 ( .A1(n19662), .A2(n19830), .B1(n19885), .B2(n19661), .ZN(
        n19656) );
  AOI22_X1 U22682 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19663), .B1(
        n19680), .B2(n19887), .ZN(n19655) );
  OAI211_X1 U22683 ( .C1(n19666), .C2(n19833), .A(n19656), .B(n19655), .ZN(
        P2_U3116) );
  AOI22_X1 U22684 ( .A1(n19680), .A2(n19893), .B1(n19891), .B2(n19661), .ZN(
        n19658) );
  AOI22_X1 U22685 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19663), .B1(
        n19662), .B2(n19834), .ZN(n19657) );
  OAI211_X1 U22686 ( .C1(n19666), .C2(n19837), .A(n19658), .B(n19657), .ZN(
        P2_U3117) );
  AOI22_X1 U22687 ( .A1(n19662), .A2(n19838), .B1(n19897), .B2(n19661), .ZN(
        n19660) );
  AOI22_X1 U22688 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19663), .B1(
        n19680), .B2(n19899), .ZN(n19659) );
  OAI211_X1 U22689 ( .C1(n19666), .C2(n19841), .A(n19660), .B(n19659), .ZN(
        P2_U3118) );
  AOI22_X1 U22690 ( .A1(n19680), .A2(n19907), .B1(n19904), .B2(n19661), .ZN(
        n19665) );
  AOI22_X1 U22691 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19663), .B1(
        n19662), .B2(n19843), .ZN(n19664) );
  OAI211_X1 U22692 ( .C1(n19666), .C2(n19849), .A(n19665), .B(n19664), .ZN(
        P2_U3119) );
  AOI22_X1 U22693 ( .A1(n19680), .A2(n19808), .B1(n19855), .B2(n19692), .ZN(
        n19677) );
  NAND2_X1 U22694 ( .A1(n20010), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19858) );
  OAI21_X1 U22695 ( .B1(n19858), .B2(n19667), .A(n20006), .ZN(n19675) );
  NAND2_X1 U22696 ( .A1(n20033), .A2(n19720), .ZN(n19674) );
  INV_X1 U22697 ( .A(n19674), .ZN(n19671) );
  INV_X1 U22698 ( .A(n19672), .ZN(n19669) );
  INV_X1 U22699 ( .A(n19692), .ZN(n19668) );
  OAI211_X1 U22700 ( .C1(n19669), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n20002), 
        .B(n19668), .ZN(n19670) );
  OAI211_X1 U22701 ( .C1(n19675), .C2(n19671), .A(n19861), .B(n19670), .ZN(
        n19694) );
  OAI21_X1 U22702 ( .B1(n19672), .B2(n19692), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19673) );
  AOI22_X1 U22703 ( .A1(P2_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n19694), .B1(
        n19856), .B2(n19693), .ZN(n19676) );
  OAI211_X1 U22704 ( .C1(n19728), .C2(n19683), .A(n19677), .B(n19676), .ZN(
        P2_U3120) );
  AOI22_X1 U22705 ( .A1(n19710), .A2(n19869), .B1(n19867), .B2(n19692), .ZN(
        n19679) );
  AOI22_X1 U22706 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19694), .B1(
        n19868), .B2(n19693), .ZN(n19678) );
  OAI211_X1 U22707 ( .C1(n19872), .C2(n19697), .A(n19679), .B(n19678), .ZN(
        P2_U3121) );
  AOI22_X1 U22708 ( .A1(n19680), .A2(n19822), .B1(n9966), .B2(n19692), .ZN(
        n19682) );
  AOI22_X1 U22709 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19694), .B1(
        n19874), .B2(n19693), .ZN(n19681) );
  OAI211_X1 U22710 ( .C1(n19755), .C2(n19683), .A(n19682), .B(n19681), .ZN(
        P2_U3122) );
  AOI22_X1 U22711 ( .A1(n19710), .A2(n19881), .B1(n19879), .B2(n19692), .ZN(
        n19685) );
  AOI22_X1 U22712 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19694), .B1(
        n19880), .B2(n19693), .ZN(n19684) );
  OAI211_X1 U22713 ( .C1(n19884), .C2(n19697), .A(n19685), .B(n19684), .ZN(
        P2_U3123) );
  AOI22_X1 U22714 ( .A1(n19710), .A2(n19887), .B1(n19885), .B2(n19692), .ZN(
        n19687) );
  AOI22_X1 U22715 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19694), .B1(
        n19886), .B2(n19693), .ZN(n19686) );
  OAI211_X1 U22716 ( .C1(n19890), .C2(n19697), .A(n19687), .B(n19686), .ZN(
        P2_U3124) );
  AOI22_X1 U22717 ( .A1(n19710), .A2(n19893), .B1(n19891), .B2(n19692), .ZN(
        n19689) );
  AOI22_X1 U22718 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19694), .B1(
        n19892), .B2(n19693), .ZN(n19688) );
  OAI211_X1 U22719 ( .C1(n19896), .C2(n19697), .A(n19689), .B(n19688), .ZN(
        P2_U3125) );
  AOI22_X1 U22720 ( .A1(n19710), .A2(n19899), .B1(n19897), .B2(n19692), .ZN(
        n19691) );
  AOI22_X1 U22721 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19694), .B1(
        n19898), .B2(n19693), .ZN(n19690) );
  OAI211_X1 U22722 ( .C1(n19902), .C2(n19697), .A(n19691), .B(n19690), .ZN(
        P2_U3126) );
  AOI22_X1 U22723 ( .A1(n19710), .A2(n19907), .B1(n19904), .B2(n19692), .ZN(
        n19696) );
  AOI22_X1 U22724 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19694), .B1(
        n19905), .B2(n19693), .ZN(n19695) );
  OAI211_X1 U22725 ( .C1(n19913), .C2(n19697), .A(n19696), .B(n19695), .ZN(
        P2_U3127) );
  AOI22_X1 U22726 ( .A1(n19709), .A2(n19874), .B1(n19708), .B2(n9966), .ZN(
        n19699) );
  AOI22_X1 U22727 ( .A1(n19710), .A2(n19822), .B1(n19737), .B2(n19875), .ZN(
        n19698) );
  OAI211_X1 U22728 ( .C1(n19714), .C2(n10769), .A(n19699), .B(n19698), .ZN(
        P2_U3130) );
  AOI22_X1 U22729 ( .A1(n19709), .A2(n19880), .B1(n19708), .B2(n19879), .ZN(
        n19701) );
  AOI22_X1 U22730 ( .A1(n19737), .A2(n19881), .B1(n19710), .B2(n19826), .ZN(
        n19700) );
  OAI211_X1 U22731 ( .C1(n19714), .C2(n21213), .A(n19701), .B(n19700), .ZN(
        P2_U3131) );
  AOI22_X1 U22732 ( .A1(n19709), .A2(n19886), .B1(n19708), .B2(n19885), .ZN(
        n19703) );
  AOI22_X1 U22733 ( .A1(n19710), .A2(n19830), .B1(n19737), .B2(n19887), .ZN(
        n19702) );
  OAI211_X1 U22734 ( .C1(n19714), .C2(n10805), .A(n19703), .B(n19702), .ZN(
        P2_U3132) );
  AOI22_X1 U22735 ( .A1(n19709), .A2(n19892), .B1(n19708), .B2(n19891), .ZN(
        n19705) );
  AOI22_X1 U22736 ( .A1(n19737), .A2(n19893), .B1(n19710), .B2(n19834), .ZN(
        n19704) );
  OAI211_X1 U22737 ( .C1(n19714), .C2(n10828), .A(n19705), .B(n19704), .ZN(
        P2_U3133) );
  AOI22_X1 U22738 ( .A1(n19709), .A2(n19898), .B1(n19708), .B2(n19897), .ZN(
        n19707) );
  AOI22_X1 U22739 ( .A1(n19710), .A2(n19838), .B1(n19737), .B2(n19899), .ZN(
        n19706) );
  OAI211_X1 U22740 ( .C1(n19714), .C2(n11242), .A(n19707), .B(n19706), .ZN(
        P2_U3134) );
  AOI22_X1 U22741 ( .A1(n19709), .A2(n19905), .B1(n19708), .B2(n19904), .ZN(
        n19712) );
  AOI22_X1 U22742 ( .A1(n19737), .A2(n19907), .B1(n19710), .B2(n19843), .ZN(
        n19711) );
  OAI211_X1 U22743 ( .C1(n19714), .C2(n19713), .A(n19712), .B(n19711), .ZN(
        P2_U3135) );
  INV_X1 U22744 ( .A(n19715), .ZN(n19719) );
  NOR2_X1 U22745 ( .A1(n19717), .A2(n19716), .ZN(n19744) );
  NOR2_X1 U22746 ( .A1(n19744), .A2(n20034), .ZN(n19718) );
  NAND2_X1 U22747 ( .A1(n19719), .A2(n19718), .ZN(n19723) );
  NAND2_X1 U22748 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19720), .ZN(
        n19722) );
  OAI21_X1 U22749 ( .B1(n19722), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n20034), 
        .ZN(n19721) );
  AOI22_X1 U22750 ( .A1(n19745), .A2(n19856), .B1(n19855), .B2(n19744), .ZN(
        n19727) );
  OAI21_X1 U22751 ( .B1(n19858), .B2(n20004), .A(n19722), .ZN(n19724) );
  AND2_X1 U22752 ( .A1(n19724), .A2(n19723), .ZN(n19725) );
  OAI211_X1 U22753 ( .C1(n19744), .C2(n20036), .A(n19725), .B(n19861), .ZN(
        n19746) );
  AOI22_X1 U22754 ( .A1(P2_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19746), .B1(
        n19737), .B2(n19808), .ZN(n19726) );
  OAI211_X1 U22755 ( .C1(n19728), .C2(n19763), .A(n19727), .B(n19726), .ZN(
        P2_U3136) );
  AOI22_X1 U22756 ( .A1(n19745), .A2(n19868), .B1(n19867), .B2(n19744), .ZN(
        n19730) );
  AOI22_X1 U22757 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19746), .B1(
        n19737), .B2(n19818), .ZN(n19729) );
  OAI211_X1 U22758 ( .C1(n19731), .C2(n19763), .A(n19730), .B(n19729), .ZN(
        P2_U3137) );
  AOI22_X1 U22759 ( .A1(n19745), .A2(n19874), .B1(n9966), .B2(n19744), .ZN(
        n19733) );
  AOI22_X1 U22760 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19746), .B1(
        n19737), .B2(n19822), .ZN(n19732) );
  OAI211_X1 U22761 ( .C1(n19755), .C2(n19763), .A(n19733), .B(n19732), .ZN(
        P2_U3138) );
  AOI22_X1 U22762 ( .A1(n19745), .A2(n19880), .B1(n19879), .B2(n19744), .ZN(
        n19735) );
  AOI22_X1 U22763 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19746), .B1(
        n19737), .B2(n19826), .ZN(n19734) );
  OAI211_X1 U22764 ( .C1(n19736), .C2(n19763), .A(n19735), .B(n19734), .ZN(
        P2_U3139) );
  AOI22_X1 U22765 ( .A1(n19745), .A2(n19886), .B1(n19885), .B2(n19744), .ZN(
        n19739) );
  AOI22_X1 U22766 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19746), .B1(
        n19769), .B2(n19887), .ZN(n19738) );
  OAI211_X1 U22767 ( .C1(n19890), .C2(n19749), .A(n19739), .B(n19738), .ZN(
        P2_U3140) );
  AOI22_X1 U22768 ( .A1(n19745), .A2(n19892), .B1(n19891), .B2(n19744), .ZN(
        n19741) );
  AOI22_X1 U22769 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19746), .B1(
        n19769), .B2(n19893), .ZN(n19740) );
  OAI211_X1 U22770 ( .C1(n19896), .C2(n19749), .A(n19741), .B(n19740), .ZN(
        P2_U3141) );
  AOI22_X1 U22771 ( .A1(n19745), .A2(n19898), .B1(n19897), .B2(n19744), .ZN(
        n19743) );
  AOI22_X1 U22772 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19746), .B1(
        n19769), .B2(n19899), .ZN(n19742) );
  OAI211_X1 U22773 ( .C1(n19902), .C2(n19749), .A(n19743), .B(n19742), .ZN(
        P2_U3142) );
  AOI22_X1 U22774 ( .A1(n19745), .A2(n19905), .B1(n19904), .B2(n19744), .ZN(
        n19748) );
  AOI22_X1 U22775 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19746), .B1(
        n19769), .B2(n19907), .ZN(n19747) );
  OAI211_X1 U22776 ( .C1(n19913), .C2(n19749), .A(n19748), .B(n19747), .ZN(
        P2_U3143) );
  AOI22_X1 U22777 ( .A1(n19768), .A2(n19868), .B1(n19867), .B2(n19767), .ZN(
        n19752) );
  INV_X1 U22778 ( .A(n19750), .ZN(n19770) );
  AOI22_X1 U22779 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n19770), .B1(
        n19760), .B2(n19869), .ZN(n19751) );
  OAI211_X1 U22780 ( .C1(n19872), .C2(n19763), .A(n19752), .B(n19751), .ZN(
        P2_U3145) );
  AOI22_X1 U22781 ( .A1(n19768), .A2(n19874), .B1(n19767), .B2(n9966), .ZN(
        n19754) );
  AOI22_X1 U22782 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n19770), .B1(
        n19769), .B2(n19822), .ZN(n19753) );
  OAI211_X1 U22783 ( .C1(n19755), .C2(n19801), .A(n19754), .B(n19753), .ZN(
        P2_U3146) );
  AOI22_X1 U22784 ( .A1(n19768), .A2(n19880), .B1(n19767), .B2(n19879), .ZN(
        n19757) );
  AOI22_X1 U22785 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n19770), .B1(
        n19760), .B2(n19881), .ZN(n19756) );
  OAI211_X1 U22786 ( .C1(n19884), .C2(n19763), .A(n19757), .B(n19756), .ZN(
        P2_U3147) );
  AOI22_X1 U22787 ( .A1(n19768), .A2(n19886), .B1(n19767), .B2(n19885), .ZN(
        n19759) );
  AOI22_X1 U22788 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n19770), .B1(
        n19760), .B2(n19887), .ZN(n19758) );
  OAI211_X1 U22789 ( .C1(n19890), .C2(n19763), .A(n19759), .B(n19758), .ZN(
        P2_U3148) );
  AOI22_X1 U22790 ( .A1(n19768), .A2(n19892), .B1(n19767), .B2(n19891), .ZN(
        n19762) );
  AOI22_X1 U22791 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19770), .B1(
        n19760), .B2(n19893), .ZN(n19761) );
  OAI211_X1 U22792 ( .C1(n19896), .C2(n19763), .A(n19762), .B(n19761), .ZN(
        P2_U3149) );
  AOI22_X1 U22793 ( .A1(n19768), .A2(n19898), .B1(n19767), .B2(n19897), .ZN(
        n19765) );
  AOI22_X1 U22794 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n19770), .B1(
        n19769), .B2(n19838), .ZN(n19764) );
  OAI211_X1 U22795 ( .C1(n19766), .C2(n19801), .A(n19765), .B(n19764), .ZN(
        P2_U3150) );
  AOI22_X1 U22796 ( .A1(n19768), .A2(n19905), .B1(n19767), .B2(n19904), .ZN(
        n19772) );
  AOI22_X1 U22797 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n19770), .B1(
        n19769), .B2(n19843), .ZN(n19771) );
  OAI211_X1 U22798 ( .C1(n19773), .C2(n19801), .A(n19772), .B(n19771), .ZN(
        P2_U3151) );
  NOR2_X1 U22799 ( .A1(n20043), .A2(n19779), .ZN(n19806) );
  NOR3_X1 U22800 ( .A1(n11209), .A2(n19806), .A3(n20034), .ZN(n19776) );
  INV_X1 U22801 ( .A(n19779), .ZN(n19774) );
  AOI21_X1 U22802 ( .B1(n20013), .B2(n19774), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19775) );
  AOI22_X1 U22803 ( .A1(n19797), .A2(n19856), .B1(n19855), .B2(n19806), .ZN(
        n19784) );
  INV_X1 U22804 ( .A(n19776), .ZN(n19777) );
  OAI211_X1 U22805 ( .C1(n20036), .C2(n19806), .A(n19777), .B(n19861), .ZN(
        n19778) );
  AOI221_X1 U22806 ( .B1(n19779), .B2(n19781), .C1(n19779), .C2(n19858), .A(
        n19778), .ZN(n19780) );
  AOI22_X1 U22807 ( .A1(P2_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n19798), .B1(
        n19844), .B2(n19863), .ZN(n19783) );
  OAI211_X1 U22808 ( .C1(n19866), .C2(n19801), .A(n19784), .B(n19783), .ZN(
        P2_U3152) );
  AOI22_X1 U22809 ( .A1(n19797), .A2(n19868), .B1(n19867), .B2(n19806), .ZN(
        n19786) );
  AOI22_X1 U22810 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19798), .B1(
        n19844), .B2(n19869), .ZN(n19785) );
  OAI211_X1 U22811 ( .C1(n19872), .C2(n19801), .A(n19786), .B(n19785), .ZN(
        P2_U3153) );
  AOI22_X1 U22812 ( .A1(n19797), .A2(n19874), .B1(n9966), .B2(n19806), .ZN(
        n19788) );
  AOI22_X1 U22813 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19798), .B1(
        n19844), .B2(n19875), .ZN(n19787) );
  OAI211_X1 U22814 ( .C1(n19878), .C2(n19801), .A(n19788), .B(n19787), .ZN(
        P2_U3154) );
  AOI22_X1 U22815 ( .A1(n19797), .A2(n19880), .B1(n19879), .B2(n19806), .ZN(
        n19790) );
  AOI22_X1 U22816 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19798), .B1(
        n19844), .B2(n19881), .ZN(n19789) );
  OAI211_X1 U22817 ( .C1(n19884), .C2(n19801), .A(n19790), .B(n19789), .ZN(
        P2_U3155) );
  AOI22_X1 U22818 ( .A1(n19797), .A2(n19886), .B1(n19885), .B2(n19806), .ZN(
        n19792) );
  AOI22_X1 U22819 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19798), .B1(
        n19844), .B2(n19887), .ZN(n19791) );
  OAI211_X1 U22820 ( .C1(n19890), .C2(n19801), .A(n19792), .B(n19791), .ZN(
        P2_U3156) );
  AOI22_X1 U22821 ( .A1(n19797), .A2(n19892), .B1(n19891), .B2(n19806), .ZN(
        n19794) );
  AOI22_X1 U22822 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19798), .B1(
        n19844), .B2(n19893), .ZN(n19793) );
  OAI211_X1 U22823 ( .C1(n19896), .C2(n19801), .A(n19794), .B(n19793), .ZN(
        P2_U3157) );
  AOI22_X1 U22824 ( .A1(n19797), .A2(n19898), .B1(n19897), .B2(n19806), .ZN(
        n19796) );
  AOI22_X1 U22825 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19798), .B1(
        n19844), .B2(n19899), .ZN(n19795) );
  OAI211_X1 U22826 ( .C1(n19902), .C2(n19801), .A(n19796), .B(n19795), .ZN(
        P2_U3158) );
  AOI22_X1 U22827 ( .A1(n19797), .A2(n19905), .B1(n19904), .B2(n19806), .ZN(
        n19800) );
  AOI22_X1 U22828 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n19798), .B1(
        n19844), .B2(n19907), .ZN(n19799) );
  OAI211_X1 U22829 ( .C1(n19913), .C2(n19801), .A(n19800), .B(n19799), .ZN(
        P2_U3159) );
  NAND3_X1 U22830 ( .A1(n19912), .A2(n19803), .A3(n20006), .ZN(n19805) );
  NAND2_X1 U22831 ( .A1(n19805), .A2(n19804), .ZN(n19809) );
  NAND3_X1 U22832 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19853), .A3(
        n20043), .ZN(n19810) );
  INV_X1 U22833 ( .A(n19810), .ZN(n19842) );
  OR2_X1 U22834 ( .A1(n19842), .A2(n19806), .ZN(n19813) );
  INV_X1 U22835 ( .A(n11223), .ZN(n19811) );
  AOI21_X1 U22836 ( .B1(n19811), .B2(n19810), .A(n20034), .ZN(n19807) );
  AOI22_X1 U22837 ( .A1(n19844), .A2(n19808), .B1(n19855), .B2(n19842), .ZN(
        n19816) );
  INV_X1 U22838 ( .A(n19809), .ZN(n19814) );
  OAI211_X1 U22839 ( .C1(n19811), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19810), 
        .B(n20002), .ZN(n19812) );
  OAI211_X1 U22840 ( .C1(n19814), .C2(n19813), .A(n19861), .B(n19812), .ZN(
        n19846) );
  AOI22_X1 U22841 ( .A1(P2_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n19846), .B1(
        n19845), .B2(n19863), .ZN(n19815) );
  OAI211_X1 U22842 ( .C1(n19850), .C2(n19817), .A(n19816), .B(n19815), .ZN(
        P2_U3160) );
  AOI22_X1 U22843 ( .A1(n19844), .A2(n19818), .B1(n19867), .B2(n19842), .ZN(
        n19820) );
  AOI22_X1 U22844 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n19846), .B1(
        n19845), .B2(n19869), .ZN(n19819) );
  OAI211_X1 U22845 ( .C1(n19850), .C2(n19821), .A(n19820), .B(n19819), .ZN(
        P2_U3161) );
  AOI22_X1 U22846 ( .A1(n19845), .A2(n19875), .B1(n9966), .B2(n19842), .ZN(
        n19824) );
  AOI22_X1 U22847 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n19846), .B1(
        n19844), .B2(n19822), .ZN(n19823) );
  OAI211_X1 U22848 ( .C1(n19850), .C2(n19825), .A(n19824), .B(n19823), .ZN(
        P2_U3162) );
  AOI22_X1 U22849 ( .A1(n19845), .A2(n19881), .B1(n19879), .B2(n19842), .ZN(
        n19828) );
  AOI22_X1 U22850 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n19846), .B1(
        n19844), .B2(n19826), .ZN(n19827) );
  OAI211_X1 U22851 ( .C1(n19850), .C2(n19829), .A(n19828), .B(n19827), .ZN(
        P2_U3163) );
  AOI22_X1 U22852 ( .A1(n19845), .A2(n19887), .B1(n19885), .B2(n19842), .ZN(
        n19832) );
  AOI22_X1 U22853 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n19846), .B1(
        n19844), .B2(n19830), .ZN(n19831) );
  OAI211_X1 U22854 ( .C1(n19850), .C2(n19833), .A(n19832), .B(n19831), .ZN(
        P2_U3164) );
  AOI22_X1 U22855 ( .A1(n19844), .A2(n19834), .B1(n19891), .B2(n19842), .ZN(
        n19836) );
  AOI22_X1 U22856 ( .A1(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n19846), .B1(
        n19845), .B2(n19893), .ZN(n19835) );
  OAI211_X1 U22857 ( .C1(n19850), .C2(n19837), .A(n19836), .B(n19835), .ZN(
        P2_U3165) );
  AOI22_X1 U22858 ( .A1(n19845), .A2(n19899), .B1(n19897), .B2(n19842), .ZN(
        n19840) );
  AOI22_X1 U22859 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n19846), .B1(
        n19844), .B2(n19838), .ZN(n19839) );
  OAI211_X1 U22860 ( .C1(n19850), .C2(n19841), .A(n19840), .B(n19839), .ZN(
        P2_U3166) );
  AOI22_X1 U22861 ( .A1(n19844), .A2(n19843), .B1(n19904), .B2(n19842), .ZN(
        n19848) );
  AOI22_X1 U22862 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n19846), .B1(
        n19845), .B2(n19907), .ZN(n19847) );
  OAI211_X1 U22863 ( .C1(n19850), .C2(n19849), .A(n19848), .B(n19847), .ZN(
        P2_U3167) );
  INV_X1 U22864 ( .A(n11210), .ZN(n19852) );
  NOR2_X1 U22865 ( .A1(n19903), .A2(n20034), .ZN(n19851) );
  NAND2_X1 U22866 ( .A1(n19852), .A2(n19851), .ZN(n19859) );
  NAND2_X1 U22867 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19853), .ZN(
        n19857) );
  OAI21_X1 U22868 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19857), .A(n20034), 
        .ZN(n19854) );
  AND2_X1 U22869 ( .A1(n19859), .A2(n19854), .ZN(n19906) );
  AOI22_X1 U22870 ( .A1(n19906), .A2(n19856), .B1(n19855), .B2(n19903), .ZN(
        n19865) );
  OAI21_X1 U22871 ( .B1(n19858), .B2(n20001), .A(n19857), .ZN(n19860) );
  AND2_X1 U22872 ( .A1(n19860), .A2(n19859), .ZN(n19862) );
  OAI211_X1 U22873 ( .C1(n19903), .C2(n20036), .A(n19862), .B(n19861), .ZN(
        n19909) );
  AOI22_X1 U22874 ( .A1(P2_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n19909), .B1(
        n19908), .B2(n19863), .ZN(n19864) );
  OAI211_X1 U22875 ( .C1(n19866), .C2(n19912), .A(n19865), .B(n19864), .ZN(
        P2_U3168) );
  AOI22_X1 U22876 ( .A1(n19906), .A2(n19868), .B1(n19867), .B2(n19903), .ZN(
        n19871) );
  AOI22_X1 U22877 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n19909), .B1(
        n19908), .B2(n19869), .ZN(n19870) );
  OAI211_X1 U22878 ( .C1(n19872), .C2(n19912), .A(n19871), .B(n19870), .ZN(
        P2_U3169) );
  AOI22_X1 U22879 ( .A1(n19906), .A2(n19874), .B1(n9966), .B2(n19903), .ZN(
        n19877) );
  AOI22_X1 U22880 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n19909), .B1(
        n19908), .B2(n19875), .ZN(n19876) );
  OAI211_X1 U22881 ( .C1(n19878), .C2(n19912), .A(n19877), .B(n19876), .ZN(
        P2_U3170) );
  AOI22_X1 U22882 ( .A1(n19906), .A2(n19880), .B1(n19879), .B2(n19903), .ZN(
        n19883) );
  AOI22_X1 U22883 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n19909), .B1(
        n19908), .B2(n19881), .ZN(n19882) );
  OAI211_X1 U22884 ( .C1(n19884), .C2(n19912), .A(n19883), .B(n19882), .ZN(
        P2_U3171) );
  AOI22_X1 U22885 ( .A1(n19906), .A2(n19886), .B1(n19885), .B2(n19903), .ZN(
        n19889) );
  AOI22_X1 U22886 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n19909), .B1(
        n19908), .B2(n19887), .ZN(n19888) );
  OAI211_X1 U22887 ( .C1(n19890), .C2(n19912), .A(n19889), .B(n19888), .ZN(
        P2_U3172) );
  AOI22_X1 U22888 ( .A1(n19906), .A2(n19892), .B1(n19891), .B2(n19903), .ZN(
        n19895) );
  AOI22_X1 U22889 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n19909), .B1(
        n19908), .B2(n19893), .ZN(n19894) );
  OAI211_X1 U22890 ( .C1(n19896), .C2(n19912), .A(n19895), .B(n19894), .ZN(
        P2_U3173) );
  AOI22_X1 U22891 ( .A1(n19906), .A2(n19898), .B1(n19897), .B2(n19903), .ZN(
        n19901) );
  AOI22_X1 U22892 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n19909), .B1(
        n19908), .B2(n19899), .ZN(n19900) );
  OAI211_X1 U22893 ( .C1(n19902), .C2(n19912), .A(n19901), .B(n19900), .ZN(
        P2_U3174) );
  AOI22_X1 U22894 ( .A1(n19906), .A2(n19905), .B1(n19904), .B2(n19903), .ZN(
        n19911) );
  AOI22_X1 U22895 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n19909), .B1(
        n19908), .B2(n19907), .ZN(n19910) );
  OAI211_X1 U22896 ( .C1(n19913), .C2(n19912), .A(n19911), .B(n19910), .ZN(
        P2_U3175) );
  AND2_X1 U22897 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n19914), .ZN(
        P2_U3179) );
  AND2_X1 U22898 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n19914), .ZN(
        P2_U3180) );
  AND2_X1 U22899 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n19914), .ZN(
        P2_U3181) );
  AND2_X1 U22900 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n19914), .ZN(
        P2_U3182) );
  AND2_X1 U22901 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n19914), .ZN(
        P2_U3183) );
  AND2_X1 U22902 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n19914), .ZN(
        P2_U3184) );
  AND2_X1 U22903 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n19914), .ZN(
        P2_U3185) );
  AND2_X1 U22904 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n19914), .ZN(
        P2_U3186) );
  AND2_X1 U22905 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n19914), .ZN(
        P2_U3187) );
  AND2_X1 U22906 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n19914), .ZN(
        P2_U3188) );
  AND2_X1 U22907 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n19914), .ZN(
        P2_U3189) );
  AND2_X1 U22908 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n19914), .ZN(
        P2_U3190) );
  AND2_X1 U22909 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n19914), .ZN(
        P2_U3191) );
  AND2_X1 U22910 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n19914), .ZN(
        P2_U3192) );
  AND2_X1 U22911 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n19914), .ZN(
        P2_U3193) );
  AND2_X1 U22912 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n19914), .ZN(
        P2_U3194) );
  AND2_X1 U22913 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n19914), .ZN(
        P2_U3195) );
  AND2_X1 U22914 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n19914), .ZN(
        P2_U3196) );
  AND2_X1 U22915 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n19914), .ZN(
        P2_U3197) );
  AND2_X1 U22916 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n19914), .ZN(
        P2_U3198) );
  AND2_X1 U22917 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n19914), .ZN(
        P2_U3199) );
  AND2_X1 U22918 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n19914), .ZN(
        P2_U3200) );
  AND2_X1 U22919 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n19914), .ZN(P2_U3201) );
  INV_X1 U22920 ( .A(P2_DATAWIDTH_REG_8__SCAN_IN), .ZN(n21303) );
  NOR2_X1 U22921 ( .A1(n21303), .A2(n20000), .ZN(P2_U3202) );
  AND2_X1 U22922 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n19914), .ZN(P2_U3203) );
  AND2_X1 U22923 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n19914), .ZN(P2_U3204) );
  AND2_X1 U22924 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n19914), .ZN(P2_U3205) );
  AND2_X1 U22925 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n19914), .ZN(P2_U3206) );
  AND2_X1 U22926 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n19914), .ZN(P2_U3207) );
  AND2_X1 U22927 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n19914), .ZN(P2_U3208) );
  NOR2_X1 U22928 ( .A1(n19915), .A2(n20069), .ZN(n19926) );
  INV_X1 U22929 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n20073) );
  OR3_X1 U22930 ( .A1(n19926), .A2(n20073), .A3(n21257), .ZN(n19917) );
  AOI211_X1 U22931 ( .C1(n20920), .C2(P2_REQUESTPENDING_REG_SCAN_IN), .A(
        n19927), .B(n19994), .ZN(n19916) );
  NOR2_X1 U22932 ( .A1(n20924), .A2(n19919), .ZN(n19932) );
  AOI211_X1 U22933 ( .C1(n19933), .C2(n19917), .A(n19916), .B(n19932), .ZN(
        n19918) );
  INV_X1 U22934 ( .A(n19918), .ZN(P2_U3209) );
  AOI21_X1 U22935 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(n20920), .A(n19933), 
        .ZN(n19923) );
  NOR2_X1 U22936 ( .A1(n20073), .A2(n19923), .ZN(n19920) );
  AOI21_X1 U22937 ( .B1(n19920), .B2(n19919), .A(n19926), .ZN(n19921) );
  OAI211_X1 U22938 ( .C1(n20920), .C2(n19922), .A(n19921), .B(n20063), .ZN(
        P2_U3210) );
  AOI21_X1 U22939 ( .B1(n19925), .B2(n19924), .A(n19923), .ZN(n19931) );
  AOI22_X1 U22940 ( .A1(n20073), .A2(n19927), .B1(n20924), .B2(n19926), .ZN(
        n19928) );
  INV_X1 U22941 ( .A(n19928), .ZN(n19929) );
  OAI211_X1 U22942 ( .C1(P2_REQUESTPENDING_REG_SCAN_IN), .C2(HOLD), .A(
        P2_STATE_REG_0__SCAN_IN), .B(n19929), .ZN(n19930) );
  OAI21_X1 U22943 ( .B1(n19932), .B2(n19931), .A(n19930), .ZN(P2_U3211) );
  NAND2_X2 U22944 ( .A1(n19994), .A2(n19933), .ZN(n19987) );
  NAND2_X2 U22945 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(n19994), .ZN(n19983) );
  OAI222_X1 U22946 ( .A1(n19987), .A2(n19936), .B1(n19935), .B2(n19994), .C1(
        n19934), .C2(n19983), .ZN(P2_U3212) );
  OAI222_X1 U22947 ( .A1(n19987), .A2(n19938), .B1(n19937), .B2(n19994), .C1(
        n19936), .C2(n19983), .ZN(P2_U3213) );
  OAI222_X1 U22948 ( .A1(n19987), .A2(n21299), .B1(n19939), .B2(n19994), .C1(
        n19938), .C2(n19983), .ZN(P2_U3214) );
  INV_X1 U22949 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n19941) );
  OAI222_X1 U22950 ( .A1(n19987), .A2(n19941), .B1(n19940), .B2(n19994), .C1(
        n21299), .C2(n19983), .ZN(P2_U3215) );
  OAI222_X1 U22951 ( .A1(n19987), .A2(n19943), .B1(n19942), .B2(n19994), .C1(
        n19941), .C2(n19983), .ZN(P2_U3216) );
  OAI222_X1 U22952 ( .A1(n19987), .A2(n19945), .B1(n19944), .B2(n19994), .C1(
        n19943), .C2(n19983), .ZN(P2_U3217) );
  OAI222_X1 U22953 ( .A1(n19987), .A2(n14167), .B1(n19946), .B2(n19994), .C1(
        n19945), .C2(n19983), .ZN(P2_U3218) );
  OAI222_X1 U22954 ( .A1(n19987), .A2(n19948), .B1(n19947), .B2(n19994), .C1(
        n14167), .C2(n19983), .ZN(P2_U3219) );
  OAI222_X1 U22955 ( .A1(n19987), .A2(n14180), .B1(n19949), .B2(n19994), .C1(
        n19948), .C2(n19983), .ZN(P2_U3220) );
  OAI222_X1 U22956 ( .A1(n19987), .A2(n15860), .B1(n19950), .B2(n19994), .C1(
        n14180), .C2(n19983), .ZN(P2_U3221) );
  OAI222_X1 U22957 ( .A1(n19987), .A2(n19952), .B1(n19951), .B2(n19994), .C1(
        n15860), .C2(n19983), .ZN(P2_U3222) );
  OAI222_X1 U22958 ( .A1(n19987), .A2(n15855), .B1(n19953), .B2(n19994), .C1(
        n19952), .C2(n19983), .ZN(P2_U3223) );
  OAI222_X1 U22959 ( .A1(n19987), .A2(n10868), .B1(n19954), .B2(n19994), .C1(
        n15855), .C2(n19983), .ZN(P2_U3224) );
  OAI222_X1 U22960 ( .A1(n19987), .A2(n19956), .B1(n19955), .B2(n19994), .C1(
        n10868), .C2(n19983), .ZN(P2_U3225) );
  OAI222_X1 U22961 ( .A1(n19987), .A2(n16011), .B1(n19957), .B2(n19994), .C1(
        n19956), .C2(n19983), .ZN(P2_U3226) );
  OAI222_X1 U22962 ( .A1(n19987), .A2(n19959), .B1(n19958), .B2(n19994), .C1(
        n16011), .C2(n19983), .ZN(P2_U3227) );
  OAI222_X1 U22963 ( .A1(n19987), .A2(n15994), .B1(n19960), .B2(n19994), .C1(
        n19959), .C2(n19983), .ZN(P2_U3228) );
  OAI222_X1 U22964 ( .A1(n19987), .A2(n19962), .B1(n19961), .B2(n19994), .C1(
        n15994), .C2(n19983), .ZN(P2_U3229) );
  OAI222_X1 U22965 ( .A1(n19987), .A2(n19964), .B1(n19963), .B2(n19994), .C1(
        n19962), .C2(n19983), .ZN(P2_U3230) );
  OAI222_X1 U22966 ( .A1(n19987), .A2(n19966), .B1(n19965), .B2(n19994), .C1(
        n19964), .C2(n19983), .ZN(P2_U3231) );
  INV_X1 U22967 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n19968) );
  OAI222_X1 U22968 ( .A1(n19987), .A2(n19968), .B1(n19967), .B2(n19994), .C1(
        n19966), .C2(n19983), .ZN(P2_U3232) );
  OAI222_X1 U22969 ( .A1(n19987), .A2(n19970), .B1(n19969), .B2(n19994), .C1(
        n19968), .C2(n19983), .ZN(P2_U3233) );
  OAI222_X1 U22970 ( .A1(n19987), .A2(n19972), .B1(n19971), .B2(n19994), .C1(
        n19970), .C2(n19983), .ZN(P2_U3234) );
  OAI222_X1 U22971 ( .A1(n19987), .A2(n19973), .B1(n21195), .B2(n19994), .C1(
        n19972), .C2(n19983), .ZN(P2_U3235) );
  INV_X1 U22972 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n19975) );
  OAI222_X1 U22973 ( .A1(n19987), .A2(n19975), .B1(n19974), .B2(n19994), .C1(
        n19973), .C2(n19983), .ZN(P2_U3236) );
  OAI222_X1 U22974 ( .A1(n19987), .A2(n19978), .B1(n19976), .B2(n19994), .C1(
        n19975), .C2(n19983), .ZN(P2_U3237) );
  INV_X1 U22975 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n19979) );
  OAI222_X1 U22976 ( .A1(n19983), .A2(n19978), .B1(n19977), .B2(n19994), .C1(
        n19979), .C2(n19987), .ZN(P2_U3238) );
  OAI222_X1 U22977 ( .A1(n19987), .A2(n19981), .B1(n19980), .B2(n19994), .C1(
        n19979), .C2(n19983), .ZN(P2_U3239) );
  INV_X1 U22978 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n19984) );
  OAI222_X1 U22979 ( .A1(n19987), .A2(n19984), .B1(n19982), .B2(n19994), .C1(
        n19981), .C2(n19983), .ZN(P2_U3240) );
  INV_X1 U22980 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n19986) );
  OAI222_X1 U22981 ( .A1(n19987), .A2(n19986), .B1(n19985), .B2(n19994), .C1(
        n19984), .C2(n19983), .ZN(P2_U3241) );
  INV_X1 U22982 ( .A(P2_BE_N_REG_3__SCAN_IN), .ZN(n19988) );
  AOI22_X1 U22983 ( .A1(n19994), .A2(n19989), .B1(n19988), .B2(n20075), .ZN(
        P2_U3585) );
  INV_X1 U22984 ( .A(P2_BE_N_REG_2__SCAN_IN), .ZN(n19990) );
  AOI22_X1 U22985 ( .A1(n19994), .A2(n19991), .B1(n19990), .B2(n20075), .ZN(
        P2_U3586) );
  INV_X1 U22986 ( .A(P2_BE_N_REG_1__SCAN_IN), .ZN(n19992) );
  AOI22_X1 U22987 ( .A1(n19994), .A2(n19993), .B1(n19992), .B2(n20075), .ZN(
        P2_U3587) );
  INV_X1 U22988 ( .A(P2_BE_N_REG_0__SCAN_IN), .ZN(n19995) );
  AOI22_X1 U22989 ( .A1(n19994), .A2(n19996), .B1(n19995), .B2(n20075), .ZN(
        P2_U3588) );
  OAI21_X1 U22990 ( .B1(n20000), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .A(n19998), 
        .ZN(n19997) );
  INV_X1 U22991 ( .A(n19997), .ZN(P2_U3591) );
  OAI21_X1 U22992 ( .B1(n20000), .B2(n19999), .A(n19998), .ZN(P2_U3592) );
  INV_X1 U22993 ( .A(n20041), .ZN(n20044) );
  OR3_X1 U22994 ( .A1(n20003), .A2(n20002), .A3(n20001), .ZN(n20012) );
  OR2_X1 U22995 ( .A1(n20004), .A2(n20028), .ZN(n20009) );
  NAND2_X1 U22996 ( .A1(n20029), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n20007) );
  AOI21_X1 U22997 ( .B1(n20007), .B2(n20006), .A(n20005), .ZN(n20008) );
  NAND2_X1 U22998 ( .A1(n20009), .A2(n20008), .ZN(n20020) );
  NAND2_X1 U22999 ( .A1(n20020), .A2(n20010), .ZN(n20011) );
  OAI211_X1 U23000 ( .C1(n20014), .C2(n20013), .A(n20012), .B(n20011), .ZN(
        n20015) );
  INV_X1 U23001 ( .A(n20015), .ZN(n20016) );
  AOI22_X1 U23002 ( .A1(n20044), .A2(n20017), .B1(n20016), .B2(n20041), .ZN(
        P2_U3602) );
  OAI21_X1 U23003 ( .B1(n20026), .B2(n20028), .A(n20018), .ZN(n20019) );
  AOI22_X1 U23004 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n20021), .B1(n20020), 
        .B2(n20019), .ZN(n20022) );
  AOI22_X1 U23005 ( .A1(n20044), .A2(n20023), .B1(n20022), .B2(n20041), .ZN(
        P2_U3603) );
  INV_X1 U23006 ( .A(n20039), .ZN(n20025) );
  OR3_X1 U23007 ( .A1(n20026), .A2(n20025), .A3(n20024), .ZN(n20027) );
  OAI21_X1 U23008 ( .B1(n20029), .B2(n20028), .A(n20027), .ZN(n20030) );
  AOI21_X1 U23009 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n20031), .A(n20030), 
        .ZN(n20032) );
  AOI22_X1 U23010 ( .A1(n20044), .A2(n20033), .B1(n20032), .B2(n20041), .ZN(
        P2_U3604) );
  NOR2_X1 U23011 ( .A1(n20035), .A2(n20034), .ZN(n20038) );
  NOR2_X1 U23012 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20036), .ZN(
        n20037) );
  AOI211_X1 U23013 ( .C1(n20040), .C2(n20039), .A(n20038), .B(n20037), .ZN(
        n20042) );
  AOI22_X1 U23014 ( .A1(n20044), .A2(n20043), .B1(n20042), .B2(n20041), .ZN(
        P2_U3605) );
  INV_X1 U23015 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n20045) );
  AOI22_X1 U23016 ( .A1(n19994), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n20045), 
        .B2(n20075), .ZN(P2_U3608) );
  INV_X1 U23017 ( .A(n20046), .ZN(n20053) );
  INV_X1 U23018 ( .A(n20047), .ZN(n20051) );
  AOI22_X1 U23019 ( .A1(n20051), .A2(n20050), .B1(n20049), .B2(n20048), .ZN(
        n20052) );
  NAND2_X1 U23020 ( .A1(n20053), .A2(n20052), .ZN(n20055) );
  MUX2_X1 U23021 ( .A(P2_MORE_REG_SCAN_IN), .B(n20055), .S(n20054), .Z(
        P2_U3609) );
  AOI21_X1 U23022 ( .B1(n20057), .B2(n20069), .A(n20056), .ZN(n20058) );
  OAI21_X1 U23023 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n20059), .A(n20058), 
        .ZN(n20074) );
  OAI21_X1 U23024 ( .B1(n20061), .B2(n20063), .A(n20060), .ZN(n20066) );
  NAND3_X1 U23025 ( .A1(n20064), .A2(n20063), .A3(n20062), .ZN(n20065) );
  AOI21_X1 U23026 ( .B1(n20066), .B2(n20065), .A(n14298), .ZN(n20071) );
  NOR2_X1 U23027 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n20067), .ZN(n20068) );
  AOI21_X1 U23028 ( .B1(P2_STATE2_REG_2__SCAN_IN), .B2(n20069), .A(n20068), 
        .ZN(n20070) );
  OAI21_X1 U23029 ( .B1(n20071), .B2(n20070), .A(n20074), .ZN(n20072) );
  OAI21_X1 U23030 ( .B1(n20074), .B2(n20073), .A(n20072), .ZN(P2_U3610) );
  OAI22_X1 U23031 ( .A1(n20075), .A2(P2_MEMORYFETCH_REG_SCAN_IN), .B1(
        P2_M_IO_N_REG_SCAN_IN), .B2(n19994), .ZN(n20076) );
  INV_X1 U23032 ( .A(n20076), .ZN(P2_U3611) );
  NAND2_X1 U23033 ( .A1(n20928), .A2(P1_STATE_REG_1__SCAN_IN), .ZN(n20918) );
  AND2_X1 U23034 ( .A1(n20918), .A2(P1_STATE_REG_0__SCAN_IN), .ZN(n20079) );
  INV_X1 U23035 ( .A(P1_ADS_N_REG_SCAN_IN), .ZN(n20078) );
  INV_X2 U23036 ( .A(n20997), .ZN(n21013) );
  AOI21_X1 U23037 ( .B1(n20079), .B2(n20078), .A(n21013), .ZN(P1_U2802) );
  NAND2_X1 U23038 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n20080), .ZN(n20083) );
  OAI21_X1 U23039 ( .B1(n20081), .B2(n20086), .A(P1_CODEFETCH_REG_SCAN_IN), 
        .ZN(n20082) );
  OAI21_X1 U23040 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n20083), .A(n20082), 
        .ZN(P1_U2803) );
  NOR2_X1 U23041 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(P1_STATE_REG_0__SCAN_IN), 
        .ZN(n20085) );
  OAI21_X1 U23042 ( .B1(n20085), .B2(P1_D_C_N_REG_SCAN_IN), .A(n20997), .ZN(
        n20084) );
  OAI21_X1 U23043 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(n20997), .A(n20084), 
        .ZN(P1_U2804) );
  OAI21_X1 U23044 ( .B1(BS16), .B2(n20085), .A(n20989), .ZN(n20987) );
  OAI21_X1 U23045 ( .B1(n20989), .B2(n21000), .A(n20987), .ZN(P1_U2805) );
  NOR2_X1 U23046 ( .A1(n20087), .A2(n20086), .ZN(n21399) );
  OAI21_X1 U23047 ( .B1(n21399), .B2(n20089), .A(n20088), .ZN(P1_U2806) );
  NOR4_X1 U23048 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_21__SCAN_IN), .A3(P1_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_23__SCAN_IN), .ZN(n20093) );
  NOR4_X1 U23049 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_17__SCAN_IN), .A3(P1_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_19__SCAN_IN), .ZN(n20092) );
  NOR4_X1 U23050 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_29__SCAN_IN), .A3(P1_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_31__SCAN_IN), .ZN(n20091) );
  NOR4_X1 U23051 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_25__SCAN_IN), .A3(P1_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_27__SCAN_IN), .ZN(n20090) );
  NAND4_X1 U23052 ( .A1(n20093), .A2(n20092), .A3(n20091), .A4(n20090), .ZN(
        n20099) );
  NOR4_X1 U23053 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_5__SCAN_IN), .A3(P1_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_7__SCAN_IN), .ZN(n20097) );
  AOI211_X1 U23054 ( .C1(P1_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A(P1_DATAWIDTH_REG_2__SCAN_IN), .B(
        P1_DATAWIDTH_REG_3__SCAN_IN), .ZN(n20096) );
  NOR4_X1 U23055 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_13__SCAN_IN), .A3(P1_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_15__SCAN_IN), .ZN(n20095) );
  NOR4_X1 U23056 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_9__SCAN_IN), .A3(P1_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_11__SCAN_IN), .ZN(n20094) );
  NAND4_X1 U23057 ( .A1(n20097), .A2(n20096), .A3(n20095), .A4(n20094), .ZN(
        n20098) );
  NOR2_X1 U23058 ( .A1(n20099), .A2(n20098), .ZN(n20996) );
  INV_X1 U23059 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n20982) );
  NOR3_X1 U23060 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A3(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n20101) );
  OAI21_X1 U23061 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n20101), .A(n20996), .ZN(
        n20100) );
  OAI21_X1 U23062 ( .B1(n20996), .B2(n20982), .A(n20100), .ZN(P1_U2807) );
  INV_X1 U23063 ( .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20988) );
  AOI21_X1 U23064 ( .B1(n13576), .B2(n20988), .A(n20101), .ZN(n20102) );
  INV_X1 U23065 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n20980) );
  INV_X1 U23066 ( .A(n20996), .ZN(n20991) );
  AOI22_X1 U23067 ( .A1(n20996), .A2(n20102), .B1(n20980), .B2(n20991), .ZN(
        P1_U2808) );
  AOI22_X1 U23068 ( .A1(n20103), .A2(n20149), .B1(n20147), .B2(
        P1_EBX_REG_9__SCAN_IN), .ZN(n20111) );
  OAI22_X1 U23069 ( .A1(P1_REIP_REG_9__SCAN_IN), .A2(n20105), .B1(n20104), 
        .B2(n20158), .ZN(n20106) );
  AOI211_X1 U23070 ( .C1(n20154), .C2(n20107), .A(n20280), .B(n20106), .ZN(
        n20110) );
  AOI22_X1 U23071 ( .A1(n20167), .A2(n20131), .B1(P1_REIP_REG_9__SCAN_IN), 
        .B2(n20108), .ZN(n20109) );
  NAND3_X1 U23072 ( .A1(n20111), .A2(n20110), .A3(n20109), .ZN(P1_U2831) );
  AOI22_X1 U23073 ( .A1(n20170), .A2(n20149), .B1(n20147), .B2(
        P1_EBX_REG_7__SCAN_IN), .ZN(n20121) );
  NOR2_X1 U23074 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(n20112), .ZN(n20116) );
  NOR2_X1 U23075 ( .A1(n20151), .A2(n20136), .ZN(n20139) );
  INV_X1 U23076 ( .A(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n20114) );
  OAI22_X1 U23077 ( .A1(n20114), .A2(n20158), .B1(n20113), .B2(n20143), .ZN(
        n20115) );
  AOI21_X1 U23078 ( .B1(n20116), .B2(n20139), .A(n20115), .ZN(n20120) );
  OAI21_X1 U23079 ( .B1(n20151), .B2(n20118), .A(n20117), .ZN(n20130) );
  AOI22_X1 U23080 ( .A1(n20172), .A2(n20131), .B1(P1_REIP_REG_7__SCAN_IN), 
        .B2(n20130), .ZN(n20119) );
  NAND4_X1 U23081 ( .A1(n20121), .A2(n20120), .A3(n20119), .A4(n20256), .ZN(
        P1_U2833) );
  OAI22_X1 U23082 ( .A1(n20125), .A2(n20124), .B1(n20123), .B2(n20122), .ZN(
        n20129) );
  INV_X1 U23083 ( .A(P1_REIP_REG_6__SCAN_IN), .ZN(n21198) );
  NAND3_X1 U23084 ( .A1(P1_REIP_REG_5__SCAN_IN), .A2(n20139), .A3(n21198), 
        .ZN(n20126) );
  OAI211_X1 U23085 ( .C1(n20143), .C2(n20127), .A(n20256), .B(n20126), .ZN(
        n20128) );
  AOI211_X1 U23086 ( .C1(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .C2(n20140), .A(
        n20129), .B(n20128), .ZN(n20134) );
  AOI22_X1 U23087 ( .A1(n20132), .A2(n20131), .B1(P1_REIP_REG_6__SCAN_IN), 
        .B2(n20130), .ZN(n20133) );
  NAND2_X1 U23088 ( .A1(n20134), .A2(n20133), .ZN(P1_U2834) );
  AOI21_X1 U23089 ( .B1(n20137), .B2(n20136), .A(n20135), .ZN(n20164) );
  INV_X1 U23090 ( .A(P1_REIP_REG_5__SCAN_IN), .ZN(n20935) );
  AOI22_X1 U23091 ( .A1(n20149), .A2(n20138), .B1(n20147), .B2(
        P1_EBX_REG_5__SCAN_IN), .ZN(n20146) );
  AOI22_X1 U23092 ( .A1(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n20140), .B1(
        n20139), .B2(n20935), .ZN(n20141) );
  OAI211_X1 U23093 ( .C1(n20143), .C2(n20142), .A(n20141), .B(n20256), .ZN(
        n20144) );
  AOI21_X1 U23094 ( .B1(n20179), .B2(n20161), .A(n20144), .ZN(n20145) );
  OAI211_X1 U23095 ( .C1(n20164), .C2(n20935), .A(n20146), .B(n20145), .ZN(
        P1_U2835) );
  INV_X1 U23096 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n20933) );
  INV_X1 U23097 ( .A(n20257), .ZN(n20148) );
  AOI22_X1 U23098 ( .A1(n20149), .A2(n20148), .B1(n20147), .B2(
        P1_EBX_REG_4__SCAN_IN), .ZN(n20163) );
  NAND3_X1 U23099 ( .A1(P1_REIP_REG_3__SCAN_IN), .A2(P1_REIP_REG_1__SCAN_IN), 
        .A3(P1_REIP_REG_2__SCAN_IN), .ZN(n20150) );
  NOR3_X1 U23100 ( .A1(n20151), .A2(P1_REIP_REG_4__SCAN_IN), .A3(n20150), .ZN(
        n20160) );
  INV_X1 U23101 ( .A(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n20157) );
  AOI22_X1 U23102 ( .A1(n20155), .A2(n20154), .B1(n20153), .B2(n20152), .ZN(
        n20156) );
  OAI211_X1 U23103 ( .C1(n20158), .C2(n20157), .A(n20156), .B(n20256), .ZN(
        n20159) );
  AOI211_X1 U23104 ( .C1(n20247), .C2(n20161), .A(n20160), .B(n20159), .ZN(
        n20162) );
  OAI211_X1 U23105 ( .C1(n20164), .C2(n20933), .A(n20163), .B(n20162), .ZN(
        P1_U2836) );
  NOR2_X1 U23106 ( .A1(n20165), .A2(n20175), .ZN(n20166) );
  AOI21_X1 U23107 ( .B1(n20167), .B2(n20178), .A(n20166), .ZN(n20168) );
  OAI21_X1 U23108 ( .B1(n20182), .B2(n20169), .A(n20168), .ZN(P1_U2863) );
  INV_X1 U23109 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n20174) );
  AOI22_X1 U23110 ( .A1(n20172), .A2(n20178), .B1(n20171), .B2(n20170), .ZN(
        n20173) );
  OAI21_X1 U23111 ( .B1(n20182), .B2(n20174), .A(n20173), .ZN(P1_U2865) );
  INV_X1 U23112 ( .A(P1_EBX_REG_5__SCAN_IN), .ZN(n20181) );
  NOR2_X1 U23113 ( .A1(n20176), .A2(n20175), .ZN(n20177) );
  AOI21_X1 U23114 ( .B1(n20179), .B2(n20178), .A(n20177), .ZN(n20180) );
  OAI21_X1 U23115 ( .B1(n20182), .B2(n20181), .A(n20180), .ZN(P1_U2867) );
  AOI22_X1 U23116 ( .A1(P1_EAX_REG_15__SCAN_IN), .A2(n20187), .B1(n20204), 
        .B2(P1_DATAO_REG_15__SCAN_IN), .ZN(n20183) );
  OAI21_X1 U23117 ( .B1(n20184), .B2(n20189), .A(n20183), .ZN(P1_U2921) );
  AOI22_X1 U23118 ( .A1(P1_LWORD_REG_14__SCAN_IN), .A2(n13910), .B1(n20204), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n20185) );
  OAI21_X1 U23119 ( .B1(n15110), .B2(n20208), .A(n20185), .ZN(P1_U2922) );
  AOI22_X1 U23120 ( .A1(P1_LWORD_REG_13__SCAN_IN), .A2(n13910), .B1(n20204), 
        .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n20186) );
  OAI21_X1 U23121 ( .B1(n15112), .B2(n20208), .A(n20186), .ZN(P1_U2923) );
  INV_X1 U23122 ( .A(P1_LWORD_REG_12__SCAN_IN), .ZN(n21240) );
  AOI22_X1 U23123 ( .A1(P1_EAX_REG_12__SCAN_IN), .A2(n20187), .B1(
        P1_DATAO_REG_12__SCAN_IN), .B2(n20204), .ZN(n20188) );
  OAI21_X1 U23124 ( .B1(n21240), .B2(n20189), .A(n20188), .ZN(P1_U2924) );
  AOI22_X1 U23125 ( .A1(P1_LWORD_REG_11__SCAN_IN), .A2(n13910), .B1(n20204), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n20190) );
  OAI21_X1 U23126 ( .B1(n15115), .B2(n20208), .A(n20190), .ZN(P1_U2925) );
  AOI22_X1 U23127 ( .A1(P1_LWORD_REG_10__SCAN_IN), .A2(n13910), .B1(n20204), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n20191) );
  OAI21_X1 U23128 ( .B1(n14493), .B2(n20208), .A(n20191), .ZN(P1_U2926) );
  AOI22_X1 U23129 ( .A1(P1_LWORD_REG_9__SCAN_IN), .A2(n13910), .B1(n20204), 
        .B2(P1_DATAO_REG_9__SCAN_IN), .ZN(n20192) );
  OAI21_X1 U23130 ( .B1(n14497), .B2(n20208), .A(n20192), .ZN(P1_U2927) );
  AOI22_X1 U23131 ( .A1(P1_LWORD_REG_8__SCAN_IN), .A2(n13910), .B1(n20204), 
        .B2(P1_DATAO_REG_8__SCAN_IN), .ZN(n20193) );
  OAI21_X1 U23132 ( .B1(n14400), .B2(n20208), .A(n20193), .ZN(P1_U2928) );
  AOI22_X1 U23133 ( .A1(P1_LWORD_REG_7__SCAN_IN), .A2(n13910), .B1(n20204), 
        .B2(P1_DATAO_REG_7__SCAN_IN), .ZN(n20194) );
  OAI21_X1 U23134 ( .B1(n12035), .B2(n20208), .A(n20194), .ZN(P1_U2929) );
  AOI22_X1 U23135 ( .A1(P1_LWORD_REG_6__SCAN_IN), .A2(n13910), .B1(n20204), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n20195) );
  OAI21_X1 U23136 ( .B1(n12029), .B2(n20208), .A(n20195), .ZN(P1_U2930) );
  AOI22_X1 U23137 ( .A1(P1_DATAO_REG_5__SCAN_IN), .A2(n20204), .B1(
        P1_LWORD_REG_5__SCAN_IN), .B2(n13910), .ZN(n20196) );
  OAI21_X1 U23138 ( .B1(n20197), .B2(n20208), .A(n20196), .ZN(P1_U2931) );
  INV_X1 U23139 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n20199) );
  AOI22_X1 U23140 ( .A1(P1_LWORD_REG_4__SCAN_IN), .A2(n13910), .B1(n20204), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .ZN(n20198) );
  OAI21_X1 U23141 ( .B1(n20199), .B2(n20208), .A(n20198), .ZN(P1_U2932) );
  AOI22_X1 U23142 ( .A1(P1_LWORD_REG_3__SCAN_IN), .A2(n13910), .B1(n20204), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n20200) );
  OAI21_X1 U23143 ( .B1(n20201), .B2(n20208), .A(n20200), .ZN(P1_U2933) );
  AOI22_X1 U23144 ( .A1(P1_LWORD_REG_2__SCAN_IN), .A2(n13910), .B1(n20204), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n20202) );
  OAI21_X1 U23145 ( .B1(n20203), .B2(n20208), .A(n20202), .ZN(P1_U2934) );
  AOI22_X1 U23146 ( .A1(P1_DATAO_REG_1__SCAN_IN), .A2(n20204), .B1(
        P1_LWORD_REG_1__SCAN_IN), .B2(n13910), .ZN(n20205) );
  OAI21_X1 U23147 ( .B1(n20206), .B2(n20208), .A(n20205), .ZN(P1_U2935) );
  AOI22_X1 U23148 ( .A1(P1_LWORD_REG_0__SCAN_IN), .A2(n13910), .B1(n20204), 
        .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n20207) );
  OAI21_X1 U23149 ( .B1(n20209), .B2(n20208), .A(n20207), .ZN(P1_U2936) );
  AOI22_X1 U23150 ( .A1(n20239), .A2(P1_EAX_REG_24__SCAN_IN), .B1(n20238), 
        .B2(P1_UWORD_REG_8__SCAN_IN), .ZN(n20212) );
  INV_X1 U23151 ( .A(n20210), .ZN(n20211) );
  NAND2_X1 U23152 ( .A1(n20224), .A2(n20211), .ZN(n20226) );
  NAND2_X1 U23153 ( .A1(n20212), .A2(n20226), .ZN(P1_U2945) );
  AOI22_X1 U23154 ( .A1(n20239), .A2(P1_EAX_REG_25__SCAN_IN), .B1(n20238), 
        .B2(P1_UWORD_REG_9__SCAN_IN), .ZN(n20215) );
  INV_X1 U23155 ( .A(n20213), .ZN(n20214) );
  NAND2_X1 U23156 ( .A1(n20224), .A2(n20214), .ZN(n20228) );
  NAND2_X1 U23157 ( .A1(n20215), .A2(n20228), .ZN(P1_U2946) );
  AOI22_X1 U23158 ( .A1(n20239), .A2(P1_EAX_REG_26__SCAN_IN), .B1(n20238), 
        .B2(P1_UWORD_REG_10__SCAN_IN), .ZN(n20218) );
  INV_X1 U23159 ( .A(n20216), .ZN(n20217) );
  NAND2_X1 U23160 ( .A1(n20224), .A2(n20217), .ZN(n20230) );
  NAND2_X1 U23161 ( .A1(n20218), .A2(n20230), .ZN(P1_U2947) );
  AOI22_X1 U23162 ( .A1(n20239), .A2(P1_EAX_REG_28__SCAN_IN), .B1(n20238), 
        .B2(P1_UWORD_REG_12__SCAN_IN), .ZN(n20221) );
  INV_X1 U23163 ( .A(n20219), .ZN(n20220) );
  NAND2_X1 U23164 ( .A1(n20224), .A2(n20220), .ZN(n20234) );
  NAND2_X1 U23165 ( .A1(n20221), .A2(n20234), .ZN(P1_U2949) );
  AOI22_X1 U23166 ( .A1(n20239), .A2(P1_EAX_REG_29__SCAN_IN), .B1(n20238), 
        .B2(P1_UWORD_REG_13__SCAN_IN), .ZN(n20225) );
  INV_X1 U23167 ( .A(n20222), .ZN(n20223) );
  NAND2_X1 U23168 ( .A1(n20224), .A2(n20223), .ZN(n20236) );
  NAND2_X1 U23169 ( .A1(n20225), .A2(n20236), .ZN(P1_U2950) );
  AOI22_X1 U23170 ( .A1(n20239), .A2(P1_EAX_REG_8__SCAN_IN), .B1(n20238), .B2(
        P1_LWORD_REG_8__SCAN_IN), .ZN(n20227) );
  NAND2_X1 U23171 ( .A1(n20227), .A2(n20226), .ZN(P1_U2960) );
  AOI22_X1 U23172 ( .A1(n20239), .A2(P1_EAX_REG_9__SCAN_IN), .B1(n20238), .B2(
        P1_LWORD_REG_9__SCAN_IN), .ZN(n20229) );
  NAND2_X1 U23173 ( .A1(n20229), .A2(n20228), .ZN(P1_U2961) );
  AOI22_X1 U23174 ( .A1(n20239), .A2(P1_EAX_REG_10__SCAN_IN), .B1(n20238), 
        .B2(P1_LWORD_REG_10__SCAN_IN), .ZN(n20231) );
  NAND2_X1 U23175 ( .A1(n20231), .A2(n20230), .ZN(P1_U2962) );
  AOI22_X1 U23176 ( .A1(n20239), .A2(P1_EAX_REG_11__SCAN_IN), .B1(n20238), 
        .B2(P1_LWORD_REG_11__SCAN_IN), .ZN(n20233) );
  NAND2_X1 U23177 ( .A1(n20233), .A2(n20232), .ZN(P1_U2963) );
  AOI22_X1 U23178 ( .A1(n20239), .A2(P1_EAX_REG_12__SCAN_IN), .B1(n20238), 
        .B2(P1_LWORD_REG_12__SCAN_IN), .ZN(n20235) );
  NAND2_X1 U23179 ( .A1(n20235), .A2(n20234), .ZN(P1_U2964) );
  AOI22_X1 U23180 ( .A1(n20239), .A2(P1_EAX_REG_13__SCAN_IN), .B1(n20238), 
        .B2(P1_LWORD_REG_13__SCAN_IN), .ZN(n20237) );
  NAND2_X1 U23181 ( .A1(n20237), .A2(n20236), .ZN(P1_U2965) );
  AOI22_X1 U23182 ( .A1(n20239), .A2(P1_EAX_REG_14__SCAN_IN), .B1(n20238), 
        .B2(P1_LWORD_REG_14__SCAN_IN), .ZN(n20241) );
  NAND2_X1 U23183 ( .A1(n20241), .A2(n20240), .ZN(P1_U2966) );
  AOI22_X1 U23184 ( .A1(n20242), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .B1(
        n20296), .B2(P1_REIP_REG_4__SCAN_IN), .ZN(n20250) );
  OAI21_X1 U23185 ( .B1(n20245), .B2(n20244), .A(n9833), .ZN(n20246) );
  INV_X1 U23186 ( .A(n20246), .ZN(n20265) );
  AOI22_X1 U23187 ( .A1(n20265), .A2(n20248), .B1(n16325), .B2(n20247), .ZN(
        n20249) );
  OAI211_X1 U23188 ( .C1(n20252), .C2(n20251), .A(n20250), .B(n20249), .ZN(
        P1_U2995) );
  OAI22_X1 U23189 ( .A1(n20254), .A2(n20260), .B1(n20253), .B2(n20261), .ZN(
        n20255) );
  NOR2_X1 U23190 ( .A1(n20277), .A2(n20255), .ZN(n20272) );
  OAI22_X1 U23191 ( .A1(n20292), .A2(n20257), .B1(n20933), .B2(n20256), .ZN(
        n20264) );
  INV_X1 U23192 ( .A(n20258), .ZN(n20259) );
  AOI22_X1 U23193 ( .A1(n20289), .A2(n20261), .B1(n20260), .B2(n20259), .ZN(
        n20274) );
  AOI211_X1 U23194 ( .C1(n20267), .C2(n20273), .A(n20274), .B(n20262), .ZN(
        n20263) );
  AOI211_X1 U23195 ( .C1(n20265), .C2(n20278), .A(n20264), .B(n20263), .ZN(
        n20266) );
  OAI21_X1 U23196 ( .B1(n20272), .B2(n20267), .A(n20266), .ZN(P1_U3027) );
  INV_X1 U23197 ( .A(n20268), .ZN(n20269) );
  AOI222_X1 U23198 ( .A1(P1_REIP_REG_3__SCAN_IN), .A2(n20280), .B1(n20282), 
        .B2(n20270), .C1(n20278), .C2(n20269), .ZN(n20271) );
  OAI221_X1 U23199 ( .B1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n20274), .C1(
        n20273), .C2(n20272), .A(n20271), .ZN(P1_U3028) );
  NAND2_X1 U23200 ( .A1(n20276), .A2(n20275), .ZN(n20287) );
  AOI21_X1 U23201 ( .B1(n20289), .B2(n13535), .A(n20277), .ZN(n20299) );
  NAND3_X1 U23202 ( .A1(n20279), .A2(n13579), .A3(n20278), .ZN(n20284) );
  AOI22_X1 U23203 ( .A1(n20282), .A2(n20281), .B1(n20280), .B2(
        P1_REIP_REG_1__SCAN_IN), .ZN(n20283) );
  AND2_X1 U23204 ( .A1(n20284), .A2(n20283), .ZN(n20285) );
  OAI221_X1 U23205 ( .B1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n20287), .C1(
        n20286), .C2(n20299), .A(n20285), .ZN(P1_U3030) );
  NOR3_X1 U23206 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n20289), .A3(
        n20288), .ZN(n20300) );
  INV_X1 U23207 ( .A(n20290), .ZN(n20294) );
  OAI22_X1 U23208 ( .A1(n20294), .A2(n20293), .B1(n20292), .B2(n20291), .ZN(
        n20295) );
  AOI21_X1 U23209 ( .B1(n20296), .B2(P1_REIP_REG_0__SCAN_IN), .A(n20295), .ZN(
        n20297) );
  OAI221_X1 U23210 ( .B1(n20300), .B2(n20299), .C1(n20300), .C2(n20298), .A(
        n20297), .ZN(P1_U3031) );
  NOR2_X1 U23211 ( .A1(n20302), .A2(n20301), .ZN(P1_U3032) );
  NOR2_X2 U23212 ( .A1(n20303), .A2(n20306), .ZN(n20304) );
  AOI22_X1 U23213 ( .A1(DATAI_16_), .A2(n20304), .B1(BUF1_REG_16__SCAN_IN), 
        .B2(n20345), .ZN(n20809) );
  AOI22_X1 U23214 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n20345), .B1(DATAI_24_), 
        .B2(n20304), .ZN(n20862) );
  INV_X1 U23215 ( .A(n20862), .ZN(n20806) );
  INV_X1 U23216 ( .A(n20732), .ZN(n20308) );
  NAND2_X1 U23217 ( .A1(n20387), .A2(n20598), .ZN(n20421) );
  INV_X1 U23218 ( .A(n20421), .ZN(n20419) );
  NAND2_X1 U23219 ( .A1(n20308), .A2(n20419), .ZN(n20314) );
  INV_X1 U23220 ( .A(n20314), .ZN(n20351) );
  NAND2_X1 U23221 ( .A1(n20341), .A2(n11644), .ZN(n20659) );
  AOI22_X1 U23222 ( .A1(n20904), .A2(n20806), .B1(n20351), .B2(n20853), .ZN(
        n20324) );
  OR2_X1 U23223 ( .A1(n20599), .A2(n20656), .ZN(n20320) );
  INV_X1 U23224 ( .A(n20320), .ZN(n20461) );
  OR2_X1 U23225 ( .A1(n20318), .A2(n20999), .ZN(n20796) );
  INV_X1 U23226 ( .A(n20904), .ZN(n20311) );
  NAND3_X1 U23227 ( .A1(n20311), .A2(n20769), .A3(n20378), .ZN(n20312) );
  NAND2_X1 U23228 ( .A1(n20769), .A2(n21000), .ZN(n20727) );
  NAND2_X1 U23229 ( .A1(n20312), .A2(n20727), .ZN(n20317) );
  NAND2_X1 U23230 ( .A1(n9946), .A2(n13838), .ZN(n20321) );
  AOI22_X1 U23231 ( .A1(n20317), .A2(n20321), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20314), .ZN(n20315) );
  NAND2_X1 U23232 ( .A1(n20316), .A2(n20353), .ZN(n20741) );
  INV_X1 U23233 ( .A(n20317), .ZN(n20322) );
  INV_X1 U23234 ( .A(n20318), .ZN(n20319) );
  NOR2_X1 U23235 ( .A1(n20319), .A2(n20999), .ZN(n20657) );
  INV_X1 U23236 ( .A(n20657), .ZN(n20601) );
  AOI22_X1 U23237 ( .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n20355), .B1(
        n20852), .B2(n20354), .ZN(n20323) );
  OAI211_X1 U23238 ( .C1(n20809), .C2(n20378), .A(n20324), .B(n20323), .ZN(
        P1_U3033) );
  AOI22_X1 U23239 ( .A1(DATAI_17_), .A2(n20304), .B1(BUF1_REG_17__SCAN_IN), 
        .B2(n20345), .ZN(n20813) );
  AOI22_X1 U23240 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n20345), .B1(DATAI_25_), 
        .B2(n20304), .ZN(n20868) );
  INV_X1 U23241 ( .A(n20868), .ZN(n20810) );
  NOR2_X2 U23242 ( .A1(n20350), .A2(n11633), .ZN(n20864) );
  AOI22_X1 U23243 ( .A1(n20904), .A2(n20810), .B1(n20351), .B2(n20864), .ZN(
        n20327) );
  NAND2_X1 U23244 ( .A1(n20325), .A2(n20353), .ZN(n20744) );
  AOI22_X1 U23245 ( .A1(P1_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n20355), .B1(
        n20863), .B2(n20354), .ZN(n20326) );
  OAI211_X1 U23246 ( .C1(n20813), .C2(n20378), .A(n20327), .B(n20326), .ZN(
        P1_U3034) );
  AOI22_X1 U23247 ( .A1(DATAI_18_), .A2(n20304), .B1(BUF1_REG_18__SCAN_IN), 
        .B2(n20345), .ZN(n20817) );
  AOI22_X1 U23248 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n20345), .B1(DATAI_26_), 
        .B2(n20304), .ZN(n20874) );
  INV_X1 U23249 ( .A(n20874), .ZN(n20814) );
  NAND2_X1 U23250 ( .A1(n20341), .A2(n11640), .ZN(n20671) );
  AOI22_X1 U23251 ( .A1(n20904), .A2(n20814), .B1(n20351), .B2(n20869), .ZN(
        n20330) );
  NOR2_X2 U23252 ( .A1(n20328), .A2(n20469), .ZN(n20870) );
  AOI22_X1 U23253 ( .A1(P1_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n20355), .B1(
        n20870), .B2(n20354), .ZN(n20329) );
  OAI211_X1 U23254 ( .C1(n20817), .C2(n20378), .A(n20330), .B(n20329), .ZN(
        P1_U3035) );
  AOI22_X1 U23255 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n20345), .B1(DATAI_19_), 
        .B2(n20304), .ZN(n20821) );
  AOI22_X1 U23256 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n20345), .B1(DATAI_27_), 
        .B2(n20304), .ZN(n20880) );
  INV_X1 U23257 ( .A(n20880), .ZN(n20818) );
  NAND2_X1 U23258 ( .A1(n20341), .A2(n20331), .ZN(n20675) );
  AOI22_X1 U23259 ( .A1(n20904), .A2(n20818), .B1(n20351), .B2(n20876), .ZN(
        n20334) );
  NAND2_X1 U23260 ( .A1(n20332), .A2(n20353), .ZN(n20750) );
  AOI22_X1 U23261 ( .A1(P1_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n20355), .B1(
        n20875), .B2(n20354), .ZN(n20333) );
  OAI211_X1 U23262 ( .C1(n20821), .C2(n20378), .A(n20334), .B(n20333), .ZN(
        P1_U3036) );
  AOI22_X1 U23263 ( .A1(DATAI_20_), .A2(n20304), .B1(BUF1_REG_20__SCAN_IN), 
        .B2(n20345), .ZN(n20825) );
  AOI22_X1 U23264 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n20345), .B1(DATAI_28_), 
        .B2(n20304), .ZN(n20886) );
  INV_X1 U23265 ( .A(n20886), .ZN(n20822) );
  NOR2_X2 U23266 ( .A1(n20350), .A2(n11679), .ZN(n20882) );
  AOI22_X1 U23267 ( .A1(n20904), .A2(n20822), .B1(n20351), .B2(n20882), .ZN(
        n20337) );
  NAND2_X1 U23268 ( .A1(n20335), .A2(n20353), .ZN(n20753) );
  AOI22_X1 U23269 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n20355), .B1(
        n20881), .B2(n20354), .ZN(n20336) );
  OAI211_X1 U23270 ( .C1(n20825), .C2(n20378), .A(n20337), .B(n20336), .ZN(
        P1_U3037) );
  AOI22_X1 U23271 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n20345), .B1(DATAI_21_), 
        .B2(n20304), .ZN(n20829) );
  AOI22_X1 U23272 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n20345), .B1(DATAI_29_), 
        .B2(n20304), .ZN(n20892) );
  INV_X1 U23273 ( .A(n20892), .ZN(n20826) );
  NOR2_X2 U23274 ( .A1(n20350), .A2(n11641), .ZN(n20887) );
  AOI22_X1 U23275 ( .A1(n20904), .A2(n20826), .B1(n20351), .B2(n20887), .ZN(
        n20340) );
  AOI22_X1 U23276 ( .A1(P1_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n20355), .B1(
        n20888), .B2(n20354), .ZN(n20339) );
  OAI211_X1 U23277 ( .C1(n20829), .C2(n20378), .A(n20340), .B(n20339), .ZN(
        P1_U3038) );
  AOI22_X1 U23278 ( .A1(DATAI_22_), .A2(n20304), .B1(BUF1_REG_22__SCAN_IN), 
        .B2(n20345), .ZN(n20833) );
  AOI22_X1 U23279 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n20345), .B1(DATAI_30_), 
        .B2(n20304), .ZN(n20898) );
  INV_X1 U23280 ( .A(n20898), .ZN(n20830) );
  NAND2_X1 U23281 ( .A1(n20341), .A2(n12766), .ZN(n20684) );
  AOI22_X1 U23282 ( .A1(n20904), .A2(n20830), .B1(n20351), .B2(n20893), .ZN(
        n20344) );
  AOI22_X1 U23283 ( .A1(P1_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n20355), .B1(
        n20894), .B2(n20354), .ZN(n20343) );
  OAI211_X1 U23284 ( .C1(n20833), .C2(n20378), .A(n20344), .B(n20343), .ZN(
        P1_U3039) );
  AOI22_X1 U23285 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n20345), .B1(DATAI_23_), 
        .B2(n20304), .ZN(n20841) );
  INV_X1 U23286 ( .A(DATAI_31_), .ZN(n21300) );
  INV_X1 U23287 ( .A(n20304), .ZN(n20348) );
  INV_X1 U23288 ( .A(n20345), .ZN(n20346) );
  OAI22_X1 U23289 ( .A1(n21300), .A2(n20348), .B1(n20347), .B2(n20346), .ZN(
        n20836) );
  NOR2_X2 U23290 ( .A1(n20350), .A2(n20349), .ZN(n20900) );
  AOI22_X1 U23291 ( .A1(n20904), .A2(n20836), .B1(n20351), .B2(n20900), .ZN(
        n20357) );
  AOI22_X1 U23292 ( .A1(P1_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n20355), .B1(
        n20902), .B2(n20354), .ZN(n20356) );
  OAI211_X1 U23293 ( .C1(n20841), .C2(n20378), .A(n20357), .B(n20356), .ZN(
        P1_U3040) );
  INV_X1 U23294 ( .A(n20358), .ZN(n20625) );
  NOR3_X2 U23295 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20767), .A3(
        n20421), .ZN(n20379) );
  AOI21_X1 U23296 ( .B1(n9946), .B2(n20625), .A(n20379), .ZN(n20360) );
  NOR2_X1 U23297 ( .A1(n20421), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n20362) );
  INV_X1 U23298 ( .A(n20362), .ZN(n20359) );
  OAI22_X1 U23299 ( .A1(n20360), .A2(n20848), .B1(n20359), .B2(n20999), .ZN(
        n20380) );
  AOI22_X1 U23300 ( .A1(n20380), .A2(n20852), .B1(n20853), .B2(n20379), .ZN(
        n20364) );
  OAI21_X1 U23301 ( .B1(n20425), .B2(n20628), .A(n20360), .ZN(n20361) );
  OAI221_X1 U23302 ( .B1(n20769), .B2(n20362), .C1(n20848), .C2(n20361), .A(
        n20856), .ZN(n20382) );
  INV_X1 U23303 ( .A(n20378), .ZN(n20381) );
  AOI22_X1 U23304 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n20382), .B1(
        n20381), .B2(n20806), .ZN(n20363) );
  OAI211_X1 U23305 ( .C1(n20809), .C2(n20418), .A(n20364), .B(n20363), .ZN(
        P1_U3041) );
  AOI22_X1 U23306 ( .A1(n20380), .A2(n20863), .B1(n20864), .B2(n20379), .ZN(
        n20366) );
  INV_X1 U23307 ( .A(n20813), .ZN(n20865) );
  AOI22_X1 U23308 ( .A1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n20382), .B1(
        n20375), .B2(n20865), .ZN(n20365) );
  OAI211_X1 U23309 ( .C1(n20868), .C2(n20378), .A(n20366), .B(n20365), .ZN(
        P1_U3042) );
  AOI22_X1 U23310 ( .A1(n20380), .A2(n20870), .B1(n20869), .B2(n20379), .ZN(
        n20368) );
  INV_X1 U23311 ( .A(n20817), .ZN(n20871) );
  AOI22_X1 U23312 ( .A1(P1_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n20382), .B1(
        n20375), .B2(n20871), .ZN(n20367) );
  OAI211_X1 U23313 ( .C1(n20874), .C2(n20378), .A(n20368), .B(n20367), .ZN(
        P1_U3043) );
  AOI22_X1 U23314 ( .A1(n20380), .A2(n20875), .B1(n20876), .B2(n20379), .ZN(
        n20370) );
  AOI22_X1 U23315 ( .A1(P1_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n20382), .B1(
        n20381), .B2(n20818), .ZN(n20369) );
  OAI211_X1 U23316 ( .C1(n20821), .C2(n20418), .A(n20370), .B(n20369), .ZN(
        P1_U3044) );
  AOI22_X1 U23317 ( .A1(n20380), .A2(n20881), .B1(n20882), .B2(n20379), .ZN(
        n20372) );
  INV_X1 U23318 ( .A(n20825), .ZN(n20883) );
  AOI22_X1 U23319 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n20382), .B1(
        n20375), .B2(n20883), .ZN(n20371) );
  OAI211_X1 U23320 ( .C1(n20886), .C2(n20378), .A(n20372), .B(n20371), .ZN(
        P1_U3045) );
  AOI22_X1 U23321 ( .A1(n20380), .A2(n20888), .B1(n20887), .B2(n20379), .ZN(
        n20374) );
  INV_X1 U23322 ( .A(n20829), .ZN(n20889) );
  AOI22_X1 U23323 ( .A1(P1_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n20382), .B1(
        n20375), .B2(n20889), .ZN(n20373) );
  OAI211_X1 U23324 ( .C1(n20892), .C2(n20378), .A(n20374), .B(n20373), .ZN(
        P1_U3046) );
  AOI22_X1 U23325 ( .A1(n20380), .A2(n20894), .B1(n20893), .B2(n20379), .ZN(
        n20377) );
  INV_X1 U23326 ( .A(n20833), .ZN(n20895) );
  AOI22_X1 U23327 ( .A1(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n20382), .B1(
        n20375), .B2(n20895), .ZN(n20376) );
  OAI211_X1 U23328 ( .C1(n20898), .C2(n20378), .A(n20377), .B(n20376), .ZN(
        P1_U3047) );
  AOI22_X1 U23329 ( .A1(n20380), .A2(n20902), .B1(n20900), .B2(n20379), .ZN(
        n20384) );
  AOI22_X1 U23330 ( .A1(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n20382), .B1(
        n20381), .B2(n20836), .ZN(n20383) );
  OAI211_X1 U23331 ( .C1(n20841), .C2(n20418), .A(n20384), .B(n20383), .ZN(
        P1_U3048) );
  OR3_X1 U23332 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20846), .A3(
        n20421), .ZN(n20412) );
  OAI22_X1 U23333 ( .A1(n20418), .A2(n20862), .B1(n20412), .B2(n20659), .ZN(
        n20385) );
  INV_X1 U23334 ( .A(n20385), .ZN(n20393) );
  NAND3_X1 U23335 ( .A1(n20459), .A2(n20418), .A3(n20769), .ZN(n20386) );
  NAND2_X1 U23336 ( .A1(n20386), .A2(n20727), .ZN(n20389) );
  NAND2_X1 U23337 ( .A1(n9946), .A2(n20799), .ZN(n20390) );
  AOI22_X1 U23338 ( .A1(n20389), .A2(n20390), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20412), .ZN(n20388) );
  NAND2_X1 U23339 ( .A1(n20656), .A2(n20387), .ZN(n20527) );
  NAND2_X1 U23340 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20527), .ZN(n20524) );
  NAND3_X1 U23341 ( .A1(n20663), .A2(n20388), .A3(n20524), .ZN(n20415) );
  INV_X1 U23342 ( .A(n20389), .ZN(n20391) );
  AOI22_X1 U23343 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n20415), .B1(
        n20852), .B2(n20414), .ZN(n20392) );
  OAI211_X1 U23344 ( .C1(n20809), .C2(n20459), .A(n20393), .B(n20392), .ZN(
        P1_U3049) );
  INV_X1 U23345 ( .A(n20864), .ZN(n20532) );
  OAI22_X1 U23346 ( .A1(n20418), .A2(n20868), .B1(n20412), .B2(n20532), .ZN(
        n20394) );
  INV_X1 U23347 ( .A(n20394), .ZN(n20396) );
  AOI22_X1 U23348 ( .A1(P1_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n20415), .B1(
        n20863), .B2(n20414), .ZN(n20395) );
  OAI211_X1 U23349 ( .C1(n20813), .C2(n20459), .A(n20396), .B(n20395), .ZN(
        P1_U3050) );
  OAI22_X1 U23350 ( .A1(n20418), .A2(n20874), .B1(n20412), .B2(n20671), .ZN(
        n20397) );
  INV_X1 U23351 ( .A(n20397), .ZN(n20399) );
  AOI22_X1 U23352 ( .A1(P1_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n20415), .B1(
        n20870), .B2(n20414), .ZN(n20398) );
  OAI211_X1 U23353 ( .C1(n20817), .C2(n20459), .A(n20399), .B(n20398), .ZN(
        P1_U3051) );
  OAI22_X1 U23354 ( .A1(n20418), .A2(n20880), .B1(n20412), .B2(n20675), .ZN(
        n20400) );
  INV_X1 U23355 ( .A(n20400), .ZN(n20402) );
  AOI22_X1 U23356 ( .A1(P1_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n20415), .B1(
        n20875), .B2(n20414), .ZN(n20401) );
  OAI211_X1 U23357 ( .C1(n20821), .C2(n20459), .A(n20402), .B(n20401), .ZN(
        P1_U3052) );
  INV_X1 U23358 ( .A(n20882), .ZN(n20542) );
  OAI22_X1 U23359 ( .A1(n20418), .A2(n20886), .B1(n20412), .B2(n20542), .ZN(
        n20403) );
  INV_X1 U23360 ( .A(n20403), .ZN(n20405) );
  AOI22_X1 U23361 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n20415), .B1(
        n20881), .B2(n20414), .ZN(n20404) );
  OAI211_X1 U23362 ( .C1(n20825), .C2(n20459), .A(n20405), .B(n20404), .ZN(
        P1_U3053) );
  INV_X1 U23363 ( .A(n20887), .ZN(n20546) );
  OAI22_X1 U23364 ( .A1(n20459), .A2(n20829), .B1(n20546), .B2(n20412), .ZN(
        n20406) );
  INV_X1 U23365 ( .A(n20406), .ZN(n20408) );
  AOI22_X1 U23366 ( .A1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n20415), .B1(
        n20888), .B2(n20414), .ZN(n20407) );
  OAI211_X1 U23367 ( .C1(n20892), .C2(n20418), .A(n20408), .B(n20407), .ZN(
        P1_U3054) );
  OAI22_X1 U23368 ( .A1(n20459), .A2(n20833), .B1(n20412), .B2(n20684), .ZN(
        n20409) );
  INV_X1 U23369 ( .A(n20409), .ZN(n20411) );
  AOI22_X1 U23370 ( .A1(P1_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n20415), .B1(
        n20894), .B2(n20414), .ZN(n20410) );
  OAI211_X1 U23371 ( .C1(n20898), .C2(n20418), .A(n20411), .B(n20410), .ZN(
        P1_U3055) );
  INV_X1 U23372 ( .A(n20836), .ZN(n20909) );
  INV_X1 U23373 ( .A(n20900), .ZN(n20554) );
  OAI22_X1 U23374 ( .A1(n20459), .A2(n20841), .B1(n20412), .B2(n20554), .ZN(
        n20413) );
  INV_X1 U23375 ( .A(n20413), .ZN(n20417) );
  AOI22_X1 U23376 ( .A1(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n20415), .B1(
        n20902), .B2(n20414), .ZN(n20416) );
  OAI211_X1 U23377 ( .C1(n20909), .C2(n20418), .A(n20417), .B(n20416), .ZN(
        P1_U3056) );
  NAND2_X1 U23378 ( .A1(n20843), .A2(n20419), .ZN(n20453) );
  OAI22_X1 U23379 ( .A1(n20459), .A2(n20862), .B1(n20659), .B2(n20453), .ZN(
        n20420) );
  INV_X1 U23380 ( .A(n20420), .ZN(n20434) );
  NOR2_X1 U23381 ( .A1(n20846), .A2(n20421), .ZN(n20429) );
  AND2_X1 U23382 ( .A1(n20423), .A2(n20422), .ZN(n20844) );
  INV_X1 U23383 ( .A(n20453), .ZN(n20424) );
  AOI21_X1 U23384 ( .B1(n9946), .B2(n20844), .A(n20424), .ZN(n20432) );
  OR2_X1 U23385 ( .A1(n20425), .A2(n20700), .ZN(n20426) );
  AND2_X1 U23386 ( .A1(n20426), .A2(n20769), .ZN(n20428) );
  NAND2_X1 U23387 ( .A1(n20432), .A2(n20428), .ZN(n20427) );
  OAI211_X1 U23388 ( .C1(n20769), .C2(n20429), .A(n20856), .B(n20427), .ZN(
        n20456) );
  INV_X1 U23389 ( .A(n20428), .ZN(n20431) );
  INV_X1 U23390 ( .A(n20429), .ZN(n20430) );
  OAI22_X1 U23391 ( .A1(n20432), .A2(n20431), .B1(n20999), .B2(n20430), .ZN(
        n20455) );
  AOI22_X1 U23392 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n20456), .B1(
        n20852), .B2(n20455), .ZN(n20433) );
  OAI211_X1 U23393 ( .C1(n20809), .C2(n20465), .A(n20434), .B(n20433), .ZN(
        P1_U3057) );
  OAI22_X1 U23394 ( .A1(n20459), .A2(n20868), .B1(n20453), .B2(n20532), .ZN(
        n20435) );
  INV_X1 U23395 ( .A(n20435), .ZN(n20437) );
  AOI22_X1 U23396 ( .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n20456), .B1(
        n20863), .B2(n20455), .ZN(n20436) );
  OAI211_X1 U23397 ( .C1(n20813), .C2(n20465), .A(n20437), .B(n20436), .ZN(
        P1_U3058) );
  OAI22_X1 U23398 ( .A1(n20465), .A2(n20817), .B1(n20453), .B2(n20671), .ZN(
        n20438) );
  INV_X1 U23399 ( .A(n20438), .ZN(n20440) );
  AOI22_X1 U23400 ( .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n20456), .B1(
        n20870), .B2(n20455), .ZN(n20439) );
  OAI211_X1 U23401 ( .C1(n20874), .C2(n20459), .A(n20440), .B(n20439), .ZN(
        P1_U3059) );
  OAI22_X1 U23402 ( .A1(n20459), .A2(n20880), .B1(n20453), .B2(n20675), .ZN(
        n20441) );
  INV_X1 U23403 ( .A(n20441), .ZN(n20443) );
  AOI22_X1 U23404 ( .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20456), .B1(
        n20875), .B2(n20455), .ZN(n20442) );
  OAI211_X1 U23405 ( .C1(n20821), .C2(n20465), .A(n20443), .B(n20442), .ZN(
        P1_U3060) );
  OAI22_X1 U23406 ( .A1(n20465), .A2(n20825), .B1(n20453), .B2(n20542), .ZN(
        n20444) );
  INV_X1 U23407 ( .A(n20444), .ZN(n20446) );
  AOI22_X1 U23408 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n20456), .B1(
        n20881), .B2(n20455), .ZN(n20445) );
  OAI211_X1 U23409 ( .C1(n20886), .C2(n20459), .A(n20446), .B(n20445), .ZN(
        P1_U3061) );
  OAI22_X1 U23410 ( .A1(n20465), .A2(n20829), .B1(n20546), .B2(n20453), .ZN(
        n20447) );
  INV_X1 U23411 ( .A(n20447), .ZN(n20449) );
  AOI22_X1 U23412 ( .A1(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n20456), .B1(
        n20888), .B2(n20455), .ZN(n20448) );
  OAI211_X1 U23413 ( .C1(n20892), .C2(n20459), .A(n20449), .B(n20448), .ZN(
        P1_U3062) );
  OAI22_X1 U23414 ( .A1(n20465), .A2(n20833), .B1(n20684), .B2(n20453), .ZN(
        n20450) );
  INV_X1 U23415 ( .A(n20450), .ZN(n20452) );
  AOI22_X1 U23416 ( .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20456), .B1(
        n20894), .B2(n20455), .ZN(n20451) );
  OAI211_X1 U23417 ( .C1(n20898), .C2(n20459), .A(n20452), .B(n20451), .ZN(
        P1_U3063) );
  OAI22_X1 U23418 ( .A1(n20465), .A2(n20841), .B1(n20554), .B2(n20453), .ZN(
        n20454) );
  INV_X1 U23419 ( .A(n20454), .ZN(n20458) );
  AOI22_X1 U23420 ( .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n20456), .B1(
        n20902), .B2(n20455), .ZN(n20457) );
  OAI211_X1 U23421 ( .C1(n20909), .C2(n20459), .A(n20458), .B(n20457), .ZN(
        P1_U3064) );
  OR2_X1 U23422 ( .A1(n20732), .A2(n20520), .ZN(n20478) );
  NOR2_X1 U23423 ( .A1(n13553), .A2(n20460), .ZN(n20561) );
  NAND3_X1 U23424 ( .A1(n20561), .A2(n20769), .A3(n13838), .ZN(n20463) );
  INV_X1 U23425 ( .A(n20796), .ZN(n20731) );
  NAND2_X1 U23426 ( .A1(n20461), .A2(n20731), .ZN(n20462) );
  NAND2_X1 U23427 ( .A1(n20463), .A2(n20462), .ZN(n20489) );
  INV_X1 U23428 ( .A(n20489), .ZN(n20477) );
  OAI22_X1 U23429 ( .A1(n20659), .A2(n20478), .B1(n20741), .B2(n20477), .ZN(
        n20464) );
  INV_X1 U23430 ( .A(n20464), .ZN(n20472) );
  INV_X1 U23431 ( .A(n20561), .ZN(n20468) );
  INV_X1 U23432 ( .A(n20519), .ZN(n20466) );
  OAI21_X1 U23433 ( .B1(n20490), .B2(n20466), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20467) );
  OAI21_X1 U23434 ( .B1(n20799), .B2(n20468), .A(n20467), .ZN(n20470) );
  AOI22_X1 U23435 ( .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n20491), .B1(
        n20490), .B2(n20806), .ZN(n20471) );
  OAI211_X1 U23436 ( .C1(n20809), .C2(n20519), .A(n20472), .B(n20471), .ZN(
        P1_U3065) );
  AOI22_X1 U23437 ( .A1(n20864), .A2(n20488), .B1(n20863), .B2(n20489), .ZN(
        n20474) );
  AOI22_X1 U23438 ( .A1(P1_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n20491), .B1(
        n20490), .B2(n20810), .ZN(n20473) );
  OAI211_X1 U23439 ( .C1(n20813), .C2(n20519), .A(n20474), .B(n20473), .ZN(
        P1_U3066) );
  AOI22_X1 U23440 ( .A1(n20870), .A2(n20489), .B1(n20869), .B2(n20488), .ZN(
        n20476) );
  AOI22_X1 U23441 ( .A1(P1_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n20491), .B1(
        n20490), .B2(n20814), .ZN(n20475) );
  OAI211_X1 U23442 ( .C1(n20817), .C2(n20519), .A(n20476), .B(n20475), .ZN(
        P1_U3067) );
  OAI22_X1 U23443 ( .A1(n20675), .A2(n20478), .B1(n20750), .B2(n20477), .ZN(
        n20479) );
  INV_X1 U23444 ( .A(n20479), .ZN(n20481) );
  AOI22_X1 U23445 ( .A1(P1_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n20491), .B1(
        n20490), .B2(n20818), .ZN(n20480) );
  OAI211_X1 U23446 ( .C1(n20821), .C2(n20519), .A(n20481), .B(n20480), .ZN(
        P1_U3068) );
  AOI22_X1 U23447 ( .A1(n20882), .A2(n20488), .B1(n20881), .B2(n20489), .ZN(
        n20483) );
  AOI22_X1 U23448 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n20491), .B1(
        n20490), .B2(n20822), .ZN(n20482) );
  OAI211_X1 U23449 ( .C1(n20825), .C2(n20519), .A(n20483), .B(n20482), .ZN(
        P1_U3069) );
  AOI22_X1 U23450 ( .A1(n20888), .A2(n20489), .B1(n20887), .B2(n20488), .ZN(
        n20485) );
  AOI22_X1 U23451 ( .A1(P1_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n20491), .B1(
        n20490), .B2(n20826), .ZN(n20484) );
  OAI211_X1 U23452 ( .C1(n20829), .C2(n20519), .A(n20485), .B(n20484), .ZN(
        P1_U3070) );
  AOI22_X1 U23453 ( .A1(n20894), .A2(n20489), .B1(n20893), .B2(n20488), .ZN(
        n20487) );
  AOI22_X1 U23454 ( .A1(P1_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n20491), .B1(
        n20490), .B2(n20830), .ZN(n20486) );
  OAI211_X1 U23455 ( .C1(n20833), .C2(n20519), .A(n20487), .B(n20486), .ZN(
        P1_U3071) );
  AOI22_X1 U23456 ( .A1(n20902), .A2(n20489), .B1(n20900), .B2(n20488), .ZN(
        n20493) );
  AOI22_X1 U23457 ( .A1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n20491), .B1(
        n20490), .B2(n20836), .ZN(n20492) );
  OAI211_X1 U23458 ( .C1(n20841), .C2(n20519), .A(n20493), .B(n20492), .ZN(
        P1_U3072) );
  NOR2_X1 U23459 ( .A1(n20520), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n20498) );
  INV_X1 U23460 ( .A(n20498), .ZN(n20494) );
  NOR2_X1 U23461 ( .A1(n20767), .A2(n20494), .ZN(n20513) );
  AOI21_X1 U23462 ( .B1(n20561), .B2(n20625), .A(n20513), .ZN(n20495) );
  OAI22_X1 U23463 ( .A1(n20495), .A2(n20848), .B1(n20494), .B2(n20999), .ZN(
        n20514) );
  AOI22_X1 U23464 ( .A1(n20853), .A2(n20513), .B1(n20514), .B2(n20852), .ZN(
        n20500) );
  OAI21_X1 U23465 ( .B1(n20496), .B2(n20628), .A(n20495), .ZN(n20497) );
  OAI221_X1 U23466 ( .B1(n20769), .B2(n20498), .C1(n20848), .C2(n20497), .A(
        n20856), .ZN(n20516) );
  INV_X1 U23467 ( .A(n20809), .ZN(n20859) );
  AOI22_X1 U23468 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n20516), .B1(
        n20515), .B2(n20859), .ZN(n20499) );
  OAI211_X1 U23469 ( .C1(n20862), .C2(n20519), .A(n20500), .B(n20499), .ZN(
        P1_U3073) );
  AOI22_X1 U23470 ( .A1(n20514), .A2(n20863), .B1(n20864), .B2(n20513), .ZN(
        n20502) );
  AOI22_X1 U23471 ( .A1(P1_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n20516), .B1(
        n20515), .B2(n20865), .ZN(n20501) );
  OAI211_X1 U23472 ( .C1(n20868), .C2(n20519), .A(n20502), .B(n20501), .ZN(
        P1_U3074) );
  AOI22_X1 U23473 ( .A1(n20870), .A2(n20514), .B1(n20869), .B2(n20513), .ZN(
        n20504) );
  AOI22_X1 U23474 ( .A1(P1_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n20516), .B1(
        n20515), .B2(n20871), .ZN(n20503) );
  OAI211_X1 U23475 ( .C1(n20874), .C2(n20519), .A(n20504), .B(n20503), .ZN(
        P1_U3075) );
  AOI22_X1 U23476 ( .A1(n20876), .A2(n20513), .B1(n20514), .B2(n20875), .ZN(
        n20506) );
  INV_X1 U23477 ( .A(n20821), .ZN(n20877) );
  AOI22_X1 U23478 ( .A1(P1_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n20516), .B1(
        n20515), .B2(n20877), .ZN(n20505) );
  OAI211_X1 U23479 ( .C1(n20880), .C2(n20519), .A(n20506), .B(n20505), .ZN(
        P1_U3076) );
  AOI22_X1 U23480 ( .A1(n20514), .A2(n20881), .B1(n20882), .B2(n20513), .ZN(
        n20508) );
  AOI22_X1 U23481 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n20516), .B1(
        n20515), .B2(n20883), .ZN(n20507) );
  OAI211_X1 U23482 ( .C1(n20886), .C2(n20519), .A(n20508), .B(n20507), .ZN(
        P1_U3077) );
  AOI22_X1 U23483 ( .A1(n20888), .A2(n20514), .B1(n20887), .B2(n20513), .ZN(
        n20510) );
  AOI22_X1 U23484 ( .A1(P1_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n20516), .B1(
        n20515), .B2(n20889), .ZN(n20509) );
  OAI211_X1 U23485 ( .C1(n20892), .C2(n20519), .A(n20510), .B(n20509), .ZN(
        P1_U3078) );
  AOI22_X1 U23486 ( .A1(n20894), .A2(n20514), .B1(n20893), .B2(n20513), .ZN(
        n20512) );
  AOI22_X1 U23487 ( .A1(P1_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n20516), .B1(
        n20515), .B2(n20895), .ZN(n20511) );
  OAI211_X1 U23488 ( .C1(n20898), .C2(n20519), .A(n20512), .B(n20511), .ZN(
        P1_U3079) );
  AOI22_X1 U23489 ( .A1(n20902), .A2(n20514), .B1(n20900), .B2(n20513), .ZN(
        n20518) );
  INV_X1 U23490 ( .A(n20841), .ZN(n20903) );
  AOI22_X1 U23491 ( .A1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n20516), .B1(
        n20515), .B2(n20903), .ZN(n20517) );
  OAI211_X1 U23492 ( .C1(n20909), .C2(n20519), .A(n20518), .B(n20517), .ZN(
        P1_U3080) );
  NOR2_X1 U23493 ( .A1(n20846), .A2(n20520), .ZN(n20568) );
  INV_X1 U23494 ( .A(n20568), .ZN(n20521) );
  OR2_X1 U23495 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20521), .ZN(
        n20553) );
  OAI22_X1 U23496 ( .A1(n20560), .A2(n20862), .B1(n20659), .B2(n20553), .ZN(
        n20522) );
  INV_X1 U23497 ( .A(n20522), .ZN(n20531) );
  NAND3_X1 U23498 ( .A1(n20592), .A2(n20560), .A3(n20769), .ZN(n20523) );
  NAND2_X1 U23499 ( .A1(n20523), .A2(n20727), .ZN(n20526) );
  NAND2_X1 U23500 ( .A1(n20561), .A2(n20799), .ZN(n20528) );
  AOI22_X1 U23501 ( .A1(n20526), .A2(n20528), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20553), .ZN(n20525) );
  NAND3_X1 U23502 ( .A1(n20803), .A2(n20525), .A3(n20524), .ZN(n20557) );
  INV_X1 U23503 ( .A(n20526), .ZN(n20529) );
  AOI22_X1 U23504 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n20557), .B1(
        n20852), .B2(n20556), .ZN(n20530) );
  OAI211_X1 U23505 ( .C1(n20809), .C2(n20592), .A(n20531), .B(n20530), .ZN(
        P1_U3081) );
  OAI22_X1 U23506 ( .A1(n20592), .A2(n20813), .B1(n20532), .B2(n20553), .ZN(
        n20533) );
  INV_X1 U23507 ( .A(n20533), .ZN(n20535) );
  AOI22_X1 U23508 ( .A1(P1_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n20557), .B1(
        n20863), .B2(n20556), .ZN(n20534) );
  OAI211_X1 U23509 ( .C1(n20868), .C2(n20560), .A(n20535), .B(n20534), .ZN(
        P1_U3082) );
  OAI22_X1 U23510 ( .A1(n20592), .A2(n20817), .B1(n20671), .B2(n20553), .ZN(
        n20536) );
  INV_X1 U23511 ( .A(n20536), .ZN(n20538) );
  AOI22_X1 U23512 ( .A1(P1_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n20557), .B1(
        n20870), .B2(n20556), .ZN(n20537) );
  OAI211_X1 U23513 ( .C1(n20874), .C2(n20560), .A(n20538), .B(n20537), .ZN(
        P1_U3083) );
  OAI22_X1 U23514 ( .A1(n20560), .A2(n20880), .B1(n20675), .B2(n20553), .ZN(
        n20539) );
  INV_X1 U23515 ( .A(n20539), .ZN(n20541) );
  AOI22_X1 U23516 ( .A1(P1_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n20557), .B1(
        n20875), .B2(n20556), .ZN(n20540) );
  OAI211_X1 U23517 ( .C1(n20821), .C2(n20592), .A(n20541), .B(n20540), .ZN(
        P1_U3084) );
  OAI22_X1 U23518 ( .A1(n20592), .A2(n20825), .B1(n20542), .B2(n20553), .ZN(
        n20543) );
  INV_X1 U23519 ( .A(n20543), .ZN(n20545) );
  AOI22_X1 U23520 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n20557), .B1(
        n20881), .B2(n20556), .ZN(n20544) );
  OAI211_X1 U23521 ( .C1(n20886), .C2(n20560), .A(n20545), .B(n20544), .ZN(
        P1_U3085) );
  OAI22_X1 U23522 ( .A1(n20592), .A2(n20829), .B1(n20546), .B2(n20553), .ZN(
        n20547) );
  INV_X1 U23523 ( .A(n20547), .ZN(n20549) );
  AOI22_X1 U23524 ( .A1(P1_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n20557), .B1(
        n20888), .B2(n20556), .ZN(n20548) );
  OAI211_X1 U23525 ( .C1(n20892), .C2(n20560), .A(n20549), .B(n20548), .ZN(
        P1_U3086) );
  OAI22_X1 U23526 ( .A1(n20560), .A2(n20898), .B1(n20684), .B2(n20553), .ZN(
        n20550) );
  INV_X1 U23527 ( .A(n20550), .ZN(n20552) );
  AOI22_X1 U23528 ( .A1(P1_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n20557), .B1(
        n20894), .B2(n20556), .ZN(n20551) );
  OAI211_X1 U23529 ( .C1(n20833), .C2(n20592), .A(n20552), .B(n20551), .ZN(
        P1_U3087) );
  OAI22_X1 U23530 ( .A1(n20592), .A2(n20841), .B1(n20554), .B2(n20553), .ZN(
        n20555) );
  INV_X1 U23531 ( .A(n20555), .ZN(n20559) );
  AOI22_X1 U23532 ( .A1(P1_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n20557), .B1(
        n20902), .B2(n20556), .ZN(n20558) );
  OAI211_X1 U23533 ( .C1(n20909), .C2(n20560), .A(n20559), .B(n20558), .ZN(
        P1_U3088) );
  INV_X1 U23534 ( .A(n20562), .ZN(n20587) );
  NAND2_X1 U23535 ( .A1(n20561), .A2(n20844), .ZN(n20563) );
  NAND2_X1 U23536 ( .A1(n20563), .A2(n20562), .ZN(n20564) );
  NAND2_X1 U23537 ( .A1(n20564), .A2(n20769), .ZN(n20566) );
  NAND2_X1 U23538 ( .A1(n20568), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20565) );
  NAND2_X1 U23539 ( .A1(n20566), .A2(n20565), .ZN(n20588) );
  AOI22_X1 U23540 ( .A1(n20853), .A2(n20587), .B1(n20852), .B2(n20588), .ZN(
        n20572) );
  OAI21_X1 U23541 ( .B1(n20568), .B2(n20567), .A(n20856), .ZN(n20589) );
  INV_X1 U23542 ( .A(n20703), .ZN(n20569) );
  NAND2_X1 U23543 ( .A1(n20570), .A2(n20569), .ZN(n20586) );
  AOI22_X1 U23544 ( .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n20589), .B1(
        n20621), .B2(n20859), .ZN(n20571) );
  OAI211_X1 U23545 ( .C1(n20862), .C2(n20592), .A(n20572), .B(n20571), .ZN(
        P1_U3089) );
  AOI22_X1 U23546 ( .A1(n20864), .A2(n20587), .B1(n20588), .B2(n20863), .ZN(
        n20574) );
  AOI22_X1 U23547 ( .A1(P1_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n20589), .B1(
        n20621), .B2(n20865), .ZN(n20573) );
  OAI211_X1 U23548 ( .C1(n20868), .C2(n20592), .A(n20574), .B(n20573), .ZN(
        P1_U3090) );
  AOI22_X1 U23549 ( .A1(n20870), .A2(n20588), .B1(n20869), .B2(n20587), .ZN(
        n20576) );
  AOI22_X1 U23550 ( .A1(P1_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n20589), .B1(
        n20621), .B2(n20871), .ZN(n20575) );
  OAI211_X1 U23551 ( .C1(n20874), .C2(n20592), .A(n20576), .B(n20575), .ZN(
        P1_U3091) );
  AOI22_X1 U23552 ( .A1(n20876), .A2(n20587), .B1(n20875), .B2(n20588), .ZN(
        n20578) );
  AOI22_X1 U23553 ( .A1(P1_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n20589), .B1(
        n20621), .B2(n20877), .ZN(n20577) );
  OAI211_X1 U23554 ( .C1(n20880), .C2(n20592), .A(n20578), .B(n20577), .ZN(
        P1_U3092) );
  AOI22_X1 U23555 ( .A1(n20882), .A2(n20587), .B1(n20588), .B2(n20881), .ZN(
        n20580) );
  AOI22_X1 U23556 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n20589), .B1(
        n20621), .B2(n20883), .ZN(n20579) );
  OAI211_X1 U23557 ( .C1(n20886), .C2(n20592), .A(n20580), .B(n20579), .ZN(
        P1_U3093) );
  AOI22_X1 U23558 ( .A1(n20888), .A2(n20588), .B1(n20887), .B2(n20587), .ZN(
        n20582) );
  AOI22_X1 U23559 ( .A1(P1_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n20589), .B1(
        n20621), .B2(n20889), .ZN(n20581) );
  OAI211_X1 U23560 ( .C1(n20892), .C2(n20592), .A(n20582), .B(n20581), .ZN(
        P1_U3094) );
  AOI22_X1 U23561 ( .A1(n20894), .A2(n20588), .B1(n20893), .B2(n20587), .ZN(
        n20585) );
  INV_X1 U23562 ( .A(n20592), .ZN(n20583) );
  AOI22_X1 U23563 ( .A1(P1_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n20589), .B1(
        n20583), .B2(n20830), .ZN(n20584) );
  OAI211_X1 U23564 ( .C1(n20833), .C2(n20586), .A(n20585), .B(n20584), .ZN(
        P1_U3095) );
  AOI22_X1 U23565 ( .A1(n20902), .A2(n20588), .B1(n20900), .B2(n20587), .ZN(
        n20591) );
  AOI22_X1 U23566 ( .A1(P1_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n20589), .B1(
        n20621), .B2(n20903), .ZN(n20590) );
  OAI211_X1 U23567 ( .C1(n20909), .C2(n20592), .A(n20591), .B(n20590), .ZN(
        P1_U3096) );
  INV_X1 U23568 ( .A(n20704), .ZN(n20596) );
  NAND2_X1 U23569 ( .A1(n20597), .A2(n13553), .ZN(n20655) );
  INV_X1 U23570 ( .A(n20655), .ZN(n20697) );
  NAND2_X1 U23571 ( .A1(n20598), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20695) );
  AOI21_X1 U23572 ( .B1(n20697), .B2(n13838), .A(n10375), .ZN(n20603) );
  INV_X1 U23573 ( .A(n20599), .ZN(n20600) );
  NOR2_X1 U23574 ( .A1(n20600), .A2(n20656), .ZN(n20730) );
  INV_X1 U23575 ( .A(n20730), .ZN(n20734) );
  OAI22_X1 U23576 ( .A1(n20603), .A2(n20848), .B1(n20601), .B2(n20734), .ZN(
        n20620) );
  AOI22_X1 U23577 ( .A1(n20620), .A2(n20852), .B1(n10375), .B2(n20853), .ZN(
        n20607) );
  INV_X1 U23578 ( .A(n20651), .ZN(n20602) );
  OAI21_X1 U23579 ( .B1(n20602), .B2(n20621), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20604) );
  NAND2_X1 U23580 ( .A1(n20604), .A2(n20603), .ZN(n20605) );
  AOI22_X1 U23581 ( .A1(P1_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n20622), .B1(
        n20621), .B2(n20806), .ZN(n20606) );
  OAI211_X1 U23582 ( .C1(n20809), .C2(n20651), .A(n20607), .B(n20606), .ZN(
        P1_U3097) );
  AOI22_X1 U23583 ( .A1(n20620), .A2(n20863), .B1(n10375), .B2(n20864), .ZN(
        n20609) );
  AOI22_X1 U23584 ( .A1(P1_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n20622), .B1(
        n20621), .B2(n20810), .ZN(n20608) );
  OAI211_X1 U23585 ( .C1(n20813), .C2(n20651), .A(n20609), .B(n20608), .ZN(
        P1_U3098) );
  AOI22_X1 U23586 ( .A1(n20620), .A2(n20870), .B1(n10375), .B2(n20869), .ZN(
        n20611) );
  AOI22_X1 U23587 ( .A1(P1_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n20622), .B1(
        n20621), .B2(n20814), .ZN(n20610) );
  OAI211_X1 U23588 ( .C1(n20817), .C2(n20651), .A(n20611), .B(n20610), .ZN(
        P1_U3099) );
  AOI22_X1 U23589 ( .A1(n20620), .A2(n20875), .B1(n10375), .B2(n20876), .ZN(
        n20613) );
  AOI22_X1 U23590 ( .A1(P1_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n20622), .B1(
        n20621), .B2(n20818), .ZN(n20612) );
  OAI211_X1 U23591 ( .C1(n20821), .C2(n20651), .A(n20613), .B(n20612), .ZN(
        P1_U3100) );
  AOI22_X1 U23592 ( .A1(n20620), .A2(n20881), .B1(n10375), .B2(n20882), .ZN(
        n20615) );
  AOI22_X1 U23593 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n20622), .B1(
        n20621), .B2(n20822), .ZN(n20614) );
  OAI211_X1 U23594 ( .C1(n20825), .C2(n20651), .A(n20615), .B(n20614), .ZN(
        P1_U3101) );
  AOI22_X1 U23595 ( .A1(n20620), .A2(n20888), .B1(n10375), .B2(n20887), .ZN(
        n20617) );
  AOI22_X1 U23596 ( .A1(P1_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n20622), .B1(
        n20621), .B2(n20826), .ZN(n20616) );
  OAI211_X1 U23597 ( .C1(n20829), .C2(n20651), .A(n20617), .B(n20616), .ZN(
        P1_U3102) );
  AOI22_X1 U23598 ( .A1(n20620), .A2(n20894), .B1(n10375), .B2(n20893), .ZN(
        n20619) );
  AOI22_X1 U23599 ( .A1(P1_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n20622), .B1(
        n20621), .B2(n20830), .ZN(n20618) );
  OAI211_X1 U23600 ( .C1(n20833), .C2(n20651), .A(n20619), .B(n20618), .ZN(
        P1_U3103) );
  AOI22_X1 U23601 ( .A1(n20620), .A2(n20902), .B1(n10375), .B2(n20900), .ZN(
        n20624) );
  AOI22_X1 U23602 ( .A1(P1_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n20622), .B1(
        n20621), .B2(n20836), .ZN(n20623) );
  OAI211_X1 U23603 ( .C1(n20841), .C2(n20651), .A(n20624), .B(n20623), .ZN(
        P1_U3104) );
  NOR2_X1 U23604 ( .A1(n20695), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n20630) );
  INV_X1 U23605 ( .A(n20630), .ZN(n20626) );
  NOR2_X1 U23606 ( .A1(n20767), .A2(n20626), .ZN(n20646) );
  AOI21_X1 U23607 ( .B1(n20697), .B2(n20625), .A(n20646), .ZN(n20627) );
  OAI22_X1 U23608 ( .A1(n20627), .A2(n20848), .B1(n20626), .B2(n20999), .ZN(
        n20647) );
  AOI22_X1 U23609 ( .A1(n20647), .A2(n20852), .B1(n20853), .B2(n20646), .ZN(
        n20633) );
  OAI21_X1 U23610 ( .B1(n20704), .B2(n20628), .A(n20627), .ZN(n20629) );
  OAI221_X1 U23611 ( .B1(n20769), .B2(n20630), .C1(n20848), .C2(n20629), .A(
        n20856), .ZN(n20648) );
  AOI22_X1 U23612 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n20648), .B1(
        n20689), .B2(n20859), .ZN(n20632) );
  OAI211_X1 U23613 ( .C1(n20862), .C2(n20651), .A(n20633), .B(n20632), .ZN(
        P1_U3105) );
  AOI22_X1 U23614 ( .A1(n20647), .A2(n20863), .B1(n20864), .B2(n20646), .ZN(
        n20635) );
  AOI22_X1 U23615 ( .A1(P1_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n20648), .B1(
        n20689), .B2(n20865), .ZN(n20634) );
  OAI211_X1 U23616 ( .C1(n20868), .C2(n20651), .A(n20635), .B(n20634), .ZN(
        P1_U3106) );
  AOI22_X1 U23617 ( .A1(n20647), .A2(n20870), .B1(n20869), .B2(n20646), .ZN(
        n20637) );
  AOI22_X1 U23618 ( .A1(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n20648), .B1(
        n20689), .B2(n20871), .ZN(n20636) );
  OAI211_X1 U23619 ( .C1(n20874), .C2(n20651), .A(n20637), .B(n20636), .ZN(
        P1_U3107) );
  AOI22_X1 U23620 ( .A1(n20647), .A2(n20875), .B1(n20876), .B2(n20646), .ZN(
        n20639) );
  AOI22_X1 U23621 ( .A1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n20648), .B1(
        n20689), .B2(n20877), .ZN(n20638) );
  OAI211_X1 U23622 ( .C1(n20880), .C2(n20651), .A(n20639), .B(n20638), .ZN(
        P1_U3108) );
  AOI22_X1 U23623 ( .A1(n20647), .A2(n20881), .B1(n20882), .B2(n20646), .ZN(
        n20641) );
  AOI22_X1 U23624 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n20648), .B1(
        n20689), .B2(n20883), .ZN(n20640) );
  OAI211_X1 U23625 ( .C1(n20886), .C2(n20651), .A(n20641), .B(n20640), .ZN(
        P1_U3109) );
  AOI22_X1 U23626 ( .A1(n20647), .A2(n20888), .B1(n20887), .B2(n20646), .ZN(
        n20643) );
  AOI22_X1 U23627 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n20648), .B1(
        n20689), .B2(n20889), .ZN(n20642) );
  OAI211_X1 U23628 ( .C1(n20892), .C2(n20651), .A(n20643), .B(n20642), .ZN(
        P1_U3110) );
  AOI22_X1 U23629 ( .A1(n20647), .A2(n20894), .B1(n20893), .B2(n20646), .ZN(
        n20645) );
  AOI22_X1 U23630 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n20648), .B1(
        n20689), .B2(n20895), .ZN(n20644) );
  OAI211_X1 U23631 ( .C1(n20898), .C2(n20651), .A(n20645), .B(n20644), .ZN(
        P1_U3111) );
  AOI22_X1 U23632 ( .A1(n20647), .A2(n20902), .B1(n20900), .B2(n20646), .ZN(
        n20650) );
  AOI22_X1 U23633 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n20648), .B1(
        n20689), .B2(n20903), .ZN(n20649) );
  OAI211_X1 U23634 ( .C1(n20909), .C2(n20651), .A(n20650), .B(n20649), .ZN(
        P1_U3112) );
  NAND3_X1 U23635 ( .A1(n20724), .A2(n20653), .A3(n20769), .ZN(n20654) );
  NAND2_X1 U23636 ( .A1(n20654), .A2(n20727), .ZN(n20661) );
  NOR2_X1 U23637 ( .A1(n20655), .A2(n13838), .ZN(n20665) );
  NAND2_X1 U23638 ( .A1(n20656), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20797) );
  INV_X1 U23639 ( .A(n20797), .ZN(n20658) );
  NOR2_X1 U23640 ( .A1(n20846), .A2(n20695), .ZN(n20702) );
  INV_X1 U23641 ( .A(n20702), .ZN(n20698) );
  NOR2_X1 U23642 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20698), .ZN(
        n20688) );
  INV_X1 U23643 ( .A(n20688), .ZN(n20683) );
  OAI22_X1 U23644 ( .A1(n20724), .A2(n20809), .B1(n20659), .B2(n20683), .ZN(
        n20660) );
  INV_X1 U23645 ( .A(n20660), .ZN(n20668) );
  INV_X1 U23646 ( .A(n20661), .ZN(n20666) );
  NAND2_X1 U23647 ( .A1(n20797), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20802) );
  OAI21_X1 U23648 ( .B1(n20738), .B2(n20688), .A(n20802), .ZN(n20662) );
  INV_X1 U23649 ( .A(n20662), .ZN(n20664) );
  AOI22_X1 U23650 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n20691), .B1(
        n20689), .B2(n20806), .ZN(n20667) );
  OAI211_X1 U23651 ( .C1(n20694), .C2(n20741), .A(n20668), .B(n20667), .ZN(
        P1_U3113) );
  AOI22_X1 U23652 ( .A1(n20689), .A2(n20810), .B1(n20864), .B2(n20688), .ZN(
        n20670) );
  INV_X1 U23653 ( .A(n20724), .ZN(n20690) );
  AOI22_X1 U23654 ( .A1(P1_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n20691), .B1(
        n20690), .B2(n20865), .ZN(n20669) );
  OAI211_X1 U23655 ( .C1(n20694), .C2(n20744), .A(n20670), .B(n20669), .ZN(
        P1_U3114) );
  INV_X1 U23656 ( .A(n20870), .ZN(n20747) );
  OAI22_X1 U23657 ( .A1(n20724), .A2(n20817), .B1(n20671), .B2(n20683), .ZN(
        n20672) );
  INV_X1 U23658 ( .A(n20672), .ZN(n20674) );
  AOI22_X1 U23659 ( .A1(P1_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n20691), .B1(
        n20689), .B2(n20814), .ZN(n20673) );
  OAI211_X1 U23660 ( .C1(n20694), .C2(n20747), .A(n20674), .B(n20673), .ZN(
        P1_U3115) );
  OAI22_X1 U23661 ( .A1(n20724), .A2(n20821), .B1(n20675), .B2(n20683), .ZN(
        n20676) );
  INV_X1 U23662 ( .A(n20676), .ZN(n20678) );
  AOI22_X1 U23663 ( .A1(P1_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n20691), .B1(
        n20689), .B2(n20818), .ZN(n20677) );
  OAI211_X1 U23664 ( .C1(n20694), .C2(n20750), .A(n20678), .B(n20677), .ZN(
        P1_U3116) );
  AOI22_X1 U23665 ( .A1(n20689), .A2(n20822), .B1(n20882), .B2(n20688), .ZN(
        n20680) );
  AOI22_X1 U23666 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n20691), .B1(
        n20690), .B2(n20883), .ZN(n20679) );
  OAI211_X1 U23667 ( .C1(n20694), .C2(n20753), .A(n20680), .B(n20679), .ZN(
        P1_U3117) );
  INV_X1 U23668 ( .A(n20888), .ZN(n20756) );
  AOI22_X1 U23669 ( .A1(n20689), .A2(n20826), .B1(n20887), .B2(n20688), .ZN(
        n20682) );
  AOI22_X1 U23670 ( .A1(P1_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n20691), .B1(
        n20690), .B2(n20889), .ZN(n20681) );
  OAI211_X1 U23671 ( .C1(n20694), .C2(n20756), .A(n20682), .B(n20681), .ZN(
        P1_U3118) );
  INV_X1 U23672 ( .A(n20894), .ZN(n20759) );
  OAI22_X1 U23673 ( .A1(n20724), .A2(n20833), .B1(n20684), .B2(n20683), .ZN(
        n20685) );
  INV_X1 U23674 ( .A(n20685), .ZN(n20687) );
  AOI22_X1 U23675 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n20691), .B1(
        n20689), .B2(n20830), .ZN(n20686) );
  OAI211_X1 U23676 ( .C1(n20694), .C2(n20759), .A(n20687), .B(n20686), .ZN(
        P1_U3119) );
  INV_X1 U23677 ( .A(n20902), .ZN(n20764) );
  AOI22_X1 U23678 ( .A1(n20689), .A2(n20836), .B1(n20900), .B2(n20688), .ZN(
        n20693) );
  AOI22_X1 U23679 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n20691), .B1(
        n20690), .B2(n20903), .ZN(n20692) );
  OAI211_X1 U23680 ( .C1(n20694), .C2(n20764), .A(n20693), .B(n20692), .ZN(
        P1_U3120) );
  NOR2_X1 U23681 ( .A1(n20696), .A2(n20695), .ZN(n20719) );
  AOI21_X1 U23682 ( .B1(n20697), .B2(n20844), .A(n20719), .ZN(n20699) );
  OAI22_X1 U23683 ( .A1(n20699), .A2(n20848), .B1(n20698), .B2(n20999), .ZN(
        n20720) );
  AOI22_X1 U23684 ( .A1(n20720), .A2(n20852), .B1(n20853), .B2(n20719), .ZN(
        n20706) );
  OAI21_X1 U23685 ( .B1(n20704), .B2(n20700), .A(n20699), .ZN(n20701) );
  OAI221_X1 U23686 ( .B1(n20769), .B2(n20702), .C1(n20848), .C2(n20701), .A(
        n20856), .ZN(n20721) );
  AOI22_X1 U23687 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n20721), .B1(
        n20760), .B2(n20859), .ZN(n20705) );
  OAI211_X1 U23688 ( .C1(n20862), .C2(n20724), .A(n20706), .B(n20705), .ZN(
        P1_U3121) );
  AOI22_X1 U23689 ( .A1(n20720), .A2(n20863), .B1(n20864), .B2(n20719), .ZN(
        n20708) );
  AOI22_X1 U23690 ( .A1(P1_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n20721), .B1(
        n20760), .B2(n20865), .ZN(n20707) );
  OAI211_X1 U23691 ( .C1(n20868), .C2(n20724), .A(n20708), .B(n20707), .ZN(
        P1_U3122) );
  AOI22_X1 U23692 ( .A1(n20720), .A2(n20870), .B1(n20869), .B2(n20719), .ZN(
        n20710) );
  AOI22_X1 U23693 ( .A1(P1_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n20721), .B1(
        n20760), .B2(n20871), .ZN(n20709) );
  OAI211_X1 U23694 ( .C1(n20874), .C2(n20724), .A(n20710), .B(n20709), .ZN(
        P1_U3123) );
  AOI22_X1 U23695 ( .A1(n20720), .A2(n20875), .B1(n20876), .B2(n20719), .ZN(
        n20712) );
  AOI22_X1 U23696 ( .A1(P1_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n20721), .B1(
        n20760), .B2(n20877), .ZN(n20711) );
  OAI211_X1 U23697 ( .C1(n20880), .C2(n20724), .A(n20712), .B(n20711), .ZN(
        P1_U3124) );
  AOI22_X1 U23698 ( .A1(n20720), .A2(n20881), .B1(n20882), .B2(n20719), .ZN(
        n20714) );
  AOI22_X1 U23699 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n20721), .B1(
        n20760), .B2(n20883), .ZN(n20713) );
  OAI211_X1 U23700 ( .C1(n20886), .C2(n20724), .A(n20714), .B(n20713), .ZN(
        P1_U3125) );
  AOI22_X1 U23701 ( .A1(n20720), .A2(n20888), .B1(n20887), .B2(n20719), .ZN(
        n20716) );
  AOI22_X1 U23702 ( .A1(P1_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n20721), .B1(
        n20760), .B2(n20889), .ZN(n20715) );
  OAI211_X1 U23703 ( .C1(n20892), .C2(n20724), .A(n20716), .B(n20715), .ZN(
        P1_U3126) );
  AOI22_X1 U23704 ( .A1(n20720), .A2(n20894), .B1(n20893), .B2(n20719), .ZN(
        n20718) );
  AOI22_X1 U23705 ( .A1(P1_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n20721), .B1(
        n20760), .B2(n20895), .ZN(n20717) );
  OAI211_X1 U23706 ( .C1(n20898), .C2(n20724), .A(n20718), .B(n20717), .ZN(
        P1_U3127) );
  AOI22_X1 U23707 ( .A1(n20720), .A2(n20902), .B1(n20900), .B2(n20719), .ZN(
        n20723) );
  AOI22_X1 U23708 ( .A1(P1_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n20721), .B1(
        n20760), .B2(n20903), .ZN(n20722) );
  OAI211_X1 U23709 ( .C1(n20909), .C2(n20724), .A(n20723), .B(n20722), .ZN(
        P1_U3128) );
  INV_X1 U23710 ( .A(n20790), .ZN(n20726) );
  NAND2_X1 U23711 ( .A1(n20726), .A2(n20769), .ZN(n20728) );
  OAI21_X1 U23712 ( .B1(n20728), .B2(n20760), .A(n20727), .ZN(n20736) );
  OR2_X1 U23713 ( .A1(n13553), .A2(n20729), .ZN(n20768) );
  NOR2_X1 U23714 ( .A1(n20768), .A2(n20799), .ZN(n20733) );
  NAND2_X1 U23715 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20845) );
  AOI22_X1 U23716 ( .A1(n20790), .A2(n20859), .B1(n20853), .B2(n10377), .ZN(
        n20740) );
  INV_X1 U23717 ( .A(n20733), .ZN(n20735) );
  AOI22_X1 U23718 ( .A1(n20736), .A2(n20735), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n20734), .ZN(n20737) );
  AOI22_X1 U23719 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n20761), .B1(
        n20760), .B2(n20806), .ZN(n20739) );
  OAI211_X1 U23720 ( .C1(n20765), .C2(n20741), .A(n20740), .B(n20739), .ZN(
        P1_U3129) );
  AOI22_X1 U23721 ( .A1(n20790), .A2(n20865), .B1(n20864), .B2(n10377), .ZN(
        n20743) );
  AOI22_X1 U23722 ( .A1(P1_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n20761), .B1(
        n20760), .B2(n20810), .ZN(n20742) );
  OAI211_X1 U23723 ( .C1(n20765), .C2(n20744), .A(n20743), .B(n20742), .ZN(
        P1_U3130) );
  AOI22_X1 U23724 ( .A1(n20790), .A2(n20871), .B1(n20869), .B2(n10377), .ZN(
        n20746) );
  AOI22_X1 U23725 ( .A1(P1_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n20761), .B1(
        n20760), .B2(n20814), .ZN(n20745) );
  OAI211_X1 U23726 ( .C1(n20765), .C2(n20747), .A(n20746), .B(n20745), .ZN(
        P1_U3131) );
  AOI22_X1 U23727 ( .A1(n20790), .A2(n20877), .B1(n20876), .B2(n10377), .ZN(
        n20749) );
  AOI22_X1 U23728 ( .A1(P1_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n20761), .B1(
        n20760), .B2(n20818), .ZN(n20748) );
  OAI211_X1 U23729 ( .C1(n20765), .C2(n20750), .A(n20749), .B(n20748), .ZN(
        P1_U3132) );
  AOI22_X1 U23730 ( .A1(n20790), .A2(n20883), .B1(n20882), .B2(n10377), .ZN(
        n20752) );
  AOI22_X1 U23731 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n20761), .B1(
        n20760), .B2(n20822), .ZN(n20751) );
  OAI211_X1 U23732 ( .C1(n20765), .C2(n20753), .A(n20752), .B(n20751), .ZN(
        P1_U3133) );
  AOI22_X1 U23733 ( .A1(n20790), .A2(n20889), .B1(n20887), .B2(n10377), .ZN(
        n20755) );
  AOI22_X1 U23734 ( .A1(P1_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n20761), .B1(
        n20760), .B2(n20826), .ZN(n20754) );
  OAI211_X1 U23735 ( .C1(n20765), .C2(n20756), .A(n20755), .B(n20754), .ZN(
        P1_U3134) );
  AOI22_X1 U23736 ( .A1(n20790), .A2(n20895), .B1(n20893), .B2(n10377), .ZN(
        n20758) );
  AOI22_X1 U23737 ( .A1(P1_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n20761), .B1(
        n20760), .B2(n20830), .ZN(n20757) );
  OAI211_X1 U23738 ( .C1(n20765), .C2(n20759), .A(n20758), .B(n20757), .ZN(
        P1_U3135) );
  AOI22_X1 U23739 ( .A1(n20790), .A2(n20903), .B1(n20900), .B2(n10377), .ZN(
        n20763) );
  AOI22_X1 U23740 ( .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n20761), .B1(
        n20760), .B2(n20836), .ZN(n20762) );
  OAI211_X1 U23741 ( .C1(n20765), .C2(n20764), .A(n20763), .B(n20762), .ZN(
        P1_U3136) );
  NOR3_X2 U23742 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20767), .A3(
        n20845), .ZN(n20788) );
  INV_X1 U23743 ( .A(n20788), .ZN(n20771) );
  NOR2_X1 U23744 ( .A1(n20845), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n20772) );
  INV_X1 U23745 ( .A(n20772), .ZN(n20770) );
  INV_X1 U23746 ( .A(n20768), .ZN(n20800) );
  NAND2_X1 U23747 ( .A1(n20800), .A2(n20769), .ZN(n20851) );
  OAI222_X1 U23748 ( .A1(n20771), .A2(n20848), .B1(n20999), .B2(n20770), .C1(
        n20358), .C2(n20851), .ZN(n20789) );
  AOI22_X1 U23749 ( .A1(n20789), .A2(n20852), .B1(n20853), .B2(n20788), .ZN(
        n20775) );
  AOI22_X1 U23750 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n20791), .B1(
        n20790), .B2(n20806), .ZN(n20774) );
  OAI211_X1 U23751 ( .C1(n20809), .C2(n20805), .A(n20775), .B(n20774), .ZN(
        P1_U3137) );
  AOI22_X1 U23752 ( .A1(n20789), .A2(n20863), .B1(n20864), .B2(n20788), .ZN(
        n20777) );
  AOI22_X1 U23753 ( .A1(P1_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n20791), .B1(
        n20790), .B2(n20810), .ZN(n20776) );
  OAI211_X1 U23754 ( .C1(n20813), .C2(n20805), .A(n20777), .B(n20776), .ZN(
        P1_U3138) );
  AOI22_X1 U23755 ( .A1(n20870), .A2(n20789), .B1(n20869), .B2(n20788), .ZN(
        n20779) );
  AOI22_X1 U23756 ( .A1(P1_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n20791), .B1(
        n20790), .B2(n20814), .ZN(n20778) );
  OAI211_X1 U23757 ( .C1(n20817), .C2(n20805), .A(n20779), .B(n20778), .ZN(
        P1_U3139) );
  AOI22_X1 U23758 ( .A1(n20789), .A2(n20875), .B1(n20876), .B2(n20788), .ZN(
        n20781) );
  AOI22_X1 U23759 ( .A1(P1_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n20791), .B1(
        n20790), .B2(n20818), .ZN(n20780) );
  OAI211_X1 U23760 ( .C1(n20821), .C2(n20805), .A(n20781), .B(n20780), .ZN(
        P1_U3140) );
  AOI22_X1 U23761 ( .A1(n20789), .A2(n20881), .B1(n20882), .B2(n20788), .ZN(
        n20783) );
  AOI22_X1 U23762 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n20791), .B1(
        n20790), .B2(n20822), .ZN(n20782) );
  OAI211_X1 U23763 ( .C1(n20825), .C2(n20805), .A(n20783), .B(n20782), .ZN(
        P1_U3141) );
  AOI22_X1 U23764 ( .A1(n20789), .A2(n20888), .B1(n20887), .B2(n20788), .ZN(
        n20785) );
  AOI22_X1 U23765 ( .A1(P1_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n20791), .B1(
        n20790), .B2(n20826), .ZN(n20784) );
  OAI211_X1 U23766 ( .C1(n20829), .C2(n20805), .A(n20785), .B(n20784), .ZN(
        P1_U3142) );
  AOI22_X1 U23767 ( .A1(n20789), .A2(n20894), .B1(n20893), .B2(n20788), .ZN(
        n20787) );
  AOI22_X1 U23768 ( .A1(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n20791), .B1(
        n20790), .B2(n20830), .ZN(n20786) );
  OAI211_X1 U23769 ( .C1(n20833), .C2(n20805), .A(n20787), .B(n20786), .ZN(
        P1_U3143) );
  AOI22_X1 U23770 ( .A1(n20789), .A2(n20902), .B1(n20900), .B2(n20788), .ZN(
        n20793) );
  AOI22_X1 U23771 ( .A1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n20791), .B1(
        n20790), .B2(n20836), .ZN(n20792) );
  OAI211_X1 U23772 ( .C1(n20841), .C2(n20805), .A(n20793), .B(n20792), .ZN(
        P1_U3144) );
  NOR3_X2 U23773 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20846), .A3(
        n20845), .ZN(n20834) );
  OAI22_X1 U23774 ( .A1(n20851), .A2(n13838), .B1(n20797), .B2(n20796), .ZN(
        n20835) );
  AOI22_X1 U23775 ( .A1(n20853), .A2(n20834), .B1(n20852), .B2(n20835), .ZN(
        n20808) );
  AOI21_X1 U23776 ( .B1(n20805), .B2(n20908), .A(n21000), .ZN(n20798) );
  AOI21_X1 U23777 ( .B1(n20800), .B2(n20799), .A(n20798), .ZN(n20801) );
  NOR2_X1 U23778 ( .A1(n20801), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20804) );
  AOI22_X1 U23779 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n20838), .B1(
        n20837), .B2(n20806), .ZN(n20807) );
  OAI211_X1 U23780 ( .C1(n20809), .C2(n20908), .A(n20808), .B(n20807), .ZN(
        P1_U3145) );
  AOI22_X1 U23781 ( .A1(n20864), .A2(n20834), .B1(n20835), .B2(n20863), .ZN(
        n20812) );
  AOI22_X1 U23782 ( .A1(P1_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n20838), .B1(
        n20837), .B2(n20810), .ZN(n20811) );
  OAI211_X1 U23783 ( .C1(n20813), .C2(n20908), .A(n20812), .B(n20811), .ZN(
        P1_U3146) );
  AOI22_X1 U23784 ( .A1(n20870), .A2(n20835), .B1(n20869), .B2(n20834), .ZN(
        n20816) );
  AOI22_X1 U23785 ( .A1(P1_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n20838), .B1(
        n20837), .B2(n20814), .ZN(n20815) );
  OAI211_X1 U23786 ( .C1(n20817), .C2(n20908), .A(n20816), .B(n20815), .ZN(
        P1_U3147) );
  AOI22_X1 U23787 ( .A1(n20876), .A2(n20834), .B1(n20875), .B2(n20835), .ZN(
        n20820) );
  AOI22_X1 U23788 ( .A1(P1_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n20838), .B1(
        n20837), .B2(n20818), .ZN(n20819) );
  OAI211_X1 U23789 ( .C1(n20821), .C2(n20908), .A(n20820), .B(n20819), .ZN(
        P1_U3148) );
  AOI22_X1 U23790 ( .A1(n20882), .A2(n20834), .B1(n20835), .B2(n20881), .ZN(
        n20824) );
  AOI22_X1 U23791 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n20838), .B1(
        n20837), .B2(n20822), .ZN(n20823) );
  OAI211_X1 U23792 ( .C1(n20825), .C2(n20908), .A(n20824), .B(n20823), .ZN(
        P1_U3149) );
  AOI22_X1 U23793 ( .A1(n20888), .A2(n20835), .B1(n20887), .B2(n20834), .ZN(
        n20828) );
  AOI22_X1 U23794 ( .A1(P1_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n20838), .B1(
        n20837), .B2(n20826), .ZN(n20827) );
  OAI211_X1 U23795 ( .C1(n20829), .C2(n20908), .A(n20828), .B(n20827), .ZN(
        P1_U3150) );
  AOI22_X1 U23796 ( .A1(n20894), .A2(n20835), .B1(n20893), .B2(n20834), .ZN(
        n20832) );
  AOI22_X1 U23797 ( .A1(P1_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n20838), .B1(
        n20837), .B2(n20830), .ZN(n20831) );
  OAI211_X1 U23798 ( .C1(n20833), .C2(n20908), .A(n20832), .B(n20831), .ZN(
        P1_U3151) );
  AOI22_X1 U23799 ( .A1(n20902), .A2(n20835), .B1(n20900), .B2(n20834), .ZN(
        n20840) );
  AOI22_X1 U23800 ( .A1(P1_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n20838), .B1(
        n20837), .B2(n20836), .ZN(n20839) );
  OAI211_X1 U23801 ( .C1(n20841), .C2(n20908), .A(n20840), .B(n20839), .ZN(
        P1_U3152) );
  INV_X1 U23802 ( .A(n20845), .ZN(n20842) );
  NAND2_X1 U23803 ( .A1(n20843), .A2(n20842), .ZN(n20847) );
  INV_X1 U23804 ( .A(n20847), .ZN(n20899) );
  INV_X1 U23805 ( .A(n20844), .ZN(n20850) );
  NOR2_X1 U23806 ( .A1(n20846), .A2(n20845), .ZN(n20857) );
  INV_X1 U23807 ( .A(n20857), .ZN(n20849) );
  OAI222_X1 U23808 ( .A1(n20851), .A2(n20850), .B1(n20999), .B2(n20849), .C1(
        n20848), .C2(n20847), .ZN(n20901) );
  AOI22_X1 U23809 ( .A1(n20853), .A2(n20899), .B1(n20852), .B2(n20901), .ZN(
        n20861) );
  NOR2_X1 U23810 ( .A1(n20855), .A2(n20854), .ZN(n20858) );
  AOI22_X1 U23811 ( .A1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n20905), .B1(
        n20904), .B2(n20859), .ZN(n20860) );
  OAI211_X1 U23812 ( .C1(n20862), .C2(n20908), .A(n20861), .B(n20860), .ZN(
        P1_U3153) );
  AOI22_X1 U23813 ( .A1(n20864), .A2(n20899), .B1(n20901), .B2(n20863), .ZN(
        n20867) );
  AOI22_X1 U23814 ( .A1(P1_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n20905), .B1(
        n20904), .B2(n20865), .ZN(n20866) );
  OAI211_X1 U23815 ( .C1(n20868), .C2(n20908), .A(n20867), .B(n20866), .ZN(
        P1_U3154) );
  AOI22_X1 U23816 ( .A1(n20870), .A2(n20901), .B1(n20869), .B2(n20899), .ZN(
        n20873) );
  AOI22_X1 U23817 ( .A1(P1_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n20905), .B1(
        n20904), .B2(n20871), .ZN(n20872) );
  OAI211_X1 U23818 ( .C1(n20874), .C2(n20908), .A(n20873), .B(n20872), .ZN(
        P1_U3155) );
  AOI22_X1 U23819 ( .A1(n20876), .A2(n20899), .B1(n20875), .B2(n20901), .ZN(
        n20879) );
  AOI22_X1 U23820 ( .A1(P1_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n20905), .B1(
        n20904), .B2(n20877), .ZN(n20878) );
  OAI211_X1 U23821 ( .C1(n20880), .C2(n20908), .A(n20879), .B(n20878), .ZN(
        P1_U3156) );
  AOI22_X1 U23822 ( .A1(n20882), .A2(n20899), .B1(n20901), .B2(n20881), .ZN(
        n20885) );
  AOI22_X1 U23823 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n20905), .B1(
        n20904), .B2(n20883), .ZN(n20884) );
  OAI211_X1 U23824 ( .C1(n20886), .C2(n20908), .A(n20885), .B(n20884), .ZN(
        P1_U3157) );
  AOI22_X1 U23825 ( .A1(n20888), .A2(n20901), .B1(n20887), .B2(n20899), .ZN(
        n20891) );
  AOI22_X1 U23826 ( .A1(P1_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n20905), .B1(
        n20904), .B2(n20889), .ZN(n20890) );
  OAI211_X1 U23827 ( .C1(n20892), .C2(n20908), .A(n20891), .B(n20890), .ZN(
        P1_U3158) );
  AOI22_X1 U23828 ( .A1(n20894), .A2(n20901), .B1(n20893), .B2(n20899), .ZN(
        n20897) );
  AOI22_X1 U23829 ( .A1(P1_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n20905), .B1(
        n20904), .B2(n20895), .ZN(n20896) );
  OAI211_X1 U23830 ( .C1(n20898), .C2(n20908), .A(n20897), .B(n20896), .ZN(
        P1_U3159) );
  AOI22_X1 U23831 ( .A1(n20902), .A2(n20901), .B1(n20900), .B2(n20899), .ZN(
        n20907) );
  AOI22_X1 U23832 ( .A1(P1_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n20905), .B1(
        n20904), .B2(n20903), .ZN(n20906) );
  OAI211_X1 U23833 ( .C1(n20909), .C2(n20908), .A(n20907), .B(n20906), .ZN(
        P1_U3160) );
  OAI211_X1 U23834 ( .C1(n20912), .C2(n20999), .A(n20911), .B(n20910), .ZN(
        P1_U3163) );
  INV_X1 U23835 ( .A(n20989), .ZN(n20985) );
  AND2_X1 U23836 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n20985), .ZN(
        P1_U3164) );
  AND2_X1 U23837 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n20985), .ZN(
        P1_U3165) );
  AND2_X1 U23838 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n20985), .ZN(
        P1_U3166) );
  AND2_X1 U23839 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n20985), .ZN(
        P1_U3167) );
  AND2_X1 U23840 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n20985), .ZN(
        P1_U3168) );
  AND2_X1 U23841 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n20985), .ZN(
        P1_U3169) );
  AND2_X1 U23842 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n20985), .ZN(
        P1_U3170) );
  AND2_X1 U23843 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n20985), .ZN(
        P1_U3171) );
  AND2_X1 U23844 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n20985), .ZN(
        P1_U3172) );
  AND2_X1 U23845 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n20985), .ZN(
        P1_U3173) );
  AND2_X1 U23846 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n20985), .ZN(
        P1_U3174) );
  AND2_X1 U23847 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n20985), .ZN(
        P1_U3175) );
  AND2_X1 U23848 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n20985), .ZN(
        P1_U3176) );
  AND2_X1 U23849 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n20985), .ZN(
        P1_U3177) );
  AND2_X1 U23850 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n20985), .ZN(
        P1_U3178) );
  AND2_X1 U23851 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n20985), .ZN(
        P1_U3179) );
  AND2_X1 U23852 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n20985), .ZN(
        P1_U3180) );
  AND2_X1 U23853 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n20985), .ZN(
        P1_U3181) );
  AND2_X1 U23854 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(n20985), .ZN(
        P1_U3182) );
  AND2_X1 U23855 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n20985), .ZN(
        P1_U3183) );
  AND2_X1 U23856 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(n20985), .ZN(
        P1_U3184) );
  AND2_X1 U23857 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n20985), .ZN(
        P1_U3185) );
  AND2_X1 U23858 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n20985), .ZN(P1_U3186) );
  AND2_X1 U23859 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n20985), .ZN(P1_U3187) );
  AND2_X1 U23860 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n20985), .ZN(P1_U3188) );
  AND2_X1 U23861 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n20985), .ZN(P1_U3189) );
  AND2_X1 U23862 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n20985), .ZN(P1_U3190) );
  AND2_X1 U23863 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n20985), .ZN(P1_U3191) );
  AND2_X1 U23864 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n20985), .ZN(P1_U3192) );
  AND2_X1 U23865 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n20985), .ZN(P1_U3193) );
  NAND2_X1 U23866 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n20913), .ZN(n20923) );
  INV_X1 U23867 ( .A(n20923), .ZN(n20917) );
  OAI21_X1 U23868 ( .B1(P1_STATE_REG_0__SCAN_IN), .B2(n20924), .A(
        P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n20914) );
  AOI211_X1 U23869 ( .C1(HOLD), .C2(P1_STATE_REG_1__SCAN_IN), .A(n20915), .B(
        n20914), .ZN(n20916) );
  OAI22_X1 U23870 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20917), .B1(n21013), 
        .B2(n20916), .ZN(P1_U3194) );
  AOI21_X1 U23871 ( .B1(n20919), .B2(n20924), .A(n20918), .ZN(n20927) );
  AOI21_X1 U23872 ( .B1(P1_REQUESTPENDING_REG_SCAN_IN), .B2(n20928), .A(n20920), .ZN(n20922) );
  OAI221_X1 U23873 ( .B1(n20922), .B2(P1_REQUESTPENDING_REG_SCAN_IN), .C1(
        n20922), .C2(n20921), .A(P1_STATE_REG_0__SCAN_IN), .ZN(n20926) );
  OAI211_X1 U23874 ( .C1(P1_STATE_REG_1__SCAN_IN), .C2(n20924), .A(
        P1_STATE_REG_2__SCAN_IN), .B(n20923), .ZN(n20925) );
  OAI21_X1 U23875 ( .B1(n20927), .B2(n20926), .A(n20925), .ZN(P1_U3196) );
  NAND2_X1 U23876 ( .A1(n21013), .A2(n20928), .ZN(n20973) );
  INV_X1 U23877 ( .A(P1_ADDRESS_REG_0__SCAN_IN), .ZN(n20929) );
  OAI222_X1 U23878 ( .A1(n20973), .A2(n13929), .B1(n20929), .B2(n21013), .C1(
        n13576), .C2(n20970), .ZN(P1_U3197) );
  INV_X1 U23879 ( .A(P1_ADDRESS_REG_1__SCAN_IN), .ZN(n20930) );
  OAI222_X1 U23880 ( .A1(n20970), .A2(n13929), .B1(n20930), .B2(n21013), .C1(
        n20932), .C2(n20973), .ZN(P1_U3198) );
  OAI222_X1 U23881 ( .A1(n20970), .A2(n20932), .B1(n20931), .B2(n21013), .C1(
        n20933), .C2(n20973), .ZN(P1_U3199) );
  INV_X1 U23882 ( .A(P1_ADDRESS_REG_3__SCAN_IN), .ZN(n21172) );
  OAI222_X1 U23883 ( .A1(n20973), .A2(n20935), .B1(n21172), .B2(n21013), .C1(
        n20933), .C2(n20970), .ZN(P1_U3200) );
  INV_X1 U23884 ( .A(P1_ADDRESS_REG_4__SCAN_IN), .ZN(n20934) );
  OAI222_X1 U23885 ( .A1(n20970), .A2(n20935), .B1(n20934), .B2(n21013), .C1(
        n21198), .C2(n20973), .ZN(P1_U3201) );
  INV_X1 U23886 ( .A(n20973), .ZN(n20976) );
  AOI22_X1 U23887 ( .A1(P1_ADDRESS_REG_5__SCAN_IN), .A2(n20997), .B1(
        P1_REIP_REG_7__SCAN_IN), .B2(n20976), .ZN(n20936) );
  OAI21_X1 U23888 ( .B1(n21198), .B2(n20970), .A(n20936), .ZN(P1_U3202) );
  AOI22_X1 U23889 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(n20997), .B1(
        P1_REIP_REG_7__SCAN_IN), .B2(n20977), .ZN(n20937) );
  OAI21_X1 U23890 ( .B1(n21260), .B2(n20973), .A(n20937), .ZN(P1_U3203) );
  INV_X1 U23891 ( .A(P1_ADDRESS_REG_7__SCAN_IN), .ZN(n20938) );
  OAI222_X1 U23892 ( .A1(n20973), .A2(n20940), .B1(n20938), .B2(n21013), .C1(
        n21260), .C2(n20970), .ZN(P1_U3204) );
  INV_X1 U23893 ( .A(P1_ADDRESS_REG_8__SCAN_IN), .ZN(n20939) );
  OAI222_X1 U23894 ( .A1(n20970), .A2(n20940), .B1(n20939), .B2(n21013), .C1(
        n20942), .C2(n20973), .ZN(P1_U3205) );
  INV_X1 U23895 ( .A(P1_ADDRESS_REG_9__SCAN_IN), .ZN(n20941) );
  INV_X1 U23896 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n21231) );
  OAI222_X1 U23897 ( .A1(n20970), .A2(n20942), .B1(n20941), .B2(n21013), .C1(
        n21231), .C2(n20973), .ZN(P1_U3206) );
  INV_X1 U23898 ( .A(P1_ADDRESS_REG_10__SCAN_IN), .ZN(n20943) );
  OAI222_X1 U23899 ( .A1(n20970), .A2(n21231), .B1(n20943), .B2(n21013), .C1(
        n20944), .C2(n20973), .ZN(P1_U3207) );
  INV_X1 U23900 ( .A(P1_ADDRESS_REG_11__SCAN_IN), .ZN(n20945) );
  OAI222_X1 U23901 ( .A1(n20973), .A2(n20947), .B1(n20945), .B2(n21013), .C1(
        n20944), .C2(n20970), .ZN(P1_U3208) );
  AOI22_X1 U23902 ( .A1(P1_ADDRESS_REG_12__SCAN_IN), .A2(n20997), .B1(
        P1_REIP_REG_14__SCAN_IN), .B2(n20976), .ZN(n20946) );
  OAI21_X1 U23903 ( .B1(n20947), .B2(n20970), .A(n20946), .ZN(P1_U3209) );
  INV_X1 U23904 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n20950) );
  AOI22_X1 U23905 ( .A1(P1_ADDRESS_REG_13__SCAN_IN), .A2(n20997), .B1(
        P1_REIP_REG_14__SCAN_IN), .B2(n20977), .ZN(n20948) );
  OAI21_X1 U23906 ( .B1(n20950), .B2(n20973), .A(n20948), .ZN(P1_U3210) );
  AOI22_X1 U23907 ( .A1(P1_ADDRESS_REG_14__SCAN_IN), .A2(n20997), .B1(
        P1_REIP_REG_16__SCAN_IN), .B2(n20976), .ZN(n20949) );
  OAI21_X1 U23908 ( .B1(n20950), .B2(n20970), .A(n20949), .ZN(P1_U3211) );
  AOI22_X1 U23909 ( .A1(P1_ADDRESS_REG_15__SCAN_IN), .A2(n20997), .B1(
        P1_REIP_REG_16__SCAN_IN), .B2(n20977), .ZN(n20951) );
  OAI21_X1 U23910 ( .B1(n20952), .B2(n20973), .A(n20951), .ZN(P1_U3212) );
  INV_X1 U23911 ( .A(P1_ADDRESS_REG_16__SCAN_IN), .ZN(n20953) );
  OAI222_X1 U23912 ( .A1(n20973), .A2(n20955), .B1(n20953), .B2(n21013), .C1(
        n20952), .C2(n20970), .ZN(P1_U3213) );
  INV_X1 U23913 ( .A(P1_ADDRESS_REG_17__SCAN_IN), .ZN(n20954) );
  OAI222_X1 U23914 ( .A1(n20970), .A2(n20955), .B1(n20954), .B2(n21013), .C1(
        n20957), .C2(n20973), .ZN(P1_U3214) );
  INV_X1 U23915 ( .A(P1_ADDRESS_REG_18__SCAN_IN), .ZN(n20956) );
  OAI222_X1 U23916 ( .A1(n20970), .A2(n20957), .B1(n20956), .B2(n21013), .C1(
        n20959), .C2(n20973), .ZN(P1_U3215) );
  AOI22_X1 U23917 ( .A1(P1_ADDRESS_REG_19__SCAN_IN), .A2(n20997), .B1(
        P1_REIP_REG_21__SCAN_IN), .B2(n20976), .ZN(n20958) );
  OAI21_X1 U23918 ( .B1(n20959), .B2(n20970), .A(n20958), .ZN(P1_U3216) );
  AOI22_X1 U23919 ( .A1(P1_ADDRESS_REG_20__SCAN_IN), .A2(n20997), .B1(
        P1_REIP_REG_21__SCAN_IN), .B2(n20977), .ZN(n20960) );
  OAI21_X1 U23920 ( .B1(n20962), .B2(n20973), .A(n20960), .ZN(P1_U3217) );
  AOI22_X1 U23921 ( .A1(P1_ADDRESS_REG_21__SCAN_IN), .A2(n20997), .B1(
        P1_REIP_REG_23__SCAN_IN), .B2(n20976), .ZN(n20961) );
  OAI21_X1 U23922 ( .B1(n20962), .B2(n20970), .A(n20961), .ZN(P1_U3218) );
  AOI22_X1 U23923 ( .A1(P1_ADDRESS_REG_22__SCAN_IN), .A2(n20997), .B1(
        P1_REIP_REG_23__SCAN_IN), .B2(n20977), .ZN(n20963) );
  OAI21_X1 U23924 ( .B1(n20965), .B2(n20973), .A(n20963), .ZN(P1_U3219) );
  AOI22_X1 U23925 ( .A1(P1_REIP_REG_25__SCAN_IN), .A2(n20976), .B1(
        P1_ADDRESS_REG_23__SCAN_IN), .B2(n20997), .ZN(n20964) );
  OAI21_X1 U23926 ( .B1(n20965), .B2(n20970), .A(n20964), .ZN(P1_U3220) );
  AOI22_X1 U23927 ( .A1(P1_REIP_REG_25__SCAN_IN), .A2(n20977), .B1(
        P1_ADDRESS_REG_24__SCAN_IN), .B2(n20997), .ZN(n20966) );
  OAI21_X1 U23928 ( .B1(n20968), .B2(n20973), .A(n20966), .ZN(P1_U3221) );
  INV_X1 U23929 ( .A(P1_ADDRESS_REG_25__SCAN_IN), .ZN(n20967) );
  OAI222_X1 U23930 ( .A1(n20970), .A2(n20968), .B1(n20967), .B2(n21013), .C1(
        n20971), .C2(n20973), .ZN(P1_U3222) );
  AOI22_X1 U23931 ( .A1(P1_REIP_REG_28__SCAN_IN), .A2(n20976), .B1(
        P1_ADDRESS_REG_26__SCAN_IN), .B2(n20997), .ZN(n20969) );
  OAI21_X1 U23932 ( .B1(n20971), .B2(n20970), .A(n20969), .ZN(P1_U3223) );
  AOI22_X1 U23933 ( .A1(P1_REIP_REG_28__SCAN_IN), .A2(n20977), .B1(
        P1_ADDRESS_REG_27__SCAN_IN), .B2(n20997), .ZN(n20972) );
  OAI21_X1 U23934 ( .B1(n20974), .B2(n20973), .A(n20972), .ZN(P1_U3224) );
  AOI222_X1 U23935 ( .A1(n20976), .A2(P1_REIP_REG_30__SCAN_IN), .B1(
        P1_ADDRESS_REG_28__SCAN_IN), .B2(n20997), .C1(P1_REIP_REG_29__SCAN_IN), 
        .C2(n20977), .ZN(n20975) );
  INV_X1 U23936 ( .A(n20975), .ZN(P1_U3225) );
  AOI222_X1 U23937 ( .A1(n20977), .A2(P1_REIP_REG_30__SCAN_IN), .B1(
        P1_ADDRESS_REG_29__SCAN_IN), .B2(n20997), .C1(P1_REIP_REG_31__SCAN_IN), 
        .C2(n20976), .ZN(n20978) );
  INV_X1 U23938 ( .A(n20978), .ZN(P1_U3226) );
  INV_X1 U23939 ( .A(P1_BE_N_REG_3__SCAN_IN), .ZN(n20979) );
  AOI22_X1 U23940 ( .A1(n21013), .A2(n20980), .B1(n20979), .B2(n20997), .ZN(
        P1_U3458) );
  INV_X1 U23941 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n20992) );
  INV_X1 U23942 ( .A(P1_BE_N_REG_2__SCAN_IN), .ZN(n21290) );
  AOI22_X1 U23943 ( .A1(n21013), .A2(n20992), .B1(n21290), .B2(n20997), .ZN(
        P1_U3459) );
  INV_X1 U23944 ( .A(P1_BE_N_REG_1__SCAN_IN), .ZN(n20981) );
  AOI22_X1 U23945 ( .A1(n21013), .A2(n20982), .B1(n20981), .B2(n20997), .ZN(
        P1_U3460) );
  INV_X1 U23946 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n20995) );
  INV_X1 U23947 ( .A(P1_BE_N_REG_0__SCAN_IN), .ZN(n20983) );
  AOI22_X1 U23948 ( .A1(n21013), .A2(n20995), .B1(n20983), .B2(n20997), .ZN(
        P1_U3461) );
  INV_X1 U23949 ( .A(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(n20986) );
  INV_X1 U23950 ( .A(n20987), .ZN(n20984) );
  AOI21_X1 U23951 ( .B1(n20986), .B2(n20985), .A(n20984), .ZN(P1_U3464) );
  OAI21_X1 U23952 ( .B1(n20989), .B2(n20988), .A(n20987), .ZN(P1_U3465) );
  AOI21_X1 U23953 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n20990) );
  AOI22_X1 U23954 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_0__SCAN_IN), 
        .B1(n20990), .B2(n13576), .ZN(n20993) );
  AOI22_X1 U23955 ( .A1(n20996), .A2(n20993), .B1(n20992), .B2(n20991), .ZN(
        P1_U3481) );
  OAI21_X1 U23956 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(P1_REIP_REG_0__SCAN_IN), 
        .A(n20996), .ZN(n20994) );
  OAI21_X1 U23957 ( .B1(n20996), .B2(n20995), .A(n20994), .ZN(P1_U3482) );
  AOI22_X1 U23958 ( .A1(n21013), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n20998), 
        .B2(n20997), .ZN(P1_U3483) );
  AOI21_X1 U23959 ( .B1(n21001), .B2(n21000), .A(n20999), .ZN(n21006) );
  INV_X1 U23960 ( .A(n21002), .ZN(n21003) );
  NAND2_X1 U23961 ( .A1(n21004), .A2(n21003), .ZN(n21005) );
  AOI21_X1 U23962 ( .B1(n21007), .B2(n21006), .A(n21005), .ZN(n21012) );
  AOI211_X1 U23963 ( .C1(n13910), .C2(n21010), .A(n21009), .B(n21008), .ZN(
        n21011) );
  MUX2_X1 U23964 ( .A(n21012), .B(P1_REQUESTPENDING_REG_SCAN_IN), .S(n21011), 
        .Z(P1_U3485) );
  MUX2_X1 U23965 ( .A(P1_M_IO_N_REG_SCAN_IN), .B(P1_MEMORYFETCH_REG_SCAN_IN), 
        .S(n21013), .Z(P1_U3486) );
  AOI22_X1 U23966 ( .A1(P1_BE_N_REG_2__SCAN_IN), .A2(keyinput195), .B1(
        P3_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(keyinput234), .ZN(n21014) );
  OAI221_X1 U23967 ( .B1(P1_BE_N_REG_2__SCAN_IN), .B2(keyinput195), .C1(
        P3_PHYADDRPOINTER_REG_14__SCAN_IN), .C2(keyinput234), .A(n21014), .ZN(
        n21021) );
  AOI22_X1 U23968 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(keyinput146), 
        .B1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B2(keyinput230), .ZN(n21015) );
  OAI221_X1 U23969 ( .B1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B2(keyinput146), 
        .C1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .C2(keyinput230), .A(n21015), 
        .ZN(n21020) );
  AOI22_X1 U23970 ( .A1(P2_EAX_REG_29__SCAN_IN), .A2(keyinput244), .B1(
        P2_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(keyinput157), .ZN(n21016) );
  OAI221_X1 U23971 ( .B1(P2_EAX_REG_29__SCAN_IN), .B2(keyinput244), .C1(
        P2_INSTADDRPOINTER_REG_14__SCAN_IN), .C2(keyinput157), .A(n21016), 
        .ZN(n21019) );
  AOI22_X1 U23972 ( .A1(P3_EAX_REG_26__SCAN_IN), .A2(keyinput247), .B1(
        P1_EAX_REG_16__SCAN_IN), .B2(keyinput148), .ZN(n21017) );
  OAI221_X1 U23973 ( .B1(P3_EAX_REG_26__SCAN_IN), .B2(keyinput247), .C1(
        P1_EAX_REG_16__SCAN_IN), .C2(keyinput148), .A(n21017), .ZN(n21018) );
  NOR4_X1 U23974 ( .A1(n21021), .A2(n21020), .A3(n21019), .A4(n21018), .ZN(
        n21049) );
  AOI22_X1 U23975 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(keyinput179), 
        .B1(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B2(keyinput173), .ZN(n21022) );
  OAI221_X1 U23976 ( .B1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(keyinput179), 
        .C1(P1_INSTQUEUE_REG_6__7__SCAN_IN), .C2(keyinput173), .A(n21022), 
        .ZN(n21029) );
  AOI22_X1 U23977 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(keyinput245), .B1(
        P1_REIP_REG_11__SCAN_IN), .B2(keyinput203), .ZN(n21023) );
  OAI221_X1 U23978 ( .B1(P3_EAX_REG_12__SCAN_IN), .B2(keyinput245), .C1(
        P1_REIP_REG_11__SCAN_IN), .C2(keyinput203), .A(n21023), .ZN(n21028) );
  AOI22_X1 U23979 ( .A1(P3_UWORD_REG_4__SCAN_IN), .A2(keyinput233), .B1(
        P3_INSTQUEUE_REG_7__3__SCAN_IN), .B2(keyinput155), .ZN(n21024) );
  OAI221_X1 U23980 ( .B1(P3_UWORD_REG_4__SCAN_IN), .B2(keyinput233), .C1(
        P3_INSTQUEUE_REG_7__3__SCAN_IN), .C2(keyinput155), .A(n21024), .ZN(
        n21027) );
  AOI22_X1 U23981 ( .A1(DATAI_31_), .A2(keyinput172), .B1(
        P2_INSTQUEUE_REG_14__3__SCAN_IN), .B2(keyinput215), .ZN(n21025) );
  OAI221_X1 U23982 ( .B1(DATAI_31_), .B2(keyinput172), .C1(
        P2_INSTQUEUE_REG_14__3__SCAN_IN), .C2(keyinput215), .A(n21025), .ZN(
        n21026) );
  NOR4_X1 U23983 ( .A1(n21029), .A2(n21028), .A3(n21027), .A4(n21026), .ZN(
        n21048) );
  AOI22_X1 U23984 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(keyinput168), 
        .B1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B2(keyinput130), .ZN(n21030) );
  OAI221_X1 U23985 ( .B1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(keyinput168), 
        .C1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .C2(keyinput130), .A(n21030), 
        .ZN(n21037) );
  AOI22_X1 U23986 ( .A1(P3_ADDRESS_REG_22__SCAN_IN), .A2(keyinput196), .B1(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(keyinput137), .ZN(n21031) );
  OAI221_X1 U23987 ( .B1(P3_ADDRESS_REG_22__SCAN_IN), .B2(keyinput196), .C1(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .C2(keyinput137), .A(n21031), 
        .ZN(n21036) );
  AOI22_X1 U23988 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(keyinput199), .B1(
        P2_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(keyinput221), .ZN(n21032) );
  OAI221_X1 U23989 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(keyinput199), .C1(
        P2_INSTADDRPOINTER_REG_23__SCAN_IN), .C2(keyinput221), .A(n21032), 
        .ZN(n21035) );
  AOI22_X1 U23990 ( .A1(DATAI_0_), .A2(keyinput235), .B1(
        P2_INSTQUEUE_REG_15__5__SCAN_IN), .B2(keyinput189), .ZN(n21033) );
  OAI221_X1 U23991 ( .B1(DATAI_0_), .B2(keyinput235), .C1(
        P2_INSTQUEUE_REG_15__5__SCAN_IN), .C2(keyinput189), .A(n21033), .ZN(
        n21034) );
  NOR4_X1 U23992 ( .A1(n21037), .A2(n21036), .A3(n21035), .A4(n21034), .ZN(
        n21047) );
  AOI22_X1 U23993 ( .A1(P3_EBX_REG_30__SCAN_IN), .A2(keyinput131), .B1(
        P2_INSTQUEUE_REG_1__4__SCAN_IN), .B2(keyinput153), .ZN(n21038) );
  OAI221_X1 U23994 ( .B1(P3_EBX_REG_30__SCAN_IN), .B2(keyinput131), .C1(
        P2_INSTQUEUE_REG_1__4__SCAN_IN), .C2(keyinput153), .A(n21038), .ZN(
        n21045) );
  AOI22_X1 U23995 ( .A1(P2_DATAWIDTH_REG_1__SCAN_IN), .A2(keyinput211), .B1(
        P2_INSTQUEUE_REG_8__2__SCAN_IN), .B2(keyinput198), .ZN(n21039) );
  OAI221_X1 U23996 ( .B1(P2_DATAWIDTH_REG_1__SCAN_IN), .B2(keyinput211), .C1(
        P2_INSTQUEUE_REG_8__2__SCAN_IN), .C2(keyinput198), .A(n21039), .ZN(
        n21044) );
  AOI22_X1 U23997 ( .A1(DATAI_2_), .A2(keyinput178), .B1(
        P1_INSTQUEUE_REG_13__3__SCAN_IN), .B2(keyinput143), .ZN(n21040) );
  OAI221_X1 U23998 ( .B1(DATAI_2_), .B2(keyinput178), .C1(
        P1_INSTQUEUE_REG_13__3__SCAN_IN), .C2(keyinput143), .A(n21040), .ZN(
        n21043) );
  AOI22_X1 U23999 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(keyinput150), 
        .B1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B2(keyinput142), .ZN(n21041) );
  OAI221_X1 U24000 ( .B1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B2(keyinput150), 
        .C1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .C2(keyinput142), .A(n21041), 
        .ZN(n21042) );
  NOR4_X1 U24001 ( .A1(n21045), .A2(n21044), .A3(n21043), .A4(n21042), .ZN(
        n21046) );
  NAND4_X1 U24002 ( .A1(n21049), .A2(n21048), .A3(n21047), .A4(n21046), .ZN(
        n21187) );
  AOI22_X1 U24003 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(keyinput152), 
        .B1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B2(keyinput133), .ZN(n21050) );
  OAI221_X1 U24004 ( .B1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B2(keyinput152), 
        .C1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .C2(keyinput133), .A(n21050), 
        .ZN(n21057) );
  AOI22_X1 U24005 ( .A1(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(keyinput186), 
        .B1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B2(keyinput141), .ZN(n21051) );
  OAI221_X1 U24006 ( .B1(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(keyinput186), 
        .C1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .C2(keyinput141), .A(n21051), 
        .ZN(n21056) );
  AOI22_X1 U24007 ( .A1(P2_LWORD_REG_15__SCAN_IN), .A2(keyinput176), .B1(
        P2_ADDRESS_REG_10__SCAN_IN), .B2(keyinput212), .ZN(n21052) );
  OAI221_X1 U24008 ( .B1(P2_LWORD_REG_15__SCAN_IN), .B2(keyinput176), .C1(
        P2_ADDRESS_REG_10__SCAN_IN), .C2(keyinput212), .A(n21052), .ZN(n21055)
         );
  AOI22_X1 U24009 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(keyinput208), .B1(
        P1_INSTQUEUE_REG_7__1__SCAN_IN), .B2(keyinput238), .ZN(n21053) );
  OAI221_X1 U24010 ( .B1(P1_REIP_REG_8__SCAN_IN), .B2(keyinput208), .C1(
        P1_INSTQUEUE_REG_7__1__SCAN_IN), .C2(keyinput238), .A(n21053), .ZN(
        n21054) );
  NOR4_X1 U24011 ( .A1(n21057), .A2(n21056), .A3(n21055), .A4(n21054), .ZN(
        n21085) );
  AOI22_X1 U24012 ( .A1(P3_EAX_REG_1__SCAN_IN), .A2(keyinput252), .B1(
        P2_EAX_REG_10__SCAN_IN), .B2(keyinput197), .ZN(n21058) );
  OAI221_X1 U24013 ( .B1(P3_EAX_REG_1__SCAN_IN), .B2(keyinput252), .C1(
        P2_EAX_REG_10__SCAN_IN), .C2(keyinput197), .A(n21058), .ZN(n21065) );
  AOI22_X1 U24014 ( .A1(BUF1_REG_18__SCAN_IN), .A2(keyinput167), .B1(
        P2_INSTQUEUE_REG_4__2__SCAN_IN), .B2(keyinput194), .ZN(n21059) );
  OAI221_X1 U24015 ( .B1(BUF1_REG_18__SCAN_IN), .B2(keyinput167), .C1(
        P2_INSTQUEUE_REG_4__2__SCAN_IN), .C2(keyinput194), .A(n21059), .ZN(
        n21064) );
  AOI22_X1 U24016 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(keyinput202), 
        .B1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B2(keyinput213), .ZN(n21060) );
  OAI221_X1 U24017 ( .B1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B2(keyinput202), 
        .C1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .C2(keyinput213), .A(n21060), 
        .ZN(n21063) );
  AOI22_X1 U24018 ( .A1(P2_UWORD_REG_0__SCAN_IN), .A2(keyinput181), .B1(
        P2_REIP_REG_14__SCAN_IN), .B2(keyinput239), .ZN(n21061) );
  OAI221_X1 U24019 ( .B1(P2_UWORD_REG_0__SCAN_IN), .B2(keyinput181), .C1(
        P2_REIP_REG_14__SCAN_IN), .C2(keyinput239), .A(n21061), .ZN(n21062) );
  NOR4_X1 U24020 ( .A1(n21065), .A2(n21064), .A3(n21063), .A4(n21062), .ZN(
        n21084) );
  AOI22_X1 U24021 ( .A1(P3_CODEFETCH_REG_SCAN_IN), .A2(keyinput228), .B1(
        P3_EBX_REG_3__SCAN_IN), .B2(keyinput255), .ZN(n21066) );
  OAI221_X1 U24022 ( .B1(P3_CODEFETCH_REG_SCAN_IN), .B2(keyinput228), .C1(
        P3_EBX_REG_3__SCAN_IN), .C2(keyinput255), .A(n21066), .ZN(n21073) );
  AOI22_X1 U24023 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(keyinput249), .B1(
        P2_LWORD_REG_10__SCAN_IN), .B2(keyinput175), .ZN(n21067) );
  OAI221_X1 U24024 ( .B1(P3_DATAWIDTH_REG_6__SCAN_IN), .B2(keyinput249), .C1(
        P2_LWORD_REG_10__SCAN_IN), .C2(keyinput175), .A(n21067), .ZN(n21072)
         );
  AOI22_X1 U24025 ( .A1(P1_LWORD_REG_0__SCAN_IN), .A2(keyinput251), .B1(
        P3_REIP_REG_14__SCAN_IN), .B2(keyinput226), .ZN(n21068) );
  OAI221_X1 U24026 ( .B1(P1_LWORD_REG_0__SCAN_IN), .B2(keyinput251), .C1(
        P3_REIP_REG_14__SCAN_IN), .C2(keyinput226), .A(n21068), .ZN(n21071) );
  AOI22_X1 U24027 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(keyinput184), 
        .B1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B2(keyinput174), .ZN(n21069) );
  OAI221_X1 U24028 ( .B1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B2(keyinput184), 
        .C1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .C2(keyinput174), .A(n21069), 
        .ZN(n21070) );
  NOR4_X1 U24029 ( .A1(n21073), .A2(n21072), .A3(n21071), .A4(n21070), .ZN(
        n21083) );
  AOI22_X1 U24030 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(keyinput149), .B1(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .B2(keyinput128), .ZN(n21074) );
  OAI221_X1 U24031 ( .B1(P2_DATAWIDTH_REG_8__SCAN_IN), .B2(keyinput149), .C1(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .C2(keyinput128), .A(n21074), 
        .ZN(n21081) );
  AOI22_X1 U24032 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(keyinput163), .B1(
        P3_EAX_REG_7__SCAN_IN), .B2(keyinput253), .ZN(n21075) );
  OAI221_X1 U24033 ( .B1(P3_EAX_REG_13__SCAN_IN), .B2(keyinput163), .C1(
        P3_EAX_REG_7__SCAN_IN), .C2(keyinput253), .A(n21075), .ZN(n21080) );
  AOI22_X1 U24034 ( .A1(P1_DATAO_REG_12__SCAN_IN), .A2(keyinput225), .B1(
        P1_REIP_REG_29__SCAN_IN), .B2(keyinput232), .ZN(n21076) );
  OAI221_X1 U24035 ( .B1(P1_DATAO_REG_12__SCAN_IN), .B2(keyinput225), .C1(
        P1_REIP_REG_29__SCAN_IN), .C2(keyinput232), .A(n21076), .ZN(n21079) );
  AOI22_X1 U24036 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(keyinput229), 
        .B1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B2(keyinput187), .ZN(n21077) );
  OAI221_X1 U24037 ( .B1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B2(keyinput229), 
        .C1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .C2(keyinput187), .A(n21077), 
        .ZN(n21078) );
  NOR4_X1 U24038 ( .A1(n21081), .A2(n21080), .A3(n21079), .A4(n21078), .ZN(
        n21082) );
  NAND4_X1 U24039 ( .A1(n21085), .A2(n21084), .A3(n21083), .A4(n21082), .ZN(
        n21186) );
  AOI22_X1 U24040 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(keyinput188), 
        .B1(n21285), .B2(keyinput151), .ZN(n21086) );
  OAI221_X1 U24041 ( .B1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B2(keyinput188), 
        .C1(n21285), .C2(keyinput151), .A(n21086), .ZN(n21097) );
  AOI22_X1 U24042 ( .A1(n21299), .A2(keyinput209), .B1(keyinput158), .B2(
        n21277), .ZN(n21087) );
  OAI221_X1 U24043 ( .B1(n21299), .B2(keyinput209), .C1(n21277), .C2(
        keyinput158), .A(n21087), .ZN(n21096) );
  AOI22_X1 U24044 ( .A1(n21090), .A2(keyinput250), .B1(n21089), .B2(
        keyinput185), .ZN(n21088) );
  OAI221_X1 U24045 ( .B1(n21090), .B2(keyinput250), .C1(n21089), .C2(
        keyinput185), .A(n21088), .ZN(n21095) );
  AOI22_X1 U24046 ( .A1(n21093), .A2(keyinput210), .B1(n21092), .B2(
        keyinput237), .ZN(n21091) );
  OAI221_X1 U24047 ( .B1(n21093), .B2(keyinput210), .C1(n21092), .C2(
        keyinput237), .A(n21091), .ZN(n21094) );
  NOR4_X1 U24048 ( .A1(n21097), .A2(n21096), .A3(n21095), .A4(n21094), .ZN(
        n21136) );
  INV_X1 U24049 ( .A(P3_DATAO_REG_26__SCAN_IN), .ZN(n21287) );
  AOI22_X1 U24050 ( .A1(n21196), .A2(keyinput164), .B1(keyinput227), .B2(
        n21287), .ZN(n21098) );
  OAI221_X1 U24051 ( .B1(n21196), .B2(keyinput164), .C1(n21287), .C2(
        keyinput227), .A(n21098), .ZN(n21107) );
  INV_X1 U24052 ( .A(DATAI_22_), .ZN(n21100) );
  AOI22_X1 U24053 ( .A1(n21101), .A2(keyinput159), .B1(keyinput135), .B2(
        n21100), .ZN(n21099) );
  OAI221_X1 U24054 ( .B1(n21101), .B2(keyinput159), .C1(n21100), .C2(
        keyinput135), .A(n21099), .ZN(n21106) );
  INV_X1 U24055 ( .A(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n21230) );
  AOI22_X1 U24056 ( .A1(n21289), .A2(keyinput248), .B1(n21230), .B2(
        keyinput217), .ZN(n21102) );
  OAI221_X1 U24057 ( .B1(n21289), .B2(keyinput248), .C1(n21230), .C2(
        keyinput217), .A(n21102), .ZN(n21105) );
  AOI22_X1 U24058 ( .A1(n21274), .A2(keyinput139), .B1(n21198), .B2(
        keyinput136), .ZN(n21103) );
  OAI221_X1 U24059 ( .B1(n21274), .B2(keyinput139), .C1(n21198), .C2(
        keyinput136), .A(n21103), .ZN(n21104) );
  NOR4_X1 U24060 ( .A1(n21107), .A2(n21106), .A3(n21105), .A4(n21104), .ZN(
        n21135) );
  AOI22_X1 U24061 ( .A1(n13022), .A2(keyinput134), .B1(keyinput166), .B2(
        n21109), .ZN(n21108) );
  OAI221_X1 U24062 ( .B1(n13022), .B2(keyinput134), .C1(n21109), .C2(
        keyinput166), .A(n21108), .ZN(n21119) );
  INV_X1 U24063 ( .A(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n21111) );
  AOI22_X1 U24064 ( .A1(n21195), .A2(keyinput140), .B1(keyinput240), .B2(
        n21111), .ZN(n21110) );
  OAI221_X1 U24065 ( .B1(n21195), .B2(keyinput140), .C1(n21111), .C2(
        keyinput240), .A(n21110), .ZN(n21118) );
  INV_X1 U24066 ( .A(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n21113) );
  AOI22_X1 U24067 ( .A1(n21239), .A2(keyinput224), .B1(n21113), .B2(
        keyinput218), .ZN(n21112) );
  OAI221_X1 U24068 ( .B1(n21239), .B2(keyinput224), .C1(n21113), .C2(
        keyinput218), .A(n21112), .ZN(n21117) );
  AOI22_X1 U24069 ( .A1(n21115), .A2(keyinput160), .B1(keyinput241), .B2(
        n21302), .ZN(n21114) );
  OAI221_X1 U24070 ( .B1(n21115), .B2(keyinput160), .C1(n21302), .C2(
        keyinput241), .A(n21114), .ZN(n21116) );
  NOR4_X1 U24071 ( .A1(n21119), .A2(n21118), .A3(n21117), .A4(n21116), .ZN(
        n21134) );
  INV_X1 U24072 ( .A(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n21121) );
  AOI22_X1 U24073 ( .A1(n21305), .A2(keyinput216), .B1(n21121), .B2(
        keyinput162), .ZN(n21120) );
  OAI221_X1 U24074 ( .B1(n21305), .B2(keyinput216), .C1(n21121), .C2(
        keyinput162), .A(n21120), .ZN(n21125) );
  XOR2_X1 U24075 ( .A(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B(keyinput170), .Z(
        n21124) );
  XNOR2_X1 U24076 ( .A(n21122), .B(keyinput145), .ZN(n21123) );
  OR3_X1 U24077 ( .A1(n21125), .A2(n21124), .A3(n21123), .ZN(n21132) );
  AOI22_X1 U24078 ( .A1(n13669), .A2(keyinput177), .B1(keyinput144), .B2(
        n21127), .ZN(n21126) );
  OAI221_X1 U24079 ( .B1(n13669), .B2(keyinput177), .C1(n21127), .C2(
        keyinput144), .A(n21126), .ZN(n21131) );
  AOI22_X1 U24080 ( .A1(n21309), .A2(keyinput243), .B1(keyinput231), .B2(
        n21129), .ZN(n21128) );
  OAI221_X1 U24081 ( .B1(n21309), .B2(keyinput243), .C1(n21129), .C2(
        keyinput231), .A(n21128), .ZN(n21130) );
  NOR3_X1 U24082 ( .A1(n21132), .A2(n21131), .A3(n21130), .ZN(n21133) );
  NAND4_X1 U24083 ( .A1(n21136), .A2(n21135), .A3(n21134), .A4(n21133), .ZN(
        n21185) );
  AOI22_X1 U24084 ( .A1(n21221), .A2(keyinput191), .B1(n21192), .B2(
        keyinput200), .ZN(n21137) );
  OAI221_X1 U24085 ( .B1(n21221), .B2(keyinput191), .C1(n21192), .C2(
        keyinput200), .A(n21137), .ZN(n21146) );
  INV_X1 U24086 ( .A(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n21262) );
  AOI22_X1 U24087 ( .A1(n21262), .A2(keyinput236), .B1(keyinput182), .B2(
        n21236), .ZN(n21138) );
  OAI221_X1 U24088 ( .B1(n21262), .B2(keyinput236), .C1(n21236), .C2(
        keyinput182), .A(n21138), .ZN(n21145) );
  AOI22_X1 U24089 ( .A1(n21140), .A2(keyinput171), .B1(n21308), .B2(
        keyinput219), .ZN(n21139) );
  OAI221_X1 U24090 ( .B1(n21140), .B2(keyinput171), .C1(n21308), .C2(
        keyinput219), .A(n21139), .ZN(n21144) );
  INV_X1 U24091 ( .A(P1_UWORD_REG_0__SCAN_IN), .ZN(n21244) );
  AOI22_X1 U24092 ( .A1(n21244), .A2(keyinput201), .B1(n21142), .B2(
        keyinput220), .ZN(n21141) );
  OAI221_X1 U24093 ( .B1(n21244), .B2(keyinput201), .C1(n21142), .C2(
        keyinput220), .A(n21141), .ZN(n21143) );
  NOR4_X1 U24094 ( .A1(n21146), .A2(n21145), .A3(n21144), .A4(n21143), .ZN(
        n21183) );
  AOI22_X1 U24095 ( .A1(n21257), .A2(keyinput138), .B1(keyinput129), .B2(
        n21148), .ZN(n21147) );
  OAI221_X1 U24096 ( .B1(n21257), .B2(keyinput138), .C1(n21148), .C2(
        keyinput129), .A(n21147), .ZN(n21158) );
  AOI22_X1 U24097 ( .A1(n21150), .A2(keyinput156), .B1(n21275), .B2(
        keyinput246), .ZN(n21149) );
  OAI221_X1 U24098 ( .B1(n21150), .B2(keyinput156), .C1(n21275), .C2(
        keyinput246), .A(n21149), .ZN(n21157) );
  AOI22_X1 U24099 ( .A1(n21152), .A2(keyinput204), .B1(n13362), .B2(
        keyinput161), .ZN(n21151) );
  OAI221_X1 U24100 ( .B1(n21152), .B2(keyinput204), .C1(n13362), .C2(
        keyinput161), .A(n21151), .ZN(n21156) );
  XNOR2_X1 U24101 ( .A(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B(keyinput193), .ZN(
        n21154) );
  XNOR2_X1 U24102 ( .A(P1_EBX_REG_21__SCAN_IN), .B(keyinput242), .ZN(n21153)
         );
  NAND2_X1 U24103 ( .A1(n21154), .A2(n21153), .ZN(n21155) );
  NOR4_X1 U24104 ( .A1(n21158), .A2(n21157), .A3(n21156), .A4(n21155), .ZN(
        n21182) );
  AOI22_X1 U24105 ( .A1(n21336), .A2(keyinput207), .B1(keyinput169), .B2(
        n21160), .ZN(n21159) );
  OAI221_X1 U24106 ( .B1(n21336), .B2(keyinput207), .C1(n21160), .C2(
        keyinput169), .A(n21159), .ZN(n21169) );
  INV_X1 U24107 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n21243) );
  AOI22_X1 U24108 ( .A1(n21162), .A2(keyinput223), .B1(keyinput222), .B2(
        n21243), .ZN(n21161) );
  OAI221_X1 U24109 ( .B1(n21162), .B2(keyinput223), .C1(n21243), .C2(
        keyinput222), .A(n21161), .ZN(n21168) );
  INV_X1 U24110 ( .A(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n21189) );
  AOI22_X1 U24111 ( .A1(n21189), .A2(keyinput183), .B1(n10505), .B2(
        keyinput132), .ZN(n21163) );
  OAI221_X1 U24112 ( .B1(n21189), .B2(keyinput183), .C1(n10505), .C2(
        keyinput132), .A(n21163), .ZN(n21167) );
  XNOR2_X1 U24113 ( .A(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B(keyinput147), .ZN(
        n21165) );
  XNOR2_X1 U24114 ( .A(DATAI_5_), .B(keyinput254), .ZN(n21164) );
  NAND2_X1 U24115 ( .A1(n21165), .A2(n21164), .ZN(n21166) );
  NOR4_X1 U24116 ( .A1(n21169), .A2(n21168), .A3(n21167), .A4(n21166), .ZN(
        n21181) );
  AOI22_X1 U24117 ( .A1(n21240), .A2(keyinput214), .B1(n13935), .B2(
        keyinput190), .ZN(n21170) );
  OAI221_X1 U24118 ( .B1(n21240), .B2(keyinput214), .C1(n13935), .C2(
        keyinput190), .A(n21170), .ZN(n21179) );
  AOI22_X1 U24119 ( .A1(n21269), .A2(keyinput192), .B1(n21172), .B2(
        keyinput206), .ZN(n21171) );
  OAI221_X1 U24120 ( .B1(n21269), .B2(keyinput192), .C1(n21172), .C2(
        keyinput206), .A(n21171), .ZN(n21178) );
  INV_X1 U24121 ( .A(P1_LWORD_REG_6__SCAN_IN), .ZN(n21256) );
  AOI22_X1 U24122 ( .A1(n21256), .A2(keyinput165), .B1(n21174), .B2(
        keyinput154), .ZN(n21173) );
  OAI221_X1 U24123 ( .B1(n21256), .B2(keyinput165), .C1(n21174), .C2(
        keyinput154), .A(n21173), .ZN(n21177) );
  INV_X1 U24124 ( .A(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n21199) );
  AOI22_X1 U24125 ( .A1(n21199), .A2(keyinput205), .B1(keyinput180), .B2(
        n21242), .ZN(n21175) );
  OAI221_X1 U24126 ( .B1(n21199), .B2(keyinput205), .C1(n21242), .C2(
        keyinput180), .A(n21175), .ZN(n21176) );
  NOR4_X1 U24127 ( .A1(n21179), .A2(n21178), .A3(n21177), .A4(n21176), .ZN(
        n21180) );
  NAND4_X1 U24128 ( .A1(n21183), .A2(n21182), .A3(n21181), .A4(n21180), .ZN(
        n21184) );
  NOR4_X1 U24129 ( .A1(n21187), .A2(n21186), .A3(n21185), .A4(n21184), .ZN(
        n21396) );
  INV_X1 U24130 ( .A(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n21190) );
  AOI22_X1 U24131 ( .A1(n21190), .A2(keyinput5), .B1(keyinput55), .B2(n21189), 
        .ZN(n21188) );
  OAI221_X1 U24132 ( .B1(n21190), .B2(keyinput5), .C1(n21189), .C2(keyinput55), 
        .A(n21188), .ZN(n21203) );
  INV_X1 U24133 ( .A(P1_LWORD_REG_0__SCAN_IN), .ZN(n21193) );
  AOI22_X1 U24134 ( .A1(n21193), .A2(keyinput123), .B1(n21192), .B2(keyinput72), .ZN(n21191) );
  OAI221_X1 U24135 ( .B1(n21193), .B2(keyinput123), .C1(n21192), .C2(
        keyinput72), .A(n21191), .ZN(n21202) );
  AOI22_X1 U24136 ( .A1(n21196), .A2(keyinput36), .B1(n21195), .B2(keyinput12), 
        .ZN(n21194) );
  OAI221_X1 U24137 ( .B1(n21196), .B2(keyinput36), .C1(n21195), .C2(keyinput12), .A(n21194), .ZN(n21201) );
  AOI22_X1 U24138 ( .A1(n21199), .A2(keyinput77), .B1(keyinput8), .B2(n21198), 
        .ZN(n21197) );
  OAI221_X1 U24139 ( .B1(n21199), .B2(keyinput77), .C1(n21198), .C2(keyinput8), 
        .A(n21197), .ZN(n21200) );
  NOR4_X1 U24140 ( .A1(n21203), .A2(n21202), .A3(n21201), .A4(n21200), .ZN(
        n21254) );
  INV_X1 U24141 ( .A(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n21206) );
  INV_X1 U24142 ( .A(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n21205) );
  AOI22_X1 U24143 ( .A1(n21206), .A2(keyinput15), .B1(n21205), .B2(keyinput46), 
        .ZN(n21204) );
  OAI221_X1 U24144 ( .B1(n21206), .B2(keyinput15), .C1(n21205), .C2(keyinput46), .A(n21204), .ZN(n21218) );
  AOI22_X1 U24145 ( .A1(n10789), .A2(keyinput87), .B1(keyinput27), .B2(n21208), 
        .ZN(n21207) );
  OAI221_X1 U24146 ( .B1(n10789), .B2(keyinput87), .C1(n21208), .C2(keyinput27), .A(n21207), .ZN(n21217) );
  INV_X1 U24147 ( .A(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n21211) );
  AOI22_X1 U24148 ( .A1(n21211), .A2(keyinput25), .B1(keyinput35), .B2(n21210), 
        .ZN(n21209) );
  OAI221_X1 U24149 ( .B1(n21211), .B2(keyinput25), .C1(n21210), .C2(keyinput35), .A(n21209), .ZN(n21216) );
  INV_X1 U24150 ( .A(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n21214) );
  AOI22_X1 U24151 ( .A1(n21214), .A2(keyinput102), .B1(n21213), .B2(keyinput56), .ZN(n21212) );
  OAI221_X1 U24152 ( .B1(n21214), .B2(keyinput102), .C1(n21213), .C2(
        keyinput56), .A(n21212), .ZN(n21215) );
  NOR4_X1 U24153 ( .A1(n21218), .A2(n21217), .A3(n21216), .A4(n21215), .ZN(
        n21253) );
  AOI22_X1 U24154 ( .A1(n21221), .A2(keyinput63), .B1(n21220), .B2(keyinput0), 
        .ZN(n21219) );
  OAI221_X1 U24155 ( .B1(n21221), .B2(keyinput63), .C1(n21220), .C2(keyinput0), 
        .A(n21219), .ZN(n21225) );
  XNOR2_X1 U24156 ( .A(n21222), .B(keyinput48), .ZN(n21224) );
  XOR2_X1 U24157 ( .A(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B(keyinput24), .Z(
        n21223) );
  OR3_X1 U24158 ( .A1(n21225), .A2(n21224), .A3(n21223), .ZN(n21234) );
  AOI22_X1 U24159 ( .A1(n21228), .A2(keyinput98), .B1(keyinput119), .B2(n21227), .ZN(n21226) );
  OAI221_X1 U24160 ( .B1(n21228), .B2(keyinput98), .C1(n21227), .C2(
        keyinput119), .A(n21226), .ZN(n21233) );
  AOI22_X1 U24161 ( .A1(n21231), .A2(keyinput75), .B1(n21230), .B2(keyinput89), 
        .ZN(n21229) );
  OAI221_X1 U24162 ( .B1(n21231), .B2(keyinput75), .C1(n21230), .C2(keyinput89), .A(n21229), .ZN(n21232) );
  NOR3_X1 U24163 ( .A1(n21234), .A2(n21233), .A3(n21232), .ZN(n21252) );
  AOI22_X1 U24164 ( .A1(n21237), .A2(keyinput85), .B1(keyinput54), .B2(n21236), 
        .ZN(n21235) );
  OAI221_X1 U24165 ( .B1(n21237), .B2(keyinput85), .C1(n21236), .C2(keyinput54), .A(n21235), .ZN(n21250) );
  AOI22_X1 U24166 ( .A1(n21240), .A2(keyinput86), .B1(n21239), .B2(keyinput96), 
        .ZN(n21238) );
  OAI221_X1 U24167 ( .B1(n21240), .B2(keyinput86), .C1(n21239), .C2(keyinput96), .A(n21238), .ZN(n21249) );
  AOI22_X1 U24168 ( .A1(n21243), .A2(keyinput94), .B1(keyinput52), .B2(n21242), 
        .ZN(n21241) );
  OAI221_X1 U24169 ( .B1(n21243), .B2(keyinput94), .C1(n21242), .C2(keyinput52), .A(n21241), .ZN(n21248) );
  XOR2_X1 U24170 ( .A(n21244), .B(keyinput73), .Z(n21246) );
  XNOR2_X1 U24171 ( .A(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B(keyinput65), .ZN(
        n21245) );
  NAND2_X1 U24172 ( .A1(n21246), .A2(n21245), .ZN(n21247) );
  NOR4_X1 U24173 ( .A1(n21250), .A2(n21249), .A3(n21248), .A4(n21247), .ZN(
        n21251) );
  NAND4_X1 U24174 ( .A1(n21254), .A2(n21253), .A3(n21252), .A4(n21251), .ZN(
        n21395) );
  AOI22_X1 U24175 ( .A1(n21257), .A2(keyinput10), .B1(keyinput37), .B2(n21256), 
        .ZN(n21255) );
  OAI221_X1 U24176 ( .B1(n21257), .B2(keyinput10), .C1(n21256), .C2(keyinput37), .A(n21255), .ZN(n21267) );
  AOI22_X1 U24177 ( .A1(n21260), .A2(keyinput80), .B1(n21259), .B2(keyinput58), 
        .ZN(n21258) );
  OAI221_X1 U24178 ( .B1(n21260), .B2(keyinput80), .C1(n21259), .C2(keyinput58), .A(n21258), .ZN(n21266) );
  AOI22_X1 U24179 ( .A1(n21262), .A2(keyinput108), .B1(n10868), .B2(
        keyinput111), .ZN(n21261) );
  OAI221_X1 U24180 ( .B1(n21262), .B2(keyinput108), .C1(n10868), .C2(
        keyinput111), .A(n21261), .ZN(n21265) );
  AOI22_X1 U24181 ( .A1(n14569), .A2(keyinput59), .B1(n14563), .B2(keyinput61), 
        .ZN(n21263) );
  OAI221_X1 U24182 ( .B1(n14569), .B2(keyinput59), .C1(n14563), .C2(keyinput61), .A(n21263), .ZN(n21264) );
  NOR4_X1 U24183 ( .A1(n21267), .A2(n21266), .A3(n21265), .A4(n21264), .ZN(
        n21393) );
  OAI22_X1 U24184 ( .A1(n21270), .A2(keyinput20), .B1(n21269), .B2(keyinput64), 
        .ZN(n21268) );
  AOI221_X1 U24185 ( .B1(n21270), .B2(keyinput20), .C1(keyinput64), .C2(n21269), .A(n21268), .ZN(n21282) );
  OAI22_X1 U24186 ( .A1(n13935), .A2(keyinput62), .B1(n21272), .B2(keyinput100), .ZN(n21271) );
  AOI221_X1 U24187 ( .B1(n13935), .B2(keyinput62), .C1(keyinput100), .C2(
        n21272), .A(n21271), .ZN(n21281) );
  OAI22_X1 U24188 ( .A1(n21275), .A2(keyinput118), .B1(n21274), .B2(keyinput11), .ZN(n21273) );
  AOI221_X1 U24189 ( .B1(n21275), .B2(keyinput118), .C1(keyinput11), .C2(
        n21274), .A(n21273), .ZN(n21280) );
  OAI22_X1 U24190 ( .A1(n21278), .A2(keyinput93), .B1(n21277), .B2(keyinput30), 
        .ZN(n21276) );
  AOI221_X1 U24191 ( .B1(n21278), .B2(keyinput93), .C1(keyinput30), .C2(n21277), .A(n21276), .ZN(n21279) );
  NAND4_X1 U24192 ( .A1(n21282), .A2(n21281), .A3(n21280), .A4(n21279), .ZN(
        n21316) );
  OAI22_X1 U24193 ( .A1(n21285), .A2(keyinput23), .B1(n21284), .B2(keyinput47), 
        .ZN(n21283) );
  AOI221_X1 U24194 ( .B1(n21285), .B2(keyinput23), .C1(keyinput47), .C2(n21284), .A(n21283), .ZN(n21297) );
  OAI22_X1 U24195 ( .A1(n10505), .A2(keyinput4), .B1(n21287), .B2(keyinput99), 
        .ZN(n21286) );
  AOI221_X1 U24196 ( .B1(n10505), .B2(keyinput4), .C1(keyinput99), .C2(n21287), 
        .A(n21286), .ZN(n21296) );
  OAI22_X1 U24197 ( .A1(n21290), .A2(keyinput67), .B1(n21289), .B2(keyinput120), .ZN(n21288) );
  AOI221_X1 U24198 ( .B1(n21290), .B2(keyinput67), .C1(keyinput120), .C2(
        n21289), .A(n21288), .ZN(n21295) );
  OAI22_X1 U24199 ( .A1(n21293), .A2(keyinput101), .B1(n21292), .B2(
        keyinput117), .ZN(n21291) );
  AOI221_X1 U24200 ( .B1(n21293), .B2(keyinput101), .C1(keyinput117), .C2(
        n21292), .A(n21291), .ZN(n21294) );
  NAND4_X1 U24201 ( .A1(n21297), .A2(n21296), .A3(n21295), .A4(n21294), .ZN(
        n21315) );
  AOI22_X1 U24202 ( .A1(n21300), .A2(keyinput44), .B1(n21299), .B2(keyinput81), 
        .ZN(n21298) );
  OAI221_X1 U24203 ( .B1(n21300), .B2(keyinput44), .C1(n21299), .C2(keyinput81), .A(n21298), .ZN(n21314) );
  OAI22_X1 U24204 ( .A1(n21303), .A2(keyinput21), .B1(n21302), .B2(keyinput113), .ZN(n21301) );
  AOI221_X1 U24205 ( .B1(n21303), .B2(keyinput21), .C1(keyinput113), .C2(
        n21302), .A(n21301), .ZN(n21312) );
  OAI22_X1 U24206 ( .A1(n21306), .A2(keyinput74), .B1(n21305), .B2(keyinput88), 
        .ZN(n21304) );
  AOI221_X1 U24207 ( .B1(n21306), .B2(keyinput74), .C1(keyinput88), .C2(n21305), .A(n21304), .ZN(n21311) );
  OAI22_X1 U24208 ( .A1(n21309), .A2(keyinput115), .B1(n21308), .B2(keyinput91), .ZN(n21307) );
  AOI221_X1 U24209 ( .B1(n21309), .B2(keyinput115), .C1(keyinput91), .C2(
        n21308), .A(n21307), .ZN(n21310) );
  NAND3_X1 U24210 ( .A1(n21312), .A2(n21311), .A3(n21310), .ZN(n21313) );
  NOR4_X1 U24211 ( .A1(n21316), .A2(n21315), .A3(n21314), .A4(n21313), .ZN(
        n21392) );
  OAI22_X1 U24212 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(keyinput2), .B1(
        keyinput127), .B2(P3_EBX_REG_3__SCAN_IN), .ZN(n21317) );
  AOI221_X1 U24213 ( .B1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B2(keyinput2), .C1(
        P3_EBX_REG_3__SCAN_IN), .C2(keyinput127), .A(n21317), .ZN(n21324) );
  OAI22_X1 U24214 ( .A1(DATAI_5_), .A2(keyinput126), .B1(keyinput3), .B2(
        P3_EBX_REG_30__SCAN_IN), .ZN(n21318) );
  AOI221_X1 U24215 ( .B1(DATAI_5_), .B2(keyinput126), .C1(
        P3_EBX_REG_30__SCAN_IN), .C2(keyinput3), .A(n21318), .ZN(n21323) );
  OAI22_X1 U24216 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(keyinput49), .B1(
        P3_INSTQUEUE_REG_0__1__SCAN_IN), .B2(keyinput122), .ZN(n21319) );
  AOI221_X1 U24217 ( .B1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B2(keyinput49), 
        .C1(keyinput122), .C2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A(n21319), 
        .ZN(n21322) );
  OAI22_X1 U24218 ( .A1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A2(keyinput112), 
        .B1(keyinput34), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n21320) );
  AOI221_X1 U24219 ( .B1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B2(keyinput112), 
        .C1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .C2(keyinput34), .A(n21320), .ZN(
        n21321) );
  NAND4_X1 U24220 ( .A1(n21324), .A2(n21323), .A3(n21322), .A4(n21321), .ZN(
        n21353) );
  OAI22_X1 U24221 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(keyinput40), 
        .B1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B2(keyinput42), .ZN(n21325) );
  AOI221_X1 U24222 ( .B1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(keyinput40), 
        .C1(keyinput42), .C2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A(n21325), .ZN(
        n21332) );
  OAI22_X1 U24223 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(keyinput22), 
        .B1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B2(keyinput76), .ZN(n21326) );
  AOI221_X1 U24224 ( .B1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B2(keyinput22), 
        .C1(keyinput76), .C2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A(n21326), .ZN(
        n21331) );
  OAI22_X1 U24225 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(keyinput18), 
        .B1(P2_DATAWIDTH_REG_1__SCAN_IN), .B2(keyinput83), .ZN(n21327) );
  AOI221_X1 U24226 ( .B1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B2(keyinput18), 
        .C1(keyinput83), .C2(P2_DATAWIDTH_REG_1__SCAN_IN), .A(n21327), .ZN(
        n21330) );
  OAI22_X1 U24227 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(keyinput33), .B1(
        P2_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(keyinput29), .ZN(n21328) );
  AOI221_X1 U24228 ( .B1(P2_STATE2_REG_1__SCAN_IN), .B2(keyinput33), .C1(
        keyinput29), .C2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A(n21328), .ZN(
        n21329) );
  NAND4_X1 U24229 ( .A1(n21332), .A2(n21331), .A3(n21330), .A4(n21329), .ZN(
        n21352) );
  OAI22_X1 U24230 ( .A1(P1_INSTQUEUE_REG_5__5__SCAN_IN), .A2(keyinput92), .B1(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(keyinput9), .ZN(n21333) );
  AOI221_X1 U24231 ( .B1(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B2(keyinput92), 
        .C1(keyinput9), .C2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A(n21333), 
        .ZN(n21341) );
  OAI22_X1 U24232 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(keyinput66), .B1(
        keyinput51), .B2(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n21334) );
  AOI221_X1 U24233 ( .B1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B2(keyinput66), 
        .C1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .C2(keyinput51), .A(n21334), 
        .ZN(n21340) );
  OAI22_X1 U24234 ( .A1(n21336), .A2(keyinput79), .B1(keyinput70), .B2(
        P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n21335) );
  AOI221_X1 U24235 ( .B1(n21336), .B2(keyinput79), .C1(
        P2_INSTQUEUE_REG_8__2__SCAN_IN), .C2(keyinput70), .A(n21335), .ZN(
        n21339) );
  OAI22_X1 U24236 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(keyinput19), .B1(
        keyinput124), .B2(P3_EAX_REG_1__SCAN_IN), .ZN(n21337) );
  AOI221_X1 U24237 ( .B1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B2(keyinput19), 
        .C1(P3_EAX_REG_1__SCAN_IN), .C2(keyinput124), .A(n21337), .ZN(n21338)
         );
  NAND4_X1 U24238 ( .A1(n21341), .A2(n21340), .A3(n21339), .A4(n21338), .ZN(
        n21351) );
  OAI22_X1 U24239 ( .A1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .A2(keyinput57), .B1(
        keyinput1), .B2(P3_EBX_REG_19__SCAN_IN), .ZN(n21342) );
  AOI221_X1 U24240 ( .B1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B2(keyinput57), 
        .C1(P3_EBX_REG_19__SCAN_IN), .C2(keyinput1), .A(n21342), .ZN(n21349)
         );
  OAI22_X1 U24241 ( .A1(P2_EAX_REG_29__SCAN_IN), .A2(keyinput116), .B1(
        keyinput17), .B2(P2_DATAO_REG_0__SCAN_IN), .ZN(n21343) );
  AOI221_X1 U24242 ( .B1(P2_EAX_REG_29__SCAN_IN), .B2(keyinput116), .C1(
        P2_DATAO_REG_0__SCAN_IN), .C2(keyinput17), .A(n21343), .ZN(n21348) );
  OAI22_X1 U24243 ( .A1(P1_EAX_REG_30__SCAN_IN), .A2(keyinput6), .B1(
        keyinput97), .B2(P1_DATAO_REG_12__SCAN_IN), .ZN(n21344) );
  AOI221_X1 U24244 ( .B1(P1_EAX_REG_30__SCAN_IN), .B2(keyinput6), .C1(
        P1_DATAO_REG_12__SCAN_IN), .C2(keyinput97), .A(n21344), .ZN(n21347) );
  OAI22_X1 U24245 ( .A1(P1_INSTQUEUE_REG_6__7__SCAN_IN), .A2(keyinput45), .B1(
        keyinput50), .B2(DATAI_2_), .ZN(n21345) );
  AOI221_X1 U24246 ( .B1(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B2(keyinput45), 
        .C1(DATAI_2_), .C2(keyinput50), .A(n21345), .ZN(n21346) );
  NAND4_X1 U24247 ( .A1(n21349), .A2(n21348), .A3(n21347), .A4(n21346), .ZN(
        n21350) );
  NOR4_X1 U24248 ( .A1(n21353), .A2(n21352), .A3(n21351), .A4(n21350), .ZN(
        n21391) );
  OAI22_X1 U24249 ( .A1(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(keyinput106), 
        .B1(P3_ADDRESS_REG_22__SCAN_IN), .B2(keyinput68), .ZN(n21354) );
  AOI221_X1 U24250 ( .B1(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(keyinput106), 
        .C1(keyinput68), .C2(P3_ADDRESS_REG_22__SCAN_IN), .A(n21354), .ZN(
        n21361) );
  OAI22_X1 U24251 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(keyinput90), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(keyinput95), .ZN(n21355) );
  AOI221_X1 U24252 ( .B1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B2(keyinput90), 
        .C1(keyinput95), .C2(P2_DATAO_REG_16__SCAN_IN), .A(n21355), .ZN(n21360) );
  OAI22_X1 U24253 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(keyinput13), .B1(
        keyinput110), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n21356) );
  AOI221_X1 U24254 ( .B1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B2(keyinput13), 
        .C1(P1_INSTQUEUE_REG_7__1__SCAN_IN), .C2(keyinput110), .A(n21356), 
        .ZN(n21359) );
  OAI22_X1 U24255 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(keyinput71), .B1(
        keyinput16), .B2(P3_EAX_REG_4__SCAN_IN), .ZN(n21357) );
  AOI221_X1 U24256 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(keyinput71), .C1(
        P3_EAX_REG_4__SCAN_IN), .C2(keyinput16), .A(n21357), .ZN(n21358) );
  NAND4_X1 U24257 ( .A1(n21361), .A2(n21360), .A3(n21359), .A4(n21358), .ZN(
        n21389) );
  OAI22_X1 U24258 ( .A1(BUF1_REG_18__SCAN_IN), .A2(keyinput39), .B1(
        P3_ADDRESS_REG_13__SCAN_IN), .B2(keyinput103), .ZN(n21362) );
  AOI221_X1 U24259 ( .B1(BUF1_REG_18__SCAN_IN), .B2(keyinput39), .C1(
        keyinput103), .C2(P3_ADDRESS_REG_13__SCAN_IN), .A(n21362), .ZN(n21369)
         );
  OAI22_X1 U24260 ( .A1(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(keyinput32), 
        .B1(keyinput31), .B2(DATAI_12_), .ZN(n21363) );
  AOI221_X1 U24261 ( .B1(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(keyinput32), 
        .C1(DATAI_12_), .C2(keyinput31), .A(n21363), .ZN(n21368) );
  OAI22_X1 U24262 ( .A1(P3_ADDRESS_REG_26__SCAN_IN), .A2(keyinput82), .B1(
        P3_DATAWIDTH_REG_20__SCAN_IN), .B2(keyinput28), .ZN(n21364) );
  AOI221_X1 U24263 ( .B1(P3_ADDRESS_REG_26__SCAN_IN), .B2(keyinput82), .C1(
        keyinput28), .C2(P3_DATAWIDTH_REG_20__SCAN_IN), .A(n21364), .ZN(n21367) );
  OAI22_X1 U24264 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(keyinput43), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(keyinput41), .ZN(n21365) );
  AOI221_X1 U24265 ( .B1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B2(keyinput43), 
        .C1(keyinput41), .C2(P3_UWORD_REG_12__SCAN_IN), .A(n21365), .ZN(n21366) );
  NAND4_X1 U24266 ( .A1(n21369), .A2(n21368), .A3(n21367), .A4(n21366), .ZN(
        n21388) );
  OAI22_X1 U24267 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(keyinput60), .B1(
        keyinput121), .B2(P3_DATAWIDTH_REG_6__SCAN_IN), .ZN(n21370) );
  AOI221_X1 U24268 ( .B1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B2(keyinput60), 
        .C1(P3_DATAWIDTH_REG_6__SCAN_IN), .C2(keyinput121), .A(n21370), .ZN(
        n21377) );
  OAI22_X1 U24269 ( .A1(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(keyinput109), 
        .B1(DATAI_0_), .B2(keyinput107), .ZN(n21371) );
  AOI221_X1 U24270 ( .B1(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(keyinput109), 
        .C1(keyinput107), .C2(DATAI_0_), .A(n21371), .ZN(n21376) );
  OAI22_X1 U24271 ( .A1(P1_ADDRESS_REG_3__SCAN_IN), .A2(keyinput78), .B1(
        keyinput26), .B2(DATAI_11_), .ZN(n21372) );
  AOI221_X1 U24272 ( .B1(P1_ADDRESS_REG_3__SCAN_IN), .B2(keyinput78), .C1(
        DATAI_11_), .C2(keyinput26), .A(n21372), .ZN(n21375) );
  OAI22_X1 U24273 ( .A1(P1_EBX_REG_21__SCAN_IN), .A2(keyinput114), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(keyinput105), .ZN(n21373) );
  AOI221_X1 U24274 ( .B1(P1_EBX_REG_21__SCAN_IN), .B2(keyinput114), .C1(
        keyinput105), .C2(P3_UWORD_REG_4__SCAN_IN), .A(n21373), .ZN(n21374) );
  NAND4_X1 U24275 ( .A1(n21377), .A2(n21376), .A3(n21375), .A4(n21374), .ZN(
        n21387) );
  OAI22_X1 U24276 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(keyinput125), .B1(
        P3_DATAWIDTH_REG_1__SCAN_IN), .B2(keyinput38), .ZN(n21378) );
  AOI221_X1 U24277 ( .B1(P3_EAX_REG_7__SCAN_IN), .B2(keyinput125), .C1(
        keyinput38), .C2(P3_DATAWIDTH_REG_1__SCAN_IN), .A(n21378), .ZN(n21385)
         );
  OAI22_X1 U24278 ( .A1(DATAI_22_), .A2(keyinput7), .B1(
        P2_UWORD_REG_0__SCAN_IN), .B2(keyinput53), .ZN(n21379) );
  AOI221_X1 U24279 ( .B1(DATAI_22_), .B2(keyinput7), .C1(keyinput53), .C2(
        P2_UWORD_REG_0__SCAN_IN), .A(n21379), .ZN(n21384) );
  OAI22_X1 U24280 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(keyinput14), .B1(
        P2_ADDRESS_REG_10__SCAN_IN), .B2(keyinput84), .ZN(n21380) );
  AOI221_X1 U24281 ( .B1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B2(keyinput14), 
        .C1(keyinput84), .C2(P2_ADDRESS_REG_10__SCAN_IN), .A(n21380), .ZN(
        n21383) );
  OAI22_X1 U24282 ( .A1(P2_EAX_REG_10__SCAN_IN), .A2(keyinput69), .B1(
        keyinput104), .B2(P1_REIP_REG_29__SCAN_IN), .ZN(n21381) );
  AOI221_X1 U24283 ( .B1(P2_EAX_REG_10__SCAN_IN), .B2(keyinput69), .C1(
        P1_REIP_REG_29__SCAN_IN), .C2(keyinput104), .A(n21381), .ZN(n21382) );
  NAND4_X1 U24284 ( .A1(n21385), .A2(n21384), .A3(n21383), .A4(n21382), .ZN(
        n21386) );
  NOR4_X1 U24285 ( .A1(n21389), .A2(n21388), .A3(n21387), .A4(n21386), .ZN(
        n21390) );
  NAND4_X1 U24286 ( .A1(n21393), .A2(n21392), .A3(n21391), .A4(n21390), .ZN(
        n21394) );
  NOR3_X1 U24287 ( .A1(n21396), .A2(n21395), .A3(n21394), .ZN(n21401) );
  NAND2_X1 U24288 ( .A1(n21397), .A2(n21399), .ZN(n21398) );
  OAI21_X1 U24289 ( .B1(n21399), .B2(P1_MORE_REG_SCAN_IN), .A(n21398), .ZN(
        n21400) );
  XNOR2_X1 U24290 ( .A(n21401), .B(n21400), .ZN(P1_U3484) );
  NOR2_X2 U11266 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10308) );
  CLKBUF_X1 U11297 ( .A(n11716), .Z(n12185) );
  CLKBUF_X1 U11304 ( .A(n12929), .Z(n9856) );
  CLKBUF_X1 U11388 ( .A(n11149), .Z(n11167) );
  CLKBUF_X1 U11416 ( .A(n11457), .Z(n11459) );
  CLKBUF_X1 U11902 ( .A(n12857), .Z(n16195) );
  CLKBUF_X3 U12516 ( .A(n11907), .Z(n9845) );
  CLKBUF_X1 U12765 ( .A(n11657), .Z(n13521) );
  CLKBUF_X1 U14685 ( .A(n16000), .Z(n16020) );
endmodule

