

module b20_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, P2_WR_REG_SCAN_IN, SI_31_, 
        SI_30_, SI_29_, SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, 
        SI_21_, SI_20_, SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, 
        SI_12_, SI_11_, SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, 
        SI_3_, SI_2_, SI_1_, SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, ADD_1068_U4, 
        ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58, ADD_1068_U59, 
        ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63, ADD_1068_U47, 
        ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51, ADD_1068_U52, 
        ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46, U126, U123, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439, P1_U3440, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462, P1_U3465, P1_U3468, 
        P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, 
        P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3509, 
        P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, 
        P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, 
        P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, 
        P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, 
        P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, 
        P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, 
        P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3554, P1_U3555, 
        P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, 
        P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, 
        P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, 
        P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, 
        P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U3973, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376, P2_U3377, P2_U3263, 
        P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, 
        P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, 
        P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, 
        P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, 
        P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399, P2_U3402, P2_U3405, 
        P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420, P2_U3423, P2_U3426, 
        P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441, P2_U3444, P2_U3446, 
        P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451, P2_U3452, P2_U3453, 
        P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458, P2_U3459, P2_U3460, 
        P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465, P2_U3466, P2_U3467, 
        P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472, P2_U3473, P2_U3474, 
        P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479, P2_U3480, P2_U3481, 
        P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486, P2_U3487, P2_U3488, 
        P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, 
        P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, 
        P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, 
        P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3491, P2_U3492, 
        P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, 
        P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, 
        P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, 
        P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, 
        P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180, P2_U3179, P2_U3178, 
        P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, P2_U3171, 
        P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, P2_U3164, 
        P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, P2_U3157, 
        P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151, P2_U3150, P2_U3893
 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_,
         SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_,
         SI_20_, SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_,
         SI_12_, SI_11_, SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_,
         SI_3_, SI_2_, SI_1_, SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_REG3_REG_7__SCAN_IN, P2_REG3_REG_27__SCAN_IN,
         P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_23__SCAN_IN,
         P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_3__SCAN_IN,
         P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_28__SCAN_IN,
         P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_1__SCAN_IN,
         P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_12__SCAN_IN,
         P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_16__SCAN_IN,
         P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_17__SCAN_IN,
         P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_4__SCAN_IN,
         P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN,
         P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN,
         P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN,
         P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN,
         P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN,
         P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950,
         n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960,
         n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970,
         n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980,
         n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990,
         n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000,
         n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010,
         n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020,
         n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030,
         n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040,
         n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050,
         n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060,
         n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070,
         n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080,
         n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090,
         n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100,
         n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110,
         n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120,
         n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130,
         n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140,
         n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150,
         n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160,
         n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170,
         n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180,
         n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190,
         n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200,
         n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210,
         n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220,
         n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230,
         n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240,
         n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250,
         n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260,
         n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270,
         n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280,
         n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290,
         n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300,
         n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310,
         n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320,
         n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330,
         n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340,
         n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350,
         n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360,
         n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370,
         n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380,
         n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390,
         n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400,
         n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410,
         n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420,
         n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430,
         n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440,
         n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450,
         n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460,
         n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470,
         n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480,
         n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490,
         n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500,
         n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510,
         n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520,
         n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530,
         n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540,
         n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550,
         n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560,
         n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570,
         n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580,
         n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590,
         n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600,
         n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610,
         n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620,
         n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630,
         n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640,
         n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650,
         n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660,
         n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670,
         n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680,
         n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690,
         n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700,
         n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710,
         n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720,
         n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730,
         n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740,
         n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750,
         n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760,
         n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770,
         n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780,
         n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790,
         n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800,
         n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810,
         n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820,
         n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830,
         n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840,
         n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850,
         n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860,
         n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870,
         n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880,
         n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890,
         n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900,
         n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910,
         n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920,
         n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930,
         n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940,
         n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950,
         n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960,
         n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970,
         n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980,
         n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990,
         n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000,
         n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010,
         n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020,
         n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030,
         n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040,
         n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050,
         n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060,
         n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070,
         n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080,
         n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090,
         n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100,
         n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110,
         n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120,
         n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130,
         n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140,
         n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150,
         n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160,
         n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170,
         n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180,
         n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190,
         n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200,
         n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210,
         n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220,
         n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230,
         n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240,
         n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250,
         n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260,
         n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270,
         n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280,
         n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290,
         n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300,
         n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310,
         n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320,
         n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330,
         n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340,
         n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350,
         n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360,
         n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370,
         n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380,
         n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390,
         n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400,
         n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410,
         n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420,
         n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430,
         n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440,
         n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450,
         n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460,
         n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470,
         n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480,
         n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490,
         n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500,
         n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510,
         n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520,
         n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530,
         n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540,
         n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550,
         n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560,
         n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570,
         n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580,
         n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590,
         n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600,
         n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610,
         n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620,
         n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630,
         n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640,
         n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650,
         n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660,
         n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670,
         n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680,
         n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690,
         n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700,
         n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710,
         n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720,
         n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730,
         n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740,
         n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750,
         n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760,
         n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770,
         n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780,
         n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790,
         n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800,
         n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810,
         n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820,
         n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830,
         n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840,
         n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850,
         n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860,
         n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870,
         n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880,
         n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890,
         n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900,
         n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910,
         n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920,
         n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930,
         n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940,
         n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950,
         n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960,
         n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970,
         n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980,
         n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990,
         n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000,
         n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010,
         n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020,
         n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030,
         n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040,
         n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050,
         n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060,
         n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070,
         n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080,
         n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090,
         n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100,
         n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110,
         n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120,
         n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130,
         n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140,
         n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150,
         n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160,
         n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170,
         n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180,
         n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190,
         n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200,
         n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210,
         n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220,
         n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230,
         n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240,
         n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250,
         n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260,
         n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270,
         n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280,
         n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290,
         n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300,
         n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310,
         n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320,
         n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330,
         n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340,
         n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350,
         n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360,
         n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370,
         n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380,
         n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390,
         n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400,
         n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410,
         n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420,
         n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430,
         n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440,
         n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450,
         n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460,
         n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470,
         n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480,
         n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490,
         n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500,
         n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510,
         n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520,
         n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530,
         n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540,
         n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550,
         n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560,
         n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570,
         n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580,
         n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590,
         n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600,
         n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610,
         n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620,
         n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630,
         n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640,
         n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650,
         n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660,
         n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670,
         n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680,
         n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690,
         n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700,
         n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710,
         n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720,
         n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730,
         n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740,
         n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750,
         n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760,
         n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770,
         n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780,
         n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790,
         n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800,
         n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810,
         n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820,
         n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830,
         n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840,
         n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850,
         n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860,
         n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870,
         n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880,
         n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890,
         n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900,
         n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910,
         n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920,
         n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930,
         n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940,
         n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950,
         n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960,
         n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970,
         n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980,
         n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990,
         n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000,
         n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010,
         n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020,
         n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030,
         n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040,
         n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050,
         n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060,
         n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070,
         n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080,
         n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090,
         n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101,
         n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111,
         n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121,
         n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131,
         n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141,
         n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151,
         n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161,
         n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171,
         n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181,
         n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191,
         n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201,
         n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211,
         n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221,
         n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231,
         n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241,
         n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251,
         n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261,
         n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271,
         n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281,
         n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291,
         n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301,
         n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311,
         n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321,
         n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331,
         n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341,
         n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351,
         n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361,
         n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371,
         n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381,
         n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391,
         n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401,
         n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411,
         n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421,
         n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431,
         n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441,
         n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451,
         n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461,
         n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471,
         n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481,
         n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491,
         n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501,
         n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511,
         n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521,
         n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531,
         n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541,
         n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551,
         n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561,
         n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571,
         n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581,
         n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591,
         n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601,
         n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611,
         n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621,
         n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631,
         n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641,
         n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651,
         n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661,
         n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671,
         n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681,
         n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691,
         n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701,
         n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711,
         n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721,
         n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731,
         n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741,
         n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751,
         n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761,
         n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771,
         n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781,
         n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791,
         n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801,
         n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811,
         n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821,
         n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831,
         n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841,
         n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851,
         n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861,
         n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871,
         n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881,
         n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891,
         n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901,
         n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911,
         n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921,
         n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931,
         n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941,
         n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951,
         n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961,
         n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971,
         n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981,
         n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991,
         n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001,
         n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011,
         n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021,
         n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031,
         n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041,
         n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051,
         n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061,
         n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071,
         n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081,
         n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091,
         n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101,
         n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111,
         n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121,
         n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131,
         n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141,
         n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151,
         n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161,
         n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171,
         n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181,
         n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191,
         n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201,
         n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211,
         n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221,
         n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231,
         n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241,
         n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251,
         n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261,
         n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271,
         n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281,
         n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291,
         n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301,
         n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311,
         n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321,
         n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331,
         n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341,
         n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351,
         n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361,
         n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371,
         n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381,
         n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391,
         n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401,
         n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411,
         n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421,
         n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431,
         n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441,
         n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451,
         n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461,
         n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471,
         n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481,
         n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491,
         n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501,
         n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511,
         n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521,
         n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531,
         n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541,
         n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551,
         n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561,
         n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571,
         n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581,
         n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591,
         n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601,
         n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611,
         n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621,
         n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631,
         n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641,
         n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651,
         n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661,
         n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671,
         n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681,
         n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691,
         n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701,
         n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711,
         n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721,
         n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731,
         n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741,
         n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751,
         n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761,
         n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771,
         n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781,
         n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791,
         n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801,
         n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811,
         n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821,
         n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831,
         n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841,
         n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851,
         n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861,
         n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871,
         n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881,
         n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891,
         n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901,
         n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911,
         n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921,
         n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931,
         n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941,
         n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951,
         n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961,
         n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971,
         n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981,
         n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991,
         n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
         n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
         n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
         n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
         n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
         n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
         n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280,
         n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288,
         n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296,
         n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304,
         n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
         n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320,
         n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328,
         n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336,
         n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344,
         n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352,
         n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360,
         n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368,
         n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376,
         n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384,
         n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392,
         n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400,
         n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408,
         n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416,
         n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424,
         n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432,
         n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440,
         n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448,
         n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456,
         n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464,
         n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472,
         n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480,
         n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488,
         n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496,
         n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504,
         n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512,
         n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520,
         n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528,
         n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536,
         n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544,
         n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552,
         n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560,
         n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568,
         n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576,
         n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584,
         n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592,
         n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600,
         n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608,
         n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616,
         n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624,
         n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632,
         n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640,
         n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648,
         n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656,
         n10657, n10658, n10659, n10660, n10661, n10662, n10663, n10664,
         n10665, n10666, n10667, n10668, n10669, n10670, n10671, n10672,
         n10673, n10674, n10675, n10676, n10677, n10678, n10679, n10680,
         n10681, n10682, n10683, n10684, n10685, n10686, n10687, n10688,
         n10689, n10690, n10691, n10692, n10693, n10694, n10695;

  NAND2_X1 U5005 ( .A1(n6749), .A2(n6748), .ZN(n9581) );
  INV_X2 U5006 ( .A(n7170), .ZN(n7140) );
  CLKBUF_X2 U5007 ( .A(n6983), .Z(n7168) );
  CLKBUF_X2 U5009 ( .A(n6526), .Z(n8851) );
  CLKBUF_X1 U5010 ( .A(n5655), .Z(n6018) );
  CLKBUF_X2 U5011 ( .A(n6667), .Z(n8848) );
  CLKBUF_X1 U5012 ( .A(n10619), .Z(n4941) );
  AND2_X1 U5013 ( .A1(n7830), .A2(n10606), .ZN(n10619) );
  INV_X1 U5014 ( .A(n10296), .ZN(n4942) );
  INV_X1 U5015 ( .A(n4942), .ZN(n4943) );
  NAND2_X1 U5016 ( .A1(n6963), .A2(n6981), .ZN(n6983) );
  NOR2_X1 U5017 ( .A1(n9581), .A2(n9585), .ZN(n9027) );
  NOR2_X1 U5018 ( .A1(n9062), .A2(n6924), .ZN(n6928) );
  NAND2_X1 U5019 ( .A1(n9596), .A2(n9007), .ZN(n9505) );
  INV_X1 U5020 ( .A(n7018), .ZN(n7170) );
  INV_X1 U5021 ( .A(n6981), .ZN(n7163) );
  INV_X1 U5022 ( .A(n6963), .ZN(n7166) );
  INV_X1 U5023 ( .A(n9060), .ZN(n9053) );
  NAND2_X1 U5024 ( .A1(n6860), .A2(n8964), .ZN(n8888) );
  BUF_X1 U5025 ( .A(n10650), .Z(n4944) );
  INV_X1 U5026 ( .A(n5436), .ZN(n7864) );
  OAI21_X2 U5027 ( .B1(n7962), .B2(n6856), .A(n8950), .ZN(n8062) );
  NAND2_X2 U5028 ( .A1(n6855), .A2(n8946), .ZN(n7962) );
  INV_X2 U5029 ( .A(n8246), .ZN(n5343) );
  NAND2_X2 U5030 ( .A1(n6483), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6480) );
  OAI21_X1 U5033 ( .B1(n7465), .B2(n6018), .A(n5765), .ZN(n10650) );
  NAND2_X1 U5034 ( .A1(n9667), .A2(n9664), .ZN(n6509) );
  NAND4_X4 U5035 ( .A1(n5611), .A2(n5610), .A3(n5609), .A4(n5608), .ZN(n6960)
         );
  XNOR2_X2 U5036 ( .A(n5662), .B(P1_IR_REG_2__SCAN_IN), .ZN(n9831) );
  AOI22_X1 U5037 ( .A1(n8847), .A2(n8849), .B1(n8848), .B2(
        P1_DATAO_REG_31__SCAN_IN), .ZN(n9630) );
  OAI21_X1 U5038 ( .B1(n8801), .B2(n5453), .A(n5825), .ZN(n5452) );
  INV_X1 U5039 ( .A(n9563), .ZN(n9245) );
  NOR2_X2 U5040 ( .A1(n8115), .A2(n6987), .ZN(n7951) );
  NAND2_X1 U5041 ( .A1(n8922), .A2(n8931), .ZN(n6851) );
  INV_X1 U5042 ( .A(n9288), .ZN(n7961) );
  NAND2_X1 U5043 ( .A1(n9291), .A2(n10586), .ZN(n8922) );
  INV_X1 U5044 ( .A(n9287), .ZN(n6575) );
  INV_X1 U5045 ( .A(n9290), .ZN(n7792) );
  CLKBUF_X3 U5046 ( .A(n5633), .Z(n6171) );
  INV_X1 U5047 ( .A(n7831), .ZN(n7857) );
  OR2_X1 U5048 ( .A1(n5602), .A2(n5601), .ZN(n5625) );
  INV_X1 U5049 ( .A(n7523), .ZN(n6508) );
  NOR2_X1 U5050 ( .A1(n7491), .A2(n7199), .ZN(P2_U3893) );
  NAND2_X2 U5051 ( .A1(n5618), .A2(n7435), .ZN(n5655) );
  INV_X2 U5052 ( .A(n7271), .ZN(n9074) );
  NAND2_X2 U5053 ( .A1(n6845), .A2(n6846), .ZN(n6515) );
  NAND2_X1 U5054 ( .A1(n6481), .A2(n6479), .ZN(n6483) );
  NAND2_X1 U5055 ( .A1(n5726), .A2(n5571), .ZN(n5733) );
  NOR2_X1 U5057 ( .A1(P2_IR_REG_4__SCAN_IN), .A2(P2_IR_REG_5__SCAN_IN), .ZN(
        n6471) );
  NOR2_X1 U5058 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n6472) );
  AOI21_X1 U5059 ( .B1(n10552), .B2(n9965), .A(n9971), .ZN(n6115) );
  OR2_X1 U5060 ( .A1(n5214), .A2(n9080), .ZN(n5208) );
  NAND2_X1 U5061 ( .A1(n5126), .A2(n10667), .ZN(n5125) );
  INV_X1 U5062 ( .A(n9973), .ZN(n5126) );
  OR2_X1 U5063 ( .A1(n8859), .A2(n9065), .ZN(n8860) );
  AND2_X1 U5064 ( .A1(n9748), .A2(n9747), .ZN(n9751) );
  NAND2_X1 U5065 ( .A1(n5239), .A2(n5238), .ZN(n9417) );
  OR2_X1 U5066 ( .A1(n8863), .A2(n8862), .ZN(n9064) );
  INV_X1 U5067 ( .A(n8863), .ZN(n9633) );
  AND2_X1 U5068 ( .A1(n5403), .A2(n6211), .ZN(n4948) );
  NAND2_X1 U5069 ( .A1(n8846), .A2(n8845), .ZN(n8863) );
  NAND2_X1 U5070 ( .A1(n5160), .A2(n5159), .ZN(n9452) );
  NAND2_X1 U5071 ( .A1(n5455), .A2(n5454), .ZN(n10025) );
  AND2_X1 U5072 ( .A1(n8839), .A2(n9273), .ZN(n9062) );
  XNOR2_X1 U5073 ( .A(n6216), .B(n6215), .ZN(n9663) );
  NAND2_X1 U5074 ( .A1(n7096), .A2(n5011), .ZN(n9770) );
  OAI21_X1 U5075 ( .B1(n9648), .B2(n9580), .A(n9461), .ZN(n5160) );
  NAND2_X1 U5076 ( .A1(n5276), .A2(n8874), .ZN(n5275) );
  NOR2_X1 U5077 ( .A1(n9499), .A2(n9504), .ZN(n9497) );
  NAND2_X1 U5078 ( .A1(n6501), .A2(n6500), .ZN(n9564) );
  NAND2_X1 U5079 ( .A1(n9541), .A2(n4957), .ZN(n9596) );
  NAND2_X1 U5080 ( .A1(n8786), .A2(n5516), .ZN(n5847) );
  OAI21_X1 U5081 ( .B1(n8808), .B2(n4960), .A(n5345), .ZN(n10123) );
  NAND2_X1 U5082 ( .A1(n5997), .A2(n5996), .ZN(n10181) );
  NAND2_X1 U5083 ( .A1(n5313), .A2(n5312), .ZN(n8775) );
  NAND2_X1 U5084 ( .A1(n9648), .A2(n9580), .ZN(n5159) );
  NAND2_X1 U5085 ( .A1(n6778), .A2(n6777), .ZN(n9215) );
  NAND2_X1 U5086 ( .A1(n6768), .A2(n6767), .ZN(n9572) );
  OR2_X1 U5087 ( .A1(n5347), .A2(n5351), .ZN(n4960) );
  NAND2_X1 U5088 ( .A1(n5932), .A2(n5931), .ZN(n10200) );
  NAND2_X1 U5089 ( .A1(n8311), .A2(n6862), .ZN(n8390) );
  NAND2_X1 U5090 ( .A1(n6740), .A2(n6739), .ZN(n9586) );
  NAND2_X1 U5091 ( .A1(n6787), .A2(n6786), .ZN(n9446) );
  NAND2_X1 U5092 ( .A1(n5839), .A2(n5838), .ZN(n10225) );
  AND2_X1 U5093 ( .A1(n6637), .A2(n6862), .ZN(n8890) );
  NAND2_X1 U5094 ( .A1(n5811), .A2(n5810), .ZN(n10235) );
  NAND2_X1 U5095 ( .A1(n5172), .A2(n5174), .ZN(n5831) );
  NAND2_X1 U5096 ( .A1(n6612), .A2(n6611), .ZN(n8359) );
  OR2_X1 U5097 ( .A1(n7002), .A2(n5056), .ZN(n5054) );
  INV_X1 U5098 ( .A(n8080), .ZN(n4945) );
  INV_X1 U5099 ( .A(n5757), .ZN(n4946) );
  NAND2_X1 U5100 ( .A1(n6603), .A2(n6602), .ZN(n8241) );
  NAND2_X1 U5101 ( .A1(n5219), .A2(n6594), .ZN(n10637) );
  NAND2_X1 U5102 ( .A1(n5109), .A2(n5115), .ZN(n5761) );
  NAND2_X1 U5103 ( .A1(n5746), .A2(n5745), .ZN(n5109) );
  NAND2_X1 U5104 ( .A1(n7497), .A2(n7496), .ZN(n9266) );
  NAND2_X1 U5105 ( .A1(n5205), .A2(n5554), .ZN(n5746) );
  NAND2_X2 U5106 ( .A1(n7838), .A2(n10593), .ZN(n6390) );
  NAND2_X1 U5107 ( .A1(n5723), .A2(n5722), .ZN(n5725) );
  XNOR2_X1 U5108 ( .A(n6965), .B(n6960), .ZN(n5436) );
  INV_X2 U5109 ( .A(n9110), .ZN(n9115) );
  AND4_X1 U5110 ( .A1(n5708), .A2(n5707), .A3(n5706), .A4(n5705), .ZN(n8136)
         );
  NAND3_X1 U5111 ( .A1(n5629), .A2(n5628), .A3(n5627), .ZN(n7932) );
  NAND4_X2 U5112 ( .A1(n5638), .A2(n5637), .A3(n5636), .A4(n5635), .ZN(n6970)
         );
  INV_X1 U5113 ( .A(n5667), .ZN(n10593) );
  AND3_X1 U5114 ( .A1(n6537), .A2(n6536), .A3(n6535), .ZN(n7725) );
  CLKBUF_X3 U5115 ( .A(n5686), .Z(n6221) );
  NAND2_X1 U5116 ( .A1(n10274), .A2(n10273), .ZN(n10296) );
  OAI211_X1 U5117 ( .C1(n6509), .C2(P2_REG3_REG_3__SCAN_IN), .A(n5339), .B(
        n6530), .ZN(n9290) );
  INV_X1 U5118 ( .A(n5625), .ZN(n5686) );
  AND3_X1 U5119 ( .A1(n5648), .A2(n5647), .A3(n5646), .ZN(n6971) );
  OAI211_X1 U5120 ( .C1(n6756), .C2(n7439), .A(n6523), .B(n6522), .ZN(n7558)
         );
  INV_X1 U5121 ( .A(n5420), .ZN(n5419) );
  CLKBUF_X1 U5122 ( .A(n8848), .Z(n8844) );
  NAND2_X2 U5123 ( .A1(n6141), .A2(n6140), .ZN(n6951) );
  INV_X2 U5124 ( .A(n6756), .ZN(n8849) );
  AND2_X1 U5125 ( .A1(n6486), .A2(n6485), .ZN(n6527) );
  OAI21_X1 U5126 ( .B1(n5428), .B2(n5421), .A(n5564), .ZN(n5420) );
  MUX2_X1 U5127 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5591), .S(
        P1_IR_REG_29__SCAN_IN), .Z(n5594) );
  NAND2_X1 U5128 ( .A1(n5595), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5597) );
  NAND2_X2 U5129 ( .A1(n6515), .A2(n7427), .ZN(n6756) );
  INV_X1 U5130 ( .A(n5422), .ZN(n5421) );
  AND2_X1 U5131 ( .A1(n6515), .A2(n7435), .ZN(n6667) );
  XNOR2_X1 U5132 ( .A(n6124), .B(n6123), .ZN(n8733) );
  XNOR2_X1 U5133 ( .A(n6142), .B(P1_IR_REG_22__SCAN_IN), .ZN(n6065) );
  MUX2_X1 U5134 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6482), .S(
        P2_IR_REG_29__SCAN_IN), .Z(n6484) );
  NAND2_X1 U5135 ( .A1(n6495), .A2(n6494), .ZN(n6845) );
  MUX2_X1 U5136 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6497), .S(
        P2_IR_REG_27__SCAN_IN), .Z(n6499) );
  MUX2_X1 U5137 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6493), .S(
        P2_IR_REG_28__SCAN_IN), .Z(n6495) );
  NAND2_X1 U5138 ( .A1(n6120), .A2(n6123), .ZN(n5589) );
  NAND2_X1 U5139 ( .A1(n6728), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6829) );
  INV_X1 U5140 ( .A(n5733), .ZN(n5573) );
  AND2_X1 U5141 ( .A1(n5191), .A2(n5579), .ZN(n5190) );
  NAND2_X2 U5142 ( .A1(n7427), .A2(P2_U3151), .ZN(n9676) );
  AND2_X2 U5143 ( .A1(n6713), .A2(n6476), .ZN(n6727) );
  NAND2_X1 U5144 ( .A1(n5519), .A2(SI_2_), .ZN(n5527) );
  INV_X1 U5145 ( .A(n5528), .ZN(n7427) );
  NOR2_X1 U5146 ( .A1(n5445), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n5083) );
  NOR2_X1 U5147 ( .A1(n5501), .A2(n4972), .ZN(n5499) );
  NAND4_X1 U5148 ( .A1(n6474), .A2(n6473), .A3(n6472), .A4(n6471), .ZN(n6592)
         );
  NAND2_X1 U5149 ( .A1(n5570), .A2(n5446), .ZN(n5445) );
  INV_X1 U5150 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n5869) );
  INV_X1 U5151 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n9920) );
  INV_X1 U5152 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n5867) );
  INV_X1 U5153 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n5866) );
  NOR2_X1 U5154 ( .A1(P2_IR_REG_23__SCAN_IN), .A2(P2_IR_REG_22__SCAN_IN), .ZN(
        n5502) );
  INV_X1 U5155 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n5596) );
  NOR2_X1 U5156 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n5569) );
  INV_X4 U5157 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  NOR3_X1 U5158 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), .A3(
        P2_IR_REG_21__SCAN_IN), .ZN(n6477) );
  INV_X1 U5159 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n5446) );
  INV_X1 U5160 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n5570) );
  NOR2_X1 U5161 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n6465) );
  NOR2_X1 U5162 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), .ZN(
        n6466) );
  NOR2_X1 U5163 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n5871) );
  NOR2_X1 U5164 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n5868) );
  NOR2_X1 U5165 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n6473) );
  NOR2_X1 U5166 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), .ZN(
        n6474) );
  AND4_X4 U5167 ( .A1(n6505), .A2(n6504), .A3(n6503), .A4(n6502), .ZN(n7503)
         );
  INV_X1 U5168 ( .A(n6509), .ZN(n6519) );
  INV_X2 U5169 ( .A(n5618), .ZN(n5645) );
  OAI21_X1 U5170 ( .B1(n9046), .B2(n4992), .A(n5224), .ZN(n5223) );
  INV_X2 U5171 ( .A(n7503), .ZN(n7527) );
  OAI21_X2 U5172 ( .B1(n6919), .B2(n9116), .A(n6918), .ZN(n8861) );
  NAND2_X1 U5173 ( .A1(n8062), .A2(n8885), .ZN(n8295) );
  AOI21_X2 U5174 ( .B1(n8295), .B2(n6858), .A(n8918), .ZN(n8194) );
  OR2_X1 U5175 ( .A1(n6322), .A2(n5082), .ZN(n6330) );
  OR2_X1 U5176 ( .A1(n6321), .A2(n6339), .ZN(n5082) );
  NAND2_X1 U5177 ( .A1(n6239), .A2(n8173), .ZN(n6079) );
  NAND2_X1 U5178 ( .A1(n6166), .A2(n6165), .ZN(n6196) );
  NOR2_X1 U5179 ( .A1(n9492), .A2(n5323), .ZN(n5322) );
  INV_X1 U5180 ( .A(n9015), .ZN(n5323) );
  OR2_X1 U5181 ( .A1(n10131), .A2(n10144), .ZN(n6300) );
  NAND2_X1 U5182 ( .A1(n6070), .A2(n7176), .ZN(n6948) );
  XNOR2_X1 U5183 ( .A(n5886), .B(n5865), .ZN(n5887) );
  OR2_X1 U5184 ( .A1(n6813), .A2(n6814), .ZN(n5505) );
  NAND2_X1 U5185 ( .A1(n5461), .A2(n5460), .ZN(n10077) );
  AOI21_X1 U5186 ( .B1(n5465), .B2(n5463), .A(n4962), .ZN(n5460) );
  NAND2_X1 U5187 ( .A1(n5080), .A2(n6359), .ZN(n5079) );
  NAND2_X1 U5188 ( .A1(n6331), .A2(n5081), .ZN(n5080) );
  OAI21_X1 U5189 ( .B1(n6330), .B2(n6324), .A(n6323), .ZN(n5081) );
  NAND3_X1 U5190 ( .A1(n9920), .A2(n5397), .A3(n5398), .ZN(n5396) );
  INV_X1 U5191 ( .A(P1_RD_REG_SCAN_IN), .ZN(n5397) );
  NAND2_X1 U5192 ( .A1(n10423), .A2(n5182), .ZN(n7248) );
  OR2_X1 U5193 ( .A1(n10414), .A2(n7247), .ZN(n5182) );
  NOR2_X1 U5194 ( .A1(n10419), .A2(n7212), .ZN(n7213) );
  NOR2_X1 U5195 ( .A1(n10414), .A2(n7965), .ZN(n7212) );
  NOR2_X1 U5196 ( .A1(n9538), .A2(n4967), .ZN(n5264) );
  NOR2_X1 U5197 ( .A1(n4967), .A2(n5266), .ZN(n5265) );
  INV_X1 U5198 ( .A(n6700), .ZN(n5266) );
  OAI21_X1 U5199 ( .B1(n6928), .B2(n5250), .A(n5249), .ZN(n5248) );
  NAND2_X1 U5200 ( .A1(n6927), .A2(n5251), .ZN(n5180) );
  NOR2_X1 U5201 ( .A1(n4951), .A2(n5258), .ZN(n5250) );
  OR2_X1 U5202 ( .A1(n6927), .A2(n5253), .ZN(n5252) );
  NAND2_X1 U5203 ( .A1(n6928), .A2(n4951), .ZN(n5253) );
  AOI21_X2 U5204 ( .B1(n5256), .B2(n5255), .A(n6935), .ZN(n5254) );
  INV_X1 U5205 ( .A(n7775), .ZN(n5255) );
  AND2_X1 U5206 ( .A1(n9215), .A2(n9446), .ZN(n6788) );
  NAND2_X1 U5207 ( .A1(n9643), .A2(n9165), .ZN(n6789) );
  INV_X1 U5208 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n6476) );
  INV_X1 U5209 ( .A(n5303), .ZN(n5299) );
  AND2_X1 U5210 ( .A1(n6951), .A2(n6947), .ZN(n7018) );
  INV_X1 U5211 ( .A(n7025), .ZN(n5041) );
  AND2_X1 U5212 ( .A1(n5038), .A2(n5286), .ZN(n5037) );
  NAND2_X1 U5213 ( .A1(n5040), .A2(n7026), .ZN(n5038) );
  INV_X1 U5214 ( .A(n5287), .ZN(n5286) );
  OAI21_X1 U5215 ( .B1(n5290), .B2(n5288), .A(n8765), .ZN(n5287) );
  OAI21_X1 U5216 ( .B1(n8847), .B2(n5406), .A(n5404), .ZN(n6341) );
  NOR2_X1 U5217 ( .A1(n5408), .A2(n5405), .ZN(n5404) );
  NOR2_X1 U5218 ( .A1(n5406), .A2(n6217), .ZN(n5405) );
  AND2_X1 U5219 ( .A1(n5408), .A2(n6211), .ZN(n5402) );
  OR2_X1 U5220 ( .A1(n10161), .A2(n8281), .ZN(n6367) );
  NOR2_X1 U5221 ( .A1(n10161), .A2(n5197), .ZN(n5196) );
  INV_X1 U5222 ( .A(n5198), .ZN(n5197) );
  OR2_X1 U5223 ( .A1(n10249), .A2(n9996), .ZN(n6359) );
  OR2_X1 U5224 ( .A1(n10222), .A2(n10125), .ZN(n6297) );
  OR2_X1 U5225 ( .A1(n8665), .A2(n8763), .ZN(n6282) );
  INV_X1 U5226 ( .A(n6079), .ZN(n5342) );
  NAND2_X1 U5227 ( .A1(n6162), .A2(n6161), .ZN(n6176) );
  INV_X1 U5228 ( .A(n5733), .ZN(n5875) );
  NOR2_X1 U5229 ( .A1(n5873), .A2(n5872), .ZN(n5874) );
  INV_X1 U5230 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n5899) );
  NAND2_X1 U5231 ( .A1(n5725), .A2(n4986), .ZN(n5205) );
  INV_X1 U5232 ( .A(n7709), .ZN(n7708) );
  OR2_X1 U5233 ( .A1(n6750), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n6759) );
  NAND2_X1 U5234 ( .A1(n9185), .A2(n9186), .ZN(n5479) );
  XNOR2_X1 U5235 ( .A(n7210), .B(n10404), .ZN(n10401) );
  INV_X1 U5236 ( .A(n7210), .ZN(n7209) );
  INV_X1 U5237 ( .A(n6846), .ZN(n7271) );
  OAI21_X1 U5238 ( .B1(n9417), .B2(n4958), .A(n4998), .ZN(n5237) );
  AOI21_X1 U5239 ( .B1(n8899), .B2(n5268), .A(n9027), .ZN(n5280) );
  INV_X1 U5240 ( .A(n6747), .ZN(n5268) );
  AOI21_X1 U5241 ( .B1(n5319), .B2(n5321), .A(n4991), .ZN(n5317) );
  NOR2_X1 U5242 ( .A1(n9497), .A2(n6738), .ZN(n9483) );
  AND2_X1 U5243 ( .A1(n9169), .A2(n9484), .ZN(n6738) );
  AND2_X1 U5244 ( .A1(n5302), .A2(n9728), .ZN(n5301) );
  NAND2_X1 U5245 ( .A1(n9679), .A2(n5303), .ZN(n5302) );
  AND2_X1 U5246 ( .A1(n7836), .A2(n7837), .ZN(n5284) );
  AND2_X1 U5247 ( .A1(n9696), .A2(n5013), .ZN(n9746) );
  NAND2_X1 U5248 ( .A1(n6069), .A2(n6068), .ZN(n7176) );
  OAI21_X1 U5249 ( .B1(n6031), .B2(n5443), .A(n4961), .ZN(n5444) );
  INV_X1 U5250 ( .A(n7353), .ZN(n5443) );
  NAND2_X1 U5251 ( .A1(n7353), .A2(n5442), .ZN(n5441) );
  NAND2_X1 U5252 ( .A1(n5444), .A2(n7360), .ZN(n9944) );
  NAND2_X1 U5253 ( .A1(n10123), .A2(n10121), .ZN(n6098) );
  AOI21_X1 U5254 ( .B1(n5467), .B2(n5469), .A(n5001), .ZN(n5466) );
  AND2_X1 U5255 ( .A1(n10222), .A2(n9723), .ZN(n5469) );
  OR2_X1 U5256 ( .A1(n4978), .A2(n5581), .ZN(n5439) );
  OR2_X1 U5257 ( .A1(n6116), .A2(n4978), .ZN(n5438) );
  NAND2_X1 U5258 ( .A1(n6072), .A2(n7176), .ZN(n7854) );
  XNOR2_X1 U5259 ( .A(n6118), .B(P1_IR_REG_26__SCAN_IN), .ZN(n6141) );
  NAND2_X1 U5260 ( .A1(n6117), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6118) );
  NAND2_X1 U5261 ( .A1(n5409), .A2(n5414), .ZN(n5888) );
  NAND2_X1 U5262 ( .A1(n5831), .A2(n5410), .ZN(n5409) );
  INV_X1 U5263 ( .A(n5416), .ZN(n5410) );
  NAND2_X1 U5264 ( .A1(n5849), .A2(n5848), .ZN(n5864) );
  NAND2_X1 U5265 ( .A1(n9172), .A2(n9171), .ZN(n9170) );
  NAND2_X1 U5266 ( .A1(n5378), .A2(n5377), .ZN(n9310) );
  NAND2_X1 U5267 ( .A1(n7223), .A2(n5382), .ZN(n5377) );
  OR2_X1 U5268 ( .A1(n9294), .A2(n5379), .ZN(n5378) );
  NAND2_X1 U5269 ( .A1(n5382), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n5379) );
  AOI21_X1 U5270 ( .B1(n6849), .B2(n9532), .A(n6848), .ZN(n9147) );
  AOI21_X1 U5271 ( .B1(n8913), .B2(n8919), .A(n9060), .ZN(n5221) );
  NAND2_X1 U5272 ( .A1(n6239), .A2(n6401), .ZN(n6268) );
  NOR2_X1 U5273 ( .A1(n5225), .A2(n9412), .ZN(n5224) );
  INV_X1 U5274 ( .A(n9051), .ZN(n5225) );
  OR2_X1 U5275 ( .A1(n9083), .A2(n9617), .ZN(n8990) );
  NOR2_X1 U5276 ( .A1(n8359), .A2(n8353), .ZN(n8960) );
  NOR2_X1 U5277 ( .A1(n10637), .A2(n8192), .ZN(n8914) );
  INV_X1 U5278 ( .A(n5289), .ZN(n5288) );
  OAI211_X1 U5279 ( .C1(n6333), .C2(n5370), .A(n7356), .B(n6332), .ZN(n6335)
         );
  NAND2_X1 U5280 ( .A1(n5079), .A2(n5077), .ZN(n6333) );
  NAND2_X1 U5281 ( .A1(n5078), .A2(n6339), .ZN(n5077) );
  NAND2_X1 U5282 ( .A1(n6338), .A2(n6337), .ZN(n5051) );
  OR2_X1 U5283 ( .A1(n9124), .A2(n9939), .ZN(n6228) );
  INV_X1 U5284 ( .A(n7945), .ZN(n6087) );
  NAND2_X1 U5285 ( .A1(n6061), .A2(n5085), .ZN(n5310) );
  INV_X1 U5286 ( .A(SI_16_), .ZN(n8535) );
  INV_X1 U5287 ( .A(n5568), .ZN(n5178) );
  XNOR2_X1 U5288 ( .A(n7523), .B(n7551), .ZN(n7504) );
  INV_X1 U5289 ( .A(n8001), .ZN(n5484) );
  INV_X1 U5290 ( .A(n8126), .ZN(n5132) );
  INV_X1 U5291 ( .A(n9664), .ZN(n6486) );
  NOR2_X1 U5292 ( .A1(n10456), .A2(n5091), .ZN(n7216) );
  NOR2_X1 U5293 ( .A1(n10447), .A2(n5092), .ZN(n5091) );
  AOI21_X1 U5294 ( .B1(P2_REG1_REG_10__SCAN_IN), .B2(n7463), .A(n10488), .ZN(
        n7219) );
  NAND2_X1 U5295 ( .A1(n8628), .A2(n7256), .ZN(n7257) );
  OR2_X1 U5296 ( .A1(n9555), .A2(n6814), .ZN(n8870) );
  INV_X1 U5297 ( .A(n5327), .ZN(n5158) );
  INV_X1 U5298 ( .A(n5328), .ZN(n5326) );
  NAND2_X1 U5299 ( .A1(n6463), .A2(n8596), .ZN(n6795) );
  INV_X1 U5300 ( .A(n6781), .ZN(n6463) );
  INV_X1 U5301 ( .A(n9034), .ZN(n5274) );
  NOR2_X1 U5302 ( .A1(n5277), .A2(n9034), .ZN(n5272) );
  INV_X1 U5303 ( .A(n6741), .ZN(n6460) );
  OR2_X1 U5304 ( .A1(n9524), .A2(n9604), .ZN(n9007) );
  NAND2_X1 U5305 ( .A1(n8773), .A2(n8993), .ZN(n5267) );
  INV_X1 U5306 ( .A(n6866), .ZN(n5316) );
  OR2_X1 U5307 ( .A1(n8987), .A2(n5316), .ZN(n5315) );
  OR2_X1 U5308 ( .A1(n9611), .A2(n9264), .ZN(n8998) );
  INV_X1 U5309 ( .A(n6663), .ZN(n5236) );
  AND2_X1 U5310 ( .A1(n8990), .A2(n8989), .ZN(n8894) );
  INV_X1 U5311 ( .A(n8960), .ZN(n6860) );
  NOR2_X1 U5312 ( .A1(n8241), .A2(n8267), .ZN(n8961) );
  NAND2_X1 U5313 ( .A1(n5246), .A2(n5245), .ZN(n5244) );
  NAND2_X1 U5314 ( .A1(n7523), .A2(n7503), .ZN(n8928) );
  OR2_X1 U5315 ( .A1(n9145), .A2(n9408), .ZN(n6915) );
  INV_X1 U5316 ( .A(n5012), .ZN(n5300) );
  NAND2_X1 U5317 ( .A1(n6983), .A2(n7831), .ZN(n5067) );
  NAND2_X1 U5318 ( .A1(n5075), .A2(n9720), .ZN(n5074) );
  INV_X1 U5319 ( .A(n7080), .ZN(n5075) );
  INV_X1 U5320 ( .A(n9720), .ZN(n5076) );
  NAND2_X1 U5321 ( .A1(n4989), .A2(n5401), .ZN(n5400) );
  INV_X1 U5322 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n6066) );
  NAND2_X1 U5323 ( .A1(n5369), .A2(n9980), .ZN(n5365) );
  OR2_X1 U5324 ( .A1(n7329), .A2(n9984), .ZN(n7358) );
  OR2_X1 U5325 ( .A1(n10174), .A2(n10015), .ZN(n6029) );
  OR2_X1 U5326 ( .A1(n10174), .A2(n9732), .ZN(n6358) );
  AND2_X1 U5327 ( .A1(n6427), .A2(n6426), .ZN(n5362) );
  OR2_X1 U5328 ( .A1(n10070), .A2(n10081), .ZN(n6427) );
  OR2_X1 U5329 ( .A1(n10200), .A2(n10097), .ZN(n6426) );
  OR2_X1 U5330 ( .A1(n10210), .A2(n10124), .ZN(n6421) );
  INV_X1 U5331 ( .A(n8809), .ZN(n6096) );
  NAND2_X1 U5332 ( .A1(n5341), .A2(n5340), .ZN(n6082) );
  NOR2_X1 U5333 ( .A1(n4945), .A2(n5449), .ZN(n5448) );
  NAND2_X1 U5334 ( .A1(n9808), .A2(n10613), .ZN(n6395) );
  NAND2_X1 U5335 ( .A1(n6447), .A2(n6070), .ZN(n6949) );
  INV_X1 U5336 ( .A(n10273), .ZN(n6138) );
  NAND2_X1 U5337 ( .A1(n6200), .A2(n6199), .ZN(n6216) );
  INV_X1 U5338 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n6076) );
  OAI21_X1 U5339 ( .B1(n6013), .B2(n5432), .A(n5430), .ZN(n6158) );
  INV_X1 U5340 ( .A(n5431), .ZN(n5430) );
  OAI21_X1 U5341 ( .B1(n5434), .B2(n5432), .A(n6047), .ZN(n5431) );
  INV_X1 U5342 ( .A(n5310), .ZN(n5308) );
  INV_X1 U5343 ( .A(SI_22_), .ZN(n8527) );
  NAND2_X1 U5344 ( .A1(n5875), .A2(n5874), .ZN(n5897) );
  NAND2_X1 U5345 ( .A1(n5642), .A2(n5527), .ZN(n5657) );
  NAND2_X1 U5346 ( .A1(n5170), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n5169) );
  NAND2_X1 U5347 ( .A1(n5166), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n5167) );
  INV_X1 U5348 ( .A(n5396), .ZN(n5166) );
  INV_X1 U5349 ( .A(n5167), .ZN(n5165) );
  NAND2_X1 U5350 ( .A1(n7873), .A2(n7872), .ZN(n7876) );
  NAND2_X1 U5351 ( .A1(n5476), .A2(n9155), .ZN(n5475) );
  INV_X1 U5352 ( .A(n5507), .ZN(n5476) );
  AND2_X1 U5353 ( .A1(n9111), .A2(n5014), .ZN(n5478) );
  OR2_X1 U5354 ( .A1(n9246), .A2(n9563), .ZN(n9111) );
  AOI21_X1 U5355 ( .B1(n5483), .B2(n7875), .A(n5482), .ZN(n5481) );
  INV_X1 U5356 ( .A(n8123), .ZN(n5482) );
  NAND2_X1 U5357 ( .A1(n5139), .A2(n4947), .ZN(n5137) );
  NAND2_X1 U5358 ( .A1(n4947), .A2(n9097), .ZN(n5138) );
  NAND2_X1 U5359 ( .A1(n7554), .A2(n7555), .ZN(n7675) );
  AND2_X1 U5360 ( .A1(n4973), .A2(n4953), .ZN(n5141) );
  NAND2_X1 U5361 ( .A1(n5145), .A2(n4985), .ZN(n5144) );
  NAND2_X1 U5362 ( .A1(n5146), .A2(n9192), .ZN(n5145) );
  NAND2_X1 U5363 ( .A1(n5127), .A2(n5470), .ZN(n7765) );
  INV_X1 U5364 ( .A(n5471), .ZN(n5127) );
  OAI21_X1 U5365 ( .B1(n7708), .B2(n5472), .A(n7732), .ZN(n5471) );
  AOI21_X1 U5366 ( .B1(n7294), .B2(n7432), .A(n7577), .ZN(n10363) );
  NAND2_X1 U5367 ( .A1(n10425), .A2(n10424), .ZN(n10423) );
  OR2_X1 U5368 ( .A1(n10401), .A2(n5006), .ZN(n5099) );
  INV_X1 U5369 ( .A(n10420), .ZN(n5101) );
  XNOR2_X1 U5370 ( .A(n7248), .B(n10431), .ZN(n10433) );
  XNOR2_X1 U5371 ( .A(n7213), .B(n10431), .ZN(n10441) );
  XNOR2_X1 U5372 ( .A(n7216), .B(n10463), .ZN(n10473) );
  NAND2_X1 U5373 ( .A1(n5383), .A2(n5090), .ZN(n10488) );
  NAND2_X1 U5374 ( .A1(n7217), .A2(n5387), .ZN(n5383) );
  OR2_X1 U5375 ( .A1(n10473), .A2(n5384), .ZN(n5090) );
  NAND2_X1 U5376 ( .A1(n5387), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n5384) );
  OR2_X1 U5377 ( .A1(n10473), .A2(n10472), .ZN(n5386) );
  NAND2_X1 U5378 ( .A1(n10484), .A2(n10485), .ZN(n10483) );
  NAND2_X1 U5379 ( .A1(n8633), .A2(n8634), .ZN(n8632) );
  NAND2_X1 U5380 ( .A1(n8629), .A2(n8630), .ZN(n8628) );
  XNOR2_X1 U5381 ( .A(n7219), .B(n10496), .ZN(n10509) );
  XNOR2_X1 U5382 ( .A(n7257), .B(n7279), .ZN(n9297) );
  NOR2_X1 U5383 ( .A1(n8626), .A2(n5093), .ZN(n7222) );
  NOR2_X1 U5384 ( .A1(n7281), .A2(n5094), .ZN(n5093) );
  NAND2_X1 U5385 ( .A1(n9351), .A2(n9352), .ZN(n9350) );
  INV_X1 U5386 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n5398) );
  NAND2_X1 U5387 ( .A1(n9364), .A2(n7264), .ZN(n9382) );
  OR2_X1 U5388 ( .A1(n9252), .A2(n9245), .ZN(n9409) );
  OR2_X1 U5389 ( .A1(n9564), .A2(n9275), .ZN(n5238) );
  NAND2_X1 U5390 ( .A1(n9427), .A2(n4988), .ZN(n5239) );
  NAND2_X1 U5391 ( .A1(n8872), .A2(n5329), .ZN(n5328) );
  NAND2_X1 U5392 ( .A1(n4965), .A2(n9038), .ZN(n5329) );
  NOR2_X1 U5393 ( .A1(n9039), .A2(n9453), .ZN(n5331) );
  AND2_X1 U5394 ( .A1(n5280), .A2(n8874), .ZN(n5277) );
  INV_X1 U5395 ( .A(n5278), .ZN(n5276) );
  AOI21_X1 U5396 ( .B1(n5280), .B2(n9478), .A(n5279), .ZN(n5278) );
  INV_X1 U5397 ( .A(n8873), .ZN(n5279) );
  AND2_X1 U5398 ( .A1(n6868), .A2(n5320), .ZN(n5319) );
  NAND2_X1 U5399 ( .A1(n5322), .A2(n9092), .ZN(n5320) );
  INV_X1 U5400 ( .A(n5322), .ZN(n5321) );
  OR2_X1 U5401 ( .A1(n9586), .A2(n9468), .ZN(n6747) );
  NAND2_X1 U5402 ( .A1(n9503), .A2(n9015), .ZN(n9491) );
  INV_X1 U5403 ( .A(n9017), .ZN(n9492) );
  OR2_X1 U5404 ( .A1(n9524), .A2(n9277), .ZN(n6725) );
  INV_X1 U5405 ( .A(n5263), .ZN(n5262) );
  INV_X1 U5406 ( .A(n8894), .ZN(n8983) );
  OAI21_X1 U5407 ( .B1(n8386), .B2(n8385), .A(n6651), .ZN(n8696) );
  OR2_X1 U5408 ( .A1(n6645), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n6657) );
  NAND2_X1 U5409 ( .A1(n8194), .A2(n8891), .ZN(n5338) );
  OR2_X1 U5410 ( .A1(n6595), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n6613) );
  NOR2_X1 U5411 ( .A1(n7963), .A2(n6575), .ZN(n5246) );
  NAND2_X1 U5412 ( .A1(n7963), .A2(n6575), .ZN(n5245) );
  OAI22_X1 U5413 ( .A1(n7726), .A2(n6538), .B1(n7725), .B2(n7792), .ZN(n7791)
         );
  NAND2_X1 U5414 ( .A1(n7792), .A2(n7783), .ZN(n8943) );
  AND2_X1 U5415 ( .A1(n8943), .A2(n8936), .ZN(n8875) );
  INV_X1 U5416 ( .A(n9515), .ZN(n9534) );
  NAND2_X1 U5417 ( .A1(n5247), .A2(n5179), .ZN(n8843) );
  NAND2_X1 U5418 ( .A1(n5254), .A2(n9498), .ZN(n5247) );
  INV_X1 U5419 ( .A(n9609), .ZN(n9616) );
  NOR2_X1 U5420 ( .A1(n6940), .A2(n9618), .ZN(n7514) );
  NAND2_X1 U5421 ( .A1(n6887), .A2(n6886), .ZN(n7339) );
  INV_X1 U5422 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5335) );
  INV_X1 U5423 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n6872) );
  NAND2_X1 U5424 ( .A1(n6878), .A2(n6872), .ZN(n6874) );
  NAND2_X1 U5425 ( .A1(n5152), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6878) );
  NAND2_X1 U5426 ( .A1(n6727), .A2(n5500), .ZN(n5152) );
  INV_X1 U5427 ( .A(n5501), .ZN(n5500) );
  XNOR2_X1 U5428 ( .A(n6837), .B(P2_IR_REG_22__SCAN_IN), .ZN(n9078) );
  NAND2_X1 U5429 ( .A1(n6830), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6835) );
  INV_X1 U5430 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n6828) );
  INV_X1 U5431 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n6834) );
  AND2_X1 U5432 ( .A1(n6571), .A2(n6559), .ZN(n7290) );
  NOR2_X1 U5433 ( .A1(n4956), .A2(n4983), .ZN(n5062) );
  OR3_X1 U5434 ( .A1(n9751), .A2(n9746), .A3(n4959), .ZN(n5298) );
  INV_X1 U5435 ( .A(n8827), .ZN(n5304) );
  NOR2_X1 U5436 ( .A1(n7068), .A2(n8827), .ZN(n5305) );
  AOI21_X1 U5437 ( .B1(n5037), .B2(n5039), .A(n5000), .ZN(n5035) );
  INV_X1 U5438 ( .A(n5037), .ZN(n5036) );
  NAND2_X1 U5439 ( .A1(n8335), .A2(n8336), .ZN(n5289) );
  OR2_X1 U5440 ( .A1(n8335), .A2(n8336), .ZN(n5290) );
  AND2_X1 U5441 ( .A1(n6978), .A2(n6979), .ZN(n9763) );
  OAI211_X1 U5442 ( .C1(n5284), .C2(n5283), .A(n5281), .B(n6997), .ZN(n8048)
         );
  INV_X1 U5443 ( .A(n6994), .ZN(n5283) );
  NAND2_X1 U5444 ( .A1(n5292), .A2(n5291), .ZN(n9780) );
  NAND2_X1 U5445 ( .A1(n5294), .A2(n5296), .ZN(n5291) );
  NAND2_X1 U5446 ( .A1(n9678), .A2(n5293), .ZN(n5292) );
  NAND2_X1 U5447 ( .A1(n5030), .A2(n7062), .ZN(n8816) );
  INV_X1 U5448 ( .A(n7060), .ZN(n5030) );
  AOI21_X1 U5449 ( .B1(n5046), .B2(n6341), .A(n5045), .ZN(n6378) );
  AND2_X1 U5450 ( .A1(n6340), .A2(n6339), .ZN(n5045) );
  NAND2_X1 U5451 ( .A1(n5048), .A2(n5047), .ZN(n5046) );
  AOI21_X1 U5452 ( .B1(n6371), .B2(n6370), .A(n6435), .ZN(n6373) );
  AOI21_X1 U5453 ( .B1(n8229), .B2(P1_REG2_REG_14__SCAN_IN), .A(n8223), .ZN(
        n9865) );
  NAND2_X1 U5454 ( .A1(n6169), .A2(n6168), .ZN(n10161) );
  AND4_X1 U5455 ( .A1(n6043), .A2(n6042), .A3(n6041), .A4(n6040), .ZN(n9996)
         );
  AND2_X1 U5456 ( .A1(n10013), .A2(n6351), .ZN(n5121) );
  NOR2_X1 U5457 ( .A1(n10027), .A2(n5120), .ZN(n10014) );
  INV_X1 U5458 ( .A(n6351), .ZN(n5120) );
  NAND2_X1 U5459 ( .A1(n6354), .A2(n6355), .ZN(n10010) );
  AND4_X1 U5460 ( .A1(n6004), .A2(n6003), .A3(n6002), .A4(n6001), .ZN(n10031)
         );
  OR2_X1 U5461 ( .A1(n10190), .A2(n10065), .ZN(n6230) );
  AND2_X1 U5462 ( .A1(n10041), .A2(n4966), .ZN(n5456) );
  AND2_X1 U5463 ( .A1(n6427), .A2(n6313), .ZN(n10062) );
  OR2_X1 U5464 ( .A1(n10058), .A2(n10062), .ZN(n5457) );
  NAND2_X1 U5465 ( .A1(n10093), .A2(n6423), .ZN(n10079) );
  OAI21_X1 U5466 ( .B1(n5466), .B2(n10108), .A(n4996), .ZN(n5465) );
  NOR2_X1 U5467 ( .A1(n5468), .A2(n10121), .ZN(n5467) );
  NOR2_X1 U5468 ( .A1(n10137), .A2(n5469), .ZN(n5468) );
  NAND2_X1 U5469 ( .A1(n5349), .A2(n6096), .ZN(n5351) );
  NAND2_X1 U5470 ( .A1(n5350), .A2(n5349), .ZN(n5348) );
  INV_X1 U5471 ( .A(n6280), .ZN(n5350) );
  INV_X1 U5472 ( .A(n5361), .ZN(n5358) );
  AOI21_X1 U5473 ( .B1(n5361), .B2(n5122), .A(n5357), .ZN(n5356) );
  INV_X1 U5474 ( .A(n6284), .ZN(n5357) );
  INV_X1 U5475 ( .A(n8660), .ZN(n5360) );
  INV_X1 U5476 ( .A(n6282), .ZN(n5359) );
  AND2_X1 U5477 ( .A1(n8687), .A2(n6282), .ZN(n5361) );
  AND2_X1 U5478 ( .A1(n6408), .A2(n6284), .ZN(n8687) );
  NAND2_X1 U5479 ( .A1(n8662), .A2(n8661), .ZN(n8660) );
  INV_X1 U5480 ( .A(n5122), .ZN(n8661) );
  OR2_X1 U5481 ( .A1(n8771), .A2(n9804), .ZN(n5786) );
  INV_X1 U5482 ( .A(n5660), .ZN(n5902) );
  OR2_X1 U5483 ( .A1(n5757), .A2(n5343), .ZN(n5758) );
  OR2_X1 U5484 ( .A1(n8167), .A2(n8176), .ZN(n8173) );
  NAND2_X1 U5485 ( .A1(n8135), .A2(n8137), .ZN(n8134) );
  AND4_X1 U5486 ( .A1(n5721), .A2(n5720), .A3(n5719), .A4(n5718), .ZN(n8029)
         );
  NAND2_X1 U5487 ( .A1(n9821), .A2(n7398), .ZN(n10145) );
  OAI211_X1 U5488 ( .C1(n6018), .C2(n7445), .A(n5666), .B(n5665), .ZN(n5667)
         );
  XNOR2_X1 U5489 ( .A(n6970), .B(n6971), .ZN(n10549) );
  OR2_X1 U5490 ( .A1(n10663), .A2(n6070), .ZN(n7178) );
  INV_X1 U5491 ( .A(n10145), .ZN(n10558) );
  NOR2_X1 U5492 ( .A1(n7932), .A2(n7857), .ZN(n7863) );
  OR2_X1 U5493 ( .A1(n10163), .A2(n10162), .ZN(n5512) );
  XNOR2_X1 U5494 ( .A(n6176), .B(n6177), .ZN(n9669) );
  XNOR2_X1 U5495 ( .A(n6158), .B(n6157), .ZN(n9672) );
  NAND2_X1 U5496 ( .A1(n6033), .A2(n6032), .ZN(n6049) );
  NOR2_X1 U5497 ( .A1(n5458), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n5191) );
  XNOR2_X1 U5498 ( .A(n6144), .B(n6143), .ZN(n7397) );
  OAI21_X1 U5499 ( .B1(n6142), .B2(P1_IR_REG_22__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n6144) );
  NAND2_X1 U5500 ( .A1(n5086), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5900) );
  NAND2_X1 U5501 ( .A1(n5900), .A2(n5899), .ZN(n5914) );
  NAND2_X1 U5502 ( .A1(n5172), .A2(n5171), .ZN(n5849) );
  AND2_X1 U5503 ( .A1(n5174), .A2(n5418), .ZN(n5171) );
  NOR2_X1 U5504 ( .A1(n5787), .A2(n5423), .ZN(n5422) );
  INV_X1 U5505 ( .A(n5425), .ZN(n5423) );
  NAND2_X1 U5506 ( .A1(n5107), .A2(n5105), .ZN(n5424) );
  AOI21_X1 U5507 ( .B1(n5111), .B2(n5115), .A(n5106), .ZN(n5105) );
  INV_X1 U5508 ( .A(n5428), .ZN(n5106) );
  NAND2_X1 U5509 ( .A1(n5427), .A2(n5426), .ZN(n5425) );
  INV_X1 U5510 ( .A(n5562), .ZN(n5427) );
  NOR2_X1 U5511 ( .A1(n5114), .A2(n5556), .ZN(n5113) );
  NAND2_X1 U5512 ( .A1(n5725), .A2(n5550), .ZN(n5732) );
  INV_X1 U5513 ( .A(n5530), .ZN(n5531) );
  NAND2_X1 U5514 ( .A1(n5657), .A2(n5656), .ZN(n5659) );
  NAND2_X1 U5515 ( .A1(n6669), .A2(n6668), .ZN(n8728) );
  NAND3_X1 U5516 ( .A1(n7675), .A2(n7674), .A3(n7678), .ZN(n7707) );
  INV_X1 U5517 ( .A(n7677), .ZN(n7678) );
  OR2_X1 U5518 ( .A1(n9090), .A2(n9604), .ZN(n9091) );
  INV_X1 U5519 ( .A(n9280), .ZN(n8718) );
  OAI22_X1 U5520 ( .A1(n9210), .A2(n9211), .B1(n9108), .B2(n9446), .ZN(n9185)
         );
  NAND2_X1 U5521 ( .A1(n6706), .A2(n6705), .ZN(n9602) );
  INV_X1 U5522 ( .A(n9275), .ZN(n9438) );
  NAND2_X1 U5523 ( .A1(n5147), .A2(n7731), .ZN(n7709) );
  AND2_X1 U5524 ( .A1(n6775), .A2(n6774), .ZN(n9459) );
  INV_X1 U5525 ( .A(n9408), .ZN(n9554) );
  INV_X1 U5526 ( .A(n9459), .ZN(n9276) );
  OAI211_X1 U5527 ( .C1(n6842), .C2(n9474), .A(n6753), .B(n6752), .ZN(n9585)
         );
  XNOR2_X1 U5528 ( .A(n6572), .B(P2_IR_REG_6__SCAN_IN), .ZN(n10414) );
  XNOR2_X1 U5529 ( .A(n7222), .B(n7279), .ZN(n9294) );
  OR2_X1 U5530 ( .A1(n9294), .A2(n9295), .ZN(n5381) );
  OAI211_X1 U5531 ( .C1(n9310), .C2(n5027), .A(n5103), .B(n5102), .ZN(n9328)
         );
  NAND2_X1 U5532 ( .A1(n5021), .A2(n5104), .ZN(n5103) );
  NAND2_X1 U5533 ( .A1(n9310), .A2(n5104), .ZN(n5102) );
  NOR2_X1 U5534 ( .A1(n9328), .A2(n9329), .ZN(n9327) );
  AOI21_X1 U5535 ( .B1(n9391), .B2(n9383), .A(n9385), .ZN(n7314) );
  AND2_X1 U5536 ( .A1(n10355), .A2(n9074), .ZN(n10370) );
  AND2_X1 U5537 ( .A1(n6921), .A2(n6920), .ZN(n8839) );
  OR2_X1 U5538 ( .A1(n9149), .A2(n10585), .ZN(n9509) );
  OR2_X1 U5539 ( .A1(n9142), .A2(n9615), .ZN(n6871) );
  INV_X1 U5540 ( .A(n9145), .ZN(n9052) );
  INV_X1 U5541 ( .A(n8799), .ZN(n7470) );
  NOR2_X1 U5542 ( .A1(n8759), .A2(n8733), .ZN(n6140) );
  AND2_X1 U5543 ( .A1(n7397), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7377) );
  NAND2_X1 U5544 ( .A1(n5042), .A2(n7025), .ZN(n8338) );
  NAND2_X1 U5545 ( .A1(n5044), .A2(n5043), .ZN(n5042) );
  INV_X1 U5546 ( .A(n8282), .ZN(n5044) );
  INV_X1 U5547 ( .A(n5058), .ZN(n5061) );
  OAI21_X1 U5548 ( .B1(n7692), .B2(n7691), .A(n7696), .ZN(n7698) );
  AND4_X1 U5549 ( .A1(n5885), .A2(n5884), .A3(n5883), .A4(n5882), .ZN(n10144)
         );
  NAND2_X1 U5550 ( .A1(n5853), .A2(n5852), .ZN(n10222) );
  AND2_X1 U5551 ( .A1(n7175), .A2(n7162), .ZN(n9784) );
  INV_X1 U5552 ( .A(n10125), .ZN(n9723) );
  NAND4_X1 U5553 ( .A1(n5674), .A2(n5673), .A3(n5672), .A4(n5671), .ZN(n6987)
         );
  NOR2_X1 U5554 ( .A1(n9915), .A2(n9914), .ZN(n9917) );
  INV_X1 U5555 ( .A(n6070), .ZN(n9923) );
  AOI21_X1 U5556 ( .B1(n5353), .B2(n10127), .A(n5352), .ZN(n9954) );
  NAND2_X1 U5557 ( .A1(n9944), .A2(n9943), .ZN(n9946) );
  NAND2_X1 U5558 ( .A1(n7366), .A2(n9795), .ZN(n9943) );
  OAI211_X1 U5559 ( .C1(n6018), .C2(n7443), .A(n5682), .B(n5681), .ZN(n8022)
         );
  OR2_X1 U5560 ( .A1(n10619), .A2(n7855), .ZN(n10573) );
  AND2_X1 U5561 ( .A1(n9964), .A2(n9956), .ZN(n7368) );
  INV_X1 U5562 ( .A(n8921), .ZN(n8924) );
  NAND2_X1 U5563 ( .A1(n5220), .A2(n5218), .ZN(n8915) );
  NAND2_X1 U5564 ( .A1(n8914), .A2(n9060), .ZN(n5218) );
  INV_X1 U5565 ( .A(n5221), .ZN(n5220) );
  NOR2_X1 U5566 ( .A1(n8975), .A2(n8974), .ZN(n5226) );
  INV_X1 U5567 ( .A(n6359), .ZN(n5078) );
  AND2_X1 U5568 ( .A1(n8397), .A2(n8388), .ZN(n8965) );
  NOR2_X1 U5569 ( .A1(n6928), .A2(n5258), .ZN(n5251) );
  NAND2_X1 U5570 ( .A1(n6928), .A2(n5257), .ZN(n5249) );
  INV_X1 U5571 ( .A(n8073), .ZN(n5340) );
  AND2_X1 U5572 ( .A1(n5203), .A2(n5202), .ZN(n5201) );
  NOR2_X1 U5573 ( .A1(n10200), .A2(n10102), .ZN(n5203) );
  NOR2_X1 U5574 ( .A1(n4944), .A2(n5757), .ZN(n5193) );
  INV_X1 U5575 ( .A(SI_28_), .ZN(n8418) );
  NAND2_X1 U5576 ( .A1(n5433), .A2(n6032), .ZN(n5432) );
  INV_X1 U5577 ( .A(n6048), .ZN(n5433) );
  INV_X1 U5578 ( .A(SI_27_), .ZN(n8523) );
  INV_X1 U5579 ( .A(SI_19_), .ZN(n8511) );
  INV_X1 U5580 ( .A(SI_20_), .ZN(n8512) );
  INV_X1 U5581 ( .A(n9086), .ZN(n5146) );
  NAND2_X1 U5582 ( .A1(n5223), .A2(n5222), .ZN(n9056) );
  INV_X1 U5583 ( .A(n9050), .ZN(n5222) );
  NAND2_X1 U5584 ( .A1(n7203), .A2(n7202), .ZN(n7204) );
  AND2_X1 U5585 ( .A1(n7562), .A2(n5394), .ZN(n7206) );
  NAND2_X1 U5586 ( .A1(n7432), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5394) );
  NAND2_X1 U5587 ( .A1(n5098), .A2(n7434), .ZN(n5097) );
  INV_X1 U5588 ( .A(n7206), .ZN(n5098) );
  OR2_X1 U5589 ( .A1(n10377), .A2(n7208), .ZN(n7210) );
  INV_X1 U5590 ( .A(n10489), .ZN(n5387) );
  NAND2_X1 U5591 ( .A1(n10448), .A2(n7250), .ZN(n7251) );
  OAI21_X1 U5592 ( .B1(n9373), .B2(n7310), .A(n9366), .ZN(n7313) );
  OR2_X1 U5593 ( .A1(n6805), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n6821) );
  AND2_X1 U5594 ( .A1(n9581), .A2(n9585), .ZN(n9029) );
  OR2_X1 U5595 ( .A1(n9169), .A2(n9517), .ZN(n9015) );
  OAI21_X1 U5596 ( .B1(n5264), .B2(n5265), .A(n5506), .ZN(n5263) );
  NOR2_X1 U5597 ( .A1(n8895), .A2(n5264), .ZN(n5260) );
  NAND2_X1 U5598 ( .A1(n6458), .A2(n9195), .ZN(n6707) );
  INV_X1 U5599 ( .A(n6694), .ZN(n6458) );
  NAND2_X1 U5600 ( .A1(n6456), .A2(n6455), .ZN(n6670) );
  INV_X1 U5601 ( .A(n6657), .ZN(n6456) );
  NOR2_X1 U5602 ( .A1(n6622), .A2(n8213), .ZN(n6623) );
  INV_X1 U5603 ( .A(n8965), .ZN(n6862) );
  NAND2_X1 U5604 ( .A1(n6454), .A2(n6453), .ZN(n6631) );
  INV_X1 U5605 ( .A(n6613), .ZN(n6454) );
  NAND2_X1 U5606 ( .A1(n8891), .A2(n6620), .ZN(n6621) );
  NAND2_X1 U5607 ( .A1(n8241), .A2(n8267), .ZN(n8919) );
  OR2_X1 U5608 ( .A1(n6565), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n6576) );
  NAND2_X1 U5609 ( .A1(n4975), .A2(n6548), .ZN(n5240) );
  OR2_X1 U5610 ( .A1(n9053), .A2(n6904), .ZN(n7489) );
  OR2_X1 U5611 ( .A1(n6884), .A2(n6898), .ZN(n7338) );
  NAND2_X1 U5612 ( .A1(n5513), .A2(n7544), .ZN(n8926) );
  INV_X1 U5613 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5336) );
  NAND2_X1 U5614 ( .A1(n6477), .A2(n5502), .ZN(n5501) );
  OR2_X1 U5615 ( .A1(n6641), .A2(P2_IR_REG_11__SCAN_IN), .ZN(n6642) );
  AND2_X1 U5616 ( .A1(n9739), .A2(n7101), .ZN(n5064) );
  INV_X1 U5617 ( .A(n7104), .ZN(n5065) );
  NAND2_X1 U5618 ( .A1(n9762), .A2(n6979), .ZN(n5058) );
  AND2_X1 U5619 ( .A1(n6994), .A2(n7811), .ZN(n5282) );
  NOR2_X1 U5620 ( .A1(n4959), .A2(n7149), .ZN(n5293) );
  INV_X1 U5621 ( .A(n9703), .ZN(n5297) );
  NAND2_X1 U5622 ( .A1(n5052), .A2(n5049), .ZN(n5048) );
  NOR2_X1 U5623 ( .A1(n5051), .A2(n5050), .ZN(n5049) );
  INV_X1 U5624 ( .A(n6336), .ZN(n5050) );
  AND2_X1 U5625 ( .A1(n5401), .A2(n4984), .ZN(n5047) );
  NOR2_X1 U5626 ( .A1(n7366), .A2(n7329), .ZN(n5198) );
  INV_X1 U5627 ( .A(n6030), .ZN(n5442) );
  OAI21_X1 U5628 ( .B1(n10044), .B2(n5119), .A(n5117), .ZN(n9992) );
  AOI21_X1 U5629 ( .B1(n5121), .B2(n5355), .A(n5118), .ZN(n5117) );
  INV_X1 U5630 ( .A(n5121), .ZN(n5119) );
  INV_X1 U5631 ( .A(n6354), .ZN(n5118) );
  NAND2_X1 U5632 ( .A1(n10181), .A2(n10031), .ZN(n6355) );
  AND2_X1 U5633 ( .A1(n4952), .A2(n5463), .ZN(n5462) );
  AND2_X1 U5634 ( .A1(n10146), .A2(n10268), .ZN(n10112) );
  INV_X1 U5635 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n5812) );
  OR2_X1 U5636 ( .A1(n5813), .A2(n5812), .ZN(n5815) );
  NAND2_X1 U5637 ( .A1(n6277), .A2(n6282), .ZN(n5122) );
  INV_X1 U5638 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5440) );
  NAND2_X1 U5639 ( .A1(n5032), .A2(n9805), .ZN(n6401) );
  INV_X1 U5640 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n5737) );
  OR2_X1 U5641 ( .A1(n5738), .A2(n5737), .ZN(n5751) );
  NOR2_X1 U5642 ( .A1(n7951), .A2(n6087), .ZN(n6088) );
  INV_X1 U5643 ( .A(n6948), .ZN(n6145) );
  NOR2_X1 U5644 ( .A1(n10181), .A2(n10032), .ZN(n10018) );
  OR2_X1 U5645 ( .A1(n6101), .A2(n10051), .ZN(n10032) );
  NAND2_X1 U5646 ( .A1(n10113), .A2(n5199), .ZN(n10051) );
  NOR2_X1 U5647 ( .A1(n10190), .A2(n5200), .ZN(n5199) );
  INV_X1 U5648 ( .A(n5201), .ZN(n5200) );
  NAND2_X1 U5649 ( .A1(n10113), .A2(n5203), .ZN(n10082) );
  NAND2_X1 U5650 ( .A1(n8253), .A2(n5193), .ZN(n8329) );
  NAND2_X1 U5651 ( .A1(n6065), .A2(n9923), .ZN(n6323) );
  AND2_X1 U5652 ( .A1(n7993), .A2(n8115), .ZN(n7995) );
  AND2_X1 U5653 ( .A1(n10551), .A2(n10593), .ZN(n7993) );
  NOR2_X1 U5654 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(P1_IR_REG_25__SCAN_IN), .ZN(
        n5587) );
  NOR2_X1 U5655 ( .A1(n6015), .A2(n5435), .ZN(n5434) );
  INV_X1 U5656 ( .A(n6012), .ZN(n5435) );
  AND2_X1 U5657 ( .A1(n5960), .A2(n5947), .ZN(n5959) );
  NAND2_X1 U5658 ( .A1(n5941), .A2(n5940), .ZN(n5399) );
  INV_X1 U5659 ( .A(SI_18_), .ZN(n8432) );
  INV_X1 U5660 ( .A(n5415), .ZN(n5414) );
  OAI21_X1 U5661 ( .B1(n5418), .B2(n5416), .A(n5862), .ZN(n5415) );
  NAND2_X1 U5662 ( .A1(n5417), .A2(n5848), .ZN(n5416) );
  INV_X1 U5663 ( .A(n5863), .ZN(n5417) );
  NAND2_X1 U5664 ( .A1(n5173), .A2(n5177), .ZN(n5172) );
  AOI21_X1 U5665 ( .B1(n5176), .B2(n5177), .A(n5175), .ZN(n5174) );
  NOR2_X1 U5666 ( .A1(n5826), .A2(SI_14_), .ZN(n5175) );
  INV_X1 U5667 ( .A(n5804), .ZN(n5176) );
  NAND2_X1 U5668 ( .A1(n5459), .A2(n5870), .ZN(n5458) );
  INV_X1 U5669 ( .A(n5574), .ZN(n5459) );
  NOR2_X1 U5670 ( .A1(n5773), .A2(n5429), .ZN(n5428) );
  INV_X1 U5671 ( .A(n5561), .ZN(n5429) );
  AND2_X1 U5672 ( .A1(n5115), .A2(n5554), .ZN(n5108) );
  INV_X1 U5673 ( .A(SI_9_), .ZN(n8549) );
  OAI211_X1 U5674 ( .C1(n5396), .C2(P2_DATAO_REG_3__SCAN_IN), .A(n5069), .B(
        n5068), .ZN(n5530) );
  NAND2_X1 U5675 ( .A1(n5170), .A2(n5070), .ZN(n5068) );
  INV_X1 U5676 ( .A(n5527), .ZN(n5156) );
  OR2_X1 U5677 ( .A1(n9112), .A2(n9245), .ZN(n5507) );
  OR2_X1 U5678 ( .A1(n8717), .A2(n8718), .ZN(n5497) );
  NOR2_X1 U5679 ( .A1(n8722), .A2(n5494), .ZN(n5493) );
  INV_X1 U5680 ( .A(n5497), .ZN(n5494) );
  NAND2_X1 U5681 ( .A1(n5496), .A2(n5498), .ZN(n5495) );
  OR2_X1 U5682 ( .A1(n6733), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n6741) );
  AND2_X1 U5683 ( .A1(n7505), .A2(n7552), .ZN(n7506) );
  OR2_X1 U5684 ( .A1(n7504), .A2(n7503), .ZN(n7505) );
  OAI21_X1 U5685 ( .B1(n7544), .B2(n7551), .A(n8926), .ZN(n7507) );
  XNOR2_X1 U5686 ( .A(n9110), .B(n5150), .ZN(n5149) );
  NAND2_X1 U5687 ( .A1(n9170), .A2(n4969), .ZN(n9218) );
  INV_X1 U5688 ( .A(n6759), .ZN(n6462) );
  OAI21_X1 U5689 ( .B1(n5480), .B2(n5132), .A(n5130), .ZN(n8347) );
  INV_X1 U5690 ( .A(n5131), .ZN(n5130) );
  OAI21_X1 U5691 ( .B1(n5481), .B2(n5132), .A(n8262), .ZN(n5131) );
  OR2_X1 U5692 ( .A1(n6707), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n6718) );
  NAND2_X1 U5693 ( .A1(n6459), .A2(n9237), .ZN(n6733) );
  INV_X1 U5694 ( .A(n6718), .ZN(n6459) );
  AND2_X1 U5695 ( .A1(n6847), .A2(n6515), .ZN(n7520) );
  INV_X1 U5696 ( .A(n9240), .ZN(n9261) );
  INV_X1 U5697 ( .A(n5489), .ZN(n5488) );
  OAI21_X1 U5698 ( .B1(n5492), .B2(n5491), .A(n9258), .ZN(n5489) );
  NOR2_X1 U5699 ( .A1(n8719), .A2(n4954), .ZN(n5492) );
  NAND2_X1 U5700 ( .A1(n6457), .A2(n8723), .ZN(n6681) );
  INV_X1 U5701 ( .A(n6670), .ZN(n6457) );
  OR2_X1 U5702 ( .A1(n6681), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n6694) );
  INV_X1 U5703 ( .A(n9056), .ZN(n9059) );
  OR2_X1 U5704 ( .A1(n7590), .A2(n7723), .ZN(n7592) );
  NAND2_X1 U5705 ( .A1(n7592), .A2(n7205), .ZN(n7563) );
  NAND2_X1 U5706 ( .A1(n7564), .A2(n7563), .ZN(n7562) );
  AND2_X1 U5707 ( .A1(n5097), .A2(n5096), .ZN(n10368) );
  NAND2_X1 U5708 ( .A1(n7206), .A2(n10360), .ZN(n5096) );
  AND2_X1 U5709 ( .A1(n7295), .A2(n10361), .ZN(n10386) );
  AOI21_X1 U5710 ( .B1(n10368), .B2(P2_REG1_REG_3__SCAN_IN), .A(n5095), .ZN(
        n10379) );
  INV_X1 U5711 ( .A(n5097), .ZN(n5095) );
  NAND2_X1 U5712 ( .A1(n10398), .A2(n7246), .ZN(n10425) );
  NAND2_X1 U5713 ( .A1(n10415), .A2(n7299), .ZN(n10435) );
  OR2_X1 U5714 ( .A1(n6545), .A2(P2_IR_REG_3__SCAN_IN), .ZN(n6586) );
  INV_X1 U5715 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n6584) );
  NAND2_X1 U5716 ( .A1(n10432), .A2(n7249), .ZN(n10449) );
  NAND2_X1 U5717 ( .A1(n10449), .A2(n10450), .ZN(n10448) );
  NAND2_X1 U5718 ( .A1(n5390), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n5389) );
  NAND2_X1 U5719 ( .A1(n7214), .A2(n5390), .ZN(n5388) );
  INV_X1 U5720 ( .A(n10457), .ZN(n5390) );
  NOR2_X1 U5721 ( .A1(n10441), .A2(n10440), .ZN(n10439) );
  XNOR2_X1 U5722 ( .A(n7251), .B(n10463), .ZN(n10465) );
  NAND2_X1 U5723 ( .A1(n10483), .A2(n7303), .ZN(n10501) );
  NAND2_X1 U5724 ( .A1(n10498), .A2(n7255), .ZN(n8629) );
  INV_X1 U5725 ( .A(n8627), .ZN(n5376) );
  NAND2_X1 U5726 ( .A1(n8632), .A2(n7305), .ZN(n9300) );
  NAND2_X1 U5727 ( .A1(n9296), .A2(n7258), .ZN(n9313) );
  NAND2_X1 U5728 ( .A1(n9313), .A2(n9314), .ZN(n9312) );
  INV_X1 U5729 ( .A(n9311), .ZN(n5382) );
  NAND2_X1 U5730 ( .A1(n9312), .A2(n5181), .ZN(n7260) );
  OR2_X1 U5731 ( .A1(n7277), .A2(n7259), .ZN(n5181) );
  NAND2_X1 U5732 ( .A1(n9346), .A2(n7262), .ZN(n7263) );
  NAND2_X1 U5733 ( .A1(n9350), .A2(n7309), .ZN(n9367) );
  AOI21_X1 U5734 ( .B1(P2_REG1_REG_16__SCAN_IN), .B2(n9356), .A(n9343), .ZN(
        n7227) );
  NAND2_X1 U5735 ( .A1(n6915), .A2(n6918), .ZN(n9116) );
  OAI21_X1 U5736 ( .B1(n9452), .B2(n5157), .A(n5325), .ZN(n5324) );
  AOI21_X1 U5737 ( .B1(n5326), .B2(n9043), .A(n9044), .ZN(n5325) );
  NAND2_X1 U5738 ( .A1(n5158), .A2(n5331), .ZN(n5157) );
  OR2_X1 U5739 ( .A1(n6769), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6779) );
  OR2_X1 U5740 ( .A1(n6779), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n6781) );
  AOI21_X1 U5741 ( .B1(n5272), .B2(n5275), .A(n5271), .ZN(n5270) );
  NAND2_X1 U5742 ( .A1(n5275), .A2(n5274), .ZN(n5273) );
  NOR2_X1 U5743 ( .A1(n9572), .A2(n9276), .ZN(n5271) );
  OR2_X1 U5744 ( .A1(n9452), .A2(n9453), .ZN(n5332) );
  NAND2_X1 U5745 ( .A1(n9505), .A2(n9504), .ZN(n9503) );
  INV_X1 U5746 ( .A(n5261), .ZN(n9513) );
  AOI21_X1 U5747 ( .B1(n5267), .B2(n5265), .A(n5264), .ZN(n5261) );
  AOI21_X1 U5748 ( .B1(n4955), .B2(n5316), .A(n8992), .ZN(n5313) );
  OR2_X1 U5749 ( .A1(n5233), .A2(n8987), .ZN(n5232) );
  NAND2_X1 U5750 ( .A1(n4974), .A2(n5236), .ZN(n5233) );
  OR2_X1 U5751 ( .A1(n6631), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6645) );
  OR2_X1 U5752 ( .A1(n8385), .A2(n8384), .ZN(n8976) );
  AND2_X1 U5753 ( .A1(n6860), .A2(n6859), .ZN(n5337) );
  NAND2_X1 U5754 ( .A1(n6452), .A2(n8573), .ZN(n6595) );
  INV_X1 U5755 ( .A(n6576), .ZN(n6452) );
  AND2_X1 U5756 ( .A1(n8954), .A2(n5244), .ZN(n5243) );
  AND2_X1 U5757 ( .A1(n6857), .A2(n8913), .ZN(n8886) );
  AND2_X1 U5758 ( .A1(n8938), .A2(n8943), .ZN(n5333) );
  AND2_X1 U5759 ( .A1(n8946), .A2(n8940), .ZN(n8879) );
  NAND2_X1 U5760 ( .A1(n5231), .A2(n7544), .ZN(n7718) );
  INV_X1 U5761 ( .A(n6850), .ZN(n7719) );
  INV_X1 U5762 ( .A(n8926), .ZN(n7717) );
  AND2_X1 U5763 ( .A1(n9070), .A2(n8090), .ZN(n6904) );
  AND4_X1 U5764 ( .A1(n6600), .A2(n6599), .A3(n6598), .A4(n6597), .ZN(n8192)
         );
  XNOR2_X1 U5765 ( .A(n6899), .B(n6478), .ZN(n7490) );
  AND2_X1 U5766 ( .A1(n5067), .A2(n6953), .ZN(n6958) );
  INV_X1 U5767 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n7803) );
  NAND2_X1 U5768 ( .A1(n9712), .A2(n7080), .ZN(n9719) );
  AND2_X1 U5769 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n5685) );
  NAND2_X1 U5770 ( .A1(n5067), .A2(n5066), .ZN(n7686) );
  AND2_X1 U5771 ( .A1(n6953), .A2(n6954), .ZN(n5066) );
  NAND2_X1 U5772 ( .A1(n7685), .A2(n7686), .ZN(n7684) );
  NAND2_X1 U5773 ( .A1(n8282), .A2(n5040), .ZN(n5034) );
  AOI21_X1 U5774 ( .B1(n4950), .B2(n5076), .A(n5011), .ZN(n5073) );
  INV_X1 U5775 ( .A(n7095), .ZN(n7096) );
  INV_X1 U5776 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n5702) );
  XNOR2_X1 U5777 ( .A(n7065), .B(n7166), .ZN(n8826) );
  NAND2_X1 U5778 ( .A1(n4971), .A2(n5407), .ZN(n6381) );
  INV_X1 U5779 ( .A(n6982), .ZN(n7838) );
  INV_X1 U5780 ( .A(n5624), .ZN(n5634) );
  AOI21_X1 U5781 ( .B1(n7631), .B2(P1_REG2_REG_8__SCAN_IN), .A(n7625), .ZN(
        n7535) );
  NOR2_X1 U5782 ( .A1(n9867), .A2(n9866), .ZN(n9870) );
  NOR2_X1 U5783 ( .A1(n9124), .A2(n5195), .ZN(n5194) );
  INV_X1 U5784 ( .A(n5196), .ZN(n5195) );
  AND2_X1 U5785 ( .A1(n7361), .A2(n5365), .ZN(n5364) );
  AND4_X1 U5786 ( .A1(n6059), .A2(n6058), .A3(n6057), .A4(n6056), .ZN(n9984)
         );
  AND2_X1 U5787 ( .A1(n6358), .A2(n6325), .ZN(n9993) );
  AOI21_X1 U5788 ( .B1(n5456), .B2(n10062), .A(n4990), .ZN(n5454) );
  NAND2_X1 U5789 ( .A1(n10079), .A2(n6426), .ZN(n10061) );
  AND4_X1 U5790 ( .A1(n5939), .A2(n5938), .A3(n5937), .A4(n5936), .ZN(n10097)
         );
  AND2_X1 U5791 ( .A1(n10117), .A2(n10112), .ZN(n10113) );
  NAND2_X1 U5792 ( .A1(n10113), .A2(n10262), .ZN(n10090) );
  NOR2_X1 U5793 ( .A1(n10147), .A2(n10222), .ZN(n10146) );
  INV_X1 U5794 ( .A(n5346), .ZN(n5345) );
  OAI21_X1 U5795 ( .B1(n5348), .B2(n5347), .A(n6297), .ZN(n5346) );
  NOR2_X1 U5796 ( .A1(n5855), .A2(n5854), .ZN(n5880) );
  INV_X1 U5797 ( .A(n5452), .ZN(n8786) );
  AND2_X1 U5798 ( .A1(n10230), .A2(n9801), .ZN(n5453) );
  NAND2_X1 U5799 ( .A1(n6097), .A2(n6096), .ZN(n8806) );
  NAND3_X1 U5800 ( .A1(n4976), .A2(n5821), .A3(n8253), .ZN(n8803) );
  AND2_X1 U5801 ( .A1(n5766), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n5780) );
  OR2_X1 U5802 ( .A1(n8074), .A2(n6398), .ZN(n6091) );
  AND2_X1 U5803 ( .A1(n8142), .A2(n5744), .ZN(n8253) );
  NAND2_X1 U5804 ( .A1(n5447), .A2(n5450), .ZN(n8180) );
  AOI21_X1 U5805 ( .B1(n5451), .B2(n8080), .A(n4993), .ZN(n5450) );
  INV_X1 U5806 ( .A(n5730), .ZN(n5451) );
  OR2_X1 U5807 ( .A1(n8034), .A2(n8038), .ZN(n8143) );
  NOR2_X1 U5808 ( .A1(n8143), .A2(n8271), .ZN(n8142) );
  AND4_X1 U5809 ( .A1(n5690), .A2(n5689), .A3(n5688), .A4(n5687), .ZN(n8030)
         );
  NOR2_X1 U5810 ( .A1(n10571), .A2(n10550), .ZN(n10551) );
  NAND2_X1 U5811 ( .A1(n6965), .A2(n7857), .ZN(n10550) );
  NAND2_X1 U5812 ( .A1(n6139), .A2(n10276), .ZN(n7161) );
  AND3_X1 U5813 ( .A1(n7159), .A2(n7178), .A3(n7158), .ZN(n6153) );
  NAND2_X1 U5814 ( .A1(n6141), .A2(n6126), .ZN(n10273) );
  AND2_X1 U5815 ( .A1(n6951), .A2(n7377), .ZN(n10274) );
  OAI21_X1 U5816 ( .B1(n6216), .B2(n6215), .A(n6206), .ZN(n6210) );
  XNOR2_X1 U5817 ( .A(n6195), .B(n6167), .ZN(n9666) );
  XNOR2_X1 U5818 ( .A(n6077), .B(n6076), .ZN(n9821) );
  NAND2_X1 U5819 ( .A1(n6116), .A2(n5581), .ZN(n6075) );
  INV_X1 U5820 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n6119) );
  INV_X1 U5821 ( .A(n5307), .ZN(n5306) );
  OAI21_X1 U5822 ( .B1(n5308), .B2(n5590), .A(n6064), .ZN(n5307) );
  AND2_X1 U5823 ( .A1(n5978), .A2(n5964), .ZN(n5965) );
  NAND2_X1 U5824 ( .A1(n6068), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6063) );
  AOI21_X1 U5825 ( .B1(n5831), .B2(n5412), .A(n5411), .ZN(n5893) );
  NOR2_X1 U5826 ( .A1(n5416), .A2(n5413), .ZN(n5412) );
  OAI21_X1 U5827 ( .B1(n5414), .B2(n5413), .A(n4994), .ZN(n5411) );
  INV_X1 U5828 ( .A(n5887), .ZN(n5413) );
  OR2_X1 U5829 ( .A1(n5833), .A2(P1_IR_REG_14__SCAN_IN), .ZN(n5834) );
  INV_X1 U5830 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n5571) );
  NAND2_X1 U5831 ( .A1(n5712), .A2(n5546), .ZN(n5723) );
  NAND2_X1 U5832 ( .A1(n5678), .A2(n5537), .ZN(n5692) );
  NAND2_X1 U5833 ( .A1(n5165), .A2(SI_1_), .ZN(n5164) );
  INV_X4 U5834 ( .A(n7427), .ZN(n7435) );
  NAND2_X1 U5835 ( .A1(n5485), .A2(n7874), .ZN(n8002) );
  INV_X1 U5836 ( .A(n7876), .ZN(n5485) );
  NAND2_X1 U5837 ( .A1(n5151), .A2(n5507), .ZN(n9156) );
  NAND2_X1 U5838 ( .A1(n5479), .A2(n5478), .ZN(n5151) );
  NAND2_X1 U5839 ( .A1(n5495), .A2(n5497), .ZN(n8721) );
  NAND2_X1 U5840 ( .A1(n7675), .A2(n7674), .ZN(n7676) );
  AOI21_X1 U5841 ( .B1(n5479), .B2(n5477), .A(n5474), .ZN(n9118) );
  AND2_X1 U5842 ( .A1(n9155), .A2(n5478), .ZN(n5477) );
  NAND2_X1 U5843 ( .A1(n5475), .A2(n5018), .ZN(n5474) );
  NAND2_X1 U5844 ( .A1(n8002), .A2(n8001), .ZN(n8125) );
  NAND2_X1 U5845 ( .A1(n6532), .A2(n7203), .ZN(n6506) );
  NAND2_X1 U5846 ( .A1(n9218), .A2(n9097), .ZN(n9178) );
  AOI21_X1 U5847 ( .B1(n8369), .B2(n8368), .A(n8367), .ZN(n8645) );
  AND2_X1 U5848 ( .A1(n8366), .A2(n8388), .ZN(n8367) );
  NAND2_X1 U5849 ( .A1(n9257), .A2(n9086), .ZN(n9193) );
  AOI21_X1 U5850 ( .B1(n5486), .B2(n4973), .A(n5144), .ZN(n9203) );
  AOI22_X1 U5851 ( .A1(n9162), .A2(n9459), .B1(n9106), .B2(n9105), .ZN(n9210)
         );
  INV_X1 U5852 ( .A(n7710), .ZN(n5473) );
  NAND2_X1 U5853 ( .A1(n5480), .A2(n5481), .ZN(n8127) );
  NAND2_X1 U5854 ( .A1(n8127), .A2(n8126), .ZN(n8263) );
  NAND2_X1 U5855 ( .A1(n9170), .A2(n9094), .ZN(n9220) );
  NAND2_X1 U5856 ( .A1(n5136), .A2(n5134), .ZN(n9227) );
  AOI21_X1 U5857 ( .B1(n5137), .B2(n5138), .A(n5135), .ZN(n5134) );
  INV_X1 U5858 ( .A(n9228), .ZN(n5135) );
  NAND2_X1 U5859 ( .A1(n5133), .A2(n5137), .ZN(n9229) );
  OR2_X1 U5860 ( .A1(n9170), .A2(n5138), .ZN(n5133) );
  NAND2_X1 U5861 ( .A1(n5143), .A2(n5142), .ZN(n9236) );
  OAI21_X1 U5862 ( .B1(n5144), .B2(n4977), .A(n4953), .ZN(n5142) );
  NAND2_X1 U5863 ( .A1(n7765), .A2(n7764), .ZN(n7873) );
  NAND2_X1 U5864 ( .A1(n7516), .A2(n10677), .ZN(n9251) );
  NAND2_X1 U5865 ( .A1(n6792), .A2(n6791), .ZN(n9252) );
  INV_X1 U5866 ( .A(n9238), .ZN(n9263) );
  NAND2_X1 U5867 ( .A1(n5486), .A2(n5488), .ZN(n9257) );
  NAND2_X1 U5868 ( .A1(n5487), .A2(n5490), .ZN(n9259) );
  NAND2_X1 U5869 ( .A1(n5496), .A2(n5492), .ZN(n5487) );
  INV_X1 U5870 ( .A(n9254), .ZN(n9256) );
  NAND2_X1 U5871 ( .A1(n9072), .A2(n9073), .ZN(n5214) );
  AND2_X1 U5872 ( .A1(n9070), .A2(n8090), .ZN(n5207) );
  INV_X1 U5873 ( .A(n5210), .ZN(n5209) );
  OAI21_X1 U5874 ( .B1(n5211), .B2(n9080), .A(n9079), .ZN(n5210) );
  NAND2_X1 U5875 ( .A1(n6492), .A2(n6491), .ZN(n9275) );
  AND2_X1 U5876 ( .A1(n6528), .A2(n6529), .ZN(n5339) );
  INV_X2 U5877 ( .A(P2_U3893), .ZN(n9292) );
  INV_X1 U5878 ( .A(n5231), .ZN(n5513) );
  NAND3_X1 U5879 ( .A1(n5089), .A2(n5088), .A3(n5087), .ZN(n7203) );
  NAND3_X1 U5880 ( .A1(n5187), .A2(P2_IR_REG_31__SCAN_IN), .A3(
        P2_IR_REG_0__SCAN_IN), .ZN(n5088) );
  NAND2_X1 U5881 ( .A1(n6609), .A2(P2_IR_REG_1__SCAN_IN), .ZN(n5089) );
  NAND2_X1 U5882 ( .A1(n7236), .A2(P2_IR_REG_1__SCAN_IN), .ZN(n5087) );
  NAND3_X1 U5883 ( .A1(n5185), .A2(n5184), .A3(n5183), .ZN(n7582) );
  OAI211_X1 U5884 ( .C1(P2_IR_REG_0__SCAN_IN), .C2(P2_IR_REG_1__SCAN_IN), .A(
        n5186), .B(P2_IR_REG_31__SCAN_IN), .ZN(n5183) );
  NAND2_X1 U5885 ( .A1(n6609), .A2(P2_IR_REG_2__SCAN_IN), .ZN(n5185) );
  NOR2_X1 U5886 ( .A1(n5029), .A2(n7211), .ZN(n10421) );
  INV_X1 U5887 ( .A(n5386), .ZN(n10471) );
  INV_X1 U5888 ( .A(n7217), .ZN(n5385) );
  INV_X1 U5889 ( .A(n5375), .ZN(n10507) );
  OR2_X1 U5890 ( .A1(n10509), .A2(n10508), .ZN(n5375) );
  INV_X1 U5891 ( .A(n7220), .ZN(n5374) );
  NAND2_X1 U5892 ( .A1(n5371), .A2(n5372), .ZN(n8626) );
  NAND2_X1 U5893 ( .A1(n7220), .A2(n5376), .ZN(n5372) );
  OR2_X1 U5894 ( .A1(n10509), .A2(n5373), .ZN(n5371) );
  NAND2_X1 U5895 ( .A1(n5376), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n5373) );
  INV_X1 U5896 ( .A(n7223), .ZN(n5380) );
  XNOR2_X1 U5897 ( .A(n7260), .B(n7275), .ZN(n9331) );
  NOR2_X1 U5898 ( .A1(n9327), .A2(n7225), .ZN(n9345) );
  NOR2_X1 U5899 ( .A1(n9310), .A2(n5021), .ZN(n7224) );
  XNOR2_X1 U5900 ( .A(n7263), .B(n7272), .ZN(n9365) );
  NAND2_X1 U5901 ( .A1(n9365), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n9364) );
  XNOR2_X1 U5902 ( .A(n7227), .B(n7272), .ZN(n9362) );
  NOR2_X1 U5903 ( .A1(n9362), .A2(n9363), .ZN(n9361) );
  OAI21_X1 U5904 ( .B1(n9362), .B2(n5392), .A(n5391), .ZN(n9378) );
  NAND2_X1 U5905 ( .A1(n5393), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n5392) );
  NAND2_X1 U5906 ( .A1(n7228), .A2(n5393), .ZN(n5391) );
  INV_X1 U5907 ( .A(n9379), .ZN(n5393) );
  INV_X1 U5908 ( .A(n7270), .ZN(n5189) );
  NAND2_X1 U5909 ( .A1(n6818), .A2(n6817), .ZN(n9145) );
  AND2_X1 U5910 ( .A1(n6827), .A2(n6826), .ZN(n9408) );
  NAND2_X1 U5911 ( .A1(n6804), .A2(n6803), .ZN(n9555) );
  NAND2_X1 U5912 ( .A1(n6802), .A2(n6801), .ZN(n9563) );
  INV_X1 U5913 ( .A(n5331), .ZN(n5330) );
  NAND2_X1 U5914 ( .A1(n5269), .A2(n5275), .ZN(n9445) );
  NAND2_X1 U5915 ( .A1(n9482), .A2(n5277), .ZN(n5269) );
  OAI21_X1 U5916 ( .B1(n9482), .B2(n9478), .A(n5280), .ZN(n9457) );
  OAI21_X1 U5917 ( .B1(n9505), .B2(n5321), .A(n5319), .ZN(n9477) );
  AND2_X1 U5918 ( .A1(n9482), .A2(n6747), .ZN(n9467) );
  NAND2_X1 U5919 ( .A1(n9541), .A2(n6867), .ZN(n9526) );
  NAND2_X1 U5920 ( .A1(n6717), .A2(n6716), .ZN(n9524) );
  NAND2_X1 U5921 ( .A1(n6693), .A2(n6692), .ZN(n9611) );
  NAND2_X1 U5922 ( .A1(n5314), .A2(n6866), .ZN(n8746) );
  NAND2_X1 U5923 ( .A1(n8672), .A2(n8987), .ZN(n5314) );
  NAND2_X1 U5924 ( .A1(n6680), .A2(n6679), .ZN(n9083) );
  NAND2_X1 U5925 ( .A1(n5235), .A2(n6663), .ZN(n8674) );
  NAND2_X1 U5926 ( .A1(n8696), .A2(n8974), .ZN(n5235) );
  AND4_X1 U5927 ( .A1(n6650), .A2(n6649), .A3(n6648), .A4(n6647), .ZN(n8698)
         );
  INV_X1 U5928 ( .A(n9282), .ZN(n8388) );
  NAND2_X1 U5929 ( .A1(n5338), .A2(n6859), .ZN(n8217) );
  OAI21_X1 U5930 ( .B1(n7959), .B2(n5246), .A(n5245), .ZN(n8060) );
  INV_X1 U5931 ( .A(n9509), .ZN(n10636) );
  AND2_X1 U5932 ( .A1(n9060), .A2(n6904), .ZN(n9150) );
  NAND2_X1 U5933 ( .A1(n7514), .A2(n10679), .ZN(n10677) );
  INV_X1 U5934 ( .A(n9252), .ZN(n9638) );
  INV_X1 U5935 ( .A(n9215), .ZN(n9643) );
  OR3_X1 U5936 ( .A1(n9607), .A2(n9606), .A3(n9605), .ZN(n9657) );
  NAND2_X1 U5937 ( .A1(n7454), .A2(n8849), .ZN(n5219) );
  AND2_X1 U5938 ( .A1(n7491), .A2(n7468), .ZN(n9659) );
  AND2_X1 U5939 ( .A1(n7490), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7468) );
  INV_X1 U5940 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n6479) );
  XNOR2_X1 U5941 ( .A(n6880), .B(n6879), .ZN(n8799) );
  INV_X1 U5942 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n6879) );
  INV_X1 U5943 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n6875) );
  NAND2_X1 U5944 ( .A1(n6874), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6876) );
  OR2_X1 U5945 ( .A1(n6878), .A2(n6872), .ZN(n6873) );
  AND2_X1 U5946 ( .A1(n7435), .A2(P2_U3151), .ZN(n9674) );
  INV_X1 U5947 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n6832) );
  XNOR2_X1 U5948 ( .A(n6835), .B(n6834), .ZN(n9070) );
  INV_X1 U5949 ( .A(n7273), .ZN(n9356) );
  INV_X1 U5950 ( .A(n10479), .ZN(n7463) );
  INV_X1 U5951 ( .A(n7290), .ZN(n10404) );
  NAND2_X1 U5952 ( .A1(n8048), .A2(n7002), .ZN(n5055) );
  OAI21_X1 U5953 ( .B1(n9780), .B2(n7324), .A(n7325), .ZN(n7326) );
  AOI21_X1 U5954 ( .B1(n10230), .B2(n7140), .A(n7059), .ZN(n8817) );
  NOR3_X1 U5955 ( .A1(n9780), .A2(n7324), .A3(n7325), .ZN(n7328) );
  AND4_X1 U5956 ( .A1(n5785), .A2(n5784), .A3(n5783), .A4(n5782), .ZN(n8706)
         );
  NAND2_X1 U5957 ( .A1(n6020), .A2(n6019), .ZN(n10174) );
  OR2_X1 U5958 ( .A1(n8785), .A2(n6018), .ZN(n6020) );
  NAND2_X1 U5959 ( .A1(n5298), .A2(n4970), .ZN(n9704) );
  NAND2_X1 U5960 ( .A1(n7835), .A2(n6994), .ZN(n7924) );
  OAI211_X1 U5961 ( .C1(n6018), .C2(n7447), .A(n5701), .B(n5700), .ZN(n7928)
         );
  NAND2_X1 U5962 ( .A1(n5879), .A2(n5878), .ZN(n10131) );
  INV_X1 U5963 ( .A(n10047), .ZN(n9753) );
  OAI21_X1 U5964 ( .B1(n9678), .B2(n9679), .A(n5303), .ZN(n9730) );
  NAND2_X1 U5965 ( .A1(n8700), .A2(n7051), .ZN(n8735) );
  AND4_X1 U5966 ( .A1(n5957), .A2(n5956), .A3(n5955), .A4(n5954), .ZN(n10081)
         );
  NAND2_X1 U5967 ( .A1(n8338), .A2(n5290), .ZN(n5285) );
  INV_X1 U5968 ( .A(n9787), .ZN(n9775) );
  NAND2_X1 U5969 ( .A1(n5905), .A2(n5904), .ZN(n10210) );
  AND2_X1 U5970 ( .A1(n6054), .A2(n6039), .ZN(n9977) );
  AND2_X1 U5971 ( .A1(n7688), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9788) );
  AND2_X1 U5972 ( .A1(n7182), .A2(n10287), .ZN(n9786) );
  INV_X1 U5973 ( .A(n9780), .ZN(n9785) );
  INV_X1 U5974 ( .A(n9786), .ZN(n9754) );
  NAND2_X1 U5975 ( .A1(n7180), .A2(n10606), .ZN(n9789) );
  INV_X1 U5976 ( .A(n6065), .ZN(n6447) );
  INV_X1 U5977 ( .A(n9996), .ZN(n9797) );
  NOR2_X1 U5978 ( .A1(n5925), .A2(n5924), .ZN(n10111) );
  INV_X1 U5979 ( .A(n8029), .ZN(n9806) );
  INV_X1 U5980 ( .A(n8136), .ZN(n9807) );
  INV_X1 U5981 ( .A(n8030), .ZN(n9808) );
  INV_X1 U5982 ( .A(P1_U3973), .ZN(n9825) );
  NAND2_X1 U5983 ( .A1(n5796), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5628) );
  AOI21_X1 U5984 ( .B1(n10527), .B2(P1_REG2_REG_4__SCAN_IN), .A(n10522), .ZN(
        n7638) );
  AOI21_X1 U5985 ( .B1(P1_REG2_REG_6__SCAN_IN), .B2(n7619), .A(n7613), .ZN(
        n7602) );
  AOI21_X1 U5986 ( .B1(n7662), .B2(P1_REG2_REG_10__SCAN_IN), .A(n7656), .ZN(
        n7748) );
  AOI21_X1 U5987 ( .B1(P1_REG2_REG_13__SCAN_IN), .B2(n8108), .A(n8102), .ZN(
        n8224) );
  AOI21_X1 U5988 ( .B1(P1_REG2_REG_16__SCAN_IN), .B2(n9881), .A(n9876), .ZN(
        n9877) );
  NOR2_X1 U5989 ( .A1(n7478), .A2(n7474), .ZN(n10524) );
  AND2_X1 U5990 ( .A1(n7355), .A2(n9944), .ZN(n9955) );
  INV_X1 U5991 ( .A(n5444), .ZN(n7354) );
  AND2_X1 U5992 ( .A1(n6107), .A2(n6055), .ZN(n9966) );
  NOR2_X1 U5993 ( .A1(n9979), .A2(n6324), .ZN(n6104) );
  NAND2_X1 U5994 ( .A1(n10026), .A2(n5121), .ZN(n10012) );
  NAND2_X1 U5995 ( .A1(n10044), .A2(n6230), .ZN(n10028) );
  NAND2_X1 U5996 ( .A1(n5457), .A2(n5456), .ZN(n10040) );
  AND2_X1 U5997 ( .A1(n5457), .A2(n4966), .ZN(n10042) );
  AOI21_X1 U5998 ( .B1(n10138), .B2(n4952), .A(n5465), .ZN(n10098) );
  NAND2_X1 U5999 ( .A1(n5464), .A2(n5466), .ZN(n10107) );
  NAND2_X1 U6000 ( .A1(n10138), .A2(n5467), .ZN(n5464) );
  AOI21_X1 U6001 ( .B1(n10138), .B2(n10137), .A(n5469), .ZN(n10120) );
  NAND2_X1 U6002 ( .A1(n5344), .A2(n5348), .ZN(n10140) );
  OR2_X1 U6003 ( .A1(n8808), .A2(n5351), .ZN(n5344) );
  NAND2_X1 U6004 ( .A1(n8660), .A2(n5361), .ZN(n8685) );
  NOR2_X1 U6005 ( .A1(n5360), .A2(n5359), .ZN(n8686) );
  INV_X1 U6006 ( .A(n10235), .ZN(n5821) );
  NAND2_X1 U6007 ( .A1(n8081), .A2(n8080), .ZN(n8079) );
  NAND2_X1 U6008 ( .A1(n8134), .A2(n5730), .ZN(n8081) );
  NAND2_X1 U6009 ( .A1(n10573), .A2(n7980), .ZN(n10615) );
  INV_X1 U6010 ( .A(n10606), .ZN(n10572) );
  INV_X1 U6011 ( .A(n10612), .ZN(n10570) );
  AND2_X1 U6012 ( .A1(n10576), .A2(n10552), .ZN(n10002) );
  AND2_X1 U6013 ( .A1(n9930), .A2(n10155), .ZN(n9131) );
  AND2_X1 U6014 ( .A1(n9954), .A2(n10165), .ZN(n10166) );
  AND2_X1 U6015 ( .A1(n10164), .A2(n5512), .ZN(n10165) );
  NAND2_X1 U6016 ( .A1(n6035), .A2(n6034), .ZN(n10249) );
  INV_X1 U6017 ( .A(n10131), .ZN(n10268) );
  INV_X1 U6018 ( .A(n7928), .ZN(n10613) );
  INV_X1 U6019 ( .A(n9821), .ZN(n10287) );
  INV_X1 U6020 ( .A(n6072), .ZN(n8320) );
  NAND2_X1 U6021 ( .A1(n5914), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5033) );
  NAND2_X1 U6022 ( .A1(n5424), .A2(n5422), .ZN(n5789) );
  NAND2_X1 U6023 ( .A1(n5424), .A2(n5425), .ZN(n5788) );
  NAND2_X1 U6024 ( .A1(n5111), .A2(n5116), .ZN(n5110) );
  NAND2_X1 U6025 ( .A1(n5659), .A2(n5533), .ZN(n5676) );
  INV_X1 U6026 ( .A(n5381), .ZN(n9293) );
  XNOR2_X1 U6027 ( .A(n7268), .B(n5189), .ZN(n5188) );
  OAI21_X1 U6028 ( .B1(n8839), .B2(n9509), .A(n6943), .ZN(n6944) );
  NOR2_X1 U6029 ( .A1(n6907), .A2(n6909), .ZN(n6910) );
  INV_X1 U6030 ( .A(n7377), .ZN(n7378) );
  NAND2_X1 U6031 ( .A1(n7810), .A2(n5059), .ZN(n7817) );
  AND2_X1 U6032 ( .A1(n7376), .A2(n7375), .ZN(n5504) );
  NAND2_X1 U6033 ( .A1(n5511), .A2(n5508), .ZN(n7371) );
  NAND2_X1 U6034 ( .A1(n6154), .A2(n10674), .ZN(n5124) );
  NAND2_X1 U6035 ( .A1(n10671), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n5123) );
  NAND2_X1 U6036 ( .A1(n5795), .A2(n5794), .ZN(n8665) );
  NAND2_X1 U6037 ( .A1(n9098), .A2(n9488), .ZN(n4947) );
  OR2_X1 U6038 ( .A1(n5747), .A2(n5458), .ZN(n4949) );
  INV_X1 U6039 ( .A(n5401), .ZN(n6435) );
  AND2_X1 U6040 ( .A1(n9722), .A2(n5074), .ZN(n4950) );
  OR2_X1 U6041 ( .A1(n9145), .A2(n9554), .ZN(n4951) );
  AND2_X1 U6042 ( .A1(n7153), .A2(n7152), .ZN(n7324) );
  AND2_X1 U6043 ( .A1(n10106), .A2(n5467), .ZN(n4952) );
  NAND2_X1 U6044 ( .A1(n9089), .A2(n9516), .ZN(n4953) );
  AND2_X1 U6045 ( .A1(n5479), .A2(n5014), .ZN(n9244) );
  AND2_X1 U6046 ( .A1(n9082), .A2(n9081), .ZN(n4954) );
  AND2_X1 U6047 ( .A1(n5315), .A2(n8894), .ZN(n4955) );
  OAI211_X2 U6048 ( .C1(n6756), .C2(n7437), .A(n6507), .B(n6506), .ZN(n7523)
         );
  INV_X1 U6049 ( .A(n10650), .ZN(n5032) );
  AND2_X1 U6050 ( .A1(n9739), .A2(n5065), .ZN(n4956) );
  AND2_X1 U6051 ( .A1(n9003), .A2(n6867), .ZN(n4957) );
  AND2_X1 U6052 ( .A1(n9638), .A2(n9245), .ZN(n4958) );
  NAND2_X1 U6053 ( .A1(n6758), .A2(n6757), .ZN(n9099) );
  INV_X1 U6054 ( .A(n9099), .ZN(n9648) );
  OR2_X1 U6055 ( .A1(n5300), .A2(n5299), .ZN(n4959) );
  AND2_X1 U6056 ( .A1(n5002), .A2(n5441), .ZN(n4961) );
  NOR2_X1 U6057 ( .A1(n10262), .A2(n10111), .ZN(n4962) );
  AND2_X1 U6058 ( .A1(n5193), .A2(n5192), .ZN(n4963) );
  INV_X1 U6059 ( .A(n7329), .ZN(n9969) );
  NAND2_X1 U6060 ( .A1(n6051), .A2(n6050), .ZN(n7329) );
  AOI21_X1 U6061 ( .B1(n9795), .B2(n10557), .A(n9940), .ZN(n9941) );
  INV_X1 U6062 ( .A(n7275), .ZN(n5104) );
  NAND2_X1 U6063 ( .A1(n4976), .A2(n8253), .ZN(n4964) );
  INV_X1 U6064 ( .A(n8719), .ZN(n5498) );
  INV_X1 U6065 ( .A(n6227), .ZN(n5408) );
  NAND3_X2 U6066 ( .A1(n6951), .A2(n7854), .A3(n6949), .ZN(n6963) );
  INV_X1 U6067 ( .A(n5796), .ZN(n5920) );
  NAND2_X1 U6068 ( .A1(n9572), .A2(n9459), .ZN(n4965) );
  AND2_X4 U6069 ( .A1(n5618), .A2(n7427), .ZN(n5660) );
  INV_X1 U6070 ( .A(n7551), .ZN(n9110) );
  NAND2_X1 U6071 ( .A1(n7502), .A2(n7501), .ZN(n7551) );
  INV_X1 U6072 ( .A(n5745), .ZN(n5111) );
  OR2_X1 U6073 ( .A1(n9099), .A2(n9580), .ZN(n8874) );
  INV_X1 U6074 ( .A(n7846), .ZN(n5150) );
  NAND2_X1 U6075 ( .A1(n5981), .A2(n5980), .ZN(n6101) );
  NAND2_X1 U6076 ( .A1(n10070), .A2(n10048), .ZN(n4966) );
  AND2_X1 U6077 ( .A1(n5560), .A2(n5116), .ZN(n5115) );
  AND2_X1 U6078 ( .A1(n9602), .A2(n9608), .ZN(n4967) );
  INV_X1 U6079 ( .A(n5258), .ZN(n5257) );
  INV_X1 U6080 ( .A(n5830), .ZN(n5418) );
  AND2_X1 U6081 ( .A1(n7236), .A2(n5187), .ZN(n4968) );
  AND2_X1 U6082 ( .A1(n9095), .A2(n9094), .ZN(n4969) );
  NOR2_X1 U6083 ( .A1(n5493), .A2(n4954), .ZN(n5491) );
  OR2_X1 U6084 ( .A1(n5301), .A2(n5300), .ZN(n4970) );
  AND4_X1 U6085 ( .A1(n9945), .A2(n7356), .A3(n6194), .A4(n6193), .ZN(n4971)
         );
  NAND2_X1 U6086 ( .A1(n5917), .A2(n5916), .ZN(n10102) );
  OR3_X1 U6087 ( .A1(P2_IR_REG_25__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), .A3(
        P2_IR_REG_26__SCAN_IN), .ZN(n4972) );
  AND2_X1 U6088 ( .A1(n5488), .A2(n9192), .ZN(n4973) );
  NAND2_X1 U6089 ( .A1(n9687), .A2(n7104), .ZN(n9738) );
  OAI21_X1 U6090 ( .B1(n9452), .B2(n5330), .A(n5328), .ZN(n9425) );
  INV_X1 U6091 ( .A(n8137), .ZN(n5449) );
  OR2_X1 U6092 ( .A1(n8974), .A2(n5236), .ZN(n4974) );
  NOR2_X1 U6093 ( .A1(n6853), .A2(n5150), .ZN(n4975) );
  AND2_X1 U6094 ( .A1(n4963), .A2(n10662), .ZN(n4976) );
  INV_X1 U6095 ( .A(n10376), .ZN(n7429) );
  XNOR2_X1 U6096 ( .A(n6556), .B(P2_IR_REG_4__SCAN_IN), .ZN(n10376) );
  AND2_X1 U6097 ( .A1(n9201), .A2(n9608), .ZN(n4977) );
  OR2_X1 U6098 ( .A1(n6076), .A2(n5440), .ZN(n4978) );
  NAND2_X1 U6099 ( .A1(n6727), .A2(n6477), .ZN(n6836) );
  INV_X1 U6100 ( .A(n6288), .ZN(n5349) );
  NAND2_X1 U6101 ( .A1(n5573), .A2(n5572), .ZN(n5747) );
  NAND2_X1 U6102 ( .A1(n5084), .A2(n5570), .ZN(n5695) );
  NAND2_X1 U6103 ( .A1(n7527), .A2(n6508), .ZN(n8921) );
  AND4_X1 U6104 ( .A1(n5756), .A2(n5755), .A3(n5754), .A4(n5753), .ZN(n8246)
         );
  NAND2_X1 U6105 ( .A1(n10044), .A2(n5354), .ZN(n10026) );
  NOR2_X1 U6106 ( .A1(n8359), .A2(n9283), .ZN(n4979) );
  INV_X1 U6107 ( .A(n9092), .ZN(n9504) );
  NOR2_X1 U6108 ( .A1(n7129), .A2(n7128), .ZN(n4980) );
  AND2_X1 U6109 ( .A1(n5298), .A2(n5295), .ZN(n4981) );
  AND4_X1 U6110 ( .A1(n5771), .A2(n5770), .A3(n5769), .A4(n5768), .ZN(n8290)
         );
  INV_X1 U6111 ( .A(n8290), .ZN(n9805) );
  NOR2_X1 U6112 ( .A1(n9361), .A2(n7228), .ZN(n4982) );
  NAND2_X1 U6113 ( .A1(n5969), .A2(n5968), .ZN(n10190) );
  AND2_X1 U6114 ( .A1(n7111), .A2(n7110), .ZN(n4983) );
  AND2_X1 U6115 ( .A1(n6362), .A2(n9935), .ZN(n7356) );
  OR2_X1 U6116 ( .A1(n6337), .A2(n6339), .ZN(n4984) );
  INV_X1 U6117 ( .A(n9097), .ZN(n5140) );
  NOR2_X1 U6118 ( .A1(n5827), .A2(n5178), .ZN(n5177) );
  INV_X1 U6119 ( .A(n9980), .ZN(n5366) );
  NAND2_X1 U6120 ( .A1(n6359), .A2(n6326), .ZN(n9980) );
  NAND2_X1 U6121 ( .A1(n9088), .A2(n9535), .ZN(n4985) );
  AND2_X1 U6122 ( .A1(n5551), .A2(n5550), .ZN(n4986) );
  INV_X1 U6123 ( .A(n9124), .ZN(n10245) );
  NAND2_X1 U6124 ( .A1(n6219), .A2(n6218), .ZN(n9124) );
  NAND2_X1 U6125 ( .A1(n8189), .A2(n6620), .ZN(n4987) );
  OR2_X1 U6126 ( .A1(n9431), .A2(n9438), .ZN(n4988) );
  INV_X1 U6127 ( .A(n5355), .ZN(n5354) );
  NAND2_X1 U6128 ( .A1(n6102), .A2(n6230), .ZN(n5355) );
  NOR2_X1 U6129 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), .ZN(
        n5586) );
  AND3_X1 U6130 ( .A1(n5622), .A2(n5621), .A3(n5620), .ZN(n6965) );
  INV_X1 U6131 ( .A(n6965), .ZN(n7861) );
  NAND2_X1 U6132 ( .A1(n9124), .A2(n9939), .ZN(n4989) );
  AND2_X1 U6133 ( .A1(n7358), .A2(n6344), .ZN(n6194) );
  INV_X1 U6134 ( .A(n6194), .ZN(n5370) );
  INV_X1 U6135 ( .A(n8176), .ZN(n8286) );
  AND4_X1 U6136 ( .A1(n5743), .A2(n5742), .A3(n5741), .A4(n5740), .ZN(n8176)
         );
  INV_X1 U6137 ( .A(n7026), .ZN(n5043) );
  NAND2_X1 U6138 ( .A1(n5063), .A2(n5062), .ZN(n9694) );
  AND2_X1 U6139 ( .A1(n5977), .A2(n10065), .ZN(n4990) );
  NOR2_X1 U6140 ( .A1(n9581), .A2(n9488), .ZN(n4991) );
  INV_X1 U6141 ( .A(n5296), .ZN(n5295) );
  NAND2_X1 U6142 ( .A1(n4970), .A2(n5297), .ZN(n5296) );
  NAND3_X1 U6143 ( .A1(n10516), .A2(P2_ADDR_REG_19__SCAN_IN), .A3(
        P1_ADDR_REG_19__SCAN_IN), .ZN(n5395) );
  INV_X1 U6144 ( .A(n5395), .ZN(n5170) );
  INV_X1 U6145 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n5870) );
  OR2_X1 U6146 ( .A1(n9045), .A2(n9419), .ZN(n4992) );
  AND2_X1 U6147 ( .A1(n8176), .A2(n5744), .ZN(n4993) );
  OR2_X1 U6148 ( .A1(n5886), .A2(SI_17_), .ZN(n4994) );
  AND2_X1 U6149 ( .A1(n5112), .A2(n5110), .ZN(n4995) );
  NAND2_X1 U6150 ( .A1(n10210), .A2(n9799), .ZN(n4996) );
  INV_X1 U6151 ( .A(n7149), .ZN(n5294) );
  OR2_X1 U6152 ( .A1(n7154), .A2(n6971), .ZN(n4997) );
  INV_X1 U6153 ( .A(n5368), .ZN(n9979) );
  NAND2_X1 U6154 ( .A1(n5367), .A2(n5366), .ZN(n5368) );
  INV_X1 U6155 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n5572) );
  NAND2_X1 U6156 ( .A1(n9252), .A2(n9563), .ZN(n4998) );
  AND2_X1 U6157 ( .A1(n6262), .A2(n8071), .ZN(n4999) );
  NAND2_X1 U6158 ( .A1(n8702), .A2(n8767), .ZN(n5000) );
  INV_X1 U6159 ( .A(n5679), .ZN(n5084) );
  OR2_X1 U6160 ( .A1(n9215), .A2(n9165), .ZN(n8872) );
  NOR2_X1 U6161 ( .A1(n10268), .A2(n10144), .ZN(n5001) );
  OAI21_X1 U6162 ( .B1(n4969), .B2(n5140), .A(n9179), .ZN(n5139) );
  OR2_X1 U6163 ( .A1(n7352), .A2(n7351), .ZN(n5002) );
  INV_X1 U6164 ( .A(n9003), .ZN(n9525) );
  AND2_X1 U6165 ( .A1(n9007), .A2(n9009), .ZN(n9003) );
  INV_X1 U6166 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n6609) );
  INV_X1 U6167 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n5070) );
  INV_X1 U6168 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n5187) );
  NAND2_X1 U6169 ( .A1(n9083), .A2(n9617), .ZN(n8989) );
  OR2_X1 U6170 ( .A1(n9564), .A2(n9438), .ZN(n9043) );
  INV_X1 U6171 ( .A(n9043), .ZN(n5327) );
  AND2_X1 U6172 ( .A1(n6367), .A2(n6432), .ZN(n9945) );
  AND2_X1 U6173 ( .A1(n5332), .A2(n4965), .ZN(n5003) );
  AND2_X1 U6174 ( .A1(n5581), .A2(n5586), .ZN(n5004) );
  AND2_X1 U6175 ( .A1(n5874), .A2(n5085), .ZN(n5005) );
  INV_X1 U6176 ( .A(n5554), .ZN(n5114) );
  NOR2_X1 U6177 ( .A1(n6324), .A2(n5370), .ZN(n5369) );
  OR2_X1 U6178 ( .A1(n10420), .A2(n10402), .ZN(n5006) );
  AND2_X1 U6179 ( .A1(n5180), .A2(n5248), .ZN(n5007) );
  NOR2_X1 U6180 ( .A1(n8124), .A2(n5484), .ZN(n5483) );
  AND2_X1 U6181 ( .A1(n5252), .A2(n5007), .ZN(n5008) );
  AND2_X1 U6182 ( .A1(n5336), .A2(n5335), .ZN(n5009) );
  INV_X1 U6183 ( .A(n5491), .ZN(n5490) );
  INV_X1 U6184 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5085) );
  NOR2_X1 U6185 ( .A1(n5747), .A2(n5574), .ZN(n5010) );
  AND2_X1 U6186 ( .A1(n6422), .A2(n6423), .ZN(n6306) );
  INV_X1 U6187 ( .A(n6306), .ZN(n5463) );
  XNOR2_X1 U6188 ( .A(n6063), .B(P1_IR_REG_21__SCAN_IN), .ZN(n6072) );
  NAND2_X1 U6189 ( .A1(n5034), .A2(n5037), .ZN(n8701) );
  INV_X1 U6190 ( .A(n10447), .ZN(n7457) );
  NAND2_X1 U6191 ( .A1(n5824), .A2(n5823), .ZN(n8801) );
  NAND2_X1 U6192 ( .A1(n5031), .A2(n8816), .ZN(n8825) );
  NAND2_X1 U6193 ( .A1(n5267), .A2(n6700), .ZN(n9530) );
  XOR2_X1 U6194 ( .A(n7092), .B(n7166), .Z(n5011) );
  INV_X1 U6195 ( .A(n6413), .ZN(n5347) );
  OR2_X1 U6196 ( .A1(n7137), .A2(n7136), .ZN(n5012) );
  AND2_X2 U6197 ( .A1(n8866), .A2(n9078), .ZN(n9060) );
  AND2_X1 U6198 ( .A1(n7129), .A2(n7128), .ZN(n5013) );
  NAND2_X1 U6199 ( .A1(n5285), .A2(n5289), .ZN(n8764) );
  NAND2_X1 U6200 ( .A1(n5311), .A2(n9770), .ZN(n9686) );
  NAND2_X1 U6201 ( .A1(n9109), .A2(n9438), .ZN(n5014) );
  NAND2_X1 U6202 ( .A1(n7060), .A2(n7061), .ZN(n8815) );
  NAND2_X1 U6203 ( .A1(n6766), .A2(n6765), .ZN(n9580) );
  AND2_X1 U6204 ( .A1(n9719), .A2(n9720), .ZN(n5015) );
  NAND2_X1 U6205 ( .A1(n10113), .A2(n5201), .ZN(n5204) );
  AND2_X1 U6206 ( .A1(n5381), .A2(n5380), .ZN(n5016) );
  AND2_X1 U6207 ( .A1(n5495), .A2(n5493), .ZN(n5017) );
  NAND2_X1 U6208 ( .A1(n4999), .A2(n5342), .ZN(n6398) );
  INV_X1 U6209 ( .A(n6398), .ZN(n5341) );
  INV_X1 U6210 ( .A(n6527), .ZN(n6540) );
  NAND2_X1 U6211 ( .A1(n9114), .A2(n9274), .ZN(n5018) );
  INV_X1 U6212 ( .A(n7366), .ZN(n9959) );
  NAND2_X1 U6213 ( .A1(n6179), .A2(n6178), .ZN(n7366) );
  INV_X1 U6214 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n7782) );
  INV_X1 U6215 ( .A(n8808), .ZN(n6097) );
  AND2_X1 U6216 ( .A1(n6156), .A2(n5123), .ZN(n5019) );
  AND2_X1 U6217 ( .A1(n5959), .A2(n5944), .ZN(n5020) );
  INV_X1 U6218 ( .A(SI_11_), .ZN(n5426) );
  NAND2_X1 U6219 ( .A1(n5949), .A2(n5948), .ZN(n10070) );
  INV_X1 U6220 ( .A(n10070), .ZN(n5202) );
  NAND2_X1 U6221 ( .A1(n5128), .A2(n8799), .ZN(n6884) );
  AND2_X1 U6222 ( .A1(n9322), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n5021) );
  AND2_X1 U6223 ( .A1(n5473), .A2(n7708), .ZN(n5022) );
  INV_X1 U6224 ( .A(n6883), .ZN(n7500) );
  AND2_X1 U6225 ( .A1(n8253), .A2(n4963), .ZN(n5023) );
  OAI21_X1 U6226 ( .B1(n8282), .B2(n5036), .A(n5035), .ZN(n8700) );
  NAND2_X1 U6227 ( .A1(n5057), .A2(n7012), .ZN(n8159) );
  INV_X1 U6228 ( .A(n6555), .ZN(n7936) );
  NAND2_X1 U6229 ( .A1(n5334), .A2(n8943), .ZN(n7790) );
  NAND2_X1 U6230 ( .A1(n5055), .A2(n8049), .ZN(n8149) );
  INV_X1 U6231 ( .A(n7281), .ZN(n8638) );
  AND2_X1 U6232 ( .A1(n6859), .A2(n8919), .ZN(n8891) );
  XNOR2_X1 U6233 ( .A(n6876), .B(n6875), .ZN(n6885) );
  OR2_X1 U6234 ( .A1(n6836), .A2(P2_IR_REG_22__SCAN_IN), .ZN(n5024) );
  NAND2_X1 U6235 ( .A1(n5284), .A2(n7810), .ZN(n7835) );
  INV_X1 U6236 ( .A(n5040), .ZN(n5039) );
  NOR2_X1 U6237 ( .A1(n5288), .A2(n5041), .ZN(n5040) );
  AND2_X1 U6238 ( .A1(n5375), .A2(n5374), .ZN(n5025) );
  AND2_X1 U6239 ( .A1(n5386), .A2(n5385), .ZN(n5026) );
  NOR2_X1 U6240 ( .A1(n8803), .A2(n10230), .ZN(n8787) );
  OR2_X1 U6241 ( .A1(n5021), .A2(n5104), .ZN(n5027) );
  NAND2_X1 U6242 ( .A1(n5309), .A2(n5306), .ZN(n6142) );
  NAND2_X1 U6243 ( .A1(n5779), .A2(n5778), .ZN(n8771) );
  INV_X1 U6244 ( .A(n8771), .ZN(n5192) );
  INV_X1 U6245 ( .A(n10561), .ZN(n10127) );
  INV_X1 U6246 ( .A(n8927), .ZN(n8866) );
  XNOR2_X1 U6247 ( .A(n6833), .B(n6832), .ZN(n8927) );
  INV_X1 U6248 ( .A(n10667), .ZN(n10239) );
  NAND2_X1 U6249 ( .A1(n6838), .A2(n7336), .ZN(n9532) );
  INV_X1 U6250 ( .A(n9532), .ZN(n9498) );
  INV_X1 U6251 ( .A(n6211), .ZN(n5406) );
  NAND2_X1 U6252 ( .A1(n5230), .A2(n6516), .ZN(n7741) );
  INV_X1 U6253 ( .A(n8049), .ZN(n5056) );
  AND2_X1 U6254 ( .A1(n7698), .A2(n7695), .ZN(n9761) );
  NAND2_X1 U6255 ( .A1(n6075), .A2(P1_IR_REG_27__SCAN_IN), .ZN(n6443) );
  NAND2_X1 U6256 ( .A1(n5149), .A2(n6853), .ZN(n7731) );
  INV_X1 U6257 ( .A(n7731), .ZN(n5472) );
  NOR2_X1 U6258 ( .A1(n10439), .A2(n7214), .ZN(n5028) );
  NOR2_X1 U6259 ( .A1(n10401), .A2(n10402), .ZN(n5029) );
  INV_X1 U6260 ( .A(n9073), .ZN(n8090) );
  XNOR2_X1 U6261 ( .A(n6829), .B(P2_IR_REG_19__SCAN_IN), .ZN(n9073) );
  INV_X1 U6262 ( .A(n9080), .ZN(n5215) );
  INV_X1 U6263 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n5071) );
  INV_X1 U6264 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n5094) );
  INV_X1 U6265 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n5092) );
  NAND2_X1 U6266 ( .A1(n5692), .A2(n5691), .ZN(n5694) );
  OAI21_X1 U6267 ( .B1(n5930), .B2(n5929), .A(n5928), .ZN(n5941) );
  INV_X1 U6268 ( .A(n5237), .ZN(n9404) );
  NAND2_X1 U6269 ( .A1(n5399), .A2(n5944), .ZN(n5958) );
  NAND2_X1 U6270 ( .A1(n5254), .A2(n5008), .ZN(n5179) );
  OAI21_X1 U6271 ( .B1(n9482), .B2(n5273), .A(n5270), .ZN(n9436) );
  NAND2_X1 U6272 ( .A1(n10416), .A2(n10417), .ZN(n10415) );
  OAI211_X1 U6273 ( .C1(n5188), .C2(n7566), .A(n7322), .B(n7323), .ZN(P2_U3201) );
  NAND2_X1 U6274 ( .A1(n5318), .A2(n5317), .ZN(n9461) );
  INV_X1 U6275 ( .A(n8840), .ZN(n5256) );
  INV_X1 U6276 ( .A(n9667), .ZN(n6485) );
  INV_X1 U6277 ( .A(n5324), .ZN(n6912) );
  NAND2_X1 U6278 ( .A1(n6513), .A2(n5518), .ZN(n5231) );
  NAND2_X1 U6279 ( .A1(n8875), .A2(n7724), .ZN(n5334) );
  OAI22_X1 U6280 ( .A1(n8825), .A2(n5305), .B1(n5304), .B2(n8826), .ZN(n9711)
         );
  NAND2_X1 U6281 ( .A1(n8815), .A2(n8817), .ZN(n5031) );
  XNOR2_X2 U6282 ( .A(n5033), .B(n5915), .ZN(n6070) );
  NAND3_X1 U6283 ( .A1(n6335), .A2(n9945), .A3(n6334), .ZN(n5052) );
  OAI21_X1 U6284 ( .B1(n8048), .B2(n5056), .A(n5053), .ZN(n5057) );
  AND2_X1 U6285 ( .A1(n5054), .A2(n8150), .ZN(n5053) );
  NAND2_X1 U6286 ( .A1(n5282), .A2(n5058), .ZN(n5281) );
  NAND2_X1 U6287 ( .A1(n5058), .A2(n7811), .ZN(n7810) );
  NAND2_X1 U6288 ( .A1(n5061), .A2(n5060), .ZN(n5059) );
  INV_X1 U6289 ( .A(n7811), .ZN(n5060) );
  NAND3_X1 U6290 ( .A1(n5311), .A2(n9770), .A3(n5064), .ZN(n5063) );
  NAND3_X1 U6291 ( .A1(n5311), .A2(n7101), .A3(n9770), .ZN(n9687) );
  NAND3_X1 U6292 ( .A1(n5396), .A2(n5395), .A3(n5071), .ZN(n5069) );
  NAND2_X1 U6293 ( .A1(n9712), .A2(n4950), .ZN(n5072) );
  OAI21_X1 U6294 ( .B1(n9712), .B2(n5076), .A(n4950), .ZN(n7095) );
  NAND2_X1 U6295 ( .A1(n5072), .A2(n5073), .ZN(n9769) );
  AND2_X2 U6296 ( .A1(n5084), .A2(n5083), .ZN(n5726) );
  NOR2_X1 U6297 ( .A1(n9751), .A2(n9746), .ZN(n9678) );
  NAND2_X1 U6298 ( .A1(n5875), .A2(n5005), .ZN(n5086) );
  NAND2_X1 U6299 ( .A1(n5100), .A2(n5099), .ZN(n10419) );
  NAND2_X1 U6300 ( .A1(n7211), .A2(n5101), .ZN(n5100) );
  NAND2_X1 U6301 ( .A1(n5205), .A2(n5108), .ZN(n5107) );
  NAND2_X1 U6302 ( .A1(n5205), .A2(n5113), .ZN(n5112) );
  INV_X1 U6303 ( .A(n5556), .ZN(n5116) );
  NAND2_X1 U6304 ( .A1(n5124), .A2(n5019), .ZN(P1_U3517) );
  NAND2_X1 U6305 ( .A1(n6115), .A2(n5125), .ZN(n6154) );
  OAI21_X1 U6306 ( .B1(n6884), .B2(P2_D_REG_0__SCAN_IN), .A(n6882), .ZN(n6883)
         );
  NAND2_X1 U6307 ( .A1(n6885), .A2(n5129), .ZN(n5128) );
  XNOR2_X1 U6308 ( .A(n6881), .B(P2_B_REG_SCAN_IN), .ZN(n5129) );
  XNOR2_X1 U6309 ( .A(n8347), .B(n8348), .ZN(n8349) );
  NAND2_X1 U6310 ( .A1(n9170), .A2(n5137), .ZN(n5136) );
  NAND2_X1 U6311 ( .A1(n5486), .A2(n5141), .ZN(n5143) );
  NAND2_X1 U6312 ( .A1(n9289), .A2(n5148), .ZN(n5147) );
  INV_X1 U6313 ( .A(n5149), .ZN(n5148) );
  OR2_X2 U6314 ( .A1(n9539), .A2(n9538), .ZN(n9541) );
  OAI21_X2 U6315 ( .B1(n8775), .B2(n8993), .A(n8998), .ZN(n9539) );
  NAND2_X1 U6316 ( .A1(n5642), .A2(n5155), .ZN(n5153) );
  INV_X1 U6317 ( .A(n5216), .ZN(n5154) );
  NAND2_X1 U6318 ( .A1(n5154), .A2(n5153), .ZN(n5678) );
  NOR2_X1 U6319 ( .A1(n5217), .A2(n5156), .ZN(n5155) );
  NAND2_X1 U6320 ( .A1(n5162), .A2(SI_1_), .ZN(n5161) );
  NAND2_X1 U6321 ( .A1(n5169), .A2(n5168), .ZN(n5162) );
  NAND3_X1 U6322 ( .A1(n5396), .A2(n5395), .A3(P1_DATAO_REG_1__SCAN_IN), .ZN(
        n5168) );
  OAI21_X1 U6323 ( .B1(n5165), .B2(n5162), .A(SI_1_), .ZN(n5525) );
  NAND3_X1 U6324 ( .A1(n5164), .A2(n5163), .A3(n5161), .ZN(n5614) );
  NAND4_X1 U6325 ( .A1(n5167), .A2(n5169), .A3(n5168), .A4(n8455), .ZN(n5163)
         );
  INV_X1 U6326 ( .A(n5805), .ZN(n5173) );
  NAND2_X1 U6327 ( .A1(n5805), .A2(n5804), .ZN(n5807) );
  NAND3_X1 U6328 ( .A1(n7236), .A2(n5187), .A3(P2_IR_REG_2__SCAN_IN), .ZN(
        n5184) );
  INV_X1 U6329 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n5186) );
  AND2_X2 U6330 ( .A1(n5573), .A2(n5190), .ZN(n6120) );
  AND2_X1 U6331 ( .A1(n6074), .A2(n5196), .ZN(n9947) );
  NAND2_X1 U6332 ( .A1(n6074), .A2(n5194), .ZN(n9931) );
  NAND2_X1 U6333 ( .A1(n6074), .A2(n5198), .ZN(n9948) );
  AND2_X1 U6334 ( .A1(n6074), .A2(n9969), .ZN(n7367) );
  INV_X1 U6335 ( .A(n5204), .ZN(n10069) );
  OAI211_X1 U6336 ( .C1(n9071), .C2(n5208), .A(n5209), .B(n5206), .ZN(P2_U3296) );
  NAND3_X1 U6337 ( .A1(n9071), .A2(n5207), .A3(n5215), .ZN(n5206) );
  OAI22_X1 U6338 ( .A1(n5213), .A2(n5212), .B1(n9072), .B2(n8090), .ZN(n5211)
         );
  NOR2_X1 U6339 ( .A1(n9070), .A2(n8090), .ZN(n5212) );
  INV_X1 U6340 ( .A(n9072), .ZN(n5213) );
  OAI21_X1 U6341 ( .B1(n5656), .B2(n5217), .A(n5675), .ZN(n5216) );
  INV_X1 U6342 ( .A(n5533), .ZN(n5217) );
  AOI21_X1 U6343 ( .B1(n5227), .B2(n5226), .A(n8981), .ZN(n8988) );
  NAND3_X1 U6344 ( .A1(n5229), .A2(n5228), .A3(n8976), .ZN(n5227) );
  OAI21_X1 U6345 ( .B1(n8958), .B2(n8965), .A(n9060), .ZN(n5228) );
  OAI21_X1 U6346 ( .B1(n8970), .B2(n8969), .A(n9053), .ZN(n5229) );
  NAND2_X1 U6347 ( .A1(n6850), .A2(n7718), .ZN(n5230) );
  INV_X1 U6348 ( .A(n7544), .ZN(n9148) );
  NAND3_X1 U6349 ( .A1(n5234), .A2(n8982), .A3(n5232), .ZN(n8747) );
  NAND3_X1 U6350 ( .A1(n8673), .A2(n8696), .A3(n4974), .ZN(n5234) );
  NAND2_X1 U6351 ( .A1(n7791), .A2(n6548), .ZN(n5241) );
  NAND3_X1 U6352 ( .A1(n5241), .A2(n7961), .A3(n5240), .ZN(n6562) );
  OAI21_X1 U6353 ( .B1(n7791), .B2(n4975), .A(n6548), .ZN(n6555) );
  NAND2_X1 U6354 ( .A1(n7959), .A2(n5245), .ZN(n5242) );
  NAND2_X1 U6355 ( .A1(n5242), .A2(n5243), .ZN(n6591) );
  XNOR2_X2 U6356 ( .A(n6480), .B(P2_IR_REG_30__SCAN_IN), .ZN(n9664) );
  AND2_X2 U6357 ( .A1(n6484), .A2(n6483), .ZN(n9667) );
  NOR2_X1 U6358 ( .A1(n9052), .A2(n9408), .ZN(n5258) );
  NAND2_X1 U6359 ( .A1(n8773), .A2(n5260), .ZN(n5259) );
  NAND2_X1 U6360 ( .A1(n5259), .A2(n5262), .ZN(n6726) );
  AOI21_X1 U6361 ( .B1(n6790), .B2(n6789), .A(n6788), .ZN(n9427) );
  MUX2_X1 U6362 ( .A(P2_IR_REG_0__SCAN_IN), .B(n9677), .S(n6515), .Z(n7544) );
  NAND2_X1 U6363 ( .A1(n6564), .A2(n6563), .ZN(n7959) );
  NAND2_X1 U6364 ( .A1(n6525), .A2(n6524), .ZN(n7726) );
  NAND2_X1 U6365 ( .A1(n6640), .A2(n6639), .ZN(n8386) );
  INV_X1 U6366 ( .A(n9436), .ZN(n6790) );
  NOR2_X1 U6367 ( .A1(n6623), .A2(n4979), .ZN(n6624) );
  OR2_X1 U6368 ( .A1(n7134), .A2(n7133), .ZN(n5303) );
  INV_X1 U6369 ( .A(n9711), .ZN(n7079) );
  OAI21_X1 U6370 ( .B1(n5897), .B2(n5310), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n6067) );
  NAND2_X1 U6371 ( .A1(n5897), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5309) );
  NAND2_X1 U6372 ( .A1(n9769), .A2(n9772), .ZN(n5311) );
  NAND2_X1 U6373 ( .A1(n8672), .A2(n4955), .ZN(n5312) );
  NAND2_X1 U6374 ( .A1(n9505), .A2(n5319), .ZN(n5318) );
  INV_X1 U6375 ( .A(n5332), .ZN(n9451) );
  NAND2_X1 U6376 ( .A1(n5334), .A2(n5333), .ZN(n7934) );
  AND3_X2 U6377 ( .A1(n6727), .A2(n5009), .A3(n5499), .ZN(n6481) );
  NAND2_X1 U6378 ( .A1(n6727), .A2(n5499), .ZN(n6496) );
  NAND3_X1 U6379 ( .A1(n6727), .A2(n5499), .A3(n5336), .ZN(n6498) );
  NAND2_X1 U6380 ( .A1(n5338), .A2(n5337), .ZN(n6861) );
  INV_X2 U6381 ( .A(n6509), .ZN(n6720) );
  NAND2_X1 U6382 ( .A1(n4946), .A2(n5343), .ZN(n6239) );
  INV_X1 U6383 ( .A(n9941), .ZN(n5352) );
  XNOR2_X1 U6384 ( .A(n9937), .B(n9945), .ZN(n5353) );
  NAND2_X2 U6385 ( .A1(n10046), .A2(n10045), .ZN(n10044) );
  OAI21_X2 U6386 ( .B1(n8662), .B2(n5358), .A(n5356), .ZN(n8808) );
  NAND2_X1 U6387 ( .A1(n10079), .A2(n5362), .ZN(n6345) );
  INV_X1 U6388 ( .A(n9981), .ZN(n5367) );
  NAND2_X1 U6389 ( .A1(n9981), .A2(n5369), .ZN(n5363) );
  NAND2_X1 U6390 ( .A1(n5363), .A2(n5364), .ZN(n9936) );
  NAND2_X1 U6391 ( .A1(n5368), .A2(n5369), .ZN(n7362) );
  OAI21_X1 U6392 ( .B1(n10441), .B2(n5389), .A(n5388), .ZN(n10456) );
  NAND2_X1 U6393 ( .A1(n5399), .A2(n5020), .ZN(n5961) );
  NOR2_X1 U6394 ( .A1(n5400), .A2(n6383), .ZN(n5407) );
  NAND2_X1 U6395 ( .A1(n5403), .A2(n5402), .ZN(n5401) );
  NAND2_X1 U6396 ( .A1(n6217), .A2(n8847), .ZN(n5403) );
  NAND2_X1 U6397 ( .A1(n6341), .A2(n6228), .ZN(n6383) );
  NAND2_X1 U6398 ( .A1(n5761), .A2(n5561), .ZN(n5774) );
  OAI21_X2 U6399 ( .B1(n5761), .B2(n5421), .A(n5419), .ZN(n5805) );
  NAND2_X1 U6400 ( .A1(n6013), .A2(n5434), .ZN(n6033) );
  NAND2_X1 U6401 ( .A1(n6013), .A2(n6012), .ZN(n6016) );
  NAND2_X1 U6402 ( .A1(n5436), .A2(n7853), .ZN(n5632) );
  AND3_X2 U6403 ( .A1(n5438), .A2(n5439), .A3(n5437), .ZN(n5618) );
  NAND2_X1 U6404 ( .A1(n6116), .A2(n5004), .ZN(n5437) );
  NAND2_X1 U6405 ( .A1(n6031), .A2(n6030), .ZN(n9974) );
  NOR2_X1 U6406 ( .A1(n5679), .A2(n5445), .ZN(n5697) );
  NAND2_X1 U6407 ( .A1(n8135), .A2(n5448), .ZN(n5447) );
  NAND2_X1 U6408 ( .A1(n10058), .A2(n5456), .ZN(n5455) );
  INV_X1 U6409 ( .A(n5457), .ZN(n10059) );
  NAND2_X1 U6410 ( .A1(n10138), .A2(n5462), .ZN(n5461) );
  NAND2_X1 U6411 ( .A1(n7710), .A2(n7731), .ZN(n5470) );
  NAND2_X1 U6412 ( .A1(n7876), .A2(n5483), .ZN(n5480) );
  INV_X1 U6413 ( .A(n8720), .ZN(n5496) );
  NAND2_X1 U6414 ( .A1(n8720), .A2(n5490), .ZN(n5486) );
  AOI21_X1 U6415 ( .B1(n7373), .B2(n10674), .A(n7371), .ZN(n7372) );
  NAND2_X1 U6416 ( .A1(n5633), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n5627) );
  NAND2_X1 U6417 ( .A1(n8912), .A2(n8911), .ZN(n9072) );
  NAND2_X1 U6418 ( .A1(n7369), .A2(n7368), .ZN(n7373) );
  NAND2_X1 U6419 ( .A1(n9955), .A2(n10667), .ZN(n7369) );
  INV_X1 U6420 ( .A(n8787), .ZN(n8802) );
  NAND2_X1 U6421 ( .A1(n7373), .A2(n10646), .ZN(n7376) );
  NAND2_X1 U6422 ( .A1(n7344), .A2(n9627), .ZN(n6911) );
  CLKBUF_X1 U6423 ( .A(n7838), .Z(n10559) );
  NOR2_X2 U6425 ( .A1(n5523), .A2(n8566), .ZN(n5612) );
  XNOR2_X1 U6426 ( .A(n6116), .B(n6119), .ZN(n8759) );
  OAI21_X1 U6427 ( .B1(n6375), .B2(n6374), .A(n6070), .ZN(n6376) );
  NAND2_X1 U6428 ( .A1(n6382), .A2(n7184), .ZN(n6441) );
  NAND2_X1 U6429 ( .A1(n5601), .A2(n5600), .ZN(n5624) );
  INV_X1 U6430 ( .A(n5601), .ZN(n10280) );
  AOI21_X1 U6431 ( .B1(n6917), .B2(n6918), .A(n6916), .ZN(n6926) );
  NAND2_X1 U6432 ( .A1(n8787), .A2(n8790), .ZN(n10147) );
  AOI21_X2 U6433 ( .B1(n9410), .B2(n6869), .A(n9049), .ZN(n6919) );
  XNOR2_X1 U6434 ( .A(n9104), .B(n9105), .ZN(n9162) );
  AND2_X2 U6435 ( .A1(n7348), .A2(n9659), .ZN(n10695) );
  NAND2_X2 U6436 ( .A1(n9149), .A2(n10677), .ZN(n10641) );
  NOR2_X1 U6437 ( .A1(n9052), .A2(n9594), .ZN(n6907) );
  INV_X1 U6438 ( .A(n7176), .ZN(n7184) );
  INV_X1 U6439 ( .A(n10646), .ZN(n10669) );
  AND2_X2 U6440 ( .A1(n6153), .A2(n6146), .ZN(n10646) );
  INV_X1 U6441 ( .A(n10414), .ZN(n7441) );
  AND2_X1 U6442 ( .A1(n7347), .A2(n7346), .ZN(n5503) );
  INV_X1 U6443 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n6450) );
  AND4_X1 U6444 ( .A1(n6112), .A2(n6111), .A3(n6110), .A4(n6109), .ZN(n9942)
         );
  OR2_X1 U6445 ( .A1(n9598), .A2(n9604), .ZN(n5506) );
  INV_X1 U6446 ( .A(n10065), .ZN(n9798) );
  AND4_X1 U6447 ( .A1(n5976), .A2(n5975), .A3(n5974), .A4(n5973), .ZN(n10065)
         );
  OR2_X1 U6448 ( .A1(n10674), .A2(n7370), .ZN(n5508) );
  OR2_X1 U6449 ( .A1(n9052), .A2(n9654), .ZN(n5509) );
  OR2_X1 U6450 ( .A1(n9959), .A2(n10219), .ZN(n5510) );
  OR2_X1 U6451 ( .A1(n9959), .A2(n10267), .ZN(n5511) );
  INV_X1 U6452 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n6455) );
  INV_X1 U6453 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n5520) );
  NAND2_X1 U6454 ( .A1(n10287), .A2(n7398), .ZN(n10143) );
  INV_X1 U6455 ( .A(n10143), .ZN(n10557) );
  INV_X1 U6456 ( .A(n10267), .ZN(n6155) );
  AND2_X1 U6457 ( .A1(n7822), .A2(n6948), .ZN(n10649) );
  OR2_X1 U6458 ( .A1(n9807), .A2(n8038), .ZN(n5514) );
  OAI211_X1 U6459 ( .C1(n6540), .C2(n6745), .A(n6744), .B(n6743), .ZN(n9468)
         );
  INV_X1 U6460 ( .A(n8323), .ZN(n6094) );
  INV_X1 U6461 ( .A(n8167), .ZN(n5744) );
  OR2_X1 U6462 ( .A1(n7498), .A2(n9078), .ZN(n5515) );
  OR2_X1 U6463 ( .A1(n10225), .A2(n9800), .ZN(n5516) );
  AND2_X1 U6464 ( .A1(n6518), .A2(n6517), .ZN(n5517) );
  AND3_X1 U6465 ( .A1(n6512), .A2(n6511), .A3(n6510), .ZN(n5518) );
  INV_X1 U6466 ( .A(n8928), .ZN(n8929) );
  MUX2_X1 U6467 ( .A(n6347), .B(n6352), .S(n6339), .Z(n6319) );
  INV_X1 U6468 ( .A(n8839), .ZN(n6923) );
  INV_X1 U6469 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n7207) );
  INV_X1 U6470 ( .A(n9802), .ZN(n5820) );
  INV_X1 U6471 ( .A(n9100), .ZN(n9102) );
  NOR2_X1 U6472 ( .A1(n10376), .A2(n7207), .ZN(n7208) );
  INV_X1 U6473 ( .A(n6381), .ZN(n6375) );
  INV_X1 U6474 ( .A(n10029), .ZN(n6102) );
  INV_X1 U6475 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n5750) );
  OR4_X1 U6476 ( .A1(P1_D_REG_31__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_29__SCAN_IN), .A4(P1_D_REG_28__SCAN_IN), .ZN(n6132) );
  NAND2_X1 U6477 ( .A1(n9102), .A2(n9580), .ZN(n9103) );
  NAND2_X1 U6478 ( .A1(n8868), .A2(n8867), .ZN(n8909) );
  INV_X1 U6479 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n8493) );
  INV_X1 U6480 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n8723) );
  INV_X1 U6481 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n9195) );
  INV_X1 U6482 ( .A(n9274), .ZN(n6814) );
  NAND2_X1 U6483 ( .A1(n6621), .A2(n4987), .ZN(n8213) );
  INV_X1 U6484 ( .A(n9714), .ZN(n7078) );
  INV_X1 U6485 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n5598) );
  NOR2_X1 U6486 ( .A1(n5907), .A2(n5906), .ZN(n5921) );
  NOR2_X1 U6487 ( .A1(n5751), .A2(n5750), .ZN(n5766) );
  OR2_X1 U6488 ( .A1(n5655), .A2(n7439), .ZN(n5647) );
  INV_X1 U6489 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n6062) );
  INV_X1 U6490 ( .A(SI_13_), .ZN(n8544) );
  INV_X1 U6491 ( .A(SI_8_), .ZN(n8557) );
  INV_X1 U6492 ( .A(n9221), .ZN(n9095) );
  INV_X1 U6493 ( .A(n9070), .ZN(n8911) );
  NAND2_X1 U6494 ( .A1(n6794), .A2(n6793), .ZN(n6805) );
  NAND2_X1 U6495 ( .A1(n6460), .A2(n8493), .ZN(n6750) );
  INV_X1 U6496 ( .A(n6929), .ZN(n6842) );
  OAI21_X1 U6497 ( .B1(n8159), .B2(n8161), .A(n8160), .ZN(n7017) );
  OR2_X1 U6498 ( .A1(n9781), .A2(n9782), .ZN(n7149) );
  NOR2_X1 U6499 ( .A1(n7819), .A2(n7161), .ZN(n7183) );
  NOR2_X1 U6500 ( .A1(n5815), .A2(n5598), .ZN(n5840) );
  OR2_X1 U6501 ( .A1(n5797), .A2(n7803), .ZN(n5813) );
  AND2_X1 U6502 ( .A1(n6170), .A2(n6108), .ZN(n9957) );
  NAND2_X1 U6503 ( .A1(n5032), .A2(n8290), .ZN(n5772) );
  OR2_X1 U6504 ( .A1(n6372), .A2(n6145), .ZN(n7187) );
  INV_X1 U6505 ( .A(n6372), .ZN(n7398) );
  INV_X1 U6506 ( .A(SI_24_), .ZN(n6010) );
  INV_X1 U6507 ( .A(SI_17_), .ZN(n5865) );
  AND2_X1 U6508 ( .A1(n5532), .A2(n5533), .ZN(n5656) );
  INV_X1 U6509 ( .A(n9446), .ZN(n9165) );
  NAND2_X1 U6510 ( .A1(n9096), .A2(n9500), .ZN(n9097) );
  NAND2_X1 U6511 ( .A1(n9085), .A2(n9278), .ZN(n9086) );
  NAND2_X1 U6512 ( .A1(n9093), .A2(n9484), .ZN(n9094) );
  NAND2_X1 U6513 ( .A1(n6462), .A2(n6461), .ZN(n6769) );
  INV_X1 U6514 ( .A(n9608), .ZN(n9516) );
  INV_X1 U6515 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n7711) );
  INV_X1 U6516 ( .A(n7498), .ZN(n10679) );
  INV_X1 U6517 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n6908) );
  OR2_X1 U6518 ( .A1(n9060), .A2(n6903), .ZN(n6937) );
  OAI22_X1 U6519 ( .A1(n8840), .A2(n5515), .B1(n9618), .B2(n8839), .ZN(n8841)
         );
  INV_X1 U6520 ( .A(n9277), .ZN(n9604) );
  INV_X1 U6521 ( .A(n9278), .ZN(n9617) );
  INV_X1 U6522 ( .A(n9284), .ZN(n8267) );
  INV_X1 U6523 ( .A(n9286), .ZN(n8010) );
  NAND2_X1 U6524 ( .A1(n7520), .A2(n9060), .ZN(n9515) );
  XNOR2_X1 U6525 ( .A(n6986), .B(n6963), .ZN(n6993) );
  AND4_X1 U6526 ( .A1(n5859), .A2(n5858), .A3(n5857), .A4(n5856), .ZN(n10125)
         );
  AND2_X1 U6527 ( .A1(n6253), .A2(n6395), .ZN(n7946) );
  OR2_X1 U6528 ( .A1(n10619), .A2(n7829), .ZN(n10612) );
  OR2_X1 U6529 ( .A1(n7654), .A2(n7184), .ZN(n10663) );
  AND2_X1 U6530 ( .A1(n6103), .A2(n6342), .ZN(n10561) );
  OAI22_X1 U6531 ( .A1(n7944), .A2(n7946), .B1(n7928), .B2(n9808), .ZN(n8026)
         );
  OR2_X1 U6532 ( .A1(n6323), .A2(n7184), .ZN(n10539) );
  INV_X1 U6533 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n6143) );
  INV_X1 U6534 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5915) );
  AND2_X1 U6535 ( .A1(n5568), .A2(n5567), .ZN(n5804) );
  INV_X1 U6536 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n9237) );
  INV_X1 U6537 ( .A(n5639), .ZN(n5641) );
  INV_X1 U6538 ( .A(n9283), .ZN(n8353) );
  OR2_X1 U6539 ( .A1(n6942), .A2(n6509), .ZN(n8857) );
  AND3_X1 U6540 ( .A1(n6737), .A2(n6736), .A3(n6735), .ZN(n9517) );
  AND2_X1 U6541 ( .A1(P2_U3893), .A2(n6845), .ZN(n10504) );
  INV_X1 U6542 ( .A(n10412), .ZN(n10495) );
  INV_X1 U6543 ( .A(n7566), .ZN(n10505) );
  OR2_X1 U6544 ( .A1(n9618), .A2(n10679), .ZN(n10585) );
  INV_X1 U6545 ( .A(n10677), .ZN(n10634) );
  INV_X1 U6546 ( .A(n9493), .ZN(n9547) );
  NAND2_X1 U6547 ( .A1(n8927), .A2(n8346), .ZN(n9618) );
  NOR2_X1 U6548 ( .A1(n7335), .A2(n6900), .ZN(n6939) );
  AND2_X1 U6549 ( .A1(n7775), .A2(n5515), .ZN(n9615) );
  INV_X1 U6550 ( .A(n9615), .ZN(n9623) );
  INV_X1 U6551 ( .A(n7326), .ZN(n7327) );
  AND2_X1 U6552 ( .A1(n7182), .A2(n9821), .ZN(n9787) );
  AOI21_X1 U6553 ( .B1(n6439), .B2(n7176), .A(n8381), .ZN(n6440) );
  INV_X1 U6554 ( .A(n10031), .ZN(n9706) );
  AND4_X1 U6555 ( .A1(n5911), .A2(n5910), .A3(n5909), .A4(n5908), .ZN(n10124)
         );
  INV_X1 U6556 ( .A(n9926), .ZN(n10519) );
  INV_X1 U6557 ( .A(n10524), .ZN(n9894) );
  INV_X1 U6558 ( .A(n10663), .ZN(n10552) );
  AND2_X1 U6559 ( .A1(n6426), .A2(n10060), .ZN(n10078) );
  AND2_X1 U6560 ( .A1(n6300), .A2(n6417), .ZN(n10121) );
  NAND2_X1 U6561 ( .A1(n10274), .A2(n7179), .ZN(n10606) );
  NAND2_X1 U6562 ( .A1(n8028), .A2(n10539), .ZN(n10667) );
  AND2_X1 U6563 ( .A1(n6152), .A2(n7161), .ZN(n7820) );
  INV_X1 U6564 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n6123) );
  AND2_X1 U6565 ( .A1(n5809), .A2(n5833), .ZN(n8108) );
  AND2_X1 U6566 ( .A1(n5699), .A2(n5698), .ZN(n7643) );
  OR3_X1 U6567 ( .A1(n6885), .A2(n6881), .A3(n7470), .ZN(n7491) );
  NAND2_X1 U6568 ( .A1(n7511), .A2(n9659), .ZN(n9254) );
  INV_X1 U6569 ( .A(n9251), .ZN(n9270) );
  NAND2_X1 U6570 ( .A1(n6812), .A2(n6811), .ZN(n9274) );
  INV_X1 U6571 ( .A(n8698), .ZN(n9281) );
  OR2_X1 U6572 ( .A1(P2_U3150), .A2(n7318), .ZN(n10412) );
  INV_X1 U6573 ( .A(n10370), .ZN(n10511) );
  NAND2_X1 U6574 ( .A1(n10641), .A2(n10683), .ZN(n9493) );
  OR2_X1 U6575 ( .A1(n9624), .A2(n9618), .ZN(n9594) );
  INV_X1 U6576 ( .A(n9624), .ZN(n9627) );
  NAND2_X2 U6577 ( .A1(n6939), .A2(n6906), .ZN(n9624) );
  OR2_X1 U6578 ( .A1(n9600), .A2(n9599), .ZN(n9656) );
  INV_X1 U6579 ( .A(n10695), .ZN(n10692) );
  NAND2_X1 U6580 ( .A1(n6884), .A2(n9659), .ZN(n7467) );
  INV_X1 U6581 ( .A(n7277), .ZN(n9322) );
  OR2_X1 U6582 ( .A1(n7328), .A2(n7173), .ZN(n7198) );
  INV_X1 U6583 ( .A(n8665), .ZN(n10662) );
  INV_X1 U6584 ( .A(n9789), .ZN(n8745) );
  INV_X1 U6585 ( .A(n9784), .ZN(n9778) );
  AND4_X1 U6586 ( .A1(n6175), .A2(n6174), .A3(n6173), .A4(n6172), .ZN(n8281)
         );
  INV_X1 U6587 ( .A(n10124), .ZN(n9799) );
  OR2_X1 U6588 ( .A1(n7421), .A2(n7419), .ZN(n7478) );
  NAND2_X1 U6589 ( .A1(n7416), .A2(n10294), .ZN(n9926) );
  INV_X1 U6590 ( .A(n10615), .ZN(n10154) );
  NAND2_X1 U6591 ( .A1(n7329), .A2(n6148), .ZN(n6149) );
  NAND2_X1 U6592 ( .A1(n10646), .A2(n10649), .ZN(n10219) );
  INV_X1 U6593 ( .A(n10102), .ZN(n10262) );
  NAND2_X1 U6594 ( .A1(n10674), .A2(n10649), .ZN(n10267) );
  NAND2_X1 U6595 ( .A1(n6153), .A2(n7820), .ZN(n10671) );
  INV_X2 U6596 ( .A(n10671), .ZN(n10674) );
  INV_X1 U6597 ( .A(n6141), .ZN(n8838) );
  INV_X1 U6598 ( .A(n10286), .ZN(n10290) );
  NAND2_X1 U6599 ( .A1(n6911), .A2(n6910), .ZN(P2_U3487) );
  INV_X1 U6600 ( .A(n7372), .ZN(P1_U3518) );
  MUX2_X1 U6601 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .S(n5528), .Z(n5519) );
  OAI21_X1 U6602 ( .B1(n5519), .B2(SI_2_), .A(n5527), .ZN(n5640) );
  INV_X1 U6603 ( .A(n5640), .ZN(n5526) );
  INV_X1 U6604 ( .A(SI_1_), .ZN(n8455) );
  INV_X1 U6605 ( .A(n5614), .ZN(n5524) );
  INV_X1 U6606 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5522) );
  INV_X1 U6607 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5521) );
  MUX2_X1 U6608 ( .A(n5522), .B(n5521), .S(n5528), .Z(n5523) );
  NAND2_X1 U6609 ( .A1(n5524), .A2(n5612), .ZN(n5616) );
  NAND2_X1 U6610 ( .A1(n5616), .A2(n5525), .ZN(n5639) );
  NAND2_X1 U6611 ( .A1(n5526), .A2(n5639), .ZN(n5642) );
  INV_X1 U6612 ( .A(SI_3_), .ZN(n5529) );
  NAND2_X1 U6613 ( .A1(n5530), .A2(n5529), .ZN(n5532) );
  NAND2_X1 U6614 ( .A1(n5531), .A2(SI_3_), .ZN(n5533) );
  MUX2_X1 U6615 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .S(n5528), .Z(n5534) );
  NAND2_X1 U6616 ( .A1(n5534), .A2(SI_4_), .ZN(n5537) );
  INV_X1 U6617 ( .A(n5534), .ZN(n5535) );
  INV_X1 U6618 ( .A(SI_4_), .ZN(n8448) );
  NAND2_X1 U6619 ( .A1(n5535), .A2(n8448), .ZN(n5536) );
  AND2_X1 U6620 ( .A1(n5537), .A2(n5536), .ZN(n5675) );
  MUX2_X1 U6621 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .S(n5528), .Z(n5538) );
  NAND2_X1 U6622 ( .A1(n5538), .A2(SI_5_), .ZN(n5542) );
  INV_X1 U6623 ( .A(n5538), .ZN(n5540) );
  INV_X1 U6624 ( .A(SI_5_), .ZN(n5539) );
  NAND2_X1 U6625 ( .A1(n5540), .A2(n5539), .ZN(n5541) );
  AND2_X1 U6626 ( .A1(n5542), .A2(n5541), .ZN(n5691) );
  NAND2_X1 U6627 ( .A1(n5694), .A2(n5542), .ZN(n5710) );
  MUX2_X1 U6628 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n7435), .Z(n5543) );
  NAND2_X1 U6629 ( .A1(n5543), .A2(SI_6_), .ZN(n5546) );
  INV_X1 U6630 ( .A(n5543), .ZN(n5544) );
  INV_X1 U6631 ( .A(SI_6_), .ZN(n8556) );
  NAND2_X1 U6632 ( .A1(n5544), .A2(n8556), .ZN(n5545) );
  AND2_X1 U6633 ( .A1(n5546), .A2(n5545), .ZN(n5709) );
  NAND2_X1 U6634 ( .A1(n5710), .A2(n5709), .ZN(n5712) );
  MUX2_X1 U6635 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n7435), .Z(n5547) );
  NAND2_X1 U6636 ( .A1(n5547), .A2(SI_7_), .ZN(n5550) );
  INV_X1 U6637 ( .A(n5547), .ZN(n5548) );
  INV_X1 U6638 ( .A(SI_7_), .ZN(n8548) );
  NAND2_X1 U6639 ( .A1(n5548), .A2(n8548), .ZN(n5549) );
  AND2_X1 U6640 ( .A1(n5550), .A2(n5549), .ZN(n5722) );
  MUX2_X1 U6641 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(P2_DATAO_REG_8__SCAN_IN), 
        .S(n7435), .Z(n5552) );
  XNOR2_X1 U6642 ( .A(n5552), .B(SI_8_), .ZN(n5731) );
  INV_X1 U6643 ( .A(n5731), .ZN(n5551) );
  INV_X1 U6644 ( .A(n5552), .ZN(n5553) );
  NAND2_X1 U6645 ( .A1(n5553), .A2(n8557), .ZN(n5554) );
  MUX2_X1 U6646 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(P2_DATAO_REG_9__SCAN_IN), 
        .S(n7435), .Z(n5555) );
  XNOR2_X1 U6647 ( .A(n5555), .B(n8549), .ZN(n5745) );
  NOR2_X1 U6648 ( .A1(n5555), .A2(SI_9_), .ZN(n5556) );
  MUX2_X1 U6649 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .S(n7435), .Z(n5557) );
  NAND2_X1 U6650 ( .A1(n5557), .A2(SI_10_), .ZN(n5561) );
  INV_X1 U6651 ( .A(n5557), .ZN(n5558) );
  INV_X1 U6652 ( .A(SI_10_), .ZN(n8547) );
  NAND2_X1 U6653 ( .A1(n5558), .A2(n8547), .ZN(n5559) );
  NAND2_X1 U6654 ( .A1(n5561), .A2(n5559), .ZN(n5759) );
  INV_X1 U6655 ( .A(n5759), .ZN(n5560) );
  MUX2_X1 U6656 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .S(n7435), .Z(n5562) );
  XNOR2_X1 U6657 ( .A(n5562), .B(SI_11_), .ZN(n5773) );
  MUX2_X1 U6658 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .S(n7435), .Z(n5563) );
  NAND2_X1 U6659 ( .A1(n5563), .A2(SI_12_), .ZN(n5564) );
  OAI21_X1 U6660 ( .B1(n5563), .B2(SI_12_), .A(n5564), .ZN(n5787) );
  MUX2_X1 U6661 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n7435), .Z(n5565) );
  NAND2_X1 U6662 ( .A1(n5565), .A2(SI_13_), .ZN(n5568) );
  INV_X1 U6663 ( .A(n5565), .ZN(n5566) );
  NAND2_X1 U6664 ( .A1(n5566), .A2(n8544), .ZN(n5567) );
  MUX2_X1 U6665 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n7435), .Z(n5826) );
  XNOR2_X1 U6666 ( .A(n5826), .B(SI_14_), .ZN(n5827) );
  NOR2_X2 U6667 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5644) );
  NAND2_X1 U6668 ( .A1(n5644), .A2(n5569), .ZN(n5679) );
  NAND3_X1 U6669 ( .A1(n5867), .A2(n5866), .A3(n5869), .ZN(n5574) );
  NOR2_X1 U6670 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), .ZN(
        n5576) );
  NOR2_X1 U6671 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_20__SCAN_IN), .ZN(
        n5575) );
  NAND4_X1 U6672 ( .A1(n5868), .A2(n5576), .A3(n5575), .A4(n5899), .ZN(n5578)
         );
  NAND3_X1 U6673 ( .A1(n5871), .A2(n5085), .A3(n6062), .ZN(n5577) );
  NOR2_X1 U6674 ( .A1(n5578), .A2(n5577), .ZN(n5579) );
  NAND2_X2 U6675 ( .A1(n5589), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6116) );
  INV_X1 U6676 ( .A(n5587), .ZN(n5580) );
  NAND2_X1 U6677 ( .A1(n5580), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5581) );
  INV_X4 U6678 ( .A(n5655), .ZN(n6217) );
  NAND2_X1 U6679 ( .A1(n7668), .A2(n6217), .ZN(n5585) );
  INV_X1 U6680 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n7669) );
  OR2_X1 U6681 ( .A1(n4949), .A2(P1_IR_REG_13__SCAN_IN), .ZN(n5833) );
  NAND2_X1 U6682 ( .A1(n5833), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5582) );
  XNOR2_X1 U6683 ( .A(n5582), .B(P1_IR_REG_14__SCAN_IN), .ZN(n8229) );
  INV_X1 U6684 ( .A(n8229), .ZN(n7670) );
  OAI22_X1 U6685 ( .A1(n5902), .A2(n7669), .B1(n5618), .B2(n7670), .ZN(n5583)
         );
  INV_X1 U6686 ( .A(n5583), .ZN(n5584) );
  NAND2_X2 U6687 ( .A1(n5585), .A2(n5584), .ZN(n10230) );
  NAND2_X1 U6688 ( .A1(n5587), .A2(n5586), .ZN(n5588) );
  NOR2_X2 U6689 ( .A1(n5589), .A2(n5588), .ZN(n5593) );
  INV_X1 U6690 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n5590) );
  OR2_X1 U6691 ( .A1(n5593), .A2(n5590), .ZN(n5591) );
  INV_X1 U6692 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n5592) );
  NAND2_X1 U6693 ( .A1(n5593), .A2(n5592), .ZN(n5595) );
  NAND2_X2 U6694 ( .A1(n5594), .A2(n5595), .ZN(n5600) );
  INV_X1 U6695 ( .A(n5600), .ZN(n10283) );
  XNOR2_X2 U6696 ( .A(n5597), .B(n5596), .ZN(n5601) );
  AND2_X4 U6697 ( .A1(n10283), .A2(n5601), .ZN(n5796) );
  NAND2_X1 U6698 ( .A1(n6220), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n5606) );
  NAND2_X1 U6699 ( .A1(n5685), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n5703) );
  NOR2_X1 U6700 ( .A1(n5703), .A2(n5702), .ZN(n5716) );
  NAND2_X1 U6701 ( .A1(n5716), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5738) );
  NAND2_X1 U6702 ( .A1(n5780), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n5797) );
  AND2_X1 U6703 ( .A1(n5815), .A2(n5598), .ZN(n5599) );
  NOR2_X1 U6704 ( .A1(n5840), .A2(n5599), .ZN(n8819) );
  NAND2_X1 U6705 ( .A1(n6171), .A2(n8819), .ZN(n5605) );
  NAND2_X1 U6706 ( .A1(n6222), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5604) );
  INV_X1 U6707 ( .A(n5600), .ZN(n5602) );
  NAND2_X1 U6708 ( .A1(n6221), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n5603) );
  NAND4_X1 U6709 ( .A1(n5606), .A2(n5605), .A3(n5604), .A4(n5603), .ZN(n9801)
         );
  NAND2_X1 U6710 ( .A1(n5634), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n5611) );
  NAND2_X1 U6711 ( .A1(n5633), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n5610) );
  INV_X1 U6712 ( .A(n5625), .ZN(n5607) );
  NAND2_X1 U6713 ( .A1(n5607), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5609) );
  NAND2_X1 U6714 ( .A1(n5796), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n5608) );
  INV_X1 U6715 ( .A(n5612), .ZN(n5613) );
  NAND2_X1 U6716 ( .A1(n5614), .A2(n5613), .ZN(n5615) );
  NAND2_X1 U6717 ( .A1(n5616), .A2(n5615), .ZN(n7437) );
  INV_X1 U6718 ( .A(n7437), .ZN(n5617) );
  NAND2_X1 U6719 ( .A1(n6217), .A2(n5617), .ZN(n5622) );
  NAND2_X1 U6720 ( .A1(n5660), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n5621) );
  NAND2_X1 U6721 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5619) );
  XNOR2_X1 U6722 ( .A(n5619), .B(P1_IR_REG_1__SCAN_IN), .ZN(n9812) );
  NAND2_X1 U6723 ( .A1(n5645), .A2(n9812), .ZN(n5620) );
  INV_X1 U6724 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n9820) );
  INV_X1 U6725 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n5623) );
  OAI22_X1 U6726 ( .A1(n5625), .A2(n9820), .B1(n5624), .B2(n5623), .ZN(n5626)
         );
  INV_X1 U6727 ( .A(n5626), .ZN(n5629) );
  NAND2_X1 U6728 ( .A1(n7435), .A2(SI_0_), .ZN(n5630) );
  XNOR2_X1 U6729 ( .A(n5630), .B(P2_DATAO_REG_0__SCAN_IN), .ZN(n10295) );
  MUX2_X1 U6730 ( .A(n10295), .B(P1_IR_REG_0__SCAN_IN), .S(n5645), .Z(n7831)
         );
  NAND2_X1 U6731 ( .A1(n7932), .A2(n7831), .ZN(n7853) );
  INV_X1 U6732 ( .A(n6960), .ZN(n6083) );
  NAND2_X1 U6733 ( .A1(n6083), .A2(n6965), .ZN(n5631) );
  NAND2_X1 U6734 ( .A1(n5632), .A2(n5631), .ZN(n10548) );
  NAND2_X1 U6735 ( .A1(n5796), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5638) );
  NAND2_X1 U6736 ( .A1(n5633), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n5637) );
  NAND2_X1 U6737 ( .A1(n5686), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5636) );
  NAND2_X1 U6738 ( .A1(n5634), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5635) );
  NAND2_X1 U6739 ( .A1(n5660), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n5648) );
  NAND2_X1 U6740 ( .A1(n5641), .A2(n5640), .ZN(n5643) );
  NAND2_X1 U6741 ( .A1(n5643), .A2(n5642), .ZN(n7439) );
  OR2_X1 U6742 ( .A1(n5644), .A2(n5590), .ZN(n5662) );
  NAND2_X1 U6743 ( .A1(n5645), .A2(n9831), .ZN(n5646) );
  NAND2_X1 U6744 ( .A1(n10548), .A2(n10549), .ZN(n5650) );
  INV_X1 U6745 ( .A(n6970), .ZN(n6085) );
  NAND2_X1 U6746 ( .A1(n6085), .A2(n6971), .ZN(n5649) );
  NAND2_X1 U6747 ( .A1(n5650), .A2(n5649), .ZN(n7982) );
  INV_X1 U6748 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n7812) );
  NAND2_X1 U6749 ( .A1(n6171), .A2(n7812), .ZN(n5654) );
  NAND2_X1 U6750 ( .A1(n5796), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n5653) );
  NAND2_X1 U6751 ( .A1(n5686), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5652) );
  INV_X2 U6752 ( .A(n5624), .ZN(n6222) );
  NAND2_X1 U6753 ( .A1(n6222), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n5651) );
  AND4_X2 U6754 ( .A1(n5654), .A2(n5653), .A3(n5652), .A4(n5651), .ZN(n6982)
         );
  OR2_X1 U6755 ( .A1(n5657), .A2(n5656), .ZN(n5658) );
  AND2_X1 U6756 ( .A1(n5659), .A2(n5658), .ZN(n6531) );
  INV_X1 U6757 ( .A(n6531), .ZN(n7445) );
  NAND2_X1 U6758 ( .A1(n5660), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n5666) );
  INV_X1 U6759 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5661) );
  NAND2_X1 U6760 ( .A1(n5662), .A2(n5661), .ZN(n5663) );
  NAND2_X1 U6761 ( .A1(n5663), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5664) );
  XNOR2_X1 U6762 ( .A(n5664), .B(P1_IR_REG_3__SCAN_IN), .ZN(n9848) );
  NAND2_X1 U6763 ( .A1(n5645), .A2(n9848), .ZN(n5665) );
  NAND2_X1 U6764 ( .A1(n6982), .A2(n5667), .ZN(n7945) );
  NAND2_X1 U6765 ( .A1(n7982), .A2(n7981), .ZN(n5669) );
  NAND2_X1 U6766 ( .A1(n6982), .A2(n10593), .ZN(n5668) );
  NAND2_X1 U6767 ( .A1(n5669), .A2(n5668), .ZN(n7989) );
  NAND2_X1 U6768 ( .A1(n5796), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5674) );
  NOR2_X1 U6769 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n5670) );
  NOR2_X1 U6770 ( .A1(n5685), .A2(n5670), .ZN(n8015) );
  NAND2_X1 U6771 ( .A1(n6171), .A2(n8015), .ZN(n5673) );
  NAND2_X1 U6772 ( .A1(n5686), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n5672) );
  NAND2_X1 U6773 ( .A1(n6222), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5671) );
  OR2_X1 U6774 ( .A1(n5676), .A2(n5675), .ZN(n5677) );
  NAND2_X1 U6775 ( .A1(n5678), .A2(n5677), .ZN(n7443) );
  NAND2_X1 U6776 ( .A1(n5660), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n5682) );
  NAND2_X1 U6777 ( .A1(n5679), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5680) );
  XNOR2_X1 U6778 ( .A(n5680), .B(P1_IR_REG_4__SCAN_IN), .ZN(n10527) );
  NAND2_X1 U6779 ( .A1(n5645), .A2(n10527), .ZN(n5681) );
  NOR2_X1 U6780 ( .A1(n6987), .A2(n8022), .ZN(n5684) );
  NAND2_X1 U6781 ( .A1(n6987), .A2(n8022), .ZN(n5683) );
  OAI21_X2 U6782 ( .B1(n7989), .B2(n5684), .A(n5683), .ZN(n7944) );
  NAND2_X1 U6783 ( .A1(n6222), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n5690) );
  NAND2_X1 U6784 ( .A1(n5796), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5689) );
  OAI21_X1 U6785 ( .B1(n5685), .B2(P1_REG3_REG_5__SCAN_IN), .A(n5703), .ZN(
        n10607) );
  INV_X1 U6786 ( .A(n10607), .ZN(n7925) );
  NAND2_X1 U6787 ( .A1(n6171), .A2(n7925), .ZN(n5688) );
  NAND2_X1 U6788 ( .A1(n5686), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n5687) );
  OR2_X1 U6789 ( .A1(n5692), .A2(n5691), .ZN(n5693) );
  NAND2_X1 U6790 ( .A1(n5694), .A2(n5693), .ZN(n7447) );
  NAND2_X1 U6791 ( .A1(n5660), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n5701) );
  NAND2_X1 U6792 ( .A1(n5695), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5696) );
  MUX2_X1 U6793 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5696), .S(
        P1_IR_REG_5__SCAN_IN), .Z(n5699) );
  INV_X1 U6794 ( .A(n5697), .ZN(n5698) );
  NAND2_X1 U6795 ( .A1(n5645), .A2(n7643), .ZN(n5700) );
  NAND2_X1 U6796 ( .A1(n8030), .A2(n7928), .ZN(n6253) );
  NAND2_X1 U6797 ( .A1(n5796), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n5708) );
  NAND2_X1 U6798 ( .A1(n6221), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n5707) );
  AND2_X1 U6799 ( .A1(n5703), .A2(n5702), .ZN(n5704) );
  NOR2_X1 U6800 ( .A1(n5716), .A2(n5704), .ZN(n8053) );
  NAND2_X1 U6801 ( .A1(n6171), .A2(n8053), .ZN(n5706) );
  NAND2_X1 U6802 ( .A1(n6222), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5705) );
  OR2_X1 U6803 ( .A1(n5710), .A2(n5709), .ZN(n5711) );
  NAND2_X1 U6804 ( .A1(n5712), .A2(n5711), .ZN(n7449) );
  NAND2_X1 U6805 ( .A1(n5660), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n5715) );
  OR2_X1 U6806 ( .A1(n5697), .A2(n5590), .ZN(n5713) );
  XNOR2_X1 U6807 ( .A(n5713), .B(P1_IR_REG_6__SCAN_IN), .ZN(n7619) );
  NAND2_X1 U6808 ( .A1(n5645), .A2(n7619), .ZN(n5714) );
  OAI211_X1 U6809 ( .C1(n7449), .C2(n6018), .A(n5715), .B(n5714), .ZN(n8038)
         );
  NAND2_X1 U6810 ( .A1(n8136), .A2(n8038), .ZN(n8073) );
  INV_X1 U6811 ( .A(n8038), .ZN(n10623) );
  NAND2_X1 U6812 ( .A1(n9807), .A2(n10623), .ZN(n8071) );
  NAND2_X1 U6813 ( .A1(n8073), .A2(n8071), .ZN(n8027) );
  NAND2_X1 U6814 ( .A1(n8026), .A2(n8027), .ZN(n8025) );
  NAND2_X1 U6815 ( .A1(n8025), .A2(n5514), .ZN(n8135) );
  INV_X2 U6816 ( .A(n5920), .ZN(n6220) );
  NAND2_X1 U6817 ( .A1(n6220), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n5721) );
  NAND2_X1 U6818 ( .A1(n6221), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n5720) );
  OR2_X1 U6819 ( .A1(n5716), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5717) );
  AND2_X1 U6820 ( .A1(n5738), .A2(n5717), .ZN(n8151) );
  NAND2_X1 U6821 ( .A1(n6171), .A2(n8151), .ZN(n5719) );
  NAND2_X1 U6822 ( .A1(n6222), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5718) );
  OR2_X1 U6823 ( .A1(n5723), .A2(n5722), .ZN(n5724) );
  NAND2_X1 U6824 ( .A1(n5725), .A2(n5724), .ZN(n7453) );
  OR2_X1 U6825 ( .A1(n7453), .A2(n6018), .ZN(n5729) );
  OR2_X1 U6826 ( .A1(n5726), .A2(n5590), .ZN(n5727) );
  XNOR2_X1 U6827 ( .A(n5727), .B(P1_IR_REG_7__SCAN_IN), .ZN(n7607) );
  AOI22_X1 U6828 ( .A1(n5660), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n7607), .B2(
        n5645), .ZN(n5728) );
  NAND2_X1 U6829 ( .A1(n5729), .A2(n5728), .ZN(n8271) );
  NAND2_X1 U6830 ( .A1(n8029), .A2(n8271), .ZN(n6261) );
  INV_X1 U6831 ( .A(n8271), .ZN(n8153) );
  NAND2_X1 U6832 ( .A1(n8153), .A2(n9806), .ZN(n6262) );
  NAND2_X1 U6833 ( .A1(n6261), .A2(n6262), .ZN(n8137) );
  NAND2_X1 U6834 ( .A1(n8029), .A2(n8153), .ZN(n5730) );
  XNOR2_X1 U6835 ( .A(n5732), .B(n5731), .ZN(n7454) );
  NAND2_X1 U6836 ( .A1(n7454), .A2(n6217), .ZN(n5736) );
  NAND2_X1 U6837 ( .A1(n5733), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5734) );
  XNOR2_X1 U6838 ( .A(n5734), .B(P1_IR_REG_8__SCAN_IN), .ZN(n7631) );
  AOI22_X1 U6839 ( .A1(n5660), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n7631), .B2(
        n5645), .ZN(n5735) );
  NAND2_X1 U6840 ( .A1(n5736), .A2(n5735), .ZN(n8167) );
  NAND2_X1 U6841 ( .A1(n6220), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5743) );
  NAND2_X1 U6842 ( .A1(n6222), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n5742) );
  NAND2_X1 U6843 ( .A1(n5738), .A2(n5737), .ZN(n5739) );
  AND2_X1 U6844 ( .A1(n5751), .A2(n5739), .ZN(n8163) );
  NAND2_X1 U6845 ( .A1(n6171), .A2(n8163), .ZN(n5741) );
  NAND2_X1 U6846 ( .A1(n6221), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n5740) );
  NAND2_X1 U6847 ( .A1(n8167), .A2(n8176), .ZN(n6078) );
  NAND2_X1 U6848 ( .A1(n8173), .A2(n6078), .ZN(n8080) );
  XNOR2_X2 U6849 ( .A(n5746), .B(n5745), .ZN(n8623) );
  NAND2_X1 U6850 ( .A1(n8623), .A2(n6217), .ZN(n5749) );
  NAND2_X1 U6851 ( .A1(n5747), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5762) );
  XNOR2_X1 U6852 ( .A(n5762), .B(P1_IR_REG_9__SCAN_IN), .ZN(n8621) );
  AOI22_X1 U6853 ( .A1(n5660), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n8621), .B2(
        n5645), .ZN(n5748) );
  NAND2_X2 U6854 ( .A1(n5749), .A2(n5748), .ZN(n5757) );
  NAND2_X1 U6855 ( .A1(n6222), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5756) );
  NAND2_X1 U6856 ( .A1(n6220), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n5755) );
  AND2_X1 U6857 ( .A1(n5751), .A2(n5750), .ZN(n5752) );
  NOR2_X1 U6858 ( .A1(n5766), .A2(n5752), .ZN(n8287) );
  NAND2_X1 U6859 ( .A1(n6171), .A2(n8287), .ZN(n5754) );
  NAND2_X1 U6860 ( .A1(n6221), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n5753) );
  NAND2_X1 U6861 ( .A1(n5757), .A2(n8246), .ZN(n6241) );
  NAND2_X1 U6862 ( .A1(n6239), .A2(n6241), .ZN(n8179) );
  NAND2_X1 U6863 ( .A1(n8180), .A2(n8179), .ZN(n8178) );
  NAND2_X1 U6864 ( .A1(n8178), .A2(n5758), .ZN(n8251) );
  NAND2_X1 U6865 ( .A1(n4995), .A2(n5759), .ZN(n5760) );
  NAND2_X1 U6866 ( .A1(n5761), .A2(n5760), .ZN(n7465) );
  INV_X1 U6867 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n7464) );
  NAND2_X1 U6868 ( .A1(n5762), .A2(n5867), .ZN(n5763) );
  NAND2_X1 U6869 ( .A1(n5763), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5775) );
  XNOR2_X1 U6870 ( .A(n5775), .B(P1_IR_REG_10__SCAN_IN), .ZN(n7662) );
  INV_X1 U6871 ( .A(n7662), .ZN(n7466) );
  OAI22_X1 U6872 ( .A1(n5902), .A2(n7464), .B1(n5618), .B2(n7466), .ZN(n5764)
         );
  INV_X1 U6873 ( .A(n5764), .ZN(n5765) );
  NAND2_X1 U6874 ( .A1(n6222), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5771) );
  NAND2_X1 U6875 ( .A1(n5796), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n5770) );
  NOR2_X1 U6876 ( .A1(n5766), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n5767) );
  OR2_X1 U6877 ( .A1(n5780), .A2(n5767), .ZN(n8252) );
  INV_X1 U6878 ( .A(n8252), .ZN(n8339) );
  NAND2_X1 U6879 ( .A1(n6171), .A2(n8339), .ZN(n5769) );
  NAND2_X1 U6880 ( .A1(n6221), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n5768) );
  NAND2_X1 U6881 ( .A1(n4944), .A2(n8290), .ZN(n6266) );
  NAND2_X1 U6882 ( .A1(n6401), .A2(n6266), .ZN(n8250) );
  NAND2_X1 U6883 ( .A1(n8251), .A2(n8250), .ZN(n8249) );
  NAND2_X1 U6884 ( .A1(n8249), .A2(n5772), .ZN(n8322) );
  XNOR2_X1 U6885 ( .A(n5774), .B(n5773), .ZN(n7480) );
  NAND2_X1 U6886 ( .A1(n7480), .A2(n6217), .ZN(n5779) );
  NAND2_X1 U6887 ( .A1(n5775), .A2(n5866), .ZN(n5776) );
  NAND2_X1 U6888 ( .A1(n5776), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5777) );
  XNOR2_X1 U6889 ( .A(n5777), .B(P1_IR_REG_11__SCAN_IN), .ZN(n7752) );
  AOI22_X1 U6890 ( .A1(n5660), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n7752), .B2(
        n5645), .ZN(n5778) );
  NAND2_X1 U6891 ( .A1(n5796), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n5785) );
  NAND2_X1 U6892 ( .A1(n6222), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5784) );
  OR2_X1 U6893 ( .A1(n5780), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n5781) );
  AND2_X1 U6894 ( .A1(n5797), .A2(n5781), .ZN(n8760) );
  NAND2_X1 U6895 ( .A1(n6171), .A2(n8760), .ZN(n5783) );
  NAND2_X1 U6896 ( .A1(n6221), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n5782) );
  OR2_X1 U6897 ( .A1(n8771), .A2(n8706), .ZN(n6273) );
  NAND2_X1 U6898 ( .A1(n8771), .A2(n8706), .ZN(n6240) );
  NAND2_X1 U6899 ( .A1(n6273), .A2(n6240), .ZN(n8323) );
  NAND2_X1 U6900 ( .A1(n8322), .A2(n8323), .ZN(n8321) );
  INV_X1 U6901 ( .A(n8706), .ZN(n9804) );
  NAND2_X1 U6902 ( .A1(n8321), .A2(n5786), .ZN(n8659) );
  NAND2_X1 U6903 ( .A1(n5788), .A2(n5787), .ZN(n5790) );
  NAND2_X1 U6904 ( .A1(n5790), .A2(n5789), .ZN(n7487) );
  OR2_X1 U6905 ( .A1(n7487), .A2(n6018), .ZN(n5795) );
  INV_X1 U6906 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n7486) );
  OR2_X1 U6907 ( .A1(n5010), .A2(n5590), .ZN(n5791) );
  MUX2_X1 U6908 ( .A(n5791), .B(P1_IR_REG_31__SCAN_IN), .S(n5870), .Z(n5792)
         );
  AND2_X1 U6909 ( .A1(n5792), .A2(n4949), .ZN(n7414) );
  INV_X1 U6910 ( .A(n7414), .ZN(n7806) );
  OAI22_X1 U6911 ( .A1(n5902), .A2(n7486), .B1(n5618), .B2(n7806), .ZN(n5793)
         );
  INV_X1 U6912 ( .A(n5793), .ZN(n5794) );
  NAND2_X1 U6913 ( .A1(n5796), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n5802) );
  NAND2_X1 U6914 ( .A1(n5797), .A2(n7803), .ZN(n5798) );
  AND2_X1 U6915 ( .A1(n5813), .A2(n5798), .ZN(n8705) );
  NAND2_X1 U6916 ( .A1(n6171), .A2(n8705), .ZN(n5801) );
  NAND2_X1 U6917 ( .A1(n6221), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n5800) );
  NAND2_X1 U6918 ( .A1(n6222), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5799) );
  NAND4_X1 U6919 ( .A1(n5802), .A2(n5801), .A3(n5800), .A4(n5799), .ZN(n9803)
         );
  NAND2_X1 U6920 ( .A1(n8665), .A2(n9803), .ZN(n5803) );
  INV_X1 U6921 ( .A(n9803), .ZN(n8763) );
  AOI22_X1 U6922 ( .A1(n8659), .A2(n5803), .B1(n10662), .B2(n8763), .ZN(n8682)
         );
  OR2_X1 U6923 ( .A1(n5805), .A2(n5804), .ZN(n5806) );
  NAND2_X1 U6924 ( .A1(n5807), .A2(n5806), .ZN(n7650) );
  OR2_X1 U6925 ( .A1(n7650), .A2(n6018), .ZN(n5811) );
  NAND2_X1 U6926 ( .A1(n4949), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5808) );
  MUX2_X1 U6927 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5808), .S(
        P1_IR_REG_13__SCAN_IN), .Z(n5809) );
  AOI22_X1 U6928 ( .A1(n5660), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n8108), .B2(
        n5645), .ZN(n5810) );
  NAND2_X1 U6929 ( .A1(n6220), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n5819) );
  NAND2_X1 U6930 ( .A1(n5813), .A2(n5812), .ZN(n5814) );
  AND2_X1 U6931 ( .A1(n5815), .A2(n5814), .ZN(n8739) );
  NAND2_X1 U6932 ( .A1(n6171), .A2(n8739), .ZN(n5818) );
  NAND2_X1 U6933 ( .A1(n6222), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n5817) );
  NAND2_X1 U6934 ( .A1(n6221), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n5816) );
  NAND4_X1 U6935 ( .A1(n5819), .A2(n5818), .A3(n5817), .A4(n5816), .ZN(n9802)
         );
  NAND2_X1 U6936 ( .A1(n5821), .A2(n5820), .ZN(n5822) );
  NAND2_X1 U6937 ( .A1(n8682), .A2(n5822), .ZN(n5824) );
  NAND2_X1 U6938 ( .A1(n10235), .A2(n9802), .ZN(n5823) );
  INV_X1 U6939 ( .A(n10230), .ZN(n8805) );
  INV_X1 U6940 ( .A(n9801), .ZN(n8832) );
  NAND2_X1 U6941 ( .A1(n8805), .A2(n8832), .ZN(n5825) );
  MUX2_X1 U6942 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .S(n7435), .Z(n5829) );
  NAND2_X1 U6943 ( .A1(n5829), .A2(SI_15_), .ZN(n5848) );
  OAI21_X1 U6944 ( .B1(n5829), .B2(SI_15_), .A(n5848), .ZN(n5830) );
  NAND2_X1 U6945 ( .A1(n5831), .A2(n5830), .ZN(n5832) );
  NAND2_X1 U6946 ( .A1(n5832), .A2(n5849), .ZN(n7704) );
  OR2_X1 U6947 ( .A1(n7704), .A2(n6018), .ZN(n5839) );
  INV_X1 U6948 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n7703) );
  NAND2_X1 U6949 ( .A1(n5834), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5836) );
  INV_X1 U6950 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n5835) );
  NAND2_X1 U6951 ( .A1(n5836), .A2(n5835), .ZN(n5850) );
  OAI21_X1 U6952 ( .B1(n5836), .B2(n5835), .A(n5850), .ZN(n9864) );
  OAI22_X1 U6953 ( .A1(n5902), .A2(n7703), .B1(n5618), .B2(n9864), .ZN(n5837)
         );
  INV_X1 U6954 ( .A(n5837), .ZN(n5838) );
  NAND2_X1 U6955 ( .A1(n6220), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n5845) );
  NAND2_X1 U6956 ( .A1(n5840), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n5855) );
  OR2_X1 U6957 ( .A1(n5840), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n5841) );
  AND2_X1 U6958 ( .A1(n5855), .A2(n5841), .ZN(n8829) );
  NAND2_X1 U6959 ( .A1(n6171), .A2(n8829), .ZN(n5844) );
  NAND2_X1 U6960 ( .A1(n6222), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n5843) );
  NAND2_X1 U6961 ( .A1(n6221), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n5842) );
  NAND4_X1 U6962 ( .A1(n5845), .A2(n5844), .A3(n5843), .A4(n5842), .ZN(n9800)
         );
  INV_X1 U6963 ( .A(n10225), .ZN(n8790) );
  INV_X1 U6964 ( .A(n9800), .ZN(n10142) );
  NAND2_X1 U6965 ( .A1(n10225), .A2(n9800), .ZN(n5846) );
  NAND2_X2 U6966 ( .A1(n5847), .A2(n5846), .ZN(n10138) );
  MUX2_X1 U6967 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(P2_DATAO_REG_16__SCAN_IN), 
        .S(n7435), .Z(n5860) );
  XNOR2_X1 U6968 ( .A(n5860), .B(SI_16_), .ZN(n5863) );
  XNOR2_X1 U6969 ( .A(n5864), .B(n5863), .ZN(n7758) );
  NAND2_X1 U6970 ( .A1(n7758), .A2(n6217), .ZN(n5853) );
  NAND2_X1 U6971 ( .A1(n5850), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5851) );
  XNOR2_X1 U6972 ( .A(n5851), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9881) );
  AOI22_X1 U6973 ( .A1(n5660), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n9881), .B2(
        n5645), .ZN(n5852) );
  NAND2_X1 U6974 ( .A1(n6222), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n5859) );
  NAND2_X1 U6975 ( .A1(n6220), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n5858) );
  INV_X1 U6976 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n5854) );
  AOI21_X1 U6977 ( .B1(n5855), .B2(n5854), .A(n5880), .ZN(n10148) );
  NAND2_X1 U6978 ( .A1(n6171), .A2(n10148), .ZN(n5857) );
  NAND2_X1 U6979 ( .A1(n6221), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n5856) );
  NAND2_X1 U6980 ( .A1(n10222), .A2(n10125), .ZN(n6413) );
  NAND2_X1 U6981 ( .A1(n6297), .A2(n6413), .ZN(n10137) );
  INV_X1 U6982 ( .A(n5860), .ZN(n5861) );
  NAND2_X1 U6983 ( .A1(n5861), .A2(n8535), .ZN(n5862) );
  MUX2_X1 U6984 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(P2_DATAO_REG_17__SCAN_IN), 
        .S(n7435), .Z(n5886) );
  XNOR2_X1 U6985 ( .A(n5888), .B(n5887), .ZN(n7885) );
  NAND2_X1 U6986 ( .A1(n7885), .A2(n6217), .ZN(n5879) );
  INV_X1 U6987 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n7917) );
  NAND4_X1 U6988 ( .A1(n5868), .A2(n5572), .A3(n5867), .A4(n5866), .ZN(n5873)
         );
  NAND3_X1 U6989 ( .A1(n5871), .A2(n5870), .A3(n5869), .ZN(n5872) );
  NAND2_X1 U6990 ( .A1(n5897), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5876) );
  XNOR2_X1 U6991 ( .A(n5876), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9898) );
  INV_X1 U6992 ( .A(n9898), .ZN(n9886) );
  OAI22_X1 U6993 ( .A1(n5902), .A2(n7917), .B1(n5618), .B2(n9886), .ZN(n5877)
         );
  INV_X1 U6994 ( .A(n5877), .ZN(n5878) );
  NAND2_X1 U6995 ( .A1(n5634), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n5885) );
  NAND2_X1 U6996 ( .A1(n6221), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n5884) );
  NAND2_X1 U6997 ( .A1(n5880), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n5907) );
  OAI21_X1 U6998 ( .B1(n5880), .B2(P1_REG3_REG_17__SCAN_IN), .A(n5907), .ZN(
        n5881) );
  INV_X1 U6999 ( .A(n5881), .ZN(n10130) );
  NAND2_X1 U7000 ( .A1(n6171), .A2(n10130), .ZN(n5883) );
  NAND2_X1 U7001 ( .A1(n6220), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n5882) );
  NAND2_X1 U7002 ( .A1(n10131), .A2(n10144), .ZN(n6417) );
  MUX2_X1 U7003 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n7435), .Z(n5889) );
  NAND2_X1 U7004 ( .A1(n5889), .A2(SI_18_), .ZN(n5912) );
  INV_X1 U7005 ( .A(n5889), .ZN(n5890) );
  NAND2_X1 U7006 ( .A1(n5890), .A2(n8432), .ZN(n5891) );
  NAND2_X1 U7007 ( .A1(n5912), .A2(n5891), .ZN(n5894) );
  INV_X1 U7008 ( .A(n5894), .ZN(n5892) );
  NAND2_X1 U7009 ( .A1(n5893), .A2(n5892), .ZN(n5913) );
  INV_X1 U7010 ( .A(n5893), .ZN(n5895) );
  NAND2_X1 U7011 ( .A1(n5895), .A2(n5894), .ZN(n5896) );
  NAND2_X1 U7012 ( .A1(n5913), .A2(n5896), .ZN(n7919) );
  OR2_X1 U7013 ( .A1(n7919), .A2(n6018), .ZN(n5905) );
  INV_X1 U7014 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n7896) );
  INV_X1 U7015 ( .A(n5900), .ZN(n5898) );
  NAND2_X1 U7016 ( .A1(n5898), .A2(P1_IR_REG_18__SCAN_IN), .ZN(n5901) );
  NAND2_X1 U7017 ( .A1(n5901), .A2(n5914), .ZN(n9893) );
  OAI22_X1 U7018 ( .A1(n5902), .A2(n7896), .B1(n5618), .B2(n9893), .ZN(n5903)
         );
  INV_X1 U7019 ( .A(n5903), .ZN(n5904) );
  INV_X1 U7020 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n5906) );
  AOI21_X1 U7021 ( .B1(n5907), .B2(n5906), .A(n5921), .ZN(n10114) );
  NAND2_X1 U7022 ( .A1(n6171), .A2(n10114), .ZN(n5911) );
  NAND2_X1 U7023 ( .A1(n6220), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n5910) );
  NAND2_X1 U7024 ( .A1(n6222), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n5909) );
  NAND2_X1 U7025 ( .A1(n6221), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n5908) );
  NAND2_X1 U7026 ( .A1(n10210), .A2(n10124), .ZN(n6416) );
  NAND2_X1 U7027 ( .A1(n6421), .A2(n6416), .ZN(n10106) );
  NAND2_X1 U7028 ( .A1(n5913), .A2(n5912), .ZN(n5930) );
  MUX2_X1 U7029 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(P2_DATAO_REG_19__SCAN_IN), 
        .S(n7435), .Z(n5926) );
  XNOR2_X1 U7030 ( .A(n5926), .B(SI_19_), .ZN(n5929) );
  XNOR2_X1 U7031 ( .A(n5930), .B(n5929), .ZN(n8088) );
  NAND2_X1 U7032 ( .A1(n8088), .A2(n6217), .ZN(n5917) );
  AOI22_X1 U7033 ( .A1(n5660), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n9923), .B2(
        n5645), .ZN(n5916) );
  INV_X1 U7034 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n10206) );
  NAND2_X1 U7035 ( .A1(n6222), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n5919) );
  NAND2_X1 U7036 ( .A1(n6221), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n5918) );
  OAI211_X1 U7037 ( .C1(n5920), .C2(n10206), .A(n5919), .B(n5918), .ZN(n5925)
         );
  OR2_X1 U7038 ( .A1(n5921), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n5922) );
  NAND2_X1 U7039 ( .A1(n5921), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n5933) );
  NAND2_X1 U7040 ( .A1(n5922), .A2(n5933), .ZN(n10099) );
  INV_X1 U7041 ( .A(n6171), .ZN(n5923) );
  NOR2_X1 U7042 ( .A1(n10099), .A2(n5923), .ZN(n5924) );
  OR2_X1 U7043 ( .A1(n10102), .A2(n10111), .ZN(n6422) );
  NAND2_X1 U7044 ( .A1(n10102), .A2(n10111), .ZN(n6423) );
  INV_X1 U7045 ( .A(n5926), .ZN(n5927) );
  NAND2_X1 U7046 ( .A1(n5927), .A2(n8511), .ZN(n5928) );
  MUX2_X1 U7047 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(P2_DATAO_REG_20__SCAN_IN), 
        .S(n7435), .Z(n5942) );
  XNOR2_X1 U7048 ( .A(n5942), .B(n8512), .ZN(n5940) );
  XNOR2_X1 U7049 ( .A(n5941), .B(n5940), .ZN(n8170) );
  NAND2_X1 U7050 ( .A1(n8170), .A2(n6217), .ZN(n5932) );
  NAND2_X1 U7051 ( .A1(n5660), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n5931) );
  NAND2_X1 U7052 ( .A1(n6222), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n5939) );
  NAND2_X1 U7053 ( .A1(n6220), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n5938) );
  INV_X1 U7054 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n9740) );
  NAND2_X1 U7055 ( .A1(n9740), .A2(n5933), .ZN(n5935) );
  INV_X1 U7056 ( .A(n5933), .ZN(n5934) );
  NAND2_X1 U7057 ( .A1(P1_REG3_REG_20__SCAN_IN), .A2(n5934), .ZN(n5952) );
  AND2_X1 U7058 ( .A1(n5935), .A2(n5952), .ZN(n10084) );
  NAND2_X1 U7059 ( .A1(n6171), .A2(n10084), .ZN(n5937) );
  NAND2_X1 U7060 ( .A1(n6221), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n5936) );
  NAND2_X1 U7061 ( .A1(n10200), .A2(n10097), .ZN(n10060) );
  INV_X1 U7062 ( .A(n10097), .ZN(n9698) );
  OAI22_X1 U7063 ( .A1(n10077), .A2(n10078), .B1(n9698), .B2(n10200), .ZN(
        n10058) );
  INV_X1 U7064 ( .A(n5942), .ZN(n5943) );
  NAND2_X1 U7065 ( .A1(n5943), .A2(n8512), .ZN(n5944) );
  MUX2_X1 U7066 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(P2_DATAO_REG_21__SCAN_IN), 
        .S(n7435), .Z(n5945) );
  NAND2_X1 U7067 ( .A1(n5945), .A2(SI_21_), .ZN(n5960) );
  INV_X1 U7068 ( .A(n5945), .ZN(n5946) );
  INV_X1 U7069 ( .A(SI_21_), .ZN(n8531) );
  NAND2_X1 U7070 ( .A1(n5946), .A2(n8531), .ZN(n5947) );
  XNOR2_X1 U7071 ( .A(n5958), .B(n5959), .ZN(n8307) );
  NAND2_X1 U7072 ( .A1(n8307), .A2(n6217), .ZN(n5949) );
  NAND2_X1 U7073 ( .A1(n5660), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n5948) );
  NAND2_X1 U7074 ( .A1(n6222), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n5957) );
  NAND2_X1 U7075 ( .A1(n6220), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n5956) );
  INV_X1 U7076 ( .A(n5952), .ZN(n5950) );
  NAND2_X1 U7077 ( .A1(n5950), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n5971) );
  INV_X1 U7078 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n5951) );
  NAND2_X1 U7079 ( .A1(n5952), .A2(n5951), .ZN(n5953) );
  AND2_X1 U7080 ( .A1(n5971), .A2(n5953), .ZN(n10071) );
  NAND2_X1 U7081 ( .A1(n6171), .A2(n10071), .ZN(n5955) );
  NAND2_X1 U7082 ( .A1(n6221), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n5954) );
  NAND2_X1 U7083 ( .A1(n10070), .A2(n10081), .ZN(n6313) );
  INV_X1 U7084 ( .A(n10081), .ZN(n10048) );
  NAND2_X1 U7085 ( .A1(n5961), .A2(n5960), .ZN(n5966) );
  MUX2_X1 U7086 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(P2_DATAO_REG_22__SCAN_IN), 
        .S(n7435), .Z(n5962) );
  NAND2_X1 U7087 ( .A1(n5962), .A2(SI_22_), .ZN(n5978) );
  INV_X1 U7088 ( .A(n5962), .ZN(n5963) );
  NAND2_X1 U7089 ( .A1(n5963), .A2(n8527), .ZN(n5964) );
  NAND2_X1 U7090 ( .A1(n5966), .A2(n5965), .ZN(n5979) );
  OR2_X1 U7091 ( .A1(n5966), .A2(n5965), .ZN(n5967) );
  NAND2_X1 U7092 ( .A1(n5979), .A2(n5967), .ZN(n8357) );
  OR2_X1 U7093 ( .A1(n8357), .A2(n6018), .ZN(n5969) );
  NAND2_X1 U7094 ( .A1(n5660), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n5968) );
  NAND2_X1 U7095 ( .A1(n6220), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n5976) );
  NAND2_X1 U7096 ( .A1(n6221), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n5975) );
  INV_X1 U7097 ( .A(n5971), .ZN(n5970) );
  NAND2_X1 U7098 ( .A1(n5970), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n5983) );
  INV_X1 U7099 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n9752) );
  NAND2_X1 U7100 ( .A1(n5971), .A2(n9752), .ZN(n5972) );
  AND2_X1 U7101 ( .A1(n5983), .A2(n5972), .ZN(n10053) );
  NAND2_X1 U7102 ( .A1(n6171), .A2(n10053), .ZN(n5974) );
  NAND2_X1 U7103 ( .A1(n6222), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n5973) );
  NAND2_X1 U7104 ( .A1(n10190), .A2(n10065), .ZN(n6229) );
  NAND2_X1 U7105 ( .A1(n6230), .A2(n6229), .ZN(n10041) );
  INV_X1 U7106 ( .A(n10190), .ZN(n5977) );
  NAND2_X1 U7107 ( .A1(n5979), .A2(n5978), .ZN(n5995) );
  MUX2_X1 U7108 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(P2_DATAO_REG_23__SCAN_IN), 
        .S(n7435), .Z(n5990) );
  XNOR2_X1 U7109 ( .A(n5990), .B(SI_23_), .ZN(n5994) );
  XNOR2_X1 U7110 ( .A(n5995), .B(n5994), .ZN(n8378) );
  NAND2_X1 U7111 ( .A1(n8378), .A2(n6217), .ZN(n5981) );
  NAND2_X1 U7112 ( .A1(n5660), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n5980) );
  NAND2_X1 U7113 ( .A1(n6220), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n5988) );
  INV_X1 U7114 ( .A(n5983), .ZN(n5982) );
  NAND2_X1 U7115 ( .A1(n5982), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n5999) );
  INV_X1 U7116 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n9680) );
  NAND2_X1 U7117 ( .A1(n5983), .A2(n9680), .ZN(n5984) );
  AND2_X1 U7118 ( .A1(n5999), .A2(n5984), .ZN(n10034) );
  NAND2_X1 U7119 ( .A1(n6171), .A2(n10034), .ZN(n5987) );
  NAND2_X1 U7120 ( .A1(n5634), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n5986) );
  NAND2_X1 U7121 ( .A1(n6221), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n5985) );
  NAND4_X1 U7122 ( .A1(n5988), .A2(n5987), .A3(n5986), .A4(n5985), .ZN(n10047)
         );
  NOR2_X1 U7123 ( .A1(n6101), .A2(n10047), .ZN(n5989) );
  INV_X1 U7124 ( .A(n6101), .ZN(n10037) );
  OAI22_X1 U7125 ( .A1(n10025), .A2(n5989), .B1(n9753), .B2(n10037), .ZN(
        n10011) );
  INV_X1 U7126 ( .A(n5990), .ZN(n5992) );
  INV_X1 U7127 ( .A(SI_23_), .ZN(n5991) );
  NAND2_X1 U7128 ( .A1(n5992), .A2(n5991), .ZN(n5993) );
  OAI21_X2 U7129 ( .B1(n5995), .B2(n5994), .A(n5993), .ZN(n6008) );
  MUX2_X1 U7130 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(P2_DATAO_REG_24__SCAN_IN), 
        .S(n7435), .Z(n6009) );
  XNOR2_X1 U7131 ( .A(n6009), .B(n6010), .ZN(n6007) );
  XNOR2_X1 U7132 ( .A(n6008), .B(n6007), .ZN(n8731) );
  NAND2_X1 U7133 ( .A1(n8731), .A2(n6217), .ZN(n5997) );
  NAND2_X1 U7134 ( .A1(n5660), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n5996) );
  NAND2_X1 U7135 ( .A1(n5634), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n6004) );
  NAND2_X1 U7136 ( .A1(n6220), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n6003) );
  INV_X1 U7137 ( .A(n5999), .ZN(n5998) );
  NAND2_X1 U7138 ( .A1(n5998), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n6023) );
  INV_X1 U7139 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n9731) );
  NAND2_X1 U7140 ( .A1(n5999), .A2(n9731), .ZN(n6000) );
  AND2_X1 U7141 ( .A1(n6023), .A2(n6000), .ZN(n10019) );
  NAND2_X1 U7142 ( .A1(n6171), .A2(n10019), .ZN(n6002) );
  NAND2_X1 U7143 ( .A1(n6221), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n6001) );
  OR2_X2 U7144 ( .A1(n10181), .A2(n10031), .ZN(n6354) );
  NAND2_X1 U7145 ( .A1(n10011), .A2(n10010), .ZN(n6006) );
  NAND2_X1 U7146 ( .A1(n10181), .A2(n9706), .ZN(n6005) );
  NAND2_X1 U7147 ( .A1(n6006), .A2(n6005), .ZN(n9991) );
  NAND2_X1 U7148 ( .A1(n6008), .A2(n6007), .ZN(n6013) );
  INV_X1 U7149 ( .A(n6009), .ZN(n6011) );
  NAND2_X1 U7150 ( .A1(n6011), .A2(n6010), .ZN(n6012) );
  MUX2_X1 U7151 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(P2_DATAO_REG_25__SCAN_IN), 
        .S(n7435), .Z(n6014) );
  NAND2_X1 U7152 ( .A1(n6014), .A2(SI_25_), .ZN(n6032) );
  OAI21_X1 U7153 ( .B1(n6014), .B2(SI_25_), .A(n6032), .ZN(n6015) );
  NAND2_X1 U7154 ( .A1(n6016), .A2(n6015), .ZN(n6017) );
  NAND2_X1 U7155 ( .A1(n6033), .A2(n6017), .ZN(n8785) );
  NAND2_X1 U7156 ( .A1(n5660), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n6019) );
  NAND2_X1 U7157 ( .A1(n6220), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n6028) );
  INV_X1 U7158 ( .A(n6023), .ZN(n6021) );
  NAND2_X1 U7159 ( .A1(n6021), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n6038) );
  INV_X1 U7160 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n6022) );
  NAND2_X1 U7161 ( .A1(n6023), .A2(n6022), .ZN(n6024) );
  AND2_X1 U7162 ( .A1(n6038), .A2(n6024), .ZN(n10003) );
  NAND2_X1 U7163 ( .A1(n6171), .A2(n10003), .ZN(n6027) );
  NAND2_X1 U7164 ( .A1(n6222), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n6026) );
  NAND2_X1 U7165 ( .A1(n6221), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n6025) );
  NAND4_X1 U7166 ( .A1(n6028), .A2(n6027), .A3(n6026), .A4(n6025), .ZN(n10015)
         );
  NAND2_X1 U7167 ( .A1(n9991), .A2(n6029), .ZN(n6031) );
  NAND2_X1 U7168 ( .A1(n10174), .A2(n10015), .ZN(n6030) );
  MUX2_X1 U7169 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(P2_DATAO_REG_26__SCAN_IN), 
        .S(n7435), .Z(n6045) );
  XNOR2_X1 U7170 ( .A(n6045), .B(SI_26_), .ZN(n6048) );
  XNOR2_X1 U7171 ( .A(n6049), .B(n6048), .ZN(n8798) );
  NAND2_X1 U7172 ( .A1(n8798), .A2(n6217), .ZN(n6035) );
  NAND2_X1 U7173 ( .A1(n5660), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n6034) );
  NAND2_X1 U7174 ( .A1(n6222), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n6043) );
  NAND2_X1 U7175 ( .A1(n6220), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n6042) );
  INV_X1 U7176 ( .A(n6038), .ZN(n6036) );
  NAND2_X1 U7177 ( .A1(n6036), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n6054) );
  INV_X1 U7178 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n6037) );
  NAND2_X1 U7179 ( .A1(n6038), .A2(n6037), .ZN(n6039) );
  NAND2_X1 U7180 ( .A1(n6171), .A2(n9977), .ZN(n6041) );
  NAND2_X1 U7181 ( .A1(n6221), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n6040) );
  NAND2_X1 U7182 ( .A1(n10249), .A2(n9996), .ZN(n6326) );
  NAND2_X1 U7183 ( .A1(n9974), .A2(n9980), .ZN(n6044) );
  NAND2_X1 U7184 ( .A1(n10249), .A2(n9797), .ZN(n7350) );
  NAND2_X1 U7185 ( .A1(n6044), .A2(n7350), .ZN(n6060) );
  INV_X1 U7186 ( .A(n6045), .ZN(n6046) );
  INV_X1 U7187 ( .A(SI_26_), .ZN(n8411) );
  NAND2_X1 U7188 ( .A1(n6046), .A2(n8411), .ZN(n6047) );
  MUX2_X1 U7189 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(P2_DATAO_REG_27__SCAN_IN), 
        .S(n7435), .Z(n6159) );
  XNOR2_X1 U7190 ( .A(n6159), .B(n8523), .ZN(n6157) );
  NAND2_X1 U7191 ( .A1(n9672), .A2(n6217), .ZN(n6051) );
  NAND2_X1 U7192 ( .A1(n5660), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n6050) );
  NAND2_X1 U7193 ( .A1(n5634), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n6059) );
  NAND2_X1 U7194 ( .A1(n6220), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n6058) );
  INV_X1 U7195 ( .A(n6054), .ZN(n6052) );
  NAND2_X1 U7196 ( .A1(n6052), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n6107) );
  INV_X1 U7197 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n6053) );
  NAND2_X1 U7198 ( .A1(n6054), .A2(n6053), .ZN(n6055) );
  NAND2_X1 U7199 ( .A1(n6171), .A2(n9966), .ZN(n6057) );
  NAND2_X1 U7200 ( .A1(n6221), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n6056) );
  NAND2_X1 U7201 ( .A1(n7329), .A2(n9984), .ZN(n6344) );
  XNOR2_X1 U7202 ( .A(n6060), .B(n5370), .ZN(n9973) );
  NOR2_X1 U7203 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), .ZN(
        n6061) );
  NAND2_X1 U7204 ( .A1(n6067), .A2(n6066), .ZN(n6068) );
  OAI21_X1 U7205 ( .B1(P1_IR_REG_21__SCAN_IN), .B2(P1_IR_REG_20__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n6064) );
  NAND2_X1 U7206 ( .A1(n8320), .A2(n6065), .ZN(n7654) );
  OR2_X1 U7207 ( .A1(n6067), .A2(n6066), .ZN(n6069) );
  NAND2_X1 U7208 ( .A1(n6949), .A2(n6948), .ZN(n6071) );
  AND2_X1 U7209 ( .A1(n7654), .A2(n6071), .ZN(n6073) );
  OR2_X1 U7210 ( .A1(n7854), .A2(n6949), .ZN(n6442) );
  NAND2_X1 U7211 ( .A1(n6073), .A2(n6442), .ZN(n8028) );
  INV_X1 U7212 ( .A(n10210), .ZN(n10117) );
  INV_X1 U7213 ( .A(n6971), .ZN(n10571) );
  INV_X1 U7214 ( .A(n8022), .ZN(n8115) );
  NAND2_X1 U7215 ( .A1(n7995), .A2(n10613), .ZN(n8034) );
  INV_X1 U7216 ( .A(n10174), .ZN(n10006) );
  NAND2_X1 U7217 ( .A1(n10018), .A2(n10006), .ZN(n9975) );
  NOR2_X2 U7218 ( .A1(n10249), .A2(n9975), .ZN(n6074) );
  INV_X1 U7219 ( .A(n6074), .ZN(n9976) );
  AOI21_X1 U7220 ( .B1(n7329), .B2(n9976), .A(n7367), .ZN(n9965) );
  OR2_X1 U7221 ( .A1(n6075), .A2(P1_IR_REG_27__SCAN_IN), .ZN(n6444) );
  NAND2_X1 U7222 ( .A1(n6444), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6077) );
  NAND2_X1 U7223 ( .A1(n6072), .A2(n6447), .ZN(n6372) );
  NAND2_X1 U7224 ( .A1(n6241), .A2(n6078), .ZN(n6265) );
  INV_X1 U7225 ( .A(n6261), .ZN(n8075) );
  OR2_X1 U7226 ( .A1(n6265), .A2(n8075), .ZN(n6183) );
  NAND2_X1 U7227 ( .A1(n6079), .A2(n6241), .ZN(n6080) );
  NAND2_X1 U7228 ( .A1(n6183), .A2(n6080), .ZN(n6081) );
  NAND2_X1 U7229 ( .A1(n6082), .A2(n6081), .ZN(n6402) );
  INV_X1 U7230 ( .A(n6402), .ZN(n6092) );
  NAND2_X1 U7231 ( .A1(n7864), .A2(n7863), .ZN(n7862) );
  NAND2_X1 U7232 ( .A1(n6083), .A2(n7861), .ZN(n6084) );
  AND2_X1 U7233 ( .A1(n7862), .A2(n6084), .ZN(n10556) );
  NAND2_X1 U7234 ( .A1(n6085), .A2(n10571), .ZN(n6086) );
  NAND2_X1 U7235 ( .A1(n10556), .A2(n6086), .ZN(n6392) );
  NAND2_X1 U7236 ( .A1(n6970), .A2(n6971), .ZN(n6389) );
  NAND2_X1 U7237 ( .A1(n6392), .A2(n6389), .ZN(n7974) );
  INV_X1 U7238 ( .A(n6390), .ZN(n6089) );
  OAI21_X1 U7239 ( .B1(n7974), .B2(n6089), .A(n6088), .ZN(n6090) );
  NAND2_X1 U7240 ( .A1(n6987), .A2(n8115), .ZN(n6394) );
  NAND2_X1 U7241 ( .A1(n6090), .A2(n6394), .ZN(n6250) );
  NAND2_X1 U7242 ( .A1(n6250), .A2(n7946), .ZN(n7954) );
  NAND2_X1 U7243 ( .A1(n7954), .A2(n6395), .ZN(n8074) );
  NAND2_X1 U7244 ( .A1(n6092), .A2(n6091), .ZN(n8245) );
  INV_X1 U7245 ( .A(n8250), .ZN(n8244) );
  NAND2_X1 U7246 ( .A1(n8245), .A2(n8244), .ZN(n6093) );
  NAND2_X1 U7247 ( .A1(n6093), .A2(n6266), .ZN(n8324) );
  INV_X1 U7248 ( .A(n8324), .ZN(n6095) );
  NAND2_X1 U7249 ( .A1(n6095), .A2(n6094), .ZN(n8326) );
  NAND2_X1 U7250 ( .A1(n8326), .A2(n6273), .ZN(n8662) );
  NAND2_X1 U7251 ( .A1(n8665), .A2(n8763), .ZN(n6277) );
  OR2_X1 U7252 ( .A1(n10235), .A2(n5820), .ZN(n6408) );
  NAND2_X1 U7253 ( .A1(n10235), .A2(n5820), .ZN(n6284) );
  OR2_X1 U7254 ( .A1(n10230), .A2(n8832), .ZN(n8791) );
  NAND2_X1 U7255 ( .A1(n10230), .A2(n8832), .ZN(n6279) );
  NAND2_X1 U7256 ( .A1(n8791), .A2(n6279), .ZN(n8809) );
  NAND2_X1 U7257 ( .A1(n8790), .A2(n9800), .ZN(n6296) );
  AND2_X1 U7258 ( .A1(n6296), .A2(n8791), .ZN(n6280) );
  AND2_X1 U7259 ( .A1(n10225), .A2(n10142), .ZN(n6288) );
  NAND2_X1 U7260 ( .A1(n6098), .A2(n6300), .ZN(n10109) );
  INV_X1 U7261 ( .A(n10106), .ZN(n10108) );
  NAND2_X1 U7262 ( .A1(n10109), .A2(n10108), .ZN(n6099) );
  NAND2_X1 U7263 ( .A1(n6099), .A2(n6421), .ZN(n10095) );
  INV_X1 U7264 ( .A(n10095), .ZN(n6100) );
  NAND2_X1 U7265 ( .A1(n6100), .A2(n6306), .ZN(n10093) );
  NAND2_X1 U7266 ( .A1(n6313), .A2(n10060), .ZN(n6309) );
  NAND2_X1 U7267 ( .A1(n6309), .A2(n6427), .ZN(n6346) );
  AND2_X2 U7268 ( .A1(n6345), .A2(n6346), .ZN(n10046) );
  INV_X1 U7269 ( .A(n10041), .ZN(n10045) );
  OR2_X1 U7270 ( .A1(n6101), .A2(n9753), .ZN(n6316) );
  NAND2_X1 U7271 ( .A1(n6101), .A2(n9753), .ZN(n6351) );
  NAND2_X1 U7272 ( .A1(n6316), .A2(n6351), .ZN(n10029) );
  INV_X1 U7273 ( .A(n10010), .ZN(n10013) );
  INV_X1 U7274 ( .A(n10015), .ZN(n9732) );
  NAND2_X1 U7275 ( .A1(n10174), .A2(n9732), .ZN(n6325) );
  NAND2_X1 U7276 ( .A1(n9992), .A2(n9993), .ZN(n9998) );
  NAND2_X1 U7277 ( .A1(n9998), .A2(n6358), .ZN(n9981) );
  NAND2_X1 U7278 ( .A1(n6072), .A2(n7184), .ZN(n6103) );
  NAND2_X1 U7279 ( .A1(n6447), .A2(n9923), .ZN(n6342) );
  OAI211_X1 U7280 ( .C1(n6194), .C2(n6104), .A(n7362), .B(n10127), .ZN(n6114)
         );
  NAND2_X1 U7281 ( .A1(n6222), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n6112) );
  NAND2_X1 U7282 ( .A1(n6220), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n6111) );
  INV_X1 U7283 ( .A(n6107), .ZN(n6105) );
  NAND2_X1 U7284 ( .A1(n6105), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n6170) );
  INV_X1 U7285 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n6106) );
  NAND2_X1 U7286 ( .A1(n6107), .A2(n6106), .ZN(n6108) );
  NAND2_X1 U7287 ( .A1(n6171), .A2(n9957), .ZN(n6110) );
  NAND2_X1 U7288 ( .A1(n6221), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n6109) );
  INV_X1 U7289 ( .A(n9942), .ZN(n9795) );
  NAND2_X1 U7290 ( .A1(n9795), .A2(n10558), .ZN(n6113) );
  OAI211_X1 U7291 ( .C1(n9996), .C2(n10143), .A(n6114), .B(n6113), .ZN(n9971)
         );
  NAND2_X1 U7292 ( .A1(n6116), .A2(n6119), .ZN(n6117) );
  NAND2_X1 U7293 ( .A1(n8759), .A2(P1_B_REG_SCAN_IN), .ZN(n6125) );
  BUF_X1 U7294 ( .A(n6120), .Z(n6121) );
  INV_X1 U7295 ( .A(n6121), .ZN(n6122) );
  NAND2_X1 U7296 ( .A1(n6122), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6124) );
  MUX2_X1 U7297 ( .A(P1_B_REG_SCAN_IN), .B(n6125), .S(n8733), .Z(n6126) );
  NAND2_X1 U7298 ( .A1(n8838), .A2(n8759), .ZN(n10275) );
  OAI21_X1 U7299 ( .B1(n10273), .B2(P1_D_REG_1__SCAN_IN), .A(n10275), .ZN(
        n7159) );
  NOR4_X1 U7300 ( .A1(P1_D_REG_27__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_25__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n6135) );
  NOR4_X1 U7301 ( .A1(P1_D_REG_23__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_21__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n6134) );
  NOR4_X1 U7302 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_13__SCAN_IN), .A4(P1_D_REG_12__SCAN_IN), .ZN(n6130) );
  NOR4_X1 U7303 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_18__SCAN_IN), .A4(P1_D_REG_16__SCAN_IN), .ZN(n6129) );
  NOR4_X1 U7304 ( .A1(P1_D_REG_7__SCAN_IN), .A2(P1_D_REG_6__SCAN_IN), .A3(
        P1_D_REG_5__SCAN_IN), .A4(P1_D_REG_2__SCAN_IN), .ZN(n6128) );
  NOR4_X1 U7305 ( .A1(P1_D_REG_11__SCAN_IN), .A2(P1_D_REG_10__SCAN_IN), .A3(
        P1_D_REG_9__SCAN_IN), .A4(P1_D_REG_8__SCAN_IN), .ZN(n6127) );
  NAND4_X1 U7306 ( .A1(n6130), .A2(n6129), .A3(n6128), .A4(n6127), .ZN(n6131)
         );
  NOR4_X1 U7307 ( .A1(P1_D_REG_4__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        n6132), .A4(n6131), .ZN(n6133) );
  NAND3_X1 U7308 ( .A1(n6135), .A2(n6134), .A3(n6133), .ZN(n6136) );
  NAND2_X1 U7309 ( .A1(n6138), .A2(n6136), .ZN(n7158) );
  INV_X1 U7310 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n6137) );
  NAND2_X1 U7311 ( .A1(n6138), .A2(n6137), .ZN(n6139) );
  NAND2_X1 U7312 ( .A1(n8838), .A2(n8733), .ZN(n10276) );
  NAND2_X1 U7313 ( .A1(n10274), .A2(n7187), .ZN(n6151) );
  NOR2_X1 U7314 ( .A1(n7161), .A2(n6151), .ZN(n6146) );
  MUX2_X1 U7315 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n6154), .S(n10646), .Z(n6147) );
  INV_X1 U7316 ( .A(n6147), .ZN(n6150) );
  INV_X1 U7317 ( .A(n7654), .ZN(n7822) );
  INV_X1 U7318 ( .A(n10219), .ZN(n6148) );
  NAND2_X1 U7319 ( .A1(n6150), .A2(n6149), .ZN(P1_U3549) );
  INV_X1 U7320 ( .A(n6151), .ZN(n6152) );
  NAND2_X1 U7321 ( .A1(n7329), .A2(n6155), .ZN(n6156) );
  INV_X2 U7322 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  NAND2_X1 U7323 ( .A1(n6158), .A2(n6157), .ZN(n6162) );
  INV_X1 U7324 ( .A(n6159), .ZN(n6160) );
  NAND2_X1 U7325 ( .A1(n6160), .A2(n8523), .ZN(n6161) );
  MUX2_X1 U7326 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(P2_DATAO_REG_28__SCAN_IN), 
        .S(n7435), .Z(n6163) );
  XNOR2_X1 U7327 ( .A(n6163), .B(n8418), .ZN(n6177) );
  NAND2_X1 U7328 ( .A1(n6176), .A2(n6177), .ZN(n6166) );
  INV_X1 U7329 ( .A(n6163), .ZN(n6164) );
  NAND2_X1 U7330 ( .A1(n6164), .A2(n8418), .ZN(n6165) );
  MUX2_X1 U7331 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .S(n7435), .Z(n6197) );
  XNOR2_X1 U7332 ( .A(n6196), .B(n6197), .ZN(n6195) );
  INV_X1 U7333 ( .A(SI_29_), .ZN(n6167) );
  NAND2_X1 U7334 ( .A1(n9666), .A2(n6217), .ZN(n6169) );
  NAND2_X1 U7335 ( .A1(n5660), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n6168) );
  NAND2_X1 U7336 ( .A1(n6222), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n6175) );
  NAND2_X1 U7337 ( .A1(n6220), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n6174) );
  INV_X1 U7338 ( .A(n6170), .ZN(n9949) );
  NAND2_X1 U7339 ( .A1(n6171), .A2(n9949), .ZN(n6173) );
  NAND2_X1 U7340 ( .A1(n6221), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n6172) );
  NAND2_X1 U7341 ( .A1(n10161), .A2(n8281), .ZN(n6432) );
  NAND2_X1 U7342 ( .A1(n9669), .A2(n6217), .ZN(n6179) );
  NAND2_X1 U7343 ( .A1(n5660), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n6178) );
  OR2_X1 U7344 ( .A1(n7366), .A2(n9942), .ZN(n6362) );
  NAND2_X1 U7345 ( .A1(n7366), .A2(n9942), .ZN(n9935) );
  INV_X1 U7346 ( .A(n10137), .ZN(n10139) );
  NAND2_X1 U7347 ( .A1(n5349), .A2(n6296), .ZN(n8792) );
  INV_X1 U7348 ( .A(n8687), .ZN(n8681) );
  AND2_X1 U7349 ( .A1(n7932), .A2(n7857), .ZN(n6386) );
  NOR2_X1 U7350 ( .A1(n7863), .A2(n6386), .ZN(n7824) );
  INV_X1 U7351 ( .A(n10549), .ZN(n10555) );
  NAND4_X1 U7352 ( .A1(n7824), .A2(n7946), .A3(n8320), .A4(n10555), .ZN(n6182)
         );
  INV_X1 U7353 ( .A(n6394), .ZN(n7947) );
  NOR2_X1 U7354 ( .A1(n7951), .A2(n7947), .ZN(n7990) );
  INV_X1 U7355 ( .A(n7981), .ZN(n6180) );
  NAND4_X1 U7356 ( .A1(n7990), .A2(n6180), .A3(n8073), .A4(n7864), .ZN(n6181)
         );
  OR3_X1 U7357 ( .A1(n8250), .A2(n6182), .A3(n6181), .ZN(n6184) );
  NOR2_X1 U7358 ( .A1(n6184), .A2(n6183), .ZN(n6185) );
  NAND4_X1 U7359 ( .A1(n8661), .A2(n5341), .A3(n6094), .A4(n6185), .ZN(n6186)
         );
  NOR4_X1 U7360 ( .A1(n8792), .A2(n8809), .A3(n8681), .A4(n6186), .ZN(n6187)
         );
  AND4_X1 U7361 ( .A1(n10108), .A2(n10121), .A3(n10139), .A4(n6187), .ZN(n6188) );
  AND2_X1 U7362 ( .A1(n6306), .A2(n6188), .ZN(n6189) );
  NAND4_X1 U7363 ( .A1(n10045), .A2(n10062), .A3(n10078), .A4(n6189), .ZN(
        n6190) );
  NOR2_X1 U7364 ( .A1(n10029), .A2(n6190), .ZN(n6191) );
  NAND3_X1 U7365 ( .A1(n9993), .A2(n10013), .A3(n6191), .ZN(n6192) );
  NOR2_X1 U7366 ( .A1(n9980), .A2(n6192), .ZN(n6193) );
  NAND2_X1 U7367 ( .A1(n6195), .A2(SI_29_), .ZN(n6200) );
  INV_X1 U7368 ( .A(n6196), .ZN(n6198) );
  NAND2_X1 U7369 ( .A1(n6198), .A2(n6197), .ZN(n6199) );
  INV_X1 U7370 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n6202) );
  INV_X1 U7371 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n6201) );
  MUX2_X1 U7372 ( .A(n6202), .B(n6201), .S(n7435), .Z(n6203) );
  INV_X1 U7373 ( .A(SI_30_), .ZN(n8517) );
  NAND2_X1 U7374 ( .A1(n6203), .A2(n8517), .ZN(n6206) );
  INV_X1 U7375 ( .A(n6203), .ZN(n6204) );
  NAND2_X1 U7376 ( .A1(n6204), .A2(SI_30_), .ZN(n6205) );
  NAND2_X1 U7377 ( .A1(n6206), .A2(n6205), .ZN(n6215) );
  MUX2_X1 U7378 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .S(n7435), .Z(n6208) );
  INV_X1 U7379 ( .A(SI_31_), .ZN(n6207) );
  XNOR2_X1 U7380 ( .A(n6208), .B(n6207), .ZN(n6209) );
  XNOR2_X2 U7381 ( .A(n6210), .B(n6209), .ZN(n8847) );
  NAND2_X1 U7382 ( .A1(n5660), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n6211) );
  NAND2_X1 U7383 ( .A1(n6220), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n6214) );
  NAND2_X1 U7384 ( .A1(n6221), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n6213) );
  NAND2_X1 U7385 ( .A1(n6222), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n6212) );
  AND3_X1 U7386 ( .A1(n6214), .A2(n6213), .A3(n6212), .ZN(n6227) );
  NAND2_X1 U7387 ( .A1(n9663), .A2(n6217), .ZN(n6219) );
  NAND2_X1 U7388 ( .A1(n5660), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n6218) );
  NAND2_X1 U7389 ( .A1(n6220), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n6225) );
  NAND2_X1 U7390 ( .A1(n6221), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n6224) );
  NAND2_X1 U7391 ( .A1(n6222), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n6223) );
  AND3_X1 U7392 ( .A1(n6225), .A2(n6224), .A3(n6223), .ZN(n9939) );
  INV_X1 U7393 ( .A(n6323), .ZN(n6339) );
  INV_X1 U7394 ( .A(n9939), .ZN(n9794) );
  NAND2_X1 U7395 ( .A1(n9794), .A2(n5408), .ZN(n6226) );
  NAND2_X1 U7396 ( .A1(n9124), .A2(n6226), .ZN(n6337) );
  OR2_X1 U7397 ( .A1(n6228), .A2(n6227), .ZN(n6338) );
  MUX2_X1 U7398 ( .A(n6432), .B(n6367), .S(n6323), .Z(n6336) );
  NAND2_X1 U7399 ( .A1(n6351), .A2(n6229), .ZN(n6347) );
  NAND2_X1 U7400 ( .A1(n6316), .A2(n6230), .ZN(n6352) );
  NAND2_X1 U7401 ( .A1(n6426), .A2(n6422), .ZN(n6232) );
  NAND2_X1 U7402 ( .A1(n10060), .A2(n6423), .ZN(n6231) );
  MUX2_X1 U7403 ( .A(n6232), .B(n6231), .S(n6323), .Z(n6233) );
  INV_X1 U7404 ( .A(n6233), .ZN(n6308) );
  NAND2_X1 U7405 ( .A1(n6421), .A2(n6339), .ZN(n6295) );
  NAND2_X1 U7406 ( .A1(n9799), .A2(n6323), .ZN(n6234) );
  OAI22_X1 U7407 ( .A1(n6416), .A2(n6323), .B1(n10210), .B2(n6234), .ZN(n6235)
         );
  INV_X1 U7408 ( .A(n6235), .ZN(n6237) );
  INV_X1 U7409 ( .A(n6300), .ZN(n6418) );
  AND2_X1 U7410 ( .A1(n6417), .A2(n6323), .ZN(n6293) );
  NAND3_X1 U7411 ( .A1(n6416), .A2(n6418), .A3(n6293), .ZN(n6236) );
  OAI211_X1 U7412 ( .C1(n6295), .C2(n6417), .A(n6237), .B(n6236), .ZN(n6238)
         );
  INV_X1 U7413 ( .A(n6238), .ZN(n6305) );
  AND2_X1 U7414 ( .A1(n6277), .A2(n6240), .ZN(n6248) );
  NAND2_X1 U7415 ( .A1(n6268), .A2(n6266), .ZN(n6245) );
  NAND2_X1 U7416 ( .A1(n6240), .A2(n6266), .ZN(n6385) );
  INV_X1 U7417 ( .A(n6241), .ZN(n6242) );
  AND2_X1 U7418 ( .A1(n6401), .A2(n6242), .ZN(n6243) );
  NOR2_X1 U7419 ( .A1(n6385), .A2(n6243), .ZN(n6244) );
  MUX2_X1 U7420 ( .A(n6245), .B(n6244), .S(n6323), .Z(n6272) );
  INV_X1 U7421 ( .A(n8173), .ZN(n6246) );
  NAND2_X1 U7422 ( .A1(n6282), .A2(n6273), .ZN(n6404) );
  AOI21_X1 U7423 ( .B1(n6272), .B2(n6246), .A(n6404), .ZN(n6247) );
  MUX2_X1 U7424 ( .A(n6248), .B(n6247), .S(n6323), .Z(n6276) );
  NAND2_X1 U7425 ( .A1(n6390), .A2(n6394), .ZN(n6249) );
  AOI21_X1 U7426 ( .B1(n7974), .B2(n7945), .A(n6249), .ZN(n6251) );
  MUX2_X1 U7427 ( .A(n6251), .B(n6250), .S(n6339), .Z(n6252) );
  NAND2_X1 U7428 ( .A1(n6252), .A2(n7946), .ZN(n6258) );
  INV_X1 U7429 ( .A(n6395), .ZN(n6255) );
  NAND2_X1 U7430 ( .A1(n7951), .A2(n6395), .ZN(n6254) );
  NAND2_X1 U7431 ( .A1(n6254), .A2(n6253), .ZN(n6397) );
  MUX2_X1 U7432 ( .A(n6255), .B(n6397), .S(n6323), .Z(n6256) );
  NOR2_X1 U7433 ( .A1(n6256), .A2(n8027), .ZN(n6257) );
  NAND2_X1 U7434 ( .A1(n6258), .A2(n6257), .ZN(n6260) );
  MUX2_X1 U7435 ( .A(n8073), .B(n8071), .S(n6323), .Z(n6259) );
  NAND3_X1 U7436 ( .A1(n6260), .A2(n5449), .A3(n6259), .ZN(n6264) );
  MUX2_X1 U7437 ( .A(n6262), .B(n6261), .S(n6323), .Z(n6263) );
  NAND3_X1 U7438 ( .A1(n6264), .A2(n4945), .A3(n6263), .ZN(n6271) );
  INV_X1 U7439 ( .A(n6265), .ZN(n6267) );
  AOI21_X1 U7440 ( .B1(n6267), .B2(n6266), .A(n6323), .ZN(n6269) );
  NOR2_X1 U7441 ( .A1(n6269), .A2(n6268), .ZN(n6270) );
  NAND2_X1 U7442 ( .A1(n6271), .A2(n6270), .ZN(n6274) );
  NAND3_X1 U7443 ( .A1(n6274), .A2(n6273), .A3(n6272), .ZN(n6275) );
  NAND2_X1 U7444 ( .A1(n6276), .A2(n6275), .ZN(n6283) );
  AND2_X1 U7445 ( .A1(n6284), .A2(n6277), .ZN(n6407) );
  INV_X1 U7446 ( .A(n6408), .ZN(n6278) );
  AOI21_X1 U7447 ( .B1(n6283), .B2(n6407), .A(n6278), .ZN(n6281) );
  INV_X1 U7448 ( .A(n6279), .ZN(n6287) );
  OAI21_X1 U7449 ( .B1(n6281), .B2(n6287), .A(n6280), .ZN(n6291) );
  NAND3_X1 U7450 ( .A1(n6283), .A2(n6408), .A3(n6282), .ZN(n6285) );
  NAND2_X1 U7451 ( .A1(n6285), .A2(n6284), .ZN(n6286) );
  NAND2_X1 U7452 ( .A1(n6286), .A2(n8791), .ZN(n6289) );
  NOR2_X1 U7453 ( .A1(n6288), .A2(n6287), .ZN(n6412) );
  NAND2_X1 U7454 ( .A1(n6289), .A2(n6412), .ZN(n6290) );
  MUX2_X1 U7455 ( .A(n6291), .B(n6290), .S(n6339), .Z(n6298) );
  NAND3_X1 U7456 ( .A1(n6298), .A2(n6413), .A3(n5349), .ZN(n6292) );
  NAND2_X1 U7457 ( .A1(n6292), .A2(n6297), .ZN(n6294) );
  NAND3_X1 U7458 ( .A1(n6294), .A2(n6293), .A3(n6416), .ZN(n6304) );
  INV_X1 U7459 ( .A(n6295), .ZN(n6302) );
  AND2_X1 U7460 ( .A1(n6297), .A2(n6296), .ZN(n6415) );
  NAND2_X1 U7461 ( .A1(n6298), .A2(n6415), .ZN(n6299) );
  NAND2_X1 U7462 ( .A1(n6299), .A2(n6413), .ZN(n6301) );
  NAND3_X1 U7463 ( .A1(n6302), .A2(n6301), .A3(n6300), .ZN(n6303) );
  NAND4_X1 U7464 ( .A1(n6306), .A2(n6305), .A3(n6304), .A4(n6303), .ZN(n6307)
         );
  NAND2_X1 U7465 ( .A1(n6308), .A2(n6307), .ZN(n6312) );
  NAND2_X1 U7466 ( .A1(n6309), .A2(n6339), .ZN(n6311) );
  OR2_X1 U7467 ( .A1(n6426), .A2(n6339), .ZN(n6310) );
  NAND4_X1 U7468 ( .A1(n6312), .A2(n6311), .A3(n6427), .A4(n6310), .ZN(n6315)
         );
  MUX2_X1 U7469 ( .A(n6313), .B(n6427), .S(n6339), .Z(n6314) );
  AOI21_X1 U7470 ( .B1(n6315), .B2(n6314), .A(n10041), .ZN(n6318) );
  MUX2_X1 U7471 ( .A(n6351), .B(n6316), .S(n6323), .Z(n6317) );
  OAI211_X1 U7472 ( .C1(n6319), .C2(n6318), .A(n10013), .B(n6317), .ZN(n6327)
         );
  INV_X1 U7473 ( .A(n6358), .ZN(n6320) );
  AOI21_X1 U7474 ( .B1(n6327), .B2(n6355), .A(n6320), .ZN(n6322) );
  INV_X1 U7475 ( .A(n6325), .ZN(n6321) );
  INV_X1 U7476 ( .A(n6326), .ZN(n6324) );
  NAND2_X1 U7477 ( .A1(n6326), .A2(n6325), .ZN(n6360) );
  INV_X1 U7478 ( .A(n6360), .ZN(n6329) );
  NAND3_X1 U7479 ( .A1(n6327), .A2(n9993), .A3(n6354), .ZN(n6328) );
  NAND3_X1 U7480 ( .A1(n6330), .A2(n6329), .A3(n6328), .ZN(n6331) );
  MUX2_X1 U7481 ( .A(n7358), .B(n6344), .S(n6339), .Z(n6332) );
  MUX2_X1 U7482 ( .A(n9935), .B(n6362), .S(n6339), .Z(n6334) );
  AND2_X1 U7483 ( .A1(n6341), .A2(n6338), .ZN(n6370) );
  INV_X1 U7484 ( .A(n6370), .ZN(n6340) );
  INV_X1 U7485 ( .A(n6378), .ZN(n6343) );
  OAI22_X1 U7486 ( .A1(n6343), .A2(n6342), .B1(n6072), .B2(n6070), .ZN(n6380)
         );
  OAI211_X1 U7487 ( .C1(n5401), .C2(n6070), .A(n6072), .B(n6065), .ZN(n6377)
         );
  AND2_X1 U7488 ( .A1(n9935), .A2(n6344), .ZN(n6365) );
  INV_X1 U7489 ( .A(n6365), .ZN(n6431) );
  INV_X1 U7490 ( .A(n6345), .ZN(n6350) );
  INV_X1 U7491 ( .A(n6346), .ZN(n6349) );
  INV_X1 U7492 ( .A(n6355), .ZN(n6348) );
  OR4_X1 U7493 ( .A1(n6360), .A2(n6349), .A3(n6348), .A4(n6347), .ZN(n6384) );
  NOR3_X1 U7494 ( .A1(n6431), .A2(n6350), .A3(n6384), .ZN(n6369) );
  NAND2_X1 U7495 ( .A1(n6352), .A2(n6351), .ZN(n6353) );
  NAND2_X1 U7496 ( .A1(n6354), .A2(n6353), .ZN(n6356) );
  NAND2_X1 U7497 ( .A1(n6356), .A2(n6355), .ZN(n6357) );
  AND2_X1 U7498 ( .A1(n6358), .A2(n6357), .ZN(n6361) );
  OAI211_X1 U7499 ( .C1(n6361), .C2(n6360), .A(n7358), .B(n6359), .ZN(n6364)
         );
  INV_X1 U7500 ( .A(n6362), .ZN(n6363) );
  AOI21_X1 U7501 ( .B1(n6365), .B2(n6364), .A(n6363), .ZN(n6366) );
  NAND2_X1 U7502 ( .A1(n6367), .A2(n6366), .ZN(n6434) );
  OAI21_X1 U7503 ( .B1(n4948), .B2(n9939), .A(n9124), .ZN(n6368) );
  OAI211_X1 U7504 ( .C1(n6369), .C2(n6434), .A(n6368), .B(n6432), .ZN(n6371)
         );
  NOR2_X1 U7505 ( .A1(n6373), .A2(n6372), .ZN(n6374) );
  OAI21_X1 U7506 ( .B1(n6378), .B2(n6377), .A(n6376), .ZN(n6379) );
  AOI21_X1 U7507 ( .B1(n6381), .B2(n6380), .A(n6379), .ZN(n6382) );
  INV_X1 U7508 ( .A(n6383), .ZN(n6437) );
  INV_X1 U7509 ( .A(n6384), .ZN(n6429) );
  INV_X1 U7510 ( .A(n6385), .ZN(n6406) );
  AOI21_X1 U7511 ( .B1(n6960), .B2(n6965), .A(n8320), .ZN(n6388) );
  INV_X1 U7512 ( .A(n6386), .ZN(n6387) );
  AND2_X1 U7513 ( .A1(n6388), .A2(n6387), .ZN(n6391) );
  OAI211_X1 U7514 ( .C1(n6392), .C2(n6391), .A(n6390), .B(n6389), .ZN(n6393)
         );
  NAND2_X1 U7515 ( .A1(n6393), .A2(n7945), .ZN(n6396) );
  NAND3_X1 U7516 ( .A1(n6396), .A2(n6395), .A3(n6394), .ZN(n6400) );
  INV_X1 U7517 ( .A(n6397), .ZN(n6399) );
  AOI21_X1 U7518 ( .B1(n6400), .B2(n6399), .A(n6398), .ZN(n6403) );
  OAI21_X1 U7519 ( .B1(n6403), .B2(n6402), .A(n6401), .ZN(n6405) );
  AOI21_X1 U7520 ( .B1(n6406), .B2(n6405), .A(n6404), .ZN(n6410) );
  INV_X1 U7521 ( .A(n6407), .ZN(n6409) );
  OAI211_X1 U7522 ( .C1(n6410), .C2(n6409), .A(n8791), .B(n6408), .ZN(n6411)
         );
  NAND2_X1 U7523 ( .A1(n6412), .A2(n6411), .ZN(n6414) );
  AOI21_X1 U7524 ( .B1(n6415), .B2(n6414), .A(n5347), .ZN(n6419) );
  OAI211_X1 U7525 ( .C1(n6419), .C2(n6418), .A(n6417), .B(n6416), .ZN(n6420)
         );
  NAND3_X1 U7526 ( .A1(n6422), .A2(n6421), .A3(n6420), .ZN(n6424) );
  NAND2_X1 U7527 ( .A1(n6424), .A2(n6423), .ZN(n6425) );
  NAND3_X1 U7528 ( .A1(n6427), .A2(n6426), .A3(n6425), .ZN(n6428) );
  NAND2_X1 U7529 ( .A1(n6429), .A2(n6428), .ZN(n6430) );
  NOR2_X1 U7530 ( .A1(n6431), .A2(n6430), .ZN(n6433) );
  OAI211_X1 U7531 ( .C1(n6434), .C2(n6433), .A(n4989), .B(n6432), .ZN(n6436)
         );
  AOI21_X1 U7532 ( .B1(n6437), .B2(n6436), .A(n6435), .ZN(n6438) );
  XNOR2_X1 U7533 ( .A(n6438), .B(n6070), .ZN(n6439) );
  OR2_X1 U7534 ( .A1(n7397), .A2(P1_U3086), .ZN(n8381) );
  NAND2_X1 U7535 ( .A1(n6441), .A2(n6440), .ZN(n6449) );
  INV_X1 U7536 ( .A(n6442), .ZN(n7823) );
  AND2_X1 U7537 ( .A1(n10274), .A2(n7823), .ZN(n7181) );
  NAND2_X1 U7538 ( .A1(n6444), .A2(n6443), .ZN(n10294) );
  OR2_X1 U7539 ( .A1(n9821), .A2(n10294), .ZN(n7474) );
  INV_X1 U7540 ( .A(n7474), .ZN(n6445) );
  NAND2_X1 U7541 ( .A1(n7181), .A2(n6445), .ZN(n6446) );
  OAI211_X1 U7542 ( .C1(n6447), .C2(n8381), .A(n6446), .B(P1_B_REG_SCAN_IN), 
        .ZN(n6448) );
  NAND2_X1 U7543 ( .A1(n6449), .A2(n6448), .ZN(P1_U3242) );
  NAND2_X1 U7544 ( .A1(n7711), .A2(n7782), .ZN(n6549) );
  INV_X1 U7545 ( .A(n6549), .ZN(n6451) );
  NAND2_X1 U7546 ( .A1(n6451), .A2(n6450), .ZN(n6565) );
  NOR2_X1 U7547 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_REG3_REG_10__SCAN_IN), 
        .ZN(n6453) );
  INV_X1 U7548 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n6461) );
  INV_X1 U7549 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n8596) );
  NAND2_X1 U7550 ( .A1(n6781), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n6464) );
  NAND2_X1 U7551 ( .A1(n6795), .A2(n6464), .ZN(n9429) );
  AND2_X1 U7552 ( .A1(n6466), .A2(n6465), .ZN(n6470) );
  NOR2_X1 U7553 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), .ZN(
        n6469) );
  NOR2_X1 U7554 ( .A1(P2_IR_REG_10__SCAN_IN), .A2(P2_IR_REG_8__SCAN_IN), .ZN(
        n6468) );
  NOR2_X1 U7555 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n6467) );
  NAND4_X1 U7556 ( .A1(n6470), .A2(n6469), .A3(n6468), .A4(n6467), .ZN(n6475)
         );
  NOR2_X2 U7557 ( .A1(n6475), .A2(n6592), .ZN(n6713) );
  INV_X1 U7558 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n6478) );
  INV_X1 U7559 ( .A(n6481), .ZN(n6494) );
  NAND2_X1 U7560 ( .A1(n6494), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6482) );
  NAND2_X1 U7561 ( .A1(n9429), .A2(n6720), .ZN(n6492) );
  INV_X1 U7562 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n6489) );
  AND2_X2 U7563 ( .A1(n9664), .A2(n6485), .ZN(n6929) );
  INV_X2 U7564 ( .A(n6842), .ZN(n8850) );
  AND2_X2 U7565 ( .A1(n9667), .A2(n6486), .ZN(n6526) );
  NAND2_X1 U7566 ( .A1(n8851), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n6488) );
  NAND2_X1 U7567 ( .A1(n8852), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n6487) );
  OAI211_X1 U7568 ( .C1(n6489), .C2(n6842), .A(n6488), .B(n6487), .ZN(n6490)
         );
  INV_X1 U7569 ( .A(n6490), .ZN(n6491) );
  NAND2_X1 U7570 ( .A1(n6498), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6493) );
  NAND2_X1 U7571 ( .A1(n6496), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6497) );
  NAND2_X1 U7572 ( .A1(n6499), .A2(n6498), .ZN(n6846) );
  OR2_X1 U7573 ( .A1(n8785), .A2(n6756), .ZN(n6501) );
  NAND2_X1 U7574 ( .A1(n8844), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n6500) );
  INV_X1 U7575 ( .A(n9564), .ZN(n9431) );
  NAND2_X1 U7576 ( .A1(n6929), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n6505) );
  NAND2_X1 U7577 ( .A1(n6527), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n6504) );
  NAND2_X1 U7578 ( .A1(n6526), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n6503) );
  NAND2_X1 U7579 ( .A1(n6519), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n6502) );
  NAND2_X1 U7580 ( .A1(n6667), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n6507) );
  INV_X4 U7581 ( .A(n6515), .ZN(n6532) );
  NAND2_X1 U7582 ( .A1(n8921), .A2(n8928), .ZN(n6850) );
  NAND2_X1 U7583 ( .A1(n6519), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n6513) );
  NAND2_X1 U7584 ( .A1(n6929), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6512) );
  NAND2_X1 U7585 ( .A1(n6526), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6511) );
  NAND2_X1 U7586 ( .A1(n6527), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n6510) );
  NAND2_X1 U7587 ( .A1(n7427), .A2(SI_0_), .ZN(n6514) );
  XNOR2_X1 U7588 ( .A(n6514), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n9677) );
  NAND2_X1 U7589 ( .A1(n7503), .A2(n6508), .ZN(n6516) );
  NAND2_X1 U7590 ( .A1(n6526), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6518) );
  NAND2_X1 U7591 ( .A1(n6527), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n6517) );
  NAND2_X1 U7592 ( .A1(n6929), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6521) );
  NAND2_X1 U7593 ( .A1(n6519), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n6520) );
  AND3_X2 U7594 ( .A1(n5517), .A2(n6521), .A3(n6520), .ZN(n7727) );
  NAND2_X1 U7595 ( .A1(n6667), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n6523) );
  NAND2_X1 U7596 ( .A1(n6532), .A2(n7582), .ZN(n6522) );
  NAND2_X1 U7597 ( .A1(n7727), .A2(n7558), .ZN(n8931) );
  INV_X1 U7598 ( .A(n7727), .ZN(n9291) );
  INV_X1 U7599 ( .A(n7558), .ZN(n10586) );
  NAND2_X1 U7600 ( .A1(n7741), .A2(n6851), .ZN(n6525) );
  NAND2_X1 U7601 ( .A1(n7727), .A2(n10586), .ZN(n6524) );
  NAND2_X1 U7602 ( .A1(n6526), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6530) );
  NAND2_X1 U7603 ( .A1(n6527), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n6529) );
  NAND2_X1 U7604 ( .A1(n6929), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n6528) );
  NAND2_X1 U7605 ( .A1(n8848), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n6537) );
  NAND2_X1 U7606 ( .A1(n8849), .A2(n6531), .ZN(n6536) );
  NAND2_X1 U7607 ( .A1(n4968), .A2(n5186), .ZN(n6545) );
  NAND2_X1 U7608 ( .A1(n6545), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6534) );
  INV_X1 U7609 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n6533) );
  XNOR2_X1 U7610 ( .A(n6534), .B(n6533), .ZN(n7434) );
  INV_X1 U7611 ( .A(n7434), .ZN(n10360) );
  NAND2_X1 U7612 ( .A1(n6532), .A2(n10360), .ZN(n6535) );
  INV_X1 U7613 ( .A(n7725), .ZN(n7783) );
  NOR2_X1 U7614 ( .A1(n9290), .A2(n7783), .ZN(n6538) );
  NAND2_X1 U7615 ( .A1(n8851), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n6544) );
  NAND2_X1 U7616 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n6539) );
  NAND2_X1 U7617 ( .A1(n6549), .A2(n6539), .ZN(n7845) );
  NAND2_X1 U7618 ( .A1(n6720), .A2(n7845), .ZN(n6543) );
  INV_X2 U7619 ( .A(n6540), .ZN(n8852) );
  NAND2_X1 U7620 ( .A1(n8852), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n6542) );
  NAND2_X1 U7621 ( .A1(n8850), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n6541) );
  AND4_X2 U7622 ( .A1(n6544), .A2(n6543), .A3(n6542), .A4(n6541), .ZN(n6853)
         );
  NAND2_X1 U7623 ( .A1(n8848), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n6547) );
  NAND2_X1 U7624 ( .A1(n6586), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6556) );
  NAND2_X1 U7625 ( .A1(n6532), .A2(n10376), .ZN(n6546) );
  OAI211_X1 U7626 ( .C1(n6756), .C2(n7443), .A(n6547), .B(n6546), .ZN(n7846)
         );
  NAND2_X1 U7627 ( .A1(n6853), .A2(n5150), .ZN(n6548) );
  NAND2_X1 U7628 ( .A1(n8851), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6554) );
  NAND2_X1 U7629 ( .A1(n6549), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n6550) );
  NAND2_X1 U7630 ( .A1(n6565), .A2(n6550), .ZN(n7939) );
  NAND2_X1 U7631 ( .A1(n6720), .A2(n7939), .ZN(n6553) );
  NAND2_X1 U7632 ( .A1(n8852), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n6552) );
  NAND2_X1 U7633 ( .A1(n8850), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n6551) );
  NAND4_X1 U7634 ( .A1(n6554), .A2(n6553), .A3(n6552), .A4(n6551), .ZN(n9288)
         );
  NAND2_X1 U7635 ( .A1(n7936), .A2(n9288), .ZN(n6564) );
  INV_X1 U7636 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n6583) );
  NAND2_X1 U7637 ( .A1(n6556), .A2(n6583), .ZN(n6557) );
  NAND2_X1 U7638 ( .A1(n6557), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6558) );
  NAND2_X1 U7639 ( .A1(n6558), .A2(n6584), .ZN(n6571) );
  OR2_X1 U7640 ( .A1(n6558), .A2(n6584), .ZN(n6559) );
  AOI22_X1 U7641 ( .A1(n8848), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n6532), .B2(
        n7290), .ZN(n6561) );
  OR2_X1 U7642 ( .A1(n7447), .A2(n6756), .ZN(n6560) );
  NAND2_X1 U7643 ( .A1(n6561), .A2(n6560), .ZN(n7940) );
  NAND2_X1 U7644 ( .A1(n6562), .A2(n7940), .ZN(n6563) );
  NAND2_X1 U7645 ( .A1(n8851), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6570) );
  NAND2_X1 U7646 ( .A1(n6565), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n6566) );
  NAND2_X1 U7647 ( .A1(n6576), .A2(n6566), .ZN(n7761) );
  NAND2_X1 U7648 ( .A1(n6720), .A2(n7761), .ZN(n6569) );
  NAND2_X1 U7649 ( .A1(n8852), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n6568) );
  NAND2_X1 U7650 ( .A1(n8850), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n6567) );
  NAND4_X1 U7651 ( .A1(n6570), .A2(n6569), .A3(n6568), .A4(n6567), .ZN(n9287)
         );
  OR2_X1 U7652 ( .A1(n7449), .A2(n6756), .ZN(n6574) );
  NAND2_X1 U7653 ( .A1(n6571), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6572) );
  AOI22_X1 U7654 ( .A1(n8848), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n6532), .B2(
        n10414), .ZN(n6573) );
  NAND2_X1 U7655 ( .A1(n6574), .A2(n6573), .ZN(n7970) );
  INV_X1 U7656 ( .A(n7970), .ZN(n7963) );
  NAND2_X1 U7657 ( .A1(n8851), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6581) );
  NAND2_X1 U7658 ( .A1(n6576), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n6577) );
  NAND2_X1 U7659 ( .A1(n6595), .A2(n6577), .ZN(n8063) );
  NAND2_X1 U7660 ( .A1(n6720), .A2(n8063), .ZN(n6580) );
  NAND2_X1 U7661 ( .A1(n8852), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n6579) );
  NAND2_X1 U7662 ( .A1(n8850), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n6578) );
  NAND4_X1 U7663 ( .A1(n6581), .A2(n6580), .A3(n6579), .A4(n6578), .ZN(n9286)
         );
  OR2_X1 U7664 ( .A1(n7453), .A2(n6756), .ZN(n6589) );
  INV_X1 U7665 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n6582) );
  NAND3_X1 U7666 ( .A1(n6584), .A2(n6583), .A3(n6582), .ZN(n6585) );
  OAI21_X1 U7667 ( .B1(n6586), .B2(n6585), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n6587) );
  XNOR2_X1 U7668 ( .A(n6587), .B(P2_IR_REG_7__SCAN_IN), .ZN(n10431) );
  AOI22_X1 U7669 ( .A1(n8848), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n6532), .B2(
        n10431), .ZN(n6588) );
  NAND2_X1 U7670 ( .A1(n6589), .A2(n6588), .ZN(n8096) );
  OR2_X1 U7671 ( .A1(n8010), .A2(n8096), .ZN(n8294) );
  NAND2_X1 U7672 ( .A1(n8096), .A2(n8010), .ZN(n8916) );
  NAND2_X1 U7673 ( .A1(n8294), .A2(n8916), .ZN(n8954) );
  OR2_X1 U7674 ( .A1(n8096), .A2(n9286), .ZN(n6590) );
  NAND2_X1 U7675 ( .A1(n6591), .A2(n6590), .ZN(n8188) );
  NAND2_X1 U7676 ( .A1(n6592), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6593) );
  XNOR2_X1 U7677 ( .A(n6593), .B(P2_IR_REG_8__SCAN_IN), .ZN(n10447) );
  AOI22_X1 U7678 ( .A1(n8848), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n6532), .B2(
        n10447), .ZN(n6594) );
  NAND2_X1 U7679 ( .A1(n8851), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n6600) );
  NAND2_X1 U7680 ( .A1(n6595), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n6596) );
  NAND2_X1 U7681 ( .A1(n6613), .A2(n6596), .ZN(n10635) );
  NAND2_X1 U7682 ( .A1(n6720), .A2(n10635), .ZN(n6599) );
  NAND2_X1 U7683 ( .A1(n8850), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n6598) );
  NAND2_X1 U7684 ( .A1(n8852), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n6597) );
  INV_X1 U7685 ( .A(n8914), .ZN(n6857) );
  NAND2_X1 U7686 ( .A1(n10637), .A2(n8192), .ZN(n8913) );
  INV_X1 U7687 ( .A(n8886), .ZN(n8297) );
  NAND2_X1 U7688 ( .A1(n8623), .A2(n8849), .ZN(n6603) );
  OR2_X1 U7689 ( .A1(n6592), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n6608) );
  NAND2_X1 U7690 ( .A1(n6608), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6601) );
  XNOR2_X1 U7691 ( .A(n6601), .B(P2_IR_REG_9__SCAN_IN), .ZN(n10463) );
  AOI22_X1 U7692 ( .A1(n8848), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6532), .B2(
        n10463), .ZN(n6602) );
  NAND2_X1 U7693 ( .A1(n8851), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n6607) );
  XNOR2_X1 U7694 ( .A(n6613), .B(P2_REG3_REG_9__SCAN_IN), .ZN(n8195) );
  NAND2_X1 U7695 ( .A1(n6720), .A2(n8195), .ZN(n6606) );
  NAND2_X1 U7696 ( .A1(n8852), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n6605) );
  NAND2_X1 U7697 ( .A1(n8850), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n6604) );
  NAND4_X1 U7698 ( .A1(n6607), .A2(n6606), .A3(n6605), .A4(n6604), .ZN(n9284)
         );
  INV_X1 U7699 ( .A(n8961), .ZN(n6859) );
  OR2_X1 U7700 ( .A1(n8241), .A2(n9284), .ZN(n6620) );
  AND2_X1 U7701 ( .A1(n8297), .A2(n6621), .ZN(n8212) );
  OR2_X1 U7702 ( .A1(n7465), .A2(n6756), .ZN(n6612) );
  NOR2_X1 U7703 ( .A1(n6608), .A2(P2_IR_REG_9__SCAN_IN), .ZN(n6627) );
  OR2_X1 U7704 ( .A1(n6627), .A2(n6609), .ZN(n6610) );
  XNOR2_X1 U7705 ( .A(n6610), .B(P2_IR_REG_10__SCAN_IN), .ZN(n10479) );
  AOI22_X1 U7706 ( .A1(n8848), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6532), .B2(
        n10479), .ZN(n6611) );
  NAND2_X1 U7707 ( .A1(n8851), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n6618) );
  OAI21_X1 U7708 ( .B1(n6613), .B2(P2_REG3_REG_9__SCAN_IN), .A(
        P2_REG3_REG_10__SCAN_IN), .ZN(n6614) );
  NAND2_X1 U7709 ( .A1(n6614), .A2(n6631), .ZN(n8264) );
  NAND2_X1 U7710 ( .A1(n6720), .A2(n8264), .ZN(n6617) );
  NAND2_X1 U7711 ( .A1(n8852), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n6616) );
  NAND2_X1 U7712 ( .A1(n8850), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n6615) );
  NAND4_X1 U7713 ( .A1(n6618), .A2(n6617), .A3(n6616), .A4(n6615), .ZN(n9283)
         );
  NAND2_X1 U7714 ( .A1(n8359), .A2(n8353), .ZN(n8964) );
  AND2_X1 U7715 ( .A1(n8212), .A2(n8888), .ZN(n6619) );
  NAND2_X1 U7716 ( .A1(n8188), .A2(n6619), .ZN(n6625) );
  INV_X1 U7717 ( .A(n8888), .ZN(n6622) );
  INV_X1 U7718 ( .A(n8192), .ZN(n9285) );
  OR2_X1 U7719 ( .A1(n10637), .A2(n9285), .ZN(n8189) );
  NAND2_X1 U7720 ( .A1(n6625), .A2(n6624), .ZN(n8309) );
  NAND2_X1 U7721 ( .A1(n7480), .A2(n8849), .ZN(n6630) );
  INV_X1 U7722 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n6626) );
  NAND2_X1 U7723 ( .A1(n6627), .A2(n6626), .ZN(n6641) );
  NAND2_X1 U7724 ( .A1(n6641), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6628) );
  XNOR2_X1 U7725 ( .A(n6628), .B(P2_IR_REG_11__SCAN_IN), .ZN(n10496) );
  AOI22_X1 U7726 ( .A1(n8848), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n6532), .B2(
        n10496), .ZN(n6629) );
  NAND2_X1 U7727 ( .A1(n6630), .A2(n6629), .ZN(n8397) );
  NAND2_X1 U7728 ( .A1(n8851), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n6636) );
  NAND2_X1 U7729 ( .A1(n6631), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6632) );
  NAND2_X1 U7730 ( .A1(n6645), .A2(n6632), .ZN(n8350) );
  NAND2_X1 U7731 ( .A1(n6720), .A2(n8350), .ZN(n6635) );
  NAND2_X1 U7732 ( .A1(n8852), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n6634) );
  NAND2_X1 U7733 ( .A1(n8850), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n6633) );
  NAND4_X1 U7734 ( .A1(n6636), .A2(n6635), .A3(n6634), .A4(n6633), .ZN(n9282)
         );
  NOR2_X1 U7735 ( .A1(n8397), .A2(n8388), .ZN(n8969) );
  INV_X1 U7736 ( .A(n8969), .ZN(n6637) );
  INV_X1 U7737 ( .A(n8890), .ZN(n6638) );
  NAND2_X1 U7738 ( .A1(n8309), .A2(n6638), .ZN(n6640) );
  OR2_X1 U7739 ( .A1(n8397), .A2(n9282), .ZN(n6639) );
  OR2_X1 U7740 ( .A1(n7487), .A2(n6756), .ZN(n6644) );
  NAND2_X1 U7741 ( .A1(n6642), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6653) );
  XNOR2_X1 U7742 ( .A(n6653), .B(P2_IR_REG_12__SCAN_IN), .ZN(n7281) );
  AOI22_X1 U7743 ( .A1(n8844), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n6532), .B2(
        n7281), .ZN(n6643) );
  NAND2_X1 U7744 ( .A1(n6644), .A2(n6643), .ZN(n8715) );
  NAND2_X1 U7745 ( .A1(n8851), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n6650) );
  NAND2_X1 U7746 ( .A1(n6645), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n6646) );
  NAND2_X1 U7747 ( .A1(n6657), .A2(n6646), .ZN(n8389) );
  NAND2_X1 U7748 ( .A1(n6720), .A2(n8389), .ZN(n6649) );
  NAND2_X1 U7749 ( .A1(n8852), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n6648) );
  NAND2_X1 U7750 ( .A1(n8850), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n6647) );
  OR2_X1 U7751 ( .A1(n8715), .A2(n9281), .ZN(n8370) );
  INV_X1 U7752 ( .A(n8370), .ZN(n8385) );
  AND2_X1 U7753 ( .A1(n8715), .A2(n9281), .ZN(n8384) );
  INV_X1 U7754 ( .A(n8384), .ZN(n6651) );
  OR2_X1 U7755 ( .A1(n7650), .A2(n6756), .ZN(n6656) );
  INV_X1 U7756 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n6652) );
  NAND2_X1 U7757 ( .A1(n6653), .A2(n6652), .ZN(n6654) );
  NAND2_X1 U7758 ( .A1(n6654), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6665) );
  XNOR2_X1 U7759 ( .A(n6665), .B(P2_IR_REG_13__SCAN_IN), .ZN(n7279) );
  AOI22_X1 U7760 ( .A1(n8848), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n6532), .B2(
        n7279), .ZN(n6655) );
  NAND2_X1 U7761 ( .A1(n6656), .A2(n6655), .ZN(n8694) );
  NAND2_X1 U7762 ( .A1(n8851), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n6662) );
  NAND2_X1 U7763 ( .A1(n6657), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n6658) );
  NAND2_X1 U7764 ( .A1(n6670), .A2(n6658), .ZN(n10676) );
  NAND2_X1 U7765 ( .A1(n6720), .A2(n10676), .ZN(n6661) );
  NAND2_X1 U7766 ( .A1(n8850), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n6660) );
  NAND2_X1 U7767 ( .A1(n8852), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n6659) );
  NAND4_X1 U7768 ( .A1(n6662), .A2(n6661), .A3(n6660), .A4(n6659), .ZN(n9280)
         );
  OR2_X1 U7769 ( .A1(n8694), .A2(n8718), .ZN(n8978) );
  NAND2_X1 U7770 ( .A1(n8694), .A2(n8718), .ZN(n8977) );
  NAND2_X1 U7771 ( .A1(n8978), .A2(n8977), .ZN(n8974) );
  NAND2_X1 U7772 ( .A1(n8694), .A2(n9280), .ZN(n6663) );
  NAND2_X1 U7773 ( .A1(n7668), .A2(n8849), .ZN(n6669) );
  INV_X1 U7774 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n6664) );
  NAND2_X1 U7775 ( .A1(n6665), .A2(n6664), .ZN(n6666) );
  NAND2_X1 U7776 ( .A1(n6666), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6677) );
  XNOR2_X1 U7777 ( .A(n6677), .B(P2_IR_REG_14__SCAN_IN), .ZN(n7277) );
  AOI22_X1 U7778 ( .A1(n6667), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n6532), .B2(
        n7277), .ZN(n6668) );
  NAND2_X1 U7779 ( .A1(n8851), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n6675) );
  NAND2_X1 U7780 ( .A1(n6670), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n6671) );
  NAND2_X1 U7781 ( .A1(n6681), .A2(n6671), .ZN(n8724) );
  NAND2_X1 U7782 ( .A1(n6720), .A2(n8724), .ZN(n6674) );
  NAND2_X1 U7783 ( .A1(n8852), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n6673) );
  NAND2_X1 U7784 ( .A1(n8850), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n6672) );
  NAND4_X1 U7785 ( .A1(n6675), .A2(n6674), .A3(n6673), .A4(n6672), .ZN(n9279)
         );
  XNOR2_X1 U7786 ( .A(n8728), .B(n9279), .ZN(n8987) );
  INV_X1 U7787 ( .A(n8987), .ZN(n8673) );
  NAND2_X1 U7788 ( .A1(n8728), .A2(n9279), .ZN(n8982) );
  OR2_X1 U7789 ( .A1(n7704), .A2(n6756), .ZN(n6680) );
  INV_X1 U7790 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n6676) );
  NAND2_X1 U7791 ( .A1(n6677), .A2(n6676), .ZN(n6678) );
  NAND2_X1 U7792 ( .A1(n6678), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6690) );
  XNOR2_X1 U7793 ( .A(n6690), .B(P2_IR_REG_15__SCAN_IN), .ZN(n7275) );
  AOI22_X1 U7794 ( .A1(n8848), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n6532), .B2(
        n7275), .ZN(n6679) );
  NAND2_X1 U7795 ( .A1(n8851), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n6686) );
  NAND2_X1 U7796 ( .A1(n6681), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n6682) );
  NAND2_X1 U7797 ( .A1(n6694), .A2(n6682), .ZN(n9267) );
  NAND2_X1 U7798 ( .A1(n6720), .A2(n9267), .ZN(n6685) );
  NAND2_X1 U7799 ( .A1(n8852), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n6684) );
  NAND2_X1 U7800 ( .A1(n8850), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n6683) );
  NAND4_X1 U7801 ( .A1(n6686), .A2(n6685), .A3(n6684), .A4(n6683), .ZN(n9278)
         );
  NAND2_X1 U7802 ( .A1(n8747), .A2(n8983), .ZN(n6688) );
  NAND2_X1 U7803 ( .A1(n9083), .A2(n9278), .ZN(n6687) );
  NAND2_X1 U7804 ( .A1(n6688), .A2(n6687), .ZN(n8773) );
  NAND2_X1 U7805 ( .A1(n7758), .A2(n8849), .ZN(n6693) );
  INV_X1 U7806 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n6689) );
  NAND2_X1 U7807 ( .A1(n6690), .A2(n6689), .ZN(n6691) );
  NAND2_X1 U7808 ( .A1(n6691), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6702) );
  XNOR2_X1 U7809 ( .A(n6702), .B(P2_IR_REG_16__SCAN_IN), .ZN(n7273) );
  AOI22_X1 U7810 ( .A1(n8844), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n7273), .B2(
        n6532), .ZN(n6692) );
  NAND2_X1 U7811 ( .A1(n8851), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n6699) );
  NAND2_X1 U7812 ( .A1(n6694), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n6695) );
  NAND2_X1 U7813 ( .A1(n6707), .A2(n6695), .ZN(n9194) );
  NAND2_X1 U7814 ( .A1(n6720), .A2(n9194), .ZN(n6698) );
  NAND2_X1 U7815 ( .A1(n8850), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n6697) );
  NAND2_X1 U7816 ( .A1(n8852), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n6696) );
  NAND4_X1 U7817 ( .A1(n6699), .A2(n6698), .A3(n6697), .A4(n6696), .ZN(n9535)
         );
  INV_X1 U7818 ( .A(n9535), .ZN(n9264) );
  NAND2_X1 U7819 ( .A1(n9611), .A2(n9264), .ZN(n8997) );
  NAND2_X1 U7820 ( .A1(n8998), .A2(n8997), .ZN(n8993) );
  NAND2_X1 U7821 ( .A1(n9611), .A2(n9535), .ZN(n6700) );
  NAND2_X1 U7822 ( .A1(n7885), .A2(n8849), .ZN(n6706) );
  INV_X1 U7823 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n6701) );
  NAND2_X1 U7824 ( .A1(n6702), .A2(n6701), .ZN(n6703) );
  NAND2_X1 U7825 ( .A1(n6703), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6704) );
  XNOR2_X1 U7826 ( .A(n6704), .B(P2_IR_REG_17__SCAN_IN), .ZN(n7272) );
  AOI22_X1 U7827 ( .A1(n7272), .A2(n6532), .B1(n8848), .B2(
        P1_DATAO_REG_17__SCAN_IN), .ZN(n6705) );
  NAND2_X1 U7828 ( .A1(n8851), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n6712) );
  NAND2_X1 U7829 ( .A1(n6707), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n6708) );
  NAND2_X1 U7830 ( .A1(n6718), .A2(n6708), .ZN(n9542) );
  NAND2_X1 U7831 ( .A1(n6720), .A2(n9542), .ZN(n6711) );
  NAND2_X1 U7832 ( .A1(n8852), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n6710) );
  NAND2_X1 U7833 ( .A1(n8850), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n6709) );
  NAND4_X1 U7834 ( .A1(n6712), .A2(n6711), .A3(n6710), .A4(n6709), .ZN(n9608)
         );
  XNOR2_X1 U7835 ( .A(n9602), .B(n9516), .ZN(n9538) );
  OR2_X1 U7836 ( .A1(n7919), .A2(n6756), .ZN(n6717) );
  INV_X1 U7837 ( .A(n6713), .ZN(n6714) );
  NAND2_X1 U7838 ( .A1(n6714), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6715) );
  XNOR2_X1 U7839 ( .A(n6715), .B(P2_IR_REG_18__SCAN_IN), .ZN(n7265) );
  AOI22_X1 U7840 ( .A1(n8844), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n6532), .B2(
        n7265), .ZN(n6716) );
  INV_X1 U7841 ( .A(n9524), .ZN(n9598) );
  NAND2_X1 U7842 ( .A1(n8851), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n6724) );
  NAND2_X1 U7843 ( .A1(n6718), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n6719) );
  NAND2_X1 U7844 ( .A1(n6733), .A2(n6719), .ZN(n9521) );
  NAND2_X1 U7845 ( .A1(n6720), .A2(n9521), .ZN(n6723) );
  NAND2_X1 U7846 ( .A1(n8852), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n6722) );
  NAND2_X1 U7847 ( .A1(n8850), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n6721) );
  NAND4_X1 U7848 ( .A1(n6724), .A2(n6723), .A3(n6722), .A4(n6721), .ZN(n9277)
         );
  NAND2_X1 U7849 ( .A1(n6726), .A2(n6725), .ZN(n9499) );
  NAND2_X1 U7850 ( .A1(n8088), .A2(n8849), .ZN(n6730) );
  INV_X1 U7851 ( .A(n6727), .ZN(n6728) );
  AOI22_X1 U7852 ( .A1(n8844), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n9073), .B2(
        n6532), .ZN(n6729) );
  NAND2_X1 U7853 ( .A1(n6730), .A2(n6729), .ZN(n9169) );
  NAND2_X1 U7854 ( .A1(n8851), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n6732) );
  NAND2_X1 U7855 ( .A1(n6929), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n6731) );
  AND2_X1 U7856 ( .A1(n6732), .A2(n6731), .ZN(n6737) );
  NAND2_X1 U7857 ( .A1(n6733), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n6734) );
  NAND2_X1 U7858 ( .A1(n6741), .A2(n6734), .ZN(n9507) );
  NAND2_X1 U7859 ( .A1(n9507), .A2(n6720), .ZN(n6736) );
  NAND2_X1 U7860 ( .A1(n8852), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n6735) );
  NAND2_X1 U7861 ( .A1(n9169), .A2(n9517), .ZN(n9016) );
  NAND2_X1 U7862 ( .A1(n9015), .A2(n9016), .ZN(n9092) );
  INV_X1 U7863 ( .A(n9517), .ZN(n9484) );
  NAND2_X1 U7864 ( .A1(n8170), .A2(n8849), .ZN(n6740) );
  NAND2_X1 U7865 ( .A1(n8844), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n6739) );
  INV_X1 U7866 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n6745) );
  NAND2_X1 U7867 ( .A1(n6741), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n6742) );
  NAND2_X1 U7868 ( .A1(n6750), .A2(n6742), .ZN(n9486) );
  NAND2_X1 U7869 ( .A1(n9486), .A2(n6720), .ZN(n6744) );
  AOI22_X1 U7870 ( .A1(n8851), .A2(P2_REG1_REG_20__SCAN_IN), .B1(n8850), .B2(
        P2_REG2_REG_20__SCAN_IN), .ZN(n6743) );
  NAND2_X1 U7871 ( .A1(n9586), .A2(n9468), .ZN(n6746) );
  NAND2_X1 U7872 ( .A1(n6747), .A2(n6746), .ZN(n9017) );
  NAND2_X1 U7873 ( .A1(n9483), .A2(n9492), .ZN(n9482) );
  NAND2_X1 U7874 ( .A1(n8307), .A2(n8849), .ZN(n6749) );
  NAND2_X1 U7875 ( .A1(n8844), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n6748) );
  INV_X1 U7876 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n9474) );
  NAND2_X1 U7877 ( .A1(n6750), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n6751) );
  NAND2_X1 U7878 ( .A1(n6759), .A2(n6751), .ZN(n9471) );
  NAND2_X1 U7879 ( .A1(n9471), .A2(n6720), .ZN(n6753) );
  AOI22_X1 U7880 ( .A1(n8851), .A2(P2_REG1_REG_21__SCAN_IN), .B1(n8852), .B2(
        P2_REG0_REG_21__SCAN_IN), .ZN(n6752) );
  INV_X1 U7881 ( .A(n9027), .ZN(n6755) );
  INV_X1 U7882 ( .A(n9029), .ZN(n6754) );
  NAND2_X1 U7883 ( .A1(n6755), .A2(n6754), .ZN(n9478) );
  OR2_X1 U7884 ( .A1(n8357), .A2(n6756), .ZN(n6758) );
  NAND2_X1 U7885 ( .A1(n8848), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n6757) );
  NAND2_X1 U7886 ( .A1(n6759), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6760) );
  NAND2_X1 U7887 ( .A1(n6769), .A2(n6760), .ZN(n9462) );
  NAND2_X1 U7888 ( .A1(n9462), .A2(n6720), .ZN(n6766) );
  INV_X1 U7889 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n6763) );
  NAND2_X1 U7890 ( .A1(n8851), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n6762) );
  NAND2_X1 U7891 ( .A1(n8852), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n6761) );
  OAI211_X1 U7892 ( .C1(n6763), .C2(n6842), .A(n6762), .B(n6761), .ZN(n6764)
         );
  INV_X1 U7893 ( .A(n6764), .ZN(n6765) );
  NAND2_X1 U7894 ( .A1(n9099), .A2(n9580), .ZN(n8873) );
  NAND2_X1 U7895 ( .A1(n8378), .A2(n8849), .ZN(n6768) );
  NAND2_X1 U7896 ( .A1(n8844), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n6767) );
  INV_X1 U7897 ( .A(n9572), .ZN(n6776) );
  NAND2_X1 U7898 ( .A1(n6769), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6770) );
  NAND2_X1 U7899 ( .A1(n6779), .A2(n6770), .ZN(n9448) );
  NAND2_X1 U7900 ( .A1(n9448), .A2(n6720), .ZN(n6775) );
  INV_X1 U7901 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n9449) );
  NAND2_X1 U7902 ( .A1(n8851), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n6772) );
  NAND2_X1 U7903 ( .A1(n8852), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n6771) );
  OAI211_X1 U7904 ( .C1(n9449), .C2(n6842), .A(n6772), .B(n6771), .ZN(n6773)
         );
  INV_X1 U7905 ( .A(n6773), .ZN(n6774) );
  NOR2_X1 U7906 ( .A1(n6776), .A2(n9459), .ZN(n9034) );
  NAND2_X1 U7907 ( .A1(n8731), .A2(n8849), .ZN(n6778) );
  NAND2_X1 U7908 ( .A1(n8844), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n6777) );
  NAND2_X1 U7909 ( .A1(n6779), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n6780) );
  NAND2_X1 U7910 ( .A1(n6781), .A2(n6780), .ZN(n9440) );
  NAND2_X1 U7911 ( .A1(n9440), .A2(n6720), .ZN(n6787) );
  INV_X1 U7912 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n6784) );
  NAND2_X1 U7913 ( .A1(n8851), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n6783) );
  NAND2_X1 U7914 ( .A1(n8852), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n6782) );
  OAI211_X1 U7915 ( .C1(n6784), .C2(n6842), .A(n6783), .B(n6782), .ZN(n6785)
         );
  INV_X1 U7916 ( .A(n6785), .ZN(n6786) );
  NAND2_X1 U7917 ( .A1(n8798), .A2(n8849), .ZN(n6792) );
  NAND2_X1 U7918 ( .A1(n8848), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n6791) );
  INV_X1 U7919 ( .A(n6795), .ZN(n6794) );
  INV_X1 U7920 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n6793) );
  NAND2_X1 U7921 ( .A1(n6795), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n6796) );
  NAND2_X1 U7922 ( .A1(n6805), .A2(n6796), .ZN(n9420) );
  NAND2_X1 U7923 ( .A1(n9420), .A2(n6720), .ZN(n6802) );
  INV_X1 U7924 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n6799) );
  NAND2_X1 U7925 ( .A1(n8851), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n6798) );
  NAND2_X1 U7926 ( .A1(n8852), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n6797) );
  OAI211_X1 U7927 ( .C1(n6799), .C2(n6842), .A(n6798), .B(n6797), .ZN(n6800)
         );
  INV_X1 U7928 ( .A(n6800), .ZN(n6801) );
  NAND2_X1 U7929 ( .A1(n9672), .A2(n8849), .ZN(n6804) );
  NAND2_X1 U7930 ( .A1(n8844), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n6803) );
  INV_X1 U7931 ( .A(n9555), .ZN(n6813) );
  NAND2_X1 U7932 ( .A1(n6805), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n6806) );
  NAND2_X1 U7933 ( .A1(n6821), .A2(n6806), .ZN(n9406) );
  NAND2_X1 U7934 ( .A1(n9406), .A2(n6720), .ZN(n6812) );
  INV_X1 U7935 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n6809) );
  NAND2_X1 U7936 ( .A1(n8851), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n6808) );
  NAND2_X1 U7937 ( .A1(n8852), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n6807) );
  OAI211_X1 U7938 ( .C1(n6809), .C2(n6842), .A(n6808), .B(n6807), .ZN(n6810)
         );
  INV_X1 U7939 ( .A(n6810), .ZN(n6811) );
  NAND2_X1 U7940 ( .A1(n9404), .A2(n5505), .ZN(n6816) );
  NAND2_X1 U7941 ( .A1(n6813), .A2(n6814), .ZN(n6815) );
  NAND2_X1 U7942 ( .A1(n6816), .A2(n6815), .ZN(n6927) );
  NAND2_X1 U7943 ( .A1(n9669), .A2(n8849), .ZN(n6818) );
  NAND2_X1 U7944 ( .A1(n8844), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n6817) );
  INV_X1 U7945 ( .A(n6821), .ZN(n6820) );
  INV_X1 U7946 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n6819) );
  NAND2_X1 U7947 ( .A1(n6820), .A2(n6819), .ZN(n6942) );
  NAND2_X1 U7948 ( .A1(n6821), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n6822) );
  NAND2_X1 U7949 ( .A1(n6942), .A2(n6822), .ZN(n9139) );
  NAND2_X1 U7950 ( .A1(n9139), .A2(n6720), .ZN(n6827) );
  INV_X1 U7951 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n9140) );
  NAND2_X1 U7952 ( .A1(n8851), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n6824) );
  NAND2_X1 U7953 ( .A1(n8852), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n6823) );
  OAI211_X1 U7954 ( .C1(n9140), .C2(n6842), .A(n6824), .B(n6823), .ZN(n6825)
         );
  INV_X1 U7955 ( .A(n6825), .ZN(n6826) );
  NAND2_X1 U7956 ( .A1(n9145), .A2(n9408), .ZN(n6918) );
  XNOR2_X1 U7957 ( .A(n6927), .B(n9116), .ZN(n6849) );
  NAND2_X1 U7958 ( .A1(n6829), .A2(n6828), .ZN(n6830) );
  NAND2_X1 U7959 ( .A1(n6835), .A2(n6834), .ZN(n6831) );
  NAND2_X1 U7960 ( .A1(n6831), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6833) );
  OR2_X1 U7961 ( .A1(n8927), .A2(n9070), .ZN(n6838) );
  NAND2_X1 U7962 ( .A1(n6836), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6837) );
  NAND2_X1 U7963 ( .A1(n9078), .A2(n9073), .ZN(n7336) );
  INV_X1 U7964 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n6841) );
  NAND2_X1 U7965 ( .A1(n8851), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n6840) );
  NAND2_X1 U7966 ( .A1(n8852), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n6839) );
  OAI211_X1 U7967 ( .C1(n6842), .C2(n6841), .A(n6840), .B(n6839), .ZN(n6843)
         );
  INV_X1 U7968 ( .A(n6843), .ZN(n6844) );
  NAND2_X1 U7969 ( .A1(n8857), .A2(n6844), .ZN(n9273) );
  INV_X1 U7970 ( .A(n9273), .ZN(n6922) );
  INV_X1 U7971 ( .A(n6845), .ZN(n9075) );
  NAND2_X1 U7972 ( .A1(n9075), .A2(n7271), .ZN(n6847) );
  NOR2_X2 U7973 ( .A1(n7520), .A2(n9053), .ZN(n9609) );
  OAI22_X1 U7974 ( .A1(n6922), .A2(n9616), .B1(n6814), .B2(n9515), .ZN(n6848)
         );
  INV_X1 U7975 ( .A(n9580), .ZN(n9101) );
  INV_X1 U7976 ( .A(n9585), .ZN(n9488) );
  NAND2_X1 U7977 ( .A1(n7719), .A2(n7717), .ZN(n7716) );
  NAND2_X1 U7978 ( .A1(n7716), .A2(n8928), .ZN(n7740) );
  INV_X1 U7979 ( .A(n6851), .ZN(n7739) );
  NAND2_X1 U7980 ( .A1(n7740), .A2(n7739), .ZN(n6852) );
  NAND2_X1 U7981 ( .A1(n6852), .A2(n8931), .ZN(n7724) );
  NAND2_X1 U7982 ( .A1(n9290), .A2(n7725), .ZN(n8936) );
  NAND2_X1 U7983 ( .A1(n6853), .A2(n7846), .ZN(n8938) );
  OR2_X1 U7984 ( .A1(n6853), .A2(n7846), .ZN(n8937) );
  INV_X1 U7985 ( .A(n7940), .ZN(n8043) );
  NAND2_X1 U7986 ( .A1(n9288), .A2(n8043), .ZN(n8940) );
  NAND2_X1 U7987 ( .A1(n8937), .A2(n8940), .ZN(n8948) );
  INV_X1 U7988 ( .A(n8948), .ZN(n6854) );
  NAND2_X1 U7989 ( .A1(n7934), .A2(n6854), .ZN(n6855) );
  NAND2_X1 U7990 ( .A1(n7961), .A2(n7940), .ZN(n8946) );
  NAND2_X1 U7991 ( .A1(n6575), .A2(n7970), .ZN(n8947) );
  INV_X1 U7992 ( .A(n8947), .ZN(n6856) );
  NAND2_X1 U7993 ( .A1(n7963), .A2(n9287), .ZN(n8950) );
  INV_X1 U7994 ( .A(n8954), .ZN(n8885) );
  NAND2_X1 U7995 ( .A1(n6857), .A2(n8294), .ZN(n8962) );
  INV_X1 U7996 ( .A(n8962), .ZN(n6858) );
  INV_X1 U7997 ( .A(n8913), .ZN(n8918) );
  NAND2_X1 U7998 ( .A1(n6861), .A2(n8964), .ZN(n8312) );
  NAND2_X1 U7999 ( .A1(n8312), .A2(n8890), .ZN(n8311) );
  NOR2_X1 U8000 ( .A1(n8715), .A2(n8698), .ZN(n8973) );
  INV_X1 U8001 ( .A(n8973), .ZN(n6863) );
  NAND2_X1 U8002 ( .A1(n8390), .A2(n6863), .ZN(n6864) );
  NAND2_X1 U8003 ( .A1(n8715), .A2(n8698), .ZN(n8971) );
  NAND2_X1 U8004 ( .A1(n6864), .A2(n8971), .ZN(n8692) );
  INV_X1 U8005 ( .A(n8974), .ZN(n8693) );
  NAND2_X1 U8006 ( .A1(n8692), .A2(n8693), .ZN(n6865) );
  NAND2_X1 U8007 ( .A1(n6865), .A2(n8977), .ZN(n8672) );
  INV_X1 U8008 ( .A(n9279), .ZN(n9081) );
  NAND2_X1 U8009 ( .A1(n8728), .A2(n9081), .ZN(n6866) );
  NAND2_X1 U8010 ( .A1(n9602), .A2(n9516), .ZN(n6867) );
  NAND2_X1 U8011 ( .A1(n9524), .A2(n9604), .ZN(n9009) );
  INV_X1 U8012 ( .A(n9468), .ZN(n9500) );
  NAND2_X1 U8013 ( .A1(n9586), .A2(n9500), .ZN(n9476) );
  AND2_X1 U8014 ( .A1(n9478), .A2(n9476), .ZN(n6868) );
  XNOR2_X1 U8015 ( .A(n9572), .B(n9276), .ZN(n9444) );
  INV_X1 U8016 ( .A(n9444), .ZN(n9453) );
  NAND2_X1 U8017 ( .A1(n9215), .A2(n9165), .ZN(n9038) );
  INV_X1 U8018 ( .A(n8872), .ZN(n9039) );
  NAND2_X1 U8019 ( .A1(n9564), .A2(n9438), .ZN(n8871) );
  INV_X1 U8020 ( .A(n8871), .ZN(n9044) );
  NAND2_X1 U8021 ( .A1(n9252), .A2(n9245), .ZN(n9047) );
  NAND2_X1 U8022 ( .A1(n6912), .A2(n9047), .ZN(n9410) );
  INV_X1 U8023 ( .A(n8870), .ZN(n9048) );
  INV_X1 U8024 ( .A(n9409), .ZN(n6913) );
  NOR2_X1 U8025 ( .A1(n9048), .A2(n6913), .ZN(n6869) );
  NAND2_X1 U8026 ( .A1(n9555), .A2(n6814), .ZN(n8869) );
  INV_X1 U8027 ( .A(n8869), .ZN(n9049) );
  INV_X1 U8028 ( .A(n9116), .ZN(n8904) );
  XNOR2_X1 U8029 ( .A(n6919), .B(n8904), .ZN(n9142) );
  AND2_X1 U8030 ( .A1(n9078), .A2(n8090), .ZN(n6901) );
  INV_X1 U8031 ( .A(n9078), .ZN(n8346) );
  OAI21_X1 U8032 ( .B1(n6904), .B2(n6901), .A(n9618), .ZN(n6870) );
  OR2_X1 U8033 ( .A1(n9150), .A2(n6870), .ZN(n7775) );
  NAND2_X1 U8034 ( .A1(n9070), .A2(n9073), .ZN(n7498) );
  NAND2_X1 U8035 ( .A1(n9147), .A2(n6871), .ZN(n7344) );
  NAND2_X1 U8036 ( .A1(n6873), .A2(n6874), .ZN(n6881) );
  OAI21_X1 U8037 ( .B1(P2_IR_REG_25__SCAN_IN), .B2(P2_IR_REG_24__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n6877) );
  NAND2_X1 U8038 ( .A1(n6878), .A2(n6877), .ZN(n6880) );
  NAND2_X1 U8039 ( .A1(n7470), .A2(n6881), .ZN(n6882) );
  OR2_X1 U8040 ( .A1(n6884), .A2(P2_D_REG_1__SCAN_IN), .ZN(n6887) );
  NAND2_X1 U8041 ( .A1(n6885), .A2(n7470), .ZN(n6886) );
  INV_X1 U8042 ( .A(n7339), .ZN(n9660) );
  AND2_X1 U8043 ( .A1(n7500), .A2(n9660), .ZN(n7335) );
  NOR2_X1 U8044 ( .A1(P2_D_REG_31__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .ZN(
        n6891) );
  NOR4_X1 U8045 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_29__SCAN_IN), .A4(P2_D_REG_28__SCAN_IN), .ZN(n6890) );
  NOR4_X1 U8046 ( .A1(P2_D_REG_23__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .A3(
        P2_D_REG_21__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n6889) );
  NOR4_X1 U8047 ( .A1(P2_D_REG_27__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_25__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n6888) );
  NAND4_X1 U8048 ( .A1(n6891), .A2(n6890), .A3(n6889), .A4(n6888), .ZN(n6897)
         );
  NOR4_X1 U8049 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n6895) );
  NOR4_X1 U8050 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_18__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n6894) );
  NOR4_X1 U8051 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n6893) );
  NOR4_X1 U8052 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n6892) );
  NAND4_X1 U8053 ( .A1(n6895), .A2(n6894), .A3(n6893), .A4(n6892), .ZN(n6896)
         );
  NOR2_X1 U8054 ( .A1(n6897), .A2(n6896), .ZN(n6898) );
  NAND2_X1 U8055 ( .A1(n5024), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6899) );
  NAND2_X1 U8056 ( .A1(n7338), .A2(n9659), .ZN(n6900) );
  OAI21_X1 U8057 ( .B1(n7498), .B2(n9618), .A(n7500), .ZN(n6905) );
  INV_X1 U8058 ( .A(n6901), .ZN(n6902) );
  NOR2_X1 U8059 ( .A1(n6902), .A2(n9070), .ZN(n6903) );
  NAND2_X1 U8060 ( .A1(n6937), .A2(n7489), .ZN(n6936) );
  AOI22_X1 U8061 ( .A1(n6905), .A2(n6936), .B1(n7339), .B2(n6937), .ZN(n6906)
         );
  NOR2_X1 U8062 ( .A1(n9627), .A2(n6908), .ZN(n6909) );
  OAI211_X1 U8063 ( .C1(n6912), .C2(n6913), .A(n8869), .B(n9047), .ZN(n6914)
         );
  NAND2_X1 U8064 ( .A1(n6914), .A2(n8870), .ZN(n6917) );
  INV_X1 U8065 ( .A(n6915), .ZN(n6916) );
  INV_X1 U8066 ( .A(n8861), .ZN(n6925) );
  NAND2_X1 U8067 ( .A1(n9666), .A2(n8849), .ZN(n6921) );
  NAND2_X1 U8068 ( .A1(n8844), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n6920) );
  NAND2_X1 U8069 ( .A1(n6923), .A2(n6922), .ZN(n8858) );
  INV_X1 U8070 ( .A(n8858), .ZN(n6924) );
  MUX2_X2 U8071 ( .A(n6926), .B(n6925), .S(n6928), .Z(n8840) );
  OR2_X1 U8072 ( .A1(n8927), .A2(n7498), .ZN(n7774) );
  NAND2_X1 U8073 ( .A1(n6929), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n6932) );
  NAND2_X1 U8074 ( .A1(n8851), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n6931) );
  NAND2_X1 U8075 ( .A1(n8852), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n6930) );
  AND3_X1 U8076 ( .A1(n6932), .A2(n6931), .A3(n6930), .ZN(n6933) );
  NAND2_X1 U8077 ( .A1(n8857), .A2(n6933), .ZN(n9272) );
  INV_X1 U8078 ( .A(n9272), .ZN(n8862) );
  NAND2_X1 U8079 ( .A1(n6515), .A2(P2_B_REG_SCAN_IN), .ZN(n6934) );
  NAND2_X1 U8080 ( .A1(n9609), .A2(n6934), .ZN(n9398) );
  OAI22_X1 U8081 ( .A1(n9408), .A2(n9515), .B1(n8862), .B2(n9398), .ZN(n6935)
         );
  OAI21_X1 U8082 ( .B1(n8840), .B2(n7774), .A(n8843), .ZN(n6941) );
  AOI22_X1 U8083 ( .A1(n6883), .A2(n6937), .B1(n7339), .B2(n6936), .ZN(n6938)
         );
  NAND2_X1 U8084 ( .A1(n6939), .A2(n6938), .ZN(n9149) );
  INV_X1 U8085 ( .A(n9659), .ZN(n6940) );
  NAND2_X1 U8086 ( .A1(n6941), .A2(n10641), .ZN(n6946) );
  INV_X2 U8087 ( .A(n10641), .ZN(n10687) );
  NOR2_X1 U8088 ( .A1(n6942), .A2(n10677), .ZN(n9400) );
  AOI21_X1 U8089 ( .B1(n10687), .B2(P2_REG2_REG_29__SCAN_IN), .A(n9400), .ZN(
        n6943) );
  INV_X1 U8090 ( .A(n6944), .ZN(n6945) );
  NAND2_X1 U8091 ( .A1(n6946), .A2(n6945), .ZN(P2_U3204) );
  INV_X1 U8092 ( .A(n7854), .ZN(n6947) );
  NAND2_X1 U8093 ( .A1(n7932), .A2(n7018), .ZN(n6953) );
  NAND2_X1 U8094 ( .A1(n6948), .A2(n7854), .ZN(n6950) );
  NAND2_X1 U8095 ( .A1(n6950), .A2(n6949), .ZN(n6952) );
  NAND2_X2 U8096 ( .A1(n6952), .A2(n6951), .ZN(n6981) );
  INV_X1 U8097 ( .A(n6951), .ZN(n6955) );
  NAND2_X1 U8098 ( .A1(n6955), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6954) );
  NAND2_X1 U8099 ( .A1(n7932), .A2(n7163), .ZN(n6957) );
  AOI22_X1 U8100 ( .A1(n7831), .A2(n7018), .B1(n6955), .B2(
        P1_IR_REG_0__SCAN_IN), .ZN(n6956) );
  NAND2_X1 U8101 ( .A1(n6957), .A2(n6956), .ZN(n7685) );
  NAND2_X1 U8102 ( .A1(n6958), .A2(n7166), .ZN(n6959) );
  NAND2_X1 U8103 ( .A1(n7684), .A2(n6959), .ZN(n7692) );
  NAND2_X1 U8104 ( .A1(n6960), .A2(n7018), .ZN(n6962) );
  NAND2_X1 U8105 ( .A1(n7861), .A2(n6983), .ZN(n6961) );
  NAND2_X1 U8106 ( .A1(n6962), .A2(n6961), .ZN(n6964) );
  XNOR2_X1 U8107 ( .A(n6964), .B(n6963), .ZN(n7691) );
  NAND2_X1 U8108 ( .A1(n6960), .A2(n7163), .ZN(n6967) );
  OR2_X1 U8109 ( .A1(n6965), .A2(n7170), .ZN(n6966) );
  NAND2_X1 U8110 ( .A1(n6967), .A2(n6966), .ZN(n7696) );
  NAND2_X1 U8111 ( .A1(n7692), .A2(n7691), .ZN(n7695) );
  INV_X1 U8112 ( .A(n6983), .ZN(n7154) );
  NAND2_X1 U8113 ( .A1(n6970), .A2(n7018), .ZN(n6968) );
  NAND2_X1 U8114 ( .A1(n4997), .A2(n6968), .ZN(n6969) );
  XNOR2_X1 U8115 ( .A(n6969), .B(n7166), .ZN(n6977) );
  INV_X1 U8116 ( .A(n6977), .ZN(n6975) );
  NAND2_X1 U8117 ( .A1(n6970), .A2(n7163), .ZN(n6973) );
  OR2_X1 U8118 ( .A1(n6971), .A2(n7170), .ZN(n6972) );
  AND2_X1 U8119 ( .A1(n6973), .A2(n6972), .ZN(n6976) );
  INV_X1 U8120 ( .A(n6976), .ZN(n6974) );
  NAND2_X1 U8121 ( .A1(n6975), .A2(n6974), .ZN(n6978) );
  NAND2_X1 U8122 ( .A1(n6977), .A2(n6976), .ZN(n6979) );
  NAND2_X1 U8123 ( .A1(n9761), .A2(n9763), .ZN(n9762) );
  OAI22_X1 U8124 ( .A1(n6982), .A2(n7170), .B1(n10593), .B2(n7154), .ZN(n6980)
         );
  XNOR2_X1 U8125 ( .A(n6980), .B(n7166), .ZN(n6990) );
  OAI22_X1 U8126 ( .A1(n6982), .A2(n6981), .B1(n10593), .B2(n7170), .ZN(n6988)
         );
  XNOR2_X1 U8127 ( .A(n6990), .B(n6988), .ZN(n7811) );
  NAND2_X1 U8128 ( .A1(n6987), .A2(n7018), .ZN(n6985) );
  NAND2_X1 U8129 ( .A1(n8022), .A2(n7168), .ZN(n6984) );
  NAND2_X1 U8130 ( .A1(n6985), .A2(n6984), .ZN(n6986) );
  AOI22_X1 U8131 ( .A1(n6987), .A2(n7163), .B1(n7018), .B2(n8022), .ZN(n6991)
         );
  XNOR2_X1 U8132 ( .A(n6993), .B(n6991), .ZN(n7836) );
  INV_X1 U8133 ( .A(n6988), .ZN(n6989) );
  NAND2_X1 U8134 ( .A1(n6990), .A2(n6989), .ZN(n7837) );
  INV_X1 U8135 ( .A(n6991), .ZN(n6992) );
  NAND2_X1 U8136 ( .A1(n6993), .A2(n6992), .ZN(n6994) );
  OAI22_X1 U8137 ( .A1(n8030), .A2(n7170), .B1(n10613), .B2(n7154), .ZN(n6995)
         );
  XNOR2_X1 U8138 ( .A(n6995), .B(n7166), .ZN(n7922) );
  AND2_X1 U8139 ( .A1(n7928), .A2(n7018), .ZN(n6996) );
  AOI21_X1 U8140 ( .B1(n9808), .B2(n7163), .A(n6996), .ZN(n6999) );
  NAND2_X1 U8141 ( .A1(n7922), .A2(n6999), .ZN(n6997) );
  OAI22_X1 U8142 ( .A1(n8136), .A2(n7170), .B1(n10623), .B2(n7154), .ZN(n6998)
         );
  XNOR2_X1 U8143 ( .A(n6998), .B(n6963), .ZN(n7003) );
  OAI22_X1 U8144 ( .A1(n8136), .A2(n6981), .B1(n10623), .B2(n7170), .ZN(n7004)
         );
  AND2_X1 U8145 ( .A1(n7003), .A2(n7004), .ZN(n8050) );
  INV_X1 U8146 ( .A(n8050), .ZN(n7001) );
  INV_X1 U8147 ( .A(n7922), .ZN(n7000) );
  INV_X1 U8148 ( .A(n6999), .ZN(n7921) );
  NAND2_X1 U8149 ( .A1(n7000), .A2(n7921), .ZN(n8047) );
  AND2_X1 U8150 ( .A1(n7001), .A2(n8047), .ZN(n7002) );
  INV_X1 U8151 ( .A(n7003), .ZN(n7006) );
  INV_X1 U8152 ( .A(n7004), .ZN(n7005) );
  NAND2_X1 U8153 ( .A1(n7006), .A2(n7005), .ZN(n8049) );
  NAND2_X1 U8154 ( .A1(n8271), .A2(n7168), .ZN(n7007) );
  OAI21_X1 U8155 ( .B1(n8029), .B2(n7170), .A(n7007), .ZN(n7008) );
  XNOR2_X1 U8156 ( .A(n7008), .B(n6963), .ZN(n7009) );
  AOI22_X1 U8157 ( .A1(n9806), .A2(n7163), .B1(n7140), .B2(n8271), .ZN(n7010)
         );
  XNOR2_X1 U8158 ( .A(n7009), .B(n7010), .ZN(n8150) );
  INV_X1 U8159 ( .A(n7009), .ZN(n7011) );
  NAND2_X1 U8160 ( .A1(n7011), .A2(n7010), .ZN(n7012) );
  NAND2_X1 U8161 ( .A1(n8167), .A2(n7168), .ZN(n7014) );
  NAND2_X1 U8162 ( .A1(n8286), .A2(n7140), .ZN(n7013) );
  NAND2_X1 U8163 ( .A1(n7014), .A2(n7013), .ZN(n7015) );
  XNOR2_X1 U8164 ( .A(n7015), .B(n7166), .ZN(n8161) );
  AOI22_X1 U8165 ( .A1(n8167), .A2(n7140), .B1(n8286), .B2(n7163), .ZN(n8160)
         );
  NAND2_X1 U8166 ( .A1(n8159), .A2(n8161), .ZN(n7016) );
  NAND2_X1 U8167 ( .A1(n7017), .A2(n7016), .ZN(n8282) );
  NAND2_X1 U8168 ( .A1(n5757), .A2(n7168), .ZN(n7020) );
  NAND2_X1 U8169 ( .A1(n5343), .A2(n7140), .ZN(n7019) );
  NAND2_X1 U8170 ( .A1(n7020), .A2(n7019), .ZN(n7021) );
  XNOR2_X1 U8171 ( .A(n7021), .B(n7166), .ZN(n8284) );
  NOR2_X1 U8172 ( .A1(n8246), .A2(n6981), .ZN(n7022) );
  AOI21_X1 U8173 ( .B1(n5757), .B2(n7140), .A(n7022), .ZN(n8283) );
  AND2_X1 U8174 ( .A1(n8284), .A2(n8283), .ZN(n7026) );
  INV_X1 U8175 ( .A(n8284), .ZN(n7024) );
  INV_X1 U8176 ( .A(n8283), .ZN(n7023) );
  NAND2_X1 U8177 ( .A1(n7024), .A2(n7023), .ZN(n7025) );
  NAND2_X1 U8178 ( .A1(n4944), .A2(n7140), .ZN(n7028) );
  NAND2_X1 U8179 ( .A1(n9805), .A2(n7163), .ZN(n7027) );
  NAND2_X1 U8180 ( .A1(n7028), .A2(n7027), .ZN(n8336) );
  NAND2_X1 U8181 ( .A1(n4944), .A2(n7168), .ZN(n7030) );
  NAND2_X1 U8182 ( .A1(n9805), .A2(n7140), .ZN(n7029) );
  NAND2_X1 U8183 ( .A1(n7030), .A2(n7029), .ZN(n7031) );
  XNOR2_X1 U8184 ( .A(n7031), .B(n6963), .ZN(n8335) );
  NAND2_X1 U8185 ( .A1(n8771), .A2(n7168), .ZN(n7033) );
  NAND2_X1 U8186 ( .A1(n9804), .A2(n7140), .ZN(n7032) );
  NAND2_X1 U8187 ( .A1(n7033), .A2(n7032), .ZN(n7034) );
  XNOR2_X1 U8188 ( .A(n7034), .B(n7166), .ZN(n7040) );
  NOR2_X1 U8189 ( .A1(n8706), .A2(n6981), .ZN(n7035) );
  AOI21_X1 U8190 ( .B1(n8771), .B2(n7140), .A(n7035), .ZN(n7041) );
  NAND2_X1 U8191 ( .A1(n7040), .A2(n7041), .ZN(n8765) );
  NAND2_X1 U8192 ( .A1(n8665), .A2(n7168), .ZN(n7037) );
  NAND2_X1 U8193 ( .A1(n9803), .A2(n7140), .ZN(n7036) );
  NAND2_X1 U8194 ( .A1(n7037), .A2(n7036), .ZN(n7038) );
  XNOR2_X1 U8195 ( .A(n7038), .B(n6963), .ZN(n7048) );
  AND2_X1 U8196 ( .A1(n9803), .A2(n7163), .ZN(n7039) );
  AOI21_X1 U8197 ( .B1(n8665), .B2(n7140), .A(n7039), .ZN(n7049) );
  XNOR2_X1 U8198 ( .A(n7048), .B(n7049), .ZN(n8702) );
  INV_X1 U8199 ( .A(n7040), .ZN(n7043) );
  INV_X1 U8200 ( .A(n7041), .ZN(n7042) );
  NAND2_X1 U8201 ( .A1(n7043), .A2(n7042), .ZN(n8767) );
  NAND2_X1 U8202 ( .A1(n10235), .A2(n7168), .ZN(n7045) );
  NAND2_X1 U8203 ( .A1(n9802), .A2(n7140), .ZN(n7044) );
  NAND2_X1 U8204 ( .A1(n7045), .A2(n7044), .ZN(n7046) );
  XNOR2_X1 U8205 ( .A(n7046), .B(n6963), .ZN(n7054) );
  AND2_X1 U8206 ( .A1(n9802), .A2(n7163), .ZN(n7047) );
  AOI21_X1 U8207 ( .B1(n10235), .B2(n7140), .A(n7047), .ZN(n7052) );
  XNOR2_X1 U8208 ( .A(n7054), .B(n7052), .ZN(n8736) );
  INV_X1 U8209 ( .A(n7048), .ZN(n7050) );
  NAND2_X1 U8210 ( .A1(n7050), .A2(n7049), .ZN(n8734) );
  AND2_X1 U8211 ( .A1(n8736), .A2(n8734), .ZN(n7051) );
  INV_X1 U8212 ( .A(n7052), .ZN(n7053) );
  NAND2_X1 U8213 ( .A1(n7054), .A2(n7053), .ZN(n7055) );
  NAND2_X1 U8214 ( .A1(n8735), .A2(n7055), .ZN(n7060) );
  NAND2_X1 U8215 ( .A1(n10230), .A2(n7168), .ZN(n7057) );
  NAND2_X1 U8216 ( .A1(n9801), .A2(n7140), .ZN(n7056) );
  NAND2_X1 U8217 ( .A1(n7057), .A2(n7056), .ZN(n7058) );
  XNOR2_X1 U8218 ( .A(n7058), .B(n6963), .ZN(n7061) );
  AND2_X1 U8219 ( .A1(n9801), .A2(n7163), .ZN(n7059) );
  INV_X1 U8220 ( .A(n7061), .ZN(n7062) );
  NAND2_X1 U8221 ( .A1(n10225), .A2(n7168), .ZN(n7064) );
  NAND2_X1 U8222 ( .A1(n9800), .A2(n7140), .ZN(n7063) );
  NAND2_X1 U8223 ( .A1(n7064), .A2(n7063), .ZN(n7065) );
  NAND2_X1 U8224 ( .A1(n10225), .A2(n7140), .ZN(n7067) );
  NAND2_X1 U8225 ( .A1(n9800), .A2(n7163), .ZN(n7066) );
  NAND2_X1 U8226 ( .A1(n7067), .A2(n7066), .ZN(n8827) );
  INV_X1 U8227 ( .A(n8826), .ZN(n7068) );
  NAND2_X1 U8228 ( .A1(n10222), .A2(n7168), .ZN(n7070) );
  NAND2_X1 U8229 ( .A1(n9723), .A2(n7140), .ZN(n7069) );
  NAND2_X1 U8230 ( .A1(n7070), .A2(n7069), .ZN(n7071) );
  XNOR2_X1 U8231 ( .A(n7071), .B(n7166), .ZN(n7073) );
  NOR2_X1 U8232 ( .A1(n10125), .A2(n6981), .ZN(n7072) );
  AOI21_X1 U8233 ( .B1(n10222), .B2(n7140), .A(n7072), .ZN(n7074) );
  NAND2_X1 U8234 ( .A1(n7073), .A2(n7074), .ZN(n7080) );
  INV_X1 U8235 ( .A(n7073), .ZN(n7076) );
  INV_X1 U8236 ( .A(n7074), .ZN(n7075) );
  NAND2_X1 U8237 ( .A1(n7076), .A2(n7075), .ZN(n7077) );
  NAND2_X1 U8238 ( .A1(n7080), .A2(n7077), .ZN(n9714) );
  NAND2_X1 U8239 ( .A1(n7079), .A2(n7078), .ZN(n9712) );
  NAND2_X1 U8240 ( .A1(n10131), .A2(n7168), .ZN(n7082) );
  INV_X1 U8241 ( .A(n10144), .ZN(n9773) );
  NAND2_X1 U8242 ( .A1(n9773), .A2(n7140), .ZN(n7081) );
  NAND2_X1 U8243 ( .A1(n7082), .A2(n7081), .ZN(n7083) );
  XNOR2_X1 U8244 ( .A(n7083), .B(n6963), .ZN(n7086) );
  NAND2_X1 U8245 ( .A1(n10131), .A2(n7140), .ZN(n7085) );
  NAND2_X1 U8246 ( .A1(n9773), .A2(n7163), .ZN(n7084) );
  NAND2_X1 U8247 ( .A1(n7085), .A2(n7084), .ZN(n7087) );
  NAND2_X1 U8248 ( .A1(n7086), .A2(n7087), .ZN(n9720) );
  INV_X1 U8249 ( .A(n7086), .ZN(n7089) );
  INV_X1 U8250 ( .A(n7087), .ZN(n7088) );
  NAND2_X1 U8251 ( .A1(n7089), .A2(n7088), .ZN(n9722) );
  NAND2_X1 U8252 ( .A1(n10210), .A2(n7168), .ZN(n7091) );
  NAND2_X1 U8253 ( .A1(n9799), .A2(n7140), .ZN(n7090) );
  NAND2_X1 U8254 ( .A1(n7091), .A2(n7090), .ZN(n7092) );
  NAND2_X1 U8255 ( .A1(n10210), .A2(n7140), .ZN(n7094) );
  NAND2_X1 U8256 ( .A1(n9799), .A2(n7163), .ZN(n7093) );
  NAND2_X1 U8257 ( .A1(n7094), .A2(n7093), .ZN(n9772) );
  NAND2_X1 U8258 ( .A1(n10102), .A2(n7168), .ZN(n7098) );
  OR2_X1 U8259 ( .A1(n10111), .A2(n7170), .ZN(n7097) );
  NAND2_X1 U8260 ( .A1(n7098), .A2(n7097), .ZN(n7099) );
  XNOR2_X1 U8261 ( .A(n7099), .B(n7166), .ZN(n7103) );
  NOR2_X1 U8262 ( .A1(n10111), .A2(n6981), .ZN(n7100) );
  AOI21_X1 U8263 ( .B1(n10102), .B2(n7140), .A(n7100), .ZN(n7102) );
  XNOR2_X1 U8264 ( .A(n7103), .B(n7102), .ZN(n9689) );
  INV_X1 U8265 ( .A(n9689), .ZN(n7101) );
  NAND2_X1 U8266 ( .A1(n7103), .A2(n7102), .ZN(n7104) );
  NAND2_X1 U8267 ( .A1(n10200), .A2(n7168), .ZN(n7106) );
  NAND2_X1 U8268 ( .A1(n9698), .A2(n7140), .ZN(n7105) );
  NAND2_X1 U8269 ( .A1(n7106), .A2(n7105), .ZN(n7107) );
  XNOR2_X1 U8270 ( .A(n7107), .B(n6963), .ZN(n7109) );
  NOR2_X1 U8271 ( .A1(n10097), .A2(n6981), .ZN(n7108) );
  AOI21_X1 U8272 ( .B1(n10200), .B2(n7140), .A(n7108), .ZN(n7110) );
  XNOR2_X1 U8273 ( .A(n7109), .B(n7110), .ZN(n9739) );
  INV_X1 U8274 ( .A(n7109), .ZN(n7111) );
  NAND2_X1 U8275 ( .A1(n10070), .A2(n7168), .ZN(n7113) );
  NAND2_X1 U8276 ( .A1(n10048), .A2(n7140), .ZN(n7112) );
  NAND2_X1 U8277 ( .A1(n7113), .A2(n7112), .ZN(n7114) );
  XNOR2_X1 U8278 ( .A(n7114), .B(n7166), .ZN(n7120) );
  NOR2_X1 U8279 ( .A1(n10081), .A2(n6981), .ZN(n7115) );
  AOI21_X1 U8280 ( .B1(n10070), .B2(n7140), .A(n7115), .ZN(n7121) );
  XNOR2_X1 U8281 ( .A(n7120), .B(n7121), .ZN(n9695) );
  NAND2_X1 U8282 ( .A1(n10190), .A2(n7168), .ZN(n7117) );
  NAND2_X1 U8283 ( .A1(n9798), .A2(n7140), .ZN(n7116) );
  NAND2_X1 U8284 ( .A1(n7117), .A2(n7116), .ZN(n7118) );
  XOR2_X1 U8285 ( .A(n7118), .B(n6963), .Z(n7129) );
  OR2_X1 U8286 ( .A1(n9695), .A2(n7129), .ZN(n7119) );
  NOR2_X1 U8287 ( .A1(n9694), .A2(n7119), .ZN(n7124) );
  INV_X1 U8288 ( .A(n7120), .ZN(n7123) );
  INV_X1 U8289 ( .A(n7121), .ZN(n7122) );
  NAND2_X1 U8290 ( .A1(n7123), .A2(n7122), .ZN(n7128) );
  NOR2_X1 U8291 ( .A1(n7124), .A2(n4980), .ZN(n9748) );
  NOR2_X1 U8292 ( .A1(n10065), .A2(n6981), .ZN(n7125) );
  AOI21_X1 U8293 ( .B1(n10190), .B2(n7018), .A(n7125), .ZN(n9747) );
  INV_X1 U8294 ( .A(n9694), .ZN(n7127) );
  INV_X1 U8295 ( .A(n9695), .ZN(n7126) );
  NAND2_X1 U8296 ( .A1(n7127), .A2(n7126), .ZN(n9696) );
  NAND2_X1 U8297 ( .A1(n6101), .A2(n7168), .ZN(n7131) );
  NAND2_X1 U8298 ( .A1(n10047), .A2(n7140), .ZN(n7130) );
  NAND2_X1 U8299 ( .A1(n7131), .A2(n7130), .ZN(n7132) );
  XNOR2_X1 U8300 ( .A(n7132), .B(n6963), .ZN(n7134) );
  OAI22_X1 U8301 ( .A1(n10037), .A2(n7170), .B1(n9753), .B2(n6981), .ZN(n7133)
         );
  XNOR2_X1 U8302 ( .A(n7134), .B(n7133), .ZN(n9679) );
  AOI22_X1 U8303 ( .A1(n10181), .A2(n7168), .B1(n7140), .B2(n9706), .ZN(n7135)
         );
  XOR2_X1 U8304 ( .A(n6963), .B(n7135), .Z(n7137) );
  INV_X1 U8305 ( .A(n10181), .ZN(n10022) );
  OAI22_X1 U8306 ( .A1(n10022), .A2(n7170), .B1(n10031), .B2(n6981), .ZN(n7136) );
  NAND2_X1 U8307 ( .A1(n7137), .A2(n7136), .ZN(n9728) );
  AOI22_X1 U8308 ( .A1(n10174), .A2(n7168), .B1(n7140), .B2(n10015), .ZN(n7138) );
  XNOR2_X1 U8309 ( .A(n7138), .B(n6963), .ZN(n7145) );
  AND2_X1 U8310 ( .A1(n10015), .A2(n7163), .ZN(n7139) );
  AOI21_X1 U8311 ( .B1(n10174), .B2(n7018), .A(n7139), .ZN(n7146) );
  XNOR2_X1 U8312 ( .A(n7145), .B(n7146), .ZN(n9703) );
  NAND2_X1 U8313 ( .A1(n10249), .A2(n7168), .ZN(n7142) );
  NAND2_X1 U8314 ( .A1(n9797), .A2(n7140), .ZN(n7141) );
  NAND2_X1 U8315 ( .A1(n7142), .A2(n7141), .ZN(n7143) );
  XNOR2_X1 U8316 ( .A(n7143), .B(n7166), .ZN(n7150) );
  NOR2_X1 U8317 ( .A1(n9996), .A2(n6981), .ZN(n7144) );
  AOI21_X1 U8318 ( .B1(n10249), .B2(n7018), .A(n7144), .ZN(n7151) );
  XNOR2_X1 U8319 ( .A(n7150), .B(n7151), .ZN(n9781) );
  INV_X1 U8320 ( .A(n7145), .ZN(n7148) );
  INV_X1 U8321 ( .A(n7146), .ZN(n7147) );
  NOR2_X1 U8322 ( .A1(n7148), .A2(n7147), .ZN(n9782) );
  INV_X1 U8323 ( .A(n7150), .ZN(n7153) );
  INV_X1 U8324 ( .A(n7151), .ZN(n7152) );
  OAI22_X1 U8325 ( .A1(n9969), .A2(n7154), .B1(n9984), .B2(n7170), .ZN(n7155)
         );
  XOR2_X1 U8326 ( .A(n6963), .B(n7155), .Z(n7157) );
  INV_X1 U8327 ( .A(n9984), .ZN(n9796) );
  AOI22_X1 U8328 ( .A1(n7329), .A2(n7140), .B1(n7163), .B2(n9796), .ZN(n7156)
         );
  NAND2_X1 U8329 ( .A1(n7157), .A2(n7156), .ZN(n7193) );
  OAI21_X1 U8330 ( .B1(n7157), .B2(n7156), .A(n7193), .ZN(n7325) );
  INV_X1 U8331 ( .A(n7158), .ZN(n7160) );
  OR2_X1 U8332 ( .A1(n7160), .A2(n7159), .ZN(n7819) );
  AND2_X1 U8333 ( .A1(n7183), .A2(n10274), .ZN(n7175) );
  NOR2_X1 U8334 ( .A1(n10649), .A2(n7398), .ZN(n7162) );
  NAND2_X1 U8335 ( .A1(n7366), .A2(n7140), .ZN(n7165) );
  NAND2_X1 U8336 ( .A1(n9795), .A2(n7163), .ZN(n7164) );
  NAND2_X1 U8337 ( .A1(n7165), .A2(n7164), .ZN(n7167) );
  XNOR2_X1 U8338 ( .A(n7167), .B(n7166), .ZN(n7172) );
  NAND2_X1 U8339 ( .A1(n7366), .A2(n7168), .ZN(n7169) );
  OAI21_X1 U8340 ( .B1(n9942), .B2(n7170), .A(n7169), .ZN(n7171) );
  XNOR2_X1 U8341 ( .A(n7172), .B(n7171), .ZN(n7174) );
  INV_X1 U8342 ( .A(n7174), .ZN(n7192) );
  NAND3_X1 U8343 ( .A1(n7193), .A2(n9784), .A3(n7192), .ZN(n7173) );
  NAND3_X1 U8344 ( .A1(n7328), .A2(n7174), .A3(n9784), .ZN(n7197) );
  INV_X1 U8345 ( .A(n7175), .ZN(n7177) );
  OR2_X1 U8346 ( .A1(n7654), .A2(n7176), .ZN(n7829) );
  OR2_X1 U8347 ( .A1(n7177), .A2(n7829), .ZN(n7180) );
  INV_X1 U8348 ( .A(n7178), .ZN(n7179) );
  AND2_X1 U8349 ( .A1(n7183), .A2(n7181), .ZN(n7182) );
  AOI22_X1 U8350 ( .A1(n9786), .A2(n9796), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3086), .ZN(n7191) );
  INV_X1 U8351 ( .A(n7183), .ZN(n7186) );
  NAND2_X1 U8352 ( .A1(n7184), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8172) );
  NAND2_X1 U8353 ( .A1(n10649), .A2(n8172), .ZN(n7185) );
  NAND2_X1 U8354 ( .A1(n7186), .A2(n7185), .ZN(n7189) );
  AND3_X1 U8355 ( .A1(n6951), .A2(n7397), .A3(n7187), .ZN(n7188) );
  NAND2_X1 U8356 ( .A1(n7189), .A2(n7188), .ZN(n7688) );
  NAND2_X1 U8357 ( .A1(n9788), .A2(n9957), .ZN(n7190) );
  OAI211_X1 U8358 ( .C1(n9775), .C2(n8281), .A(n7191), .B(n7190), .ZN(n7195)
         );
  NOR3_X1 U8359 ( .A1(n7193), .A2(n7192), .A3(n9778), .ZN(n7194) );
  AOI211_X1 U8360 ( .C1(n7366), .C2(n9789), .A(n7195), .B(n7194), .ZN(n7196)
         );
  NAND3_X1 U8361 ( .A1(n7198), .A2(n7197), .A3(n7196), .ZN(P1_U3220) );
  INV_X1 U8362 ( .A(n7468), .ZN(n7199) );
  NAND2_X1 U8363 ( .A1(n7491), .A2(n9053), .ZN(n7200) );
  NAND2_X1 U8364 ( .A1(n7200), .A2(n7490), .ZN(n7316) );
  NAND2_X1 U8365 ( .A1(n7316), .A2(n6515), .ZN(n7201) );
  NAND2_X1 U8366 ( .A1(n7201), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3150) );
  INV_X1 U8367 ( .A(n7582), .ZN(n7432) );
  INV_X1 U8368 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n7236) );
  NAND2_X1 U8369 ( .A1(n7236), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n7202) );
  NAND2_X1 U8370 ( .A1(n4968), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n7205) );
  NAND2_X1 U8371 ( .A1(n7204), .A2(n7205), .ZN(n7590) );
  INV_X1 U8372 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n7723) );
  XNOR2_X1 U8373 ( .A(n7582), .B(P2_REG1_REG_2__SCAN_IN), .ZN(n7564) );
  AOI22_X1 U8374 ( .A1(n10376), .A2(P2_REG1_REG_4__SCAN_IN), .B1(n7207), .B2(
        n7429), .ZN(n10378) );
  NOR2_X1 U8375 ( .A1(n10379), .A2(n10378), .ZN(n10377) );
  NOR2_X1 U8376 ( .A1(n7290), .A2(n7209), .ZN(n7211) );
  INV_X1 U8377 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n10402) );
  MUX2_X1 U8378 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n7965), .S(n10414), .Z(n10420) );
  INV_X1 U8379 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n10440) );
  NOR2_X1 U8380 ( .A1(n10431), .A2(n7213), .ZN(n7214) );
  NAND2_X1 U8381 ( .A1(P2_REG1_REG_8__SCAN_IN), .A2(n7457), .ZN(n7215) );
  OAI21_X1 U8382 ( .B1(n7457), .B2(P2_REG1_REG_8__SCAN_IN), .A(n7215), .ZN(
        n10457) );
  NOR2_X1 U8383 ( .A1(n10463), .A2(n7216), .ZN(n7217) );
  INV_X1 U8384 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n10472) );
  NAND2_X1 U8385 ( .A1(P2_REG1_REG_10__SCAN_IN), .A2(n7463), .ZN(n7218) );
  OAI21_X1 U8386 ( .B1(n7463), .B2(P2_REG1_REG_10__SCAN_IN), .A(n7218), .ZN(
        n10489) );
  NOR2_X1 U8387 ( .A1(n10496), .A2(n7219), .ZN(n7220) );
  INV_X1 U8388 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n10508) );
  NAND2_X1 U8389 ( .A1(P2_REG1_REG_12__SCAN_IN), .A2(n8638), .ZN(n7221) );
  OAI21_X1 U8390 ( .B1(P2_REG1_REG_12__SCAN_IN), .B2(n8638), .A(n7221), .ZN(
        n8627) );
  NOR2_X1 U8391 ( .A1(n7279), .A2(n7222), .ZN(n7223) );
  INV_X1 U8392 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n9295) );
  INV_X1 U8393 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n9626) );
  AOI22_X1 U8394 ( .A1(n7277), .A2(P2_REG1_REG_14__SCAN_IN), .B1(n9626), .B2(
        n9322), .ZN(n9311) );
  NOR2_X1 U8395 ( .A1(n7275), .A2(n7224), .ZN(n7225) );
  INV_X1 U8396 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n9329) );
  NAND2_X1 U8397 ( .A1(P2_REG1_REG_16__SCAN_IN), .A2(n9356), .ZN(n7226) );
  OAI21_X1 U8398 ( .B1(P2_REG1_REG_16__SCAN_IN), .B2(n9356), .A(n7226), .ZN(
        n9344) );
  NOR2_X1 U8399 ( .A1(n9345), .A2(n9344), .ZN(n9343) );
  NOR2_X1 U8400 ( .A1(n7272), .A2(n7227), .ZN(n7228) );
  INV_X1 U8401 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n9363) );
  INV_X1 U8402 ( .A(n7265), .ZN(n9391) );
  NAND2_X1 U8403 ( .A1(n9391), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n7229) );
  OAI21_X1 U8404 ( .B1(n9391), .B2(P2_REG1_REG_18__SCAN_IN), .A(n7229), .ZN(
        n9379) );
  INV_X1 U8405 ( .A(n7229), .ZN(n7230) );
  NOR2_X1 U8406 ( .A1(n9378), .A2(n7230), .ZN(n7231) );
  XNOR2_X1 U8407 ( .A(n8090), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n7269) );
  XNOR2_X1 U8408 ( .A(n7231), .B(n7269), .ZN(n7232) );
  NOR2_X1 U8409 ( .A1(n6845), .A2(P2_U3151), .ZN(n9670) );
  AND2_X1 U8410 ( .A1(n9670), .A2(n7316), .ZN(n10355) );
  NAND2_X1 U8411 ( .A1(n7232), .A2(n10370), .ZN(n7323) );
  INV_X1 U8412 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n7233) );
  MUX2_X1 U8413 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n7233), .S(n9073), .Z(n7270)
         );
  INV_X1 U8414 ( .A(n7272), .ZN(n9373) );
  NAND2_X1 U8415 ( .A1(P2_REG2_REG_16__SCAN_IN), .A2(n9356), .ZN(n7262) );
  INV_X1 U8416 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n7234) );
  AOI22_X1 U8417 ( .A1(n7273), .A2(n7234), .B1(P2_REG2_REG_16__SCAN_IN), .B2(
        n9356), .ZN(n9348) );
  INV_X1 U8418 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n7259) );
  AOI22_X1 U8419 ( .A1(n7277), .A2(n7259), .B1(P2_REG2_REG_14__SCAN_IN), .B2(
        n9322), .ZN(n9314) );
  INV_X1 U8420 ( .A(n7279), .ZN(n9305) );
  NAND2_X1 U8421 ( .A1(P2_REG2_REG_12__SCAN_IN), .A2(n8638), .ZN(n7256) );
  INV_X1 U8422 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n8391) );
  AOI22_X1 U8423 ( .A1(P2_REG2_REG_12__SCAN_IN), .A2(n8638), .B1(n7281), .B2(
        n8391), .ZN(n8630) );
  INV_X1 U8424 ( .A(n10496), .ZN(n7482) );
  NAND2_X1 U8425 ( .A1(P2_REG2_REG_10__SCAN_IN), .A2(n7463), .ZN(n7253) );
  INV_X1 U8426 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7235) );
  AOI22_X1 U8427 ( .A1(n10479), .A2(n7235), .B1(P2_REG2_REG_10__SCAN_IN), .B2(
        n7463), .ZN(n10482) );
  INV_X1 U8428 ( .A(n10463), .ZN(n7460) );
  NAND2_X1 U8429 ( .A1(P2_REG2_REG_8__SCAN_IN), .A2(n7457), .ZN(n7250) );
  INV_X1 U8430 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n10640) );
  AOI22_X1 U8431 ( .A1(n10447), .A2(n10640), .B1(P2_REG2_REG_8__SCAN_IN), .B2(
        n7457), .ZN(n10450) );
  INV_X1 U8432 ( .A(n10431), .ZN(n7452) );
  INV_X1 U8433 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n7247) );
  AOI22_X1 U8434 ( .A1(n10414), .A2(n7247), .B1(P2_REG2_REG_6__SCAN_IN), .B2(
        n7441), .ZN(n10424) );
  INV_X1 U8435 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n7244) );
  AOI22_X1 U8436 ( .A1(n10376), .A2(n7244), .B1(P2_REG2_REG_4__SCAN_IN), .B2(
        n7429), .ZN(n10382) );
  INV_X1 U8437 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n7241) );
  MUX2_X1 U8438 ( .A(n7241), .B(P2_REG2_REG_2__SCAN_IN), .S(n7582), .Z(n7567)
         );
  AND2_X1 U8439 ( .A1(n4968), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n7238) );
  NAND2_X1 U8440 ( .A1(n7236), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n7237) );
  OAI22_X1 U8441 ( .A1(n7238), .A2(n7203), .B1(n4968), .B2(n7237), .ZN(n7589)
         );
  NAND2_X1 U8442 ( .A1(n7589), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n7240) );
  INV_X1 U8443 ( .A(n7238), .ZN(n7239) );
  NAND2_X1 U8444 ( .A1(n7240), .A2(n7239), .ZN(n7568) );
  NAND2_X1 U8445 ( .A1(n7567), .A2(n7568), .ZN(n7572) );
  OAI21_X1 U8446 ( .B1(n7582), .B2(n7241), .A(n7572), .ZN(n7242) );
  NAND2_X1 U8447 ( .A1(n7434), .A2(n7242), .ZN(n7243) );
  XOR2_X1 U8448 ( .A(n7242), .B(n7434), .Z(n10366) );
  NAND2_X1 U8449 ( .A1(P2_REG2_REG_3__SCAN_IN), .A2(n10366), .ZN(n10365) );
  NAND2_X1 U8450 ( .A1(n7243), .A2(n10365), .ZN(n10381) );
  NAND2_X1 U8451 ( .A1(n10382), .A2(n10381), .ZN(n10380) );
  OAI21_X1 U8452 ( .B1(n10376), .B2(n7244), .A(n10380), .ZN(n7245) );
  NAND2_X1 U8453 ( .A1(n10404), .A2(n7245), .ZN(n7246) );
  XNOR2_X1 U8454 ( .A(n7245), .B(n7290), .ZN(n10399) );
  NAND2_X1 U8455 ( .A1(P2_REG2_REG_5__SCAN_IN), .A2(n10399), .ZN(n10398) );
  NAND2_X1 U8456 ( .A1(n7452), .A2(n7248), .ZN(n7249) );
  NAND2_X1 U8457 ( .A1(P2_REG2_REG_7__SCAN_IN), .A2(n10433), .ZN(n10432) );
  NAND2_X1 U8458 ( .A1(n7460), .A2(n7251), .ZN(n7252) );
  NAND2_X1 U8459 ( .A1(P2_REG2_REG_9__SCAN_IN), .A2(n10465), .ZN(n10464) );
  NAND2_X1 U8460 ( .A1(n7252), .A2(n10464), .ZN(n10481) );
  NAND2_X1 U8461 ( .A1(n10482), .A2(n10481), .ZN(n10480) );
  NAND2_X1 U8462 ( .A1(n7253), .A2(n10480), .ZN(n7254) );
  NAND2_X1 U8463 ( .A1(n7482), .A2(n7254), .ZN(n7255) );
  XNOR2_X1 U8464 ( .A(n10496), .B(n7254), .ZN(n10499) );
  NAND2_X1 U8465 ( .A1(P2_REG2_REG_11__SCAN_IN), .A2(n10499), .ZN(n10498) );
  NAND2_X1 U8466 ( .A1(n9305), .A2(n7257), .ZN(n7258) );
  NAND2_X1 U8467 ( .A1(P2_REG2_REG_13__SCAN_IN), .A2(n9297), .ZN(n9296) );
  NAND2_X1 U8468 ( .A1(n5104), .A2(n7260), .ZN(n7261) );
  NAND2_X1 U8469 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n9331), .ZN(n9330) );
  NAND2_X1 U8470 ( .A1(n7261), .A2(n9330), .ZN(n9347) );
  NAND2_X1 U8471 ( .A1(n9348), .A2(n9347), .ZN(n9346) );
  NAND2_X1 U8472 ( .A1(n9373), .A2(n7263), .ZN(n7264) );
  INV_X1 U8473 ( .A(n9382), .ZN(n7266) );
  INV_X1 U8474 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n9380) );
  OAI21_X1 U8475 ( .B1(n7266), .B2(n9380), .A(n7265), .ZN(n7267) );
  OAI21_X1 U8476 ( .B1(P2_REG2_REG_18__SCAN_IN), .B2(n9382), .A(n7267), .ZN(
        n7268) );
  NAND2_X1 U8477 ( .A1(n10355), .A2(n7271), .ZN(n7566) );
  MUX2_X1 U8478 ( .A(n7270), .B(n7269), .S(n9074), .Z(n7315) );
  MUX2_X1 U8479 ( .A(P2_REG2_REG_17__SCAN_IN), .B(P2_REG1_REG_17__SCAN_IN), 
        .S(n9074), .Z(n7310) );
  XNOR2_X1 U8480 ( .A(n7272), .B(n7310), .ZN(n9368) );
  MUX2_X1 U8481 ( .A(P2_REG2_REG_16__SCAN_IN), .B(P2_REG1_REG_16__SCAN_IN), 
        .S(n9074), .Z(n7274) );
  OR2_X1 U8482 ( .A1(n7274), .A2(n9356), .ZN(n7309) );
  XNOR2_X1 U8483 ( .A(n7274), .B(n7273), .ZN(n9352) );
  MUX2_X1 U8484 ( .A(P2_REG2_REG_15__SCAN_IN), .B(P2_REG1_REG_15__SCAN_IN), 
        .S(n9074), .Z(n7276) );
  OR2_X1 U8485 ( .A1(n7276), .A2(n5104), .ZN(n7308) );
  XNOR2_X1 U8486 ( .A(n7276), .B(n7275), .ZN(n9335) );
  MUX2_X1 U8487 ( .A(P2_REG2_REG_14__SCAN_IN), .B(P2_REG1_REG_14__SCAN_IN), 
        .S(n9074), .Z(n7278) );
  OR2_X1 U8488 ( .A1(n7278), .A2(n9322), .ZN(n7307) );
  XNOR2_X1 U8489 ( .A(n7278), .B(n7277), .ZN(n9318) );
  MUX2_X1 U8490 ( .A(P2_REG2_REG_13__SCAN_IN), .B(P2_REG1_REG_13__SCAN_IN), 
        .S(n9074), .Z(n7280) );
  OR2_X1 U8491 ( .A1(n7280), .A2(n9305), .ZN(n7306) );
  XNOR2_X1 U8492 ( .A(n7280), .B(n7279), .ZN(n9301) );
  MUX2_X1 U8493 ( .A(P2_REG2_REG_12__SCAN_IN), .B(P2_REG1_REG_12__SCAN_IN), 
        .S(n9074), .Z(n7282) );
  OR2_X1 U8494 ( .A1(n7282), .A2(n8638), .ZN(n7305) );
  XNOR2_X1 U8495 ( .A(n7282), .B(n7281), .ZN(n8634) );
  MUX2_X1 U8496 ( .A(P2_REG2_REG_11__SCAN_IN), .B(P2_REG1_REG_11__SCAN_IN), 
        .S(n9074), .Z(n7283) );
  OR2_X1 U8497 ( .A1(n7283), .A2(n7482), .ZN(n7304) );
  XNOR2_X1 U8498 ( .A(n7283), .B(n10496), .ZN(n10502) );
  MUX2_X1 U8499 ( .A(P2_REG2_REG_10__SCAN_IN), .B(P2_REG1_REG_10__SCAN_IN), 
        .S(n9074), .Z(n7284) );
  OR2_X1 U8500 ( .A1(n7284), .A2(n7463), .ZN(n7303) );
  XNOR2_X1 U8501 ( .A(n7284), .B(n10479), .ZN(n10485) );
  MUX2_X1 U8502 ( .A(P2_REG2_REG_9__SCAN_IN), .B(P2_REG1_REG_9__SCAN_IN), .S(
        n9074), .Z(n7285) );
  OR2_X1 U8503 ( .A1(n7285), .A2(n7460), .ZN(n7302) );
  XNOR2_X1 U8504 ( .A(n7285), .B(n10463), .ZN(n10468) );
  MUX2_X1 U8505 ( .A(P2_REG2_REG_8__SCAN_IN), .B(P2_REG1_REG_8__SCAN_IN), .S(
        n9074), .Z(n7286) );
  OR2_X1 U8506 ( .A1(n7286), .A2(n7457), .ZN(n7301) );
  XNOR2_X1 U8507 ( .A(n7286), .B(n10447), .ZN(n10453) );
  MUX2_X1 U8508 ( .A(P2_REG2_REG_7__SCAN_IN), .B(P2_REG1_REG_7__SCAN_IN), .S(
        n9074), .Z(n7287) );
  OR2_X1 U8509 ( .A1(n7287), .A2(n7452), .ZN(n7300) );
  XNOR2_X1 U8510 ( .A(n7287), .B(n10431), .ZN(n10436) );
  MUX2_X1 U8511 ( .A(P2_REG2_REG_6__SCAN_IN), .B(P2_REG1_REG_6__SCAN_IN), .S(
        n9074), .Z(n7288) );
  OR2_X1 U8512 ( .A1(n7288), .A2(n7441), .ZN(n7299) );
  XNOR2_X1 U8513 ( .A(n7288), .B(n10414), .ZN(n10417) );
  INV_X1 U8514 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n7938) );
  MUX2_X1 U8515 ( .A(n7938), .B(n10402), .S(n9074), .Z(n7289) );
  NOR2_X1 U8516 ( .A1(n7289), .A2(n7290), .ZN(n7298) );
  AOI21_X1 U8517 ( .B1(n7290), .B2(n7289), .A(n7298), .ZN(n10395) );
  MUX2_X1 U8518 ( .A(P2_REG2_REG_4__SCAN_IN), .B(P2_REG1_REG_4__SCAN_IN), .S(
        n9074), .Z(n7296) );
  INV_X1 U8519 ( .A(n7296), .ZN(n7297) );
  MUX2_X1 U8520 ( .A(P2_REG2_REG_3__SCAN_IN), .B(P2_REG1_REG_3__SCAN_IN), .S(
        n9074), .Z(n7291) );
  OR2_X1 U8521 ( .A1(n7291), .A2(n7434), .ZN(n7295) );
  XNOR2_X1 U8522 ( .A(n7291), .B(n10360), .ZN(n10362) );
  MUX2_X1 U8523 ( .A(P2_REG2_REG_2__SCAN_IN), .B(P2_REG1_REG_2__SCAN_IN), .S(
        n9074), .Z(n7294) );
  MUX2_X1 U8524 ( .A(P2_REG2_REG_1__SCAN_IN), .B(P2_REG1_REG_1__SCAN_IN), .S(
        n9074), .Z(n7293) );
  INV_X1 U8525 ( .A(n7203), .ZN(n7430) );
  XOR2_X1 U8526 ( .A(n7203), .B(n7293), .Z(n7588) );
  INV_X1 U8527 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n7292) );
  INV_X1 U8528 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n7547) );
  MUX2_X1 U8529 ( .A(n7292), .B(n7547), .S(n9074), .Z(n10353) );
  AND2_X1 U8530 ( .A1(n10353), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n7587) );
  NOR2_X1 U8531 ( .A1(n7588), .A2(n7587), .ZN(n7585) );
  AOI21_X1 U8532 ( .B1(n7293), .B2(n7430), .A(n7585), .ZN(n7578) );
  XOR2_X1 U8533 ( .A(n7582), .B(n7294), .Z(n7579) );
  NOR2_X1 U8534 ( .A1(n7578), .A2(n7579), .ZN(n7577) );
  NAND2_X1 U8535 ( .A1(n10362), .A2(n10363), .ZN(n10361) );
  XNOR2_X1 U8536 ( .A(n7296), .B(n10376), .ZN(n10385) );
  NAND2_X1 U8537 ( .A1(n10386), .A2(n10385), .ZN(n10384) );
  OAI21_X1 U8538 ( .B1(n10376), .B2(n7297), .A(n10384), .ZN(n10394) );
  AND2_X1 U8539 ( .A1(n10394), .A2(n10395), .ZN(n10396) );
  NOR2_X1 U8540 ( .A1(n7298), .A2(n10396), .ZN(n10416) );
  NAND2_X1 U8541 ( .A1(n10436), .A2(n10435), .ZN(n10434) );
  NAND2_X1 U8542 ( .A1(n7300), .A2(n10434), .ZN(n10452) );
  NAND2_X1 U8543 ( .A1(n10453), .A2(n10452), .ZN(n10451) );
  NAND2_X1 U8544 ( .A1(n7301), .A2(n10451), .ZN(n10467) );
  NAND2_X1 U8545 ( .A1(n10468), .A2(n10467), .ZN(n10466) );
  NAND2_X1 U8546 ( .A1(n7302), .A2(n10466), .ZN(n10484) );
  NAND2_X1 U8547 ( .A1(n10502), .A2(n10501), .ZN(n10500) );
  NAND2_X1 U8548 ( .A1(n7304), .A2(n10500), .ZN(n8633) );
  NAND2_X1 U8549 ( .A1(n9301), .A2(n9300), .ZN(n9299) );
  NAND2_X1 U8550 ( .A1(n7306), .A2(n9299), .ZN(n9317) );
  NAND2_X1 U8551 ( .A1(n9318), .A2(n9317), .ZN(n9316) );
  NAND2_X1 U8552 ( .A1(n7307), .A2(n9316), .ZN(n9334) );
  NAND2_X1 U8553 ( .A1(n9335), .A2(n9334), .ZN(n9333) );
  NAND2_X1 U8554 ( .A1(n7308), .A2(n9333), .ZN(n9351) );
  NAND2_X1 U8555 ( .A1(n9368), .A2(n9367), .ZN(n9366) );
  INV_X1 U8556 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n7311) );
  MUX2_X1 U8557 ( .A(n9380), .B(n7311), .S(n9074), .Z(n7312) );
  NAND2_X1 U8558 ( .A1(n7313), .A2(n7312), .ZN(n9383) );
  NOR2_X1 U8559 ( .A1(n7313), .A2(n7312), .ZN(n9385) );
  XOR2_X1 U8560 ( .A(n7315), .B(n7314), .Z(n7321) );
  NOR2_X1 U8561 ( .A1(n9074), .A2(P2_U3151), .ZN(n9673) );
  NAND2_X1 U8562 ( .A1(n7316), .A2(n9673), .ZN(n7317) );
  MUX2_X1 U8563 ( .A(n7317), .B(n9292), .S(n9075), .Z(n10403) );
  NOR2_X1 U8564 ( .A1(n10403), .A2(n8090), .ZN(n7320) );
  INV_X1 U8565 ( .A(n7490), .ZN(n8379) );
  NOR2_X1 U8566 ( .A1(n7491), .A2(n8379), .ZN(n7318) );
  NAND2_X1 U8567 ( .A1(P2_U3151), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n9173) );
  OAI21_X1 U8568 ( .B1(n10412), .B2(n5398), .A(n9173), .ZN(n7319) );
  AOI211_X1 U8569 ( .C1(n7321), .C2(n10504), .A(n7320), .B(n7319), .ZN(n7322)
         );
  OAI21_X1 U8570 ( .B1(n7328), .B2(n7327), .A(n9784), .ZN(n7334) );
  NAND2_X1 U8571 ( .A1(n7329), .A2(n9789), .ZN(n7333) );
  AOI22_X1 U8572 ( .A1(n9788), .A2(n9966), .B1(n9787), .B2(n9795), .ZN(n7331)
         );
  AOI22_X1 U8573 ( .A1(n9786), .A2(n9797), .B1(P1_REG3_REG_27__SCAN_IN), .B2(
        P1_U3086), .ZN(n7330) );
  AND2_X1 U8574 ( .A1(n7331), .A2(n7330), .ZN(n7332) );
  NAND3_X1 U8575 ( .A1(n7334), .A2(n7333), .A3(n7332), .ZN(P1_U3214) );
  NAND2_X1 U8576 ( .A1(n7335), .A2(n7338), .ZN(n7513) );
  OR2_X1 U8577 ( .A1(n7336), .A2(n9070), .ZN(n7340) );
  NOR2_X1 U8578 ( .A1(n7340), .A2(n8866), .ZN(n7508) );
  NOR2_X1 U8579 ( .A1(n9150), .A2(n7508), .ZN(n7337) );
  OR2_X1 U8580 ( .A1(n7513), .A2(n7337), .ZN(n7343) );
  NAND3_X1 U8581 ( .A1(n6883), .A2(n7339), .A3(n7338), .ZN(n7518) );
  NAND3_X1 U8582 ( .A1(n9053), .A2(n9618), .A3(n7340), .ZN(n7510) );
  NAND2_X1 U8583 ( .A1(n7510), .A2(n10585), .ZN(n7488) );
  INV_X1 U8584 ( .A(n7488), .ZN(n7341) );
  OR2_X1 U8585 ( .A1(n7518), .A2(n7341), .ZN(n7342) );
  NAND2_X1 U8586 ( .A1(n7343), .A2(n7342), .ZN(n7348) );
  NAND2_X1 U8587 ( .A1(n7344), .A2(n10695), .ZN(n7347) );
  INV_X1 U8588 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n7345) );
  OR2_X1 U8589 ( .A1(n10695), .A2(n7345), .ZN(n7346) );
  NAND2_X1 U8590 ( .A1(n7348), .A2(n7514), .ZN(n9654) );
  NAND2_X1 U8591 ( .A1(n5503), .A2(n5509), .ZN(P2_U3455) );
  NAND2_X1 U8592 ( .A1(n9969), .A2(n9984), .ZN(n7349) );
  AND2_X1 U8593 ( .A1(n9980), .A2(n7349), .ZN(n7353) );
  INV_X1 U8594 ( .A(n7349), .ZN(n7352) );
  AND2_X1 U8595 ( .A1(n5370), .A2(n7350), .ZN(n7351) );
  NAND2_X1 U8596 ( .A1(n7354), .A2(n7356), .ZN(n7355) );
  NAND2_X1 U8597 ( .A1(n7362), .A2(n7358), .ZN(n7357) );
  INV_X1 U8598 ( .A(n7356), .ZN(n7360) );
  NAND2_X1 U8599 ( .A1(n7357), .A2(n7360), .ZN(n7363) );
  INV_X1 U8600 ( .A(n7358), .ZN(n7359) );
  NOR2_X1 U8601 ( .A1(n7360), .A2(n7359), .ZN(n7361) );
  NAND2_X1 U8602 ( .A1(n7363), .A2(n9936), .ZN(n7365) );
  OAI22_X1 U8603 ( .A1(n8281), .A2(n10145), .B1(n9984), .B2(n10143), .ZN(n7364) );
  AOI21_X1 U8604 ( .B1(n7365), .B2(n10127), .A(n7364), .ZN(n9964) );
  OAI211_X1 U8605 ( .C1(n9959), .C2(n7367), .A(n10552), .B(n9948), .ZN(n9956)
         );
  INV_X1 U8606 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n7370) );
  INV_X1 U8607 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n7374) );
  OR2_X1 U8608 ( .A1(n10646), .A2(n7374), .ZN(n7375) );
  NAND2_X1 U8609 ( .A1(n5504), .A2(n5510), .ZN(P1_U3550) );
  NOR2_X4 U8610 ( .A1(n6951), .A2(n7378), .ZN(P1_U3973) );
  NAND2_X1 U8611 ( .A1(n8108), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n7379) );
  OAI21_X1 U8612 ( .B1(n8108), .B2(P1_REG2_REG_13__SCAN_IN), .A(n7379), .ZN(
        n8103) );
  NOR2_X1 U8613 ( .A1(P1_REG2_REG_12__SCAN_IN), .A2(n7414), .ZN(n7380) );
  AOI21_X1 U8614 ( .B1(n7414), .B2(P1_REG2_REG_12__SCAN_IN), .A(n7380), .ZN(
        n7798) );
  NOR2_X1 U8615 ( .A1(P1_REG2_REG_9__SCAN_IN), .A2(n8621), .ZN(n7381) );
  AOI21_X1 U8616 ( .B1(n8621), .B2(P1_REG2_REG_9__SCAN_IN), .A(n7381), .ZN(
        n7536) );
  INV_X1 U8617 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n7382) );
  MUX2_X1 U8618 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n7382), .S(n9831), .Z(n9834)
         );
  INV_X1 U8619 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n7856) );
  MUX2_X1 U8620 ( .A(P1_REG2_REG_1__SCAN_IN), .B(n7856), .S(n9812), .Z(n9815)
         );
  AND2_X1 U8621 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n9814) );
  NAND2_X1 U8622 ( .A1(n9815), .A2(n9814), .ZN(n9813) );
  NAND2_X1 U8623 ( .A1(n9812), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n7383) );
  NAND2_X1 U8624 ( .A1(n9813), .A2(n7383), .ZN(n9833) );
  NAND2_X1 U8625 ( .A1(n9834), .A2(n9833), .ZN(n9832) );
  NAND2_X1 U8626 ( .A1(n9831), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n7384) );
  NAND2_X1 U8627 ( .A1(n9832), .A2(n7384), .ZN(n9850) );
  INV_X1 U8628 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n7385) );
  XNOR2_X1 U8629 ( .A(n9848), .B(n7385), .ZN(n9851) );
  NAND2_X1 U8630 ( .A1(n9850), .A2(n9851), .ZN(n9849) );
  NAND2_X1 U8631 ( .A1(n9848), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n7386) );
  NAND2_X1 U8632 ( .A1(n9849), .A2(n7386), .ZN(n10525) );
  OR2_X1 U8633 ( .A1(n10527), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n7388) );
  NAND2_X1 U8634 ( .A1(P1_REG2_REG_4__SCAN_IN), .A2(n10527), .ZN(n7387) );
  AND2_X1 U8635 ( .A1(n7388), .A2(n7387), .ZN(n10526) );
  AND2_X1 U8636 ( .A1(n10525), .A2(n10526), .ZN(n10522) );
  NAND2_X1 U8637 ( .A1(P1_REG2_REG_5__SCAN_IN), .A2(n7643), .ZN(n7389) );
  OAI21_X1 U8638 ( .B1(P1_REG2_REG_5__SCAN_IN), .B2(n7643), .A(n7389), .ZN(
        n7639) );
  NOR2_X1 U8639 ( .A1(n7638), .A2(n7639), .ZN(n7637) );
  AOI21_X1 U8640 ( .B1(n7643), .B2(P1_REG2_REG_5__SCAN_IN), .A(n7637), .ZN(
        n7614) );
  NAND2_X1 U8641 ( .A1(n7619), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n7390) );
  OAI21_X1 U8642 ( .B1(n7619), .B2(P1_REG2_REG_6__SCAN_IN), .A(n7390), .ZN(
        n7615) );
  NOR2_X1 U8643 ( .A1(n7614), .A2(n7615), .ZN(n7613) );
  NAND2_X1 U8644 ( .A1(n7607), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n7391) );
  OAI21_X1 U8645 ( .B1(n7607), .B2(P1_REG2_REG_7__SCAN_IN), .A(n7391), .ZN(
        n7603) );
  NOR2_X1 U8646 ( .A1(n7602), .A2(n7603), .ZN(n7601) );
  AOI21_X1 U8647 ( .B1(P1_REG2_REG_7__SCAN_IN), .B2(n7607), .A(n7601), .ZN(
        n7626) );
  NAND2_X1 U8648 ( .A1(P1_REG2_REG_8__SCAN_IN), .A2(n7631), .ZN(n7392) );
  OAI21_X1 U8649 ( .B1(P1_REG2_REG_8__SCAN_IN), .B2(n7631), .A(n7392), .ZN(
        n7627) );
  NOR2_X1 U8650 ( .A1(n7626), .A2(n7627), .ZN(n7625) );
  NAND2_X1 U8651 ( .A1(n7536), .A2(n7535), .ZN(n7534) );
  OAI21_X1 U8652 ( .B1(P1_REG2_REG_9__SCAN_IN), .B2(n8621), .A(n7534), .ZN(
        n7657) );
  INV_X1 U8653 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n7393) );
  AOI22_X1 U8654 ( .A1(P1_REG2_REG_10__SCAN_IN), .A2(n7466), .B1(n7662), .B2(
        n7393), .ZN(n7658) );
  NOR2_X1 U8655 ( .A1(n7657), .A2(n7658), .ZN(n7656) );
  NAND2_X1 U8656 ( .A1(P1_REG2_REG_11__SCAN_IN), .A2(n7752), .ZN(n7394) );
  OAI21_X1 U8657 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n7752), .A(n7394), .ZN(
        n7747) );
  NOR2_X1 U8658 ( .A1(n7748), .A2(n7747), .ZN(n7746) );
  AOI21_X1 U8659 ( .B1(n7752), .B2(P1_REG2_REG_11__SCAN_IN), .A(n7746), .ZN(
        n7797) );
  NAND2_X1 U8660 ( .A1(n7798), .A2(n7797), .ZN(n7796) );
  OAI21_X1 U8661 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(n7414), .A(n7796), .ZN(
        n8104) );
  NOR2_X1 U8662 ( .A1(n8103), .A2(n8104), .ZN(n8102) );
  INV_X1 U8663 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n7395) );
  AOI22_X1 U8664 ( .A1(P1_REG2_REG_14__SCAN_IN), .A2(n7670), .B1(n8229), .B2(
        n7395), .ZN(n8225) );
  NOR2_X1 U8665 ( .A1(n8224), .A2(n8225), .ZN(n8223) );
  XNOR2_X1 U8666 ( .A(n9864), .B(n9865), .ZN(n7401) );
  INV_X1 U8667 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n7400) );
  NOR2_X1 U8668 ( .A1(n7400), .A2(n7401), .ZN(n9866) );
  INV_X1 U8669 ( .A(n7397), .ZN(n7396) );
  OAI21_X1 U8670 ( .B1(n6951), .B2(n7396), .A(P1_STATE_REG_SCAN_IN), .ZN(n7421) );
  NAND2_X1 U8671 ( .A1(n7398), .A2(n7397), .ZN(n7399) );
  NAND2_X1 U8672 ( .A1(n5618), .A2(n7399), .ZN(n7419) );
  AOI211_X1 U8673 ( .C1(n7401), .C2(n7400), .A(n9866), .B(n9894), .ZN(n7426)
         );
  INV_X1 U8674 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n10670) );
  AOI22_X1 U8675 ( .A1(P1_REG1_REG_12__SCAN_IN), .A2(n7414), .B1(n7806), .B2(
        n10670), .ZN(n7801) );
  INV_X1 U8676 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n7402) );
  MUX2_X1 U8677 ( .A(n7402), .B(P1_REG1_REG_10__SCAN_IN), .S(n7662), .Z(n7660)
         );
  INV_X1 U8678 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n7403) );
  MUX2_X1 U8679 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n7403), .S(n8621), .Z(n7533)
         );
  INV_X1 U8680 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n10567) );
  MUX2_X1 U8681 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n10567), .S(n9831), .Z(n9837)
         );
  INV_X1 U8682 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n10545) );
  MUX2_X1 U8683 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n10545), .S(n9812), .Z(n9811)
         );
  AND2_X1 U8684 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n9810) );
  NAND2_X1 U8685 ( .A1(n9811), .A2(n9810), .ZN(n9809) );
  NAND2_X1 U8686 ( .A1(n9812), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n7404) );
  NAND2_X1 U8687 ( .A1(n9809), .A2(n7404), .ZN(n9836) );
  NAND2_X1 U8688 ( .A1(n9837), .A2(n9836), .ZN(n9835) );
  NAND2_X1 U8689 ( .A1(n9831), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n7405) );
  NAND2_X1 U8690 ( .A1(n9835), .A2(n7405), .ZN(n9843) );
  INV_X1 U8691 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n7406) );
  XNOR2_X1 U8692 ( .A(n9848), .B(n7406), .ZN(n9844) );
  NAND2_X1 U8693 ( .A1(n9843), .A2(n9844), .ZN(n9842) );
  NAND2_X1 U8694 ( .A1(n9848), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n7407) );
  NAND2_X1 U8695 ( .A1(n9842), .A2(n7407), .ZN(n10520) );
  OR2_X1 U8696 ( .A1(n10527), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n7409) );
  NAND2_X1 U8697 ( .A1(P1_REG1_REG_4__SCAN_IN), .A2(n10527), .ZN(n7408) );
  AND2_X1 U8698 ( .A1(n7409), .A2(n7408), .ZN(n10521) );
  AND2_X1 U8699 ( .A1(n10520), .A2(n10521), .ZN(n10517) );
  AOI21_X1 U8700 ( .B1(P1_REG1_REG_4__SCAN_IN), .B2(n10527), .A(n10517), .ZN(
        n7642) );
  NAND2_X1 U8701 ( .A1(P1_REG1_REG_5__SCAN_IN), .A2(n7643), .ZN(n7410) );
  OAI21_X1 U8702 ( .B1(n7643), .B2(P1_REG1_REG_5__SCAN_IN), .A(n7410), .ZN(
        n7641) );
  NOR2_X1 U8703 ( .A1(n7642), .A2(n7641), .ZN(n7640) );
  AOI21_X1 U8704 ( .B1(n7643), .B2(P1_REG1_REG_5__SCAN_IN), .A(n7640), .ZN(
        n7618) );
  NAND2_X1 U8705 ( .A1(n7619), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n7411) );
  OAI21_X1 U8706 ( .B1(n7619), .B2(P1_REG1_REG_6__SCAN_IN), .A(n7411), .ZN(
        n7617) );
  NOR2_X1 U8707 ( .A1(n7618), .A2(n7617), .ZN(n7616) );
  AOI21_X1 U8708 ( .B1(n7619), .B2(P1_REG1_REG_6__SCAN_IN), .A(n7616), .ZN(
        n7606) );
  INV_X1 U8709 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n7412) );
  MUX2_X1 U8710 ( .A(n7412), .B(P1_REG1_REG_7__SCAN_IN), .S(n7607), .Z(n7605)
         );
  NOR2_X1 U8711 ( .A1(n7606), .A2(n7605), .ZN(n7604) );
  AOI21_X1 U8712 ( .B1(n7607), .B2(P1_REG1_REG_7__SCAN_IN), .A(n7604), .ZN(
        n7630) );
  INV_X1 U8713 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n7413) );
  MUX2_X1 U8714 ( .A(n7413), .B(P1_REG1_REG_8__SCAN_IN), .S(n7631), .Z(n7629)
         );
  NOR2_X1 U8715 ( .A1(n7630), .A2(n7629), .ZN(n7628) );
  AOI21_X1 U8716 ( .B1(n7631), .B2(P1_REG1_REG_8__SCAN_IN), .A(n7628), .ZN(
        n7532) );
  NAND2_X1 U8717 ( .A1(n7533), .A2(n7532), .ZN(n7531) );
  OAI21_X1 U8718 ( .B1(n8621), .B2(P1_REG1_REG_9__SCAN_IN), .A(n7531), .ZN(
        n7661) );
  NOR2_X1 U8719 ( .A1(n7660), .A2(n7661), .ZN(n7659) );
  AOI21_X1 U8720 ( .B1(n7662), .B2(P1_REG1_REG_10__SCAN_IN), .A(n7659), .ZN(
        n7751) );
  MUX2_X1 U8721 ( .A(n8654), .B(P1_REG1_REG_11__SCAN_IN), .S(n7752), .Z(n7750)
         );
  NOR2_X1 U8722 ( .A1(n7751), .A2(n7750), .ZN(n7749) );
  AOI21_X1 U8723 ( .B1(n7752), .B2(P1_REG1_REG_11__SCAN_IN), .A(n7749), .ZN(
        n7800) );
  NAND2_X1 U8724 ( .A1(n7801), .A2(n7800), .ZN(n7799) );
  OAI21_X1 U8725 ( .B1(P1_REG1_REG_12__SCAN_IN), .B2(n7414), .A(n7799), .ZN(
        n8107) );
  INV_X1 U8726 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n7415) );
  MUX2_X1 U8727 ( .A(n7415), .B(P1_REG1_REG_13__SCAN_IN), .S(n8108), .Z(n8106)
         );
  NOR2_X1 U8728 ( .A1(n8107), .A2(n8106), .ZN(n8105) );
  AOI21_X1 U8729 ( .B1(n8108), .B2(P1_REG1_REG_13__SCAN_IN), .A(n8105), .ZN(
        n8228) );
  XNOR2_X1 U8730 ( .A(n8229), .B(P1_REG1_REG_14__SCAN_IN), .ZN(n8227) );
  NOR2_X1 U8731 ( .A1(n8228), .A2(n8227), .ZN(n8226) );
  AOI21_X1 U8732 ( .B1(n8229), .B2(P1_REG1_REG_14__SCAN_IN), .A(n8226), .ZN(
        n9855) );
  XNOR2_X1 U8733 ( .A(n9864), .B(n9855), .ZN(n7418) );
  INV_X1 U8734 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n7417) );
  NOR2_X1 U8735 ( .A1(n7417), .A2(n7418), .ZN(n9856) );
  INV_X1 U8736 ( .A(n7478), .ZN(n7416) );
  AOI211_X1 U8737 ( .C1(n7418), .C2(n7417), .A(n9856), .B(n9926), .ZN(n7425)
         );
  NOR2_X2 U8738 ( .A1(n7478), .A2(n10287), .ZN(n10528) );
  INV_X1 U8739 ( .A(n10528), .ZN(n9887) );
  NOR2_X1 U8740 ( .A1(n9887), .A2(n9864), .ZN(n7424) );
  INV_X1 U8741 ( .A(n7419), .ZN(n7420) );
  OR2_X1 U8742 ( .A1(n7421), .A2(n7420), .ZN(n9921) );
  INV_X1 U8743 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n7422) );
  NAND2_X1 U8744 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n8830) );
  OAI21_X1 U8745 ( .B1(n9921), .B2(n7422), .A(n8830), .ZN(n7423) );
  OR4_X1 U8746 ( .A1(n7426), .A2(n7425), .A3(n7424), .A4(n7423), .ZN(P1_U3258)
         );
  INV_X1 U8747 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n7428) );
  INV_X1 U8748 ( .A(n9674), .ZN(n9137) );
  OAI222_X1 U8749 ( .A1(n9676), .A2(n7443), .B1(n7429), .B2(P2_U3151), .C1(
        n7428), .C2(n9137), .ZN(P2_U3291) );
  OAI222_X1 U8750 ( .A1(n9676), .A2(n7437), .B1(n7430), .B2(P2_U3151), .C1(
        n5520), .C2(n9137), .ZN(P2_U3294) );
  INV_X1 U8751 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n7431) );
  OAI222_X1 U8752 ( .A1(n9676), .A2(n7447), .B1(n10404), .B2(P2_U3151), .C1(
        n7431), .C2(n9137), .ZN(P2_U3290) );
  INV_X1 U8753 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n7433) );
  OAI222_X1 U8754 ( .A1(n9137), .A2(n7433), .B1(n7432), .B2(P2_U3151), .C1(
        n9676), .C2(n7439), .ZN(P2_U3293) );
  OAI222_X1 U8755 ( .A1(n9137), .A2(n5071), .B1(n7434), .B2(P2_U3151), .C1(
        n9676), .C2(n7445), .ZN(P2_U3292) );
  AND2_X1 U8756 ( .A1(n7435), .A2(P1_U3086), .ZN(n8622) );
  INV_X2 U8757 ( .A(n8622), .ZN(n10293) );
  NOR2_X2 U8758 ( .A1(n7435), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10286) );
  AOI22_X1 U8759 ( .A1(n10286), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(
        P1_STATE_REG_SCAN_IN), .B2(n9812), .ZN(n7436) );
  OAI21_X1 U8760 ( .B1(n7437), .B2(n10293), .A(n7436), .ZN(P1_U3354) );
  AOI22_X1 U8761 ( .A1(n10286), .A2(P2_DATAO_REG_2__SCAN_IN), .B1(n9831), .B2(
        P1_STATE_REG_SCAN_IN), .ZN(n7438) );
  OAI21_X1 U8762 ( .B1(n7439), .B2(n10293), .A(n7438), .ZN(P1_U3353) );
  INV_X1 U8763 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n7440) );
  OAI222_X1 U8764 ( .A1(n9676), .A2(n7449), .B1(n7441), .B2(P2_U3151), .C1(
        n7440), .C2(n9137), .ZN(P2_U3289) );
  AOI22_X1 U8765 ( .A1(P2_DATAO_REG_4__SCAN_IN), .A2(n10286), .B1(n10527), 
        .B2(P1_STATE_REG_SCAN_IN), .ZN(n7442) );
  OAI21_X1 U8766 ( .B1(n7443), .B2(n10293), .A(n7442), .ZN(P1_U3351) );
  AOI22_X1 U8767 ( .A1(n9848), .A2(P1_STATE_REG_SCAN_IN), .B1(n10286), .B2(
        P2_DATAO_REG_3__SCAN_IN), .ZN(n7444) );
  OAI21_X1 U8768 ( .B1(n7445), .B2(n10293), .A(n7444), .ZN(P1_U3352) );
  AOI22_X1 U8769 ( .A1(n7643), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n10286), .ZN(n7446) );
  OAI21_X1 U8770 ( .B1(n7447), .B2(n10293), .A(n7446), .ZN(P1_U3350) );
  AOI22_X1 U8771 ( .A1(n7619), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n10286), .ZN(n7448) );
  OAI21_X1 U8772 ( .B1(n7449), .B2(n10293), .A(n7448), .ZN(P1_U3349) );
  AOI22_X1 U8773 ( .A1(n7607), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n10286), .ZN(n7450) );
  OAI21_X1 U8774 ( .B1(n7453), .B2(n10293), .A(n7450), .ZN(P1_U3348) );
  INV_X1 U8775 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n7451) );
  OAI222_X1 U8776 ( .A1(n9676), .A2(n7453), .B1(n7452), .B2(P2_U3151), .C1(
        n7451), .C2(n9137), .ZN(P2_U3288) );
  INV_X1 U8777 ( .A(n7454), .ZN(n7456) );
  AOI22_X1 U8778 ( .A1(n7631), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n10286), .ZN(n7455) );
  OAI21_X1 U8779 ( .B1(n7456), .B2(n10293), .A(n7455), .ZN(P1_U3347) );
  AND2_X1 U8780 ( .A1(n7467), .A2(P2_D_REG_8__SCAN_IN), .ZN(P2_U3257) );
  AND2_X1 U8781 ( .A1(n7467), .A2(P2_D_REG_20__SCAN_IN), .ZN(P2_U3245) );
  AND2_X1 U8782 ( .A1(n7467), .A2(P2_D_REG_23__SCAN_IN), .ZN(P2_U3242) );
  AND2_X1 U8783 ( .A1(n7467), .A2(P2_D_REG_9__SCAN_IN), .ZN(P2_U3256) );
  AND2_X1 U8784 ( .A1(n7467), .A2(P2_D_REG_29__SCAN_IN), .ZN(P2_U3236) );
  AND2_X1 U8785 ( .A1(n7467), .A2(P2_D_REG_17__SCAN_IN), .ZN(P2_U3248) );
  AND2_X1 U8786 ( .A1(n7467), .A2(P2_D_REG_14__SCAN_IN), .ZN(P2_U3251) );
  AND2_X1 U8787 ( .A1(n7467), .A2(P2_D_REG_11__SCAN_IN), .ZN(P2_U3254) );
  AND2_X1 U8788 ( .A1(n7467), .A2(P2_D_REG_6__SCAN_IN), .ZN(P2_U3259) );
  AND2_X1 U8789 ( .A1(n7467), .A2(P2_D_REG_3__SCAN_IN), .ZN(P2_U3262) );
  AND2_X1 U8790 ( .A1(n7467), .A2(P2_D_REG_26__SCAN_IN), .ZN(P2_U3239) );
  INV_X1 U8791 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n7887) );
  OAI222_X1 U8792 ( .A1(n7457), .A2(P2_U3151), .B1(n9676), .B2(n7456), .C1(
        n9137), .C2(n7887), .ZN(P2_U3287) );
  NAND2_X1 U8793 ( .A1(n9292), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n7458) );
  OAI21_X1 U8794 ( .B1(n5513), .B2(n9292), .A(n7458), .ZN(P2_U3491) );
  INV_X1 U8795 ( .A(n8623), .ZN(n7461) );
  INV_X1 U8796 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n7459) );
  OAI222_X1 U8797 ( .A1(n9676), .A2(n7461), .B1(n7460), .B2(P2_U3151), .C1(
        n7459), .C2(n9137), .ZN(P2_U3286) );
  INV_X1 U8798 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n7462) );
  OAI222_X1 U8799 ( .A1(n9676), .A2(n7465), .B1(n7463), .B2(P2_U3151), .C1(
        n7462), .C2(n9137), .ZN(P2_U3285) );
  OAI222_X1 U8800 ( .A1(P1_U3086), .A2(n7466), .B1(n10293), .B2(n7465), .C1(
        n7464), .C2(n10290), .ZN(P1_U3345) );
  INV_X1 U8801 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n7471) );
  AND2_X1 U8802 ( .A1(n7468), .A2(n6881), .ZN(n7469) );
  AOI22_X1 U8803 ( .A1(n7467), .A2(n7471), .B1(n7470), .B2(n7469), .ZN(
        P2_U3376) );
  INV_X1 U8804 ( .A(n10294), .ZN(n7472) );
  OR2_X1 U8805 ( .A1(n9821), .A2(n7472), .ZN(n9827) );
  INV_X1 U8806 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n7473) );
  OAI22_X1 U8807 ( .A1(n7474), .A2(n9820), .B1(n9827), .B2(n7473), .ZN(n7475)
         );
  XNOR2_X1 U8808 ( .A(n7475), .B(P1_IR_REG_0__SCAN_IN), .ZN(n7479) );
  NAND2_X1 U8809 ( .A1(P1_U3086), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n7477) );
  INV_X1 U8810 ( .A(n9921), .ZN(n10534) );
  NAND2_X1 U8811 ( .A1(n10534), .A2(P1_ADDR_REG_0__SCAN_IN), .ZN(n7476) );
  OAI211_X1 U8812 ( .C1(n7479), .C2(n7478), .A(n7477), .B(n7476), .ZN(P1_U3243) );
  AND2_X1 U8813 ( .A1(n7467), .A2(P2_D_REG_5__SCAN_IN), .ZN(P2_U3260) );
  AND2_X1 U8814 ( .A1(n7467), .A2(P2_D_REG_25__SCAN_IN), .ZN(P2_U3240) );
  AND2_X1 U8815 ( .A1(n7467), .A2(P2_D_REG_10__SCAN_IN), .ZN(P2_U3255) );
  AND2_X1 U8816 ( .A1(n7467), .A2(P2_D_REG_19__SCAN_IN), .ZN(P2_U3246) );
  AND2_X1 U8817 ( .A1(n7467), .A2(P2_D_REG_2__SCAN_IN), .ZN(P2_U3263) );
  AND2_X1 U8818 ( .A1(n7467), .A2(P2_D_REG_16__SCAN_IN), .ZN(P2_U3249) );
  AND2_X1 U8819 ( .A1(n7467), .A2(P2_D_REG_4__SCAN_IN), .ZN(P2_U3261) );
  AND2_X1 U8820 ( .A1(n7467), .A2(P2_D_REG_7__SCAN_IN), .ZN(P2_U3258) );
  AND2_X1 U8821 ( .A1(n7467), .A2(P2_D_REG_24__SCAN_IN), .ZN(P2_U3241) );
  AND2_X1 U8822 ( .A1(n7467), .A2(P2_D_REG_31__SCAN_IN), .ZN(P2_U3234) );
  AND2_X1 U8823 ( .A1(n7467), .A2(P2_D_REG_21__SCAN_IN), .ZN(P2_U3244) );
  AND2_X1 U8824 ( .A1(n7467), .A2(P2_D_REG_28__SCAN_IN), .ZN(P2_U3237) );
  AND2_X1 U8825 ( .A1(n7467), .A2(P2_D_REG_12__SCAN_IN), .ZN(P2_U3253) );
  AND2_X1 U8826 ( .A1(n7467), .A2(P2_D_REG_13__SCAN_IN), .ZN(P2_U3252) );
  AND2_X1 U8827 ( .A1(n7467), .A2(P2_D_REG_30__SCAN_IN), .ZN(P2_U3235) );
  AND2_X1 U8828 ( .A1(n7467), .A2(P2_D_REG_15__SCAN_IN), .ZN(P2_U3250) );
  AND2_X1 U8829 ( .A1(n7467), .A2(P2_D_REG_27__SCAN_IN), .ZN(P2_U3238) );
  AND2_X1 U8830 ( .A1(n7467), .A2(P2_D_REG_22__SCAN_IN), .ZN(P2_U3243) );
  AND2_X1 U8831 ( .A1(n7467), .A2(P2_D_REG_18__SCAN_IN), .ZN(P2_U3247) );
  INV_X1 U8832 ( .A(n7480), .ZN(n7483) );
  AOI22_X1 U8833 ( .A1(n7752), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n10286), .ZN(n7481) );
  OAI21_X1 U8834 ( .B1(n7483), .B2(n10293), .A(n7481), .ZN(P1_U3344) );
  INV_X1 U8835 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n7484) );
  OAI222_X1 U8836 ( .A1(n9137), .A2(n7484), .B1(n9676), .B2(n7483), .C1(
        P2_U3151), .C2(n7482), .ZN(P2_U3284) );
  INV_X1 U8837 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n7485) );
  OAI222_X1 U8838 ( .A1(n9676), .A2(n7487), .B1(n8638), .B2(P2_U3151), .C1(
        n7485), .C2(n9137), .ZN(P2_U3283) );
  OAI222_X1 U8839 ( .A1(P1_U3086), .A2(n7806), .B1(n10293), .B2(n7487), .C1(
        n7486), .C2(n10290), .ZN(P1_U3343) );
  NAND2_X1 U8840 ( .A1(n7513), .A2(n7488), .ZN(n7494) );
  NAND3_X1 U8841 ( .A1(n7491), .A2(n7490), .A3(n7489), .ZN(n7492) );
  AOI21_X1 U8842 ( .B1(n7518), .B2(n7508), .A(n7492), .ZN(n7493) );
  NAND2_X1 U8843 ( .A1(n7494), .A2(n7493), .ZN(n7495) );
  NAND2_X1 U8844 ( .A1(n7495), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7497) );
  NAND2_X1 U8845 ( .A1(n9659), .A2(n9150), .ZN(n7517) );
  INV_X1 U8846 ( .A(n7517), .ZN(n9076) );
  NAND2_X1 U8847 ( .A1(n7518), .A2(n9076), .ZN(n7496) );
  NOR2_X1 U8848 ( .A1(n9266), .A2(P2_U3151), .ZN(n7561) );
  INV_X1 U8849 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n7776) );
  AND2_X1 U8850 ( .A1(n8927), .A2(n7498), .ZN(n7499) );
  NAND2_X1 U8851 ( .A1(n7500), .A2(n7499), .ZN(n7502) );
  NAND2_X1 U8852 ( .A1(n8866), .A2(n9070), .ZN(n7501) );
  NAND2_X1 U8853 ( .A1(n7503), .A2(n7504), .ZN(n7552) );
  NAND2_X1 U8854 ( .A1(n7507), .A2(n7506), .ZN(n7553) );
  OAI21_X1 U8855 ( .B1(n7507), .B2(n7506), .A(n7553), .ZN(n7512) );
  INV_X1 U8856 ( .A(n7508), .ZN(n7509) );
  OAI22_X1 U8857 ( .A1(n7513), .A2(n7510), .B1(n7509), .B2(n7518), .ZN(n7511)
         );
  NAND2_X1 U8858 ( .A1(n7512), .A2(n9256), .ZN(n7525) );
  INV_X1 U8859 ( .A(n7513), .ZN(n7515) );
  NAND2_X1 U8860 ( .A1(n7515), .A2(n7514), .ZN(n7516) );
  OR2_X1 U8861 ( .A1(n7518), .A2(n7517), .ZN(n7519) );
  NOR2_X2 U8862 ( .A1(n7519), .A2(n7520), .ZN(n9238) );
  INV_X1 U8863 ( .A(n7519), .ZN(n7521) );
  NAND2_X1 U8864 ( .A1(n7521), .A2(n7520), .ZN(n9240) );
  OAI22_X1 U8865 ( .A1(n9263), .A2(n7727), .B1(n5513), .B2(n9240), .ZN(n7522)
         );
  AOI21_X1 U8866 ( .B1(n7523), .B2(n9251), .A(n7522), .ZN(n7524) );
  OAI211_X1 U8867 ( .C1(n7561), .C2(n7776), .A(n7525), .B(n7524), .ZN(P2_U3162) );
  INV_X1 U8868 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n7529) );
  NOR2_X1 U8869 ( .A1(n5513), .A2(n7544), .ZN(n8925) );
  INV_X1 U8870 ( .A(n8925), .ZN(n7526) );
  NAND2_X1 U8871 ( .A1(n7526), .A2(n8926), .ZN(n8877) );
  NAND2_X1 U8872 ( .A1(n9615), .A2(n9498), .ZN(n7528) );
  AOI22_X1 U8873 ( .A1(n8877), .A2(n7528), .B1(n9609), .B2(n7527), .ZN(n7550)
         );
  MUX2_X1 U8874 ( .A(n7529), .B(n7550), .S(n10695), .Z(n7530) );
  OAI21_X1 U8875 ( .B1(n9148), .B2(n9654), .A(n7530), .ZN(P2_U3390) );
  OAI21_X1 U8876 ( .B1(n7533), .B2(n7532), .A(n7531), .ZN(n7538) );
  OAI21_X1 U8877 ( .B1(n7536), .B2(n7535), .A(n7534), .ZN(n7537) );
  AOI22_X1 U8878 ( .A1(n10519), .A2(n7538), .B1(n10524), .B2(n7537), .ZN(n7542) );
  INV_X1 U8879 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n7539) );
  NAND2_X1 U8880 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_U3086), .ZN(n8288) );
  OAI21_X1 U8881 ( .B1(n9921), .B2(n7539), .A(n8288), .ZN(n7540) );
  AOI21_X1 U8882 ( .B1(n10528), .B2(n8621), .A(n7540), .ZN(n7541) );
  NAND2_X1 U8883 ( .A1(n7542), .A2(n7541), .ZN(P1_U3252) );
  INV_X1 U8884 ( .A(n8877), .ZN(n9151) );
  INV_X1 U8885 ( .A(n7561), .ZN(n7543) );
  NAND2_X1 U8886 ( .A1(n7543), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n7546) );
  AOI22_X1 U8887 ( .A1(n7527), .A2(n9238), .B1(n9251), .B2(n7544), .ZN(n7545)
         );
  OAI211_X1 U8888 ( .C1(n9151), .C2(n9254), .A(n7546), .B(n7545), .ZN(P2_U3172) );
  OAI22_X1 U8889 ( .A1(n9148), .A2(n9594), .B1(n9627), .B2(n7547), .ZN(n7548)
         );
  INV_X1 U8890 ( .A(n7548), .ZN(n7549) );
  OAI21_X1 U8891 ( .B1(n7550), .B2(n9624), .A(n7549), .ZN(P2_U3459) );
  INV_X1 U8892 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n10584) );
  XNOR2_X1 U8893 ( .A(n7551), .B(n7558), .ZN(n7673) );
  XNOR2_X1 U8894 ( .A(n7673), .B(n9291), .ZN(n7555) );
  NAND2_X1 U8895 ( .A1(n7553), .A2(n7552), .ZN(n7554) );
  OAI21_X1 U8896 ( .B1(n7555), .B2(n7554), .A(n7675), .ZN(n7556) );
  NAND2_X1 U8897 ( .A1(n7556), .A2(n9256), .ZN(n7560) );
  OAI22_X1 U8898 ( .A1(n9263), .A2(n7792), .B1(n7503), .B2(n9240), .ZN(n7557)
         );
  AOI21_X1 U8899 ( .B1(n7558), .B2(n9251), .A(n7557), .ZN(n7559) );
  OAI211_X1 U8900 ( .C1(n7561), .C2(n10584), .A(n7560), .B(n7559), .ZN(
        P2_U3177) );
  INV_X1 U8901 ( .A(n10403), .ZN(n10497) );
  INV_X1 U8902 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n7576) );
  OAI21_X1 U8903 ( .B1(n7564), .B2(n7563), .A(n7562), .ZN(n7565) );
  AOI22_X1 U8904 ( .A1(n10370), .A2(n7565), .B1(P2_REG3_REG_2__SCAN_IN), .B2(
        P2_U3151), .ZN(n7575) );
  INV_X1 U8905 ( .A(n7567), .ZN(n7570) );
  INV_X1 U8906 ( .A(n7568), .ZN(n7569) );
  NAND2_X1 U8907 ( .A1(n7570), .A2(n7569), .ZN(n7571) );
  NAND2_X1 U8908 ( .A1(n7572), .A2(n7571), .ZN(n7573) );
  NAND2_X1 U8909 ( .A1(n10505), .A2(n7573), .ZN(n7574) );
  OAI211_X1 U8910 ( .C1(n7576), .C2(n10412), .A(n7575), .B(n7574), .ZN(n7581)
         );
  INV_X1 U8911 ( .A(n10504), .ZN(n7586) );
  AOI211_X1 U8912 ( .C1(n7579), .C2(n7578), .A(n7586), .B(n7577), .ZN(n7580)
         );
  AOI211_X1 U8913 ( .C1(n10497), .C2(n7582), .A(n7581), .B(n7580), .ZN(n7583)
         );
  INV_X1 U8914 ( .A(n7583), .ZN(P2_U3184) );
  AOI22_X1 U8915 ( .A1(n8108), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n10286), .ZN(n7584) );
  OAI21_X1 U8916 ( .B1(n7650), .B2(n10293), .A(n7584), .ZN(P1_U3342) );
  AOI211_X1 U8917 ( .C1(n7588), .C2(n7587), .A(n7586), .B(n7585), .ZN(n7599)
         );
  INV_X1 U8918 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n7597) );
  XNOR2_X1 U8919 ( .A(n7589), .B(P2_REG2_REG_1__SCAN_IN), .ZN(n7595) );
  NOR2_X1 U8920 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7776), .ZN(n7594) );
  NAND2_X1 U8921 ( .A1(n7590), .A2(n7723), .ZN(n7591) );
  AOI21_X1 U8922 ( .B1(n7592), .B2(n7591), .A(n10511), .ZN(n7593) );
  AOI211_X1 U8923 ( .C1(n10505), .C2(n7595), .A(n7594), .B(n7593), .ZN(n7596)
         );
  OAI21_X1 U8924 ( .B1(n10412), .B2(n7597), .A(n7596), .ZN(n7598) );
  AOI211_X1 U8925 ( .C1(n10497), .C2(n7203), .A(n7599), .B(n7598), .ZN(n7600)
         );
  INV_X1 U8926 ( .A(n7600), .ZN(P2_U3183) );
  AOI211_X1 U8927 ( .C1(n7603), .C2(n7602), .A(n7601), .B(n9894), .ZN(n7612)
         );
  AOI211_X1 U8928 ( .C1(n7606), .C2(n7605), .A(n7604), .B(n9926), .ZN(n7611)
         );
  INV_X1 U8929 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n7609) );
  NAND2_X1 U8930 ( .A1(n10528), .A2(n7607), .ZN(n7608) );
  NAND2_X1 U8931 ( .A1(P1_U3086), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n8152) );
  OAI211_X1 U8932 ( .C1(n7609), .C2(n9921), .A(n7608), .B(n8152), .ZN(n7610)
         );
  OR3_X1 U8933 ( .A1(n7612), .A2(n7611), .A3(n7610), .ZN(P1_U3250) );
  AOI211_X1 U8934 ( .C1(n7615), .C2(n7614), .A(n7613), .B(n9894), .ZN(n7624)
         );
  AOI211_X1 U8935 ( .C1(n7618), .C2(n7617), .A(n7616), .B(n9926), .ZN(n7623)
         );
  INV_X1 U8936 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n7621) );
  NAND2_X1 U8937 ( .A1(n10528), .A2(n7619), .ZN(n7620) );
  NAND2_X1 U8938 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n8054) );
  OAI211_X1 U8939 ( .C1(n7621), .C2(n9921), .A(n7620), .B(n8054), .ZN(n7622)
         );
  OR3_X1 U8940 ( .A1(n7624), .A2(n7623), .A3(n7622), .ZN(P1_U3249) );
  AOI211_X1 U8941 ( .C1(n7627), .C2(n7626), .A(n7625), .B(n9894), .ZN(n7636)
         );
  AOI211_X1 U8942 ( .C1(n7630), .C2(n7629), .A(n7628), .B(n9926), .ZN(n7635)
         );
  INV_X1 U8943 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n7633) );
  NAND2_X1 U8944 ( .A1(n10528), .A2(n7631), .ZN(n7632) );
  NAND2_X1 U8945 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_U3086), .ZN(n8164) );
  OAI211_X1 U8946 ( .C1(n7633), .C2(n9921), .A(n7632), .B(n8164), .ZN(n7634)
         );
  OR3_X1 U8947 ( .A1(n7636), .A2(n7635), .A3(n7634), .ZN(P1_U3251) );
  AOI211_X1 U8948 ( .C1(n7639), .C2(n7638), .A(n7637), .B(n9894), .ZN(n7648)
         );
  AOI211_X1 U8949 ( .C1(n7642), .C2(n7641), .A(n7640), .B(n9926), .ZN(n7647)
         );
  INV_X1 U8950 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n7645) );
  NAND2_X1 U8951 ( .A1(n10528), .A2(n7643), .ZN(n7644) );
  NAND2_X1 U8952 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n7926) );
  OAI211_X1 U8953 ( .C1(n7645), .C2(n9921), .A(n7644), .B(n7926), .ZN(n7646)
         );
  OR3_X1 U8954 ( .A1(n7648), .A2(n7647), .A3(n7646), .ZN(P1_U3248) );
  INV_X1 U8955 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n7649) );
  OAI222_X1 U8956 ( .A1(n9676), .A2(n7650), .B1(n9305), .B2(P2_U3151), .C1(
        n7649), .C2(n9137), .ZN(P2_U3282) );
  INV_X1 U8957 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n8319) );
  NAND2_X1 U8958 ( .A1(n9585), .A2(P2_U3893), .ZN(n7651) );
  OAI21_X1 U8959 ( .B1(P2_U3893), .B2(n8319), .A(n7651), .ZN(P2_U3512) );
  INV_X1 U8960 ( .A(n7824), .ZN(n7652) );
  OAI21_X1 U8961 ( .B1(n10667), .B2(n10127), .A(n7652), .ZN(n7653) );
  NAND2_X1 U8962 ( .A1(n6960), .A2(n10558), .ZN(n7825) );
  OAI211_X1 U8963 ( .C1(n7654), .C2(n7857), .A(n7653), .B(n7825), .ZN(n10241)
         );
  NAND2_X1 U8964 ( .A1(n10241), .A2(n10674), .ZN(n7655) );
  OAI21_X1 U8965 ( .B1(n10674), .B2(n5623), .A(n7655), .ZN(P1_U3453) );
  AOI211_X1 U8966 ( .C1(n7658), .C2(n7657), .A(n7656), .B(n9894), .ZN(n7667)
         );
  AOI211_X1 U8967 ( .C1(n7661), .C2(n7660), .A(n7659), .B(n9926), .ZN(n7666)
         );
  INV_X1 U8968 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n7664) );
  NAND2_X1 U8969 ( .A1(n10528), .A2(n7662), .ZN(n7663) );
  NAND2_X1 U8970 ( .A1(P1_REG3_REG_10__SCAN_IN), .A2(P1_U3086), .ZN(n8340) );
  OAI211_X1 U8971 ( .C1(n7664), .C2(n9921), .A(n7663), .B(n8340), .ZN(n7665)
         );
  OR3_X1 U8972 ( .A1(n7667), .A2(n7666), .A3(n7665), .ZN(P1_U3253) );
  INV_X1 U8973 ( .A(n7668), .ZN(n7671) );
  OAI222_X1 U8974 ( .A1(n7670), .A2(P1_U3086), .B1(n10293), .B2(n7671), .C1(
        n7669), .C2(n10290), .ZN(P1_U3341) );
  INV_X1 U8975 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n7672) );
  OAI222_X1 U8976 ( .A1(n9137), .A2(n7672), .B1(n9676), .B2(n7671), .C1(
        P2_U3151), .C2(n9322), .ZN(P2_U3281) );
  INV_X1 U8977 ( .A(n9266), .ZN(n7773) );
  NAND2_X1 U8978 ( .A1(n7727), .A2(n7673), .ZN(n7674) );
  XNOR2_X1 U8979 ( .A(n7725), .B(n7551), .ZN(n7705) );
  XNOR2_X1 U8980 ( .A(n7705), .B(n9290), .ZN(n7677) );
  AOI21_X1 U8981 ( .B1(n7676), .B2(n7677), .A(n9254), .ZN(n7679) );
  NAND2_X1 U8982 ( .A1(n7679), .A2(n7707), .ZN(n7682) );
  INV_X1 U8983 ( .A(n6853), .ZN(n9289) );
  NOR2_X1 U8984 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7782), .ZN(n10359) );
  OAI22_X1 U8985 ( .A1(n9270), .A2(n7725), .B1(n7727), .B2(n9240), .ZN(n7680)
         );
  AOI211_X1 U8986 ( .C1(n9238), .C2(n9289), .A(n10359), .B(n7680), .ZN(n7681)
         );
  OAI211_X1 U8987 ( .C1(P2_REG3_REG_3__SCAN_IN), .C2(n7773), .A(n7682), .B(
        n7681), .ZN(P2_U3158) );
  INV_X1 U8988 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n7683) );
  OAI222_X1 U8989 ( .A1(n9676), .A2(n7704), .B1(n5104), .B2(P2_U3151), .C1(
        n7683), .C2(n9137), .ZN(P2_U3280) );
  OAI21_X1 U8990 ( .B1(n7686), .B2(n7685), .A(n7684), .ZN(n7687) );
  INV_X1 U8991 ( .A(n7687), .ZN(n9823) );
  AOI22_X1 U8992 ( .A1(n9823), .A2(n9784), .B1(n9787), .B2(n6960), .ZN(n7690)
         );
  OR2_X1 U8993 ( .A1(n7688), .A2(P1_U3086), .ZN(n9765) );
  AOI22_X1 U8994 ( .A1(n9789), .A2(n7831), .B1(n9765), .B2(
        P1_REG3_REG_0__SCAN_IN), .ZN(n7689) );
  NAND2_X1 U8995 ( .A1(n7690), .A2(n7689), .ZN(P1_U3232) );
  XNOR2_X1 U8996 ( .A(n7692), .B(n7691), .ZN(n7694) );
  INV_X1 U8997 ( .A(n7696), .ZN(n7693) );
  NAND2_X1 U8998 ( .A1(n7694), .A2(n7693), .ZN(n7699) );
  INV_X1 U8999 ( .A(n7695), .ZN(n7697) );
  AOI22_X1 U9000 ( .A1(n7699), .A2(n7698), .B1(n7697), .B2(n7696), .ZN(n7702)
         );
  AOI22_X1 U9001 ( .A1(n9786), .A2(n7932), .B1(n9787), .B2(n6970), .ZN(n7701)
         );
  AOI22_X1 U9002 ( .A1(n7861), .A2(n9789), .B1(n9765), .B2(
        P1_REG3_REG_1__SCAN_IN), .ZN(n7700) );
  OAI211_X1 U9003 ( .C1(n7702), .C2(n9778), .A(n7701), .B(n7700), .ZN(P1_U3222) );
  OAI222_X1 U9004 ( .A1(P1_U3086), .A2(n9864), .B1(n10293), .B2(n7704), .C1(
        n7703), .C2(n10290), .ZN(P1_U3340) );
  NAND2_X1 U9005 ( .A1(n7705), .A2(n9290), .ZN(n7706) );
  NAND2_X1 U9006 ( .A1(n7707), .A2(n7706), .ZN(n7710) );
  AOI21_X1 U9007 ( .B1(n7710), .B2(n7709), .A(n5022), .ZN(n7715) );
  NOR2_X1 U9008 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7711), .ZN(n10375) );
  OAI22_X1 U9009 ( .A1(n9270), .A2(n5150), .B1(n7792), .B2(n9240), .ZN(n7712)
         );
  AOI211_X1 U9010 ( .C1(n9238), .C2(n9288), .A(n10375), .B(n7712), .ZN(n7714)
         );
  NAND2_X1 U9011 ( .A1(n9266), .A2(n7845), .ZN(n7713) );
  OAI211_X1 U9012 ( .C1(n7715), .C2(n9254), .A(n7714), .B(n7713), .ZN(P2_U3170) );
  OAI21_X1 U9013 ( .B1(n7719), .B2(n7717), .A(n7716), .ZN(n7780) );
  NOR2_X1 U9014 ( .A1(n6508), .A2(n9618), .ZN(n7721) );
  XNOR2_X1 U9015 ( .A(n7719), .B(n7718), .ZN(n7720) );
  OAI222_X1 U9016 ( .A1(n9616), .A2(n7727), .B1(n9515), .B2(n5513), .C1(n9498), 
        .C2(n7720), .ZN(n7777) );
  AOI211_X1 U9017 ( .C1(n9623), .C2(n7780), .A(n7721), .B(n7777), .ZN(n10538)
         );
  OR2_X1 U9018 ( .A1(n10538), .A2(n9624), .ZN(n7722) );
  OAI21_X1 U9019 ( .B1(n9627), .B2(n7723), .A(n7722), .ZN(P2_U3460) );
  XNOR2_X1 U9020 ( .A(n7724), .B(n8875), .ZN(n7788) );
  OAI22_X1 U9021 ( .A1(n6853), .A2(n9616), .B1(n7725), .B2(n9618), .ZN(n7729)
         );
  XNOR2_X1 U9022 ( .A(n7726), .B(n8875), .ZN(n7728) );
  OAI22_X1 U9023 ( .A1(n7728), .A2(n9498), .B1(n7727), .B2(n9515), .ZN(n7785)
         );
  AOI211_X1 U9024 ( .C1(n7788), .C2(n9623), .A(n7729), .B(n7785), .ZN(n10600)
         );
  NAND2_X1 U9025 ( .A1(n9624), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n7730) );
  OAI21_X1 U9026 ( .B1(n10600), .B2(n9624), .A(n7730), .ZN(P2_U3462) );
  INV_X1 U9027 ( .A(n7939), .ZN(n7738) );
  XNOR2_X1 U9028 ( .A(n7940), .B(n9115), .ZN(n7762) );
  XNOR2_X1 U9029 ( .A(n7762), .B(n9288), .ZN(n7732) );
  NOR3_X1 U9030 ( .A1(n5022), .A2(n5472), .A3(n7732), .ZN(n7734) );
  INV_X1 U9031 ( .A(n7765), .ZN(n7733) );
  OAI21_X1 U9032 ( .B1(n7734), .B2(n7733), .A(n9256), .ZN(n7737) );
  NOR2_X1 U9033 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6450), .ZN(n10409) );
  OAI22_X1 U9034 ( .A1(n9270), .A2(n8043), .B1(n6853), .B2(n9240), .ZN(n7735)
         );
  AOI211_X1 U9035 ( .C1(n9238), .C2(n9287), .A(n10409), .B(n7735), .ZN(n7736)
         );
  OAI211_X1 U9036 ( .C1(n7738), .C2(n7773), .A(n7737), .B(n7736), .ZN(P2_U3167) );
  XNOR2_X1 U9037 ( .A(n7740), .B(n7739), .ZN(n10590) );
  XNOR2_X1 U9038 ( .A(n7741), .B(n6851), .ZN(n7742) );
  AOI222_X1 U9039 ( .A1(n9532), .A2(n7742), .B1(n7527), .B2(n9534), .C1(n9290), 
        .C2(n9609), .ZN(n10587) );
  OAI21_X1 U9040 ( .B1(n10586), .B2(n9618), .A(n10587), .ZN(n7743) );
  AOI21_X1 U9041 ( .B1(n10590), .B2(n9623), .A(n7743), .ZN(n10583) );
  INV_X1 U9042 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n7744) );
  OR2_X1 U9043 ( .A1(n9627), .A2(n7744), .ZN(n7745) );
  OAI21_X1 U9044 ( .B1(n10583), .B2(n9624), .A(n7745), .ZN(P2_U3461) );
  NOR2_X1 U9045 ( .A1(n10534), .A2(P1_U3973), .ZN(P1_U3085) );
  AOI211_X1 U9046 ( .C1(n7748), .C2(n7747), .A(n7746), .B(n9894), .ZN(n7757)
         );
  AOI211_X1 U9047 ( .C1(n7751), .C2(n7750), .A(n7749), .B(n9926), .ZN(n7756)
         );
  INV_X1 U9048 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n7754) );
  NAND2_X1 U9049 ( .A1(n10528), .A2(n7752), .ZN(n7753) );
  NAND2_X1 U9050 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n8761) );
  OAI211_X1 U9051 ( .C1(n7754), .C2(n9921), .A(n7753), .B(n8761), .ZN(n7755)
         );
  OR3_X1 U9052 ( .A1(n7757), .A2(n7756), .A3(n7755), .ZN(P1_U3254) );
  INV_X1 U9053 ( .A(n9881), .ZN(n9863) );
  INV_X1 U9054 ( .A(n7758), .ZN(n7760) );
  INV_X1 U9055 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n7759) );
  OAI222_X1 U9056 ( .A1(n9863), .A2(P1_U3086), .B1(n10293), .B2(n7760), .C1(
        n7759), .C2(n10290), .ZN(P1_U3339) );
  INV_X1 U9057 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n7889) );
  OAI222_X1 U9058 ( .A1(n9356), .A2(P2_U3151), .B1(n9676), .B2(n7760), .C1(
        n9137), .C2(n7889), .ZN(P2_U3279) );
  INV_X1 U9059 ( .A(n7761), .ZN(n7968) );
  NAND2_X1 U9060 ( .A1(n7762), .A2(n7961), .ZN(n7763) );
  AND2_X1 U9061 ( .A1(n7765), .A2(n7763), .ZN(n7767) );
  XNOR2_X1 U9062 ( .A(n7970), .B(n9115), .ZN(n7870) );
  XNOR2_X1 U9063 ( .A(n7870), .B(n9287), .ZN(n7766) );
  AND2_X1 U9064 ( .A1(n7766), .A2(n7763), .ZN(n7764) );
  OAI211_X1 U9065 ( .C1(n7767), .C2(n7766), .A(n7873), .B(n9256), .ZN(n7772)
         );
  NAND2_X1 U9066 ( .A1(n9238), .A2(n9286), .ZN(n7769) );
  INV_X1 U9067 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n8615) );
  NOR2_X1 U9068 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8615), .ZN(n10413) );
  INV_X1 U9069 ( .A(n10413), .ZN(n7768) );
  OAI211_X1 U9070 ( .C1(n7961), .C2(n9240), .A(n7769), .B(n7768), .ZN(n7770)
         );
  AOI21_X1 U9071 ( .B1(n7970), .B2(n9251), .A(n7770), .ZN(n7771) );
  OAI211_X1 U9072 ( .C1(n7968), .C2(n7773), .A(n7772), .B(n7771), .ZN(P2_U3179) );
  NAND2_X1 U9073 ( .A1(n7775), .A2(n7774), .ZN(n10683) );
  OAI22_X1 U9074 ( .A1(n9509), .A2(n6508), .B1(n10677), .B2(n7776), .ZN(n7779)
         );
  MUX2_X1 U9075 ( .A(n7777), .B(P2_REG2_REG_1__SCAN_IN), .S(n10687), .Z(n7778)
         );
  AOI211_X1 U9076 ( .C1(n9547), .C2(n7780), .A(n7779), .B(n7778), .ZN(n7781)
         );
  INV_X1 U9077 ( .A(n7781), .ZN(P2_U3232) );
  NAND2_X1 U9078 ( .A1(n10641), .A2(n9609), .ZN(n9545) );
  AOI22_X1 U9079 ( .A1(n10636), .A2(n7783), .B1(n10634), .B2(n7782), .ZN(n7784) );
  OAI21_X1 U9080 ( .B1(n6853), .B2(n9545), .A(n7784), .ZN(n7787) );
  MUX2_X1 U9081 ( .A(n7785), .B(P2_REG2_REG_3__SCAN_IN), .S(n10687), .Z(n7786)
         );
  AOI211_X1 U9082 ( .C1(n9547), .C2(n7788), .A(n7787), .B(n7786), .ZN(n7789)
         );
  INV_X1 U9083 ( .A(n7789), .ZN(P2_U3230) );
  XNOR2_X1 U9084 ( .A(n6853), .B(n5150), .ZN(n8878) );
  XNOR2_X1 U9085 ( .A(n7790), .B(n8878), .ZN(n7851) );
  OAI22_X1 U9086 ( .A1(n7961), .A2(n9616), .B1(n5150), .B2(n9618), .ZN(n7794)
         );
  XOR2_X1 U9087 ( .A(n7791), .B(n8878), .Z(n7793) );
  OAI22_X1 U9088 ( .A1(n7793), .A2(n9498), .B1(n7792), .B2(n9515), .ZN(n7848)
         );
  AOI211_X1 U9089 ( .C1(n9623), .C2(n7851), .A(n7794), .B(n7848), .ZN(n10602)
         );
  OR2_X1 U9090 ( .A1(n10602), .A2(n9624), .ZN(n7795) );
  OAI21_X1 U9091 ( .B1(n9627), .B2(n7207), .A(n7795), .ZN(P2_U3463) );
  OAI21_X1 U9092 ( .B1(n7798), .B2(n7797), .A(n7796), .ZN(n7808) );
  OAI21_X1 U9093 ( .B1(n7801), .B2(n7800), .A(n7799), .ZN(n7802) );
  NAND2_X1 U9094 ( .A1(n7802), .A2(n10519), .ZN(n7805) );
  NOR2_X1 U9095 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7803), .ZN(n8709) );
  AOI21_X1 U9096 ( .B1(n10534), .B2(P1_ADDR_REG_12__SCAN_IN), .A(n8709), .ZN(
        n7804) );
  OAI211_X1 U9097 ( .C1(n9887), .C2(n7806), .A(n7805), .B(n7804), .ZN(n7807)
         );
  AOI21_X1 U9098 ( .B1(n7808), .B2(n10524), .A(n7807), .ZN(n7809) );
  INV_X1 U9099 ( .A(n7809), .ZN(P1_U3255) );
  AOI22_X1 U9100 ( .A1(n9788), .A2(n7812), .B1(n9786), .B2(n6970), .ZN(n7815)
         );
  NAND2_X1 U9101 ( .A1(P1_U3086), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n9845) );
  INV_X1 U9102 ( .A(n9845), .ZN(n7813) );
  AOI21_X1 U9103 ( .B1(n9787), .B2(n6987), .A(n7813), .ZN(n7814) );
  OAI211_X1 U9104 ( .C1(n10593), .C2(n8745), .A(n7815), .B(n7814), .ZN(n7816)
         );
  AOI21_X1 U9105 ( .B1(n7817), .B2(n9784), .A(n7816), .ZN(n7818) );
  INV_X1 U9106 ( .A(n7818), .ZN(P1_U3218) );
  INV_X1 U9107 ( .A(n7819), .ZN(n7821) );
  NAND2_X1 U9108 ( .A1(n7821), .A2(n7820), .ZN(n7830) );
  INV_X1 U9109 ( .A(n10619), .ZN(n7834) );
  NOR3_X1 U9110 ( .A1(n7824), .A2(n7823), .A3(n7822), .ZN(n7828) );
  INV_X1 U9111 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n7826) );
  OAI21_X1 U9112 ( .B1(n10606), .B2(n7826), .A(n7825), .ZN(n7827) );
  OAI21_X1 U9113 ( .B1(n7828), .B2(n7827), .A(n7834), .ZN(n7833) );
  NOR2_X2 U9114 ( .A1(n7830), .A2(n9923), .ZN(n10576) );
  OAI21_X1 U9115 ( .B1(n10570), .B2(n10002), .A(n7831), .ZN(n7832) );
  OAI211_X1 U9116 ( .C1(n9820), .C2(n7834), .A(n7833), .B(n7832), .ZN(P1_U3293) );
  NAND2_X1 U9117 ( .A1(n7835), .A2(n9784), .ZN(n7844) );
  AOI21_X1 U9118 ( .B1(n7810), .B2(n7837), .A(n7836), .ZN(n7843) );
  AOI22_X1 U9119 ( .A1(n9788), .A2(n8015), .B1(n9786), .B2(n10559), .ZN(n7842)
         );
  INV_X1 U9120 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n7839) );
  NOR2_X1 U9121 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7839), .ZN(n10533) );
  NOR2_X1 U9122 ( .A1(n8745), .A2(n8115), .ZN(n7840) );
  AOI211_X1 U9123 ( .C1(n9787), .C2(n9808), .A(n10533), .B(n7840), .ZN(n7841)
         );
  OAI211_X1 U9124 ( .C1(n7844), .C2(n7843), .A(n7842), .B(n7841), .ZN(P1_U3230) );
  AOI22_X1 U9125 ( .A1(n10636), .A2(n7846), .B1(n10634), .B2(n7845), .ZN(n7847) );
  OAI21_X1 U9126 ( .B1(n7961), .B2(n9545), .A(n7847), .ZN(n7850) );
  MUX2_X1 U9127 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n7848), .S(n10641), .Z(n7849)
         );
  AOI211_X1 U9128 ( .C1(n9547), .C2(n7851), .A(n7850), .B(n7849), .ZN(n7852)
         );
  INV_X1 U9129 ( .A(n7852), .ZN(P2_U3229) );
  XNOR2_X1 U9130 ( .A(n7853), .B(n7864), .ZN(n10540) );
  OR2_X1 U9131 ( .A1(n7854), .A2(n6070), .ZN(n7855) );
  NOR2_X1 U9132 ( .A1(n7834), .A2(n7856), .ZN(n7860) );
  INV_X1 U9133 ( .A(n10576), .ZN(n10608) );
  OAI211_X1 U9134 ( .C1(n6965), .C2(n7857), .A(n10552), .B(n10550), .ZN(n10541) );
  INV_X1 U9135 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n7858) );
  OAI22_X1 U9136 ( .A1(n10608), .A2(n10541), .B1(n7858), .B2(n10606), .ZN(
        n7859) );
  AOI211_X1 U9137 ( .C1(n10570), .C2(n7861), .A(n7860), .B(n7859), .ZN(n7869)
         );
  AOI22_X1 U9138 ( .A1(n10557), .A2(n7932), .B1(n6970), .B2(n10558), .ZN(n7867) );
  OAI21_X1 U9139 ( .B1(n7864), .B2(n7863), .A(n7862), .ZN(n7865) );
  NAND2_X1 U9140 ( .A1(n7865), .A2(n10127), .ZN(n7866) );
  OAI211_X1 U9141 ( .C1(n10540), .C2(n8028), .A(n7867), .B(n7866), .ZN(n10542)
         );
  NAND2_X1 U9142 ( .A1(n10542), .A2(n7834), .ZN(n7868) );
  OAI211_X1 U9143 ( .C1(n10540), .C2(n10573), .A(n7869), .B(n7868), .ZN(
        P1_U3292) );
  INV_X1 U9144 ( .A(n7870), .ZN(n7871) );
  NAND2_X1 U9145 ( .A1(n7871), .A2(n9287), .ZN(n7872) );
  XNOR2_X1 U9146 ( .A(n8096), .B(n9110), .ZN(n7999) );
  XNOR2_X1 U9147 ( .A(n7999), .B(n9286), .ZN(n7875) );
  INV_X1 U9148 ( .A(n7875), .ZN(n7874) );
  NAND2_X1 U9149 ( .A1(n7876), .A2(n7875), .ZN(n7877) );
  AOI21_X1 U9150 ( .B1(n8002), .B2(n7877), .A(n9254), .ZN(n7884) );
  NAND2_X1 U9151 ( .A1(P2_U3151), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n10444) );
  INV_X1 U9152 ( .A(n10444), .ZN(n7878) );
  AOI21_X1 U9153 ( .B1(n9285), .B2(n9238), .A(n7878), .ZN(n7882) );
  NAND2_X1 U9154 ( .A1(n8096), .A2(n9251), .ZN(n7881) );
  NAND2_X1 U9155 ( .A1(n9266), .A2(n8063), .ZN(n7880) );
  NAND2_X1 U9156 ( .A1(n9261), .A2(n9287), .ZN(n7879) );
  NAND4_X1 U9157 ( .A1(n7882), .A2(n7881), .A3(n7880), .A4(n7879), .ZN(n7883)
         );
  OR2_X1 U9158 ( .A1(n7884), .A2(n7883), .ZN(P2_U3153) );
  INV_X1 U9159 ( .A(n7885), .ZN(n7918) );
  INV_X1 U9160 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n7891) );
  OAI222_X1 U9161 ( .A1(n9676), .A2(n7918), .B1(n9137), .B2(n7891), .C1(
        P2_U3151), .C2(n9373), .ZN(P2_U3278) );
  NAND2_X1 U9162 ( .A1(n8286), .A2(P1_U3973), .ZN(n7886) );
  OAI21_X1 U9163 ( .B1(n7887), .B2(P1_U3973), .A(n7886), .ZN(P1_U3562) );
  NAND2_X1 U9164 ( .A1(n9723), .A2(P1_U3973), .ZN(n7888) );
  OAI21_X1 U9165 ( .B1(n7889), .B2(P1_U3973), .A(n7888), .ZN(P1_U3570) );
  NAND2_X1 U9166 ( .A1(n9773), .A2(P1_U3973), .ZN(n7890) );
  OAI21_X1 U9167 ( .B1(n7891), .B2(P1_U3973), .A(n7890), .ZN(P1_U3571) );
  INV_X1 U9168 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n8210) );
  NAND2_X1 U9169 ( .A1(n9698), .A2(P1_U3973), .ZN(n7892) );
  OAI21_X1 U9170 ( .B1(n8210), .B2(P1_U3973), .A(n7892), .ZN(P1_U3574) );
  INV_X1 U9171 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n8089) );
  INV_X1 U9172 ( .A(n10111), .ZN(n7893) );
  NAND2_X1 U9173 ( .A1(n7893), .A2(P1_U3973), .ZN(n7894) );
  OAI21_X1 U9174 ( .B1(n8089), .B2(P1_U3973), .A(n7894), .ZN(P1_U3573) );
  INV_X1 U9175 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n9136) );
  NAND2_X1 U9176 ( .A1(n9706), .A2(P1_U3973), .ZN(n7895) );
  OAI21_X1 U9177 ( .B1(n9136), .B2(P1_U3973), .A(n7895), .ZN(P1_U3578) );
  OAI222_X1 U9178 ( .A1(n10290), .A2(n7896), .B1(n10293), .B2(n7919), .C1(
        P1_U3086), .C2(n9893), .ZN(P1_U3337) );
  NOR2_X1 U9179 ( .A1(P2_ADDR_REG_18__SCAN_IN), .A2(P1_ADDR_REG_18__SCAN_IN), 
        .ZN(n7897) );
  AOI21_X1 U9180 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(P2_ADDR_REG_18__SCAN_IN), 
        .A(n7897), .ZN(n10352) );
  NOR2_X1 U9181 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n7898) );
  AOI21_X1 U9182 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n7898), .ZN(n10349) );
  NOR2_X1 U9183 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n7899) );
  AOI21_X1 U9184 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n7899), .ZN(n10346) );
  NOR2_X1 U9185 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n7900) );
  AOI21_X1 U9186 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n7900), .ZN(n10343) );
  NOR2_X1 U9187 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n7901) );
  AOI21_X1 U9188 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n7901), .ZN(n10340) );
  NOR2_X1 U9189 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n7902) );
  AOI21_X1 U9190 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n7902), .ZN(n10337) );
  NOR2_X1 U9191 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n7903) );
  AOI21_X1 U9192 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n7903), .ZN(n10334) );
  NOR2_X1 U9193 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n7904) );
  AOI21_X1 U9194 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n7904), .ZN(n10331) );
  NOR2_X1 U9195 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n7905) );
  AOI21_X1 U9196 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n7905), .ZN(n10328) );
  NOR2_X1 U9197 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n7906) );
  AOI21_X1 U9198 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(P2_ADDR_REG_9__SCAN_IN), 
        .A(n7906), .ZN(n10325) );
  NOR2_X1 U9199 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n7907) );
  AOI21_X1 U9200 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(P2_ADDR_REG_8__SCAN_IN), 
        .A(n7907), .ZN(n10322) );
  NOR2_X1 U9201 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n7908) );
  AOI21_X1 U9202 ( .B1(P1_ADDR_REG_7__SCAN_IN), .B2(P2_ADDR_REG_7__SCAN_IN), 
        .A(n7908), .ZN(n10319) );
  NOR2_X1 U9203 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(P1_ADDR_REG_6__SCAN_IN), 
        .ZN(n7909) );
  AOI21_X1 U9204 ( .B1(P1_ADDR_REG_6__SCAN_IN), .B2(P2_ADDR_REG_6__SCAN_IN), 
        .A(n7909), .ZN(n10316) );
  NOR2_X1 U9205 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n7910) );
  AOI21_X1 U9206 ( .B1(P1_ADDR_REG_5__SCAN_IN), .B2(P2_ADDR_REG_5__SCAN_IN), 
        .A(n7910), .ZN(n10313) );
  NAND2_X1 U9207 ( .A1(P2_ADDR_REG_0__SCAN_IN), .A2(P1_ADDR_REG_0__SCAN_IN), 
        .ZN(n10299) );
  INV_X1 U9208 ( .A(n10299), .ZN(n7911) );
  INV_X1 U9209 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10300) );
  NAND2_X1 U9210 ( .A1(n10300), .A2(n10299), .ZN(n10298) );
  AOI22_X1 U9211 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(n7911), .B1(
        P2_ADDR_REG_1__SCAN_IN), .B2(n10298), .ZN(n10304) );
  NAND2_X1 U9212 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n7912) );
  OAI21_X1 U9213 ( .B1(P1_ADDR_REG_2__SCAN_IN), .B2(P2_ADDR_REG_2__SCAN_IN), 
        .A(n7912), .ZN(n10303) );
  NOR2_X1 U9214 ( .A1(n10304), .A2(n10303), .ZN(n10302) );
  AOI21_X1 U9215 ( .B1(P2_ADDR_REG_2__SCAN_IN), .B2(P1_ADDR_REG_2__SCAN_IN), 
        .A(n10302), .ZN(n10307) );
  NAND2_X1 U9216 ( .A1(P2_ADDR_REG_3__SCAN_IN), .A2(P1_ADDR_REG_3__SCAN_IN), 
        .ZN(n7913) );
  OAI21_X1 U9217 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(P1_ADDR_REG_3__SCAN_IN), 
        .A(n7913), .ZN(n10306) );
  NOR2_X1 U9218 ( .A1(n10307), .A2(n10306), .ZN(n10305) );
  AOI21_X1 U9219 ( .B1(P1_ADDR_REG_3__SCAN_IN), .B2(P2_ADDR_REG_3__SCAN_IN), 
        .A(n10305), .ZN(n10310) );
  NOR2_X1 U9220 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n7914) );
  AOI21_X1 U9221 ( .B1(P2_ADDR_REG_4__SCAN_IN), .B2(P1_ADDR_REG_4__SCAN_IN), 
        .A(n7914), .ZN(n10309) );
  NAND2_X1 U9222 ( .A1(n10310), .A2(n10309), .ZN(n10308) );
  OAI21_X1 U9223 ( .B1(P1_ADDR_REG_4__SCAN_IN), .B2(P2_ADDR_REG_4__SCAN_IN), 
        .A(n10308), .ZN(n10312) );
  NAND2_X1 U9224 ( .A1(n10313), .A2(n10312), .ZN(n10311) );
  OAI21_X1 U9225 ( .B1(P2_ADDR_REG_5__SCAN_IN), .B2(P1_ADDR_REG_5__SCAN_IN), 
        .A(n10311), .ZN(n10315) );
  NAND2_X1 U9226 ( .A1(n10316), .A2(n10315), .ZN(n10314) );
  OAI21_X1 U9227 ( .B1(P2_ADDR_REG_6__SCAN_IN), .B2(P1_ADDR_REG_6__SCAN_IN), 
        .A(n10314), .ZN(n10318) );
  NAND2_X1 U9228 ( .A1(n10319), .A2(n10318), .ZN(n10317) );
  OAI21_X1 U9229 ( .B1(P2_ADDR_REG_7__SCAN_IN), .B2(P1_ADDR_REG_7__SCAN_IN), 
        .A(n10317), .ZN(n10321) );
  NAND2_X1 U9230 ( .A1(n10322), .A2(n10321), .ZN(n10320) );
  OAI21_X1 U9231 ( .B1(P2_ADDR_REG_8__SCAN_IN), .B2(P1_ADDR_REG_8__SCAN_IN), 
        .A(n10320), .ZN(n10324) );
  NAND2_X1 U9232 ( .A1(n10325), .A2(n10324), .ZN(n10323) );
  OAI21_X1 U9233 ( .B1(P2_ADDR_REG_9__SCAN_IN), .B2(P1_ADDR_REG_9__SCAN_IN), 
        .A(n10323), .ZN(n10327) );
  NAND2_X1 U9234 ( .A1(n10328), .A2(n10327), .ZN(n10326) );
  OAI21_X1 U9235 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n10326), .ZN(n10330) );
  NAND2_X1 U9236 ( .A1(n10331), .A2(n10330), .ZN(n10329) );
  OAI21_X1 U9237 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n10329), .ZN(n10333) );
  NAND2_X1 U9238 ( .A1(n10334), .A2(n10333), .ZN(n10332) );
  OAI21_X1 U9239 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10332), .ZN(n10336) );
  NAND2_X1 U9240 ( .A1(n10337), .A2(n10336), .ZN(n10335) );
  OAI21_X1 U9241 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n10335), .ZN(n10339) );
  NAND2_X1 U9242 ( .A1(n10340), .A2(n10339), .ZN(n10338) );
  OAI21_X1 U9243 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10338), .ZN(n10342) );
  NAND2_X1 U9244 ( .A1(n10343), .A2(n10342), .ZN(n10341) );
  OAI21_X1 U9245 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n10341), .ZN(n10345) );
  NAND2_X1 U9246 ( .A1(n10346), .A2(n10345), .ZN(n10344) );
  OAI21_X1 U9247 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n10344), .ZN(n10348) );
  NAND2_X1 U9248 ( .A1(n10349), .A2(n10348), .ZN(n10347) );
  OAI21_X1 U9249 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10347), .ZN(n10351) );
  NAND2_X1 U9250 ( .A1(n10352), .A2(n10351), .ZN(n10350) );
  OAI21_X1 U9251 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(P1_ADDR_REG_18__SCAN_IN), 
        .A(n10350), .ZN(n7916) );
  XNOR2_X1 U9252 ( .A(n9920), .B(P2_ADDR_REG_19__SCAN_IN), .ZN(n7915) );
  XNOR2_X1 U9253 ( .A(n7916), .B(n7915), .ZN(ADD_1068_U4) );
  OAI222_X1 U9254 ( .A1(P1_U3086), .A2(n9886), .B1(n10293), .B2(n7918), .C1(
        n7917), .C2(n10290), .ZN(P1_U3338) );
  INV_X1 U9255 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n7920) );
  OAI222_X1 U9256 ( .A1(n9137), .A2(n7920), .B1(n9391), .B2(P2_U3151), .C1(
        n9676), .C2(n7919), .ZN(P2_U3277) );
  XNOR2_X1 U9257 ( .A(n7922), .B(n7921), .ZN(n7923) );
  XNOR2_X1 U9258 ( .A(n7924), .B(n7923), .ZN(n7931) );
  AOI22_X1 U9259 ( .A1(n7925), .A2(n9788), .B1(n9786), .B2(n6987), .ZN(n7930)
         );
  OAI21_X1 U9260 ( .B1(n9775), .B2(n8136), .A(n7926), .ZN(n7927) );
  AOI21_X1 U9261 ( .B1(n7928), .B2(n9789), .A(n7927), .ZN(n7929) );
  OAI211_X1 U9262 ( .C1(n7931), .C2(n9778), .A(n7930), .B(n7929), .ZN(P1_U3227) );
  NAND2_X1 U9263 ( .A1(n7932), .A2(P1_U3973), .ZN(n7933) );
  OAI21_X1 U9264 ( .B1(P1_U3973), .B2(n5522), .A(n7933), .ZN(P1_U3554) );
  NAND2_X1 U9265 ( .A1(n7934), .A2(n8937), .ZN(n7935) );
  XOR2_X1 U9266 ( .A(n8879), .B(n7935), .Z(n8045) );
  INV_X1 U9267 ( .A(n8045), .ZN(n7943) );
  XNOR2_X1 U9268 ( .A(n7936), .B(n8879), .ZN(n7937) );
  AOI222_X1 U9269 ( .A1(n9532), .A2(n7937), .B1(n9287), .B2(n9609), .C1(n9289), 
        .C2(n9534), .ZN(n8042) );
  MUX2_X1 U9270 ( .A(n7938), .B(n8042), .S(n10641), .Z(n7942) );
  AOI22_X1 U9271 ( .A1(n10636), .A2(n7940), .B1(n10634), .B2(n7939), .ZN(n7941) );
  OAI211_X1 U9272 ( .C1(n7943), .C2(n9493), .A(n7942), .B(n7941), .ZN(P2_U3228) );
  INV_X1 U9273 ( .A(n7946), .ZN(n7950) );
  XNOR2_X1 U9274 ( .A(n7944), .B(n7950), .ZN(n10605) );
  OR2_X1 U9275 ( .A1(n7974), .A2(n7981), .ZN(n7976) );
  NAND2_X1 U9276 ( .A1(n7976), .A2(n7945), .ZN(n7991) );
  INV_X1 U9277 ( .A(n7991), .ZN(n7948) );
  NOR3_X1 U9278 ( .A1(n7948), .A2(n7947), .A3(n7946), .ZN(n7949) );
  AOI211_X1 U9279 ( .C1(n7951), .C2(n7950), .A(n10561), .B(n7949), .ZN(n7955)
         );
  INV_X1 U9280 ( .A(n6987), .ZN(n7952) );
  OAI22_X1 U9281 ( .A1(n7952), .A2(n10143), .B1(n8136), .B2(n10145), .ZN(n7953) );
  AOI21_X1 U9282 ( .B1(n7955), .B2(n7954), .A(n7953), .ZN(n10618) );
  OAI211_X1 U9283 ( .C1(n7995), .C2(n10613), .A(n10552), .B(n8034), .ZN(n10609) );
  OAI211_X1 U9284 ( .C1(n10239), .C2(n10605), .A(n10618), .B(n10609), .ZN(
        n8121) );
  INV_X1 U9285 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n7956) );
  OAI22_X1 U9286 ( .A1(n10267), .A2(n10613), .B1(n10674), .B2(n7956), .ZN(
        n7957) );
  AOI21_X1 U9287 ( .B1(n8121), .B2(n10674), .A(n7957), .ZN(n7958) );
  INV_X1 U9288 ( .A(n7958), .ZN(P1_U3468) );
  NAND2_X1 U9289 ( .A1(n8950), .A2(n8947), .ZN(n8882) );
  XNOR2_X1 U9290 ( .A(n7959), .B(n8882), .ZN(n7960) );
  OAI222_X1 U9291 ( .A1(n9616), .A2(n8010), .B1(n9515), .B2(n7961), .C1(n7960), 
        .C2(n9498), .ZN(n7967) );
  XNOR2_X1 U9292 ( .A(n7962), .B(n8882), .ZN(n7973) );
  OAI22_X1 U9293 ( .A1(n7973), .A2(n9615), .B1(n7963), .B2(n9618), .ZN(n7964)
         );
  NOR2_X1 U9294 ( .A1(n7967), .A2(n7964), .ZN(n10621) );
  INV_X1 U9295 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n7965) );
  OR2_X1 U9296 ( .A1(n9627), .A2(n7965), .ZN(n7966) );
  OAI21_X1 U9297 ( .B1(n10621), .B2(n9624), .A(n7966), .ZN(P2_U3465) );
  NAND2_X1 U9298 ( .A1(n7967), .A2(n10641), .ZN(n7972) );
  OAI22_X1 U9299 ( .A1(n10641), .A2(n7247), .B1(n7968), .B2(n10677), .ZN(n7969) );
  AOI21_X1 U9300 ( .B1(n10636), .B2(n7970), .A(n7969), .ZN(n7971) );
  OAI211_X1 U9301 ( .C1(n7973), .C2(n9493), .A(n7972), .B(n7971), .ZN(P2_U3227) );
  NAND2_X1 U9302 ( .A1(n7974), .A2(n7981), .ZN(n7975) );
  NAND2_X1 U9303 ( .A1(n7976), .A2(n7975), .ZN(n7977) );
  NAND2_X1 U9304 ( .A1(n7977), .A2(n10127), .ZN(n7979) );
  AOI22_X1 U9305 ( .A1(n10558), .A2(n6987), .B1(n6970), .B2(n10557), .ZN(n7978) );
  NAND2_X1 U9306 ( .A1(n7979), .A2(n7978), .ZN(n10594) );
  INV_X1 U9307 ( .A(n10594), .ZN(n7988) );
  OR2_X1 U9308 ( .A1(n10619), .A2(n8028), .ZN(n7980) );
  XNOR2_X1 U9309 ( .A(n7982), .B(n7981), .ZN(n10596) );
  INV_X1 U9310 ( .A(n7993), .ZN(n7983) );
  OAI211_X1 U9311 ( .C1(n10593), .C2(n10551), .A(n7983), .B(n10552), .ZN(
        n10592) );
  OAI22_X1 U9312 ( .A1(n10592), .A2(n10608), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        n10606), .ZN(n7984) );
  AOI21_X1 U9313 ( .B1(P1_REG2_REG_3__SCAN_IN), .B2(n4941), .A(n7984), .ZN(
        n7985) );
  OAI21_X1 U9314 ( .B1(n10593), .B2(n10612), .A(n7985), .ZN(n7986) );
  AOI21_X1 U9315 ( .B1(n10615), .B2(n10596), .A(n7986), .ZN(n7987) );
  OAI21_X1 U9316 ( .B1(n4941), .B2(n7988), .A(n7987), .ZN(P1_U3290) );
  XNOR2_X1 U9317 ( .A(n7989), .B(n7990), .ZN(n8019) );
  XNOR2_X1 U9318 ( .A(n7991), .B(n7990), .ZN(n7992) );
  AOI222_X1 U9319 ( .A1(n10127), .A2(n7992), .B1(n10559), .B2(n10557), .C1(
        n9808), .C2(n10558), .ZN(n8024) );
  OAI21_X1 U9320 ( .B1(n7993), .B2(n8115), .A(n10552), .ZN(n7994) );
  OR2_X1 U9321 ( .A1(n7995), .A2(n7994), .ZN(n8014) );
  OAI211_X1 U9322 ( .C1(n10239), .C2(n8019), .A(n8024), .B(n8014), .ZN(n8117)
         );
  INV_X1 U9323 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n7996) );
  OAI22_X1 U9324 ( .A1(n10267), .A2(n8115), .B1(n10674), .B2(n7996), .ZN(n7997) );
  AOI21_X1 U9325 ( .B1(n8117), .B2(n10674), .A(n7997), .ZN(n7998) );
  INV_X1 U9326 ( .A(n7998), .ZN(P1_U3465) );
  INV_X1 U9327 ( .A(n7999), .ZN(n8000) );
  NAND2_X1 U9328 ( .A1(n8000), .A2(n8010), .ZN(n8001) );
  XNOR2_X1 U9329 ( .A(n10637), .B(n9115), .ZN(n8003) );
  AND2_X1 U9330 ( .A1(n8003), .A2(n8192), .ZN(n8124) );
  INV_X1 U9331 ( .A(n8124), .ZN(n8005) );
  INV_X1 U9332 ( .A(n8003), .ZN(n8004) );
  NAND2_X1 U9333 ( .A1(n8004), .A2(n9285), .ZN(n8123) );
  NAND2_X1 U9334 ( .A1(n8005), .A2(n8123), .ZN(n8006) );
  XNOR2_X1 U9335 ( .A(n8125), .B(n8006), .ZN(n8013) );
  NAND2_X1 U9336 ( .A1(n9266), .A2(n10635), .ZN(n8009) );
  NAND2_X1 U9337 ( .A1(P2_U3151), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n10460) );
  INV_X1 U9338 ( .A(n10460), .ZN(n8007) );
  AOI21_X1 U9339 ( .B1(n9238), .B2(n9284), .A(n8007), .ZN(n8008) );
  OAI211_X1 U9340 ( .C1(n8010), .C2(n9240), .A(n8009), .B(n8008), .ZN(n8011)
         );
  AOI21_X1 U9341 ( .B1(n10637), .B2(n9251), .A(n8011), .ZN(n8012) );
  OAI21_X1 U9342 ( .B1(n8013), .B2(n9254), .A(n8012), .ZN(P2_U3161) );
  INV_X1 U9343 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n8018) );
  INV_X1 U9344 ( .A(n8014), .ZN(n8016) );
  AOI22_X1 U9345 ( .A1(n8016), .A2(n10576), .B1(n8015), .B2(n10572), .ZN(n8017) );
  OAI21_X1 U9346 ( .B1(n8018), .B2(n7834), .A(n8017), .ZN(n8021) );
  NOR2_X1 U9347 ( .A1(n8019), .A2(n10154), .ZN(n8020) );
  AOI211_X1 U9348 ( .C1(n10570), .C2(n8022), .A(n8021), .B(n8020), .ZN(n8023)
         );
  OAI21_X1 U9349 ( .B1(n8024), .B2(n4941), .A(n8023), .ZN(P1_U3289) );
  OAI21_X1 U9350 ( .B1(n8026), .B2(n8027), .A(n8025), .ZN(n10626) );
  INV_X1 U9351 ( .A(n10626), .ZN(n8041) );
  XOR2_X1 U9352 ( .A(n8074), .B(n8027), .Z(n8033) );
  INV_X1 U9353 ( .A(n8028), .ZN(n10564) );
  OAI22_X1 U9354 ( .A1(n8030), .A2(n10143), .B1(n8029), .B2(n10145), .ZN(n8031) );
  AOI21_X1 U9355 ( .B1(n10626), .B2(n10564), .A(n8031), .ZN(n8032) );
  OAI21_X1 U9356 ( .B1(n8033), .B2(n10561), .A(n8032), .ZN(n10624) );
  NAND2_X1 U9357 ( .A1(n10624), .A2(n7834), .ZN(n8040) );
  INV_X1 U9358 ( .A(n8034), .ZN(n8035) );
  OAI211_X1 U9359 ( .C1(n8035), .C2(n10623), .A(n10552), .B(n8143), .ZN(n10622) );
  AOI22_X1 U9360 ( .A1(n4941), .A2(P1_REG2_REG_6__SCAN_IN), .B1(n8053), .B2(
        n10572), .ZN(n8036) );
  OAI21_X1 U9361 ( .B1(n10622), .B2(n10608), .A(n8036), .ZN(n8037) );
  AOI21_X1 U9362 ( .B1(n10570), .B2(n8038), .A(n8037), .ZN(n8039) );
  OAI211_X1 U9363 ( .C1(n8041), .C2(n10573), .A(n8040), .B(n8039), .ZN(
        P1_U3287) );
  OAI21_X1 U9364 ( .B1(n8043), .B2(n9618), .A(n8042), .ZN(n8044) );
  AOI21_X1 U9365 ( .B1(n9623), .B2(n8045), .A(n8044), .ZN(n10604) );
  NAND2_X1 U9366 ( .A1(n9624), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n8046) );
  OAI21_X1 U9367 ( .B1(n10604), .B2(n9624), .A(n8046), .ZN(P2_U3464) );
  NAND2_X1 U9368 ( .A1(n8048), .A2(n8047), .ZN(n8052) );
  NOR2_X1 U9369 ( .A1(n5056), .A2(n8050), .ZN(n8051) );
  XNOR2_X1 U9370 ( .A(n8052), .B(n8051), .ZN(n8059) );
  AOI22_X1 U9371 ( .A1(n8053), .A2(n9788), .B1(n9786), .B2(n9808), .ZN(n8058)
         );
  INV_X1 U9372 ( .A(n8054), .ZN(n8056) );
  NOR2_X1 U9373 ( .A1(n8745), .A2(n10623), .ZN(n8055) );
  AOI211_X1 U9374 ( .C1(n9787), .C2(n9806), .A(n8056), .B(n8055), .ZN(n8057)
         );
  OAI211_X1 U9375 ( .C1(n8059), .C2(n9778), .A(n8058), .B(n8057), .ZN(P1_U3239) );
  XNOR2_X1 U9376 ( .A(n8060), .B(n8885), .ZN(n8061) );
  OAI22_X1 U9377 ( .A1(n8061), .A2(n9498), .B1(n6575), .B2(n9515), .ZN(n8094)
         );
  OAI21_X1 U9378 ( .B1(n8062), .B2(n8885), .A(n8295), .ZN(n8092) );
  INV_X1 U9379 ( .A(n9545), .ZN(n9470) );
  INV_X1 U9380 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n8065) );
  INV_X1 U9381 ( .A(n8063), .ZN(n8064) );
  OAI22_X1 U9382 ( .A1(n10641), .A2(n8065), .B1(n8064), .B2(n10677), .ZN(n8066) );
  AOI21_X1 U9383 ( .B1(n9470), .B2(n9285), .A(n8066), .ZN(n8068) );
  NAND2_X1 U9384 ( .A1(n10636), .A2(n8096), .ZN(n8067) );
  OAI211_X1 U9385 ( .C1(n8092), .C2(n9493), .A(n8068), .B(n8067), .ZN(n8069)
         );
  AOI21_X1 U9386 ( .B1(n8094), .B2(n10641), .A(n8069), .ZN(n8070) );
  INV_X1 U9387 ( .A(n8070), .ZN(P2_U3226) );
  INV_X1 U9388 ( .A(n8071), .ZN(n8072) );
  AOI21_X1 U9389 ( .B1(n8074), .B2(n8073), .A(n8072), .ZN(n8138) );
  AOI21_X1 U9390 ( .B1(n8138), .B2(n5449), .A(n8075), .ZN(n8076) );
  NAND2_X1 U9391 ( .A1(n8076), .A2(n4945), .ZN(n8174) );
  OAI211_X1 U9392 ( .C1(n8076), .C2(n4945), .A(n8174), .B(n10127), .ZN(n8078)
         );
  AOI22_X1 U9393 ( .A1(n10558), .A2(n5343), .B1(n9806), .B2(n10557), .ZN(n8077) );
  NAND2_X1 U9394 ( .A1(n8078), .A2(n8077), .ZN(n8203) );
  INV_X1 U9395 ( .A(n8203), .ZN(n8087) );
  OAI21_X1 U9396 ( .B1(n8081), .B2(n8080), .A(n8079), .ZN(n8205) );
  INV_X1 U9397 ( .A(n8142), .ZN(n8082) );
  AOI211_X1 U9398 ( .C1(n8167), .C2(n8082), .A(n10663), .B(n8253), .ZN(n8204)
         );
  NAND2_X1 U9399 ( .A1(n8204), .A2(n10576), .ZN(n8084) );
  AOI22_X1 U9400 ( .A1(n10619), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n8163), .B2(
        n10572), .ZN(n8083) );
  OAI211_X1 U9401 ( .C1(n5744), .C2(n10612), .A(n8084), .B(n8083), .ZN(n8085)
         );
  AOI21_X1 U9402 ( .B1(n8205), .B2(n10615), .A(n8085), .ZN(n8086) );
  OAI21_X1 U9403 ( .B1(n8087), .B2(n4941), .A(n8086), .ZN(P1_U3285) );
  INV_X1 U9404 ( .A(n8088), .ZN(n9135) );
  OAI222_X1 U9405 ( .A1(P2_U3151), .A2(n8090), .B1(n9676), .B2(n9135), .C1(
        n9137), .C2(n8089), .ZN(P2_U3276) );
  OAI22_X1 U9406 ( .A1(n8092), .A2(n9615), .B1(n8192), .B2(n9616), .ZN(n8093)
         );
  NOR2_X1 U9407 ( .A1(n8094), .A2(n8093), .ZN(n8101) );
  INV_X1 U9408 ( .A(n9594), .ZN(n8304) );
  AOI22_X1 U9409 ( .A1(n8304), .A2(n8096), .B1(n9624), .B2(
        P2_REG1_REG_7__SCAN_IN), .ZN(n8095) );
  OAI21_X1 U9410 ( .B1(n8101), .B2(n9624), .A(n8095), .ZN(P2_U3466) );
  INV_X1 U9411 ( .A(n8096), .ZN(n8098) );
  INV_X1 U9412 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n8097) );
  OAI22_X1 U9413 ( .A1(n9654), .A2(n8098), .B1(n10695), .B2(n8097), .ZN(n8099)
         );
  INV_X1 U9414 ( .A(n8099), .ZN(n8100) );
  OAI21_X1 U9415 ( .B1(n8101), .B2(n10692), .A(n8100), .ZN(P2_U3411) );
  AOI211_X1 U9416 ( .C1(n8104), .C2(n8103), .A(n8102), .B(n9894), .ZN(n8113)
         );
  AOI211_X1 U9417 ( .C1(n8107), .C2(n8106), .A(n8105), .B(n9926), .ZN(n8112)
         );
  INV_X1 U9418 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n8110) );
  NAND2_X1 U9419 ( .A1(n10528), .A2(n8108), .ZN(n8109) );
  NAND2_X1 U9420 ( .A1(P1_U3086), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n8738) );
  OAI211_X1 U9421 ( .C1(n8110), .C2(n9921), .A(n8109), .B(n8738), .ZN(n8111)
         );
  OR3_X1 U9422 ( .A1(n8113), .A2(n8112), .A3(n8111), .ZN(P1_U3256) );
  INV_X1 U9423 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n8114) );
  OAI22_X1 U9424 ( .A1(n10219), .A2(n8115), .B1(n10646), .B2(n8114), .ZN(n8116) );
  AOI21_X1 U9425 ( .B1(n8117), .B2(n10646), .A(n8116), .ZN(n8118) );
  INV_X1 U9426 ( .A(n8118), .ZN(P1_U3526) );
  INV_X1 U9427 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n8119) );
  OAI22_X1 U9428 ( .A1(n10219), .A2(n10613), .B1(n10646), .B2(n8119), .ZN(
        n8120) );
  AOI21_X1 U9429 ( .B1(n8121), .B2(n10646), .A(n8120), .ZN(n8122) );
  INV_X1 U9430 ( .A(n8122), .ZN(P1_U3527) );
  INV_X1 U9431 ( .A(n8241), .ZN(n8133) );
  XNOR2_X1 U9432 ( .A(n8241), .B(n9115), .ZN(n8260) );
  XNOR2_X1 U9433 ( .A(n8260), .B(n9284), .ZN(n8126) );
  OAI211_X1 U9434 ( .C1(n8127), .C2(n8126), .A(n8263), .B(n9256), .ZN(n8132)
         );
  NAND2_X1 U9435 ( .A1(P2_U3151), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n10476) );
  INV_X1 U9436 ( .A(n10476), .ZN(n8128) );
  AOI21_X1 U9437 ( .B1(n9238), .B2(n9283), .A(n8128), .ZN(n8129) );
  OAI21_X1 U9438 ( .B1(n8192), .B2(n9240), .A(n8129), .ZN(n8130) );
  AOI21_X1 U9439 ( .B1(n8195), .B2(n9266), .A(n8130), .ZN(n8131) );
  OAI211_X1 U9440 ( .C1(n8133), .C2(n9270), .A(n8132), .B(n8131), .ZN(P2_U3171) );
  OAI21_X1 U9441 ( .B1(n8135), .B2(n8137), .A(n8134), .ZN(n8145) );
  OAI22_X1 U9442 ( .A1(n8136), .A2(n10143), .B1(n8176), .B2(n10145), .ZN(n8141) );
  XNOR2_X1 U9443 ( .A(n8138), .B(n8137), .ZN(n8139) );
  NOR2_X1 U9444 ( .A1(n8139), .A2(n10561), .ZN(n8140) );
  AOI211_X1 U9445 ( .C1(n10564), .C2(n8145), .A(n8141), .B(n8140), .ZN(n8274)
         );
  AOI21_X1 U9446 ( .B1(n8271), .B2(n8143), .A(n8142), .ZN(n8272) );
  AOI22_X1 U9447 ( .A1(n10619), .A2(P1_REG2_REG_7__SCAN_IN), .B1(n8151), .B2(
        n10572), .ZN(n8144) );
  OAI21_X1 U9448 ( .B1(n10612), .B2(n8153), .A(n8144), .ZN(n8147) );
  INV_X1 U9449 ( .A(n8145), .ZN(n8275) );
  NOR2_X1 U9450 ( .A1(n8275), .A2(n10573), .ZN(n8146) );
  AOI211_X1 U9451 ( .C1(n8272), .C2(n10002), .A(n8147), .B(n8146), .ZN(n8148)
         );
  OAI21_X1 U9452 ( .B1(n8274), .B2(n4941), .A(n8148), .ZN(P1_U3286) );
  XOR2_X1 U9453 ( .A(n8149), .B(n8150), .Z(n8158) );
  AOI22_X1 U9454 ( .A1(n8151), .A2(n9788), .B1(n9786), .B2(n9807), .ZN(n8157)
         );
  INV_X1 U9455 ( .A(n8152), .ZN(n8155) );
  NOR2_X1 U9456 ( .A1(n8745), .A2(n8153), .ZN(n8154) );
  AOI211_X1 U9457 ( .C1(n9787), .C2(n8286), .A(n8155), .B(n8154), .ZN(n8156)
         );
  OAI211_X1 U9458 ( .C1(n8158), .C2(n9778), .A(n8157), .B(n8156), .ZN(P1_U3213) );
  XNOR2_X1 U9459 ( .A(n8161), .B(n8160), .ZN(n8162) );
  XNOR2_X1 U9460 ( .A(n8159), .B(n8162), .ZN(n8169) );
  AOI22_X1 U9461 ( .A1(n9788), .A2(n8163), .B1(n9786), .B2(n9806), .ZN(n8165)
         );
  OAI211_X1 U9462 ( .C1(n8246), .C2(n9775), .A(n8165), .B(n8164), .ZN(n8166)
         );
  AOI21_X1 U9463 ( .B1(n8167), .B2(n9789), .A(n8166), .ZN(n8168) );
  OAI21_X1 U9464 ( .B1(n8169), .B2(n9778), .A(n8168), .ZN(P1_U3221) );
  INV_X1 U9465 ( .A(n8170), .ZN(n8211) );
  NAND2_X1 U9466 ( .A1(n10286), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n8171) );
  OAI211_X1 U9467 ( .C1(n8211), .C2(n10293), .A(n8172), .B(n8171), .ZN(
        P1_U3335) );
  NAND2_X1 U9468 ( .A1(n8174), .A2(n8173), .ZN(n8175) );
  XOR2_X1 U9469 ( .A(n8179), .B(n8175), .Z(n8177) );
  OAI22_X1 U9470 ( .A1(n8177), .A2(n10561), .B1(n8176), .B2(n10143), .ZN(
        n10643) );
  INV_X1 U9471 ( .A(n10643), .ZN(n8187) );
  OAI21_X1 U9472 ( .B1(n8180), .B2(n8179), .A(n8178), .ZN(n10645) );
  XNOR2_X1 U9473 ( .A(n8253), .B(n5757), .ZN(n8182) );
  NOR2_X1 U9474 ( .A1(n8290), .A2(n10145), .ZN(n8181) );
  AOI21_X1 U9475 ( .B1(n8182), .B2(n10552), .A(n8181), .ZN(n10642) );
  AOI22_X1 U9476 ( .A1(n4941), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n8287), .B2(
        n10572), .ZN(n8184) );
  NAND2_X1 U9477 ( .A1(n10570), .A2(n5757), .ZN(n8183) );
  OAI211_X1 U9478 ( .C1(n10642), .C2(n10608), .A(n8184), .B(n8183), .ZN(n8185)
         );
  AOI21_X1 U9479 ( .B1(n10645), .B2(n10615), .A(n8185), .ZN(n8186) );
  OAI21_X1 U9480 ( .B1(n8187), .B2(n4941), .A(n8186), .ZN(P1_U3284) );
  NAND2_X1 U9481 ( .A1(n8188), .A2(n8297), .ZN(n8190) );
  NAND2_X1 U9482 ( .A1(n8190), .A2(n8189), .ZN(n8191) );
  XNOR2_X1 U9483 ( .A(n8191), .B(n8891), .ZN(n8193) );
  OAI22_X1 U9484 ( .A1(n8193), .A2(n9498), .B1(n8192), .B2(n9515), .ZN(n8237)
         );
  XNOR2_X1 U9485 ( .A(n8194), .B(n8891), .ZN(n8235) );
  INV_X1 U9486 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n8197) );
  INV_X1 U9487 ( .A(n8195), .ZN(n8196) );
  OAI22_X1 U9488 ( .A1(n10641), .A2(n8197), .B1(n8196), .B2(n10677), .ZN(n8198) );
  AOI21_X1 U9489 ( .B1(n9470), .B2(n9283), .A(n8198), .ZN(n8200) );
  NAND2_X1 U9490 ( .A1(n8241), .A2(n10636), .ZN(n8199) );
  OAI211_X1 U9491 ( .C1(n8235), .C2(n9493), .A(n8200), .B(n8199), .ZN(n8201)
         );
  AOI21_X1 U9492 ( .B1(n8237), .B2(n10641), .A(n8201), .ZN(n8202) );
  INV_X1 U9493 ( .A(n8202), .ZN(P2_U3224) );
  AOI211_X1 U9494 ( .C1(n10667), .C2(n8205), .A(n8204), .B(n8203), .ZN(n8207)
         );
  MUX2_X1 U9495 ( .A(n7413), .B(n8207), .S(n10646), .Z(n8206) );
  OAI21_X1 U9496 ( .B1(n5744), .B2(n10219), .A(n8206), .ZN(P1_U3530) );
  INV_X1 U9497 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n8208) );
  MUX2_X1 U9498 ( .A(n8208), .B(n8207), .S(n10674), .Z(n8209) );
  OAI21_X1 U9499 ( .B1(n5744), .B2(n10267), .A(n8209), .ZN(P1_U3477) );
  OAI222_X1 U9500 ( .A1(n9676), .A2(n8211), .B1(n9137), .B2(n8210), .C1(n9070), 
        .C2(P2_U3151), .ZN(P2_U3275) );
  NAND2_X1 U9501 ( .A1(n8188), .A2(n8212), .ZN(n8214) );
  NAND2_X1 U9502 ( .A1(n8214), .A2(n8213), .ZN(n8215) );
  XOR2_X1 U9503 ( .A(n8888), .B(n8215), .Z(n8216) );
  OAI22_X1 U9504 ( .A1(n8216), .A2(n9498), .B1(n8267), .B2(n9515), .ZN(n8361)
         );
  INV_X1 U9505 ( .A(n8361), .ZN(n8222) );
  XNOR2_X1 U9506 ( .A(n8217), .B(n8888), .ZN(n8363) );
  NAND2_X1 U9507 ( .A1(n8359), .A2(n10636), .ZN(n8219) );
  AOI22_X1 U9508 ( .A1(n10687), .A2(P2_REG2_REG_10__SCAN_IN), .B1(n10634), 
        .B2(n8264), .ZN(n8218) );
  OAI211_X1 U9509 ( .C1(n8388), .C2(n9545), .A(n8219), .B(n8218), .ZN(n8220)
         );
  AOI21_X1 U9510 ( .B1(n8363), .B2(n9547), .A(n8220), .ZN(n8221) );
  OAI21_X1 U9511 ( .B1(n8222), .B2(n10687), .A(n8221), .ZN(P2_U3223) );
  AOI211_X1 U9512 ( .C1(n8225), .C2(n8224), .A(n8223), .B(n9894), .ZN(n8234)
         );
  AOI211_X1 U9513 ( .C1(n8228), .C2(n8227), .A(n8226), .B(n9926), .ZN(n8233)
         );
  INV_X1 U9514 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n8231) );
  NAND2_X1 U9515 ( .A1(n10528), .A2(n8229), .ZN(n8230) );
  NAND2_X1 U9516 ( .A1(P1_U3086), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n8820) );
  OAI211_X1 U9517 ( .C1(n8231), .C2(n9921), .A(n8230), .B(n8820), .ZN(n8232)
         );
  OR3_X1 U9518 ( .A1(n8234), .A2(n8233), .A3(n8232), .ZN(P1_U3257) );
  OAI22_X1 U9519 ( .A1(n8235), .A2(n9615), .B1(n8353), .B2(n9616), .ZN(n8236)
         );
  NOR2_X1 U9520 ( .A1(n8237), .A2(n8236), .ZN(n8243) );
  AOI22_X1 U9521 ( .A1(n8241), .A2(n8304), .B1(n9624), .B2(
        P2_REG1_REG_9__SCAN_IN), .ZN(n8238) );
  OAI21_X1 U9522 ( .B1(n8243), .B2(n9624), .A(n8238), .ZN(P2_U3468) );
  INV_X1 U9523 ( .A(n9654), .ZN(n8299) );
  INV_X1 U9524 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n8239) );
  NOR2_X1 U9525 ( .A1(n10695), .A2(n8239), .ZN(n8240) );
  AOI21_X1 U9526 ( .B1(n8241), .B2(n8299), .A(n8240), .ZN(n8242) );
  OAI21_X1 U9527 ( .B1(n8243), .B2(n10692), .A(n8242), .ZN(P2_U3417) );
  XNOR2_X1 U9528 ( .A(n8245), .B(n8244), .ZN(n8248) );
  OAI22_X1 U9529 ( .A1(n8706), .A2(n10145), .B1(n8246), .B2(n10143), .ZN(n8247) );
  AOI21_X1 U9530 ( .B1(n8248), .B2(n10127), .A(n8247), .ZN(n10652) );
  OAI21_X1 U9531 ( .B1(n8251), .B2(n8250), .A(n8249), .ZN(n10655) );
  NAND2_X1 U9532 ( .A1(n10655), .A2(n10615), .ZN(n8259) );
  OAI22_X1 U9533 ( .A1(n7834), .A2(n7393), .B1(n8252), .B2(n10606), .ZN(n8257)
         );
  INV_X1 U9534 ( .A(n8253), .ZN(n8254) );
  OAI21_X1 U9535 ( .B1(n8254), .B2(n5757), .A(n4944), .ZN(n8255) );
  NAND2_X1 U9536 ( .A1(n8255), .A2(n8329), .ZN(n10653) );
  INV_X1 U9537 ( .A(n10002), .ZN(n8668) );
  NOR2_X1 U9538 ( .A1(n10653), .A2(n8668), .ZN(n8256) );
  AOI211_X1 U9539 ( .C1(n10570), .C2(n4944), .A(n8257), .B(n8256), .ZN(n8258)
         );
  OAI211_X1 U9540 ( .C1(n4941), .C2(n10652), .A(n8259), .B(n8258), .ZN(
        P1_U3283) );
  INV_X1 U9541 ( .A(n8260), .ZN(n8261) );
  NAND2_X1 U9542 ( .A1(n8261), .A2(n9284), .ZN(n8262) );
  XOR2_X1 U9543 ( .A(n9115), .B(n8359), .Z(n8348) );
  XNOR2_X1 U9544 ( .A(n8349), .B(n8353), .ZN(n8270) );
  NAND2_X1 U9545 ( .A1(n9266), .A2(n8264), .ZN(n8266) );
  AOI22_X1 U9546 ( .A1(n9238), .A2(n9282), .B1(P2_REG3_REG_10__SCAN_IN), .B2(
        P2_U3151), .ZN(n8265) );
  OAI211_X1 U9547 ( .C1(n8267), .C2(n9240), .A(n8266), .B(n8265), .ZN(n8268)
         );
  AOI21_X1 U9548 ( .B1(n8359), .B2(n9251), .A(n8268), .ZN(n8269) );
  OAI21_X1 U9549 ( .B1(n8270), .B2(n9254), .A(n8269), .ZN(P2_U3157) );
  AOI22_X1 U9550 ( .A1(n8272), .A2(n10552), .B1(n10649), .B2(n8271), .ZN(n8273) );
  OAI211_X1 U9551 ( .C1(n8275), .C2(n10539), .A(n8274), .B(n8273), .ZN(n8277)
         );
  NAND2_X1 U9552 ( .A1(n8277), .A2(n10646), .ZN(n8276) );
  OAI21_X1 U9553 ( .B1(n10646), .B2(n7412), .A(n8276), .ZN(P1_U3529) );
  INV_X1 U9554 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n8279) );
  NAND2_X1 U9555 ( .A1(n8277), .A2(n10674), .ZN(n8278) );
  OAI21_X1 U9556 ( .B1(n10674), .B2(n8279), .A(n8278), .ZN(P1_U3474) );
  NAND2_X1 U9557 ( .A1(n9825), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n8280) );
  OAI21_X1 U9558 ( .B1(n8281), .B2(n9825), .A(n8280), .ZN(P1_U3583) );
  XNOR2_X1 U9559 ( .A(n8284), .B(n8283), .ZN(n8285) );
  XNOR2_X1 U9560 ( .A(n8282), .B(n8285), .ZN(n8293) );
  AOI22_X1 U9561 ( .A1(n8287), .A2(n9788), .B1(n9786), .B2(n8286), .ZN(n8289)
         );
  OAI211_X1 U9562 ( .C1(n8290), .C2(n9775), .A(n8289), .B(n8288), .ZN(n8291)
         );
  AOI21_X1 U9563 ( .B1(n5757), .B2(n9789), .A(n8291), .ZN(n8292) );
  OAI21_X1 U9564 ( .B1(n8293), .B2(n9778), .A(n8292), .ZN(P1_U3231) );
  INV_X1 U9565 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n8302) );
  NAND2_X1 U9566 ( .A1(n8295), .A2(n8294), .ZN(n8296) );
  XNOR2_X1 U9567 ( .A(n8296), .B(n8886), .ZN(n10632) );
  XNOR2_X1 U9568 ( .A(n8188), .B(n8297), .ZN(n8298) );
  AOI222_X1 U9569 ( .A1(n9532), .A2(n8298), .B1(n9284), .B2(n9609), .C1(n9286), 
        .C2(n9534), .ZN(n10631) );
  OAI21_X1 U9570 ( .B1(n9615), .B2(n10632), .A(n10631), .ZN(n8303) );
  NAND2_X1 U9571 ( .A1(n8303), .A2(n10695), .ZN(n8301) );
  NAND2_X1 U9572 ( .A1(n8299), .A2(n10637), .ZN(n8300) );
  OAI211_X1 U9573 ( .C1(n10695), .C2(n8302), .A(n8301), .B(n8300), .ZN(
        P2_U3414) );
  NAND2_X1 U9574 ( .A1(n8303), .A2(n9627), .ZN(n8306) );
  NAND2_X1 U9575 ( .A1(n10637), .A2(n8304), .ZN(n8305) );
  OAI211_X1 U9576 ( .C1(n9627), .C2(n5092), .A(n8306), .B(n8305), .ZN(P2_U3467) );
  INV_X1 U9577 ( .A(n8307), .ZN(n8318) );
  INV_X1 U9578 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n8308) );
  OAI222_X1 U9579 ( .A1(n9676), .A2(n8318), .B1(P2_U3151), .B2(n8927), .C1(
        n8308), .C2(n9137), .ZN(P2_U3274) );
  XNOR2_X1 U9580 ( .A(n8309), .B(n8890), .ZN(n8310) );
  OAI22_X1 U9581 ( .A1(n8310), .A2(n9498), .B1(n8353), .B2(n9515), .ZN(n8398)
         );
  INV_X1 U9582 ( .A(n8398), .ZN(n8317) );
  OAI21_X1 U9583 ( .B1(n8312), .B2(n8890), .A(n8311), .ZN(n8400) );
  NAND2_X1 U9584 ( .A1(n8397), .A2(n10636), .ZN(n8314) );
  AOI22_X1 U9585 ( .A1(n10687), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n10634), 
        .B2(n8350), .ZN(n8313) );
  OAI211_X1 U9586 ( .C1(n8698), .C2(n9545), .A(n8314), .B(n8313), .ZN(n8315)
         );
  AOI21_X1 U9587 ( .B1(n8400), .B2(n9547), .A(n8315), .ZN(n8316) );
  OAI21_X1 U9588 ( .B1(n8317), .B2(n10687), .A(n8316), .ZN(P2_U3222) );
  OAI222_X1 U9589 ( .A1(n8320), .A2(P1_U3086), .B1(n10290), .B2(n8319), .C1(
        n8318), .C2(n10293), .ZN(P1_U3334) );
  OAI21_X1 U9590 ( .B1(n8322), .B2(n8323), .A(n8321), .ZN(n8653) );
  INV_X1 U9591 ( .A(n8653), .ZN(n8334) );
  NAND2_X1 U9592 ( .A1(n8324), .A2(n8323), .ZN(n8325) );
  NAND3_X1 U9593 ( .A1(n8326), .A2(n10127), .A3(n8325), .ZN(n8328) );
  AOI22_X1 U9594 ( .A1(n9805), .A2(n10557), .B1(n10558), .B2(n9803), .ZN(n8327) );
  NAND2_X1 U9595 ( .A1(n8328), .A2(n8327), .ZN(n8651) );
  AOI211_X1 U9596 ( .C1(n8771), .C2(n8329), .A(n10663), .B(n5023), .ZN(n8652)
         );
  NAND2_X1 U9597 ( .A1(n8652), .A2(n10576), .ZN(n8331) );
  AOI22_X1 U9598 ( .A1(n10619), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n8760), .B2(
        n10572), .ZN(n8330) );
  OAI211_X1 U9599 ( .C1(n5192), .C2(n10612), .A(n8331), .B(n8330), .ZN(n8332)
         );
  AOI21_X1 U9600 ( .B1(n7834), .B2(n8651), .A(n8332), .ZN(n8333) );
  OAI21_X1 U9601 ( .B1(n8334), .B2(n10154), .A(n8333), .ZN(P1_U3282) );
  XOR2_X1 U9602 ( .A(n8336), .B(n8335), .Z(n8337) );
  XNOR2_X1 U9603 ( .A(n8338), .B(n8337), .ZN(n8344) );
  AOI22_X1 U9604 ( .A1(n8339), .A2(n9788), .B1(n9786), .B2(n5343), .ZN(n8341)
         );
  OAI211_X1 U9605 ( .C1(n8706), .C2(n9775), .A(n8341), .B(n8340), .ZN(n8342)
         );
  AOI21_X1 U9606 ( .B1(n4944), .B2(n9789), .A(n8342), .ZN(n8343) );
  OAI21_X1 U9607 ( .B1(n8344), .B2(n9778), .A(n8343), .ZN(P1_U3217) );
  INV_X1 U9608 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n8345) );
  OAI222_X1 U9609 ( .A1(n9676), .A2(n8357), .B1(P2_U3151), .B2(n8346), .C1(
        n8345), .C2(n9137), .ZN(P2_U3273) );
  OAI22_X1 U9610 ( .A1(n8349), .A2(n9283), .B1(n8348), .B2(n8347), .ZN(n8369)
         );
  XNOR2_X1 U9611 ( .A(n8397), .B(n9115), .ZN(n8366) );
  XNOR2_X1 U9612 ( .A(n8366), .B(n9282), .ZN(n8368) );
  XOR2_X1 U9613 ( .A(n8369), .B(n8368), .Z(n8356) );
  AOI22_X1 U9614 ( .A1(n9281), .A2(n9238), .B1(P2_REG3_REG_11__SCAN_IN), .B2(
        P2_U3151), .ZN(n8352) );
  NAND2_X1 U9615 ( .A1(n9266), .A2(n8350), .ZN(n8351) );
  OAI211_X1 U9616 ( .C1(n8353), .C2(n9240), .A(n8352), .B(n8351), .ZN(n8354)
         );
  AOI21_X1 U9617 ( .B1(n8397), .B2(n9251), .A(n8354), .ZN(n8355) );
  OAI21_X1 U9618 ( .B1(n8356), .B2(n9254), .A(n8355), .ZN(P2_U3176) );
  INV_X1 U9619 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n8358) );
  OAI222_X1 U9620 ( .A1(n10290), .A2(n8358), .B1(P1_U3086), .B2(n6065), .C1(
        n8357), .C2(n10293), .ZN(P1_U3333) );
  INV_X1 U9621 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n8365) );
  INV_X1 U9622 ( .A(n8359), .ZN(n8360) );
  OAI22_X1 U9623 ( .A1(n8360), .A2(n9618), .B1(n8388), .B2(n9616), .ZN(n8362)
         );
  AOI211_X1 U9624 ( .C1(n9623), .C2(n8363), .A(n8362), .B(n8361), .ZN(n10659)
         );
  OR2_X1 U9625 ( .A1(n10659), .A2(n9624), .ZN(n8364) );
  OAI21_X1 U9626 ( .B1(n9627), .B2(n8365), .A(n8364), .ZN(P2_U3469) );
  MUX2_X1 U9627 ( .A(n8370), .B(n8971), .S(n9115), .Z(n8643) );
  INV_X1 U9628 ( .A(n8643), .ZN(n8371) );
  MUX2_X1 U9629 ( .A(n8384), .B(n8973), .S(n9115), .Z(n8644) );
  NOR2_X1 U9630 ( .A1(n8371), .A2(n8644), .ZN(n8372) );
  XNOR2_X1 U9631 ( .A(n8645), .B(n8372), .ZN(n8377) );
  INV_X1 U9632 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n8594) );
  NOR2_X1 U9633 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8594), .ZN(n8631) );
  AOI21_X1 U9634 ( .B1(n9261), .B2(n9282), .A(n8631), .ZN(n8374) );
  NAND2_X1 U9635 ( .A1(n9266), .A2(n8389), .ZN(n8373) );
  OAI211_X1 U9636 ( .C1(n8718), .C2(n9263), .A(n8374), .B(n8373), .ZN(n8375)
         );
  AOI21_X1 U9637 ( .B1(n8715), .B2(n9251), .A(n8375), .ZN(n8376) );
  OAI21_X1 U9638 ( .B1(n8377), .B2(n9254), .A(n8376), .ZN(P2_U3164) );
  INV_X1 U9639 ( .A(n8378), .ZN(n8383) );
  NAND2_X1 U9640 ( .A1(n8379), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9080) );
  NAND2_X1 U9641 ( .A1(n9674), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n8380) );
  OAI211_X1 U9642 ( .C1(n8383), .C2(n9676), .A(n9080), .B(n8380), .ZN(P2_U3272) );
  NAND2_X1 U9643 ( .A1(n10286), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n8382) );
  OAI211_X1 U9644 ( .C1(n8383), .C2(n10293), .A(n8382), .B(n8381), .ZN(
        P1_U3332) );
  XNOR2_X1 U9645 ( .A(n8386), .B(n8976), .ZN(n8387) );
  OAI222_X1 U9646 ( .A1(n9515), .A2(n8388), .B1(n9616), .B2(n8718), .C1(n8387), 
        .C2(n9498), .ZN(n8713) );
  AOI21_X1 U9647 ( .B1(n10634), .B2(n8389), .A(n8713), .ZN(n8396) );
  XOR2_X1 U9648 ( .A(n8390), .B(n8976), .Z(n8712) );
  INV_X1 U9649 ( .A(n8712), .ZN(n8394) );
  INV_X1 U9650 ( .A(n8715), .ZN(n8392) );
  OAI22_X1 U9651 ( .A1(n8392), .A2(n9509), .B1(n8391), .B2(n10641), .ZN(n8393)
         );
  AOI21_X1 U9652 ( .B1(n8394), .B2(n9547), .A(n8393), .ZN(n8395) );
  OAI21_X1 U9653 ( .B1(n8396), .B2(n10687), .A(n8395), .ZN(P2_U3221) );
  INV_X1 U9654 ( .A(n8397), .ZN(n8405) );
  INV_X1 U9655 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n8401) );
  NOR2_X1 U9656 ( .A1(n8698), .A2(n9616), .ZN(n8399) );
  AOI211_X1 U9657 ( .C1(n9623), .C2(n8400), .A(n8399), .B(n8398), .ZN(n8403)
         );
  MUX2_X1 U9658 ( .A(n8401), .B(n8403), .S(n10695), .Z(n8402) );
  OAI21_X1 U9659 ( .B1(n8405), .B2(n9654), .A(n8402), .ZN(P2_U3423) );
  MUX2_X1 U9660 ( .A(n10508), .B(n8403), .S(n9627), .Z(n8404) );
  OAI21_X1 U9661 ( .B1(n8405), .B2(n9594), .A(n8404), .ZN(P2_U3470) );
  INV_X1 U9662 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n9260) );
  OAI22_X1 U9663 ( .A1(n9260), .A2(keyinput_63), .B1(keyinput_62), .B2(
        P2_REG3_REG_26__SCAN_IN), .ZN(n8406) );
  AOI221_X1 U9664 ( .B1(n9260), .B2(keyinput_63), .C1(P2_REG3_REG_26__SCAN_IN), 
        .C2(keyinput_62), .A(n8406), .ZN(n8503) );
  INV_X1 U9665 ( .A(keyinput_60), .ZN(n8501) );
  INV_X1 U9666 ( .A(keyinput_59), .ZN(n8499) );
  OAI22_X1 U9667 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(keyinput_48), .B1(
        keyinput_49), .B2(P2_REG3_REG_5__SCAN_IN), .ZN(n8407) );
  AOI221_X1 U9668 ( .B1(P2_REG3_REG_16__SCAN_IN), .B2(keyinput_48), .C1(
        P2_REG3_REG_5__SCAN_IN), .C2(keyinput_49), .A(n8407), .ZN(n8487) );
  INV_X1 U9669 ( .A(keyinput_47), .ZN(n8483) );
  INV_X1 U9670 ( .A(keyinput_46), .ZN(n8481) );
  INV_X1 U9671 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n8591) );
  INV_X1 U9672 ( .A(keyinput_45), .ZN(n8479) );
  OAI22_X1 U9673 ( .A1(P2_REG3_REG_23__SCAN_IN), .A2(keyinput_38), .B1(
        P2_REG3_REG_10__SCAN_IN), .B2(keyinput_39), .ZN(n8408) );
  AOI221_X1 U9674 ( .B1(P2_REG3_REG_23__SCAN_IN), .B2(keyinput_38), .C1(
        keyinput_39), .C2(P2_REG3_REG_10__SCAN_IN), .A(n8408), .ZN(n8470) );
  INV_X1 U9675 ( .A(keyinput_37), .ZN(n8468) );
  INV_X1 U9676 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n8576) );
  INV_X1 U9677 ( .A(keyinput_36), .ZN(n8466) );
  INV_X1 U9678 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n8573) );
  INV_X1 U9679 ( .A(keyinput_35), .ZN(n8464) );
  INV_X1 U9680 ( .A(keyinput_34), .ZN(n8462) );
  INV_X1 U9681 ( .A(keyinput_19), .ZN(n8439) );
  INV_X1 U9682 ( .A(SI_14_), .ZN(n8541) );
  INV_X1 U9683 ( .A(keyinput_18), .ZN(n8437) );
  OAI22_X1 U9684 ( .A1(SI_20_), .A2(keyinput_12), .B1(keyinput_13), .B2(SI_19_), .ZN(n8409) );
  AOI221_X1 U9685 ( .B1(SI_20_), .B2(keyinput_12), .C1(SI_19_), .C2(
        keyinput_13), .A(n8409), .ZN(n8429) );
  INV_X1 U9686 ( .A(SI_25_), .ZN(n8412) );
  AOI22_X1 U9687 ( .A1(n8412), .A2(keyinput_7), .B1(n8411), .B2(keyinput_6), 
        .ZN(n8410) );
  OAI221_X1 U9688 ( .B1(n8412), .B2(keyinput_7), .C1(n8411), .C2(keyinput_6), 
        .A(n8410), .ZN(n8422) );
  INV_X1 U9689 ( .A(keyinput_5), .ZN(n8420) );
  OAI22_X1 U9690 ( .A1(SI_31_), .A2(keyinput_1), .B1(keyinput_0), .B2(
        P2_WR_REG_SCAN_IN), .ZN(n8413) );
  AOI221_X1 U9691 ( .B1(SI_31_), .B2(keyinput_1), .C1(P2_WR_REG_SCAN_IN), .C2(
        keyinput_0), .A(n8413), .ZN(n8417) );
  OAI22_X1 U9692 ( .A1(n8517), .A2(keyinput_2), .B1(keyinput_3), .B2(SI_29_), 
        .ZN(n8414) );
  AOI221_X1 U9693 ( .B1(n8517), .B2(keyinput_2), .C1(SI_29_), .C2(keyinput_3), 
        .A(n8414), .ZN(n8415) );
  OAI21_X1 U9694 ( .B1(n8418), .B2(keyinput_4), .A(n8415), .ZN(n8416) );
  AOI211_X1 U9695 ( .C1(n8418), .C2(keyinput_4), .A(n8417), .B(n8416), .ZN(
        n8419) );
  AOI221_X1 U9696 ( .B1(SI_27_), .B2(keyinput_5), .C1(n8523), .C2(n8420), .A(
        n8419), .ZN(n8421) );
  OAI22_X1 U9697 ( .A1(n8422), .A2(n8421), .B1(SI_24_), .B2(keyinput_8), .ZN(
        n8423) );
  AOI21_X1 U9698 ( .B1(SI_24_), .B2(keyinput_8), .A(n8423), .ZN(n8426) );
  OAI22_X1 U9699 ( .A1(n8527), .A2(keyinput_10), .B1(keyinput_9), .B2(SI_23_), 
        .ZN(n8424) );
  AOI221_X1 U9700 ( .B1(n8527), .B2(keyinput_10), .C1(SI_23_), .C2(keyinput_9), 
        .A(n8424), .ZN(n8425) );
  AOI22_X1 U9701 ( .A1(n8426), .A2(n8425), .B1(keyinput_11), .B2(SI_21_), .ZN(
        n8427) );
  OAI21_X1 U9702 ( .B1(keyinput_11), .B2(SI_21_), .A(n8427), .ZN(n8428) );
  AOI22_X1 U9703 ( .A1(n8429), .A2(n8428), .B1(SI_17_), .B2(keyinput_15), .ZN(
        n8430) );
  OAI21_X1 U9704 ( .B1(SI_17_), .B2(keyinput_15), .A(n8430), .ZN(n8435) );
  AOI22_X1 U9705 ( .A1(n8535), .A2(keyinput_16), .B1(n8432), .B2(keyinput_14), 
        .ZN(n8431) );
  OAI221_X1 U9706 ( .B1(n8535), .B2(keyinput_16), .C1(n8432), .C2(keyinput_14), 
        .A(n8431), .ZN(n8434) );
  NAND2_X1 U9707 ( .A1(SI_15_), .A2(keyinput_17), .ZN(n8433) );
  OAI221_X1 U9708 ( .B1(n8435), .B2(n8434), .C1(SI_15_), .C2(keyinput_17), .A(
        n8433), .ZN(n8436) );
  OAI221_X1 U9709 ( .B1(SI_14_), .B2(keyinput_18), .C1(n8541), .C2(n8437), .A(
        n8436), .ZN(n8438) );
  OAI221_X1 U9710 ( .B1(SI_13_), .B2(n8439), .C1(n8544), .C2(keyinput_19), .A(
        n8438), .ZN(n8454) );
  AOI22_X1 U9711 ( .A1(SI_7_), .A2(keyinput_25), .B1(SI_10_), .B2(keyinput_22), 
        .ZN(n8440) );
  OAI221_X1 U9712 ( .B1(SI_7_), .B2(keyinput_25), .C1(SI_10_), .C2(keyinput_22), .A(n8440), .ZN(n8446) );
  AOI22_X1 U9713 ( .A1(n5426), .A2(keyinput_21), .B1(keyinput_23), .B2(n8549), 
        .ZN(n8441) );
  OAI221_X1 U9714 ( .B1(n5426), .B2(keyinput_21), .C1(n8549), .C2(keyinput_23), 
        .A(n8441), .ZN(n8445) );
  XOR2_X1 U9715 ( .A(n8556), .B(keyinput_26), .Z(n8444) );
  AOI22_X1 U9716 ( .A1(SI_12_), .A2(keyinput_20), .B1(n8557), .B2(keyinput_24), 
        .ZN(n8442) );
  OAI221_X1 U9717 ( .B1(SI_12_), .B2(keyinput_20), .C1(n8557), .C2(keyinput_24), .A(n8442), .ZN(n8443) );
  NOR4_X1 U9718 ( .A1(n8446), .A2(n8445), .A3(n8444), .A4(n8443), .ZN(n8453)
         );
  AOI22_X1 U9719 ( .A1(SI_5_), .A2(keyinput_27), .B1(n8448), .B2(keyinput_28), 
        .ZN(n8447) );
  OAI221_X1 U9720 ( .B1(SI_5_), .B2(keyinput_27), .C1(n8448), .C2(keyinput_28), 
        .A(n8447), .ZN(n8452) );
  XNOR2_X1 U9721 ( .A(SI_3_), .B(keyinput_29), .ZN(n8450) );
  XNOR2_X1 U9722 ( .A(SI_2_), .B(keyinput_30), .ZN(n8449) );
  NAND2_X1 U9723 ( .A1(n8450), .A2(n8449), .ZN(n8451) );
  AOI211_X1 U9724 ( .C1(n8454), .C2(n8453), .A(n8452), .B(n8451), .ZN(n8459)
         );
  AND2_X1 U9725 ( .A1(SI_0_), .A2(keyinput_32), .ZN(n8458) );
  XNOR2_X1 U9726 ( .A(n8455), .B(keyinput_31), .ZN(n8457) );
  INV_X1 U9727 ( .A(P2_RD_REG_SCAN_IN), .ZN(n10516) );
  XNOR2_X1 U9728 ( .A(keyinput_33), .B(n10516), .ZN(n8456) );
  NOR4_X1 U9729 ( .A1(n8459), .A2(n8458), .A3(n8457), .A4(n8456), .ZN(n8460)
         );
  OAI21_X1 U9730 ( .B1(SI_0_), .B2(keyinput_32), .A(n8460), .ZN(n8461) );
  OAI221_X1 U9731 ( .B1(P2_STATE_REG_SCAN_IN), .B2(keyinput_34), .C1(P2_U3151), 
        .C2(n8462), .A(n8461), .ZN(n8463) );
  OAI221_X1 U9732 ( .B1(P2_REG3_REG_7__SCAN_IN), .B2(keyinput_35), .C1(n8573), 
        .C2(n8464), .A(n8463), .ZN(n8465) );
  OAI221_X1 U9733 ( .B1(P2_REG3_REG_27__SCAN_IN), .B2(keyinput_36), .C1(n8576), 
        .C2(n8466), .A(n8465), .ZN(n8467) );
  OAI221_X1 U9734 ( .B1(P2_REG3_REG_14__SCAN_IN), .B2(n8468), .C1(n8723), .C2(
        keyinput_37), .A(n8467), .ZN(n8469) );
  OAI211_X1 U9735 ( .C1(P2_REG3_REG_3__SCAN_IN), .C2(keyinput_40), .A(n8470), 
        .B(n8469), .ZN(n8471) );
  AOI21_X1 U9736 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(keyinput_40), .A(n8471), 
        .ZN(n8477) );
  INV_X1 U9737 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n8473) );
  AOI22_X1 U9738 ( .A1(n8473), .A2(keyinput_41), .B1(n6819), .B2(keyinput_42), 
        .ZN(n8472) );
  OAI221_X1 U9739 ( .B1(n8473), .B2(keyinput_41), .C1(n6819), .C2(keyinput_42), 
        .A(n8472), .ZN(n8476) );
  OAI22_X1 U9740 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(keyinput_43), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(keyinput_44), .ZN(n8474) );
  AOI221_X1 U9741 ( .B1(P2_REG3_REG_8__SCAN_IN), .B2(keyinput_43), .C1(
        keyinput_44), .C2(P2_REG3_REG_1__SCAN_IN), .A(n8474), .ZN(n8475) );
  OAI21_X1 U9742 ( .B1(n8477), .B2(n8476), .A(n8475), .ZN(n8478) );
  OAI221_X1 U9743 ( .B1(P2_REG3_REG_21__SCAN_IN), .B2(keyinput_45), .C1(n8591), 
        .C2(n8479), .A(n8478), .ZN(n8480) );
  OAI221_X1 U9744 ( .B1(P2_REG3_REG_12__SCAN_IN), .B2(n8481), .C1(n8594), .C2(
        keyinput_46), .A(n8480), .ZN(n8482) );
  OAI221_X1 U9745 ( .B1(P2_REG3_REG_25__SCAN_IN), .B2(keyinput_47), .C1(n8596), 
        .C2(n8483), .A(n8482), .ZN(n8486) );
  INV_X1 U9746 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n9204) );
  AOI22_X1 U9747 ( .A1(P2_REG3_REG_24__SCAN_IN), .A2(keyinput_51), .B1(n9204), 
        .B2(keyinput_50), .ZN(n8484) );
  OAI221_X1 U9748 ( .B1(P2_REG3_REG_24__SCAN_IN), .B2(keyinput_51), .C1(n9204), 
        .C2(keyinput_50), .A(n8484), .ZN(n8485) );
  AOI21_X1 U9749 ( .B1(n8487), .B2(n8486), .A(n8485), .ZN(n8491) );
  OAI22_X1 U9750 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(keyinput_52), .B1(
        keyinput_54), .B2(P2_REG3_REG_0__SCAN_IN), .ZN(n8488) );
  AOI221_X1 U9751 ( .B1(P2_REG3_REG_4__SCAN_IN), .B2(keyinput_52), .C1(
        P2_REG3_REG_0__SCAN_IN), .C2(keyinput_54), .A(n8488), .ZN(n8489) );
  OAI21_X1 U9752 ( .B1(keyinput_53), .B2(P2_REG3_REG_9__SCAN_IN), .A(n8489), 
        .ZN(n8490) );
  AOI211_X1 U9753 ( .C1(keyinput_53), .C2(P2_REG3_REG_9__SCAN_IN), .A(n8491), 
        .B(n8490), .ZN(n8497) );
  AOI22_X1 U9754 ( .A1(n6455), .A2(keyinput_56), .B1(n8493), .B2(keyinput_55), 
        .ZN(n8492) );
  OAI221_X1 U9755 ( .B1(n6455), .B2(keyinput_56), .C1(n8493), .C2(keyinput_55), 
        .A(n8492), .ZN(n8496) );
  OAI22_X1 U9756 ( .A1(n6461), .A2(keyinput_57), .B1(keyinput_58), .B2(
        P2_REG3_REG_11__SCAN_IN), .ZN(n8494) );
  AOI221_X1 U9757 ( .B1(n6461), .B2(keyinput_57), .C1(P2_REG3_REG_11__SCAN_IN), 
        .C2(keyinput_58), .A(n8494), .ZN(n8495) );
  OAI21_X1 U9758 ( .B1(n8497), .B2(n8496), .A(n8495), .ZN(n8498) );
  OAI221_X1 U9759 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(keyinput_59), .C1(n10584), 
        .C2(n8499), .A(n8498), .ZN(n8500) );
  OAI221_X1 U9760 ( .B1(P2_REG3_REG_18__SCAN_IN), .B2(n8501), .C1(n9237), .C2(
        keyinput_60), .A(n8500), .ZN(n8502) );
  OAI211_X1 U9761 ( .C1(P2_REG3_REG_6__SCAN_IN), .C2(keyinput_61), .A(n8503), 
        .B(n8502), .ZN(n8504) );
  AOI21_X1 U9762 ( .B1(P2_REG3_REG_6__SCAN_IN), .B2(keyinput_61), .A(n8504), 
        .ZN(n8620) );
  INV_X1 U9763 ( .A(keyinput_124), .ZN(n8614) );
  INV_X1 U9764 ( .A(keyinput_123), .ZN(n8612) );
  OAI22_X1 U9765 ( .A1(P2_REG3_REG_20__SCAN_IN), .A2(keyinput_119), .B1(
        keyinput_120), .B2(P2_REG3_REG_13__SCAN_IN), .ZN(n8505) );
  AOI221_X1 U9766 ( .B1(P2_REG3_REG_20__SCAN_IN), .B2(keyinput_119), .C1(
        P2_REG3_REG_13__SCAN_IN), .C2(keyinput_120), .A(n8505), .ZN(n8610) );
  OAI22_X1 U9767 ( .A1(n6450), .A2(keyinput_113), .B1(keyinput_112), .B2(
        P2_REG3_REG_16__SCAN_IN), .ZN(n8506) );
  AOI221_X1 U9768 ( .B1(n6450), .B2(keyinput_113), .C1(P2_REG3_REG_16__SCAN_IN), .C2(keyinput_112), .A(n8506), .ZN(n8601) );
  INV_X1 U9769 ( .A(keyinput_111), .ZN(n8597) );
  INV_X1 U9770 ( .A(keyinput_110), .ZN(n8593) );
  INV_X1 U9771 ( .A(keyinput_109), .ZN(n8590) );
  INV_X1 U9772 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n8583) );
  INV_X1 U9773 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n8508) );
  OAI22_X1 U9774 ( .A1(n8508), .A2(keyinput_102), .B1(keyinput_104), .B2(
        P2_REG3_REG_3__SCAN_IN), .ZN(n8507) );
  AOI221_X1 U9775 ( .B1(n8508), .B2(keyinput_102), .C1(P2_REG3_REG_3__SCAN_IN), 
        .C2(keyinput_104), .A(n8507), .ZN(n8581) );
  INV_X1 U9776 ( .A(keyinput_101), .ZN(n8579) );
  INV_X1 U9777 ( .A(keyinput_100), .ZN(n8577) );
  INV_X1 U9778 ( .A(keyinput_99), .ZN(n8574) );
  INV_X1 U9779 ( .A(keyinput_98), .ZN(n8571) );
  INV_X1 U9780 ( .A(keyinput_83), .ZN(n8545) );
  INV_X1 U9781 ( .A(keyinput_82), .ZN(n8542) );
  OAI22_X1 U9782 ( .A1(SI_18_), .A2(keyinput_78), .B1(keyinput_79), .B2(SI_17_), .ZN(n8509) );
  AOI221_X1 U9783 ( .B1(SI_18_), .B2(keyinput_78), .C1(SI_17_), .C2(
        keyinput_79), .A(n8509), .ZN(n8539) );
  AOI22_X1 U9784 ( .A1(n8512), .A2(keyinput_76), .B1(keyinput_77), .B2(n8511), 
        .ZN(n8510) );
  OAI221_X1 U9785 ( .B1(n8512), .B2(keyinput_76), .C1(n8511), .C2(keyinput_77), 
        .A(n8510), .ZN(n8533) );
  AOI22_X1 U9786 ( .A1(SI_23_), .A2(keyinput_73), .B1(SI_24_), .B2(keyinput_72), .ZN(n8513) );
  OAI221_X1 U9787 ( .B1(SI_23_), .B2(keyinput_73), .C1(SI_24_), .C2(
        keyinput_72), .A(n8513), .ZN(n8529) );
  OAI22_X1 U9788 ( .A1(SI_26_), .A2(keyinput_70), .B1(keyinput_71), .B2(SI_25_), .ZN(n8514) );
  AOI221_X1 U9789 ( .B1(SI_26_), .B2(keyinput_70), .C1(SI_25_), .C2(
        keyinput_71), .A(n8514), .ZN(n8525) );
  INV_X1 U9790 ( .A(keyinput_69), .ZN(n8522) );
  OAI22_X1 U9791 ( .A1(SI_31_), .A2(keyinput_65), .B1(keyinput_64), .B2(
        P2_WR_REG_SCAN_IN), .ZN(n8515) );
  AOI221_X1 U9792 ( .B1(SI_31_), .B2(keyinput_65), .C1(P2_WR_REG_SCAN_IN), 
        .C2(keyinput_64), .A(n8515), .ZN(n8519) );
  AOI22_X1 U9793 ( .A1(SI_29_), .A2(keyinput_67), .B1(n8517), .B2(keyinput_66), 
        .ZN(n8516) );
  OAI221_X1 U9794 ( .B1(SI_29_), .B2(keyinput_67), .C1(n8517), .C2(keyinput_66), .A(n8516), .ZN(n8518) );
  AOI211_X1 U9795 ( .C1(SI_28_), .C2(keyinput_68), .A(n8519), .B(n8518), .ZN(
        n8520) );
  OAI21_X1 U9796 ( .B1(SI_28_), .B2(keyinput_68), .A(n8520), .ZN(n8521) );
  OAI221_X1 U9797 ( .B1(SI_27_), .B2(keyinput_69), .C1(n8523), .C2(n8522), .A(
        n8521), .ZN(n8524) );
  AOI22_X1 U9798 ( .A1(n8525), .A2(n8524), .B1(keyinput_74), .B2(n8527), .ZN(
        n8526) );
  OAI21_X1 U9799 ( .B1(keyinput_74), .B2(n8527), .A(n8526), .ZN(n8528) );
  OAI22_X1 U9800 ( .A1(keyinput_75), .A2(n8531), .B1(n8529), .B2(n8528), .ZN(
        n8530) );
  AOI21_X1 U9801 ( .B1(keyinput_75), .B2(n8531), .A(n8530), .ZN(n8532) );
  OAI22_X1 U9802 ( .A1(n8533), .A2(n8532), .B1(n8535), .B2(keyinput_80), .ZN(
        n8534) );
  AOI21_X1 U9803 ( .B1(n8535), .B2(keyinput_80), .A(n8534), .ZN(n8538) );
  INV_X1 U9804 ( .A(SI_15_), .ZN(n8537) );
  NOR2_X1 U9805 ( .A1(n8537), .A2(keyinput_81), .ZN(n8536) );
  AOI221_X1 U9806 ( .B1(n8539), .B2(n8538), .C1(keyinput_81), .C2(n8537), .A(
        n8536), .ZN(n8540) );
  AOI221_X1 U9807 ( .B1(SI_14_), .B2(n8542), .C1(n8541), .C2(keyinput_82), .A(
        n8540), .ZN(n8543) );
  AOI221_X1 U9808 ( .B1(SI_13_), .B2(n8545), .C1(n8544), .C2(keyinput_83), .A(
        n8543), .ZN(n8554) );
  AOI22_X1 U9809 ( .A1(n8548), .A2(keyinput_89), .B1(n8547), .B2(keyinput_86), 
        .ZN(n8546) );
  OAI221_X1 U9810 ( .B1(n8548), .B2(keyinput_89), .C1(n8547), .C2(keyinput_86), 
        .A(n8546), .ZN(n8553) );
  XOR2_X1 U9811 ( .A(n8549), .B(keyinput_87), .Z(n8552) );
  AOI22_X1 U9812 ( .A1(SI_12_), .A2(keyinput_84), .B1(n5426), .B2(keyinput_85), 
        .ZN(n8550) );
  OAI221_X1 U9813 ( .B1(SI_12_), .B2(keyinput_84), .C1(n5426), .C2(keyinput_85), .A(n8550), .ZN(n8551) );
  NOR4_X1 U9814 ( .A1(n8554), .A2(n8553), .A3(n8552), .A4(n8551), .ZN(n8564)
         );
  OAI22_X1 U9815 ( .A1(n8557), .A2(keyinput_88), .B1(n8556), .B2(keyinput_90), 
        .ZN(n8555) );
  AOI221_X1 U9816 ( .B1(n8557), .B2(keyinput_88), .C1(keyinput_90), .C2(n8556), 
        .A(n8555), .ZN(n8563) );
  AOI22_X1 U9817 ( .A1(SI_3_), .A2(keyinput_93), .B1(SI_4_), .B2(keyinput_92), 
        .ZN(n8558) );
  OAI221_X1 U9818 ( .B1(SI_3_), .B2(keyinput_93), .C1(SI_4_), .C2(keyinput_92), 
        .A(n8558), .ZN(n8562) );
  XNOR2_X1 U9819 ( .A(SI_5_), .B(keyinput_91), .ZN(n8560) );
  XNOR2_X1 U9820 ( .A(SI_2_), .B(keyinput_94), .ZN(n8559) );
  NAND2_X1 U9821 ( .A1(n8560), .A2(n8559), .ZN(n8561) );
  AOI211_X1 U9822 ( .C1(n8564), .C2(n8563), .A(n8562), .B(n8561), .ZN(n8568)
         );
  INV_X1 U9823 ( .A(SI_0_), .ZN(n8566) );
  AOI22_X1 U9824 ( .A1(n10516), .A2(keyinput_97), .B1(keyinput_96), .B2(n8566), 
        .ZN(n8565) );
  OAI221_X1 U9825 ( .B1(n10516), .B2(keyinput_97), .C1(n8566), .C2(keyinput_96), .A(n8565), .ZN(n8567) );
  AOI211_X1 U9826 ( .C1(SI_1_), .C2(keyinput_95), .A(n8568), .B(n8567), .ZN(
        n8569) );
  OAI21_X1 U9827 ( .B1(SI_1_), .B2(keyinput_95), .A(n8569), .ZN(n8570) );
  OAI221_X1 U9828 ( .B1(P2_STATE_REG_SCAN_IN), .B2(keyinput_98), .C1(P2_U3151), 
        .C2(n8571), .A(n8570), .ZN(n8572) );
  OAI221_X1 U9829 ( .B1(P2_REG3_REG_7__SCAN_IN), .B2(n8574), .C1(n8573), .C2(
        keyinput_99), .A(n8572), .ZN(n8575) );
  OAI221_X1 U9830 ( .B1(P2_REG3_REG_27__SCAN_IN), .B2(n8577), .C1(n8576), .C2(
        keyinput_100), .A(n8575), .ZN(n8578) );
  OAI221_X1 U9831 ( .B1(P2_REG3_REG_14__SCAN_IN), .B2(keyinput_101), .C1(n8723), .C2(n8579), .A(n8578), .ZN(n8580) );
  OAI211_X1 U9832 ( .C1(n8583), .C2(keyinput_103), .A(n8581), .B(n8580), .ZN(
        n8582) );
  AOI21_X1 U9833 ( .B1(n8583), .B2(keyinput_103), .A(n8582), .ZN(n8588) );
  AOI22_X1 U9834 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(keyinput_105), .B1(n6819), 
        .B2(keyinput_106), .ZN(n8584) );
  OAI221_X1 U9835 ( .B1(P2_REG3_REG_19__SCAN_IN), .B2(keyinput_105), .C1(n6819), .C2(keyinput_106), .A(n8584), .ZN(n8587) );
  OAI22_X1 U9836 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(keyinput_107), .B1(
        keyinput_108), .B2(P2_REG3_REG_1__SCAN_IN), .ZN(n8585) );
  AOI221_X1 U9837 ( .B1(P2_REG3_REG_8__SCAN_IN), .B2(keyinput_107), .C1(
        P2_REG3_REG_1__SCAN_IN), .C2(keyinput_108), .A(n8585), .ZN(n8586) );
  OAI21_X1 U9838 ( .B1(n8588), .B2(n8587), .A(n8586), .ZN(n8589) );
  OAI221_X1 U9839 ( .B1(P2_REG3_REG_21__SCAN_IN), .B2(keyinput_109), .C1(n8591), .C2(n8590), .A(n8589), .ZN(n8592) );
  OAI221_X1 U9840 ( .B1(P2_REG3_REG_12__SCAN_IN), .B2(keyinput_110), .C1(n8594), .C2(n8593), .A(n8592), .ZN(n8595) );
  OAI221_X1 U9841 ( .B1(P2_REG3_REG_25__SCAN_IN), .B2(n8597), .C1(n8596), .C2(
        keyinput_111), .A(n8595), .ZN(n8600) );
  AOI22_X1 U9842 ( .A1(P2_REG3_REG_24__SCAN_IN), .A2(keyinput_115), .B1(n9204), 
        .B2(keyinput_114), .ZN(n8598) );
  OAI221_X1 U9843 ( .B1(P2_REG3_REG_24__SCAN_IN), .B2(keyinput_115), .C1(n9204), .C2(keyinput_114), .A(n8598), .ZN(n8599) );
  AOI21_X1 U9844 ( .B1(n8601), .B2(n8600), .A(n8599), .ZN(n8605) );
  INV_X1 U9845 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n8603) );
  AOI22_X1 U9846 ( .A1(P2_REG3_REG_0__SCAN_IN), .A2(keyinput_118), .B1(n8603), 
        .B2(keyinput_117), .ZN(n8602) );
  OAI221_X1 U9847 ( .B1(P2_REG3_REG_0__SCAN_IN), .B2(keyinput_118), .C1(n8603), 
        .C2(keyinput_117), .A(n8602), .ZN(n8604) );
  AOI211_X1 U9848 ( .C1(P2_REG3_REG_4__SCAN_IN), .C2(keyinput_116), .A(n8605), 
        .B(n8604), .ZN(n8606) );
  OAI21_X1 U9849 ( .B1(P2_REG3_REG_4__SCAN_IN), .B2(keyinput_116), .A(n8606), 
        .ZN(n8609) );
  AOI22_X1 U9850 ( .A1(P2_REG3_REG_11__SCAN_IN), .A2(keyinput_122), .B1(n6461), 
        .B2(keyinput_121), .ZN(n8607) );
  OAI221_X1 U9851 ( .B1(P2_REG3_REG_11__SCAN_IN), .B2(keyinput_122), .C1(n6461), .C2(keyinput_121), .A(n8607), .ZN(n8608) );
  AOI21_X1 U9852 ( .B1(n8610), .B2(n8609), .A(n8608), .ZN(n8611) );
  AOI221_X1 U9853 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(keyinput_123), .C1(n10584), .C2(n8612), .A(n8611), .ZN(n8613) );
  AOI221_X1 U9854 ( .B1(P2_REG3_REG_18__SCAN_IN), .B2(keyinput_124), .C1(n9237), .C2(n8614), .A(n8613), .ZN(n8619) );
  XOR2_X1 U9855 ( .A(n8615), .B(keyinput_125), .Z(n8618) );
  AOI22_X1 U9856 ( .A1(n9260), .A2(keyinput_127), .B1(n6793), .B2(keyinput_126), .ZN(n8616) );
  OAI221_X1 U9857 ( .B1(n9260), .B2(keyinput_127), .C1(n6793), .C2(
        keyinput_126), .A(n8616), .ZN(n8617) );
  NOR4_X1 U9858 ( .A1(n8620), .A2(n8619), .A3(n8618), .A4(n8617), .ZN(n8625)
         );
  AOI222_X1 U9859 ( .A1(n8623), .A2(n8622), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8621), .C1(P2_DATAO_REG_9__SCAN_IN), .C2(n10286), .ZN(n8624) );
  XNOR2_X1 U9860 ( .A(n8625), .B(n8624), .ZN(P1_U3346) );
  AOI21_X1 U9861 ( .B1(n5025), .B2(n8627), .A(n8626), .ZN(n8642) );
  OAI21_X1 U9862 ( .B1(n8630), .B2(n8629), .A(n8628), .ZN(n8640) );
  AOI21_X1 U9863 ( .B1(n10495), .B2(P2_ADDR_REG_12__SCAN_IN), .A(n8631), .ZN(
        n8637) );
  OAI21_X1 U9864 ( .B1(n8634), .B2(n8633), .A(n8632), .ZN(n8635) );
  NAND2_X1 U9865 ( .A1(n8635), .A2(n10504), .ZN(n8636) );
  OAI211_X1 U9866 ( .C1(n10403), .C2(n8638), .A(n8637), .B(n8636), .ZN(n8639)
         );
  AOI21_X1 U9867 ( .B1(n8640), .B2(n10505), .A(n8639), .ZN(n8641) );
  OAI21_X1 U9868 ( .B1(n8642), .B2(n10511), .A(n8641), .ZN(P2_U3194) );
  OAI21_X1 U9869 ( .B1(n8645), .B2(n8644), .A(n8643), .ZN(n8720) );
  XNOR2_X1 U9870 ( .A(n8694), .B(n9115), .ZN(n8717) );
  XOR2_X1 U9871 ( .A(n9280), .B(n8717), .Z(n8719) );
  XNOR2_X1 U9872 ( .A(n8720), .B(n8719), .ZN(n8650) );
  NOR2_X1 U9873 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6455), .ZN(n9298) );
  AOI21_X1 U9874 ( .B1(n9281), .B2(n9261), .A(n9298), .ZN(n8647) );
  NAND2_X1 U9875 ( .A1(n9266), .A2(n10676), .ZN(n8646) );
  OAI211_X1 U9876 ( .C1(n9081), .C2(n9263), .A(n8647), .B(n8646), .ZN(n8648)
         );
  AOI21_X1 U9877 ( .B1(n8694), .B2(n9251), .A(n8648), .ZN(n8649) );
  OAI21_X1 U9878 ( .B1(n8650), .B2(n9254), .A(n8649), .ZN(P2_U3174) );
  INV_X1 U9879 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n8654) );
  AOI211_X1 U9880 ( .C1(n8653), .C2(n10667), .A(n8652), .B(n8651), .ZN(n8656)
         );
  MUX2_X1 U9881 ( .A(n8654), .B(n8656), .S(n10646), .Z(n8655) );
  OAI21_X1 U9882 ( .B1(n5192), .B2(n10219), .A(n8655), .ZN(P1_U3533) );
  INV_X1 U9883 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n8657) );
  MUX2_X1 U9884 ( .A(n8657), .B(n8656), .S(n10674), .Z(n8658) );
  OAI21_X1 U9885 ( .B1(n5192), .B2(n10267), .A(n8658), .ZN(P1_U3486) );
  XOR2_X1 U9886 ( .A(n8661), .B(n8659), .Z(n10668) );
  INV_X1 U9887 ( .A(n10668), .ZN(n8671) );
  OAI211_X1 U9888 ( .C1(n8662), .C2(n8661), .A(n8660), .B(n10127), .ZN(n8664)
         );
  AOI22_X1 U9889 ( .A1(n9804), .A2(n10557), .B1(n10558), .B2(n9802), .ZN(n8663) );
  NAND2_X1 U9890 ( .A1(n8664), .A2(n8663), .ZN(n10666) );
  OAI21_X1 U9891 ( .B1(n10662), .B2(n5023), .A(n4964), .ZN(n10664) );
  AOI22_X1 U9892 ( .A1(n4941), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n8705), .B2(
        n10572), .ZN(n8667) );
  NAND2_X1 U9893 ( .A1(n8665), .A2(n10570), .ZN(n8666) );
  OAI211_X1 U9894 ( .C1(n10664), .C2(n8668), .A(n8667), .B(n8666), .ZN(n8669)
         );
  AOI21_X1 U9895 ( .B1(n10666), .B2(n7834), .A(n8669), .ZN(n8670) );
  OAI21_X1 U9896 ( .B1(n8671), .B2(n10154), .A(n8670), .ZN(P1_U3281) );
  XNOR2_X1 U9897 ( .A(n8672), .B(n8987), .ZN(n9622) );
  INV_X1 U9898 ( .A(n9622), .ZN(n8680) );
  XNOR2_X1 U9899 ( .A(n8674), .B(n8673), .ZN(n8675) );
  OAI22_X1 U9900 ( .A1(n8675), .A2(n9498), .B1(n8718), .B2(n9515), .ZN(n9620)
         );
  INV_X1 U9901 ( .A(n8728), .ZN(n9619) );
  INV_X1 U9902 ( .A(n8724), .ZN(n8676) );
  OAI22_X1 U9903 ( .A1(n9619), .A2(n10585), .B1(n8676), .B2(n10677), .ZN(n8677) );
  OAI21_X1 U9904 ( .B1(n9620), .B2(n8677), .A(n10641), .ZN(n8679) );
  AOI22_X1 U9905 ( .A1(n9470), .A2(n9278), .B1(n10687), .B2(
        P2_REG2_REG_14__SCAN_IN), .ZN(n8678) );
  OAI211_X1 U9906 ( .C1(n8680), .C2(n9493), .A(n8679), .B(n8678), .ZN(P2_U3219) );
  XNOR2_X1 U9907 ( .A(n8682), .B(n8681), .ZN(n10240) );
  INV_X1 U9908 ( .A(n8803), .ZN(n8683) );
  AOI21_X1 U9909 ( .B1(n10235), .B2(n4964), .A(n8683), .ZN(n10236) );
  AOI22_X1 U9910 ( .A1(n10619), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n8739), .B2(
        n10572), .ZN(n8684) );
  OAI21_X1 U9911 ( .B1(n5821), .B2(n10612), .A(n8684), .ZN(n8690) );
  OAI21_X1 U9912 ( .B1(n8687), .B2(n8686), .A(n8685), .ZN(n8688) );
  AOI222_X1 U9913 ( .A1(n10127), .A2(n8688), .B1(n9801), .B2(n10558), .C1(
        n9803), .C2(n10557), .ZN(n10238) );
  NOR2_X1 U9914 ( .A1(n10238), .A2(n4941), .ZN(n8689) );
  AOI211_X1 U9915 ( .C1(n10236), .C2(n10002), .A(n8690), .B(n8689), .ZN(n8691)
         );
  OAI21_X1 U9916 ( .B1(n10154), .B2(n10240), .A(n8691), .ZN(P1_U3280) );
  XNOR2_X1 U9917 ( .A(n8692), .B(n8693), .ZN(n10684) );
  INV_X1 U9918 ( .A(n8694), .ZN(n8695) );
  NOR2_X1 U9919 ( .A1(n8695), .A2(n9618), .ZN(n10675) );
  XNOR2_X1 U9920 ( .A(n8696), .B(n8974), .ZN(n8697) );
  OAI222_X1 U9921 ( .A1(n9616), .A2(n9081), .B1(n9515), .B2(n8698), .C1(n8697), 
        .C2(n9498), .ZN(n10681) );
  AOI211_X1 U9922 ( .C1(n10684), .C2(n9623), .A(n10675), .B(n10681), .ZN(
        n10689) );
  NAND2_X1 U9923 ( .A1(n9624), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n8699) );
  OAI21_X1 U9924 ( .B1(n10689), .B2(n9624), .A(n8699), .ZN(P2_U3472) );
  INV_X1 U9925 ( .A(n8700), .ZN(n8704) );
  AOI21_X1 U9926 ( .B1(n8701), .B2(n8767), .A(n8702), .ZN(n8703) );
  OAI21_X1 U9927 ( .B1(n8704), .B2(n8703), .A(n9784), .ZN(n8711) );
  INV_X1 U9928 ( .A(n9788), .ZN(n9756) );
  INV_X1 U9929 ( .A(n8705), .ZN(n8707) );
  OAI22_X1 U9930 ( .A1(n9756), .A2(n8707), .B1(n9754), .B2(n8706), .ZN(n8708)
         );
  AOI211_X1 U9931 ( .C1(n9787), .C2(n9802), .A(n8709), .B(n8708), .ZN(n8710)
         );
  OAI211_X1 U9932 ( .C1(n10662), .C2(n8745), .A(n8711), .B(n8710), .ZN(
        P1_U3224) );
  INV_X1 U9933 ( .A(n9618), .ZN(n9610) );
  NOR2_X1 U9934 ( .A1(n8712), .A2(n9615), .ZN(n8714) );
  AOI211_X1 U9935 ( .C1(n9610), .C2(n8715), .A(n8714), .B(n8713), .ZN(n10661)
         );
  OR2_X1 U9936 ( .A1(n10661), .A2(n9624), .ZN(n8716) );
  OAI21_X1 U9937 ( .B1(n9627), .B2(n5094), .A(n8716), .ZN(P2_U3471) );
  XNOR2_X1 U9938 ( .A(n8728), .B(n9115), .ZN(n9082) );
  XOR2_X1 U9939 ( .A(n9279), .B(n9082), .Z(n8722) );
  AOI21_X1 U9940 ( .B1(n8722), .B2(n8721), .A(n5017), .ZN(n8730) );
  NOR2_X1 U9941 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8723), .ZN(n9315) );
  AOI21_X1 U9942 ( .B1(n9261), .B2(n9280), .A(n9315), .ZN(n8726) );
  NAND2_X1 U9943 ( .A1(n9266), .A2(n8724), .ZN(n8725) );
  OAI211_X1 U9944 ( .C1(n9617), .C2(n9263), .A(n8726), .B(n8725), .ZN(n8727)
         );
  AOI21_X1 U9945 ( .B1(n8728), .B2(n9251), .A(n8727), .ZN(n8729) );
  OAI21_X1 U9946 ( .B1(n8730), .B2(n9254), .A(n8729), .ZN(P2_U3155) );
  INV_X1 U9947 ( .A(n8731), .ZN(n9138) );
  INV_X1 U9948 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n8732) );
  OAI222_X1 U9949 ( .A1(n8733), .A2(P1_U3086), .B1(n10293), .B2(n9138), .C1(
        n8732), .C2(n10290), .ZN(P1_U3331) );
  AND2_X1 U9950 ( .A1(n8700), .A2(n8734), .ZN(n8737) );
  OAI211_X1 U9951 ( .C1(n8737), .C2(n8736), .A(n9784), .B(n8735), .ZN(n8744)
         );
  INV_X1 U9952 ( .A(n8738), .ZN(n8742) );
  INV_X1 U9953 ( .A(n8739), .ZN(n8740) );
  OAI22_X1 U9954 ( .A1(n9756), .A2(n8740), .B1(n9775), .B2(n8832), .ZN(n8741)
         );
  AOI211_X1 U9955 ( .C1(n9786), .C2(n9803), .A(n8742), .B(n8741), .ZN(n8743)
         );
  OAI211_X1 U9956 ( .C1(n5821), .C2(n8745), .A(n8744), .B(n8743), .ZN(P1_U3234) );
  XNOR2_X1 U9957 ( .A(n8746), .B(n8983), .ZN(n8754) );
  XNOR2_X1 U9958 ( .A(n8747), .B(n8983), .ZN(n8748) );
  OAI222_X1 U9959 ( .A1(n9515), .A2(n9081), .B1(n9616), .B2(n9264), .C1(n8748), 
        .C2(n9498), .ZN(n8756) );
  NAND2_X1 U9960 ( .A1(n8756), .A2(n10641), .ZN(n8753) );
  INV_X1 U9961 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n8750) );
  INV_X1 U9962 ( .A(n9267), .ZN(n8749) );
  OAI22_X1 U9963 ( .A1(n10641), .A2(n8750), .B1(n8749), .B2(n10677), .ZN(n8751) );
  AOI21_X1 U9964 ( .B1(n9083), .B2(n10636), .A(n8751), .ZN(n8752) );
  OAI211_X1 U9965 ( .C1(n8754), .C2(n9493), .A(n8753), .B(n8752), .ZN(P2_U3218) );
  INV_X1 U9966 ( .A(n9083), .ZN(n9271) );
  OAI22_X1 U9967 ( .A1(n8754), .A2(n9615), .B1(n9271), .B2(n9618), .ZN(n8755)
         );
  NOR2_X1 U9968 ( .A1(n8756), .A2(n8755), .ZN(n10694) );
  NAND2_X1 U9969 ( .A1(n9624), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n8757) );
  OAI21_X1 U9970 ( .B1(n10694), .B2(n9624), .A(n8757), .ZN(P2_U3474) );
  INV_X1 U9971 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n8758) );
  OAI222_X1 U9972 ( .A1(n8759), .A2(P1_U3086), .B1(n10293), .B2(n8785), .C1(
        n8758), .C2(n10290), .ZN(P1_U3330) );
  AOI22_X1 U9973 ( .A1(n9788), .A2(n8760), .B1(n9786), .B2(n9805), .ZN(n8762)
         );
  OAI211_X1 U9974 ( .C1(n8763), .C2(n9775), .A(n8762), .B(n8761), .ZN(n8770)
         );
  INV_X1 U9975 ( .A(n8701), .ZN(n8768) );
  AOI21_X1 U9976 ( .B1(n8765), .B2(n8767), .A(n8764), .ZN(n8766) );
  AOI211_X1 U9977 ( .C1(n8768), .C2(n8767), .A(n9778), .B(n8766), .ZN(n8769)
         );
  AOI211_X1 U9978 ( .C1(n8771), .C2(n9789), .A(n8770), .B(n8769), .ZN(n8772)
         );
  INV_X1 U9979 ( .A(n8772), .ZN(P1_U3236) );
  INV_X1 U9980 ( .A(n8993), .ZN(n8895) );
  XNOR2_X1 U9981 ( .A(n8773), .B(n8895), .ZN(n8774) );
  AOI22_X1 U9982 ( .A1(n8774), .A2(n9532), .B1(n9534), .B2(n9278), .ZN(n9613)
         );
  OR2_X1 U9983 ( .A1(n8775), .A2(n8993), .ZN(n8777) );
  NAND2_X1 U9984 ( .A1(n8775), .A2(n8993), .ZN(n8776) );
  NAND2_X1 U9985 ( .A1(n8777), .A2(n8776), .ZN(n9614) );
  INV_X1 U9986 ( .A(n9194), .ZN(n8778) );
  OAI22_X1 U9987 ( .A1(n10641), .A2(n7234), .B1(n8778), .B2(n10677), .ZN(n8779) );
  AOI21_X1 U9988 ( .B1(n9470), .B2(n9608), .A(n8779), .ZN(n8781) );
  NAND2_X1 U9989 ( .A1(n9611), .A2(n10636), .ZN(n8780) );
  OAI211_X1 U9990 ( .C1(n9614), .C2(n9493), .A(n8781), .B(n8780), .ZN(n8782)
         );
  INV_X1 U9991 ( .A(n8782), .ZN(n8783) );
  OAI21_X1 U9992 ( .B1(n9613), .B2(n10687), .A(n8783), .ZN(P2_U3217) );
  INV_X1 U9993 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n8784) );
  OAI222_X1 U9994 ( .A1(n9676), .A2(n8785), .B1(P2_U3151), .B2(n6885), .C1(
        n8784), .C2(n9137), .ZN(P2_U3270) );
  XNOR2_X1 U9995 ( .A(n8786), .B(n8792), .ZN(n10229) );
  INV_X1 U9996 ( .A(n10147), .ZN(n8788) );
  AOI21_X1 U9997 ( .B1(n10225), .B2(n8802), .A(n8788), .ZN(n10226) );
  AOI22_X1 U9998 ( .A1(n10619), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n8829), .B2(
        n10572), .ZN(n8789) );
  OAI21_X1 U9999 ( .B1(n8790), .B2(n10612), .A(n8789), .ZN(n8796) );
  NAND2_X1 U10000 ( .A1(n8806), .A2(n8791), .ZN(n8793) );
  XNOR2_X1 U10001 ( .A(n8793), .B(n8792), .ZN(n8794) );
  AOI222_X1 U10002 ( .A1(n10127), .A2(n8794), .B1(n9723), .B2(n10558), .C1(
        n9801), .C2(n10557), .ZN(n10228) );
  NOR2_X1 U10003 ( .A1(n10228), .A2(n4941), .ZN(n8795) );
  AOI211_X1 U10004 ( .C1(n10226), .C2(n10002), .A(n8796), .B(n8795), .ZN(n8797) );
  OAI21_X1 U10005 ( .B1(n10229), .B2(n10154), .A(n8797), .ZN(P1_U3278) );
  INV_X1 U10006 ( .A(n8798), .ZN(n8837) );
  AOI22_X1 U10007 ( .A1(n8799), .A2(P2_STATE_REG_SCAN_IN), .B1(n9674), .B2(
        P1_DATAO_REG_26__SCAN_IN), .ZN(n8800) );
  OAI21_X1 U10008 ( .B1(n8837), .B2(n9676), .A(n8800), .ZN(P2_U3269) );
  XNOR2_X1 U10009 ( .A(n8801), .B(n8809), .ZN(n10234) );
  AOI21_X1 U10010 ( .B1(n10230), .B2(n8803), .A(n8787), .ZN(n10231) );
  AOI22_X1 U10011 ( .A1(n10619), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n8819), 
        .B2(n10572), .ZN(n8804) );
  OAI21_X1 U10012 ( .B1(n8805), .B2(n10612), .A(n8804), .ZN(n8813) );
  AND2_X1 U10013 ( .A1(n9800), .A2(n10558), .ZN(n8811) );
  INV_X1 U10014 ( .A(n8806), .ZN(n8807) );
  AOI211_X1 U10015 ( .C1(n8809), .C2(n8808), .A(n10561), .B(n8807), .ZN(n8810)
         );
  AOI211_X1 U10016 ( .C1(n10557), .C2(n9802), .A(n8811), .B(n8810), .ZN(n10233) );
  NOR2_X1 U10017 ( .A1(n10233), .A2(n4941), .ZN(n8812) );
  AOI211_X1 U10018 ( .C1(n10231), .C2(n10002), .A(n8813), .B(n8812), .ZN(n8814) );
  OAI21_X1 U10019 ( .B1(n10154), .B2(n10234), .A(n8814), .ZN(P1_U3279) );
  NAND2_X1 U10020 ( .A1(n8816), .A2(n8815), .ZN(n8818) );
  XNOR2_X1 U10021 ( .A(n8818), .B(n8817), .ZN(n8824) );
  AOI22_X1 U10022 ( .A1(n8819), .A2(n9788), .B1(n9787), .B2(n9800), .ZN(n8821)
         );
  OAI211_X1 U10023 ( .C1(n5820), .C2(n9754), .A(n8821), .B(n8820), .ZN(n8822)
         );
  AOI21_X1 U10024 ( .B1(n10230), .B2(n9789), .A(n8822), .ZN(n8823) );
  OAI21_X1 U10025 ( .B1(n8824), .B2(n9778), .A(n8823), .ZN(P1_U3215) );
  XOR2_X1 U10026 ( .A(n8827), .B(n8826), .Z(n8828) );
  XNOR2_X1 U10027 ( .A(n8825), .B(n8828), .ZN(n8835) );
  AOI22_X1 U10028 ( .A1(n9788), .A2(n8829), .B1(n9787), .B2(n9723), .ZN(n8831)
         );
  OAI211_X1 U10029 ( .C1(n8832), .C2(n9754), .A(n8831), .B(n8830), .ZN(n8833)
         );
  AOI21_X1 U10030 ( .B1(n10225), .B2(n9789), .A(n8833), .ZN(n8834) );
  OAI21_X1 U10031 ( .B1(n8835), .B2(n9778), .A(n8834), .ZN(P1_U3241) );
  INV_X1 U10032 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n8836) );
  OAI222_X1 U10033 ( .A1(P1_U3086), .A2(n8838), .B1(n10293), .B2(n8837), .C1(
        n8836), .C2(n10290), .ZN(P1_U3329) );
  INV_X1 U10034 ( .A(n8841), .ZN(n8842) );
  NAND2_X1 U10035 ( .A1(n8843), .A2(n8842), .ZN(n9553) );
  MUX2_X1 U10036 ( .A(n9553), .B(P2_REG0_REG_29__SCAN_IN), .S(n10692), .Z(
        P2_U3456) );
  INV_X1 U10037 ( .A(n9062), .ZN(n8902) );
  NAND2_X1 U10038 ( .A1(n9663), .A2(n8849), .ZN(n8846) );
  NAND2_X1 U10039 ( .A1(n8844), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n8845) );
  INV_X1 U10040 ( .A(n9630), .ZN(n8864) );
  NAND2_X1 U10041 ( .A1(n8850), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n8855) );
  NAND2_X1 U10042 ( .A1(n8851), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n8854) );
  NAND2_X1 U10043 ( .A1(n8852), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n8853) );
  AND3_X1 U10044 ( .A1(n8855), .A2(n8854), .A3(n8853), .ZN(n8856) );
  NAND2_X1 U10045 ( .A1(n8857), .A2(n8856), .ZN(n9397) );
  NAND2_X1 U10046 ( .A1(n9630), .A2(n9397), .ZN(n9068) );
  OAI21_X1 U10047 ( .B1(n9633), .B2(n8864), .A(n9068), .ZN(n8859) );
  OAI21_X1 U10048 ( .B1(n9633), .B2(n9272), .A(n8858), .ZN(n9065) );
  AOI21_X1 U10049 ( .B1(n8861), .B2(n8902), .A(n8860), .ZN(n8910) );
  INV_X1 U10050 ( .A(n9064), .ZN(n8865) );
  NAND2_X1 U10051 ( .A1(n8865), .A2(n8864), .ZN(n8868) );
  NOR2_X1 U10052 ( .A1(n9630), .A2(n9397), .ZN(n9067) );
  NOR2_X1 U10053 ( .A1(n9067), .A2(n8927), .ZN(n8867) );
  INV_X1 U10054 ( .A(n9068), .ZN(n8906) );
  NAND2_X1 U10055 ( .A1(n8870), .A2(n8869), .ZN(n9412) );
  NAND2_X1 U10056 ( .A1(n9409), .A2(n9047), .ZN(n9419) );
  INV_X1 U10057 ( .A(n9419), .ZN(n9416) );
  NAND2_X1 U10058 ( .A1(n9043), .A2(n8871), .ZN(n9426) );
  NAND2_X1 U10059 ( .A1(n8872), .A2(n9038), .ZN(n9441) );
  INV_X1 U10060 ( .A(n9478), .ZN(n8899) );
  NAND2_X1 U10061 ( .A1(n8874), .A2(n8873), .ZN(n9460) );
  INV_X1 U10062 ( .A(n8875), .ZN(n8876) );
  NOR2_X1 U10063 ( .A1(n8877), .A2(n8876), .ZN(n8881) );
  NOR2_X1 U10064 ( .A1(n6850), .A2(n6851), .ZN(n8880) );
  NAND4_X1 U10065 ( .A1(n8881), .A2(n8880), .A3(n8879), .A4(n8878), .ZN(n8883)
         );
  NOR2_X1 U10066 ( .A1(n8883), .A2(n8882), .ZN(n8884) );
  NAND3_X1 U10067 ( .A1(n8886), .A2(n8885), .A3(n8884), .ZN(n8887) );
  NOR2_X1 U10068 ( .A1(n8888), .A2(n8887), .ZN(n8889) );
  NAND4_X1 U10069 ( .A1(n8891), .A2(n8890), .A3(n8976), .A4(n8889), .ZN(n8892)
         );
  NOR2_X1 U10070 ( .A1(n8892), .A2(n8974), .ZN(n8893) );
  NAND4_X1 U10071 ( .A1(n8895), .A2(n8894), .A3(n8893), .A4(n8987), .ZN(n8896)
         );
  NOR3_X1 U10072 ( .A1(n9525), .A2(n9538), .A3(n8896), .ZN(n8897) );
  NAND4_X1 U10073 ( .A1(n9460), .A2(n9504), .A3(n8897), .A4(n9017), .ZN(n8898)
         );
  NOR4_X1 U10074 ( .A1(n9426), .A2(n9441), .A3(n8899), .A4(n8898), .ZN(n8900)
         );
  NAND3_X1 U10075 ( .A1(n9416), .A2(n8900), .A3(n9444), .ZN(n8901) );
  NOR2_X1 U10076 ( .A1(n9412), .A2(n8901), .ZN(n8903) );
  NAND4_X1 U10077 ( .A1(n9064), .A2(n8904), .A3(n8903), .A4(n8902), .ZN(n8905)
         );
  NOR4_X1 U10078 ( .A1(n9067), .A2(n8906), .A3(n9065), .A4(n8905), .ZN(n8907)
         );
  NAND2_X1 U10079 ( .A1(n8907), .A2(n8927), .ZN(n8908) );
  OAI21_X1 U10080 ( .B1(n8910), .B2(n8909), .A(n8908), .ZN(n8912) );
  MUX2_X1 U10081 ( .A(n9585), .B(n9581), .S(n9060), .Z(n9026) );
  INV_X1 U10082 ( .A(n9026), .ZN(n9030) );
  OR2_X1 U10083 ( .A1(n8915), .A2(n8961), .ZN(n8959) );
  INV_X1 U10084 ( .A(n8916), .ZN(n8917) );
  NOR2_X1 U10085 ( .A1(n8918), .A2(n8917), .ZN(n8920) );
  OAI211_X1 U10086 ( .C1(n8959), .C2(n8920), .A(n8919), .B(n8964), .ZN(n8957)
         );
  AOI21_X1 U10087 ( .B1(n8925), .B2(n8928), .A(n8924), .ZN(n8923) );
  OAI211_X1 U10088 ( .C1(n8923), .C2(n6851), .A(n8922), .B(n8936), .ZN(n8934)
         );
  AOI211_X1 U10089 ( .C1(n8927), .C2(n8926), .A(n8925), .B(n8924), .ZN(n8930)
         );
  NOR2_X1 U10090 ( .A1(n8930), .A2(n8929), .ZN(n8932) );
  OAI211_X1 U10091 ( .C1(n8932), .C2(n6851), .A(n8931), .B(n8943), .ZN(n8933)
         );
  MUX2_X1 U10092 ( .A(n8934), .B(n8933), .S(n9053), .Z(n8935) );
  NAND2_X1 U10093 ( .A1(n8935), .A2(n8938), .ZN(n8945) );
  NAND2_X1 U10094 ( .A1(n8937), .A2(n8936), .ZN(n8939) );
  OAI211_X1 U10095 ( .C1(n8945), .C2(n8939), .A(n8938), .B(n8946), .ZN(n8941)
         );
  NAND3_X1 U10096 ( .A1(n8941), .A2(n8950), .A3(n8940), .ZN(n8942) );
  NAND2_X1 U10097 ( .A1(n8942), .A2(n8947), .ZN(n8953) );
  INV_X1 U10098 ( .A(n8943), .ZN(n8944) );
  NOR2_X1 U10099 ( .A1(n8945), .A2(n8944), .ZN(n8949) );
  OAI211_X1 U10100 ( .C1(n8949), .C2(n8948), .A(n8947), .B(n8946), .ZN(n8951)
         );
  NAND2_X1 U10101 ( .A1(n8951), .A2(n8950), .ZN(n8952) );
  MUX2_X1 U10102 ( .A(n8953), .B(n8952), .S(n9060), .Z(n8955) );
  NOR3_X1 U10103 ( .A1(n8955), .A2(n8954), .A3(n8959), .ZN(n8956) );
  AOI21_X1 U10104 ( .B1(n9060), .B2(n8957), .A(n8956), .ZN(n8968) );
  NOR3_X1 U10105 ( .A1(n8968), .A2(n8969), .A3(n8960), .ZN(n8958) );
  INV_X1 U10106 ( .A(n8959), .ZN(n8963) );
  AOI211_X1 U10107 ( .C1(n8963), .C2(n8962), .A(n8961), .B(n8960), .ZN(n8967)
         );
  INV_X1 U10108 ( .A(n8964), .ZN(n8966) );
  AOI211_X1 U10109 ( .C1(n8968), .C2(n8967), .A(n8966), .B(n8965), .ZN(n8970)
         );
  INV_X1 U10110 ( .A(n8971), .ZN(n8972) );
  MUX2_X1 U10111 ( .A(n8973), .B(n8972), .S(n9053), .Z(n8975) );
  INV_X1 U10112 ( .A(n8977), .ZN(n8980) );
  INV_X1 U10113 ( .A(n8978), .ZN(n8979) );
  MUX2_X1 U10114 ( .A(n8980), .B(n8979), .S(n9053), .Z(n8981) );
  NOR3_X1 U10115 ( .A1(n8988), .A2(n8983), .A3(n8982), .ZN(n8996) );
  NAND2_X1 U10116 ( .A1(n8990), .A2(n9081), .ZN(n8985) );
  NAND2_X1 U10117 ( .A1(n8989), .A2(n9619), .ZN(n8984) );
  MUX2_X1 U10118 ( .A(n8985), .B(n8984), .S(n9053), .Z(n8986) );
  AOI21_X1 U10119 ( .B1(n8988), .B2(n8987), .A(n8986), .ZN(n8995) );
  INV_X1 U10120 ( .A(n8989), .ZN(n8992) );
  INV_X1 U10121 ( .A(n8990), .ZN(n8991) );
  MUX2_X1 U10122 ( .A(n8992), .B(n8991), .S(n9053), .Z(n8994) );
  NOR4_X1 U10123 ( .A1(n8996), .A2(n8995), .A3(n8994), .A4(n8993), .ZN(n9002)
         );
  INV_X1 U10124 ( .A(n8997), .ZN(n9000) );
  INV_X1 U10125 ( .A(n8998), .ZN(n8999) );
  MUX2_X1 U10126 ( .A(n9000), .B(n8999), .S(n9060), .Z(n9001) );
  NOR2_X1 U10127 ( .A1(n9002), .A2(n9001), .ZN(n9014) );
  MUX2_X1 U10128 ( .A(n9608), .B(n9602), .S(n9053), .Z(n9006) );
  NAND2_X1 U10129 ( .A1(n9003), .A2(n9006), .ZN(n9005) );
  MUX2_X1 U10130 ( .A(n9009), .B(n9007), .S(n9060), .Z(n9004) );
  OAI211_X1 U10131 ( .C1(n9014), .C2(n9005), .A(n9504), .B(n9004), .ZN(n9020)
         );
  INV_X1 U10132 ( .A(n9006), .ZN(n9013) );
  NAND2_X1 U10133 ( .A1(n9007), .A2(n9516), .ZN(n9011) );
  INV_X1 U10134 ( .A(n9602), .ZN(n9008) );
  NAND2_X1 U10135 ( .A1(n9009), .A2(n9008), .ZN(n9010) );
  MUX2_X1 U10136 ( .A(n9011), .B(n9010), .S(n9060), .Z(n9012) );
  AOI21_X1 U10137 ( .B1(n9014), .B2(n9013), .A(n9012), .ZN(n9019) );
  MUX2_X1 U10138 ( .A(n9016), .B(n9015), .S(n9053), .Z(n9018) );
  OAI211_X1 U10139 ( .C1(n9020), .C2(n9019), .A(n9018), .B(n9017), .ZN(n9025)
         );
  NAND2_X1 U10140 ( .A1(n9586), .A2(n9053), .ZN(n9023) );
  INV_X1 U10141 ( .A(n9586), .ZN(n9021) );
  NAND2_X1 U10142 ( .A1(n9021), .A2(n9060), .ZN(n9022) );
  MUX2_X1 U10143 ( .A(n9023), .B(n9022), .S(n9468), .Z(n9024) );
  OAI211_X1 U10144 ( .C1(n9027), .C2(n9026), .A(n9025), .B(n9024), .ZN(n9028)
         );
  OAI21_X1 U10145 ( .B1(n9030), .B2(n9029), .A(n9028), .ZN(n9033) );
  NOR3_X1 U10146 ( .A1(n9648), .A2(n9053), .A3(n9580), .ZN(n9032) );
  NOR3_X1 U10147 ( .A1(n9099), .A2(n9060), .A3(n9101), .ZN(n9031) );
  AOI211_X1 U10148 ( .C1(n9033), .C2(n9460), .A(n9032), .B(n9031), .ZN(n9037)
         );
  NOR2_X1 U10149 ( .A1(n9572), .A2(n9060), .ZN(n9035) );
  AOI211_X1 U10150 ( .C1(n9459), .C2(n9060), .A(n9035), .B(n9034), .ZN(n9036)
         );
  AOI211_X1 U10151 ( .C1(n9037), .C2(n9444), .A(n9036), .B(n9441), .ZN(n9042)
         );
  INV_X1 U10152 ( .A(n9038), .ZN(n9040) );
  MUX2_X1 U10153 ( .A(n9040), .B(n9039), .S(n9053), .Z(n9041) );
  NOR3_X1 U10154 ( .A1(n9042), .A2(n9041), .A3(n9426), .ZN(n9046) );
  MUX2_X1 U10155 ( .A(n9044), .B(n5327), .S(n9060), .Z(n9045) );
  MUX2_X1 U10156 ( .A(n9047), .B(n9409), .S(n9053), .Z(n9051) );
  MUX2_X1 U10157 ( .A(n9049), .B(n9048), .S(n9060), .Z(n9050) );
  MUX2_X1 U10158 ( .A(n9408), .B(n9052), .S(n9060), .Z(n9055) );
  INV_X1 U10159 ( .A(n9055), .ZN(n9058) );
  MUX2_X1 U10160 ( .A(n9554), .B(n9145), .S(n9053), .Z(n9054) );
  OAI21_X1 U10161 ( .B1(n9056), .B2(n9055), .A(n9054), .ZN(n9057) );
  OAI21_X1 U10162 ( .B1(n9059), .B2(n9058), .A(n9057), .ZN(n9061) );
  XNOR2_X1 U10163 ( .A(n9061), .B(n9060), .ZN(n9063) );
  NOR2_X1 U10164 ( .A1(n9063), .A2(n9062), .ZN(n9066) );
  OAI21_X1 U10165 ( .B1(n9066), .B2(n9065), .A(n9064), .ZN(n9069) );
  AOI21_X1 U10166 ( .B1(n9069), .B2(n9068), .A(n9067), .ZN(n9071) );
  NAND3_X1 U10167 ( .A1(n9076), .A2(n9075), .A3(n9074), .ZN(n9077) );
  OAI211_X1 U10168 ( .C1(n9078), .C2(n9080), .A(n9077), .B(P2_B_REG_SCAN_IN), 
        .ZN(n9079) );
  XNOR2_X1 U10169 ( .A(n9083), .B(n9115), .ZN(n9084) );
  XNOR2_X1 U10170 ( .A(n9084), .B(n9278), .ZN(n9258) );
  INV_X1 U10171 ( .A(n9084), .ZN(n9085) );
  XNOR2_X1 U10172 ( .A(n9611), .B(n9115), .ZN(n9087) );
  XNOR2_X1 U10173 ( .A(n9087), .B(n9535), .ZN(n9192) );
  INV_X1 U10174 ( .A(n9087), .ZN(n9088) );
  XNOR2_X1 U10175 ( .A(n9602), .B(n9110), .ZN(n9201) );
  INV_X1 U10176 ( .A(n9201), .ZN(n9089) );
  XNOR2_X1 U10177 ( .A(n9524), .B(n9115), .ZN(n9090) );
  XNOR2_X1 U10178 ( .A(n9090), .B(n9277), .ZN(n9235) );
  NAND2_X1 U10179 ( .A1(n9236), .A2(n9235), .ZN(n9234) );
  NAND2_X1 U10180 ( .A1(n9234), .A2(n9091), .ZN(n9172) );
  XNOR2_X1 U10181 ( .A(n9092), .B(n9110), .ZN(n9171) );
  INV_X1 U10182 ( .A(n9171), .ZN(n9093) );
  XNOR2_X1 U10183 ( .A(n9586), .B(n9115), .ZN(n9096) );
  XOR2_X1 U10184 ( .A(n9468), .B(n9096), .Z(n9221) );
  XNOR2_X1 U10185 ( .A(n9581), .B(n9115), .ZN(n9098) );
  XNOR2_X1 U10186 ( .A(n9098), .B(n9585), .ZN(n9179) );
  XNOR2_X1 U10187 ( .A(n9099), .B(n9115), .ZN(n9100) );
  XNOR2_X1 U10188 ( .A(n9100), .B(n9580), .ZN(n9228) );
  NAND2_X1 U10189 ( .A1(n9227), .A2(n9103), .ZN(n9104) );
  XNOR2_X1 U10190 ( .A(n9572), .B(n9115), .ZN(n9105) );
  INV_X1 U10191 ( .A(n9104), .ZN(n9106) );
  XNOR2_X1 U10192 ( .A(n9215), .B(n9115), .ZN(n9107) );
  XOR2_X1 U10193 ( .A(n9446), .B(n9107), .Z(n9211) );
  INV_X1 U10194 ( .A(n9107), .ZN(n9108) );
  XNOR2_X1 U10195 ( .A(n9564), .B(n9115), .ZN(n9109) );
  XNOR2_X1 U10196 ( .A(n9109), .B(n9275), .ZN(n9186) );
  XNOR2_X1 U10197 ( .A(n9252), .B(n9110), .ZN(n9246) );
  INV_X1 U10198 ( .A(n9246), .ZN(n9112) );
  XNOR2_X1 U10199 ( .A(n9555), .B(n9115), .ZN(n9113) );
  XNOR2_X1 U10200 ( .A(n9113), .B(n9274), .ZN(n9155) );
  INV_X1 U10201 ( .A(n9113), .ZN(n9114) );
  XNOR2_X1 U10202 ( .A(n9116), .B(n9115), .ZN(n9117) );
  XNOR2_X1 U10203 ( .A(n9118), .B(n9117), .ZN(n9123) );
  NAND2_X1 U10204 ( .A1(n9273), .A2(n9238), .ZN(n9120) );
  AOI22_X1 U10205 ( .A1(n9139), .A2(n9266), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3151), .ZN(n9119) );
  OAI211_X1 U10206 ( .C1(n6814), .C2(n9240), .A(n9120), .B(n9119), .ZN(n9121)
         );
  AOI21_X1 U10207 ( .B1(n9145), .B2(n9251), .A(n9121), .ZN(n9122) );
  OAI21_X1 U10208 ( .B1(n9123), .B2(n9254), .A(n9122), .ZN(P2_U3160) );
  INV_X1 U10209 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n9129) );
  XNOR2_X1 U10210 ( .A(n9931), .B(n4948), .ZN(n9125) );
  NAND2_X1 U10211 ( .A1(n9125), .A2(n10552), .ZN(n9930) );
  INV_X1 U10212 ( .A(P1_B_REG_SCAN_IN), .ZN(n9126) );
  NOR2_X1 U10213 ( .A1(n10294), .A2(n9126), .ZN(n9127) );
  OR2_X1 U10214 ( .A1(n10145), .A2(n9127), .ZN(n9938) );
  INV_X1 U10215 ( .A(n9938), .ZN(n9128) );
  NAND2_X1 U10216 ( .A1(n5408), .A2(n9128), .ZN(n10155) );
  MUX2_X1 U10217 ( .A(n9129), .B(n9131), .S(n10674), .Z(n9130) );
  OAI21_X1 U10218 ( .B1(n4948), .B2(n10267), .A(n9130), .ZN(P1_U3521) );
  INV_X1 U10219 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n9132) );
  MUX2_X1 U10220 ( .A(n9132), .B(n9131), .S(n10646), .Z(n9133) );
  OAI21_X1 U10221 ( .B1(n4948), .B2(n10219), .A(n9133), .ZN(P1_U3553) );
  INV_X1 U10222 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n9134) );
  OAI222_X1 U10223 ( .A1(n6070), .A2(P1_U3086), .B1(n10293), .B2(n9135), .C1(
        n9134), .C2(n10290), .ZN(P1_U3336) );
  OAI222_X1 U10224 ( .A1(n9676), .A2(n9138), .B1(n9137), .B2(n9136), .C1(n6881), .C2(P2_U3151), .ZN(P2_U3271) );
  INV_X1 U10225 ( .A(n9139), .ZN(n9141) );
  OAI22_X1 U10226 ( .A1(n9141), .A2(n10677), .B1(n10641), .B2(n9140), .ZN(
        n9144) );
  NOR2_X1 U10227 ( .A1(n9142), .A2(n9493), .ZN(n9143) );
  AOI211_X1 U10228 ( .C1(n10636), .C2(n9145), .A(n9144), .B(n9143), .ZN(n9146)
         );
  OAI21_X1 U10229 ( .B1(n9147), .B2(n10687), .A(n9146), .ZN(P2_U3205) );
  INV_X1 U10230 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n10358) );
  OAI22_X1 U10231 ( .A1(n9509), .A2(n9148), .B1(n10358), .B2(n10677), .ZN(
        n9153) );
  NOR4_X1 U10232 ( .A1(n9151), .A2(n9150), .A3(n9610), .A4(n9149), .ZN(n9152)
         );
  AOI211_X1 U10233 ( .C1(n10687), .C2(P2_REG2_REG_0__SCAN_IN), .A(n9153), .B(
        n9152), .ZN(n9154) );
  OAI21_X1 U10234 ( .B1(n7503), .B2(n9545), .A(n9154), .ZN(P2_U3233) );
  XNOR2_X1 U10235 ( .A(n9156), .B(n9155), .ZN(n9161) );
  NAND2_X1 U10236 ( .A1(n9554), .A2(n9238), .ZN(n9158) );
  AOI22_X1 U10237 ( .A1(n9406), .A2(n9266), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3151), .ZN(n9157) );
  OAI211_X1 U10238 ( .C1(n9245), .C2(n9240), .A(n9158), .B(n9157), .ZN(n9159)
         );
  AOI21_X1 U10239 ( .B1(n9555), .B2(n9251), .A(n9159), .ZN(n9160) );
  OAI21_X1 U10240 ( .B1(n9161), .B2(n9254), .A(n9160), .ZN(P2_U3154) );
  XNOR2_X1 U10241 ( .A(n9162), .B(n9276), .ZN(n9168) );
  AOI22_X1 U10242 ( .A1(n9580), .A2(n9261), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3151), .ZN(n9164) );
  NAND2_X1 U10243 ( .A1(n9448), .A2(n9266), .ZN(n9163) );
  OAI211_X1 U10244 ( .C1(n9165), .C2(n9263), .A(n9164), .B(n9163), .ZN(n9166)
         );
  AOI21_X1 U10245 ( .B1(n9572), .B2(n9251), .A(n9166), .ZN(n9167) );
  OAI21_X1 U10246 ( .B1(n9168), .B2(n9254), .A(n9167), .ZN(P2_U3156) );
  INV_X1 U10247 ( .A(n9169), .ZN(n9655) );
  OAI211_X1 U10248 ( .C1(n9172), .C2(n9171), .A(n9170), .B(n9256), .ZN(n9177)
         );
  NAND2_X1 U10249 ( .A1(n9468), .A2(n9238), .ZN(n9174) );
  OAI211_X1 U10250 ( .C1(n9604), .C2(n9240), .A(n9174), .B(n9173), .ZN(n9175)
         );
  AOI21_X1 U10251 ( .B1(n9507), .B2(n9266), .A(n9175), .ZN(n9176) );
  OAI211_X1 U10252 ( .C1(n9655), .C2(n9270), .A(n9177), .B(n9176), .ZN(
        P2_U3159) );
  XOR2_X1 U10253 ( .A(n9179), .B(n9178), .Z(n9184) );
  AOI22_X1 U10254 ( .A1(n9580), .A2(n9238), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3151), .ZN(n9181) );
  NAND2_X1 U10255 ( .A1(n9266), .A2(n9471), .ZN(n9180) );
  OAI211_X1 U10256 ( .C1(n9500), .C2(n9240), .A(n9181), .B(n9180), .ZN(n9182)
         );
  AOI21_X1 U10257 ( .B1(n9581), .B2(n9251), .A(n9182), .ZN(n9183) );
  OAI21_X1 U10258 ( .B1(n9184), .B2(n9254), .A(n9183), .ZN(P2_U3163) );
  XOR2_X1 U10259 ( .A(n9186), .B(n9185), .Z(n9191) );
  AOI22_X1 U10260 ( .A1(n9446), .A2(n9261), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3151), .ZN(n9188) );
  NAND2_X1 U10261 ( .A1(n9429), .A2(n9266), .ZN(n9187) );
  OAI211_X1 U10262 ( .C1(n9245), .C2(n9263), .A(n9188), .B(n9187), .ZN(n9189)
         );
  AOI21_X1 U10263 ( .B1(n9564), .B2(n9251), .A(n9189), .ZN(n9190) );
  OAI21_X1 U10264 ( .B1(n9191), .B2(n9254), .A(n9190), .ZN(P2_U3165) );
  XNOR2_X1 U10265 ( .A(n9193), .B(n9192), .ZN(n9200) );
  NAND2_X1 U10266 ( .A1(n9266), .A2(n9194), .ZN(n9197) );
  NOR2_X1 U10267 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9195), .ZN(n9349) );
  AOI21_X1 U10268 ( .B1(n9238), .B2(n9608), .A(n9349), .ZN(n9196) );
  OAI211_X1 U10269 ( .C1(n9617), .C2(n9240), .A(n9197), .B(n9196), .ZN(n9198)
         );
  AOI21_X1 U10270 ( .B1(n9611), .B2(n9251), .A(n9198), .ZN(n9199) );
  OAI21_X1 U10271 ( .B1(n9200), .B2(n9254), .A(n9199), .ZN(P2_U3166) );
  XNOR2_X1 U10272 ( .A(n9201), .B(n9608), .ZN(n9202) );
  XNOR2_X1 U10273 ( .A(n9203), .B(n9202), .ZN(n9209) );
  NOR2_X1 U10274 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9204), .ZN(n9370) );
  AOI21_X1 U10275 ( .B1(n9261), .B2(n9535), .A(n9370), .ZN(n9206) );
  NAND2_X1 U10276 ( .A1(n9266), .A2(n9542), .ZN(n9205) );
  OAI211_X1 U10277 ( .C1(n9604), .C2(n9263), .A(n9206), .B(n9205), .ZN(n9207)
         );
  AOI21_X1 U10278 ( .B1(n9602), .B2(n9251), .A(n9207), .ZN(n9208) );
  OAI21_X1 U10279 ( .B1(n9209), .B2(n9254), .A(n9208), .ZN(P2_U3168) );
  XOR2_X1 U10280 ( .A(n9211), .B(n9210), .Z(n9217) );
  AOI22_X1 U10281 ( .A1(n9276), .A2(n9261), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3151), .ZN(n9213) );
  NAND2_X1 U10282 ( .A1(n9440), .A2(n9266), .ZN(n9212) );
  OAI211_X1 U10283 ( .C1(n9438), .C2(n9263), .A(n9213), .B(n9212), .ZN(n9214)
         );
  AOI21_X1 U10284 ( .B1(n9215), .B2(n9251), .A(n9214), .ZN(n9216) );
  OAI21_X1 U10285 ( .B1(n9217), .B2(n9254), .A(n9216), .ZN(P2_U3169) );
  INV_X1 U10286 ( .A(n9218), .ZN(n9219) );
  AOI21_X1 U10287 ( .B1(n9221), .B2(n9220), .A(n9219), .ZN(n9226) );
  AOI22_X1 U10288 ( .A1(n9585), .A2(n9238), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3151), .ZN(n9223) );
  NAND2_X1 U10289 ( .A1(n9266), .A2(n9486), .ZN(n9222) );
  OAI211_X1 U10290 ( .C1(n9517), .C2(n9240), .A(n9223), .B(n9222), .ZN(n9224)
         );
  AOI21_X1 U10291 ( .B1(n9586), .B2(n9251), .A(n9224), .ZN(n9225) );
  OAI21_X1 U10292 ( .B1(n9226), .B2(n9254), .A(n9225), .ZN(P2_U3173) );
  OAI211_X1 U10293 ( .C1(n9229), .C2(n9228), .A(n9227), .B(n9256), .ZN(n9233)
         );
  AOI22_X1 U10294 ( .A1(n9585), .A2(n9261), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3151), .ZN(n9230) );
  OAI21_X1 U10295 ( .B1(n9459), .B2(n9263), .A(n9230), .ZN(n9231) );
  AOI21_X1 U10296 ( .B1(n9462), .B2(n9266), .A(n9231), .ZN(n9232) );
  OAI211_X1 U10297 ( .C1(n9648), .C2(n9270), .A(n9233), .B(n9232), .ZN(
        P2_U3175) );
  OAI211_X1 U10298 ( .C1(n9236), .C2(n9235), .A(n9234), .B(n9256), .ZN(n9243)
         );
  NOR2_X1 U10299 ( .A1(n9237), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9386) );
  AOI21_X1 U10300 ( .B1(n9484), .B2(n9238), .A(n9386), .ZN(n9239) );
  OAI21_X1 U10301 ( .B1(n9516), .B2(n9240), .A(n9239), .ZN(n9241) );
  AOI21_X1 U10302 ( .B1(n9521), .B2(n9266), .A(n9241), .ZN(n9242) );
  OAI211_X1 U10303 ( .C1(n9598), .C2(n9270), .A(n9243), .B(n9242), .ZN(
        P2_U3178) );
  XNOR2_X1 U10304 ( .A(n9246), .B(n9245), .ZN(n9247) );
  XNOR2_X1 U10305 ( .A(n9244), .B(n9247), .ZN(n9255) );
  AOI22_X1 U10306 ( .A1(n9275), .A2(n9261), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3151), .ZN(n9249) );
  NAND2_X1 U10307 ( .A1(n9420), .A2(n9266), .ZN(n9248) );
  OAI211_X1 U10308 ( .C1(n6814), .C2(n9263), .A(n9249), .B(n9248), .ZN(n9250)
         );
  AOI21_X1 U10309 ( .B1(n9252), .B2(n9251), .A(n9250), .ZN(n9253) );
  OAI21_X1 U10310 ( .B1(n9255), .B2(n9254), .A(n9253), .ZN(P2_U3180) );
  OAI211_X1 U10311 ( .C1(n9259), .C2(n9258), .A(n9257), .B(n9256), .ZN(n9269)
         );
  NOR2_X1 U10312 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9260), .ZN(n9332) );
  AOI21_X1 U10313 ( .B1(n9261), .B2(n9279), .A(n9332), .ZN(n9262) );
  OAI21_X1 U10314 ( .B1(n9264), .B2(n9263), .A(n9262), .ZN(n9265) );
  AOI21_X1 U10315 ( .B1(n9267), .B2(n9266), .A(n9265), .ZN(n9268) );
  OAI211_X1 U10316 ( .C1(n9271), .C2(n9270), .A(n9269), .B(n9268), .ZN(
        P2_U3181) );
  MUX2_X1 U10317 ( .A(n9397), .B(P2_DATAO_REG_31__SCAN_IN), .S(n9292), .Z(
        P2_U3522) );
  MUX2_X1 U10318 ( .A(n9272), .B(P2_DATAO_REG_30__SCAN_IN), .S(n9292), .Z(
        P2_U3521) );
  MUX2_X1 U10319 ( .A(n9273), .B(P2_DATAO_REG_29__SCAN_IN), .S(n9292), .Z(
        P2_U3520) );
  MUX2_X1 U10320 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n9554), .S(P2_U3893), .Z(
        P2_U3519) );
  MUX2_X1 U10321 ( .A(n9274), .B(P2_DATAO_REG_27__SCAN_IN), .S(n9292), .Z(
        P2_U3518) );
  MUX2_X1 U10322 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n9563), .S(P2_U3893), .Z(
        P2_U3517) );
  MUX2_X1 U10323 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n9275), .S(P2_U3893), .Z(
        P2_U3516) );
  MUX2_X1 U10324 ( .A(n9446), .B(P2_DATAO_REG_24__SCAN_IN), .S(n9292), .Z(
        P2_U3515) );
  MUX2_X1 U10325 ( .A(n9276), .B(P2_DATAO_REG_23__SCAN_IN), .S(n9292), .Z(
        P2_U3514) );
  MUX2_X1 U10326 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n9580), .S(P2_U3893), .Z(
        P2_U3513) );
  MUX2_X1 U10327 ( .A(n9468), .B(P2_DATAO_REG_20__SCAN_IN), .S(n9292), .Z(
        P2_U3511) );
  MUX2_X1 U10328 ( .A(n9484), .B(P2_DATAO_REG_19__SCAN_IN), .S(n9292), .Z(
        P2_U3510) );
  MUX2_X1 U10329 ( .A(n9277), .B(P2_DATAO_REG_18__SCAN_IN), .S(n9292), .Z(
        P2_U3509) );
  MUX2_X1 U10330 ( .A(n9608), .B(P2_DATAO_REG_17__SCAN_IN), .S(n9292), .Z(
        P2_U3508) );
  MUX2_X1 U10331 ( .A(n9535), .B(P2_DATAO_REG_16__SCAN_IN), .S(n9292), .Z(
        P2_U3507) );
  MUX2_X1 U10332 ( .A(n9278), .B(P2_DATAO_REG_15__SCAN_IN), .S(n9292), .Z(
        P2_U3506) );
  MUX2_X1 U10333 ( .A(n9279), .B(P2_DATAO_REG_14__SCAN_IN), .S(n9292), .Z(
        P2_U3505) );
  MUX2_X1 U10334 ( .A(n9280), .B(P2_DATAO_REG_13__SCAN_IN), .S(n9292), .Z(
        P2_U3504) );
  MUX2_X1 U10335 ( .A(n9281), .B(P2_DATAO_REG_12__SCAN_IN), .S(n9292), .Z(
        P2_U3503) );
  MUX2_X1 U10336 ( .A(n9282), .B(P2_DATAO_REG_11__SCAN_IN), .S(n9292), .Z(
        P2_U3502) );
  MUX2_X1 U10337 ( .A(n9283), .B(P2_DATAO_REG_10__SCAN_IN), .S(n9292), .Z(
        P2_U3501) );
  MUX2_X1 U10338 ( .A(n9284), .B(P2_DATAO_REG_9__SCAN_IN), .S(n9292), .Z(
        P2_U3500) );
  MUX2_X1 U10339 ( .A(n9285), .B(P2_DATAO_REG_8__SCAN_IN), .S(n9292), .Z(
        P2_U3499) );
  MUX2_X1 U10340 ( .A(n9286), .B(P2_DATAO_REG_7__SCAN_IN), .S(n9292), .Z(
        P2_U3498) );
  MUX2_X1 U10341 ( .A(n9287), .B(P2_DATAO_REG_6__SCAN_IN), .S(n9292), .Z(
        P2_U3497) );
  MUX2_X1 U10342 ( .A(n9288), .B(P2_DATAO_REG_5__SCAN_IN), .S(n9292), .Z(
        P2_U3496) );
  MUX2_X1 U10343 ( .A(n9289), .B(P2_DATAO_REG_4__SCAN_IN), .S(n9292), .Z(
        P2_U3495) );
  MUX2_X1 U10344 ( .A(n9290), .B(P2_DATAO_REG_3__SCAN_IN), .S(n9292), .Z(
        P2_U3494) );
  MUX2_X1 U10345 ( .A(n9291), .B(P2_DATAO_REG_2__SCAN_IN), .S(n9292), .Z(
        P2_U3493) );
  MUX2_X1 U10346 ( .A(n7527), .B(P2_DATAO_REG_1__SCAN_IN), .S(n9292), .Z(
        P2_U3492) );
  AOI21_X1 U10347 ( .B1(n9295), .B2(n9294), .A(n9293), .ZN(n9309) );
  OAI21_X1 U10348 ( .B1(P2_REG2_REG_13__SCAN_IN), .B2(n9297), .A(n9296), .ZN(
        n9307) );
  AOI21_X1 U10349 ( .B1(n10495), .B2(P2_ADDR_REG_13__SCAN_IN), .A(n9298), .ZN(
        n9304) );
  OAI21_X1 U10350 ( .B1(n9301), .B2(n9300), .A(n9299), .ZN(n9302) );
  NAND2_X1 U10351 ( .A1(n9302), .A2(n10504), .ZN(n9303) );
  OAI211_X1 U10352 ( .C1(n10403), .C2(n9305), .A(n9304), .B(n9303), .ZN(n9306)
         );
  AOI21_X1 U10353 ( .B1(n9307), .B2(n10505), .A(n9306), .ZN(n9308) );
  OAI21_X1 U10354 ( .B1(n9309), .B2(n10511), .A(n9308), .ZN(P2_U3195) );
  AOI21_X1 U10355 ( .B1(n5016), .B2(n9311), .A(n9310), .ZN(n9326) );
  OAI21_X1 U10356 ( .B1(n9314), .B2(n9313), .A(n9312), .ZN(n9324) );
  AOI21_X1 U10357 ( .B1(n10495), .B2(P2_ADDR_REG_14__SCAN_IN), .A(n9315), .ZN(
        n9321) );
  OAI21_X1 U10358 ( .B1(n9318), .B2(n9317), .A(n9316), .ZN(n9319) );
  NAND2_X1 U10359 ( .A1(n9319), .A2(n10504), .ZN(n9320) );
  OAI211_X1 U10360 ( .C1(n10403), .C2(n9322), .A(n9321), .B(n9320), .ZN(n9323)
         );
  AOI21_X1 U10361 ( .B1(n9324), .B2(n10505), .A(n9323), .ZN(n9325) );
  OAI21_X1 U10362 ( .B1(n9326), .B2(n10511), .A(n9325), .ZN(P2_U3196) );
  AOI21_X1 U10363 ( .B1(n9329), .B2(n9328), .A(n9327), .ZN(n9342) );
  OAI21_X1 U10364 ( .B1(P2_REG2_REG_15__SCAN_IN), .B2(n9331), .A(n9330), .ZN(
        n9340) );
  AOI21_X1 U10365 ( .B1(n10495), .B2(P2_ADDR_REG_15__SCAN_IN), .A(n9332), .ZN(
        n9338) );
  OAI21_X1 U10366 ( .B1(n9335), .B2(n9334), .A(n9333), .ZN(n9336) );
  NAND2_X1 U10367 ( .A1(n9336), .A2(n10504), .ZN(n9337) );
  OAI211_X1 U10368 ( .C1(n10403), .C2(n5104), .A(n9338), .B(n9337), .ZN(n9339)
         );
  AOI21_X1 U10369 ( .B1(n9340), .B2(n10505), .A(n9339), .ZN(n9341) );
  OAI21_X1 U10370 ( .B1(n9342), .B2(n10511), .A(n9341), .ZN(P2_U3197) );
  AOI21_X1 U10371 ( .B1(n9345), .B2(n9344), .A(n9343), .ZN(n9360) );
  OAI21_X1 U10372 ( .B1(n9348), .B2(n9347), .A(n9346), .ZN(n9358) );
  AOI21_X1 U10373 ( .B1(n10495), .B2(P2_ADDR_REG_16__SCAN_IN), .A(n9349), .ZN(
        n9355) );
  OAI21_X1 U10374 ( .B1(n9352), .B2(n9351), .A(n9350), .ZN(n9353) );
  NAND2_X1 U10375 ( .A1(n9353), .A2(n10504), .ZN(n9354) );
  OAI211_X1 U10376 ( .C1(n10403), .C2(n9356), .A(n9355), .B(n9354), .ZN(n9357)
         );
  AOI21_X1 U10377 ( .B1(n9358), .B2(n10505), .A(n9357), .ZN(n9359) );
  OAI21_X1 U10378 ( .B1(n9360), .B2(n10511), .A(n9359), .ZN(P2_U3198) );
  AOI21_X1 U10379 ( .B1(n9363), .B2(n9362), .A(n9361), .ZN(n9377) );
  OAI21_X1 U10380 ( .B1(P2_REG2_REG_17__SCAN_IN), .B2(n9365), .A(n9364), .ZN(
        n9375) );
  OAI21_X1 U10381 ( .B1(n9368), .B2(n9367), .A(n9366), .ZN(n9369) );
  NAND2_X1 U10382 ( .A1(n9369), .A2(n10504), .ZN(n9372) );
  AOI21_X1 U10383 ( .B1(n10495), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n9370), .ZN(
        n9371) );
  OAI211_X1 U10384 ( .C1(n10403), .C2(n9373), .A(n9372), .B(n9371), .ZN(n9374)
         );
  AOI21_X1 U10385 ( .B1(n9375), .B2(n10505), .A(n9374), .ZN(n9376) );
  OAI21_X1 U10386 ( .B1(n9377), .B2(n10511), .A(n9376), .ZN(P2_U3199) );
  AOI21_X1 U10387 ( .B1(n4982), .B2(n9379), .A(n9378), .ZN(n9396) );
  XNOR2_X1 U10388 ( .A(n9391), .B(n9380), .ZN(n9381) );
  XNOR2_X1 U10389 ( .A(n9382), .B(n9381), .ZN(n9394) );
  INV_X1 U10390 ( .A(n9383), .ZN(n9384) );
  NOR2_X1 U10391 ( .A1(n9385), .A2(n9384), .ZN(n9387) );
  AOI21_X1 U10392 ( .B1(n9387), .B2(P2_U3893), .A(n10497), .ZN(n9392) );
  AOI21_X1 U10393 ( .B1(n10495), .B2(P2_ADDR_REG_18__SCAN_IN), .A(n9386), .ZN(
        n9390) );
  INV_X1 U10394 ( .A(n9387), .ZN(n9388) );
  NAND3_X1 U10395 ( .A1(n9388), .A2(n10504), .A3(n9391), .ZN(n9389) );
  OAI211_X1 U10396 ( .C1(n9392), .C2(n9391), .A(n9390), .B(n9389), .ZN(n9393)
         );
  AOI21_X1 U10397 ( .B1(n9394), .B2(n10505), .A(n9393), .ZN(n9395) );
  OAI21_X1 U10398 ( .B1(n9396), .B2(n10511), .A(n9395), .ZN(P2_U3200) );
  INV_X1 U10399 ( .A(n9397), .ZN(n9399) );
  NOR2_X1 U10400 ( .A1(n9399), .A2(n9398), .ZN(n9628) );
  NOR3_X1 U10401 ( .A1(n9628), .A2(n10687), .A3(n9400), .ZN(n9403) );
  NOR2_X1 U10402 ( .A1(n10641), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n9401) );
  OAI22_X1 U10403 ( .A1(n9630), .A2(n9509), .B1(n9403), .B2(n9401), .ZN(
        P2_U3202) );
  NOR2_X1 U10404 ( .A1(n10641), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n9402) );
  OAI22_X1 U10405 ( .A1(n9633), .A2(n9509), .B1(n9403), .B2(n9402), .ZN(
        P2_U3203) );
  XNOR2_X1 U10406 ( .A(n9404), .B(n9412), .ZN(n9405) );
  AOI22_X1 U10407 ( .A1(n9405), .A2(n9532), .B1(n9534), .B2(n9563), .ZN(n9557)
         );
  AOI22_X1 U10408 ( .A1(n9406), .A2(n10634), .B1(n10687), .B2(
        P2_REG2_REG_27__SCAN_IN), .ZN(n9407) );
  OAI21_X1 U10409 ( .B1(n9408), .B2(n9545), .A(n9407), .ZN(n9414) );
  NAND2_X1 U10410 ( .A1(n9410), .A2(n9409), .ZN(n9411) );
  XOR2_X1 U10411 ( .A(n9412), .B(n9411), .Z(n9558) );
  NOR2_X1 U10412 ( .A1(n9558), .A2(n9493), .ZN(n9413) );
  AOI211_X1 U10413 ( .C1(n10636), .C2(n9555), .A(n9414), .B(n9413), .ZN(n9415)
         );
  OAI21_X1 U10414 ( .B1(n9557), .B2(n10687), .A(n9415), .ZN(P2_U3206) );
  XNOR2_X1 U10415 ( .A(n9417), .B(n9416), .ZN(n9418) );
  OAI222_X1 U10416 ( .A1(n9515), .A2(n9438), .B1(n9616), .B2(n6814), .C1(n9498), .C2(n9418), .ZN(n9559) );
  INV_X1 U10417 ( .A(n9559), .ZN(n9424) );
  XNOR2_X1 U10418 ( .A(n6912), .B(n9419), .ZN(n9560) );
  AOI22_X1 U10419 ( .A1(n9420), .A2(n10634), .B1(n10687), .B2(
        P2_REG2_REG_26__SCAN_IN), .ZN(n9421) );
  OAI21_X1 U10420 ( .B1(n9638), .B2(n9509), .A(n9421), .ZN(n9422) );
  AOI21_X1 U10421 ( .B1(n9560), .B2(n9547), .A(n9422), .ZN(n9423) );
  OAI21_X1 U10422 ( .B1(n9424), .B2(n10687), .A(n9423), .ZN(P2_U3207) );
  XNOR2_X1 U10423 ( .A(n9425), .B(n9426), .ZN(n9567) );
  XNOR2_X1 U10424 ( .A(n9427), .B(n9426), .ZN(n9428) );
  AOI22_X1 U10425 ( .A1(n9428), .A2(n9532), .B1(n9534), .B2(n9446), .ZN(n9566)
         );
  INV_X1 U10426 ( .A(n9566), .ZN(n9433) );
  INV_X1 U10427 ( .A(n9429), .ZN(n9430) );
  OAI22_X1 U10428 ( .A1(n9431), .A2(n10585), .B1(n9430), .B2(n10677), .ZN(
        n9432) );
  OAI21_X1 U10429 ( .B1(n9433), .B2(n9432), .A(n10641), .ZN(n9435) );
  AOI22_X1 U10430 ( .A1(n9563), .A2(n9470), .B1(n10687), .B2(
        P2_REG2_REG_25__SCAN_IN), .ZN(n9434) );
  OAI211_X1 U10431 ( .C1(n9567), .C2(n9493), .A(n9435), .B(n9434), .ZN(
        P2_U3208) );
  NOR2_X1 U10432 ( .A1(n9643), .A2(n10585), .ZN(n9439) );
  XOR2_X1 U10433 ( .A(n9441), .B(n9436), .Z(n9437) );
  OAI222_X1 U10434 ( .A1(n9616), .A2(n9438), .B1(n9515), .B2(n9459), .C1(n9498), .C2(n9437), .ZN(n9568) );
  AOI211_X1 U10435 ( .C1(n10634), .C2(n9440), .A(n9439), .B(n9568), .ZN(n9443)
         );
  XNOR2_X1 U10436 ( .A(n5003), .B(n9441), .ZN(n9569) );
  AOI22_X1 U10437 ( .A1(n9569), .A2(n9547), .B1(P2_REG2_REG_24__SCAN_IN), .B2(
        n10687), .ZN(n9442) );
  OAI21_X1 U10438 ( .B1(n9443), .B2(n10687), .A(n9442), .ZN(P2_U3209) );
  XNOR2_X1 U10439 ( .A(n9445), .B(n9444), .ZN(n9447) );
  AOI222_X1 U10440 ( .A1(n9532), .A2(n9447), .B1(n9446), .B2(n9609), .C1(n9580), .C2(n9534), .ZN(n9574) );
  INV_X1 U10441 ( .A(n9448), .ZN(n9450) );
  OAI22_X1 U10442 ( .A1(n9450), .A2(n10677), .B1(n10641), .B2(n9449), .ZN(
        n9455) );
  AOI21_X1 U10443 ( .B1(n9453), .B2(n9452), .A(n9451), .ZN(n9575) );
  NOR2_X1 U10444 ( .A1(n9575), .A2(n9493), .ZN(n9454) );
  AOI211_X1 U10445 ( .C1(n10636), .C2(n9572), .A(n9455), .B(n9454), .ZN(n9456)
         );
  OAI21_X1 U10446 ( .B1(n9574), .B2(n10687), .A(n9456), .ZN(P2_U3210) );
  XNOR2_X1 U10447 ( .A(n9457), .B(n9460), .ZN(n9458) );
  OAI222_X1 U10448 ( .A1(n9616), .A2(n9459), .B1(n9515), .B2(n9488), .C1(n9458), .C2(n9498), .ZN(n9576) );
  INV_X1 U10449 ( .A(n9576), .ZN(n9466) );
  XOR2_X1 U10450 ( .A(n9461), .B(n9460), .Z(n9577) );
  AOI22_X1 U10451 ( .A1(n10687), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n9462), 
        .B2(n10634), .ZN(n9463) );
  OAI21_X1 U10452 ( .B1(n9648), .B2(n9509), .A(n9463), .ZN(n9464) );
  AOI21_X1 U10453 ( .B1(n9577), .B2(n9547), .A(n9464), .ZN(n9465) );
  OAI21_X1 U10454 ( .B1(n9466), .B2(n10687), .A(n9465), .ZN(P2_U3211) );
  XNOR2_X1 U10455 ( .A(n9467), .B(n9478), .ZN(n9469) );
  AOI22_X1 U10456 ( .A1(n9469), .A2(n9532), .B1(n9534), .B2(n9468), .ZN(n9583)
         );
  NAND2_X1 U10457 ( .A1(n9580), .A2(n9470), .ZN(n9473) );
  NAND2_X1 U10458 ( .A1(n9471), .A2(n10634), .ZN(n9472) );
  OAI211_X1 U10459 ( .C1(n10641), .C2(n9474), .A(n9473), .B(n9472), .ZN(n9475)
         );
  AOI21_X1 U10460 ( .B1(n9581), .B2(n10636), .A(n9475), .ZN(n9481) );
  OR2_X1 U10461 ( .A1(n9491), .A2(n9492), .ZN(n9489) );
  AND2_X1 U10462 ( .A1(n9489), .A2(n9476), .ZN(n9479) );
  OAI21_X1 U10463 ( .B1(n9479), .B2(n9478), .A(n9477), .ZN(n9584) );
  OR2_X1 U10464 ( .A1(n9584), .A2(n9493), .ZN(n9480) );
  OAI211_X1 U10465 ( .C1(n9583), .C2(n10687), .A(n9481), .B(n9480), .ZN(
        P2_U3212) );
  OAI21_X1 U10466 ( .B1(n9492), .B2(n9483), .A(n9482), .ZN(n9485) );
  AOI22_X1 U10467 ( .A1(n9485), .A2(n9532), .B1(n9534), .B2(n9484), .ZN(n9588)
         );
  AOI22_X1 U10468 ( .A1(n10687), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n10634), 
        .B2(n9486), .ZN(n9487) );
  OAI21_X1 U10469 ( .B1(n9488), .B2(n9545), .A(n9487), .ZN(n9495) );
  INV_X1 U10470 ( .A(n9489), .ZN(n9490) );
  AOI21_X1 U10471 ( .B1(n9492), .B2(n9491), .A(n9490), .ZN(n9589) );
  NOR2_X1 U10472 ( .A1(n9589), .A2(n9493), .ZN(n9494) );
  AOI211_X1 U10473 ( .C1(n10636), .C2(n9586), .A(n9495), .B(n9494), .ZN(n9496)
         );
  OAI21_X1 U10474 ( .B1(n10687), .B2(n9588), .A(n9496), .ZN(P2_U3213) );
  AOI211_X1 U10475 ( .C1(n9504), .C2(n9499), .A(n9498), .B(n9497), .ZN(n9502)
         );
  OAI22_X1 U10476 ( .A1(n9500), .A2(n9616), .B1(n9604), .B2(n9515), .ZN(n9501)
         );
  OR2_X1 U10477 ( .A1(n9502), .A2(n9501), .ZN(n9590) );
  INV_X1 U10478 ( .A(n9590), .ZN(n9512) );
  OAI21_X1 U10479 ( .B1(n9505), .B2(n9504), .A(n9503), .ZN(n9506) );
  INV_X1 U10480 ( .A(n9506), .ZN(n9591) );
  AOI22_X1 U10481 ( .A1(n10687), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n10634), 
        .B2(n9507), .ZN(n9508) );
  OAI21_X1 U10482 ( .B1(n9655), .B2(n9509), .A(n9508), .ZN(n9510) );
  AOI21_X1 U10483 ( .B1(n9591), .B2(n9547), .A(n9510), .ZN(n9511) );
  OAI21_X1 U10484 ( .B1(n9512), .B2(n10687), .A(n9511), .ZN(P2_U3214) );
  XNOR2_X1 U10485 ( .A(n9513), .B(n9525), .ZN(n9514) );
  NAND2_X1 U10486 ( .A1(n9514), .A2(n9532), .ZN(n9520) );
  OAI22_X1 U10487 ( .A1(n9517), .A2(n9616), .B1(n9516), .B2(n9515), .ZN(n9518)
         );
  INV_X1 U10488 ( .A(n9518), .ZN(n9519) );
  NAND2_X1 U10489 ( .A1(n9520), .A2(n9519), .ZN(n9600) );
  INV_X1 U10490 ( .A(n9600), .ZN(n9529) );
  INV_X1 U10491 ( .A(n9521), .ZN(n9522) );
  OAI22_X1 U10492 ( .A1(n10641), .A2(n9380), .B1(n9522), .B2(n10677), .ZN(
        n9523) );
  AOI21_X1 U10493 ( .B1(n9524), .B2(n10636), .A(n9523), .ZN(n9528) );
  NAND2_X1 U10494 ( .A1(n9526), .A2(n9525), .ZN(n9595) );
  NAND3_X1 U10495 ( .A1(n9596), .A2(n9595), .A3(n9547), .ZN(n9527) );
  OAI211_X1 U10496 ( .C1(n9529), .C2(n10687), .A(n9528), .B(n9527), .ZN(
        P2_U3215) );
  INV_X1 U10497 ( .A(n9538), .ZN(n9531) );
  XNOR2_X1 U10498 ( .A(n9530), .B(n9531), .ZN(n9533) );
  NAND2_X1 U10499 ( .A1(n9533), .A2(n9532), .ZN(n9537) );
  NAND2_X1 U10500 ( .A1(n9535), .A2(n9534), .ZN(n9536) );
  NAND2_X1 U10501 ( .A1(n9537), .A2(n9536), .ZN(n9606) );
  INV_X1 U10502 ( .A(n9606), .ZN(n9549) );
  NAND2_X1 U10503 ( .A1(n9539), .A2(n9538), .ZN(n9540) );
  NAND2_X1 U10504 ( .A1(n9541), .A2(n9540), .ZN(n9601) );
  NAND2_X1 U10505 ( .A1(n9602), .A2(n10636), .ZN(n9544) );
  AOI22_X1 U10506 ( .A1(n10687), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n10634), 
        .B2(n9542), .ZN(n9543) );
  OAI211_X1 U10507 ( .C1(n9604), .C2(n9545), .A(n9544), .B(n9543), .ZN(n9546)
         );
  AOI21_X1 U10508 ( .B1(n9601), .B2(n9547), .A(n9546), .ZN(n9548) );
  OAI21_X1 U10509 ( .B1(n9549), .B2(n10687), .A(n9548), .ZN(P2_U3216) );
  NAND2_X1 U10510 ( .A1(n9628), .A2(n9627), .ZN(n9551) );
  NAND2_X1 U10511 ( .A1(n9624), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n9550) );
  OAI211_X1 U10512 ( .C1(n9630), .C2(n9594), .A(n9551), .B(n9550), .ZN(
        P2_U3490) );
  NAND2_X1 U10513 ( .A1(n9624), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n9552) );
  OAI211_X1 U10514 ( .C1(n9633), .C2(n9594), .A(n9552), .B(n9551), .ZN(
        P2_U3489) );
  MUX2_X1 U10515 ( .A(n9553), .B(P2_REG1_REG_29__SCAN_IN), .S(n9624), .Z(
        P2_U3488) );
  AOI22_X1 U10516 ( .A1(n9555), .A2(n9610), .B1(n9609), .B2(n9554), .ZN(n9556)
         );
  OAI211_X1 U10517 ( .C1(n9615), .C2(n9558), .A(n9557), .B(n9556), .ZN(n9634)
         );
  MUX2_X1 U10518 ( .A(n9634), .B(P2_REG1_REG_27__SCAN_IN), .S(n9624), .Z(
        P2_U3486) );
  AOI21_X1 U10519 ( .B1(n9560), .B2(n9623), .A(n9559), .ZN(n9635) );
  INV_X1 U10520 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n9561) );
  MUX2_X1 U10521 ( .A(n9635), .B(n9561), .S(n9624), .Z(n9562) );
  OAI21_X1 U10522 ( .B1(n9638), .B2(n9594), .A(n9562), .ZN(P2_U3485) );
  AOI22_X1 U10523 ( .A1(n9564), .A2(n9610), .B1(n9609), .B2(n9563), .ZN(n9565)
         );
  OAI211_X1 U10524 ( .C1(n9615), .C2(n9567), .A(n9566), .B(n9565), .ZN(n9639)
         );
  MUX2_X1 U10525 ( .A(n9639), .B(P2_REG1_REG_25__SCAN_IN), .S(n9624), .Z(
        P2_U3484) );
  AOI21_X1 U10526 ( .B1(n9569), .B2(n9623), .A(n9568), .ZN(n9640) );
  INV_X1 U10527 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n9570) );
  MUX2_X1 U10528 ( .A(n9640), .B(n9570), .S(n9624), .Z(n9571) );
  OAI21_X1 U10529 ( .B1(n9643), .B2(n9594), .A(n9571), .ZN(P2_U3483) );
  NAND2_X1 U10530 ( .A1(n9572), .A2(n9610), .ZN(n9573) );
  OAI211_X1 U10531 ( .C1(n9615), .C2(n9575), .A(n9574), .B(n9573), .ZN(n9644)
         );
  MUX2_X1 U10532 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n9644), .S(n9627), .Z(
        P2_U3482) );
  INV_X1 U10533 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n9578) );
  AOI21_X1 U10534 ( .B1(n9577), .B2(n9623), .A(n9576), .ZN(n9645) );
  MUX2_X1 U10535 ( .A(n9578), .B(n9645), .S(n9627), .Z(n9579) );
  OAI21_X1 U10536 ( .B1(n9648), .B2(n9594), .A(n9579), .ZN(P2_U3481) );
  AOI22_X1 U10537 ( .A1(n9581), .A2(n9610), .B1(n9609), .B2(n9580), .ZN(n9582)
         );
  OAI211_X1 U10538 ( .C1(n9615), .C2(n9584), .A(n9583), .B(n9582), .ZN(n9649)
         );
  MUX2_X1 U10539 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n9649), .S(n9627), .Z(
        P2_U3480) );
  AOI22_X1 U10540 ( .A1(n9586), .A2(n9610), .B1(n9609), .B2(n9585), .ZN(n9587)
         );
  OAI211_X1 U10541 ( .C1(n9615), .C2(n9589), .A(n9588), .B(n9587), .ZN(n9650)
         );
  MUX2_X1 U10542 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n9650), .S(n9627), .Z(
        P2_U3479) );
  INV_X1 U10543 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n9592) );
  AOI21_X1 U10544 ( .B1(n9591), .B2(n9623), .A(n9590), .ZN(n9651) );
  MUX2_X1 U10545 ( .A(n9592), .B(n9651), .S(n9627), .Z(n9593) );
  OAI21_X1 U10546 ( .B1(n9655), .B2(n9594), .A(n9593), .ZN(P2_U3478) );
  NAND3_X1 U10547 ( .A1(n9596), .A2(n9595), .A3(n9623), .ZN(n9597) );
  OAI21_X1 U10548 ( .B1(n9598), .B2(n9618), .A(n9597), .ZN(n9599) );
  MUX2_X1 U10549 ( .A(n9656), .B(P2_REG1_REG_18__SCAN_IN), .S(n9624), .Z(
        P2_U3477) );
  AND2_X1 U10550 ( .A1(n9601), .A2(n9623), .ZN(n9607) );
  NAND2_X1 U10551 ( .A1(n9602), .A2(n9610), .ZN(n9603) );
  OAI21_X1 U10552 ( .B1(n9604), .B2(n9616), .A(n9603), .ZN(n9605) );
  MUX2_X1 U10553 ( .A(n9657), .B(P2_REG1_REG_17__SCAN_IN), .S(n9624), .Z(
        P2_U3476) );
  AOI22_X1 U10554 ( .A1(n9611), .A2(n9610), .B1(n9609), .B2(n9608), .ZN(n9612)
         );
  OAI211_X1 U10555 ( .C1(n9615), .C2(n9614), .A(n9613), .B(n9612), .ZN(n9658)
         );
  MUX2_X1 U10556 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n9658), .S(n9627), .Z(
        P2_U3475) );
  OAI22_X1 U10557 ( .A1(n9619), .A2(n9618), .B1(n9617), .B2(n9616), .ZN(n9621)
         );
  AOI211_X1 U10558 ( .C1(n9623), .C2(n9622), .A(n9621), .B(n9620), .ZN(n10691)
         );
  OR2_X1 U10559 ( .A1(n10691), .A2(n9624), .ZN(n9625) );
  OAI21_X1 U10560 ( .B1(n9627), .B2(n9626), .A(n9625), .ZN(P2_U3473) );
  NAND2_X1 U10561 ( .A1(n10692), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n9629) );
  NAND2_X1 U10562 ( .A1(n9628), .A2(n10695), .ZN(n9631) );
  OAI211_X1 U10563 ( .C1(n9630), .C2(n9654), .A(n9629), .B(n9631), .ZN(
        P2_U3458) );
  NAND2_X1 U10564 ( .A1(n10692), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n9632) );
  OAI211_X1 U10565 ( .C1(n9633), .C2(n9654), .A(n9632), .B(n9631), .ZN(
        P2_U3457) );
  MUX2_X1 U10566 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n9634), .S(n10695), .Z(
        P2_U3454) );
  INV_X1 U10567 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n9636) );
  MUX2_X1 U10568 ( .A(n9636), .B(n9635), .S(n10695), .Z(n9637) );
  OAI21_X1 U10569 ( .B1(n9638), .B2(n9654), .A(n9637), .ZN(P2_U3453) );
  MUX2_X1 U10570 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n9639), .S(n10695), .Z(
        P2_U3452) );
  INV_X1 U10571 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n9641) );
  MUX2_X1 U10572 ( .A(n9641), .B(n9640), .S(n10695), .Z(n9642) );
  OAI21_X1 U10573 ( .B1(n9643), .B2(n9654), .A(n9642), .ZN(P2_U3451) );
  MUX2_X1 U10574 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n9644), .S(n10695), .Z(
        P2_U3450) );
  INV_X1 U10575 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n9646) );
  MUX2_X1 U10576 ( .A(n9646), .B(n9645), .S(n10695), .Z(n9647) );
  OAI21_X1 U10577 ( .B1(n9648), .B2(n9654), .A(n9647), .ZN(P2_U3449) );
  MUX2_X1 U10578 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n9649), .S(n10695), .Z(
        P2_U3448) );
  MUX2_X1 U10579 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n9650), .S(n10695), .Z(
        P2_U3447) );
  INV_X1 U10580 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n9652) );
  MUX2_X1 U10581 ( .A(n9652), .B(n9651), .S(n10695), .Z(n9653) );
  OAI21_X1 U10582 ( .B1(n9655), .B2(n9654), .A(n9653), .ZN(P2_U3446) );
  MUX2_X1 U10583 ( .A(n9656), .B(P2_REG0_REG_18__SCAN_IN), .S(n10692), .Z(
        P2_U3444) );
  MUX2_X1 U10584 ( .A(n9657), .B(P2_REG0_REG_17__SCAN_IN), .S(n10692), .Z(
        P2_U3441) );
  MUX2_X1 U10585 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n9658), .S(n10695), .Z(
        P2_U3438) );
  MUX2_X1 U10586 ( .A(P2_D_REG_1__SCAN_IN), .B(n9660), .S(n9659), .Z(P2_U3377)
         );
  INV_X1 U10587 ( .A(n8847), .ZN(n10279) );
  NOR4_X1 U10588 ( .A1(n6483), .A2(P2_IR_REG_30__SCAN_IN), .A3(P2_U3151), .A4(
        n6609), .ZN(n9661) );
  AOI21_X1 U10589 ( .B1(P1_DATAO_REG_31__SCAN_IN), .B2(n9674), .A(n9661), .ZN(
        n9662) );
  OAI21_X1 U10590 ( .B1(n10279), .B2(n9676), .A(n9662), .ZN(P2_U3264) );
  INV_X1 U10591 ( .A(n9663), .ZN(n10282) );
  AOI22_X1 U10592 ( .A1(n9664), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n9674), .ZN(n9665) );
  OAI21_X1 U10593 ( .B1(n10282), .B2(n9676), .A(n9665), .ZN(P2_U3265) );
  INV_X1 U10594 ( .A(n9666), .ZN(n10285) );
  AOI22_X1 U10595 ( .A1(n9667), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_29__SCAN_IN), .B2(n9674), .ZN(n9668) );
  OAI21_X1 U10596 ( .B1(n10285), .B2(n9676), .A(n9668), .ZN(P2_U3266) );
  INV_X1 U10597 ( .A(n9669), .ZN(n10289) );
  AOI21_X1 U10598 ( .B1(P1_DATAO_REG_28__SCAN_IN), .B2(n9674), .A(n9670), .ZN(
        n9671) );
  OAI21_X1 U10599 ( .B1(n10289), .B2(n9676), .A(n9671), .ZN(P2_U3267) );
  INV_X1 U10600 ( .A(n9672), .ZN(n10292) );
  AOI21_X1 U10601 ( .B1(P1_DATAO_REG_27__SCAN_IN), .B2(n9674), .A(n9673), .ZN(
        n9675) );
  OAI21_X1 U10602 ( .B1(n10292), .B2(n9676), .A(n9675), .ZN(P2_U3268) );
  MUX2_X1 U10603 ( .A(n9677), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  XOR2_X1 U10604 ( .A(n9679), .B(n9678), .Z(n9685) );
  OAI22_X1 U10605 ( .A1(n9775), .A2(n10031), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9680), .ZN(n9683) );
  INV_X1 U10606 ( .A(n10034), .ZN(n9681) );
  OAI22_X1 U10607 ( .A1(n9756), .A2(n9681), .B1(n9754), .B2(n10065), .ZN(n9682) );
  AOI211_X1 U10608 ( .C1(n6101), .C2(n9789), .A(n9683), .B(n9682), .ZN(n9684)
         );
  OAI21_X1 U10609 ( .B1(n9685), .B2(n9778), .A(n9684), .ZN(P1_U3216) );
  INV_X1 U10610 ( .A(n9687), .ZN(n9688) );
  AOI21_X1 U10611 ( .B1(n9689), .B2(n9686), .A(n9688), .ZN(n9693) );
  NAND2_X1 U10612 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9919) );
  OAI21_X1 U10613 ( .B1(n9775), .B2(n10097), .A(n9919), .ZN(n9691) );
  OAI22_X1 U10614 ( .A1(n10099), .A2(n9756), .B1(n9754), .B2(n10124), .ZN(
        n9690) );
  AOI211_X1 U10615 ( .C1(n10102), .C2(n9789), .A(n9691), .B(n9690), .ZN(n9692)
         );
  OAI21_X1 U10616 ( .B1(n9693), .B2(n9778), .A(n9692), .ZN(P1_U3219) );
  AOI21_X1 U10617 ( .B1(n9694), .B2(n9695), .A(n9778), .ZN(n9697) );
  NAND2_X1 U10618 ( .A1(n9697), .A2(n9696), .ZN(n9702) );
  AOI22_X1 U10619 ( .A1(n9787), .A2(n9798), .B1(P1_REG3_REG_21__SCAN_IN), .B2(
        P1_U3086), .ZN(n9701) );
  AOI22_X1 U10620 ( .A1(n10071), .A2(n9788), .B1(n9786), .B2(n9698), .ZN(n9700) );
  NAND2_X1 U10621 ( .A1(n10070), .A2(n9789), .ZN(n9699) );
  NAND4_X1 U10622 ( .A1(n9702), .A2(n9701), .A3(n9700), .A4(n9699), .ZN(
        P1_U3223) );
  AOI21_X1 U10623 ( .B1(n9704), .B2(n9703), .A(n4981), .ZN(n9705) );
  OR2_X1 U10624 ( .A1(n9705), .A2(n9778), .ZN(n9710) );
  AOI22_X1 U10625 ( .A1(n9787), .A2(n9797), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3086), .ZN(n9709) );
  AOI22_X1 U10626 ( .A1(n10003), .A2(n9788), .B1(n9786), .B2(n9706), .ZN(n9708) );
  NAND2_X1 U10627 ( .A1(n10174), .A2(n9789), .ZN(n9707) );
  NAND4_X1 U10628 ( .A1(n9710), .A2(n9709), .A3(n9708), .A4(n9707), .ZN(
        P1_U3225) );
  INV_X1 U10629 ( .A(n9712), .ZN(n9713) );
  AOI21_X1 U10630 ( .B1(n9714), .B2(n9711), .A(n9713), .ZN(n9718) );
  AOI22_X1 U10631 ( .A1(n10148), .A2(n9788), .B1(n9786), .B2(n9800), .ZN(n9715) );
  NAND2_X1 U10632 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9862) );
  OAI211_X1 U10633 ( .C1(n10144), .C2(n9775), .A(n9715), .B(n9862), .ZN(n9716)
         );
  AOI21_X1 U10634 ( .B1(n10222), .B2(n9789), .A(n9716), .ZN(n9717) );
  OAI21_X1 U10635 ( .B1(n9718), .B2(n9778), .A(n9717), .ZN(P1_U3226) );
  AOI21_X1 U10636 ( .B1(n9720), .B2(n9722), .A(n9719), .ZN(n9721) );
  AOI21_X1 U10637 ( .B1(n5015), .B2(n9722), .A(n9721), .ZN(n9727) );
  AOI22_X1 U10638 ( .A1(n9788), .A2(n10130), .B1(n9786), .B2(n9723), .ZN(n9724) );
  NAND2_X1 U10639 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9885) );
  OAI211_X1 U10640 ( .C1(n10124), .C2(n9775), .A(n9724), .B(n9885), .ZN(n9725)
         );
  AOI21_X1 U10641 ( .B1(n10131), .B2(n9789), .A(n9725), .ZN(n9726) );
  OAI21_X1 U10642 ( .B1(n9727), .B2(n9778), .A(n9726), .ZN(P1_U3228) );
  NAND2_X1 U10643 ( .A1(n5012), .A2(n9728), .ZN(n9729) );
  XNOR2_X1 U10644 ( .A(n9730), .B(n9729), .ZN(n9737) );
  OAI22_X1 U10645 ( .A1(n9775), .A2(n9732), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9731), .ZN(n9735) );
  INV_X1 U10646 ( .A(n10019), .ZN(n9733) );
  OAI22_X1 U10647 ( .A1(n9733), .A2(n9756), .B1(n9754), .B2(n9753), .ZN(n9734)
         );
  AOI211_X1 U10648 ( .C1(n10181), .C2(n9789), .A(n9735), .B(n9734), .ZN(n9736)
         );
  OAI21_X1 U10649 ( .B1(n9737), .B2(n9778), .A(n9736), .ZN(P1_U3229) );
  XOR2_X1 U10650 ( .A(n9738), .B(n9739), .Z(n9745) );
  OAI22_X1 U10651 ( .A1(n9775), .A2(n10081), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9740), .ZN(n9743) );
  INV_X1 U10652 ( .A(n10084), .ZN(n9741) );
  OAI22_X1 U10653 ( .A1(n9741), .A2(n9756), .B1(n9754), .B2(n10111), .ZN(n9742) );
  AOI211_X1 U10654 ( .C1(n10200), .C2(n9789), .A(n9743), .B(n9742), .ZN(n9744)
         );
  OAI21_X1 U10655 ( .B1(n9745), .B2(n9778), .A(n9744), .ZN(P1_U3233) );
  INV_X1 U10656 ( .A(n9746), .ZN(n9750) );
  AOI21_X1 U10657 ( .B1(n9750), .B2(n9748), .A(n9747), .ZN(n9749) );
  AOI21_X1 U10658 ( .B1(n9751), .B2(n9750), .A(n9749), .ZN(n9760) );
  OAI22_X1 U10659 ( .A1(n9775), .A2(n9753), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9752), .ZN(n9758) );
  INV_X1 U10660 ( .A(n10053), .ZN(n9755) );
  OAI22_X1 U10661 ( .A1(n9756), .A2(n9755), .B1(n9754), .B2(n10081), .ZN(n9757) );
  AOI211_X1 U10662 ( .C1(n10190), .C2(n9789), .A(n9758), .B(n9757), .ZN(n9759)
         );
  OAI21_X1 U10663 ( .B1(n9760), .B2(n9778), .A(n9759), .ZN(P1_U3235) );
  OAI21_X1 U10664 ( .B1(n9761), .B2(n9763), .A(n9762), .ZN(n9764) );
  NAND2_X1 U10665 ( .A1(n9764), .A2(n9784), .ZN(n9768) );
  AOI22_X1 U10666 ( .A1(n9786), .A2(n6960), .B1(n9787), .B2(n10559), .ZN(n9767) );
  AOI22_X1 U10667 ( .A1(n10571), .A2(n9789), .B1(n9765), .B2(
        P1_REG3_REG_2__SCAN_IN), .ZN(n9766) );
  NAND3_X1 U10668 ( .A1(n9768), .A2(n9767), .A3(n9766), .ZN(P1_U3237) );
  NAND2_X1 U10669 ( .A1(n9770), .A2(n9769), .ZN(n9771) );
  XOR2_X1 U10670 ( .A(n9772), .B(n9771), .Z(n9779) );
  AOI22_X1 U10671 ( .A1(n10114), .A2(n9788), .B1(n9786), .B2(n9773), .ZN(n9774) );
  NAND2_X1 U10672 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9902) );
  OAI211_X1 U10673 ( .C1(n10111), .C2(n9775), .A(n9774), .B(n9902), .ZN(n9776)
         );
  AOI21_X1 U10674 ( .B1(n10210), .B2(n9789), .A(n9776), .ZN(n9777) );
  OAI21_X1 U10675 ( .B1(n9779), .B2(n9778), .A(n9777), .ZN(P1_U3238) );
  OAI21_X1 U10676 ( .B1(n4981), .B2(n9782), .A(n9781), .ZN(n9783) );
  NAND3_X1 U10677 ( .A1(n9785), .A2(n9784), .A3(n9783), .ZN(n9793) );
  AOI22_X1 U10678 ( .A1(n9786), .A2(n10015), .B1(P1_REG3_REG_26__SCAN_IN), 
        .B2(P1_U3086), .ZN(n9792) );
  AOI22_X1 U10679 ( .A1(n9788), .A2(n9977), .B1(n9787), .B2(n9796), .ZN(n9791)
         );
  NAND2_X1 U10680 ( .A1(n10249), .A2(n9789), .ZN(n9790) );
  NAND4_X1 U10681 ( .A1(n9793), .A2(n9792), .A3(n9791), .A4(n9790), .ZN(
        P1_U3240) );
  MUX2_X1 U10682 ( .A(n5408), .B(P1_DATAO_REG_31__SCAN_IN), .S(n9825), .Z(
        P1_U3585) );
  MUX2_X1 U10683 ( .A(n9794), .B(P1_DATAO_REG_30__SCAN_IN), .S(n9825), .Z(
        P1_U3584) );
  MUX2_X1 U10684 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9795), .S(P1_U3973), .Z(
        P1_U3582) );
  MUX2_X1 U10685 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9796), .S(P1_U3973), .Z(
        P1_U3581) );
  MUX2_X1 U10686 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9797), .S(P1_U3973), .Z(
        P1_U3580) );
  MUX2_X1 U10687 ( .A(n10015), .B(P1_DATAO_REG_25__SCAN_IN), .S(n9825), .Z(
        P1_U3579) );
  MUX2_X1 U10688 ( .A(n10047), .B(P1_DATAO_REG_23__SCAN_IN), .S(n9825), .Z(
        P1_U3577) );
  MUX2_X1 U10689 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9798), .S(P1_U3973), .Z(
        P1_U3576) );
  MUX2_X1 U10690 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n10048), .S(P1_U3973), .Z(
        P1_U3575) );
  MUX2_X1 U10691 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9799), .S(P1_U3973), .Z(
        P1_U3572) );
  MUX2_X1 U10692 ( .A(n9800), .B(P1_DATAO_REG_15__SCAN_IN), .S(n9825), .Z(
        P1_U3569) );
  MUX2_X1 U10693 ( .A(n9801), .B(P1_DATAO_REG_14__SCAN_IN), .S(n9825), .Z(
        P1_U3568) );
  MUX2_X1 U10694 ( .A(n9802), .B(P1_DATAO_REG_13__SCAN_IN), .S(n9825), .Z(
        P1_U3567) );
  MUX2_X1 U10695 ( .A(n9803), .B(P1_DATAO_REG_12__SCAN_IN), .S(n9825), .Z(
        P1_U3566) );
  MUX2_X1 U10696 ( .A(n9804), .B(P1_DATAO_REG_11__SCAN_IN), .S(n9825), .Z(
        P1_U3565) );
  MUX2_X1 U10697 ( .A(n9805), .B(P1_DATAO_REG_10__SCAN_IN), .S(n9825), .Z(
        P1_U3564) );
  MUX2_X1 U10698 ( .A(n5343), .B(P1_DATAO_REG_9__SCAN_IN), .S(n9825), .Z(
        P1_U3563) );
  MUX2_X1 U10699 ( .A(n9806), .B(P1_DATAO_REG_7__SCAN_IN), .S(n9825), .Z(
        P1_U3561) );
  MUX2_X1 U10700 ( .A(n9807), .B(P1_DATAO_REG_6__SCAN_IN), .S(n9825), .Z(
        P1_U3560) );
  MUX2_X1 U10701 ( .A(n9808), .B(P1_DATAO_REG_5__SCAN_IN), .S(n9825), .Z(
        P1_U3559) );
  MUX2_X1 U10702 ( .A(n6987), .B(P1_DATAO_REG_4__SCAN_IN), .S(n9825), .Z(
        P1_U3558) );
  MUX2_X1 U10703 ( .A(n10559), .B(P1_DATAO_REG_3__SCAN_IN), .S(n9825), .Z(
        P1_U3557) );
  MUX2_X1 U10704 ( .A(n6970), .B(P1_DATAO_REG_2__SCAN_IN), .S(n9825), .Z(
        P1_U3556) );
  MUX2_X1 U10705 ( .A(n6960), .B(P1_DATAO_REG_1__SCAN_IN), .S(n9825), .Z(
        P1_U3555) );
  OAI211_X1 U10706 ( .C1(n9811), .C2(n9810), .A(n10519), .B(n9809), .ZN(n9819)
         );
  AOI22_X1 U10707 ( .A1(n10534), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n9818) );
  NAND2_X1 U10708 ( .A1(n10528), .A2(n9812), .ZN(n9817) );
  OAI211_X1 U10709 ( .C1(n9815), .C2(n9814), .A(n10524), .B(n9813), .ZN(n9816)
         );
  NAND4_X1 U10710 ( .A1(n9819), .A2(n9818), .A3(n9817), .A4(n9816), .ZN(
        P1_U3244) );
  NOR2_X1 U10711 ( .A1(n9821), .A2(n9820), .ZN(n9822) );
  XNOR2_X1 U10712 ( .A(n9822), .B(P1_IR_REG_0__SCAN_IN), .ZN(n9826) );
  NOR2_X1 U10713 ( .A1(n9823), .A2(n9827), .ZN(n9824) );
  AOI211_X1 U10714 ( .C1(n9827), .C2(n9826), .A(n9825), .B(n9824), .ZN(n10532)
         );
  INV_X1 U10715 ( .A(n10532), .ZN(n9841) );
  INV_X1 U10716 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n9829) );
  INV_X1 U10717 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n9828) );
  OAI22_X1 U10718 ( .A1(n9921), .A2(n9829), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9828), .ZN(n9830) );
  AOI21_X1 U10719 ( .B1(n10528), .B2(n9831), .A(n9830), .ZN(n9840) );
  OAI211_X1 U10720 ( .C1(n9834), .C2(n9833), .A(n10524), .B(n9832), .ZN(n9839)
         );
  OAI211_X1 U10721 ( .C1(n9837), .C2(n9836), .A(n10519), .B(n9835), .ZN(n9838)
         );
  NAND4_X1 U10722 ( .A1(n9841), .A2(n9840), .A3(n9839), .A4(n9838), .ZN(
        P1_U3245) );
  OAI211_X1 U10723 ( .C1(n9844), .C2(n9843), .A(n10519), .B(n9842), .ZN(n9854)
         );
  INV_X1 U10724 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n9846) );
  OAI21_X1 U10725 ( .B1(n9921), .B2(n9846), .A(n9845), .ZN(n9847) );
  AOI21_X1 U10726 ( .B1(n10528), .B2(n9848), .A(n9847), .ZN(n9853) );
  OAI211_X1 U10727 ( .C1(n9851), .C2(n9850), .A(n10524), .B(n9849), .ZN(n9852)
         );
  NAND3_X1 U10728 ( .A1(n9854), .A2(n9853), .A3(n9852), .ZN(P1_U3246) );
  NOR2_X1 U10729 ( .A1(n9855), .A2(n9864), .ZN(n9857) );
  NOR2_X1 U10730 ( .A1(n9857), .A2(n9856), .ZN(n9860) );
  INV_X1 U10731 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n9858) );
  AOI22_X1 U10732 ( .A1(n9881), .A2(P1_REG1_REG_16__SCAN_IN), .B1(n9858), .B2(
        n9863), .ZN(n9859) );
  NAND2_X1 U10733 ( .A1(n9859), .A2(n9860), .ZN(n9880) );
  OAI21_X1 U10734 ( .B1(n9860), .B2(n9859), .A(n9880), .ZN(n9873) );
  NAND2_X1 U10735 ( .A1(n10534), .A2(P1_ADDR_REG_16__SCAN_IN), .ZN(n9861) );
  OAI211_X1 U10736 ( .C1(n9887), .C2(n9863), .A(n9862), .B(n9861), .ZN(n9872)
         );
  NOR2_X1 U10737 ( .A1(n9865), .A2(n9864), .ZN(n9867) );
  NAND2_X1 U10738 ( .A1(n9881), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n9868) );
  OAI21_X1 U10739 ( .B1(n9881), .B2(P1_REG2_REG_16__SCAN_IN), .A(n9868), .ZN(
        n9869) );
  NOR2_X1 U10740 ( .A1(n9870), .A2(n9869), .ZN(n9876) );
  AOI211_X1 U10741 ( .C1(n9870), .C2(n9869), .A(n9876), .B(n9894), .ZN(n9871)
         );
  AOI211_X1 U10742 ( .C1(n10519), .C2(n9873), .A(n9872), .B(n9871), .ZN(n9874)
         );
  INV_X1 U10743 ( .A(n9874), .ZN(P1_U3259) );
  NOR2_X1 U10744 ( .A1(n9898), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n9875) );
  AOI21_X1 U10745 ( .B1(P1_REG2_REG_17__SCAN_IN), .B2(n9898), .A(n9875), .ZN(
        n9878) );
  NAND2_X1 U10746 ( .A1(n9878), .A2(n9877), .ZN(n9892) );
  OAI21_X1 U10747 ( .B1(n9878), .B2(n9877), .A(n9892), .ZN(n9879) );
  NAND2_X1 U10748 ( .A1(n9879), .A2(n10524), .ZN(n9891) );
  INV_X1 U10749 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n10217) );
  AOI22_X1 U10750 ( .A1(n9898), .A2(P1_REG1_REG_17__SCAN_IN), .B1(n10217), 
        .B2(n9886), .ZN(n9883) );
  OAI21_X1 U10751 ( .B1(n9881), .B2(P1_REG1_REG_16__SCAN_IN), .A(n9880), .ZN(
        n9882) );
  NAND2_X1 U10752 ( .A1(n9883), .A2(n9882), .ZN(n9897) );
  OAI21_X1 U10753 ( .B1(n9883), .B2(n9882), .A(n9897), .ZN(n9889) );
  NAND2_X1 U10754 ( .A1(n10534), .A2(P1_ADDR_REG_17__SCAN_IN), .ZN(n9884) );
  OAI211_X1 U10755 ( .C1(n9887), .C2(n9886), .A(n9885), .B(n9884), .ZN(n9888)
         );
  AOI21_X1 U10756 ( .B1(n9889), .B2(n10519), .A(n9888), .ZN(n9890) );
  NAND2_X1 U10757 ( .A1(n9891), .A2(n9890), .ZN(P1_U3260) );
  OAI21_X1 U10758 ( .B1(n9898), .B2(P1_REG2_REG_17__SCAN_IN), .A(n9892), .ZN(
        n9896) );
  INV_X1 U10759 ( .A(n9893), .ZN(n9901) );
  NAND2_X1 U10760 ( .A1(n9901), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9913) );
  OAI21_X1 U10761 ( .B1(n9901), .B2(P1_REG2_REG_18__SCAN_IN), .A(n9913), .ZN(
        n9895) );
  NOR2_X1 U10762 ( .A1(n9896), .A2(n9895), .ZN(n9915) );
  AOI211_X1 U10763 ( .C1(n9896), .C2(n9895), .A(n9894), .B(n9915), .ZN(n9907)
         );
  NAND2_X1 U10764 ( .A1(n9901), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n9908) );
  OAI21_X1 U10765 ( .B1(n9901), .B2(P1_REG1_REG_18__SCAN_IN), .A(n9908), .ZN(
        n9900) );
  OAI21_X1 U10766 ( .B1(P1_REG1_REG_17__SCAN_IN), .B2(n9898), .A(n9897), .ZN(
        n9899) );
  NOR2_X1 U10767 ( .A1(n9899), .A2(n9900), .ZN(n9910) );
  AOI211_X1 U10768 ( .C1(n9900), .C2(n9899), .A(n9926), .B(n9910), .ZN(n9906)
         );
  INV_X1 U10769 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n9904) );
  NAND2_X1 U10770 ( .A1(n10528), .A2(n9901), .ZN(n9903) );
  OAI211_X1 U10771 ( .C1(n9904), .C2(n9921), .A(n9903), .B(n9902), .ZN(n9905)
         );
  OR3_X1 U10772 ( .A1(n9907), .A2(n9906), .A3(n9905), .ZN(P1_U3261) );
  INV_X1 U10773 ( .A(n9908), .ZN(n9909) );
  NOR2_X1 U10774 ( .A1(n9910), .A2(n9909), .ZN(n9912) );
  XNOR2_X1 U10775 ( .A(n6070), .B(n10206), .ZN(n9911) );
  XNOR2_X1 U10776 ( .A(n9912), .B(n9911), .ZN(n9927) );
  INV_X1 U10777 ( .A(n9913), .ZN(n9914) );
  XNOR2_X1 U10778 ( .A(n6070), .B(P1_REG2_REG_19__SCAN_IN), .ZN(n9916) );
  XNOR2_X1 U10779 ( .A(n9917), .B(n9916), .ZN(n9918) );
  NAND2_X1 U10780 ( .A1(n9918), .A2(n10524), .ZN(n9925) );
  OAI21_X1 U10781 ( .B1(n9921), .B2(n9920), .A(n9919), .ZN(n9922) );
  AOI21_X1 U10782 ( .B1(n10528), .B2(n9923), .A(n9922), .ZN(n9924) );
  OAI211_X1 U10783 ( .C1(n9927), .C2(n9926), .A(n9925), .B(n9924), .ZN(
        P1_U3262) );
  NOR2_X1 U10784 ( .A1(n4941), .A2(n10155), .ZN(n9933) );
  NOR2_X1 U10785 ( .A1(n4948), .A2(n10612), .ZN(n9928) );
  AOI211_X1 U10786 ( .C1(n4941), .C2(P1_REG2_REG_31__SCAN_IN), .A(n9933), .B(
        n9928), .ZN(n9929) );
  OAI21_X1 U10787 ( .B1(n9930), .B2(n10608), .A(n9929), .ZN(P1_U3263) );
  OAI211_X1 U10788 ( .C1(n10245), .C2(n9947), .A(n10552), .B(n9931), .ZN(
        n10156) );
  NOR2_X1 U10789 ( .A1(n10245), .A2(n10612), .ZN(n9932) );
  AOI211_X1 U10790 ( .C1(n4941), .C2(P1_REG2_REG_30__SCAN_IN), .A(n9933), .B(
        n9932), .ZN(n9934) );
  OAI21_X1 U10791 ( .B1(n10608), .B2(n10156), .A(n9934), .ZN(P1_U3264) );
  NAND2_X1 U10792 ( .A1(n9936), .A2(n9935), .ZN(n9937) );
  NOR2_X1 U10793 ( .A1(n9939), .A2(n9938), .ZN(n9940) );
  XNOR2_X1 U10794 ( .A(n9946), .B(n9945), .ZN(n10159) );
  NAND2_X1 U10795 ( .A1(n10159), .A2(n10615), .ZN(n9953) );
  AOI211_X1 U10796 ( .C1(n10161), .C2(n9948), .A(n10663), .B(n9947), .ZN(
        n10160) );
  AOI22_X1 U10797 ( .A1(n10619), .A2(P1_REG2_REG_29__SCAN_IN), .B1(n9949), 
        .B2(n10572), .ZN(n9950) );
  OAI21_X1 U10798 ( .B1(n10163), .B2(n10612), .A(n9950), .ZN(n9951) );
  AOI21_X1 U10799 ( .B1(n10160), .B2(n10576), .A(n9951), .ZN(n9952) );
  OAI211_X1 U10800 ( .C1(n9954), .C2(n4941), .A(n9953), .B(n9952), .ZN(
        P1_U3356) );
  NAND2_X1 U10801 ( .A1(n9955), .A2(n10615), .ZN(n9963) );
  INV_X1 U10802 ( .A(n9956), .ZN(n9961) );
  AOI22_X1 U10803 ( .A1(n10619), .A2(P1_REG2_REG_28__SCAN_IN), .B1(n9957), 
        .B2(n10572), .ZN(n9958) );
  OAI21_X1 U10804 ( .B1(n9959), .B2(n10612), .A(n9958), .ZN(n9960) );
  AOI21_X1 U10805 ( .B1(n9961), .B2(n10576), .A(n9960), .ZN(n9962) );
  OAI211_X1 U10806 ( .C1(n9964), .C2(n4941), .A(n9963), .B(n9962), .ZN(
        P1_U3265) );
  NAND2_X1 U10807 ( .A1(n9965), .A2(n10002), .ZN(n9968) );
  AOI22_X1 U10808 ( .A1(n10619), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n9966), 
        .B2(n10572), .ZN(n9967) );
  OAI211_X1 U10809 ( .C1(n9969), .C2(n10612), .A(n9968), .B(n9967), .ZN(n9970)
         );
  AOI21_X1 U10810 ( .B1(n9971), .B2(n7834), .A(n9970), .ZN(n9972) );
  OAI21_X1 U10811 ( .B1(n9973), .B2(n10154), .A(n9972), .ZN(P1_U3266) );
  XNOR2_X1 U10812 ( .A(n9974), .B(n9980), .ZN(n10170) );
  INV_X1 U10813 ( .A(n10249), .ZN(n10173) );
  INV_X1 U10814 ( .A(n9975), .ZN(n10000) );
  OAI211_X1 U10815 ( .C1(n10173), .C2(n10000), .A(n9976), .B(n10552), .ZN(
        n10168) );
  INV_X1 U10816 ( .A(n10168), .ZN(n9989) );
  AOI22_X1 U10817 ( .A1(n10619), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n9977), 
        .B2(n10572), .ZN(n9978) );
  OAI21_X1 U10818 ( .B1(n10173), .B2(n10612), .A(n9978), .ZN(n9988) );
  NAND2_X1 U10819 ( .A1(n9981), .A2(n9980), .ZN(n9982) );
  NAND2_X1 U10820 ( .A1(n5368), .A2(n9982), .ZN(n9986) );
  NAND2_X1 U10821 ( .A1(n10015), .A2(n10557), .ZN(n9983) );
  OAI21_X1 U10822 ( .B1(n9984), .B2(n10145), .A(n9983), .ZN(n9985) );
  AOI21_X1 U10823 ( .B1(n9986), .B2(n10127), .A(n9985), .ZN(n10169) );
  NOR2_X1 U10824 ( .A1(n10169), .A2(n4941), .ZN(n9987) );
  AOI211_X1 U10825 ( .C1(n9989), .C2(n10576), .A(n9988), .B(n9987), .ZN(n9990)
         );
  OAI21_X1 U10826 ( .B1(n10170), .B2(n10154), .A(n9990), .ZN(P1_U3267) );
  XOR2_X1 U10827 ( .A(n9991), .B(n9993), .Z(n10178) );
  INV_X1 U10828 ( .A(n9992), .ZN(n9995) );
  INV_X1 U10829 ( .A(n9993), .ZN(n9994) );
  AOI21_X1 U10830 ( .B1(n9995), .B2(n9994), .A(n10561), .ZN(n9999) );
  OAI22_X1 U10831 ( .A1(n10031), .A2(n10143), .B1(n9996), .B2(n10145), .ZN(
        n9997) );
  AOI21_X1 U10832 ( .B1(n9999), .B2(n9998), .A(n9997), .ZN(n10177) );
  INV_X1 U10833 ( .A(n10177), .ZN(n10008) );
  INV_X1 U10834 ( .A(n10018), .ZN(n10001) );
  AOI21_X1 U10835 ( .B1(n10174), .B2(n10001), .A(n10000), .ZN(n10175) );
  NAND2_X1 U10836 ( .A1(n10175), .A2(n10002), .ZN(n10005) );
  AOI22_X1 U10837 ( .A1(n10619), .A2(P1_REG2_REG_25__SCAN_IN), .B1(n10003), 
        .B2(n10572), .ZN(n10004) );
  OAI211_X1 U10838 ( .C1(n10006), .C2(n10612), .A(n10005), .B(n10004), .ZN(
        n10007) );
  AOI21_X1 U10839 ( .B1(n10008), .B2(n7834), .A(n10007), .ZN(n10009) );
  OAI21_X1 U10840 ( .B1(n10178), .B2(n10154), .A(n10009), .ZN(P1_U3268) );
  XNOR2_X1 U10841 ( .A(n10011), .B(n10010), .ZN(n10183) );
  OAI211_X1 U10842 ( .C1(n10014), .C2(n10013), .A(n10012), .B(n10127), .ZN(
        n10017) );
  AOI22_X1 U10843 ( .A1(n10557), .A2(n10047), .B1(n10015), .B2(n10558), .ZN(
        n10016) );
  NAND2_X1 U10844 ( .A1(n10017), .A2(n10016), .ZN(n10179) );
  AOI211_X1 U10845 ( .C1(n10181), .C2(n10032), .A(n10663), .B(n10018), .ZN(
        n10180) );
  NAND2_X1 U10846 ( .A1(n10180), .A2(n10576), .ZN(n10021) );
  AOI22_X1 U10847 ( .A1(n10619), .A2(P1_REG2_REG_24__SCAN_IN), .B1(n10019), 
        .B2(n10572), .ZN(n10020) );
  OAI211_X1 U10848 ( .C1(n10022), .C2(n10612), .A(n10021), .B(n10020), .ZN(
        n10023) );
  AOI21_X1 U10849 ( .B1(n10179), .B2(n7834), .A(n10023), .ZN(n10024) );
  OAI21_X1 U10850 ( .B1(n10183), .B2(n10154), .A(n10024), .ZN(P1_U3269) );
  XOR2_X1 U10851 ( .A(n10029), .B(n10025), .Z(n10187) );
  INV_X1 U10852 ( .A(n10026), .ZN(n10027) );
  AOI21_X1 U10853 ( .B1(n10029), .B2(n10028), .A(n10027), .ZN(n10030) );
  OAI222_X1 U10854 ( .A1(n10145), .A2(n10031), .B1(n10143), .B2(n10065), .C1(
        n10561), .C2(n10030), .ZN(n10184) );
  INV_X1 U10855 ( .A(n10032), .ZN(n10033) );
  AOI211_X1 U10856 ( .C1(n6101), .C2(n10051), .A(n10663), .B(n10033), .ZN(
        n10185) );
  NAND2_X1 U10857 ( .A1(n10185), .A2(n10576), .ZN(n10036) );
  AOI22_X1 U10858 ( .A1(n10619), .A2(P1_REG2_REG_23__SCAN_IN), .B1(n10034), 
        .B2(n10572), .ZN(n10035) );
  OAI211_X1 U10859 ( .C1(n10037), .C2(n10612), .A(n10036), .B(n10035), .ZN(
        n10038) );
  AOI21_X1 U10860 ( .B1(n10184), .B2(n7834), .A(n10038), .ZN(n10039) );
  OAI21_X1 U10861 ( .B1(n10187), .B2(n10154), .A(n10039), .ZN(P1_U3270) );
  OAI21_X1 U10862 ( .B1(n10042), .B2(n10041), .A(n10040), .ZN(n10043) );
  INV_X1 U10863 ( .A(n10043), .ZN(n10192) );
  OAI211_X1 U10864 ( .C1(n10046), .C2(n10045), .A(n10044), .B(n10127), .ZN(
        n10050) );
  AOI22_X1 U10865 ( .A1(n10048), .A2(n10557), .B1(n10558), .B2(n10047), .ZN(
        n10049) );
  NAND2_X1 U10866 ( .A1(n10050), .A2(n10049), .ZN(n10188) );
  INV_X1 U10867 ( .A(n10051), .ZN(n10052) );
  AOI211_X1 U10868 ( .C1(n10190), .C2(n5204), .A(n10663), .B(n10052), .ZN(
        n10189) );
  NAND2_X1 U10869 ( .A1(n10189), .A2(n10576), .ZN(n10055) );
  AOI22_X1 U10870 ( .A1(n10619), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n10053), 
        .B2(n10572), .ZN(n10054) );
  OAI211_X1 U10871 ( .C1(n5977), .C2(n10612), .A(n10055), .B(n10054), .ZN(
        n10056) );
  AOI21_X1 U10872 ( .B1(n10188), .B2(n7834), .A(n10056), .ZN(n10057) );
  OAI21_X1 U10873 ( .B1(n10192), .B2(n10154), .A(n10057), .ZN(P1_U3271) );
  AOI21_X1 U10874 ( .B1(n10062), .B2(n10058), .A(n10059), .ZN(n10195) );
  INV_X1 U10875 ( .A(n10195), .ZN(n10076) );
  NAND2_X1 U10876 ( .A1(n10061), .A2(n10060), .ZN(n10063) );
  XNOR2_X1 U10877 ( .A(n10063), .B(n10062), .ZN(n10064) );
  NAND2_X1 U10878 ( .A1(n10064), .A2(n10127), .ZN(n10068) );
  OAI22_X1 U10879 ( .A1(n10065), .A2(n10145), .B1(n10097), .B2(n10143), .ZN(
        n10066) );
  INV_X1 U10880 ( .A(n10066), .ZN(n10067) );
  NAND2_X1 U10881 ( .A1(n10068), .A2(n10067), .ZN(n10193) );
  AOI211_X1 U10882 ( .C1(n10070), .C2(n10082), .A(n10663), .B(n10069), .ZN(
        n10194) );
  NAND2_X1 U10883 ( .A1(n10194), .A2(n10576), .ZN(n10073) );
  AOI22_X1 U10884 ( .A1(n10619), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n10071), 
        .B2(n10572), .ZN(n10072) );
  OAI211_X1 U10885 ( .C1(n5202), .C2(n10612), .A(n10073), .B(n10072), .ZN(
        n10074) );
  AOI21_X1 U10886 ( .B1(n10193), .B2(n7834), .A(n10074), .ZN(n10075) );
  OAI21_X1 U10887 ( .B1(n10076), .B2(n10154), .A(n10075), .ZN(P1_U3272) );
  XOR2_X1 U10888 ( .A(n10077), .B(n10078), .Z(n10202) );
  XOR2_X1 U10889 ( .A(n10079), .B(n10078), .Z(n10080) );
  OAI222_X1 U10890 ( .A1(n10145), .A2(n10081), .B1(n10143), .B2(n10111), .C1(
        n10080), .C2(n10561), .ZN(n10198) );
  INV_X1 U10891 ( .A(n10200), .ZN(n10087) );
  INV_X1 U10892 ( .A(n10082), .ZN(n10083) );
  AOI211_X1 U10893 ( .C1(n10200), .C2(n10090), .A(n10663), .B(n10083), .ZN(
        n10199) );
  NAND2_X1 U10894 ( .A1(n10199), .A2(n10576), .ZN(n10086) );
  AOI22_X1 U10895 ( .A1(n10619), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n10084), 
        .B2(n10572), .ZN(n10085) );
  OAI211_X1 U10896 ( .C1(n10087), .C2(n10612), .A(n10086), .B(n10085), .ZN(
        n10088) );
  AOI21_X1 U10897 ( .B1(n10198), .B2(n7834), .A(n10088), .ZN(n10089) );
  OAI21_X1 U10898 ( .B1(n10202), .B2(n10154), .A(n10089), .ZN(P1_U3273) );
  INV_X1 U10899 ( .A(n10113), .ZN(n10092) );
  INV_X1 U10900 ( .A(n10090), .ZN(n10091) );
  AOI211_X1 U10901 ( .C1(n10102), .C2(n10092), .A(n10663), .B(n10091), .ZN(
        n10204) );
  INV_X1 U10902 ( .A(n10093), .ZN(n10094) );
  AOI21_X1 U10903 ( .B1(n5463), .B2(n10095), .A(n10094), .ZN(n10096) );
  OAI222_X1 U10904 ( .A1(n10145), .A2(n10097), .B1(n10143), .B2(n10124), .C1(
        n10561), .C2(n10096), .ZN(n10203) );
  AOI21_X1 U10905 ( .B1(n10204), .B2(n6070), .A(n10203), .ZN(n10105) );
  XNOR2_X1 U10906 ( .A(n10098), .B(n5463), .ZN(n10205) );
  NAND2_X1 U10907 ( .A1(n10205), .A2(n10615), .ZN(n10104) );
  INV_X1 U10908 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n10100) );
  OAI22_X1 U10909 ( .A1(n7834), .A2(n10100), .B1(n10099), .B2(n10606), .ZN(
        n10101) );
  AOI21_X1 U10910 ( .B1(n10102), .B2(n10570), .A(n10101), .ZN(n10103) );
  OAI211_X1 U10911 ( .C1(n4941), .C2(n10105), .A(n10104), .B(n10103), .ZN(
        P1_U3274) );
  XNOR2_X1 U10912 ( .A(n10107), .B(n10106), .ZN(n10212) );
  XNOR2_X1 U10913 ( .A(n10109), .B(n10108), .ZN(n10110) );
  OAI222_X1 U10914 ( .A1(n10145), .A2(n10111), .B1(n10143), .B2(n10144), .C1(
        n10561), .C2(n10110), .ZN(n10208) );
  INV_X1 U10915 ( .A(n10112), .ZN(n10129) );
  AOI211_X1 U10916 ( .C1(n10210), .C2(n10129), .A(n10663), .B(n10113), .ZN(
        n10209) );
  NAND2_X1 U10917 ( .A1(n10209), .A2(n10576), .ZN(n10116) );
  AOI22_X1 U10918 ( .A1(n10619), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n10114), 
        .B2(n10572), .ZN(n10115) );
  OAI211_X1 U10919 ( .C1(n10117), .C2(n10612), .A(n10116), .B(n10115), .ZN(
        n10118) );
  AOI21_X1 U10920 ( .B1(n10208), .B2(n7834), .A(n10118), .ZN(n10119) );
  OAI21_X1 U10921 ( .B1(n10212), .B2(n10154), .A(n10119), .ZN(P1_U3275) );
  XNOR2_X1 U10922 ( .A(n10120), .B(n10121), .ZN(n10215) );
  INV_X1 U10923 ( .A(n10121), .ZN(n10122) );
  XNOR2_X1 U10924 ( .A(n10123), .B(n10122), .ZN(n10128) );
  OAI22_X1 U10925 ( .A1(n10125), .A2(n10143), .B1(n10124), .B2(n10145), .ZN(
        n10126) );
  AOI21_X1 U10926 ( .B1(n10128), .B2(n10127), .A(n10126), .ZN(n10214) );
  INV_X1 U10927 ( .A(n10214), .ZN(n10135) );
  OAI211_X1 U10928 ( .C1(n10268), .C2(n10146), .A(n10129), .B(n10552), .ZN(
        n10213) );
  AOI22_X1 U10929 ( .A1(n10619), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n10572), 
        .B2(n10130), .ZN(n10133) );
  NAND2_X1 U10930 ( .A1(n10131), .A2(n10570), .ZN(n10132) );
  OAI211_X1 U10931 ( .C1(n10213), .C2(n10608), .A(n10133), .B(n10132), .ZN(
        n10134) );
  AOI21_X1 U10932 ( .B1(n10135), .B2(n7834), .A(n10134), .ZN(n10136) );
  OAI21_X1 U10933 ( .B1(n10215), .B2(n10154), .A(n10136), .ZN(P1_U3276) );
  XNOR2_X1 U10934 ( .A(n10138), .B(n10137), .ZN(n10224) );
  XNOR2_X1 U10935 ( .A(n10140), .B(n10139), .ZN(n10141) );
  OAI222_X1 U10936 ( .A1(n10145), .A2(n10144), .B1(n10143), .B2(n10142), .C1(
        n10141), .C2(n10561), .ZN(n10220) );
  INV_X1 U10937 ( .A(n10222), .ZN(n10151) );
  AOI211_X1 U10938 ( .C1(n10222), .C2(n10147), .A(n10663), .B(n10146), .ZN(
        n10221) );
  NAND2_X1 U10939 ( .A1(n10221), .A2(n10576), .ZN(n10150) );
  AOI22_X1 U10940 ( .A1(n10619), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n10148), 
        .B2(n10572), .ZN(n10149) );
  OAI211_X1 U10941 ( .C1(n10151), .C2(n10612), .A(n10150), .B(n10149), .ZN(
        n10152) );
  AOI21_X1 U10942 ( .B1(n10220), .B2(n7834), .A(n10152), .ZN(n10153) );
  OAI21_X1 U10943 ( .B1(n10224), .B2(n10154), .A(n10153), .ZN(P1_U3277) );
  INV_X1 U10944 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n10157) );
  AND2_X1 U10945 ( .A1(n10156), .A2(n10155), .ZN(n10242) );
  MUX2_X1 U10946 ( .A(n10157), .B(n10242), .S(n10646), .Z(n10158) );
  OAI21_X1 U10947 ( .B1(n10245), .B2(n10219), .A(n10158), .ZN(P1_U3552) );
  NAND2_X1 U10948 ( .A1(n10159), .A2(n10667), .ZN(n10167) );
  INV_X1 U10949 ( .A(n10160), .ZN(n10164) );
  INV_X1 U10950 ( .A(n10161), .ZN(n10163) );
  INV_X1 U10951 ( .A(n10649), .ZN(n10162) );
  NAND2_X1 U10952 ( .A1(n10167), .A2(n10166), .ZN(n10246) );
  MUX2_X1 U10953 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n10246), .S(n10646), .Z(
        P1_U3551) );
  OAI211_X1 U10954 ( .C1(n10170), .C2(n10239), .A(n10169), .B(n10168), .ZN(
        n10247) );
  MUX2_X1 U10955 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n10247), .S(n10646), .Z(
        n10171) );
  INV_X1 U10956 ( .A(n10171), .ZN(n10172) );
  OAI21_X1 U10957 ( .B1(n10173), .B2(n10219), .A(n10172), .ZN(P1_U3548) );
  AOI22_X1 U10958 ( .A1(n10175), .A2(n10552), .B1(n10649), .B2(n10174), .ZN(
        n10176) );
  OAI211_X1 U10959 ( .C1(n10178), .C2(n10239), .A(n10177), .B(n10176), .ZN(
        n10251) );
  MUX2_X1 U10960 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n10251), .S(n10646), .Z(
        P1_U3547) );
  AOI211_X1 U10961 ( .C1(n10649), .C2(n10181), .A(n10180), .B(n10179), .ZN(
        n10182) );
  OAI21_X1 U10962 ( .B1(n10183), .B2(n10239), .A(n10182), .ZN(n10252) );
  MUX2_X1 U10963 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n10252), .S(n10646), .Z(
        P1_U3546) );
  AOI211_X1 U10964 ( .C1(n10649), .C2(n6101), .A(n10185), .B(n10184), .ZN(
        n10186) );
  OAI21_X1 U10965 ( .B1(n10187), .B2(n10239), .A(n10186), .ZN(n10253) );
  MUX2_X1 U10966 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n10253), .S(n10646), .Z(
        P1_U3545) );
  AOI211_X1 U10967 ( .C1(n10649), .C2(n10190), .A(n10189), .B(n10188), .ZN(
        n10191) );
  OAI21_X1 U10968 ( .B1(n10192), .B2(n10239), .A(n10191), .ZN(n10254) );
  MUX2_X1 U10969 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n10254), .S(n10646), .Z(
        P1_U3544) );
  INV_X1 U10970 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n10196) );
  AOI211_X1 U10971 ( .C1(n10195), .C2(n10667), .A(n10194), .B(n10193), .ZN(
        n10255) );
  MUX2_X1 U10972 ( .A(n10196), .B(n10255), .S(n10646), .Z(n10197) );
  OAI21_X1 U10973 ( .B1(n5202), .B2(n10219), .A(n10197), .ZN(P1_U3543) );
  AOI211_X1 U10974 ( .C1(n10649), .C2(n10200), .A(n10199), .B(n10198), .ZN(
        n10201) );
  OAI21_X1 U10975 ( .B1(n10202), .B2(n10239), .A(n10201), .ZN(n10258) );
  MUX2_X1 U10976 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n10258), .S(n10646), .Z(
        P1_U3542) );
  AOI211_X1 U10977 ( .C1(n10205), .C2(n10667), .A(n10204), .B(n10203), .ZN(
        n10259) );
  MUX2_X1 U10978 ( .A(n10206), .B(n10259), .S(n10646), .Z(n10207) );
  OAI21_X1 U10979 ( .B1(n10262), .B2(n10219), .A(n10207), .ZN(P1_U3541) );
  AOI211_X1 U10980 ( .C1(n10649), .C2(n10210), .A(n10209), .B(n10208), .ZN(
        n10211) );
  OAI21_X1 U10981 ( .B1(n10212), .B2(n10239), .A(n10211), .ZN(n10263) );
  MUX2_X1 U10982 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n10263), .S(n10646), .Z(
        P1_U3540) );
  OAI211_X1 U10983 ( .C1(n10215), .C2(n10239), .A(n10214), .B(n10213), .ZN(
        n10216) );
  INV_X1 U10984 ( .A(n10216), .ZN(n10264) );
  MUX2_X1 U10985 ( .A(n10217), .B(n10264), .S(n10646), .Z(n10218) );
  OAI21_X1 U10986 ( .B1(n10268), .B2(n10219), .A(n10218), .ZN(P1_U3539) );
  AOI211_X1 U10987 ( .C1(n10649), .C2(n10222), .A(n10221), .B(n10220), .ZN(
        n10223) );
  OAI21_X1 U10988 ( .B1(n10224), .B2(n10239), .A(n10223), .ZN(n10269) );
  MUX2_X1 U10989 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n10269), .S(n10646), .Z(
        P1_U3538) );
  AOI22_X1 U10990 ( .A1(n10226), .A2(n10552), .B1(n10649), .B2(n10225), .ZN(
        n10227) );
  OAI211_X1 U10991 ( .C1(n10229), .C2(n10239), .A(n10228), .B(n10227), .ZN(
        n10270) );
  MUX2_X1 U10992 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n10270), .S(n10646), .Z(
        P1_U3537) );
  AOI22_X1 U10993 ( .A1(n10231), .A2(n10552), .B1(n10649), .B2(n10230), .ZN(
        n10232) );
  OAI211_X1 U10994 ( .C1(n10239), .C2(n10234), .A(n10233), .B(n10232), .ZN(
        n10271) );
  MUX2_X1 U10995 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n10271), .S(n10646), .Z(
        P1_U3536) );
  AOI22_X1 U10996 ( .A1(n10236), .A2(n10552), .B1(n10649), .B2(n10235), .ZN(
        n10237) );
  OAI211_X1 U10997 ( .C1(n10240), .C2(n10239), .A(n10238), .B(n10237), .ZN(
        n10272) );
  MUX2_X1 U10998 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n10272), .S(n10646), .Z(
        P1_U3535) );
  MUX2_X1 U10999 ( .A(P1_REG1_REG_0__SCAN_IN), .B(n10241), .S(n10646), .Z(
        P1_U3522) );
  INV_X1 U11000 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n10243) );
  MUX2_X1 U11001 ( .A(n10243), .B(n10242), .S(n10674), .Z(n10244) );
  OAI21_X1 U11002 ( .B1(n10245), .B2(n10267), .A(n10244), .ZN(P1_U3520) );
  MUX2_X1 U11003 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n10246), .S(n10674), .Z(
        P1_U3519) );
  MUX2_X1 U11004 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n10247), .S(n10674), .Z(
        n10248) );
  AOI21_X1 U11005 ( .B1(n6155), .B2(n10249), .A(n10248), .ZN(n10250) );
  INV_X1 U11006 ( .A(n10250), .ZN(P1_U3516) );
  MUX2_X1 U11007 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n10251), .S(n10674), .Z(
        P1_U3515) );
  MUX2_X1 U11008 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n10252), .S(n10674), .Z(
        P1_U3514) );
  MUX2_X1 U11009 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n10253), .S(n10674), .Z(
        P1_U3513) );
  MUX2_X1 U11010 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n10254), .S(n10674), .Z(
        P1_U3512) );
  INV_X1 U11011 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n10256) );
  MUX2_X1 U11012 ( .A(n10256), .B(n10255), .S(n10674), .Z(n10257) );
  OAI21_X1 U11013 ( .B1(n5202), .B2(n10267), .A(n10257), .ZN(P1_U3511) );
  MUX2_X1 U11014 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n10258), .S(n10674), .Z(
        P1_U3510) );
  INV_X1 U11015 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n10260) );
  MUX2_X1 U11016 ( .A(n10260), .B(n10259), .S(n10674), .Z(n10261) );
  OAI21_X1 U11017 ( .B1(n10262), .B2(n10267), .A(n10261), .ZN(P1_U3509) );
  MUX2_X1 U11018 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n10263), .S(n10674), .Z(
        P1_U3507) );
  INV_X1 U11019 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n10265) );
  MUX2_X1 U11020 ( .A(n10265), .B(n10264), .S(n10674), .Z(n10266) );
  OAI21_X1 U11021 ( .B1(n10268), .B2(n10267), .A(n10266), .ZN(P1_U3504) );
  MUX2_X1 U11022 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n10269), .S(n10674), .Z(
        P1_U3501) );
  MUX2_X1 U11023 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n10270), .S(n10674), .Z(
        P1_U3498) );
  MUX2_X1 U11024 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n10271), .S(n10674), .Z(
        P1_U3495) );
  MUX2_X1 U11025 ( .A(P1_REG0_REG_13__SCAN_IN), .B(n10272), .S(n10674), .Z(
        P1_U3492) );
  MUX2_X1 U11026 ( .A(n10275), .B(P1_D_REG_1__SCAN_IN), .S(n4943), .Z(P1_U3440) );
  MUX2_X1 U11027 ( .A(n10276), .B(P1_D_REG_0__SCAN_IN), .S(n4943), .Z(P1_U3439) );
  NOR4_X1 U11028 ( .A1(n5595), .A2(P1_IR_REG_30__SCAN_IN), .A3(P1_U3086), .A4(
        n5590), .ZN(n10277) );
  AOI21_X1 U11029 ( .B1(P2_DATAO_REG_31__SCAN_IN), .B2(n10286), .A(n10277), 
        .ZN(n10278) );
  OAI21_X1 U11030 ( .B1(n10279), .B2(n10293), .A(n10278), .ZN(P1_U3324) );
  AOI22_X1 U11031 ( .A1(n10280), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_30__SCAN_IN), .B2(n10286), .ZN(n10281) );
  OAI21_X1 U11032 ( .B1(n10282), .B2(n10293), .A(n10281), .ZN(P1_U3325) );
  AOI22_X1 U11033 ( .A1(n10283), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n10286), .ZN(n10284) );
  OAI21_X1 U11034 ( .B1(n10285), .B2(n10293), .A(n10284), .ZN(P1_U3326) );
  AOI22_X1 U11035 ( .A1(n10287), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(n10286), .ZN(n10288) );
  OAI21_X1 U11036 ( .B1(n10289), .B2(n10293), .A(n10288), .ZN(P1_U3327) );
  INV_X1 U11037 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n10291) );
  OAI222_X1 U11038 ( .A1(P1_U3086), .A2(n10294), .B1(n10293), .B2(n10292), 
        .C1(n10291), .C2(n10290), .ZN(P1_U3328) );
  MUX2_X1 U11039 ( .A(n10295), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  AND2_X1 U11040 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n4943), .ZN(P1_U3323) );
  AND2_X1 U11041 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n4943), .ZN(P1_U3322) );
  AND2_X1 U11042 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n4943), .ZN(P1_U3321) );
  AND2_X1 U11043 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n4943), .ZN(P1_U3320) );
  AND2_X1 U11044 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n4943), .ZN(P1_U3319) );
  AND2_X1 U11045 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n4943), .ZN(P1_U3318) );
  AND2_X1 U11046 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n4943), .ZN(P1_U3317) );
  AND2_X1 U11047 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n4943), .ZN(P1_U3316) );
  AND2_X1 U11048 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n4943), .ZN(P1_U3315) );
  AND2_X1 U11049 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n4943), .ZN(P1_U3314) );
  AND2_X1 U11050 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n4943), .ZN(P1_U3313) );
  AND2_X1 U11051 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n4943), .ZN(P1_U3312) );
  AND2_X1 U11052 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n4943), .ZN(P1_U3311) );
  AND2_X1 U11053 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n4943), .ZN(P1_U3310) );
  AND2_X1 U11054 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n4943), .ZN(P1_U3309) );
  AND2_X1 U11055 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n4943), .ZN(P1_U3308) );
  AND2_X1 U11056 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n4943), .ZN(P1_U3307) );
  AND2_X1 U11057 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n4943), .ZN(P1_U3306) );
  AND2_X1 U11058 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n4943), .ZN(P1_U3305) );
  AND2_X1 U11059 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n4943), .ZN(P1_U3304) );
  AND2_X1 U11060 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n4943), .ZN(P1_U3303) );
  AND2_X1 U11061 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n4943), .ZN(P1_U3302) );
  AND2_X1 U11062 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n4943), .ZN(P1_U3301) );
  AND2_X1 U11063 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n4943), .ZN(P1_U3300) );
  AND2_X1 U11064 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n4943), .ZN(P1_U3299) );
  AND2_X1 U11065 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n4943), .ZN(P1_U3298) );
  AND2_X1 U11066 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n4943), .ZN(P1_U3297) );
  AND2_X1 U11067 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n4943), .ZN(P1_U3296) );
  AND2_X1 U11068 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n4943), .ZN(P1_U3295) );
  AND2_X1 U11069 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n4943), .ZN(P1_U3294) );
  OAI21_X1 U11070 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(n10299), .ZN(n10297) );
  INV_X1 U11071 ( .A(n10297), .ZN(ADD_1068_U46) );
  OAI21_X1 U11072 ( .B1(n10300), .B2(n10299), .A(n10298), .ZN(n10301) );
  XNOR2_X1 U11073 ( .A(n10301), .B(P2_ADDR_REG_1__SCAN_IN), .ZN(ADD_1068_U5)
         );
  AOI21_X1 U11074 ( .B1(n10304), .B2(n10303), .A(n10302), .ZN(ADD_1068_U54) );
  AOI21_X1 U11075 ( .B1(n10307), .B2(n10306), .A(n10305), .ZN(ADD_1068_U53) );
  OAI21_X1 U11076 ( .B1(n10310), .B2(n10309), .A(n10308), .ZN(ADD_1068_U52) );
  OAI21_X1 U11077 ( .B1(n10313), .B2(n10312), .A(n10311), .ZN(ADD_1068_U51) );
  OAI21_X1 U11078 ( .B1(n10316), .B2(n10315), .A(n10314), .ZN(ADD_1068_U50) );
  OAI21_X1 U11079 ( .B1(n10319), .B2(n10318), .A(n10317), .ZN(ADD_1068_U49) );
  OAI21_X1 U11080 ( .B1(n10322), .B2(n10321), .A(n10320), .ZN(ADD_1068_U48) );
  OAI21_X1 U11081 ( .B1(n10325), .B2(n10324), .A(n10323), .ZN(ADD_1068_U47) );
  OAI21_X1 U11082 ( .B1(n10328), .B2(n10327), .A(n10326), .ZN(ADD_1068_U63) );
  OAI21_X1 U11083 ( .B1(n10331), .B2(n10330), .A(n10329), .ZN(ADD_1068_U62) );
  OAI21_X1 U11084 ( .B1(n10334), .B2(n10333), .A(n10332), .ZN(ADD_1068_U61) );
  OAI21_X1 U11085 ( .B1(n10337), .B2(n10336), .A(n10335), .ZN(ADD_1068_U60) );
  OAI21_X1 U11086 ( .B1(n10340), .B2(n10339), .A(n10338), .ZN(ADD_1068_U59) );
  OAI21_X1 U11087 ( .B1(n10343), .B2(n10342), .A(n10341), .ZN(ADD_1068_U58) );
  OAI21_X1 U11088 ( .B1(n10346), .B2(n10345), .A(n10344), .ZN(ADD_1068_U57) );
  OAI21_X1 U11089 ( .B1(n10349), .B2(n10348), .A(n10347), .ZN(ADD_1068_U56) );
  OAI21_X1 U11090 ( .B1(n10352), .B2(n10351), .A(n10350), .ZN(ADD_1068_U55) );
  AOI22_X1 U11091 ( .A1(n10497), .A2(P2_IR_REG_0__SCAN_IN), .B1(n10495), .B2(
        P2_ADDR_REG_0__SCAN_IN), .ZN(n10357) );
  XNOR2_X1 U11092 ( .A(n10353), .B(P2_IR_REG_0__SCAN_IN), .ZN(n10354) );
  OAI21_X1 U11093 ( .B1(n10504), .B2(n10355), .A(n10354), .ZN(n10356) );
  OAI211_X1 U11094 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n10358), .A(n10357), .B(
        n10356), .ZN(P2_U3182) );
  AOI21_X1 U11095 ( .B1(n10497), .B2(n10360), .A(n10359), .ZN(n10374) );
  OAI21_X1 U11096 ( .B1(n10363), .B2(n10362), .A(n10361), .ZN(n10364) );
  AOI22_X1 U11097 ( .A1(n10364), .A2(n10504), .B1(n10495), .B2(
        P2_ADDR_REG_3__SCAN_IN), .ZN(n10373) );
  OAI21_X1 U11098 ( .B1(P2_REG2_REG_3__SCAN_IN), .B2(n10366), .A(n10365), .ZN(
        n10367) );
  NAND2_X1 U11099 ( .A1(n10505), .A2(n10367), .ZN(n10372) );
  XNOR2_X1 U11100 ( .A(n10368), .B(P2_REG1_REG_3__SCAN_IN), .ZN(n10369) );
  NAND2_X1 U11101 ( .A1(n10370), .A2(n10369), .ZN(n10371) );
  NAND4_X1 U11102 ( .A1(n10374), .A2(n10373), .A3(n10372), .A4(n10371), .ZN(
        P2_U3185) );
  INV_X1 U11103 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n10393) );
  AOI21_X1 U11104 ( .B1(n10497), .B2(n10376), .A(n10375), .ZN(n10392) );
  AOI21_X1 U11105 ( .B1(n10379), .B2(n10378), .A(n10377), .ZN(n10389) );
  OAI21_X1 U11106 ( .B1(n10382), .B2(n10381), .A(n10380), .ZN(n10383) );
  NAND2_X1 U11107 ( .A1(n10505), .A2(n10383), .ZN(n10388) );
  OAI211_X1 U11108 ( .C1(n10386), .C2(n10385), .A(n10384), .B(n10504), .ZN(
        n10387) );
  OAI211_X1 U11109 ( .C1(n10511), .C2(n10389), .A(n10388), .B(n10387), .ZN(
        n10390) );
  INV_X1 U11110 ( .A(n10390), .ZN(n10391) );
  OAI211_X1 U11111 ( .C1(n10412), .C2(n10393), .A(n10392), .B(n10391), .ZN(
        P2_U3186) );
  INV_X1 U11112 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n10411) );
  OAI21_X1 U11113 ( .B1(n10395), .B2(n10394), .A(n10504), .ZN(n10397) );
  NOR2_X1 U11114 ( .A1(n10397), .A2(n10396), .ZN(n10408) );
  OAI21_X1 U11115 ( .B1(n10399), .B2(P2_REG2_REG_5__SCAN_IN), .A(n10398), .ZN(
        n10400) );
  AND2_X1 U11116 ( .A1(n10400), .A2(n10505), .ZN(n10407) );
  AOI21_X1 U11117 ( .B1(n10402), .B2(n10401), .A(n5029), .ZN(n10405) );
  OAI22_X1 U11118 ( .A1(n10405), .A2(n10511), .B1(n10404), .B2(n10403), .ZN(
        n10406) );
  NOR4_X1 U11119 ( .A1(n10409), .A2(n10408), .A3(n10407), .A4(n10406), .ZN(
        n10410) );
  OAI21_X1 U11120 ( .B1(n10412), .B2(n10411), .A(n10410), .ZN(P2_U3187) );
  AOI21_X1 U11121 ( .B1(n10497), .B2(n10414), .A(n10413), .ZN(n10430) );
  OAI21_X1 U11122 ( .B1(n10417), .B2(n10416), .A(n10415), .ZN(n10418) );
  AOI22_X1 U11123 ( .A1(n10418), .A2(n10504), .B1(n10495), .B2(
        P2_ADDR_REG_6__SCAN_IN), .ZN(n10429) );
  AOI21_X1 U11124 ( .B1(n10421), .B2(n10420), .A(n10419), .ZN(n10422) );
  OR2_X1 U11125 ( .A1(n10422), .A2(n10511), .ZN(n10428) );
  OAI21_X1 U11126 ( .B1(n10425), .B2(n10424), .A(n10423), .ZN(n10426) );
  NAND2_X1 U11127 ( .A1(n10426), .A2(n10505), .ZN(n10427) );
  NAND4_X1 U11128 ( .A1(n10430), .A2(n10429), .A3(n10428), .A4(n10427), .ZN(
        P2_U3188) );
  AOI22_X1 U11129 ( .A1(n10497), .A2(n10431), .B1(n10495), .B2(
        P2_ADDR_REG_7__SCAN_IN), .ZN(n10446) );
  OAI21_X1 U11130 ( .B1(P2_REG2_REG_7__SCAN_IN), .B2(n10433), .A(n10432), .ZN(
        n10438) );
  OAI21_X1 U11131 ( .B1(n10436), .B2(n10435), .A(n10434), .ZN(n10437) );
  AOI22_X1 U11132 ( .A1(n10438), .A2(n10505), .B1(n10504), .B2(n10437), .ZN(
        n10445) );
  AOI21_X1 U11133 ( .B1(n10441), .B2(n10440), .A(n10439), .ZN(n10442) );
  OR2_X1 U11134 ( .A1(n10511), .A2(n10442), .ZN(n10443) );
  NAND4_X1 U11135 ( .A1(n10446), .A2(n10445), .A3(n10444), .A4(n10443), .ZN(
        P2_U3189) );
  AOI22_X1 U11136 ( .A1(n10497), .A2(n10447), .B1(n10495), .B2(
        P2_ADDR_REG_8__SCAN_IN), .ZN(n10462) );
  OAI21_X1 U11137 ( .B1(n10450), .B2(n10449), .A(n10448), .ZN(n10455) );
  OAI21_X1 U11138 ( .B1(n10453), .B2(n10452), .A(n10451), .ZN(n10454) );
  AOI22_X1 U11139 ( .A1(n10455), .A2(n10505), .B1(n10504), .B2(n10454), .ZN(
        n10461) );
  AOI21_X1 U11140 ( .B1(n5028), .B2(n10457), .A(n10456), .ZN(n10458) );
  OR2_X1 U11141 ( .A1(n10458), .A2(n10511), .ZN(n10459) );
  NAND4_X1 U11142 ( .A1(n10462), .A2(n10461), .A3(n10460), .A4(n10459), .ZN(
        P2_U3190) );
  AOI22_X1 U11143 ( .A1(n10497), .A2(n10463), .B1(n10495), .B2(
        P2_ADDR_REG_9__SCAN_IN), .ZN(n10478) );
  OAI21_X1 U11144 ( .B1(P2_REG2_REG_9__SCAN_IN), .B2(n10465), .A(n10464), .ZN(
        n10470) );
  OAI21_X1 U11145 ( .B1(n10468), .B2(n10467), .A(n10466), .ZN(n10469) );
  AOI22_X1 U11146 ( .A1(n10470), .A2(n10505), .B1(n10504), .B2(n10469), .ZN(
        n10477) );
  AOI21_X1 U11147 ( .B1(n10473), .B2(n10472), .A(n10471), .ZN(n10474) );
  OR2_X1 U11148 ( .A1(n10511), .A2(n10474), .ZN(n10475) );
  NAND4_X1 U11149 ( .A1(n10478), .A2(n10477), .A3(n10476), .A4(n10475), .ZN(
        P2_U3191) );
  AOI22_X1 U11150 ( .A1(n10497), .A2(n10479), .B1(n10495), .B2(
        P2_ADDR_REG_10__SCAN_IN), .ZN(n10494) );
  OAI21_X1 U11151 ( .B1(n10482), .B2(n10481), .A(n10480), .ZN(n10487) );
  OAI21_X1 U11152 ( .B1(n10485), .B2(n10484), .A(n10483), .ZN(n10486) );
  AOI22_X1 U11153 ( .A1(n10487), .A2(n10505), .B1(n10504), .B2(n10486), .ZN(
        n10493) );
  NAND2_X1 U11154 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3151), .ZN(n10492)
         );
  AOI21_X1 U11155 ( .B1(n5026), .B2(n10489), .A(n10488), .ZN(n10490) );
  OR2_X1 U11156 ( .A1(n10490), .A2(n10511), .ZN(n10491) );
  NAND4_X1 U11157 ( .A1(n10494), .A2(n10493), .A3(n10492), .A4(n10491), .ZN(
        P2_U3192) );
  AOI22_X1 U11158 ( .A1(n10497), .A2(n10496), .B1(n10495), .B2(
        P2_ADDR_REG_11__SCAN_IN), .ZN(n10515) );
  OAI21_X1 U11159 ( .B1(P2_REG2_REG_11__SCAN_IN), .B2(n10499), .A(n10498), 
        .ZN(n10506) );
  OAI21_X1 U11160 ( .B1(n10502), .B2(n10501), .A(n10500), .ZN(n10503) );
  AOI22_X1 U11161 ( .A1(n10506), .A2(n10505), .B1(n10504), .B2(n10503), .ZN(
        n10514) );
  NAND2_X1 U11162 ( .A1(P2_REG3_REG_11__SCAN_IN), .A2(P2_U3151), .ZN(n10513)
         );
  AOI21_X1 U11163 ( .B1(n10509), .B2(n10508), .A(n10507), .ZN(n10510) );
  OR2_X1 U11164 ( .A1(n10511), .A2(n10510), .ZN(n10512) );
  NAND4_X1 U11165 ( .A1(n10515), .A2(n10514), .A3(n10513), .A4(n10512), .ZN(
        P2_U3193) );
  XOR2_X1 U11166 ( .A(n10516), .B(P1_RD_REG_SCAN_IN), .Z(U126) );
  INV_X1 U11167 ( .A(n10517), .ZN(n10518) );
  OAI211_X1 U11168 ( .C1(n10521), .C2(n10520), .A(n10519), .B(n10518), .ZN(
        n10531) );
  INV_X1 U11169 ( .A(n10522), .ZN(n10523) );
  OAI211_X1 U11170 ( .C1(n10526), .C2(n10525), .A(n10524), .B(n10523), .ZN(
        n10530) );
  NAND2_X1 U11171 ( .A1(n10528), .A2(n10527), .ZN(n10529) );
  AND3_X1 U11172 ( .A1(n10531), .A2(n10530), .A3(n10529), .ZN(n10536) );
  AOI211_X1 U11173 ( .C1(n10534), .C2(P1_ADDR_REG_4__SCAN_IN), .A(n10533), .B(
        n10532), .ZN(n10535) );
  NAND2_X1 U11174 ( .A1(n10536), .A2(n10535), .ZN(P1_U3247) );
  INV_X1 U11175 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n10537) );
  AOI22_X1 U11176 ( .A1(n10695), .A2(n10538), .B1(n10537), .B2(n10692), .ZN(
        P2_U3393) );
  INV_X1 U11177 ( .A(n10539), .ZN(n10627) );
  INV_X1 U11178 ( .A(n10540), .ZN(n10544) );
  OAI21_X1 U11179 ( .B1(n6965), .B2(n10162), .A(n10541), .ZN(n10543) );
  AOI211_X1 U11180 ( .C1(n10627), .C2(n10544), .A(n10543), .B(n10542), .ZN(
        n10547) );
  AOI22_X1 U11181 ( .A1(n10646), .A2(n10547), .B1(n10545), .B2(n10669), .ZN(
        P1_U3523) );
  INV_X1 U11182 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n10546) );
  AOI22_X1 U11183 ( .A1(n10674), .A2(n10547), .B1(n10546), .B2(n10671), .ZN(
        P1_U3456) );
  XNOR2_X1 U11184 ( .A(n10548), .B(n10549), .ZN(n10578) );
  INV_X1 U11185 ( .A(n10550), .ZN(n10554) );
  INV_X1 U11186 ( .A(n10551), .ZN(n10553) );
  OAI211_X1 U11187 ( .C1(n6971), .C2(n10554), .A(n10553), .B(n10552), .ZN(
        n10574) );
  OAI21_X1 U11188 ( .B1(n6971), .B2(n10162), .A(n10574), .ZN(n10566) );
  XNOR2_X1 U11189 ( .A(n10556), .B(n10555), .ZN(n10562) );
  AOI22_X1 U11190 ( .A1(n10559), .A2(n10558), .B1(n10557), .B2(n6960), .ZN(
        n10560) );
  OAI21_X1 U11191 ( .B1(n10562), .B2(n10561), .A(n10560), .ZN(n10563) );
  AOI21_X1 U11192 ( .B1(n10564), .B2(n10578), .A(n10563), .ZN(n10581) );
  INV_X1 U11193 ( .A(n10581), .ZN(n10565) );
  AOI211_X1 U11194 ( .C1(n10627), .C2(n10578), .A(n10566), .B(n10565), .ZN(
        n10569) );
  AOI22_X1 U11195 ( .A1(n10646), .A2(n10569), .B1(n10567), .B2(n10669), .ZN(
        P1_U3524) );
  INV_X1 U11196 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n10568) );
  AOI22_X1 U11197 ( .A1(n10674), .A2(n10569), .B1(n10568), .B2(n10671), .ZN(
        P1_U3459) );
  AOI222_X1 U11198 ( .A1(P1_REG2_REG_2__SCAN_IN), .A2(n4941), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(n10572), .C1(n10571), .C2(n10570), .ZN(
        n10580) );
  INV_X1 U11199 ( .A(n10573), .ZN(n10577) );
  INV_X1 U11200 ( .A(n10574), .ZN(n10575) );
  AOI22_X1 U11201 ( .A1(n10578), .A2(n10577), .B1(n10576), .B2(n10575), .ZN(
        n10579) );
  OAI211_X1 U11202 ( .C1(n4941), .C2(n10581), .A(n10580), .B(n10579), .ZN(
        P1_U3291) );
  INV_X1 U11203 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n10582) );
  AOI22_X1 U11204 ( .A1(n10695), .A2(n10583), .B1(n10582), .B2(n10692), .ZN(
        P2_U3396) );
  OAI22_X1 U11205 ( .A1(n10586), .A2(n10585), .B1(n10677), .B2(n10584), .ZN(
        n10589) );
  INV_X1 U11206 ( .A(n10587), .ZN(n10588) );
  AOI211_X1 U11207 ( .C1(n10590), .C2(n10683), .A(n10589), .B(n10588), .ZN(
        n10591) );
  AOI22_X1 U11208 ( .A1(n10687), .A2(n7241), .B1(n10591), .B2(n10641), .ZN(
        P2_U3231) );
  OAI21_X1 U11209 ( .B1(n10593), .B2(n10162), .A(n10592), .ZN(n10595) );
  AOI211_X1 U11210 ( .C1(n10667), .C2(n10596), .A(n10595), .B(n10594), .ZN(
        n10598) );
  AOI22_X1 U11211 ( .A1(n10646), .A2(n10598), .B1(n7406), .B2(n10669), .ZN(
        P1_U3525) );
  INV_X1 U11212 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n10597) );
  AOI22_X1 U11213 ( .A1(n10674), .A2(n10598), .B1(n10597), .B2(n10671), .ZN(
        P1_U3462) );
  INV_X1 U11214 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n10599) );
  AOI22_X1 U11215 ( .A1(n10695), .A2(n10600), .B1(n10599), .B2(n10692), .ZN(
        P2_U3399) );
  INV_X1 U11216 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n10601) );
  AOI22_X1 U11217 ( .A1(n10695), .A2(n10602), .B1(n10601), .B2(n10692), .ZN(
        P2_U3402) );
  INV_X1 U11218 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n10603) );
  AOI22_X1 U11219 ( .A1(n10695), .A2(n10604), .B1(n10603), .B2(n10692), .ZN(
        P2_U3405) );
  INV_X1 U11220 ( .A(n10605), .ZN(n10616) );
  OAI22_X1 U11221 ( .A1(n10609), .A2(n10608), .B1(n10607), .B2(n10606), .ZN(
        n10610) );
  AOI21_X1 U11222 ( .B1(P1_REG2_REG_5__SCAN_IN), .B2(n4941), .A(n10610), .ZN(
        n10611) );
  OAI21_X1 U11223 ( .B1(n10613), .B2(n10612), .A(n10611), .ZN(n10614) );
  AOI21_X1 U11224 ( .B1(n10616), .B2(n10615), .A(n10614), .ZN(n10617) );
  OAI21_X1 U11225 ( .B1(n4941), .B2(n10618), .A(n10617), .ZN(P1_U3288) );
  INV_X1 U11226 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10620) );
  AOI22_X1 U11227 ( .A1(n10695), .A2(n10621), .B1(n10620), .B2(n10692), .ZN(
        P2_U3408) );
  OAI21_X1 U11228 ( .B1(n10623), .B2(n10162), .A(n10622), .ZN(n10625) );
  AOI211_X1 U11229 ( .C1(n10627), .C2(n10626), .A(n10625), .B(n10624), .ZN(
        n10630) );
  INV_X1 U11230 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n10628) );
  AOI22_X1 U11231 ( .A1(n10646), .A2(n10630), .B1(n10628), .B2(n10669), .ZN(
        P1_U3528) );
  INV_X1 U11232 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n10629) );
  AOI22_X1 U11233 ( .A1(n10674), .A2(n10630), .B1(n10629), .B2(n10671), .ZN(
        P1_U3471) );
  INV_X1 U11234 ( .A(n10683), .ZN(n10633) );
  OAI21_X1 U11235 ( .B1(n10633), .B2(n10632), .A(n10631), .ZN(n10638) );
  AOI222_X1 U11236 ( .A1(n10641), .A2(n10638), .B1(n10637), .B2(n10636), .C1(
        n10635), .C2(n10634), .ZN(n10639) );
  OAI21_X1 U11237 ( .B1(n10641), .B2(n10640), .A(n10639), .ZN(P2_U3225) );
  OAI21_X1 U11238 ( .B1(n4946), .B2(n10162), .A(n10642), .ZN(n10644) );
  AOI211_X1 U11239 ( .C1(n10667), .C2(n10645), .A(n10644), .B(n10643), .ZN(
        n10648) );
  AOI22_X1 U11240 ( .A1(n10646), .A2(n10648), .B1(n7403), .B2(n10669), .ZN(
        P1_U3531) );
  INV_X1 U11241 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n10647) );
  AOI22_X1 U11242 ( .A1(n10674), .A2(n10648), .B1(n10647), .B2(n10671), .ZN(
        P1_U3480) );
  NAND2_X1 U11243 ( .A1(n4944), .A2(n10649), .ZN(n10651) );
  OAI211_X1 U11244 ( .C1(n10663), .C2(n10653), .A(n10652), .B(n10651), .ZN(
        n10654) );
  AOI21_X1 U11245 ( .B1(n10655), .B2(n10667), .A(n10654), .ZN(n10657) );
  AOI22_X1 U11246 ( .A1(n10646), .A2(n10657), .B1(n7402), .B2(n10669), .ZN(
        P1_U3532) );
  INV_X1 U11247 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n10656) );
  AOI22_X1 U11248 ( .A1(n10674), .A2(n10657), .B1(n10656), .B2(n10671), .ZN(
        P1_U3483) );
  INV_X1 U11249 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n10658) );
  AOI22_X1 U11250 ( .A1(n10695), .A2(n10659), .B1(n10658), .B2(n10692), .ZN(
        P2_U3420) );
  INV_X1 U11251 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n10660) );
  AOI22_X1 U11252 ( .A1(n10695), .A2(n10661), .B1(n10660), .B2(n10692), .ZN(
        P2_U3426) );
  OAI22_X1 U11253 ( .A1(n10664), .A2(n10663), .B1(n10662), .B2(n10162), .ZN(
        n10665) );
  AOI211_X1 U11254 ( .C1(n10668), .C2(n10667), .A(n10666), .B(n10665), .ZN(
        n10673) );
  AOI22_X1 U11255 ( .A1(n10646), .A2(n10673), .B1(n10670), .B2(n10669), .ZN(
        P1_U3534) );
  INV_X1 U11256 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n10672) );
  AOI22_X1 U11257 ( .A1(n10674), .A2(n10673), .B1(n10672), .B2(n10671), .ZN(
        P1_U3489) );
  INV_X1 U11258 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n10686) );
  INV_X1 U11259 ( .A(n10675), .ZN(n10680) );
  INV_X1 U11260 ( .A(n10676), .ZN(n10678) );
  OAI22_X1 U11261 ( .A1(n10680), .A2(n10679), .B1(n10678), .B2(n10677), .ZN(
        n10682) );
  AOI211_X1 U11262 ( .C1(n10684), .C2(n10683), .A(n10682), .B(n10681), .ZN(
        n10685) );
  AOI22_X1 U11263 ( .A1(n10687), .A2(n10686), .B1(n10685), .B2(n10641), .ZN(
        P2_U3220) );
  INV_X1 U11264 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n10688) );
  AOI22_X1 U11265 ( .A1(n10695), .A2(n10689), .B1(n10688), .B2(n10692), .ZN(
        P2_U3429) );
  INV_X1 U11266 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n10690) );
  AOI22_X1 U11267 ( .A1(n10695), .A2(n10691), .B1(n10690), .B2(n10692), .ZN(
        P2_U3432) );
  INV_X1 U11268 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n10693) );
  AOI22_X1 U11269 ( .A1(n10695), .A2(n10694), .B1(n10693), .B2(n10692), .ZN(
        P2_U3435) );
  XNOR2_X1 U11270 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  AND2_X1 U6424 ( .A1(n10280), .A2(n10283), .ZN(n5633) );
  NAND2_X1 U5032 ( .A1(n5807), .A2(n5568), .ZN(n5828) );
  XNOR2_X1 U5031 ( .A(n5828), .B(n5827), .ZN(n7668) );
  NAND2_X2 U5008 ( .A1(n5396), .A2(n5395), .ZN(n5528) );
  NAND2_X1 U5056 ( .A1(n7945), .A2(n6390), .ZN(n7981) );
endmodule

