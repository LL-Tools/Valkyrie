

module b17_C_AntiSAT_k_256_6 ( P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, 
        DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, 
        DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, 
        DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, 
        DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, 
        DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, 
        HOLD, NA, BS16, READY1, READY2, P1_READREQUEST_REG_SCAN_IN, 
        P1_ADS_N_REG_SCAN_IN, P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, 
        P1_D_C_N_REG_SCAN_IN, P1_REQUESTPENDING_REG_SCAN_IN, 
        P1_STATEBS16_REG_SCAN_IN, P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, 
        P1_W_R_N_REG_SCAN_IN, P1_BYTEENABLE_REG_0__SCAN_IN, 
        P1_BYTEENABLE_REG_1__SCAN_IN, P1_BYTEENABLE_REG_2__SCAN_IN, 
        P1_BYTEENABLE_REG_3__SCAN_IN, P1_REIP_REG_31__SCAN_IN, 
        P1_REIP_REG_30__SCAN_IN, P1_REIP_REG_29__SCAN_IN, 
        P1_REIP_REG_28__SCAN_IN, P1_REIP_REG_27__SCAN_IN, 
        P1_REIP_REG_26__SCAN_IN, P1_REIP_REG_25__SCAN_IN, 
        P1_REIP_REG_24__SCAN_IN, P1_REIP_REG_23__SCAN_IN, 
        P1_REIP_REG_22__SCAN_IN, P1_REIP_REG_21__SCAN_IN, 
        P1_REIP_REG_20__SCAN_IN, P1_REIP_REG_19__SCAN_IN, 
        P1_REIP_REG_18__SCAN_IN, P1_REIP_REG_17__SCAN_IN, 
        P1_REIP_REG_16__SCAN_IN, P1_REIP_REG_15__SCAN_IN, 
        P1_REIP_REG_14__SCAN_IN, P1_REIP_REG_13__SCAN_IN, 
        P1_REIP_REG_12__SCAN_IN, P1_REIP_REG_11__SCAN_IN, 
        P1_REIP_REG_10__SCAN_IN, P1_REIP_REG_9__SCAN_IN, 
        P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN, 
        P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, P1_REIP_REG_3__SCAN_IN, 
        P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN, 
        P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, P1_EBX_REG_29__SCAN_IN, 
        P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN, 
        P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, P1_EBX_REG_23__SCAN_IN, 
        P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN, 
        P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, P1_EBX_REG_17__SCAN_IN, 
        P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN, 
        P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, P1_EBX_REG_11__SCAN_IN, 
        P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, P1_EBX_REG_8__SCAN_IN, 
        P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, P1_EBX_REG_5__SCAN_IN, 
        P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, P1_EBX_REG_2__SCAN_IN, 
        P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, P1_EAX_REG_31__SCAN_IN, 
        P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN, 
        P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, P1_EAX_REG_25__SCAN_IN, 
        P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN, 
        P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, P1_EAX_REG_19__SCAN_IN, 
        P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN, 
        P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, P1_EAX_REG_13__SCAN_IN, 
        P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, 
        P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, 
        P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, 
        P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, 
        P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, 
        keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, 
        keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, 
        keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, 
        keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, 
        keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, 
        keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, 
        keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, 
        keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, 
        keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, 
        keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, 
        keyinput60, keyinput61, keyinput62, keyinput63, keyinput64, keyinput65, 
        keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, keyinput71, 
        keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, keyinput77, 
        keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, keyinput83, 
        keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, keyinput89, 
        keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, keyinput95, 
        keyinput96, keyinput97, keyinput98, keyinput99, keyinput100, 
        keyinput101, keyinput102, keyinput103, keyinput104, keyinput105, 
        keyinput106, keyinput107, keyinput108, keyinput109, keyinput110, 
        keyinput111, keyinput112, keyinput113, keyinput114, keyinput115, 
        keyinput116, keyinput117, keyinput118, keyinput119, keyinput120, 
        keyinput121, keyinput122, keyinput123, keyinput124, keyinput125, 
        keyinput126, keyinput127, keyinput128, keyinput129, keyinput130, 
        keyinput131, keyinput132, keyinput133, keyinput134, keyinput135, 
        keyinput136, keyinput137, keyinput138, keyinput139, keyinput140, 
        keyinput141, keyinput142, keyinput143, keyinput144, keyinput145, 
        keyinput146, keyinput147, keyinput148, keyinput149, keyinput150, 
        keyinput151, keyinput152, keyinput153, keyinput154, keyinput155, 
        keyinput156, keyinput157, keyinput158, keyinput159, keyinput160, 
        keyinput161, keyinput162, keyinput163, keyinput164, keyinput165, 
        keyinput166, keyinput167, keyinput168, keyinput169, keyinput170, 
        keyinput171, keyinput172, keyinput173, keyinput174, keyinput175, 
        keyinput176, keyinput177, keyinput178, keyinput179, keyinput180, 
        keyinput181, keyinput182, keyinput183, keyinput184, keyinput185, 
        keyinput186, keyinput187, keyinput188, keyinput189, keyinput190, 
        keyinput191, keyinput192, keyinput193, keyinput194, keyinput195, 
        keyinput196, keyinput197, keyinput198, keyinput199, keyinput200, 
        keyinput201, keyinput202, keyinput203, keyinput204, keyinput205, 
        keyinput206, keyinput207, keyinput208, keyinput209, keyinput210, 
        keyinput211, keyinput212, keyinput213, keyinput214, keyinput215, 
        keyinput216, keyinput217, keyinput218, keyinput219, keyinput220, 
        keyinput221, keyinput222, keyinput223, keyinput224, keyinput225, 
        keyinput226, keyinput227, keyinput228, keyinput229, keyinput230, 
        keyinput231, keyinput232, keyinput233, keyinput234, keyinput235, 
        keyinput236, keyinput237, keyinput238, keyinput239, keyinput240, 
        keyinput241, keyinput242, keyinput243, keyinput244, keyinput245, 
        keyinput246, keyinput247, keyinput248, keyinput249, keyinput250, 
        keyinput251, keyinput252, keyinput253, keyinput254, keyinput255, U355, 
        U356, U357, U358, U359, U360, U361, U362, U363, U364, U366, U367, U368, 
        U369, U370, U371, U372, U373, U374, U375, U347, U348, U349, U350, U351, 
        U352, U353, U354, U365, U376, U247, U246, U245, U244, U243, U242, U241, 
        U240, U239, U238, U237, U236, U235, U234, U233, U232, U231, U230, U229, 
        U228, U227, U226, U225, U224, U223, U222, U221, U220, U219, U218, U217, 
        U216, U251, U252, U253, U254, U255, U256, U257, U258, U259, U260, U261, 
        U262, U263, U264, U265, U266, U267, U268, U269, U270, U271, U272, U273, 
        U274, U275, U276, U277, U278, U279, U280, U281, U282, U212, U215, U213, 
        U214, P3_U3274, P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, 
        P3_U3059, P3_U3058, P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, 
        P3_U3052, P3_U3051, P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, 
        P3_U3045, P3_U3044, P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, 
        P3_U3038, P3_U3037, P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, 
        P3_U3031, P3_U3030, P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, 
        P3_U3026, P3_U3025, P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, 
        P3_U3019, P3_U3018, P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, 
        P3_U3012, P3_U3011, P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, 
        P3_U3005, P3_U3004, P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, 
        P3_U3282, P3_U2998, P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, 
        P3_U2992, P3_U2991, P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, 
        P3_U2985, P3_U2984, P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, 
        P3_U2978, P3_U2977, P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, 
        P3_U2971, P3_U2970, P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, 
        P3_U2964, P3_U2963, P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, 
        P3_U2957, P3_U2956, P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, 
        P3_U2950, P3_U2949, P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, 
        P3_U2943, P3_U2942, P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, 
        P3_U2936, P3_U2935, P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, 
        P3_U2929, P3_U2928, P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, 
        P3_U2922, P3_U2921, P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, 
        P3_U2915, P3_U2914, P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, 
        P3_U2908, P3_U2907, P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, 
        P3_U2901, P3_U2900, P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, 
        P3_U2894, P3_U2893, P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, 
        P3_U2887, P3_U2886, P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, 
        P3_U2880, P3_U2879, P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, 
        P3_U2873, P3_U2872, P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, 
        P3_U3285, P3_U3288, P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, 
        P3_U2864, P3_U2863, P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, 
        P3_U2857, P3_U2856, P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, 
        P3_U2850, P3_U2849, P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, 
        P3_U2843, P3_U2842, P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, 
        P3_U2836, P3_U2835, P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, 
        P3_U2829, P3_U2828, P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, 
        P3_U2822, P3_U2821, P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, 
        P3_U2815, P3_U2814, P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, 
        P3_U2808, P3_U2807, P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, 
        P3_U2801, P3_U2800, P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, 
        P3_U2794, P3_U2793, P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, 
        P3_U2787, P3_U2786, P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, 
        P3_U2780, P3_U2779, P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, 
        P3_U2773, P3_U2772, P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, 
        P3_U2766, P3_U2765, P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, 
        P3_U2759, P3_U2758, P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, 
        P3_U2752, P3_U2751, P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, 
        P3_U2745, P3_U2744, P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, 
        P3_U2738, P3_U2737, P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, 
        P3_U2731, P3_U2730, P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, 
        P3_U2724, P3_U2723, P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, 
        P3_U2717, P3_U2716, P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, 
        P3_U2710, P3_U2709, P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, 
        P3_U2703, P3_U2702, P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, 
        P3_U2696, P3_U2695, P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, 
        P3_U2689, P3_U2688, P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, 
        P3_U2682, P3_U2681, P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, 
        P3_U2675, P3_U2674, P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, 
        P3_U2668, P3_U2667, P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, 
        P3_U2661, P3_U2660, P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, 
        P3_U2654, P3_U2653, P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, 
        P3_U2647, P3_U2646, P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, 
        P3_U2640, P3_U2639, P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, 
        P3_U3295, P3_U2636, P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, 
        P3_U3298, P3_U3299, P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, 
        P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, 
        P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, 
        P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, 
        P2_U3179, P2_U3593, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, 
        P2_U3173, P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, 
        P2_U3166, P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, 
        P2_U3159, P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, 
        P2_U3152, P2_U3151, P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, 
        P2_U3145, P2_U3144, P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, 
        P2_U3138, P2_U3137, P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, 
        P2_U3131, P2_U3130, P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, 
        P2_U3124, P2_U3123, P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, 
        P2_U3117, P2_U3116, P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, 
        P2_U3110, P2_U3109, P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, 
        P2_U3103, P2_U3102, P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, 
        P2_U3096, P2_U3095, P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, 
        P2_U3089, P2_U3088, P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, 
        P2_U3082, P2_U3081, P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, 
        P2_U3075, P2_U3074, P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, 
        P2_U3068, P2_U3067, P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, 
        P2_U3061, P2_U3060, P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, 
        P2_U3054, P2_U3053, P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, 
        P2_U3595, P2_U3596, P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, 
        P2_U3603, P2_U3604, P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, 
        P2_U3042, P2_U3041, P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, 
        P2_U3035, P2_U3034, P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, 
        P2_U3028, P2_U3027, P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, 
        P2_U3021, P2_U3020, P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, 
        P2_U3014, P2_U3013, P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, 
        P2_U3007, P2_U3006, P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, 
        P2_U3000, P2_U2999, P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, 
        P2_U2993, P2_U2992, P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, 
        P2_U2986, P2_U2985, P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, 
        P2_U2979, P2_U2978, P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, 
        P2_U2972, P2_U2971, P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, 
        P2_U2965, P2_U2964, P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, 
        P2_U2958, P2_U2957, P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, 
        P2_U2951, P2_U2950, P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, 
        P2_U2944, P2_U2943, P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, 
        P2_U2937, P2_U2936, P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, 
        P2_U2930, P2_U2929, P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, 
        P2_U2923, P2_U2922, P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, 
        P2_U2916, P2_U2915, P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, 
        P2_U2909, P2_U2908, P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, 
        P2_U2902, P2_U2901, P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, 
        P2_U2895, P2_U2894, P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, 
        P2_U2888, P2_U2887, P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, 
        P2_U2881, P2_U2880, P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, 
        P2_U2874, P2_U2873, P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, 
        P2_U2867, P2_U2866, P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, 
        P2_U2860, P2_U2859, P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, 
        P2_U2853, P2_U2852, P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, 
        P2_U2846, P2_U2845, P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, 
        P2_U2839, P2_U2838, P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, 
        P2_U2832, P2_U2831, P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, 
        P2_U2825, P2_U2824, P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, 
        P2_U2819, P2_U3609, P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, 
        P2_U2815, P2_U3612, P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, 
        P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, 
        P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, 
        P1_U3212, P1_U3211, P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, 
        P1_U3205, P1_U3204, P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, 
        P1_U3198, P1_U3197, P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, 
        P1_U3193, P1_U3192, P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, 
        P1_U3186, P1_U3185, P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, 
        P1_U3179, P1_U3178, P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, 
        P1_U3172, P1_U3171, P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, 
        P1_U3165, P1_U3164, P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, 
        P1_U3159, P1_U3158, P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, 
        P1_U3152, P1_U3151, P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, 
        P1_U3145, P1_U3144, P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, 
        P1_U3138, P1_U3137, P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, 
        P1_U3131, P1_U3130, P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, 
        P1_U3124, P1_U3123, P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, 
        P1_U3117, P1_U3116, P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, 
        P1_U3110, P1_U3109, P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, 
        P1_U3103, P1_U3102, P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, 
        P1_U3096, P1_U3095, P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, 
        P1_U3089, P1_U3088, P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, 
        P1_U3082, P1_U3081, P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, 
        P1_U3075, P1_U3074, P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, 
        P1_U3068, P1_U3067, P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, 
        P1_U3061, P1_U3060, P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, 
        P1_U3054, P1_U3053, P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, 
        P1_U3047, P1_U3046, P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, 
        P1_U3040, P1_U3039, P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, 
        P1_U3033, P1_U3468, P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, 
        P1_U3475, P1_U3476, P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, 
        P1_U3028, P1_U3027, P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, 
        P1_U3021, P1_U3020, P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, 
        P1_U3014, P1_U3013, P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, 
        P1_U3007, P1_U3006, P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, 
        P1_U3000, P1_U2999, P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, 
        P1_U2993, P1_U2992, P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, 
        P1_U2986, P1_U2985, P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, 
        P1_U2979, P1_U2978, P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, 
        P1_U2972, P1_U2971, P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, 
        P1_U2965, P1_U2964, P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, 
        P1_U2958, P1_U2957, P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, 
        P1_U2951, P1_U2950, P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, 
        P1_U2944, P1_U2943, P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, 
        P1_U2937, P1_U2936, P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, 
        P1_U2930, P1_U2929, P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, 
        P1_U2923, P1_U2922, P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, 
        P1_U2916, P1_U2915, P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, 
        P1_U2909, P1_U2908, P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, 
        P1_U2902, P1_U2901, P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, 
        P1_U2895, P1_U2894, P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, 
        P1_U2888, P1_U2887, P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, 
        P1_U2881, P1_U2880, P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, 
        P1_U2874, P1_U2873, P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, 
        P1_U2867, P1_U2866, P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, 
        P1_U2860, P1_U2859, P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, 
        P1_U2853, P1_U2852, P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, 
        P1_U2846, P1_U2845, P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, 
        P1_U2839, P1_U2838, P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, 
        P1_U2832, P1_U2831, P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, 
        P1_U2825, P1_U2824, P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, 
        P1_U2818, P1_U2817, P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, 
        P1_U2811, P1_U2810, P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, 
        P1_U3483, P1_U2806, P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, 
        P1_U2803, P1_U2802, P1_U3487, P1_U2801 );
  input P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_,
         DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_,
         DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_,
         DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_,
         DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_,
         DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2,
         P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
         P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
         P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
         P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
         P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
         P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
         P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
         P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
         P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
         P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
         P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
         P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
         P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
         P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
         P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
         P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
         P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
         P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN,
         P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
         P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
         P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN,
         P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN,
         P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
         P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
         P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN,
         P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
         P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
         P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN,
         P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
         P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
         P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN,
         P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
         P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
         P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
         P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
         P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
         P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
         P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN,
         P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
         P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
         P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN,
         P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
         P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
         P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN,
         P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
         P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
         P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
         P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
         P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
         P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN, keyinput0, keyinput1, keyinput2,
         keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8,
         keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127, keyinput128, keyinput129,
         keyinput130, keyinput131, keyinput132, keyinput133, keyinput134,
         keyinput135, keyinput136, keyinput137, keyinput138, keyinput139,
         keyinput140, keyinput141, keyinput142, keyinput143, keyinput144,
         keyinput145, keyinput146, keyinput147, keyinput148, keyinput149,
         keyinput150, keyinput151, keyinput152, keyinput153, keyinput154,
         keyinput155, keyinput156, keyinput157, keyinput158, keyinput159,
         keyinput160, keyinput161, keyinput162, keyinput163, keyinput164,
         keyinput165, keyinput166, keyinput167, keyinput168, keyinput169,
         keyinput170, keyinput171, keyinput172, keyinput173, keyinput174,
         keyinput175, keyinput176, keyinput177, keyinput178, keyinput179,
         keyinput180, keyinput181, keyinput182, keyinput183, keyinput184,
         keyinput185, keyinput186, keyinput187, keyinput188, keyinput189,
         keyinput190, keyinput191, keyinput192, keyinput193, keyinput194,
         keyinput195, keyinput196, keyinput197, keyinput198, keyinput199,
         keyinput200, keyinput201, keyinput202, keyinput203, keyinput204,
         keyinput205, keyinput206, keyinput207, keyinput208, keyinput209,
         keyinput210, keyinput211, keyinput212, keyinput213, keyinput214,
         keyinput215, keyinput216, keyinput217, keyinput218, keyinput219,
         keyinput220, keyinput221, keyinput222, keyinput223, keyinput224,
         keyinput225, keyinput226, keyinput227, keyinput228, keyinput229,
         keyinput230, keyinput231, keyinput232, keyinput233, keyinput234,
         keyinput235, keyinput236, keyinput237, keyinput238, keyinput239,
         keyinput240, keyinput241, keyinput242, keyinput243, keyinput244,
         keyinput245, keyinput246, keyinput247, keyinput248, keyinput249,
         keyinput250, keyinput251, keyinput252, keyinput253, keyinput254,
         keyinput255;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9837, n9838,
         n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848,
         n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858,
         n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868,
         n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878,
         n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888,
         n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898,
         n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908,
         n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918,
         n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928,
         n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938,
         n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948,
         n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958,
         n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968,
         n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978,
         n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988,
         n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998,
         n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
         n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
         n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
         n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
         n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
         n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
         n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247,
         n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255,
         n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263,
         n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271,
         n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279,
         n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287,
         n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295,
         n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303,
         n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311,
         n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319,
         n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327,
         n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335,
         n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343,
         n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351,
         n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359,
         n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367,
         n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375,
         n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383,
         n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391,
         n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399,
         n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407,
         n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415,
         n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423,
         n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431,
         n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439,
         n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447,
         n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455,
         n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463,
         n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471,
         n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479,
         n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487,
         n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495,
         n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503,
         n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511,
         n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519,
         n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527,
         n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535,
         n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543,
         n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551,
         n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559,
         n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567,
         n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575,
         n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583,
         n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591,
         n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599,
         n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607,
         n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10615,
         n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623,
         n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631,
         n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639,
         n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647,
         n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655,
         n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663,
         n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671,
         n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679,
         n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687,
         n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695,
         n10696, n10697, n10698, n10699, n10700, n10701, n10702, n10703,
         n10704, n10705, n10706, n10707, n10708, n10709, n10710, n10711,
         n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719,
         n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727,
         n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735,
         n10736, n10737, n10738, n10739, n10740, n10741, n10742, n10743,
         n10744, n10745, n10746, n10747, n10748, n10749, n10750, n10751,
         n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759,
         n10760, n10761, n10762, n10763, n10764, n10765, n10766, n10767,
         n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10775,
         n10776, n10777, n10778, n10779, n10780, n10781, n10782, n10783,
         n10784, n10785, n10786, n10787, n10788, n10789, n10790, n10791,
         n10792, n10793, n10794, n10795, n10796, n10797, n10798, n10799,
         n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807,
         n10808, n10809, n10810, n10811, n10812, n10813, n10814, n10815,
         n10816, n10817, n10818, n10819, n10820, n10821, n10822, n10823,
         n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831,
         n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839,
         n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847,
         n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10855,
         n10856, n10857, n10858, n10859, n10860, n10861, n10862, n10863,
         n10864, n10865, n10866, n10867, n10868, n10869, n10870, n10871,
         n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879,
         n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887,
         n10888, n10889, n10890, n10891, n10892, n10893, n10894, n10895,
         n10896, n10897, n10898, n10899, n10900, n10901, n10902, n10903,
         n10904, n10905, n10906, n10907, n10908, n10909, n10910, n10911,
         n10912, n10913, n10914, n10915, n10916, n10917, n10918, n10919,
         n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927,
         n10928, n10929, n10930, n10931, n10932, n10933, n10934, n10935,
         n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10943,
         n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10951,
         n10952, n10953, n10954, n10955, n10956, n10957, n10958, n10959,
         n10960, n10961, n10962, n10963, n10964, n10965, n10966, n10967,
         n10968, n10969, n10970, n10971, n10972, n10973, n10974, n10975,
         n10976, n10977, n10978, n10979, n10980, n10981, n10982, n10983,
         n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991,
         n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999,
         n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007,
         n11008, n11009, n11010, n11011, n11012, n11013, n11014, n11015,
         n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023,
         n11024, n11025, n11026, n11027, n11028, n11029, n11030, n11031,
         n11032, n11033, n11034, n11035, n11036, n11037, n11038, n11039,
         n11040, n11041, n11042, n11043, n11044, n11045, n11046, n11047,
         n11048, n11049, n11050, n11051, n11052, n11053, n11054, n11055,
         n11056, n11057, n11058, n11059, n11060, n11061, n11062, n11063,
         n11064, n11065, n11066, n11067, n11068, n11069, n11070, n11071,
         n11072, n11073, n11074, n11075, n11076, n11077, n11078, n11079,
         n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087,
         n11088, n11089, n11090, n11091, n11092, n11093, n11094, n11095,
         n11096, n11097, n11098, n11099, n11100, n11101, n11102, n11103,
         n11104, n11105, n11106, n11107, n11108, n11109, n11110, n11111,
         n11112, n11113, n11114, n11115, n11116, n11117, n11118, n11119,
         n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11127,
         n11128, n11129, n11130, n11131, n11132, n11133, n11134, n11135,
         n11136, n11137, n11138, n11139, n11140, n11141, n11142, n11143,
         n11144, n11145, n11146, n11147, n11148, n11149, n11150, n11151,
         n11152, n11153, n11154, n11155, n11156, n11157, n11158, n11159,
         n11160, n11161, n11162, n11163, n11164, n11165, n11166, n11167,
         n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11175,
         n11176, n11177, n11178, n11179, n11180, n11181, n11182, n11183,
         n11184, n11185, n11186, n11187, n11188, n11189, n11190, n11191,
         n11192, n11193, n11194, n11195, n11196, n11197, n11198, n11199,
         n11200, n11201, n11202, n11203, n11204, n11205, n11206, n11207,
         n11208, n11209, n11210, n11211, n11212, n11213, n11214, n11215,
         n11216, n11217, n11218, n11219, n11220, n11221, n11222, n11223,
         n11224, n11225, n11226, n11227, n11228, n11229, n11230, n11231,
         n11232, n11233, n11234, n11235, n11236, n11237, n11238, n11239,
         n11240, n11241, n11242, n11243, n11244, n11245, n11246, n11247,
         n11248, n11249, n11250, n11251, n11252, n11253, n11254, n11255,
         n11256, n11257, n11258, n11259, n11260, n11261, n11262, n11263,
         n11264, n11265, n11266, n11267, n11268, n11269, n11270, n11271,
         n11272, n11273, n11274, n11275, n11276, n11277, n11278, n11279,
         n11280, n11281, n11282, n11283, n11284, n11285, n11286, n11287,
         n11288, n11289, n11290, n11291, n11292, n11293, n11294, n11295,
         n11296, n11297, n11298, n11299, n11300, n11301, n11302, n11303,
         n11304, n11305, n11306, n11307, n11308, n11309, n11310, n11311,
         n11312, n11313, n11314, n11315, n11316, n11317, n11318, n11319,
         n11320, n11321, n11322, n11323, n11324, n11325, n11326, n11327,
         n11328, n11329, n11330, n11331, n11332, n11333, n11334, n11335,
         n11336, n11337, n11338, n11339, n11340, n11341, n11342, n11343,
         n11344, n11345, n11346, n11347, n11348, n11349, n11350, n11351,
         n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359,
         n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367,
         n11368, n11369, n11370, n11371, n11372, n11373, n11374, n11375,
         n11376, n11377, n11378, n11379, n11380, n11381, n11382, n11383,
         n11384, n11385, n11386, n11387, n11388, n11389, n11390, n11391,
         n11392, n11393, n11394, n11395, n11396, n11397, n11398, n11399,
         n11400, n11401, n11402, n11403, n11404, n11405, n11406, n11407,
         n11408, n11409, n11410, n11411, n11412, n11413, n11414, n11415,
         n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423,
         n11424, n11425, n11426, n11427, n11428, n11429, n11430, n11431,
         n11432, n11433, n11434, n11435, n11436, n11437, n11438, n11439,
         n11440, n11441, n11442, n11443, n11444, n11445, n11446, n11447,
         n11448, n11449, n11450, n11451, n11452, n11453, n11454, n11455,
         n11456, n11457, n11458, n11459, n11460, n11461, n11462, n11463,
         n11464, n11465, n11466, n11467, n11468, n11469, n11470, n11471,
         n11472, n11473, n11474, n11475, n11476, n11477, n11478, n11479,
         n11480, n11481, n11482, n11483, n11484, n11485, n11486, n11487,
         n11488, n11489, n11490, n11491, n11492, n11493, n11494, n11495,
         n11496, n11497, n11498, n11499, n11500, n11501, n11502, n11503,
         n11504, n11505, n11506, n11507, n11508, n11509, n11510, n11511,
         n11512, n11513, n11514, n11515, n11516, n11517, n11518, n11519,
         n11520, n11521, n11522, n11523, n11524, n11525, n11526, n11527,
         n11528, n11529, n11530, n11531, n11532, n11533, n11534, n11535,
         n11536, n11537, n11538, n11539, n11540, n11541, n11542, n11543,
         n11544, n11545, n11546, n11547, n11548, n11549, n11550, n11551,
         n11552, n11553, n11554, n11555, n11556, n11557, n11558, n11559,
         n11560, n11561, n11562, n11563, n11564, n11565, n11566, n11567,
         n11568, n11569, n11570, n11571, n11572, n11573, n11574, n11575,
         n11576, n11577, n11578, n11579, n11580, n11581, n11582, n11583,
         n11584, n11585, n11586, n11587, n11588, n11589, n11590, n11591,
         n11592, n11593, n11594, n11595, n11596, n11597, n11598, n11599,
         n11600, n11601, n11602, n11603, n11604, n11605, n11606, n11607,
         n11608, n11609, n11610, n11611, n11612, n11613, n11614, n11615,
         n11616, n11617, n11618, n11619, n11620, n11621, n11622, n11623,
         n11624, n11625, n11626, n11627, n11628, n11629, n11630, n11631,
         n11632, n11633, n11634, n11635, n11636, n11637, n11638, n11639,
         n11640, n11641, n11642, n11643, n11644, n11645, n11646, n11647,
         n11648, n11649, n11650, n11651, n11652, n11653, n11654, n11655,
         n11656, n11657, n11658, n11659, n11660, n11661, n11662, n11663,
         n11664, n11665, n11666, n11667, n11668, n11669, n11670, n11671,
         n11672, n11673, n11674, n11675, n11676, n11677, n11678, n11679,
         n11680, n11681, n11682, n11683, n11684, n11685, n11686, n11687,
         n11688, n11689, n11690, n11691, n11692, n11693, n11694, n11695,
         n11696, n11697, n11698, n11699, n11700, n11701, n11702, n11703,
         n11704, n11705, n11706, n11707, n11708, n11709, n11710, n11711,
         n11712, n11713, n11714, n11715, n11716, n11717, n11718, n11719,
         n11720, n11721, n11722, n11723, n11724, n11725, n11726, n11727,
         n11728, n11729, n11730, n11731, n11732, n11733, n11734, n11735,
         n11736, n11737, n11738, n11739, n11740, n11741, n11742, n11743,
         n11744, n11745, n11746, n11747, n11748, n11749, n11750, n11751,
         n11752, n11753, n11754, n11755, n11756, n11757, n11758, n11759,
         n11760, n11761, n11762, n11763, n11764, n11765, n11766, n11767,
         n11768, n11769, n11770, n11771, n11772, n11773, n11774, n11775,
         n11776, n11777, n11778, n11779, n11780, n11781, n11782, n11783,
         n11784, n11785, n11786, n11787, n11788, n11789, n11790, n11791,
         n11792, n11793, n11794, n11795, n11796, n11797, n11798, n11799,
         n11800, n11801, n11802, n11803, n11804, n11805, n11806, n11807,
         n11808, n11809, n11810, n11811, n11812, n11813, n11814, n11815,
         n11816, n11817, n11818, n11819, n11820, n11821, n11822, n11823,
         n11824, n11825, n11826, n11827, n11828, n11829, n11830, n11831,
         n11832, n11833, n11834, n11835, n11836, n11837, n11838, n11839,
         n11840, n11841, n11842, n11843, n11844, n11845, n11846, n11847,
         n11848, n11849, n11850, n11851, n11852, n11853, n11854, n11855,
         n11856, n11857, n11858, n11859, n11860, n11861, n11862, n11863,
         n11864, n11865, n11866, n11867, n11868, n11869, n11870, n11871,
         n11872, n11873, n11874, n11875, n11876, n11877, n11878, n11879,
         n11880, n11881, n11882, n11883, n11884, n11885, n11886, n11887,
         n11888, n11889, n11890, n11891, n11892, n11893, n11894, n11895,
         n11896, n11897, n11898, n11899, n11900, n11901, n11902, n11903,
         n11904, n11905, n11906, n11907, n11908, n11909, n11910, n11911,
         n11912, n11913, n11914, n11915, n11916, n11917, n11918, n11919,
         n11920, n11921, n11922, n11923, n11924, n11925, n11926, n11927,
         n11928, n11929, n11930, n11931, n11932, n11933, n11934, n11935,
         n11936, n11937, n11938, n11939, n11940, n11941, n11942, n11943,
         n11944, n11945, n11946, n11947, n11948, n11949, n11950, n11951,
         n11952, n11953, n11954, n11955, n11956, n11957, n11958, n11959,
         n11960, n11961, n11962, n11963, n11964, n11965, n11966, n11967,
         n11968, n11969, n11970, n11971, n11972, n11973, n11974, n11975,
         n11976, n11977, n11978, n11979, n11980, n11981, n11982, n11983,
         n11984, n11985, n11986, n11987, n11988, n11989, n11990, n11991,
         n11992, n11993, n11994, n11995, n11996, n11997, n11998, n11999,
         n12000, n12001, n12002, n12003, n12004, n12005, n12006, n12007,
         n12008, n12009, n12010, n12011, n12012, n12013, n12014, n12015,
         n12016, n12017, n12018, n12019, n12020, n12021, n12022, n12023,
         n12024, n12025, n12026, n12027, n12028, n12029, n12030, n12031,
         n12032, n12033, n12034, n12035, n12036, n12037, n12038, n12039,
         n12040, n12041, n12042, n12043, n12044, n12045, n12046, n12047,
         n12048, n12049, n12050, n12051, n12052, n12053, n12054, n12055,
         n12056, n12057, n12058, n12059, n12060, n12061, n12062, n12063,
         n12064, n12065, n12066, n12067, n12068, n12069, n12070, n12071,
         n12072, n12073, n12074, n12075, n12076, n12077, n12078, n12079,
         n12080, n12081, n12082, n12083, n12084, n12085, n12086, n12087,
         n12088, n12089, n12090, n12091, n12092, n12093, n12094, n12095,
         n12096, n12097, n12098, n12099, n12100, n12101, n12102, n12103,
         n12104, n12105, n12106, n12107, n12108, n12109, n12110, n12111,
         n12112, n12113, n12114, n12115, n12116, n12117, n12118, n12119,
         n12120, n12121, n12122, n12123, n12124, n12125, n12126, n12127,
         n12128, n12129, n12130, n12131, n12132, n12133, n12134, n12135,
         n12136, n12137, n12138, n12139, n12140, n12141, n12142, n12143,
         n12144, n12145, n12146, n12147, n12148, n12149, n12150, n12151,
         n12152, n12153, n12154, n12155, n12156, n12157, n12158, n12159,
         n12160, n12161, n12162, n12163, n12164, n12165, n12166, n12167,
         n12168, n12169, n12170, n12171, n12172, n12173, n12174, n12175,
         n12176, n12177, n12178, n12179, n12180, n12181, n12182, n12183,
         n12184, n12185, n12186, n12187, n12188, n12189, n12190, n12191,
         n12192, n12193, n12194, n12195, n12196, n12197, n12198, n12199,
         n12200, n12201, n12202, n12203, n12204, n12205, n12206, n12207,
         n12208, n12209, n12210, n12211, n12212, n12213, n12214, n12215,
         n12216, n12217, n12218, n12219, n12220, n12221, n12222, n12223,
         n12224, n12225, n12226, n12227, n12228, n12229, n12230, n12231,
         n12232, n12233, n12234, n12235, n12236, n12237, n12238, n12239,
         n12240, n12241, n12242, n12243, n12244, n12245, n12246, n12247,
         n12248, n12249, n12250, n12251, n12252, n12253, n12254, n12255,
         n12256, n12257, n12258, n12259, n12260, n12261, n12262, n12263,
         n12264, n12265, n12266, n12267, n12268, n12269, n12270, n12271,
         n12272, n12273, n12274, n12275, n12276, n12277, n12278, n12279,
         n12280, n12281, n12282, n12283, n12284, n12285, n12286, n12287,
         n12288, n12289, n12290, n12291, n12292, n12293, n12294, n12295,
         n12296, n12297, n12298, n12299, n12300, n12301, n12302, n12303,
         n12304, n12305, n12306, n12307, n12308, n12309, n12310, n12311,
         n12312, n12313, n12314, n12315, n12316, n12317, n12318, n12319,
         n12320, n12321, n12322, n12323, n12324, n12325, n12326, n12327,
         n12328, n12329, n12330, n12331, n12332, n12333, n12334, n12335,
         n12336, n12337, n12338, n12339, n12340, n12341, n12342, n12343,
         n12344, n12345, n12346, n12347, n12348, n12349, n12350, n12351,
         n12352, n12353, n12354, n12355, n12356, n12357, n12358, n12359,
         n12360, n12361, n12362, n12363, n12364, n12365, n12366, n12367,
         n12368, n12369, n12370, n12371, n12372, n12373, n12374, n12375,
         n12376, n12377, n12378, n12379, n12380, n12381, n12382, n12383,
         n12384, n12385, n12386, n12387, n12388, n12389, n12390, n12391,
         n12392, n12393, n12394, n12395, n12396, n12397, n12398, n12399,
         n12400, n12401, n12402, n12403, n12404, n12405, n12406, n12407,
         n12408, n12409, n12410, n12411, n12412, n12413, n12414, n12415,
         n12416, n12417, n12418, n12419, n12420, n12421, n12422, n12423,
         n12424, n12425, n12426, n12427, n12428, n12429, n12430, n12431,
         n12432, n12433, n12434, n12435, n12436, n12437, n12438, n12439,
         n12440, n12441, n12442, n12443, n12444, n12445, n12446, n12447,
         n12448, n12449, n12450, n12451, n12452, n12453, n12454, n12455,
         n12456, n12457, n12458, n12459, n12460, n12461, n12462, n12463,
         n12464, n12465, n12466, n12467, n12468, n12469, n12470, n12471,
         n12472, n12473, n12474, n12475, n12476, n12477, n12478, n12479,
         n12480, n12481, n12482, n12483, n12484, n12485, n12486, n12487,
         n12488, n12489, n12490, n12491, n12492, n12493, n12494, n12495,
         n12496, n12497, n12498, n12499, n12500, n12501, n12502, n12503,
         n12504, n12505, n12506, n12507, n12508, n12509, n12510, n12511,
         n12512, n12513, n12514, n12515, n12516, n12517, n12518, n12519,
         n12520, n12521, n12522, n12523, n12524, n12525, n12526, n12527,
         n12528, n12529, n12530, n12531, n12532, n12533, n12534, n12535,
         n12536, n12537, n12538, n12539, n12540, n12541, n12542, n12543,
         n12544, n12545, n12546, n12547, n12548, n12549, n12550, n12551,
         n12552, n12553, n12554, n12555, n12556, n12557, n12558, n12559,
         n12560, n12561, n12562, n12563, n12564, n12565, n12566, n12567,
         n12568, n12569, n12570, n12571, n12572, n12573, n12574, n12575,
         n12576, n12577, n12578, n12579, n12580, n12581, n12582, n12583,
         n12584, n12585, n12586, n12587, n12588, n12589, n12590, n12591,
         n12592, n12593, n12594, n12595, n12596, n12597, n12598, n12599,
         n12600, n12601, n12602, n12603, n12604, n12605, n12606, n12607,
         n12608, n12609, n12610, n12611, n12612, n12613, n12614, n12615,
         n12616, n12617, n12618, n12619, n12620, n12621, n12622, n12623,
         n12624, n12625, n12626, n12627, n12628, n12629, n12630, n12631,
         n12632, n12633, n12634, n12635, n12636, n12637, n12638, n12639,
         n12640, n12641, n12642, n12643, n12644, n12645, n12646, n12647,
         n12648, n12649, n12650, n12651, n12652, n12653, n12654, n12655,
         n12656, n12657, n12658, n12659, n12660, n12661, n12662, n12663,
         n12664, n12665, n12666, n12667, n12668, n12669, n12670, n12671,
         n12672, n12673, n12674, n12675, n12676, n12677, n12678, n12679,
         n12680, n12681, n12682, n12683, n12684, n12685, n12686, n12687,
         n12688, n12689, n12690, n12691, n12692, n12693, n12694, n12695,
         n12696, n12697, n12698, n12699, n12700, n12701, n12702, n12703,
         n12704, n12705, n12706, n12707, n12708, n12709, n12710, n12711,
         n12712, n12713, n12714, n12715, n12716, n12717, n12718, n12719,
         n12720, n12721, n12722, n12723, n12724, n12725, n12726, n12727,
         n12728, n12729, n12730, n12731, n12732, n12733, n12734, n12735,
         n12736, n12737, n12738, n12739, n12740, n12741, n12742, n12743,
         n12744, n12745, n12746, n12747, n12748, n12749, n12750, n12751,
         n12752, n12753, n12754, n12755, n12756, n12757, n12758, n12759,
         n12760, n12761, n12762, n12763, n12764, n12765, n12766, n12767,
         n12768, n12769, n12770, n12771, n12772, n12773, n12774, n12775,
         n12776, n12777, n12778, n12779, n12780, n12781, n12782, n12783,
         n12784, n12785, n12786, n12787, n12788, n12789, n12791, n12792,
         n12793, n12794, n12795, n12796, n12797, n12798, n12799, n12800,
         n12801, n12802, n12803, n12804, n12805, n12806, n12807, n12808,
         n12809, n12810, n12811, n12812, n12813, n12814, n12815, n12816,
         n12817, n12818, n12819, n12820, n12821, n12822, n12823, n12824,
         n12825, n12826, n12827, n12828, n12829, n12830, n12831, n12832,
         n12833, n12834, n12835, n12836, n12837, n12838, n12839, n12840,
         n12841, n12842, n12843, n12844, n12845, n12846, n12847, n12848,
         n12849, n12850, n12851, n12852, n12853, n12854, n12855, n12856,
         n12857, n12858, n12859, n12860, n12861, n12862, n12863, n12864,
         n12865, n12866, n12867, n12868, n12869, n12870, n12871, n12872,
         n12873, n12874, n12875, n12876, n12877, n12878, n12879, n12880,
         n12881, n12882, n12883, n12884, n12885, n12886, n12887, n12888,
         n12889, n12890, n12891, n12892, n12893, n12894, n12895, n12896,
         n12897, n12898, n12899, n12900, n12901, n12902, n12903, n12904,
         n12905, n12906, n12907, n12908, n12909, n12910, n12911, n12912,
         n12913, n12914, n12915, n12916, n12917, n12918, n12919, n12920,
         n12921, n12922, n12923, n12924, n12925, n12926, n12927, n12928,
         n12929, n12930, n12931, n12932, n12933, n12934, n12935, n12936,
         n12937, n12938, n12939, n12940, n12941, n12942, n12943, n12944,
         n12945, n12946, n12947, n12948, n12949, n12950, n12951, n12952,
         n12953, n12954, n12955, n12956, n12957, n12958, n12959, n12960,
         n12961, n12962, n12963, n12964, n12965, n12966, n12967, n12968,
         n12969, n12970, n12971, n12972, n12973, n12974, n12975, n12976,
         n12977, n12978, n12979, n12980, n12981, n12982, n12983, n12984,
         n12985, n12986, n12987, n12988, n12989, n12990, n12991, n12992,
         n12993, n12994, n12995, n12996, n12997, n12998, n12999, n13000,
         n13001, n13002, n13003, n13004, n13005, n13006, n13007, n13008,
         n13009, n13010, n13011, n13012, n13013, n13014, n13015, n13016,
         n13017, n13018, n13019, n13020, n13021, n13022, n13023, n13024,
         n13025, n13026, n13027, n13028, n13029, n13030, n13031, n13032,
         n13033, n13034, n13035, n13036, n13037, n13038, n13039, n13040,
         n13041, n13042, n13043, n13044, n13045, n13046, n13047, n13048,
         n13049, n13050, n13051, n13052, n13053, n13054, n13055, n13056,
         n13057, n13058, n13059, n13060, n13061, n13062, n13063, n13064,
         n13065, n13066, n13067, n13068, n13069, n13070, n13071, n13072,
         n13073, n13074, n13075, n13076, n13077, n13078, n13079, n13080,
         n13081, n13082, n13083, n13084, n13085, n13086, n13087, n13088,
         n13089, n13090, n13091, n13092, n13093, n13094, n13095, n13096,
         n13097, n13098, n13099, n13100, n13101, n13102, n13103, n13104,
         n13105, n13106, n13107, n13108, n13109, n13110, n13111, n13112,
         n13113, n13114, n13115, n13116, n13117, n13118, n13119, n13120,
         n13121, n13122, n13123, n13124, n13125, n13126, n13127, n13128,
         n13129, n13130, n13131, n13132, n13133, n13134, n13135, n13136,
         n13137, n13138, n13139, n13140, n13141, n13142, n13143, n13144,
         n13145, n13146, n13147, n13148, n13149, n13150, n13151, n13152,
         n13153, n13154, n13155, n13156, n13157, n13158, n13159, n13160,
         n13161, n13162, n13163, n13164, n13165, n13166, n13167, n13168,
         n13169, n13170, n13171, n13172, n13173, n13174, n13175, n13176,
         n13177, n13178, n13179, n13180, n13181, n13182, n13183, n13184,
         n13185, n13186, n13187, n13188, n13189, n13190, n13191, n13192,
         n13193, n13194, n13195, n13196, n13197, n13198, n13199, n13200,
         n13201, n13202, n13203, n13204, n13205, n13206, n13207, n13208,
         n13209, n13210, n13211, n13212, n13213, n13214, n13215, n13216,
         n13217, n13218, n13219, n13220, n13221, n13222, n13223, n13224,
         n13225, n13226, n13227, n13228, n13229, n13230, n13231, n13232,
         n13233, n13234, n13235, n13236, n13237, n13238, n13239, n13240,
         n13241, n13242, n13243, n13244, n13245, n13246, n13247, n13248,
         n13249, n13250, n13251, n13252, n13253, n13254, n13255, n13256,
         n13257, n13258, n13259, n13260, n13261, n13262, n13263, n13264,
         n13265, n13266, n13267, n13268, n13269, n13270, n13271, n13272,
         n13273, n13274, n13275, n13276, n13277, n13278, n13279, n13280,
         n13281, n13282, n13283, n13284, n13285, n13286, n13287, n13288,
         n13289, n13290, n13291, n13292, n13293, n13294, n13295, n13296,
         n13297, n13298, n13299, n13300, n13301, n13302, n13303, n13304,
         n13305, n13306, n13307, n13308, n13309, n13310, n13311, n13312,
         n13313, n13314, n13315, n13316, n13317, n13318, n13319, n13320,
         n13321, n13322, n13323, n13324, n13325, n13326, n13327, n13328,
         n13329, n13330, n13331, n13332, n13333, n13334, n13335, n13336,
         n13337, n13338, n13339, n13340, n13341, n13342, n13343, n13344,
         n13345, n13346, n13347, n13348, n13349, n13350, n13351, n13352,
         n13353, n13354, n13355, n13356, n13357, n13358, n13359, n13360,
         n13361, n13362, n13363, n13364, n13365, n13366, n13367, n13368,
         n13369, n13370, n13371, n13372, n13373, n13374, n13375, n13376,
         n13377, n13378, n13379, n13380, n13381, n13382, n13383, n13384,
         n13385, n13386, n13387, n13388, n13389, n13390, n13391, n13392,
         n13393, n13394, n13395, n13396, n13397, n13398, n13399, n13400,
         n13401, n13402, n13403, n13404, n13405, n13406, n13407, n13408,
         n13409, n13410, n13411, n13412, n13413, n13414, n13415, n13416,
         n13417, n13418, n13419, n13420, n13421, n13422, n13423, n13424,
         n13425, n13426, n13427, n13428, n13429, n13430, n13431, n13432,
         n13433, n13434, n13435, n13436, n13437, n13438, n13439, n13440,
         n13441, n13442, n13443, n13444, n13445, n13446, n13447, n13448,
         n13449, n13450, n13451, n13452, n13453, n13454, n13455, n13456,
         n13457, n13458, n13459, n13460, n13461, n13462, n13463, n13464,
         n13465, n13466, n13467, n13468, n13469, n13470, n13471, n13472,
         n13473, n13474, n13475, n13476, n13477, n13478, n13479, n13480,
         n13481, n13482, n13483, n13484, n13485, n13486, n13487, n13488,
         n13489, n13490, n13491, n13492, n13493, n13494, n13495, n13496,
         n13497, n13498, n13499, n13500, n13501, n13502, n13503, n13504,
         n13505, n13506, n13507, n13508, n13509, n13510, n13511, n13512,
         n13513, n13514, n13515, n13516, n13517, n13518, n13519, n13520,
         n13521, n13522, n13523, n13524, n13525, n13526, n13527, n13528,
         n13529, n13530, n13531, n13532, n13533, n13534, n13535, n13536,
         n13537, n13538, n13539, n13540, n13541, n13542, n13543, n13544,
         n13545, n13546, n13547, n13548, n13549, n13550, n13551, n13552,
         n13553, n13554, n13555, n13556, n13557, n13558, n13559, n13560,
         n13561, n13562, n13563, n13564, n13565, n13566, n13567, n13568,
         n13569, n13570, n13571, n13572, n13573, n13574, n13575, n13576,
         n13577, n13578, n13579, n13580, n13581, n13582, n13583, n13584,
         n13585, n13586, n13587, n13588, n13589, n13590, n13591, n13592,
         n13593, n13594, n13595, n13596, n13597, n13598, n13599, n13600,
         n13601, n13602, n13603, n13604, n13605, n13606, n13607, n13608,
         n13609, n13610, n13611, n13612, n13613, n13614, n13615, n13616,
         n13617, n13618, n13619, n13620, n13621, n13622, n13623, n13624,
         n13625, n13626, n13627, n13628, n13629, n13630, n13631, n13632,
         n13633, n13634, n13635, n13636, n13637, n13638, n13639, n13640,
         n13641, n13642, n13643, n13644, n13645, n13646, n13647, n13648,
         n13649, n13650, n13651, n13652, n13653, n13654, n13655, n13656,
         n13657, n13658, n13659, n13660, n13661, n13662, n13663, n13664,
         n13665, n13666, n13667, n13668, n13669, n13670, n13671, n13672,
         n13673, n13674, n13675, n13676, n13677, n13678, n13679, n13680,
         n13681, n13682, n13683, n13684, n13685, n13686, n13687, n13688,
         n13689, n13690, n13691, n13692, n13693, n13694, n13695, n13696,
         n13697, n13698, n13699, n13700, n13701, n13702, n13703, n13704,
         n13705, n13706, n13707, n13708, n13709, n13710, n13711, n13712,
         n13713, n13714, n13715, n13716, n13717, n13718, n13719, n13720,
         n13721, n13722, n13723, n13724, n13725, n13726, n13727, n13728,
         n13729, n13730, n13731, n13732, n13733, n13734, n13735, n13736,
         n13737, n13738, n13739, n13740, n13741, n13742, n13743, n13744,
         n13745, n13746, n13747, n13748, n13749, n13750, n13751, n13752,
         n13753, n13754, n13755, n13756, n13757, n13758, n13759, n13760,
         n13761, n13762, n13763, n13764, n13765, n13766, n13767, n13768,
         n13769, n13770, n13771, n13772, n13773, n13774, n13775, n13776,
         n13777, n13778, n13779, n13780, n13781, n13782, n13783, n13784,
         n13785, n13786, n13787, n13788, n13789, n13790, n13791, n13792,
         n13793, n13794, n13795, n13796, n13797, n13798, n13799, n13800,
         n13801, n13802, n13803, n13804, n13805, n13806, n13807, n13808,
         n13809, n13810, n13811, n13812, n13813, n13814, n13815, n13816,
         n13817, n13818, n13819, n13820, n13821, n13822, n13823, n13824,
         n13825, n13826, n13827, n13828, n13829, n13830, n13831, n13832,
         n13833, n13834, n13835, n13836, n13837, n13838, n13839, n13840,
         n13841, n13842, n13843, n13844, n13845, n13846, n13847, n13848,
         n13849, n13850, n13851, n13852, n13853, n13854, n13855, n13856,
         n13857, n13858, n13859, n13860, n13861, n13862, n13863, n13864,
         n13865, n13866, n13867, n13868, n13869, n13870, n13871, n13872,
         n13873, n13874, n13875, n13876, n13877, n13878, n13879, n13880,
         n13881, n13882, n13883, n13884, n13885, n13886, n13887, n13888,
         n13889, n13890, n13891, n13892, n13893, n13894, n13895, n13896,
         n13897, n13898, n13899, n13900, n13901, n13902, n13903, n13904,
         n13905, n13906, n13907, n13908, n13909, n13910, n13911, n13912,
         n13913, n13914, n13915, n13916, n13917, n13918, n13919, n13920,
         n13921, n13922, n13923, n13924, n13925, n13926, n13927, n13928,
         n13929, n13930, n13931, n13932, n13933, n13934, n13935, n13936,
         n13937, n13938, n13939, n13940, n13941, n13942, n13943, n13944,
         n13945, n13946, n13947, n13948, n13949, n13950, n13951, n13952,
         n13953, n13954, n13955, n13956, n13957, n13958, n13959, n13960,
         n13961, n13962, n13963, n13964, n13965, n13966, n13967, n13968,
         n13969, n13970, n13971, n13972, n13973, n13974, n13975, n13976,
         n13977, n13978, n13979, n13980, n13981, n13982, n13983, n13984,
         n13985, n13986, n13987, n13988, n13989, n13990, n13991, n13992,
         n13993, n13994, n13995, n13996, n13997, n13998, n13999, n14000,
         n14001, n14002, n14003, n14004, n14005, n14006, n14007, n14008,
         n14009, n14010, n14011, n14012, n14013, n14014, n14015, n14016,
         n14017, n14018, n14019, n14020, n14021, n14022, n14023, n14024,
         n14025, n14026, n14027, n14028, n14029, n14030, n14031, n14032,
         n14033, n14034, n14035, n14036, n14037, n14038, n14039, n14040,
         n14041, n14042, n14043, n14044, n14045, n14046, n14047, n14048,
         n14049, n14050, n14051, n14052, n14053, n14054, n14055, n14056,
         n14057, n14058, n14059, n14060, n14061, n14062, n14063, n14064,
         n14065, n14066, n14067, n14068, n14069, n14070, n14071, n14072,
         n14073, n14074, n14075, n14076, n14077, n14078, n14079, n14080,
         n14081, n14082, n14083, n14084, n14085, n14086, n14087, n14088,
         n14089, n14090, n14091, n14092, n14093, n14094, n14095, n14096,
         n14097, n14098, n14099, n14100, n14101, n14102, n14103, n14104,
         n14105, n14106, n14107, n14108, n14109, n14110, n14111, n14112,
         n14113, n14114, n14115, n14116, n14117, n14118, n14119, n14120,
         n14121, n14122, n14123, n14124, n14125, n14126, n14127, n14128,
         n14129, n14130, n14131, n14132, n14133, n14134, n14135, n14136,
         n14137, n14138, n14139, n14140, n14141, n14142, n14143, n14144,
         n14145, n14146, n14147, n14148, n14149, n14150, n14151, n14152,
         n14153, n14154, n14155, n14156, n14157, n14158, n14159, n14160,
         n14161, n14162, n14163, n14164, n14165, n14166, n14167, n14168,
         n14169, n14170, n14171, n14172, n14173, n14174, n14175, n14176,
         n14177, n14178, n14179, n14180, n14181, n14182, n14183, n14184,
         n14185, n14186, n14187, n14188, n14189, n14190, n14191, n14192,
         n14193, n14194, n14195, n14196, n14197, n14198, n14199, n14200,
         n14201, n14202, n14203, n14204, n14205, n14206, n14207, n14208,
         n14209, n14210, n14211, n14212, n14213, n14214, n14215, n14216,
         n14217, n14218, n14219, n14220, n14221, n14222, n14223, n14224,
         n14225, n14226, n14227, n14228, n14229, n14230, n14231, n14232,
         n14233, n14234, n14235, n14236, n14237, n14238, n14239, n14240,
         n14241, n14242, n14243, n14244, n14245, n14246, n14247, n14248,
         n14249, n14250, n14251, n14252, n14253, n14254, n14255, n14256,
         n14257, n14258, n14259, n14260, n14261, n14262, n14263, n14264,
         n14265, n14266, n14267, n14268, n14269, n14270, n14271, n14272,
         n14273, n14274, n14275, n14276, n14277, n14278, n14279, n14280,
         n14281, n14282, n14283, n14284, n14285, n14286, n14287, n14288,
         n14289, n14290, n14291, n14292, n14293, n14294, n14295, n14296,
         n14297, n14298, n14299, n14300, n14301, n14302, n14303, n14304,
         n14305, n14306, n14307, n14308, n14309, n14310, n14311, n14312,
         n14313, n14314, n14315, n14316, n14317, n14318, n14319, n14320,
         n14321, n14322, n14323, n14324, n14325, n14326, n14327, n14328,
         n14329, n14330, n14331, n14332, n14333, n14334, n14335, n14336,
         n14337, n14338, n14339, n14340, n14341, n14342, n14343, n14344,
         n14345, n14346, n14347, n14348, n14349, n14350, n14351, n14352,
         n14353, n14354, n14355, n14356, n14357, n14358, n14359, n14360,
         n14361, n14362, n14363, n14364, n14365, n14366, n14367, n14368,
         n14369, n14370, n14371, n14372, n14373, n14374, n14375, n14376,
         n14377, n14378, n14379, n14380, n14381, n14382, n14383, n14384,
         n14385, n14386, n14387, n14388, n14389, n14390, n14391, n14392,
         n14393, n14394, n14395, n14396, n14397, n14398, n14399, n14400,
         n14401, n14402, n14403, n14404, n14405, n14406, n14407, n14408,
         n14409, n14410, n14411, n14412, n14413, n14414, n14415, n14416,
         n14417, n14418, n14419, n14420, n14421, n14422, n14423, n14424,
         n14425, n14426, n14427, n14428, n14429, n14430, n14431, n14432,
         n14433, n14434, n14435, n14436, n14437, n14438, n14439, n14440,
         n14441, n14442, n14443, n14444, n14445, n14446, n14447, n14448,
         n14449, n14450, n14451, n14452, n14453, n14454, n14455, n14456,
         n14457, n14458, n14459, n14460, n14461, n14462, n14463, n14464,
         n14465, n14466, n14467, n14468, n14469, n14470, n14471, n14472,
         n14473, n14474, n14475, n14476, n14477, n14478, n14479, n14480,
         n14481, n14482, n14483, n14484, n14485, n14486, n14487, n14488,
         n14489, n14490, n14491, n14492, n14493, n14494, n14495, n14496,
         n14497, n14498, n14499, n14500, n14501, n14502, n14503, n14504,
         n14505, n14506, n14507, n14508, n14509, n14510, n14511, n14512,
         n14513, n14514, n14515, n14516, n14517, n14518, n14519, n14520,
         n14521, n14522, n14523, n14524, n14525, n14526, n14527, n14528,
         n14529, n14530, n14531, n14532, n14533, n14534, n14535, n14536,
         n14537, n14538, n14539, n14540, n14541, n14542, n14543, n14544,
         n14545, n14546, n14547, n14548, n14549, n14550, n14551, n14552,
         n14553, n14554, n14555, n14556, n14557, n14558, n14559, n14560,
         n14561, n14562, n14563, n14564, n14565, n14566, n14567, n14568,
         n14569, n14570, n14571, n14572, n14573, n14574, n14575, n14576,
         n14577, n14578, n14579, n14580, n14581, n14582, n14583, n14584,
         n14585, n14586, n14587, n14588, n14589, n14590, n14591, n14592,
         n14593, n14594, n14595, n14596, n14597, n14598, n14599, n14600,
         n14601, n14602, n14603, n14604, n14605, n14606, n14607, n14608,
         n14609, n14610, n14611, n14612, n14613, n14614, n14615, n14616,
         n14617, n14618, n14619, n14620, n14621, n14622, n14623, n14624,
         n14625, n14626, n14627, n14628, n14629, n14630, n14631, n14632,
         n14633, n14634, n14635, n14636, n14637, n14638, n14639, n14640,
         n14641, n14642, n14643, n14644, n14645, n14646, n14647, n14648,
         n14649, n14650, n14651, n14652, n14653, n14654, n14655, n14656,
         n14657, n14658, n14659, n14660, n14661, n14662, n14663, n14664,
         n14665, n14666, n14667, n14668, n14669, n14670, n14671, n14672,
         n14673, n14674, n14675, n14676, n14677, n14678, n14679, n14680,
         n14681, n14682, n14683, n14684, n14685, n14686, n14687, n14688,
         n14689, n14690, n14691, n14692, n14693, n14694, n14695, n14696,
         n14697, n14698, n14699, n14700, n14701, n14702, n14703, n14704,
         n14705, n14706, n14707, n14708, n14709, n14710, n14711, n14712,
         n14713, n14714, n14715, n14716, n14717, n14718, n14719, n14720,
         n14721, n14722, n14723, n14724, n14725, n14726, n14727, n14728,
         n14729, n14730, n14731, n14732, n14733, n14734, n14735, n14736,
         n14737, n14738, n14739, n14740, n14741, n14742, n14743, n14744,
         n14745, n14746, n14747, n14748, n14749, n14750, n14751, n14752,
         n14753, n14754, n14755, n14756, n14757, n14758, n14759, n14760,
         n14761, n14762, n14763, n14764, n14765, n14766, n14767, n14768,
         n14769, n14770, n14771, n14772, n14773, n14774, n14775, n14776,
         n14777, n14778, n14779, n14780, n14781, n14782, n14783, n14784,
         n14785, n14786, n14787, n14788, n14789, n14790, n14791, n14792,
         n14793, n14794, n14795, n14796, n14797, n14798, n14799, n14800,
         n14801, n14802, n14803, n14804, n14805, n14806, n14807, n14808,
         n14809, n14810, n14811, n14812, n14813, n14814, n14815, n14816,
         n14817, n14818, n14819, n14820, n14821, n14822, n14823, n14824,
         n14825, n14826, n14827, n14828, n14829, n14830, n14831, n14832,
         n14833, n14834, n14835, n14836, n14837, n14838, n14839, n14840,
         n14841, n14842, n14843, n14844, n14845, n14846, n14847, n14848,
         n14849, n14850, n14851, n14852, n14853, n14854, n14855, n14856,
         n14857, n14858, n14859, n14860, n14861, n14862, n14863, n14864,
         n14865, n14866, n14867, n14868, n14869, n14870, n14871, n14872,
         n14873, n14874, n14875, n14876, n14877, n14878, n14879, n14880,
         n14881, n14882, n14883, n14884, n14885, n14886, n14887, n14888,
         n14889, n14890, n14891, n14892, n14893, n14894, n14895, n14896,
         n14897, n14898, n14899, n14900, n14901, n14902, n14903, n14904,
         n14905, n14906, n14907, n14908, n14909, n14910, n14911, n14912,
         n14913, n14914, n14915, n14916, n14917, n14918, n14919, n14920,
         n14921, n14922, n14923, n14924, n14925, n14926, n14927, n14928,
         n14929, n14930, n14931, n14932, n14933, n14934, n14935, n14936,
         n14937, n14938, n14939, n14940, n14941, n14942, n14943, n14944,
         n14945, n14946, n14947, n14948, n14949, n14950, n14951, n14952,
         n14953, n14954, n14955, n14956, n14957, n14958, n14959, n14960,
         n14961, n14962, n14963, n14964, n14965, n14966, n14967, n14968,
         n14969, n14970, n14971, n14972, n14973, n14974, n14975, n14976,
         n14977, n14978, n14979, n14980, n14981, n14982, n14983, n14984,
         n14985, n14986, n14987, n14988, n14989, n14990, n14991, n14992,
         n14993, n14994, n14995, n14996, n14997, n14998, n14999, n15000,
         n15001, n15002, n15003, n15004, n15005, n15006, n15007, n15008,
         n15009, n15010, n15011, n15012, n15013, n15014, n15015, n15016,
         n15017, n15018, n15019, n15020, n15021, n15022, n15023, n15024,
         n15025, n15026, n15027, n15028, n15029, n15030, n15031, n15032,
         n15033, n15034, n15035, n15036, n15037, n15038, n15039, n15040,
         n15041, n15042, n15043, n15044, n15045, n15046, n15047, n15048,
         n15049, n15050, n15051, n15052, n15053, n15054, n15055, n15056,
         n15057, n15058, n15059, n15060, n15061, n15062, n15063, n15064,
         n15065, n15066, n15067, n15068, n15069, n15070, n15071, n15072,
         n15073, n15074, n15075, n15076, n15077, n15078, n15079, n15080,
         n15081, n15082, n15083, n15084, n15085, n15086, n15087, n15088,
         n15089, n15090, n15091, n15092, n15093, n15094, n15095, n15096,
         n15097, n15098, n15099, n15100, n15101, n15102, n15103, n15104,
         n15105, n15106, n15107, n15108, n15109, n15110, n15111, n15112,
         n15113, n15114, n15115, n15116, n15117, n15118, n15119, n15120,
         n15121, n15122, n15123, n15124, n15125, n15126, n15127, n15128,
         n15129, n15130, n15131, n15132, n15133, n15134, n15135, n15136,
         n15137, n15138, n15139, n15140, n15141, n15142, n15143, n15144,
         n15145, n15146, n15147, n15148, n15149, n15150, n15151, n15152,
         n15153, n15154, n15155, n15156, n15157, n15158, n15159, n15160,
         n15161, n15162, n15163, n15164, n15165, n15166, n15167, n15168,
         n15169, n15170, n15171, n15172, n15173, n15174, n15175, n15176,
         n15177, n15178, n15179, n15180, n15181, n15182, n15183, n15184,
         n15185, n15186, n15187, n15188, n15189, n15190, n15191, n15192,
         n15193, n15194, n15195, n15196, n15197, n15198, n15199, n15200,
         n15201, n15202, n15203, n15204, n15205, n15206, n15207, n15208,
         n15209, n15210, n15211, n15212, n15213, n15214, n15215, n15216,
         n15217, n15218, n15219, n15220, n15221, n15222, n15223, n15224,
         n15225, n15226, n15227, n15228, n15229, n15230, n15231, n15232,
         n15233, n15234, n15235, n15236, n15237, n15238, n15239, n15240,
         n15241, n15242, n15243, n15244, n15245, n15246, n15247, n15248,
         n15249, n15250, n15251, n15252, n15253, n15254, n15255, n15256,
         n15257, n15258, n15259, n15260, n15261, n15262, n15263, n15264,
         n15265, n15266, n15267, n15268, n15269, n15270, n15271, n15272,
         n15273, n15274, n15275, n15276, n15277, n15278, n15279, n15280,
         n15281, n15282, n15283, n15284, n15285, n15286, n15287, n15288,
         n15289, n15290, n15291, n15292, n15293, n15294, n15295, n15296,
         n15297, n15298, n15299, n15300, n15301, n15302, n15303, n15304,
         n15305, n15306, n15307, n15308, n15309, n15310, n15311, n15312,
         n15313, n15314, n15315, n15316, n15317, n15318, n15319, n15320,
         n15321, n15322, n15323, n15324, n15325, n15326, n15327, n15328,
         n15329, n15330, n15331, n15332, n15333, n15334, n15335, n15336,
         n15337, n15338, n15339, n15340, n15341, n15342, n15343, n15344,
         n15345, n15346, n15347, n15348, n15349, n15350, n15351, n15352,
         n15353, n15354, n15355, n15356, n15357, n15358, n15359, n15360,
         n15361, n15362, n15363, n15364, n15365, n15366, n15367, n15368,
         n15369, n15370, n15371, n15372, n15373, n15374, n15375, n15376,
         n15377, n15378, n15379, n15380, n15381, n15382, n15383, n15384,
         n15385, n15386, n15387, n15388, n15389, n15390, n15391, n15392,
         n15393, n15394, n15395, n15396, n15397, n15398, n15399, n15400,
         n15401, n15402, n15403, n15404, n15405, n15406, n15407, n15408,
         n15409, n15410, n15411, n15412, n15413, n15414, n15415, n15416,
         n15417, n15418, n15419, n15420, n15421, n15422, n15423, n15424,
         n15425, n15426, n15427, n15428, n15429, n15430, n15431, n15432,
         n15433, n15434, n15435, n15436, n15437, n15438, n15439, n15440,
         n15441, n15442, n15443, n15444, n15445, n15446, n15447, n15448,
         n15449, n15450, n15451, n15452, n15453, n15454, n15455, n15456,
         n15457, n15458, n15459, n15460, n15461, n15462, n15463, n15464,
         n15465, n15466, n15467, n15468, n15469, n15470, n15471, n15472,
         n15473, n15474, n15475, n15476, n15477, n15478, n15479, n15480,
         n15481, n15482, n15483, n15484, n15485, n15486, n15487, n15488,
         n15489, n15490, n15491, n15492, n15493, n15494, n15495, n15496,
         n15497, n15498, n15499, n15500, n15501, n15502, n15503, n15504,
         n15505, n15506, n15507, n15508, n15509, n15510, n15511, n15512,
         n15513, n15514, n15515, n15516, n15517, n15518, n15519, n15520,
         n15521, n15522, n15523, n15524, n15525, n15526, n15527, n15528,
         n15529, n15530, n15531, n15532, n15533, n15534, n15535, n15536,
         n15537, n15538, n15539, n15540, n15541, n15542, n15543, n15544,
         n15545, n15546, n15547, n15548, n15549, n15550, n15551, n15552,
         n15553, n15554, n15555, n15556, n15557, n15558, n15559, n15560,
         n15561, n15562, n15563, n15564, n15565, n15566, n15567, n15568,
         n15569, n15570, n15571, n15572, n15573, n15574, n15575, n15576,
         n15577, n15578, n15579, n15580, n15581, n15582, n15583, n15584,
         n15585, n15586, n15587, n15588, n15589, n15590, n15591, n15592,
         n15593, n15594, n15595, n15596, n15597, n15598, n15599, n15600,
         n15601, n15602, n15603, n15604, n15605, n15606, n15607, n15608,
         n15609, n15610, n15611, n15612, n15613, n15614, n15615, n15616,
         n15617, n15618, n15619, n15620, n15621, n15622, n15623, n15624,
         n15625, n15626, n15627, n15628, n15629, n15630, n15631, n15632,
         n15633, n15634, n15635, n15636, n15637, n15638, n15639, n15640,
         n15641, n15642, n15643, n15644, n15645, n15646, n15647, n15648,
         n15649, n15650, n15651, n15652, n15653, n15654, n15655, n15656,
         n15657, n15658, n15659, n15660, n15661, n15662, n15663, n15664,
         n15665, n15666, n15667, n15668, n15669, n15670, n15671, n15672,
         n15673, n15674, n15675, n15676, n15677, n15678, n15679, n15680,
         n15681, n15682, n15683, n15684, n15685, n15686, n15687, n15688,
         n15689, n15690, n15691, n15692, n15693, n15694, n15695, n15696,
         n15697, n15698, n15699, n15700, n15701, n15702, n15703, n15704,
         n15705, n15706, n15707, n15708, n15709, n15710, n15711, n15712,
         n15713, n15714, n15715, n15716, n15717, n15718, n15719, n15720,
         n15721, n15722, n15723, n15724, n15725, n15726, n15727, n15728,
         n15729, n15730, n15731, n15732, n15733, n15734, n15735, n15736,
         n15737, n15738, n15739, n15740, n15741, n15742, n15743, n15744,
         n15745, n15746, n15747, n15748, n15749, n15750, n15751, n15752,
         n15753, n15754, n15755, n15756, n15757, n15758, n15759, n15760,
         n15761, n15762, n15763, n15764, n15765, n15766, n15767, n15768,
         n15769, n15770, n15771, n15772, n15773, n15774, n15775, n15776,
         n15777, n15778, n15779, n15780, n15781, n15782, n15783, n15784,
         n15785, n15786, n15787, n15788, n15789, n15790, n15791, n15792,
         n15793, n15794, n15795, n15796, n15797, n15798, n15799, n15800,
         n15801, n15802, n15803, n15804, n15805, n15806, n15807, n15808,
         n15809, n15810, n15811, n15812, n15813, n15814, n15815, n15816,
         n15817, n15818, n15819, n15820, n15821, n15822, n15823, n15824,
         n15825, n15826, n15827, n15828, n15829, n15830, n15831, n15832,
         n15833, n15834, n15835, n15836, n15837, n15838, n15839, n15840,
         n15841, n15842, n15843, n15844, n15845, n15846, n15847, n15848,
         n15849, n15850, n15851, n15852, n15853, n15854, n15855, n15856,
         n15857, n15858, n15859, n15860, n15861, n15862, n15863, n15864,
         n15865, n15866, n15867, n15868, n15869, n15870, n15871, n15872,
         n15873, n15874, n15875, n15876, n15877, n15878, n15879, n15880,
         n15881, n15882, n15883, n15884, n15885, n15886, n15887, n15888,
         n15889, n15890, n15891, n15892, n15893, n15894, n15895, n15896,
         n15897, n15898, n15899, n15900, n15901, n15902, n15903, n15904,
         n15905, n15906, n15907, n15908, n15909, n15910, n15911, n15912,
         n15913, n15914, n15915, n15916, n15917, n15918, n15919, n15920,
         n15921, n15922, n15923, n15924, n15925, n15926, n15927, n15928,
         n15929, n15930, n15931, n15932, n15933, n15934, n15935, n15936,
         n15937, n15938, n15939, n15940, n15941, n15942, n15943, n15944,
         n15945, n15946, n15947, n15948, n15949, n15950, n15951, n15952,
         n15953, n15954, n15955, n15956, n15957, n15958, n15959, n15960,
         n15961, n15962, n15963, n15964, n15965, n15966, n15967, n15968,
         n15969, n15970, n15971, n15972, n15973, n15974, n15975, n15976,
         n15977, n15978, n15979, n15980, n15981, n15982, n15983, n15984,
         n15985, n15986, n15987, n15988, n15989, n15990, n15991, n15992,
         n15993, n15994, n15995, n15996, n15997, n15998, n15999, n16000,
         n16001, n16002, n16003, n16004, n16005, n16006, n16007, n16008,
         n16009, n16010, n16011, n16012, n16013, n16014, n16015, n16016,
         n16017, n16018, n16019, n16020, n16021, n16022, n16023, n16024,
         n16025, n16026, n16027, n16028, n16029, n16030, n16031, n16032,
         n16033, n16034, n16035, n16036, n16037, n16038, n16039, n16040,
         n16041, n16042, n16043, n16044, n16045, n16046, n16047, n16048,
         n16049, n16050, n16051, n16052, n16053, n16054, n16055, n16056,
         n16057, n16058, n16059, n16060, n16061, n16062, n16063, n16064,
         n16065, n16066, n16067, n16068, n16069, n16070, n16071, n16072,
         n16073, n16074, n16075, n16076, n16077, n16078, n16079, n16080,
         n16081, n16082, n16083, n16084, n16085, n16086, n16087, n16088,
         n16089, n16090, n16091, n16092, n16093, n16094, n16095, n16096,
         n16097, n16098, n16099, n16100, n16101, n16102, n16103, n16104,
         n16105, n16106, n16107, n16108, n16109, n16110, n16111, n16112,
         n16113, n16114, n16115, n16116, n16117, n16118, n16119, n16120,
         n16121, n16122, n16123, n16124, n16125, n16126, n16127, n16128,
         n16129, n16130, n16131, n16132, n16133, n16134, n16135, n16136,
         n16137, n16138, n16139, n16140, n16141, n16142, n16143, n16144,
         n16145, n16146, n16147, n16148, n16149, n16150, n16151, n16152,
         n16153, n16154, n16155, n16156, n16157, n16158, n16159, n16160,
         n16161, n16162, n16163, n16164, n16165, n16166, n16167, n16168,
         n16169, n16170, n16171, n16172, n16173, n16174, n16175, n16176,
         n16177, n16178, n16179, n16180, n16181, n16182, n16183, n16184,
         n16185, n16186, n16187, n16188, n16189, n16190, n16191, n16192,
         n16193, n16194, n16195, n16196, n16197, n16198, n16199, n16200,
         n16201, n16202, n16203, n16204, n16205, n16206, n16207, n16208,
         n16209, n16210, n16211, n16212, n16213, n16214, n16215, n16216,
         n16217, n16218, n16219, n16220, n16221, n16222, n16223, n16224,
         n16225, n16226, n16227, n16228, n16229, n16230, n16231, n16232,
         n16233, n16234, n16235, n16236, n16237, n16238, n16239, n16240,
         n16241, n16242, n16243, n16244, n16245, n16246, n16247, n16248,
         n16249, n16250, n16251, n16252, n16253, n16254, n16255, n16256,
         n16257, n16258, n16259, n16260, n16261, n16262, n16263, n16264,
         n16265, n16266, n16267, n16268, n16269, n16270, n16271, n16272,
         n16273, n16274, n16275, n16276, n16277, n16278, n16279, n16280,
         n16281, n16282, n16283, n16284, n16285, n16286, n16287, n16288,
         n16289, n16290, n16291, n16292, n16293, n16294, n16295, n16296,
         n16297, n16298, n16299, n16300, n16301, n16302, n16303, n16304,
         n16305, n16306, n16307, n16308, n16309, n16310, n16311, n16312,
         n16313, n16314, n16315, n16316, n16317, n16318, n16319, n16320,
         n16321, n16322, n16323, n16324, n16325, n16326, n16327, n16328,
         n16329, n16330, n16331, n16332, n16333, n16334, n16335, n16336,
         n16337, n16338, n16339, n16340, n16341, n16342, n16343, n16344,
         n16345, n16346, n16347, n16348, n16349, n16350, n16351, n16352,
         n16353, n16354, n16355, n16356, n16357, n16358, n16359, n16360,
         n16361, n16362, n16363, n16364, n16365, n16366, n16367, n16368,
         n16369, n16370, n16371, n16372, n16373, n16374, n16375, n16376,
         n16377, n16378, n16379, n16380, n16381, n16382, n16383, n16384,
         n16385, n16386, n16387, n16388, n16389, n16390, n16391, n16392,
         n16393, n16394, n16395, n16396, n16397, n16398, n16399, n16400,
         n16401, n16402, n16403, n16404, n16405, n16406, n16407, n16408,
         n16409, n16410, n16411, n16412, n16413, n16414, n16415, n16416,
         n16417, n16418, n16419, n16420, n16421, n16422, n16423, n16424,
         n16425, n16426, n16427, n16428, n16429, n16430, n16431, n16432,
         n16433, n16434, n16435, n16436, n16437, n16438, n16439, n16440,
         n16441, n16442, n16443, n16444, n16445, n16446, n16447, n16448,
         n16449, n16450, n16451, n16452, n16453, n16454, n16455, n16456,
         n16457, n16458, n16459, n16460, n16461, n16462, n16463, n16464,
         n16465, n16466, n16467, n16468, n16469, n16470, n16471, n16472,
         n16473, n16474, n16475, n16476, n16477, n16478, n16479, n16480,
         n16481, n16482, n16483, n16484, n16485, n16486, n16487, n16488,
         n16489, n16490, n16491, n16492, n16493, n16494, n16495, n16496,
         n16497, n16498, n16499, n16500, n16501, n16502, n16503, n16504,
         n16505, n16506, n16507, n16508, n16509, n16510, n16511, n16512,
         n16513, n16514, n16515, n16516, n16517, n16518, n16519, n16520,
         n16521, n16522, n16523, n16524, n16525, n16526, n16527, n16528,
         n16529, n16530, n16531, n16532, n16533, n16534, n16535, n16536,
         n16537, n16538, n16539, n16540, n16541, n16542, n16543, n16544,
         n16545, n16546, n16547, n16548, n16549, n16550, n16551, n16552,
         n16553, n16554, n16555, n16556, n16557, n16558, n16559, n16560,
         n16561, n16562, n16563, n16564, n16565, n16566, n16567, n16568,
         n16569, n16570, n16571, n16572, n16573, n16574, n16575, n16576,
         n16577, n16578, n16579, n16580, n16581, n16582, n16583, n16584,
         n16585, n16586, n16587, n16588, n16589, n16590, n16591, n16592,
         n16593, n16594, n16595, n16596, n16597, n16598, n16599, n16600,
         n16601, n16602, n16603, n16604, n16605, n16606, n16607, n16608,
         n16609, n16610, n16611, n16612, n16613, n16614, n16615, n16616,
         n16617, n16618, n16619, n16620, n16621, n16622, n16623, n16624,
         n16625, n16626, n16627, n16628, n16629, n16630, n16631, n16632,
         n16633, n16634, n16635, n16636, n16637, n16638, n16639, n16640,
         n16641, n16642, n16643, n16644, n16645, n16646, n16647, n16648,
         n16649, n16650, n16651, n16652, n16653, n16654, n16655, n16656,
         n16657, n16658, n16659, n16660, n16661, n16662, n16663, n16664,
         n16665, n16666, n16667, n16668, n16669, n16670, n16671, n16672,
         n16673, n16674, n16675, n16676, n16677, n16678, n16679, n16680,
         n16681, n16682, n16683, n16684, n16685, n16686, n16687, n16688,
         n16689, n16690, n16691, n16692, n16693, n16694, n16695, n16696,
         n16697, n16698, n16699, n16700, n16701, n16702, n16703, n16704,
         n16705, n16706, n16707, n16708, n16709, n16710, n16711, n16712,
         n16713, n16714, n16715, n16716, n16717, n16718, n16719, n16720,
         n16721, n16722, n16723, n16724, n16725, n16726, n16727, n16728,
         n16729, n16730, n16731, n16732, n16733, n16734, n16735, n16736,
         n16737, n16738, n16739, n16740, n16741, n16742, n16743, n16744,
         n16745, n16746, n16747, n16748, n16749, n16750, n16751, n16752,
         n16753, n16754, n16755, n16756, n16757, n16758, n16759, n16760,
         n16761, n16762, n16763, n16764, n16765, n16766, n16767, n16768,
         n16769, n16770, n16771, n16772, n16773, n16774, n16775, n16776,
         n16777, n16778, n16779, n16780, n16781, n16782, n16783, n16784,
         n16785, n16786, n16787, n16788, n16789, n16790, n16791, n16792,
         n16793, n16794, n16795, n16796, n16797, n16798, n16799, n16800,
         n16801, n16802, n16803, n16804, n16805, n16806, n16807, n16808,
         n16809, n16810, n16811, n16812, n16813, n16814, n16815, n16816,
         n16817, n16818, n16819, n16820, n16821, n16822, n16823, n16824,
         n16825, n16826, n16827, n16828, n16829, n16830, n16831, n16832,
         n16833, n16834, n16835, n16836, n16837, n16838, n16839, n16840,
         n16841, n16842, n16843, n16844, n16845, n16846, n16847, n16848,
         n16849, n16850, n16851, n16852, n16853, n16854, n16855, n16856,
         n16857, n16858, n16859, n16860, n16861, n16862, n16863, n16864,
         n16865, n16866, n16867, n16868, n16869, n16870, n16871, n16872,
         n16873, n16874, n16875, n16876, n16877, n16878, n16879, n16880,
         n16881, n16882, n16883, n16884, n16885, n16886, n16887, n16888,
         n16889, n16890, n16891, n16892, n16893, n16894, n16895, n16896,
         n16897, n16898, n16899, n16900, n16901, n16902, n16903, n16904,
         n16905, n16906, n16907, n16908, n16909, n16910, n16911, n16912,
         n16913, n16914, n16915, n16916, n16917, n16918, n16919, n16920,
         n16921, n16922, n16923, n16924, n16925, n16926, n16927, n16928,
         n16929, n16930, n16931, n16932, n16933, n16934, n16935, n16936,
         n16937, n16938, n16939, n16940, n16941, n16942, n16943, n16944,
         n16945, n16946, n16947, n16948, n16949, n16950, n16951, n16952,
         n16953, n16954, n16955, n16956, n16957, n16958, n16959, n16960,
         n16961, n16962, n16963, n16964, n16965, n16966, n16967, n16968,
         n16969, n16970, n16971, n16972, n16973, n16974, n16975, n16976,
         n16977, n16978, n16979, n16980, n16981, n16982, n16983, n16984,
         n16985, n16986, n16987, n16988, n16989, n16990, n16991, n16992,
         n16993, n16994, n16995, n16996, n16997, n16998, n16999, n17000,
         n17001, n17002, n17003, n17004, n17005, n17006, n17007, n17008,
         n17009, n17010, n17011, n17012, n17013, n17014, n17015, n17016,
         n17017, n17018, n17019, n17020, n17021, n17022, n17023, n17024,
         n17025, n17026, n17027, n17028, n17029, n17030, n17031, n17032,
         n17033, n17034, n17035, n17036, n17037, n17038, n17039, n17040,
         n17041, n17042, n17043, n17044, n17045, n17046, n17047, n17048,
         n17049, n17050, n17051, n17052, n17053, n17054, n17055, n17056,
         n17057, n17058, n17059, n17060, n17061, n17062, n17063, n17064,
         n17065, n17066, n17067, n17068, n17069, n17070, n17071, n17072,
         n17073, n17074, n17075, n17076, n17077, n17078, n17079, n17080,
         n17081, n17082, n17083, n17084, n17085, n17086, n17087, n17088,
         n17089, n17090, n17091, n17092, n17093, n17094, n17095, n17096,
         n17097, n17098, n17099, n17100, n17101, n17102, n17103, n17104,
         n17105, n17106, n17107, n17108, n17109, n17110, n17111, n17112,
         n17113, n17114, n17115, n17116, n17117, n17118, n17119, n17120,
         n17121, n17122, n17123, n17124, n17125, n17126, n17127, n17128,
         n17129, n17130, n17131, n17132, n17133, n17134, n17135, n17136,
         n17137, n17138, n17139, n17140, n17141, n17142, n17143, n17144,
         n17145, n17146, n17147, n17148, n17149, n17150, n17151, n17152,
         n17153, n17154, n17155, n17156, n17157, n17158, n17159, n17160,
         n17161, n17162, n17163, n17164, n17165, n17166, n17167, n17168,
         n17169, n17170, n17171, n17172, n17173, n17174, n17175, n17176,
         n17177, n17178, n17179, n17180, n17181, n17182, n17183, n17184,
         n17185, n17186, n17187, n17188, n17189, n17190, n17191, n17192,
         n17193, n17194, n17195, n17196, n17197, n17198, n17199, n17200,
         n17201, n17202, n17203, n17204, n17205, n17206, n17207, n17208,
         n17209, n17210, n17211, n17212, n17213, n17214, n17215, n17216,
         n17217, n17218, n17219, n17220, n17221, n17222, n17223, n17224,
         n17225, n17226, n17227, n17228, n17229, n17230, n17231, n17232,
         n17233, n17234, n17235, n17236, n17237, n17238, n17239, n17240,
         n17241, n17242, n17243, n17244, n17245, n17246, n17247, n17248,
         n17249, n17250, n17251, n17252, n17253, n17254, n17255, n17256,
         n17257, n17258, n17259, n17260, n17261, n17262, n17263, n17264,
         n17265, n17266, n17267, n17268, n17269, n17270, n17271, n17272,
         n17273, n17274, n17275, n17276, n17277, n17278, n17279, n17280,
         n17281, n17282, n17283, n17284, n17285, n17286, n17287, n17288,
         n17289, n17290, n17291, n17292, n17293, n17294, n17295, n17296,
         n17297, n17298, n17299, n17300, n17301, n17302, n17303, n17304,
         n17305, n17306, n17307, n17308, n17309, n17310, n17311, n17312,
         n17313, n17314, n17315, n17316, n17317, n17318, n17319, n17320,
         n17321, n17322, n17323, n17324, n17325, n17326, n17327, n17328,
         n17329, n17330, n17331, n17332, n17333, n17334, n17335, n17336,
         n17337, n17338, n17339, n17340, n17341, n17342, n17343, n17344,
         n17345, n17346, n17347, n17348, n17349, n17350, n17351, n17352,
         n17353, n17354, n17355, n17356, n17357, n17358, n17359, n17360,
         n17361, n17362, n17363, n17364, n17365, n17366, n17367, n17368,
         n17369, n17370, n17371, n17372, n17373, n17374, n17375, n17376,
         n17377, n17378, n17379, n17380, n17381, n17382, n17383, n17384,
         n17385, n17386, n17387, n17388, n17389, n17390, n17391, n17392,
         n17393, n17394, n17395, n17396, n17397, n17398, n17399, n17400,
         n17401, n17402, n17403, n17404, n17405, n17406, n17407, n17408,
         n17409, n17410, n17411, n17412, n17413, n17414, n17415, n17416,
         n17417, n17418, n17419, n17420, n17421, n17422, n17423, n17424,
         n17425, n17426, n17427, n17428, n17429, n17430, n17431, n17432,
         n17433, n17434, n17435, n17436, n17437, n17438, n17439, n17440,
         n17441, n17442, n17443, n17444, n17445, n17446, n17447, n17448,
         n17449, n17450, n17451, n17452, n17453, n17454, n17455, n17456,
         n17457, n17458, n17459, n17460, n17461, n17462, n17463, n17464,
         n17465, n17466, n17467, n17468, n17469, n17470, n17471, n17472,
         n17473, n17474, n17475, n17476, n17477, n17478, n17479, n17480,
         n17481, n17482, n17483, n17484, n17485, n17486, n17487, n17488,
         n17489, n17490, n17491, n17492, n17493, n17494, n17495, n17496,
         n17497, n17498, n17499, n17500, n17501, n17502, n17503, n17504,
         n17505, n17506, n17507, n17508, n17509, n17510, n17511, n17512,
         n17513, n17514, n17515, n17516, n17517, n17518, n17519, n17520,
         n17521, n17522, n17523, n17524, n17525, n17526, n17527, n17528,
         n17529, n17530, n17531, n17532, n17533, n17534, n17535, n17536,
         n17537, n17538, n17539, n17540, n17541, n17542, n17543, n17544,
         n17545, n17546, n17547, n17548, n17549, n17550, n17551, n17552,
         n17553, n17554, n17555, n17556, n17557, n17558, n17559, n17560,
         n17561, n17562, n17563, n17564, n17565, n17566, n17567, n17568,
         n17569, n17570, n17571, n17572, n17573, n17574, n17575, n17576,
         n17577, n17578, n17579, n17580, n17581, n17582, n17583, n17584,
         n17585, n17586, n17587, n17588, n17589, n17590, n17591, n17592,
         n17593, n17594, n17595, n17596, n17597, n17598, n17599, n17600,
         n17601, n17602, n17603, n17604, n17605, n17606, n17607, n17608,
         n17609, n17610, n17611, n17612, n17613, n17614, n17615, n17616,
         n17617, n17618, n17619, n17620, n17621, n17622, n17623, n17624,
         n17625, n17626, n17627, n17628, n17629, n17630, n17631, n17632,
         n17633, n17634, n17635, n17636, n17637, n17638, n17639, n17640,
         n17641, n17642, n17643, n17644, n17645, n17646, n17647, n17648,
         n17649, n17650, n17651, n17652, n17653, n17654, n17655, n17656,
         n17657, n17658, n17659, n17660, n17661, n17662, n17663, n17664,
         n17665, n17666, n17667, n17668, n17669, n17670, n17671, n17672,
         n17673, n17674, n17675, n17676, n17677, n17678, n17679, n17680,
         n17681, n17682, n17683, n17684, n17685, n17686, n17687, n17688,
         n17689, n17690, n17691, n17692, n17693, n17694, n17695, n17696,
         n17697, n17698, n17699, n17700, n17701, n17702, n17703, n17704,
         n17705, n17706, n17707, n17708, n17709, n17710, n17711, n17712,
         n17713, n17714, n17715, n17716, n17717, n17718, n17719, n17720,
         n17721, n17722, n17723, n17724, n17725, n17726, n17727, n17728,
         n17729, n17730, n17731, n17732, n17733, n17734, n17735, n17736,
         n17737, n17738, n17739, n17740, n17741, n17742, n17743, n17744,
         n17745, n17746, n17747, n17748, n17749, n17750, n17751, n17752,
         n17753, n17754, n17755, n17756, n17757, n17758, n17759, n17760,
         n17761, n17762, n17763, n17764, n17765, n17766, n17767, n17768,
         n17769, n17770, n17771, n17772, n17773, n17774, n17775, n17776,
         n17777, n17778, n17779, n17780, n17781, n17782, n17783, n17784,
         n17785, n17786, n17787, n17788, n17789, n17790, n17791, n17792,
         n17793, n17794, n17795, n17796, n17797, n17798, n17799, n17800,
         n17801, n17802, n17803, n17804, n17805, n17806, n17807, n17808,
         n17809, n17810, n17811, n17812, n17813, n17814, n17815, n17816,
         n17817, n17818, n17819, n17820, n17821, n17822, n17823, n17824,
         n17825, n17826, n17827, n17828, n17829, n17830, n17831, n17832,
         n17833, n17834, n17835, n17836, n17837, n17838, n17839, n17840,
         n17841, n17842, n17843, n17844, n17845, n17846, n17847, n17848,
         n17849, n17850, n17851, n17852, n17853, n17854, n17855, n17856,
         n17857, n17858, n17859, n17860, n17861, n17862, n17863, n17864,
         n17865, n17866, n17867, n17868, n17869, n17870, n17871, n17872,
         n17873, n17874, n17875, n17876, n17877, n17878, n17879, n17880,
         n17881, n17882, n17883, n17884, n17885, n17886, n17887, n17888,
         n17889, n17890, n17891, n17892, n17893, n17894, n17895, n17896,
         n17897, n17898, n17899, n17900, n17901, n17902, n17903, n17904,
         n17905, n17906, n17907, n17908, n17909, n17910, n17911, n17912,
         n17913, n17914, n17915, n17916, n17917, n17918, n17919, n17920,
         n17921, n17922, n17923, n17924, n17925, n17926, n17927, n17928,
         n17929, n17930, n17931, n17932, n17933, n17934, n17935, n17936,
         n17937, n17938, n17939, n17940, n17941, n17942, n17943, n17944,
         n17945, n17946, n17947, n17948, n17949, n17950, n17951, n17952,
         n17953, n17954, n17955, n17956, n17957, n17958, n17959, n17960,
         n17961, n17962, n17963, n17964, n17965, n17966, n17967, n17968,
         n17969, n17970, n17971, n17972, n17973, n17974, n17975, n17976,
         n17977, n17978, n17979, n17980, n17981, n17982, n17983, n17984,
         n17985, n17986, n17987, n17988, n17989, n17990, n17991, n17992,
         n17993, n17994, n17995, n17996, n17997, n17998, n17999, n18000,
         n18001, n18002, n18003, n18004, n18005, n18006, n18007, n18008,
         n18009, n18010, n18011, n18012, n18013, n18014, n18015, n18016,
         n18017, n18018, n18019, n18020, n18021, n18022, n18023, n18024,
         n18025, n18026, n18027, n18028, n18029, n18030, n18031, n18032,
         n18033, n18034, n18035, n18036, n18037, n18038, n18039, n18040,
         n18041, n18042, n18043, n18044, n18045, n18046, n18047, n18048,
         n18049, n18050, n18051, n18052, n18053, n18054, n18055, n18056,
         n18057, n18058, n18059, n18060, n18061, n18062, n18063, n18064,
         n18065, n18066, n18067, n18068, n18069, n18070, n18071, n18072,
         n18073, n18074, n18075, n18076, n18077, n18078, n18079, n18080,
         n18081, n18082, n18083, n18084, n18085, n18086, n18087, n18088,
         n18089, n18090, n18091, n18092, n18093, n18094, n18095, n18096,
         n18097, n18098, n18099, n18100, n18101, n18102, n18103, n18104,
         n18105, n18106, n18107, n18108, n18109, n18110, n18111, n18112,
         n18113, n18114, n18115, n18116, n18117, n18118, n18119, n18120,
         n18121, n18122, n18123, n18124, n18125, n18126, n18127, n18128,
         n18129, n18130, n18131, n18132, n18133, n18134, n18135, n18136,
         n18137, n18138, n18139, n18140, n18141, n18142, n18143, n18144,
         n18145, n18146, n18147, n18148, n18149, n18150, n18151, n18152,
         n18153, n18154, n18155, n18156, n18157, n18158, n18159, n18160,
         n18161, n18162, n18163, n18164, n18165, n18166, n18167, n18168,
         n18169, n18170, n18171, n18172, n18173, n18174, n18175, n18176,
         n18177, n18178, n18179, n18180, n18181, n18182, n18183, n18184,
         n18185, n18186, n18187, n18188, n18189, n18190, n18191, n18192,
         n18193, n18194, n18195, n18196, n18197, n18198, n18199, n18200,
         n18201, n18202, n18203, n18204, n18205, n18206, n18207, n18208,
         n18209, n18210, n18211, n18212, n18213, n18214, n18215, n18216,
         n18217, n18218, n18219, n18220, n18221, n18222, n18223, n18224,
         n18225, n18226, n18227, n18228, n18229, n18230, n18231, n18232,
         n18233, n18234, n18235, n18236, n18237, n18238, n18239, n18240,
         n18241, n18242, n18243, n18244, n18245, n18246, n18247, n18248,
         n18249, n18250, n18251, n18252, n18253, n18254, n18255, n18256,
         n18257, n18258, n18259, n18260, n18261, n18262, n18263, n18264,
         n18265, n18266, n18267, n18268, n18269, n18270, n18271, n18272,
         n18273, n18274, n18275, n18276, n18277, n18278, n18279, n18280,
         n18281, n18282, n18283, n18284, n18285, n18286, n18287, n18288,
         n18289, n18290, n18291, n18292, n18293, n18294, n18295, n18296,
         n18297, n18298, n18299, n18300, n18301, n18302, n18303, n18304,
         n18305, n18306, n18307, n18308, n18309, n18310, n18311, n18312,
         n18313, n18314, n18315, n18316, n18317, n18318, n18319, n18320,
         n18321, n18322, n18323, n18324, n18325, n18326, n18327, n18328,
         n18329, n18330, n18331, n18332, n18333, n18334, n18335, n18336,
         n18337, n18338, n18339, n18340, n18341, n18342, n18343, n18344,
         n18345, n18346, n18347, n18348, n18349, n18350, n18351, n18352,
         n18353, n18354, n18355, n18356, n18357, n18358, n18359, n18360,
         n18361, n18362, n18363, n18364, n18365, n18366, n18367, n18368,
         n18369, n18370, n18371, n18372, n18373, n18374, n18375, n18376,
         n18377, n18378, n18379, n18380, n18381, n18382, n18383, n18384,
         n18385, n18386, n18387, n18388, n18389, n18390, n18391, n18392,
         n18393, n18394, n18395, n18396, n18397, n18398, n18399, n18400,
         n18401, n18402, n18403, n18404, n18405, n18406, n18407, n18408,
         n18409, n18410, n18411, n18412, n18413, n18414, n18415, n18416,
         n18417, n18418, n18419, n18420, n18421, n18422, n18423, n18424,
         n18425, n18426, n18427, n18428, n18429, n18430, n18431, n18432,
         n18433, n18434, n18435, n18436, n18437, n18438, n18439, n18440,
         n18441, n18442, n18443, n18444, n18445, n18446, n18447, n18448,
         n18449, n18450, n18451, n18452, n18453, n18454, n18455, n18456,
         n18457, n18458, n18459, n18460, n18461, n18462, n18463, n18464,
         n18465, n18466, n18467, n18468, n18469, n18470, n18471, n18472,
         n18473, n18474, n18475, n18476, n18477, n18478, n18479, n18480,
         n18481, n18482, n18483, n18484, n18485, n18486, n18487, n18488,
         n18489, n18490, n18491, n18492, n18493, n18494, n18495, n18496,
         n18497, n18498, n18499, n18500, n18501, n18502, n18503, n18504,
         n18505, n18506, n18507, n18508, n18509, n18510, n18511, n18512,
         n18513, n18514, n18515, n18516, n18517, n18518, n18519, n18520,
         n18521, n18522, n18523, n18524, n18525, n18526, n18527, n18528,
         n18529, n18530, n18531, n18532, n18533, n18534, n18535, n18536,
         n18537, n18538, n18539, n18540, n18541, n18542, n18543, n18544,
         n18545, n18546, n18547, n18548, n18549, n18550, n18551, n18552,
         n18553, n18554, n18555, n18556, n18557, n18558, n18559, n18560,
         n18561, n18562, n18563, n18564, n18565, n18566, n18567, n18568,
         n18569, n18570, n18571, n18572, n18573, n18574, n18575, n18576,
         n18577, n18578, n18579, n18580, n18581, n18582, n18583, n18584,
         n18585, n18586, n18587, n18588, n18589, n18590, n18591, n18592,
         n18593, n18594, n18595, n18596, n18597, n18598, n18599, n18600,
         n18601, n18602, n18603, n18604, n18605, n18606, n18607, n18608,
         n18609, n18610, n18611, n18612, n18613, n18614, n18615, n18616,
         n18617, n18618, n18619, n18620, n18621, n18622, n18623, n18624,
         n18625, n18626, n18627, n18628, n18629, n18630, n18631, n18632,
         n18633, n18634, n18635, n18636, n18637, n18638, n18639, n18640,
         n18641, n18642, n18643, n18644, n18645, n18646, n18647, n18648,
         n18649, n18650, n18651, n18652, n18653, n18654, n18655, n18656,
         n18657, n18658, n18659, n18660, n18661, n18662, n18663, n18664,
         n18665, n18666, n18667, n18668, n18669, n18670, n18671, n18672,
         n18673, n18674, n18675, n18676, n18677, n18678, n18679, n18680,
         n18681, n18682, n18683, n18684, n18685, n18686, n18687, n18688,
         n18689, n18690, n18691, n18692, n18693, n18694, n18695, n18696,
         n18697, n18698, n18699, n18700, n18701, n18702, n18703, n18704,
         n18705, n18706, n18707, n18708, n18709, n18710, n18711, n18712,
         n18713, n18714, n18715, n18716, n18717, n18718, n18719, n18720,
         n18721, n18722, n18723, n18724, n18725, n18726, n18727, n18728,
         n18729, n18730, n18731, n18732, n18733, n18734, n18735, n18736,
         n18737, n18738, n18739, n18740, n18741, n18742, n18743, n18744,
         n18745, n18746, n18747, n18748, n18749, n18750, n18751, n18752,
         n18753, n18754, n18755, n18756, n18757, n18758, n18759, n18760,
         n18761, n18762, n18763, n18764, n18765, n18766, n18767, n18768,
         n18769, n18770, n18771, n18772, n18773, n18774, n18775, n18776,
         n18777, n18778, n18779, n18780, n18781, n18782, n18783, n18784,
         n18785, n18786, n18787, n18788, n18789, n18790, n18791, n18792,
         n18793, n18794, n18795, n18796, n18797, n18798, n18799, n18800,
         n18801, n18802, n18803, n18804, n18805, n18806, n18807, n18808,
         n18809, n18810, n18811, n18812, n18813, n18814, n18815, n18816,
         n18817, n18818, n18819, n18820, n18821, n18822, n18823, n18824,
         n18825, n18826, n18827, n18828, n18829, n18830, n18831, n18832,
         n18833, n18834, n18835, n18836, n18837, n18838, n18839, n18840,
         n18841, n18842, n18843, n18844, n18845, n18846, n18847, n18848,
         n18849, n18850, n18851, n18852, n18853, n18854, n18855, n18856,
         n18857, n18858, n18859, n18860, n18861, n18862, n18863, n18864,
         n18865, n18866, n18867, n18868, n18869, n18870, n18871, n18872,
         n18873, n18874, n18875, n18876, n18877, n18878, n18879, n18880,
         n18881, n18882, n18883, n18884, n18885, n18886, n18887, n18888,
         n18889, n18890, n18891, n18892, n18893, n18894, n18895, n18896,
         n18897, n18898, n18899, n18900, n18901, n18902, n18903, n18904,
         n18905, n18906, n18907, n18908, n18909, n18910, n18911, n18912,
         n18913, n18914, n18915, n18916, n18917, n18918, n18919, n18920,
         n18921, n18922, n18923, n18924, n18925, n18926, n18927, n18928,
         n18929, n18930, n18931, n18932, n18933, n18934, n18935, n18936,
         n18937, n18938, n18939, n18940, n18941, n18942, n18943, n18944,
         n18945, n18946, n18947, n18948, n18949, n18950, n18951, n18952,
         n18953, n18954, n18955, n18956, n18957, n18958, n18959, n18960,
         n18961, n18962, n18963, n18964, n18965, n18966, n18967, n18968,
         n18969, n18970, n18971, n18972, n18973, n18974, n18975, n18976,
         n18977, n18978, n18979, n18980, n18981, n18982, n18983, n18984,
         n18985, n18986, n18987, n18988, n18989, n18990, n18991, n18992,
         n18993, n18994, n18995, n18996, n18997, n18998, n18999, n19000,
         n19001, n19002, n19003, n19004, n19005, n19006, n19007, n19008,
         n19009, n19010, n19011, n19012, n19013, n19015, n19016, n19017,
         n19018, n19019, n19020, n19021, n19022, n19023, n19024, n19025,
         n19026, n19027, n19028, n19029, n19030, n19031, n19032, n19033,
         n19034, n19035, n19036, n19037, n19038, n19039, n19040, n19041,
         n19042, n19043, n19044, n19045, n19046, n19047, n19048, n19049,
         n19050, n19051, n19052, n19053, n19054, n19055, n19056, n19057,
         n19058, n19059, n19060, n19061, n19062, n19063, n19064, n19065,
         n19066, n19067, n19068, n19069, n19070, n19071, n19072, n19073,
         n19074, n19075, n19076, n19077, n19078, n19079, n19080, n19081,
         n19082, n19083, n19084, n19085, n19086, n19087, n19088, n19089,
         n19090, n19091, n19092, n19093, n19094, n19095, n19096, n19097,
         n19098, n19099, n19100, n19101, n19102, n19103, n19104, n19105,
         n19106, n19107, n19108, n19109, n19110, n19111, n19112, n19113,
         n19114, n19115, n19116, n19117, n19118, n19119, n19120, n19121,
         n19122, n19123, n19124, n19125, n19126, n19127, n19128, n19129,
         n19130, n19131, n19132, n19133, n19134, n19135, n19136, n19137,
         n19138, n19139, n19140, n19141, n19142, n19143, n19144, n19145,
         n19146, n19147, n19148, n19149, n19150, n19151, n19152, n19153,
         n19154, n19155, n19156, n19157, n19158, n19159, n19160, n19161,
         n19162, n19163, n19164, n19165, n19166, n19167, n19168, n19169,
         n19170, n19171, n19172, n19173, n19174, n19175, n19176, n19177,
         n19178, n19179, n19180, n19181, n19182, n19183, n19184, n19185,
         n19186, n19187, n19188, n19189, n19190, n19191, n19192, n19193,
         n19194, n19195, n19196, n19197, n19198, n19199, n19200, n19201,
         n19202, n19203, n19204, n19205, n19206, n19207, n19208, n19209,
         n19210, n19211, n19212, n19213, n19214, n19215, n19216, n19217,
         n19218, n19219, n19220, n19221, n19222, n19223, n19224, n19225,
         n19226, n19227, n19228, n19229, n19230, n19231, n19232, n19233,
         n19234, n19235, n19236, n19237, n19238, n19239, n19240, n19241,
         n19242, n19243, n19244, n19245, n19246, n19247, n19248, n19249,
         n19250, n19251, n19252, n19253, n19254, n19255, n19256, n19257,
         n19258, n19259, n19260, n19261, n19262, n19263, n19264, n19265,
         n19266, n19267, n19268, n19269, n19270, n19271, n19272, n19273,
         n19274, n19275, n19276, n19277, n19278, n19279, n19280, n19281,
         n19282, n19283, n19284, n19285, n19286, n19287, n19288, n19289,
         n19290, n19291, n19292, n19293, n19294, n19295, n19296, n19297,
         n19298, n19299, n19300, n19301, n19302, n19303, n19304, n19305,
         n19306, n19307, n19308, n19309, n19310, n19311, n19312, n19313,
         n19314, n19315, n19316, n19317, n19318, n19319, n19320, n19321,
         n19322, n19323, n19324, n19325, n19326, n19327, n19328, n19329,
         n19330, n19331, n19332, n19333, n19334, n19335, n19336, n19337,
         n19338, n19339, n19340, n19341, n19342, n19343, n19344, n19345,
         n19346, n19347, n19348, n19349, n19350, n19351, n19352, n19353,
         n19354, n19355, n19356, n19357, n19358, n19359, n19360, n19361,
         n19362, n19363, n19364, n19365, n19366, n19367, n19368, n19369,
         n19370, n19371, n19372, n19373, n19374, n19375, n19376, n19377,
         n19378, n19379, n19380, n19381, n19382, n19383, n19384, n19385,
         n19386, n19387, n19388, n19389, n19390, n19391, n19392, n19393,
         n19394, n19395, n19396, n19397, n19398, n19399, n19400, n19401,
         n19402, n19403, n19404, n19405, n19406, n19407, n19408, n19409,
         n19410, n19411, n19412, n19413, n19414, n19415, n19416, n19417,
         n19418, n19419, n19420, n19421, n19422, n19423, n19424, n19425,
         n19426, n19427, n19428, n19429, n19430, n19431, n19432, n19433,
         n19434, n19435, n19436, n19437, n19438, n19439, n19440, n19441,
         n19442, n19443, n19444, n19445, n19446, n19447, n19448, n19449,
         n19450, n19451, n19452, n19453, n19454, n19455, n19456, n19457,
         n19458, n19459, n19460, n19461, n19462, n19463, n19464, n19465,
         n19466, n19467, n19468, n19469, n19470, n19471, n19472, n19473,
         n19474, n19475, n19476, n19477, n19478, n19479, n19480, n19481,
         n19482, n19483, n19484, n19485, n19486, n19487, n19488, n19489,
         n19490, n19491, n19492, n19493, n19494, n19495, n19496, n19497,
         n19498, n19499, n19500, n19501, n19502, n19503, n19504, n19505,
         n19506, n19507, n19508, n19509, n19510, n19511, n19512, n19513,
         n19514, n19515, n19516, n19517, n19518, n19519, n19520, n19521,
         n19522, n19523, n19524, n19525, n19526, n19527, n19528, n19529,
         n19530, n19531, n19532, n19533, n19534, n19535, n19536, n19537,
         n19538, n19539, n19540, n19541, n19542, n19543, n19544, n19545,
         n19546, n19547, n19548, n19549, n19550, n19551, n19552, n19553,
         n19554, n19555, n19556, n19557, n19558, n19559, n19560, n19561,
         n19562, n19563, n19564, n19565, n19566, n19567, n19568, n19569,
         n19570, n19571, n19572, n19573, n19574, n19575, n19576, n19577,
         n19578, n19579, n19580, n19581, n19582, n19583, n19584, n19585,
         n19586, n19587, n19588, n19589, n19590, n19591, n19592, n19593,
         n19594, n19595, n19596, n19597, n19598, n19599, n19600, n19601,
         n19602, n19603, n19604, n19605, n19606, n19607, n19608, n19609,
         n19610, n19611, n19612, n19613, n19614, n19615, n19616, n19617,
         n19618, n19619, n19620, n19621, n19622, n19623, n19624, n19625,
         n19626, n19627, n19628, n19629, n19630, n19631, n19632, n19633,
         n19634, n19635, n19636, n19637, n19638, n19639, n19640, n19641,
         n19642, n19643, n19644, n19645, n19646, n19647, n19648, n19649,
         n19650, n19651, n19652, n19653, n19654, n19655, n19656, n19657,
         n19658, n19659, n19660, n19661, n19662, n19663, n19664, n19665,
         n19666, n19667, n19668, n19669, n19670, n19671, n19672, n19673,
         n19674, n19675, n19676, n19677, n19678, n19679, n19680, n19681,
         n19682, n19683, n19684, n19685, n19686, n19687, n19688, n19689,
         n19690, n19691, n19692, n19693, n19694, n19695, n19696, n19697,
         n19698, n19699, n19700, n19701, n19702, n19703, n19704, n19705,
         n19706, n19707, n19708, n19709, n19710, n19711, n19712, n19713,
         n19714, n19715, n19716, n19717, n19718, n19719, n19720, n19721,
         n19722, n19723, n19724, n19725, n19726, n19727, n19728, n19729,
         n19730, n19731, n19732, n19733, n19734, n19735, n19736, n19737,
         n19738, n19739, n19740, n19741, n19742, n19743, n19744, n19745,
         n19746, n19747, n19748, n19749, n19750, n19751, n19752, n19753,
         n19754, n19755, n19756, n19757, n19758, n19759, n19760, n19761,
         n19762, n19763, n19764, n19765, n19766, n19767, n19768, n19769,
         n19770, n19771, n19772, n19773, n19774, n19775, n19776, n19777,
         n19778, n19779, n19780, n19781, n19782, n19783, n19784, n19785,
         n19786, n19787, n19788, n19789, n19790, n19791, n19792, n19793,
         n19794, n19795, n19796, n19797, n19798, n19799, n19800, n19801,
         n19802, n19803, n19804, n19805, n19806, n19807, n19808, n19809,
         n19810, n19811, n19812, n19813, n19814, n19815, n19816, n19817,
         n19818, n19819, n19820, n19821, n19822, n19823, n19824, n19825,
         n19826, n19827, n19828, n19829, n19830, n19831, n19832, n19833,
         n19834, n19835, n19836, n19837, n19838, n19839, n19840, n19841,
         n19842, n19843, n19844, n19845, n19846, n19847, n19848, n19849,
         n19850, n19851, n19852, n19853, n19854, n19855, n19856, n19857,
         n19858, n19859, n19860, n19861, n19862, n19863, n19864, n19865,
         n19866, n19867, n19868, n19869, n19870, n19871, n19872, n19873,
         n19874, n19875, n19876, n19877, n19878, n19879, n19880, n19881,
         n19882, n19883, n19884, n19885, n19886, n19887, n19888, n19889,
         n19890, n19891, n19892, n19893, n19894, n19895, n19896, n19897,
         n19898, n19899, n19900, n19901, n19902, n19903, n19904, n19905,
         n19906, n19907, n19908, n19909, n19910, n19911, n19912, n19913,
         n19914, n19915, n19916, n19917, n19918, n19919, n19920, n19921,
         n19922, n19923, n19924, n19925, n19926, n19927, n19928, n19929,
         n19930, n19931, n19932, n19933, n19934, n19935, n19936, n19937,
         n19938, n19939, n19940, n19941, n19942, n19943, n19944, n19945,
         n19946, n19947, n19948, n19949, n19950, n19951, n19952, n19953,
         n19954, n19955, n19956, n19957, n19958, n19959, n19960, n19961,
         n19962, n19963, n19964, n19965, n19966, n19967, n19968, n19969,
         n19970, n19971, n19972, n19973, n19974, n19975, n19976, n19977,
         n19978, n19979, n19980, n19981, n19982, n19983, n19984, n19985,
         n19986, n19987, n19988, n19989, n19990, n19991, n19992, n19993,
         n19994, n19995, n19996, n19997, n19998, n19999, n20000, n20001,
         n20002, n20003, n20004, n20005, n20006, n20007, n20008, n20009,
         n20010, n20011, n20012, n20013, n20014, n20015, n20016, n20017,
         n20018, n20019, n20020, n20021, n20022, n20023, n20024, n20025,
         n20026, n20027, n20028, n20029, n20030, n20031, n20032, n20033,
         n20034, n20035, n20036, n20037, n20038, n20039, n20040, n20041,
         n20042, n20043, n20044, n20045, n20046, n20047, n20048, n20049,
         n20050, n20051, n20052, n20053, n20054, n20055, n20056, n20057,
         n20058, n20059, n20060, n20061, n20062, n20063, n20064, n20065,
         n20066, n20067, n20068, n20069, n20070, n20071, n20072, n20073,
         n20074, n20075, n20076, n20077, n20078, n20079, n20080, n20081,
         n20082, n20083, n20084, n20085, n20086, n20087, n20088, n20089,
         n20090, n20091, n20092, n20093, n20094, n20095, n20096, n20097,
         n20098, n20099, n20100, n20101, n20102, n20103, n20104, n20105,
         n20106, n20107, n20108, n20109, n20110, n20111, n20112, n20113,
         n20114, n20115, n20116, n20117, n20118, n20119, n20120, n20121,
         n20122, n20123, n20124, n20125, n20126, n20127, n20128, n20129,
         n20130, n20131, n20132, n20133, n20134, n20135, n20136, n20137,
         n20138, n20139, n20140, n20141, n20142, n20143, n20144, n20145,
         n20146, n20147, n20148, n20149, n20150, n20151, n20152, n20153,
         n20154, n20155, n20156, n20157, n20158, n20159, n20160, n20161,
         n20162, n20163, n20164, n20165, n20166, n20167, n20168, n20169,
         n20170, n20171, n20172, n20173, n20174, n20175, n20176, n20177,
         n20178, n20179, n20180, n20181, n20182, n20183, n20184, n20185,
         n20186, n20187, n20188, n20189, n20190, n20191, n20192, n20193,
         n20194, n20195, n20196, n20197, n20198, n20199, n20200, n20201,
         n20202, n20203, n20204, n20205, n20206, n20207, n20208, n20209,
         n20210, n20211, n20212, n20213, n20214, n20215, n20216, n20217,
         n20218, n20219, n20220, n20221, n20222, n20223, n20224, n20225,
         n20226, n20227, n20228, n20229, n20230, n20231, n20232, n20233,
         n20234, n20235, n20236, n20237, n20238, n20239, n20240, n20241,
         n20242, n20243, n20244, n20245, n20246, n20247, n20248, n20249,
         n20250, n20251, n20252, n20253, n20254, n20255, n20256, n20257,
         n20258, n20259, n20260, n20261, n20262, n20263, n20264, n20265,
         n20266, n20267, n20268, n20269, n20270, n20271, n20272, n20273,
         n20274, n20275, n20276, n20277, n20278, n20279, n20280, n20281,
         n20282, n20283, n20284, n20285, n20286, n20287, n20288, n20289,
         n20290, n20291, n20292, n20293, n20294, n20295, n20296, n20297,
         n20298, n20299, n20300, n20301, n20302, n20303, n20304, n20305,
         n20306, n20307, n20308, n20309, n20310, n20311, n20312, n20313,
         n20314, n20315, n20316, n20317, n20318, n20319, n20320, n20321,
         n20322, n20323, n20324, n20325, n20326, n20327, n20328, n20329,
         n20330, n20331, n20332, n20333, n20334, n20335, n20336, n20337,
         n20338, n20339, n20340, n20341, n20342, n20343, n20344, n20345,
         n20346, n20347, n20348, n20349, n20350, n20351, n20352, n20353,
         n20354, n20355, n20356, n20357, n20358, n20359, n20360, n20361,
         n20362, n20363, n20364, n20365, n20366, n20367, n20368, n20369,
         n20370, n20371, n20372, n20373, n20374, n20375, n20376, n20377,
         n20378, n20379, n20380, n20381, n20382, n20383, n20384, n20385,
         n20386, n20387, n20388, n20389, n20390, n20391, n20392, n20393,
         n20394, n20395, n20396, n20397, n20398, n20399, n20400, n20401,
         n20402, n20403, n20404, n20405, n20406, n20407, n20408, n20409,
         n20410, n20411, n20412, n20413, n20414, n20415, n20416, n20417,
         n20418, n20419, n20420, n20421, n20422, n20423, n20424, n20425,
         n20426, n20427, n20428, n20429, n20430, n20431, n20432, n20433,
         n20434, n20435, n20436, n20437, n20438, n20439, n20440, n20441,
         n20442, n20443, n20444, n20445, n20446, n20447, n20448, n20449,
         n20450, n20451, n20452, n20453, n20454, n20455, n20456, n20457,
         n20458, n20459, n20460, n20461, n20462, n20463, n20464, n20465,
         n20466, n20467, n20468, n20469, n20470, n20471, n20472, n20473,
         n20474, n20475, n20476, n20477, n20478, n20479, n20480, n20481,
         n20482, n20483, n20484, n20485, n20486, n20487, n20488, n20489,
         n20490, n20491, n20492, n20493, n20494, n20495, n20496, n20497,
         n20498, n20499, n20500, n20501, n20502, n20503, n20504, n20505,
         n20506, n20507, n20508, n20509, n20510, n20511, n20512, n20513,
         n20514, n20515, n20516, n20517, n20518, n20519, n20520, n20521,
         n20522, n20523, n20524, n20525, n20526, n20527, n20528, n20529,
         n20530, n20531, n20532, n20533, n20534, n20535, n20536, n20537,
         n20538, n20539, n20540, n20541, n20542, n20543, n20544, n20545,
         n20546, n20547, n20548, n20549, n20550, n20551, n20552, n20553,
         n20554, n20555, n20556, n20557, n20558, n20559, n20560, n20561,
         n20562, n20563, n20564, n20565, n20566, n20567, n20568, n20569,
         n20570, n20571, n20572, n20573, n20574, n20575, n20576, n20577,
         n20578, n20579, n20580, n20581, n20582, n20583, n20584, n20585,
         n20586, n20587, n20588, n20589, n20590, n20591, n20592, n20593,
         n20594, n20595, n20596, n20597, n20598, n20599, n20600, n20601,
         n20602, n20603, n20604, n20605, n20606, n20607, n20608, n20609,
         n20610, n20611, n20612, n20613, n20614, n20615, n20616, n20617,
         n20618, n20619, n20620, n20621, n20622, n20623, n20624, n20625,
         n20626, n20627, n20628, n20629, n20630, n20631, n20632, n20633,
         n20634, n20635, n20636, n20637, n20638, n20639, n20640, n20641,
         n20642, n20643, n20644, n20645, n20646, n20647, n20648, n20649,
         n20650, n20651, n20652, n20653, n20654, n20655, n20656, n20657,
         n20658, n20659, n20660, n20661, n20662, n20663, n20664, n20665,
         n20666, n20667, n20668, n20669, n20671, n20672, n20673, n20674,
         n20675, n20676, n20677, n20678, n20679, n20680, n20681, n20682,
         n20683, n20684, n20685, n20686, n20687, n20688, n20689, n20690,
         n20691, n20692, n20693, n20694, n20695, n20696, n20697, n20698,
         n20699, n20700, n20701, n20702, n20703, n20704, n20705, n20706,
         n20707, n20708, n20709, n20710, n20711, n20712, n20713, n20714,
         n20715, n20716, n20717, n20718, n20719, n20720, n20721, n20722,
         n20723, n20724, n20725, n20726, n20727, n20728, n20729, n20730,
         n20731, n20732, n20733, n20734, n20735, n20736, n20737, n20738,
         n20739, n20740, n20741, n20742, n20743, n20744, n20745, n20746,
         n20747, n20748, n20749, n20750, n20751, n20752, n20753, n20754,
         n20755, n20756, n20757, n20758, n20759, n20760, n20761, n20762,
         n20763, n20764, n20765, n20766, n20767, n20768, n20769, n20770,
         n20771, n20772, n20773, n20774, n20775, n20776, n20777, n20778,
         n20779, n20780, n20781, n20782, n20783, n20784, n20785, n20786,
         n20787, n20788, n20789, n20790, n20791, n20792, n20793, n20794,
         n20795, n20796, n20797, n20798, n20799, n20800, n20801, n20802,
         n20803, n20804, n20805, n20806, n20807, n20808, n20809, n20810,
         n20811, n20812, n20813, n20814, n20815, n20816, n20817, n20818,
         n20819, n20820, n20821, n20822, n20823, n20824, n20825, n20826,
         n20827, n20828, n20829, n20830, n20831, n20832, n20833, n20834,
         n20835, n20836, n20837, n20838, n20839, n20840, n20841, n20842,
         n20843, n20844, n20845, n20846, n20847, n20848, n20849, n20850,
         n20851, n20852, n20853, n20854, n20855, n20856, n20857, n20858,
         n20859, n20860, n20861, n20862, n20863, n20864, n20865, n20866,
         n20867, n20868, n20869, n20870, n20871, n20872, n20873, n20874,
         n20875, n20876, n20877, n20878, n20879, n20880, n20881, n20882,
         n20883, n20884, n20885, n20886, n20887, n20888, n20889, n20890,
         n20891, n20892, n20893, n20894, n20895, n20896, n20897, n20898,
         n20899, n20900, n20901, n20902, n20903, n20904, n20905, n20906,
         n20907, n20908, n20909, n20910, n20911, n20912, n20913, n20914,
         n20915, n20916, n20917, n20918, n20919, n20920, n20921, n20922,
         n20923, n20924, n20925, n20926, n20927, n20928, n20929, n20930,
         n20931, n20932, n20933, n20934, n20935, n20936, n20937, n20938,
         n20939, n20940, n20941, n20942, n20943, n20944, n20945, n20946,
         n20947, n20948, n20949, n20950, n20951, n20952, n20953, n20954,
         n20955, n20956, n20957, n20958, n20959, n20960, n20961, n20962,
         n20963, n20964, n20965, n20966, n20967, n20968, n20969, n20970,
         n20971, n20972, n20973, n20974, n20975, n20976, n20977, n20978,
         n20979, n20980, n20981, n20982, n20983, n20984, n20985, n20986,
         n20987, n20988, n20989, n20990, n20991, n20992, n20993, n20994,
         n20995, n20996, n20997, n20998, n20999, n21000, n21001, n21002,
         n21003, n21004, n21005, n21006, n21007, n21008, n21009, n21010,
         n21011, n21012, n21013, n21014, n21015, n21016, n21017, n21018,
         n21019, n21020, n21021, n21022, n21023, n21024, n21025, n21026,
         n21027, n21028, n21029, n21030, n21031, n21032, n21033, n21034,
         n21035, n21036, n21037, n21038, n21039, n21040, n21041, n21042,
         n21043, n21044, n21045, n21046, n21047, n21048, n21049, n21050,
         n21051, n21052, n21053, n21054, n21055, n21056, n21057, n21058,
         n21059, n21060, n21061, n21062, n21063, n21064, n21065, n21066,
         n21067, n21068, n21069, n21070, n21071, n21072, n21073, n21074,
         n21075, n21076, n21077, n21078, n21079, n21080, n21081, n21082,
         n21083, n21084, n21085, n21086, n21087, n21088, n21089, n21090,
         n21091, n21092, n21093, n21094, n21095, n21096, n21097, n21098,
         n21099, n21100, n21101, n21102, n21103, n21104, n21105, n21106,
         n21107, n21108, n21109, n21110, n21111, n21112, n21113, n21114,
         n21115, n21116, n21117, n21118, n21119, n21120, n21121, n21122,
         n21123, n21124, n21125, n21126, n21127, n21128, n21129, n21130,
         n21131, n21132, n21133, n21134, n21135, n21136, n21137, n21138,
         n21139, n21140, n21141, n21142, n21143, n21144, n21145, n21146,
         n21147, n21148, n21149, n21150, n21151, n21152, n21153, n21154,
         n21155, n21156, n21157, n21158, n21159, n21160, n21161, n21162,
         n21163, n21164, n21165, n21166, n21167, n21168, n21169, n21170,
         n21171, n21172, n21173, n21174, n21175, n21176, n21177, n21178,
         n21179, n21180, n21181, n21182, n21183, n21184, n21185, n21186,
         n21187, n21188, n21189, n21190, n21191, n21192, n21193, n21194,
         n21195, n21196, n21197, n21198, n21199, n21200, n21201, n21202,
         n21203, n21204, n21205, n21206, n21207, n21208, n21209, n21210,
         n21211, n21212, n21213, n21214, n21215, n21216, n21217, n21218;

  AND2_X1 U11271 ( .A1(n20022), .A2(n13965), .ZN(n20034) );
  CLKBUF_X2 U11272 ( .A(n11335), .Z(n10053) );
  NAND2_X1 U11273 ( .A1(n12446), .A2(n15612), .ZN(n15613) );
  INV_X1 U11274 ( .A(n10609), .ZN(n11096) );
  NOR2_X1 U11275 ( .A1(n13167), .A2(n13166), .ZN(n18886) );
  CLKBUF_X1 U11276 ( .A(n11792), .Z(n11958) );
  BUF_X2 U11277 ( .A(n11175), .Z(n13396) );
  CLKBUF_X2 U11278 ( .A(n11250), .Z(n9835) );
  INV_X2 U11279 ( .A(n11180), .ZN(n11197) );
  NAND2_X1 U11280 ( .A1(n16751), .A2(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n16750) );
  CLKBUF_X3 U11281 ( .A(n13058), .Z(n9839) );
  AND2_X1 U11282 ( .A1(n12945), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11680) );
  AND2_X1 U11283 ( .A1(n12799), .A2(n11654), .ZN(n12789) );
  AND2_X1 U11284 ( .A1(n12929), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11727) );
  CLKBUF_X2 U11285 ( .A(n11766), .Z(n12781) );
  INV_X1 U11286 ( .A(n17136), .ZN(n17217) );
  CLKBUF_X2 U11287 ( .A(n10980), .Z(n9863) );
  CLKBUF_X2 U11288 ( .A(n10498), .Z(n11023) );
  CLKBUF_X2 U11289 ( .A(n10710), .Z(n10925) );
  CLKBUF_X2 U11290 ( .A(n10467), .Z(n11080) );
  NOR2_X1 U11291 ( .A1(n13015), .A2(n13014), .ZN(n13058) );
  CLKBUF_X2 U11292 ( .A(n10400), .Z(n11057) );
  NAND4_X1 U11293 ( .A1(n11440), .A2(n12434), .A3(n9874), .A4(n12431), .ZN(
        n11472) );
  BUF_X1 U11294 ( .A(n9894), .Z(n13781) );
  AND2_X1 U11295 ( .A1(n20177), .A2(n13376), .ZN(n13809) );
  INV_X1 U11296 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n17888) );
  CLKBUF_X3 U11297 ( .A(n10423), .Z(n9854) );
  INV_X1 U11298 ( .A(n12571), .ZN(n20177) );
  OR2_X1 U11299 ( .A1(n10299), .A2(n10298), .ZN(n10474) );
  AND2_X2 U11300 ( .A1(n10284), .A2(n13744), .ZN(n9867) );
  AND2_X1 U11301 ( .A1(n13744), .A2(n13716), .ZN(n10467) );
  AND2_X1 U11302 ( .A1(n10292), .A2(n10290), .ZN(n10387) );
  AND2_X1 U11303 ( .A1(n13744), .A2(n10291), .ZN(n10710) );
  AND2_X1 U11304 ( .A1(n10291), .A2(n10293), .ZN(n10596) );
  AND2_X1 U11305 ( .A1(n10283), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13743) );
  CLKBUF_X2 U11306 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n15752) );
  INV_X1 U11308 ( .A(n21218), .ZN(n9828) );
  AND2_X1 U11309 ( .A1(n10419), .A2(n14519), .ZN(n12560) );
  AND2_X1 U11310 ( .A1(n10474), .A2(n11106), .ZN(n11147) );
  NOR2_X2 U11311 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11655) );
  AND2_X1 U11312 ( .A1(n10290), .A2(n13716), .ZN(n10330) );
  AND2_X1 U11313 ( .A1(n10417), .A2(n14519), .ZN(n13392) );
  AND4_X1 U11314 ( .A1(n10311), .A2(n10310), .A3(n10309), .A4(n10308), .ZN(
        n10317) );
  NAND2_X1 U11315 ( .A1(n10436), .A2(n10435), .ZN(n10497) );
  AND2_X1 U11316 ( .A1(n12799), .A2(n11655), .ZN(n11668) );
  AND2_X1 U11317 ( .A1(n12828), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11771) );
  INV_X1 U11318 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11651) );
  NAND2_X1 U11319 ( .A1(n18854), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13012) );
  NOR2_X2 U11320 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10291) );
  AND2_X1 U11321 ( .A1(n12439), .A2(n11470), .ZN(n13563) );
  INV_X1 U11322 ( .A(n11451), .ZN(n12412) );
  NOR2_X1 U11323 ( .A1(n13012), .A2(n13010), .ZN(n13065) );
  AND2_X1 U11324 ( .A1(n20168), .A2(n9854), .ZN(n15891) );
  INV_X1 U11325 ( .A(n20294), .ZN(n10576) );
  INV_X1 U11327 ( .A(n19079), .ZN(n11335) );
  NAND2_X1 U11328 ( .A1(n12269), .A2(n12194), .ZN(n12192) );
  NOR2_X1 U11329 ( .A1(n14263), .A2(n11893), .ZN(n14266) );
  NAND2_X1 U11330 ( .A1(n11452), .A2(n11451), .ZN(n11794) );
  AND2_X1 U11331 ( .A1(n13568), .A2(n13569), .ZN(n13567) );
  CLKBUF_X2 U11332 ( .A(n11436), .Z(n19297) );
  NOR2_X2 U11333 ( .A1(n9854), .A2(n9858), .ZN(n13959) );
  INV_X1 U11334 ( .A(n16023), .ZN(n19992) );
  NAND2_X1 U11335 ( .A1(n10590), .A2(n10589), .ZN(n13875) );
  OR2_X1 U11336 ( .A1(n15596), .A2(n15280), .ZN(n15573) );
  NOR2_X1 U11337 ( .A1(n13863), .A2(n10179), .ZN(n14223) );
  NAND2_X1 U11338 ( .A1(n16580), .A2(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n17586) );
  NOR2_X1 U11339 ( .A1(n18024), .A2(n17783), .ZN(n17690) );
  NAND2_X1 U11340 ( .A1(n18118), .A2(n18692), .ZN(n18139) );
  XNOR2_X1 U11341 ( .A(n13113), .B(n13112), .ZN(n17878) );
  INV_X1 U11342 ( .A(n14030), .ZN(n14029) );
  AOI221_X1 U11343 ( .B1(P1_REIP_REG_23__SCAN_IN), .B2(n15951), .C1(n15950), 
        .C2(n15951), .A(n15949), .ZN(n15952) );
  INV_X1 U11344 ( .A(n20034), .ZN(n20006) );
  OAI21_X1 U11345 ( .B1(n14682), .B2(n14680), .A(n14681), .ZN(n15948) );
  INV_X1 U11346 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n19917) );
  INV_X2 U11347 ( .A(n19937), .ZN(n19940) );
  INV_X1 U11348 ( .A(n17767), .ZN(n17750) );
  INV_X1 U11349 ( .A(n17218), .ZN(n17080) );
  BUF_X1 U11350 ( .A(n11435), .Z(n14035) );
  NAND2_X1 U11351 ( .A1(n14674), .A2(n10201), .ZN(n9829) );
  AND2_X1 U11352 ( .A1(n13743), .A2(n13716), .ZN(n10400) );
  MUX2_X2 U11353 ( .A(n12328), .B(n12306), .S(n12308), .Z(n12285) );
  AND3_X2 U11354 ( .A1(n11421), .A2(n11420), .A3(n12985), .ZN(n11461) );
  NOR2_X2 U11355 ( .A1(n14697), .A2(n14698), .ZN(n9960) );
  OAI21_X1 U11356 ( .B1(n14663), .B2(n20145), .A(n10270), .ZN(n14500) );
  NAND2_X2 U11357 ( .A1(n12420), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11508) );
  OAI21_X2 U11358 ( .B1(n14476), .B2(n9919), .A(n9999), .ZN(n9998) );
  NAND2_X2 U11359 ( .A1(n13072), .A2(n10272), .ZN(n17421) );
  AND2_X2 U11360 ( .A1(n11339), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11653) );
  NAND2_X2 U11362 ( .A1(n11471), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11494) );
  NAND2_X2 U11363 ( .A1(n11466), .A2(n11465), .ZN(n11471) );
  NOR2_X1 U11364 ( .A1(n13015), .A2(n13012), .ZN(n13047) );
  AND2_X4 U11365 ( .A1(n9947), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10292) );
  AND2_X2 U11366 ( .A1(n11654), .A2(n15754), .ZN(n9830) );
  NOR2_X2 U11367 ( .A1(n15648), .A2(n11920), .ZN(n15632) );
  NAND2_X2 U11368 ( .A1(n13563), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11543) );
  AND2_X2 U11369 ( .A1(n10211), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n15743) );
  CLKBUF_X1 U11370 ( .A(n10342), .Z(n9831) );
  AND2_X1 U11371 ( .A1(n13743), .A2(n10291), .ZN(n10342) );
  CLKBUF_X1 U11372 ( .A(n10342), .Z(n11065) );
  NOR2_X1 U11374 ( .A1(n13015), .A2(n13009), .ZN(n17218) );
  XNOR2_X2 U11375 ( .A(n12176), .B(n12425), .ZN(n14330) );
  INV_X1 U11376 ( .A(n12684), .ZN(n14243) );
  INV_X1 U11377 ( .A(n14437), .ZN(n13160) );
  BUF_X8 U11378 ( .A(n13160), .Z(n9849) );
  XNOR2_X2 U11379 ( .A(n12599), .B(n12593), .ZN(n20094) );
  NAND2_X2 U11380 ( .A1(n13931), .A2(n12592), .ZN(n12599) );
  NAND2_X1 U11381 ( .A1(n15308), .A2(n9899), .ZN(n12402) );
  INV_X1 U11382 ( .A(n12338), .ZN(n12062) );
  INV_X4 U11383 ( .A(n9913), .ZN(n16081) );
  NAND2_X1 U11384 ( .A1(n10240), .A2(n10239), .ZN(n17705) );
  NAND2_X1 U11385 ( .A1(n17809), .A2(n17818), .ZN(n17817) );
  INV_X1 U11387 ( .A(n14243), .ZN(n10247) );
  AND2_X1 U11388 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n17161), .ZN(n15796) );
  AND2_X1 U11389 ( .A1(n12192), .A2(n11746), .ZN(n12213) );
  NOR2_X1 U11390 ( .A1(n18736), .A2(n16587), .ZN(n16939) );
  INV_X4 U11391 ( .A(n12102), .ZN(n12417) );
  NAND2_X1 U11392 ( .A1(n13477), .A2(n9846), .ZN(n11184) );
  NAND3_X1 U11393 ( .A1(n13249), .A2(n13248), .A3(n13247), .ZN(n13274) );
  INV_X2 U11394 ( .A(n10474), .ZN(n20182) );
  INV_X1 U11395 ( .A(n10417), .ZN(n10422) );
  INV_X4 U11396 ( .A(n16370), .ZN(n12392) );
  INV_X2 U11397 ( .A(n11451), .ZN(n11788) );
  AND4_X1 U11398 ( .A1(n10391), .A2(n10390), .A3(n10389), .A4(n10388), .ZN(
        n10408) );
  AND4_X1 U11399 ( .A1(n10395), .A2(n10394), .A3(n10393), .A4(n10392), .ZN(
        n10407) );
  AND4_X1 U11400 ( .A1(n10399), .A2(n10398), .A3(n10397), .A4(n10396), .ZN(
        n10406) );
  AND4_X1 U11401 ( .A1(n10404), .A2(n10403), .A3(n10402), .A4(n10401), .ZN(
        n10405) );
  AND2_X2 U11402 ( .A1(n11652), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11777) );
  CLKBUF_X2 U11403 ( .A(n13066), .Z(n17098) );
  BUF_X2 U11404 ( .A(n13066), .Z(n17199) );
  CLKBUF_X2 U11405 ( .A(n13088), .Z(n17192) );
  CLKBUF_X1 U11406 ( .A(n11427), .Z(n12941) );
  CLKBUF_X1 U11407 ( .A(n10510), .Z(n9833) );
  CLKBUF_X2 U11408 ( .A(n11078), .Z(n11064) );
  INV_X1 U11409 ( .A(n20814), .ZN(n9834) );
  INV_X2 U11410 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n18718) );
  NOR2_X4 U11411 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10290) );
  AND2_X2 U11413 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10293) );
  XNOR2_X1 U11414 ( .A(n12505), .B(n12504), .ZN(n12531) );
  OAI21_X1 U11415 ( .B1(n14475), .B2(n14474), .A(n10039), .ZN(n14819) );
  NAND2_X1 U11416 ( .A1(n10040), .A2(n9927), .ZN(n10039) );
  OR2_X1 U11417 ( .A1(n12534), .A2(n16295), .ZN(n12514) );
  NAND2_X1 U11418 ( .A1(n14839), .A2(n14963), .ZN(n14475) );
  INV_X1 U11419 ( .A(n10210), .ZN(n14556) );
  OAI21_X1 U11420 ( .B1(n15420), .B2(n15419), .A(n15366), .ZN(n15410) );
  AOI21_X1 U11421 ( .B1(n15300), .B2(n12403), .A(n12402), .ZN(n12407) );
  NAND2_X1 U11422 ( .A1(n14848), .A2(n14838), .ZN(n14839) );
  OAI21_X1 U11423 ( .B1(n14580), .B2(n14582), .A(n14581), .ZN(n14842) );
  NAND2_X1 U11424 ( .A1(n10006), .A2(n12651), .ZN(n14838) );
  NOR2_X1 U11425 ( .A1(n15629), .A2(n15626), .ZN(n15429) );
  OR2_X1 U11426 ( .A1(n15675), .A2(n15413), .ZN(n16241) );
  INV_X1 U11427 ( .A(n15398), .ZN(n15675) );
  AOI21_X1 U11428 ( .B1(n15170), .B2(n12919), .A(n15166), .ZN(n15161) );
  INV_X1 U11429 ( .A(n12357), .ZN(n9988) );
  NOR2_X1 U11430 ( .A1(n12902), .A2(n12904), .ZN(n15172) );
  NAND2_X2 U11431 ( .A1(n14934), .A2(n12638), .ZN(n14891) );
  OR2_X1 U11432 ( .A1(n13148), .A2(n17757), .ZN(n15907) );
  NOR2_X1 U11433 ( .A1(n12901), .A2(n12900), .ZN(n12904) );
  AND2_X1 U11434 ( .A1(n16447), .A2(n10238), .ZN(n13148) );
  NOR2_X1 U11435 ( .A1(n15177), .A2(n10268), .ZN(n12901) );
  NAND2_X1 U11436 ( .A1(n13147), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n17561) );
  NOR2_X1 U11437 ( .A1(n10273), .A2(n10148), .ZN(n10147) );
  NOR2_X1 U11438 ( .A1(n17570), .A2(n13145), .ZN(n13147) );
  NAND2_X1 U11439 ( .A1(n12349), .A2(n12348), .ZN(n14220) );
  NAND2_X1 U11440 ( .A1(n10128), .A2(n10126), .ZN(n14163) );
  NAND2_X1 U11441 ( .A1(n12124), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n14089) );
  AOI21_X1 U11442 ( .B1(n10035), .B2(n10038), .A(n10033), .ZN(n10032) );
  NAND2_X1 U11443 ( .A1(n12168), .A2(n19059), .ZN(n12176) );
  OAI21_X1 U11444 ( .B1(n10172), .B2(n15196), .A(n10171), .ZN(n12862) );
  NAND2_X1 U11445 ( .A1(n12599), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12600) );
  AND2_X1 U11446 ( .A1(n16091), .A2(n10036), .ZN(n10035) );
  NOR2_X1 U11447 ( .A1(n10130), .A2(n10131), .ZN(n10127) );
  NOR2_X1 U11448 ( .A1(n10005), .A2(n14926), .ZN(n16064) );
  NAND2_X1 U11449 ( .A1(n14101), .A2(n12417), .ZN(n12123) );
  AND2_X1 U11450 ( .A1(n9983), .A2(n12338), .ZN(n14101) );
  OR2_X1 U11451 ( .A1(n12629), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16091) );
  INV_X1 U11452 ( .A(n16099), .ZN(n10130) );
  OR2_X1 U11453 ( .A1(n14247), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12636) );
  NAND2_X1 U11454 ( .A1(n13933), .A2(n13932), .ZN(n13931) );
  OR2_X1 U11455 ( .A1(n14922), .A2(n14925), .ZN(n10005) );
  XNOR2_X1 U11456 ( .A(n12591), .B(n12584), .ZN(n13933) );
  NOR2_X1 U11457 ( .A1(n15195), .A2(n15197), .ZN(n15196) );
  NAND2_X1 U11458 ( .A1(n10235), .A2(n10228), .ZN(n10227) );
  NAND2_X2 U11459 ( .A1(n12612), .A2(n12632), .ZN(n9913) );
  OAI21_X1 U11460 ( .B1(n12247), .B2(n12246), .A(n10236), .ZN(n10235) );
  XNOR2_X1 U11461 ( .A(n12582), .B(n20135), .ZN(n13777) );
  NAND2_X1 U11462 ( .A1(n10669), .A2(n10668), .ZN(n12612) );
  AND2_X1 U11463 ( .A1(n12100), .A2(n11813), .ZN(n10245) );
  AND2_X1 U11464 ( .A1(n10541), .A2(n10558), .ZN(n13765) );
  OR3_X2 U11465 ( .A1(n12245), .A2(n15385), .A3(n15367), .ZN(n12246) );
  AND2_X1 U11466 ( .A1(n12099), .A2(n12098), .ZN(n12100) );
  NAND2_X1 U11467 ( .A1(n13704), .A2(n12577), .ZN(n12582) );
  NAND2_X1 U11468 ( .A1(n13131), .A2(n17817), .ZN(n17754) );
  AND4_X1 U11469 ( .A1(n12025), .A2(n12024), .A3(n12023), .A4(n12022), .ZN(
        n12026) );
  NAND2_X1 U11470 ( .A1(n13703), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13704) );
  NAND2_X1 U11471 ( .A1(n10576), .A2(n10577), .ZN(n10628) );
  XNOR2_X1 U11472 ( .A(n12575), .B(n13382), .ZN(n13703) );
  NAND2_X1 U11473 ( .A1(n10030), .A2(n10029), .ZN(n10537) );
  AND2_X1 U11474 ( .A1(n14733), .A2(n14732), .ZN(n14735) );
  NAND2_X1 U11475 ( .A1(n12569), .A2(n12568), .ZN(n12575) );
  NOR2_X1 U11476 ( .A1(n17816), .A2(n18144), .ZN(n17815) );
  NAND2_X1 U11477 ( .A1(n14243), .A2(n12008), .ZN(n12063) );
  NAND2_X1 U11478 ( .A1(n11988), .A2(n13628), .ZN(n19508) );
  OAI22_X1 U11479 ( .A1(n12017), .A2(n19482), .B1(n12080), .B2(n12016), .ZN(
        n12018) );
  NOR2_X1 U11480 ( .A1(n20294), .A2(n9930), .ZN(n10010) );
  NAND2_X1 U11481 ( .A1(n12008), .A2(n10247), .ZN(n12064) );
  NAND2_X1 U11482 ( .A1(n14243), .A2(n11988), .ZN(n12071) );
  NAND2_X1 U11483 ( .A1(n12021), .A2(n14243), .ZN(n12141) );
  NAND2_X1 U11484 ( .A1(n14053), .A2(n10282), .ZN(n19542) );
  CLKBUF_X1 U11485 ( .A(n12554), .Z(n14806) );
  NAND2_X1 U11486 ( .A1(n12020), .A2(n14243), .ZN(n19452) );
  NAND2_X1 U11487 ( .A1(n12020), .A2(n13628), .ZN(n14124) );
  NAND2_X1 U11488 ( .A1(n12014), .A2(n13842), .ZN(n19482) );
  NAND2_X1 U11489 ( .A1(n13842), .A2(n11994), .ZN(n19304) );
  NAND2_X1 U11490 ( .A1(n13842), .A2(n12004), .ZN(n19358) );
  XNOR2_X1 U11491 ( .A(n10533), .B(n10531), .ZN(n10542) );
  NOR2_X1 U11492 ( .A1(n20047), .A2(n20811), .ZN(n20071) );
  NAND2_X1 U11493 ( .A1(n9997), .A2(n10453), .ZN(n10462) );
  INV_X1 U11494 ( .A(n10161), .ZN(n19098) );
  NAND2_X1 U11495 ( .A1(n10190), .A2(n10189), .ZN(n10533) );
  NAND2_X1 U11496 ( .A1(n12200), .A2(n11748), .ZN(n12219) );
  INV_X2 U11497 ( .A(n17375), .ZN(n17413) );
  AND2_X1 U11498 ( .A1(n13998), .A2(n13991), .ZN(n14076) );
  NOR2_X2 U11499 ( .A1(n16589), .A2(n18139), .ZN(n18681) );
  NAND2_X1 U11500 ( .A1(n10460), .A2(n10459), .ZN(n10461) );
  NAND2_X1 U11501 ( .A1(n11486), .A2(n11485), .ZN(n11985) );
  AOI221_X1 U11502 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(n16403), .C1(n19928), .C2(
        n16403), .A(n19747), .ZN(n19925) );
  NAND2_X1 U11503 ( .A1(n11980), .A2(n11979), .ZN(n11982) );
  INV_X1 U11504 ( .A(n11968), .ZN(n11984) );
  NAND2_X1 U11505 ( .A1(n15803), .A2(n15815), .ZN(n18699) );
  AND2_X1 U11506 ( .A1(n11491), .A2(n11490), .ZN(n11968) );
  NOR2_X1 U11507 ( .A1(n12175), .A2(n10074), .ZN(n12191) );
  NAND2_X1 U11508 ( .A1(n10413), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10433) );
  NOR2_X1 U11509 ( .A1(n13813), .A2(n9953), .ZN(n9952) );
  NOR2_X1 U11510 ( .A1(n12167), .A2(n12166), .ZN(n12173) );
  NOR2_X2 U11511 ( .A1(n17393), .A2(n13126), .ZN(n17818) );
  XNOR2_X1 U11512 ( .A(n13567), .B(n11797), .ZN(n13551) );
  AND2_X1 U11513 ( .A1(n10549), .A2(n10192), .ZN(n10191) );
  AND3_X1 U11514 ( .A1(n10057), .A2(n12103), .A3(n10056), .ZN(n10055) );
  NAND2_X1 U11515 ( .A1(n10440), .A2(n10424), .ZN(n13403) );
  AND2_X1 U11516 ( .A1(n10441), .A2(n13390), .ZN(n13711) );
  NAND2_X1 U11517 ( .A1(n10420), .A2(n13618), .ZN(n10440) );
  OAI21_X1 U11518 ( .B1(n11934), .B2(n12331), .A(n11787), .ZN(n13568) );
  NAND2_X1 U11519 ( .A1(n11179), .A2(n11178), .ZN(n11183) );
  AND2_X1 U11520 ( .A1(n11800), .A2(n11786), .ZN(n11787) );
  OR2_X1 U11521 ( .A1(n11184), .A2(P1_EBX_REG_1__SCAN_IN), .ZN(n11179) );
  OR2_X1 U11522 ( .A1(n13709), .A2(n13373), .ZN(n13386) );
  CLKBUF_X2 U11524 ( .A(n11802), .Z(n11960) );
  AND2_X1 U11525 ( .A1(n13409), .A2(n13405), .ZN(n10441) );
  INV_X1 U11526 ( .A(n13809), .ZN(n13718) );
  AND2_X1 U11527 ( .A1(n11453), .A2(n11437), .ZN(n11963) );
  CLKBUF_X3 U11528 ( .A(n11443), .Z(n19271) );
  AND2_X1 U11529 ( .A1(n12376), .A2(n10253), .ZN(n11453) );
  INV_X1 U11530 ( .A(n11250), .ZN(n13477) );
  OAI211_X1 U11531 ( .C1(n13072), .C2(n13107), .A(n10220), .B(n10219), .ZN(
        n17901) );
  AND2_X2 U11532 ( .A1(n10423), .A2(n10421), .ZN(n13808) );
  OR2_X1 U11533 ( .A1(n11686), .A2(n11685), .ZN(n12059) );
  INV_X2 U11534 ( .A(n11443), .ZN(n13427) );
  AND2_X1 U11535 ( .A1(n11459), .A2(n11419), .ZN(n11420) );
  NAND4_X2 U11536 ( .A1(n11745), .A2(n11744), .A3(n11743), .A4(n11742), .ZN(
        n12102) );
  CLKBUF_X1 U11537 ( .A(n11637), .Z(n12308) );
  INV_X2 U11538 ( .A(n16509), .ZN(n16515) );
  CLKBUF_X1 U11539 ( .A(n11441), .Z(n19281) );
  INV_X1 U11540 ( .A(n11112), .ZN(n10418) );
  INV_X1 U11541 ( .A(n14519), .ZN(n20194) );
  AND2_X1 U11542 ( .A1(n11435), .A2(n11436), .ZN(n12376) );
  NAND2_X1 U11543 ( .A1(n11362), .A2(n11361), .ZN(n11441) );
  NOR2_X1 U11544 ( .A1(n13071), .A2(n13070), .ZN(n13072) );
  OR2_X1 U11545 ( .A1(n10509), .A2(n10508), .ZN(n12633) );
  NAND2_X1 U11546 ( .A1(n11350), .A2(n11349), .ZN(n11459) );
  NAND2_X1 U11547 ( .A1(n11387), .A2(n11386), .ZN(n11436) );
  OR2_X1 U11548 ( .A1(n10520), .A2(n10519), .ZN(n12570) );
  NAND4_X1 U11549 ( .A1(n10408), .A2(n10407), .A3(n10406), .A4(n10405), .ZN(
        n10421) );
  NAND4_X2 U11550 ( .A1(n10408), .A2(n10407), .A3(n10406), .A4(n10405), .ZN(
        n9858) );
  OR2_X2 U11551 ( .A1(n10364), .A2(n10363), .ZN(n14519) );
  NAND4_X1 U11552 ( .A1(n10384), .A2(n10383), .A3(n10382), .A4(n10381), .ZN(
        n10423) );
  AND4_X1 U11553 ( .A1(n10380), .A2(n10379), .A3(n10378), .A4(n10377), .ZN(
        n10381) );
  AND4_X1 U11554 ( .A1(n10307), .A2(n10306), .A3(n10305), .A4(n10304), .ZN(
        n10318) );
  AND4_X1 U11555 ( .A1(n10303), .A2(n10302), .A3(n10301), .A4(n10300), .ZN(
        n10319) );
  NOR2_X2 U11556 ( .A1(n20160), .A2(n20159), .ZN(n20161) );
  AND4_X1 U11557 ( .A1(n10368), .A2(n10367), .A3(n10366), .A4(n10365), .ZN(
        n10384) );
  AND4_X1 U11558 ( .A1(n10372), .A2(n10371), .A3(n10370), .A4(n10369), .ZN(
        n10383) );
  AND4_X1 U11559 ( .A1(n10376), .A2(n10375), .A3(n10374), .A4(n10373), .ZN(
        n10382) );
  INV_X1 U11560 ( .A(n13219), .ZN(n17216) );
  AND2_X2 U11561 ( .A1(n12954), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11723) );
  INV_X2 U11562 ( .A(n16547), .ZN(U215) );
  AND4_X1 U11563 ( .A1(n10315), .A2(n10314), .A3(n10313), .A4(n10312), .ZN(
        n10316) );
  AND4_X1 U11564 ( .A1(n11431), .A2(n11430), .A3(n11429), .A4(n11428), .ZN(
        n11432) );
  AND2_X2 U11565 ( .A1(n12944), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12782) );
  NAND2_X1 U11566 ( .A1(n11652), .A2(n11651), .ZN(n10264) );
  INV_X1 U11567 ( .A(n13063), .ZN(n13219) );
  BUF_X2 U11568 ( .A(n10335), .Z(n11059) );
  BUF_X2 U11569 ( .A(n10387), .Z(n11085) );
  NAND2_X2 U11570 ( .A1(n19940), .A2(n19830), .ZN(n19875) );
  INV_X1 U11572 ( .A(n13047), .ZN(n13161) );
  NOR2_X1 U11573 ( .A1(n18236), .A2(n17909), .ZN(n18881) );
  INV_X1 U11574 ( .A(n13011), .ZN(n17136) );
  BUF_X4 U11575 ( .A(n12797), .Z(n12954) );
  AND2_X2 U11576 ( .A1(n12953), .A2(n11651), .ZN(n12783) );
  NOR3_X2 U11577 ( .A1(n18745), .A2(n18718), .A3(n18366), .ZN(n18337) );
  BUF_X4 U11578 ( .A(n12949), .Z(n12944) );
  INV_X2 U11579 ( .A(n12801), .ZN(n11652) );
  BUF_X4 U11580 ( .A(n13077), .Z(n9837) );
  OR2_X1 U11581 ( .A1(n13009), .A2(n16947), .ZN(n14437) );
  BUF_X4 U11582 ( .A(n13027), .Z(n9838) );
  CLKBUF_X1 U11583 ( .A(n12828), .Z(n12950) );
  BUF_X2 U11584 ( .A(n11646), .Z(n12953) );
  AND2_X2 U11585 ( .A1(n10284), .A2(n10293), .ZN(n10595) );
  CLKBUF_X3 U11586 ( .A(n11078), .Z(n10930) );
  BUF_X2 U11587 ( .A(n10330), .Z(n11058) );
  INV_X2 U11588 ( .A(n16552), .ZN(n9840) );
  NAND2_X2 U11590 ( .A1(n20802), .A2(n20208), .ZN(n10609) );
  AND2_X2 U11591 ( .A1(n11654), .A2(n15754), .ZN(n12828) );
  NAND2_X1 U11592 ( .A1(n18844), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13014) );
  NAND2_X1 U11593 ( .A1(n18862), .A2(n18870), .ZN(n16947) );
  NAND2_X1 U11594 ( .A1(n18844), .A2(n18854), .ZN(n13009) );
  NAND3_X2 U11595 ( .A1(n18902), .A2(n18891), .A3(n18901), .ZN(n18218) );
  INV_X2 U11596 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10581) );
  NAND2_X1 U11597 ( .A1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n11329) );
  INV_X2 U11598 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n9947) );
  INV_X1 U11599 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n18844) );
  INV_X1 U11600 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n15737) );
  INV_X1 U11601 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n18862) );
  INV_X2 U11602 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n18854) );
  NAND2_X1 U11603 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n18705) );
  AND3_X1 U11604 ( .A1(n11442), .A2(n12426), .A3(n12392), .ZN(n12443) );
  AND2_X1 U11605 ( .A1(n10284), .A2(n10290), .ZN(n9864) );
  AND2_X1 U11606 ( .A1(n10284), .A2(n13743), .ZN(n9841) );
  AND2_X1 U11607 ( .A1(n10284), .A2(n13743), .ZN(n9842) );
  BUF_X4 U11608 ( .A(n16913), .Z(n9843) );
  XOR2_X1 U11609 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .B(n13315), .Z(
        n16913) );
  AND2_X1 U11610 ( .A1(n10284), .A2(n13743), .ZN(n10980) );
  AND2_X1 U11611 ( .A1(n15743), .A2(n15754), .ZN(n9844) );
  AND2_X1 U11612 ( .A1(n15743), .A2(n15754), .ZN(n9845) );
  AND2_X1 U11613 ( .A1(n9854), .A2(n10421), .ZN(n9846) );
  INV_X1 U11614 ( .A(n10433), .ZN(n10452) );
  AND2_X1 U11615 ( .A1(n11653), .A2(n15752), .ZN(n9847) );
  AND2_X1 U11616 ( .A1(n11653), .A2(n15752), .ZN(n9848) );
  NOR2_X4 U11617 ( .A1(n11443), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n11792) );
  AND2_X2 U11618 ( .A1(n20177), .A2(n9854), .ZN(n11180) );
  NOR2_X2 U11619 ( .A1(n13487), .A2(n20194), .ZN(n13371) );
  AND2_X1 U11620 ( .A1(n12290), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n9850) );
  AND3_X4 U11621 ( .A1(n15754), .A2(n10246), .A3(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11427) );
  INV_X2 U11622 ( .A(n9887), .ZN(n9851) );
  OR2_X1 U11623 ( .A1(n13016), .A2(n18705), .ZN(n9887) );
  AND2_X1 U11624 ( .A1(n11654), .A2(n15754), .ZN(n9852) );
  AND2_X1 U11625 ( .A1(n11654), .A2(n15754), .ZN(n9853) );
  AND2_X1 U11626 ( .A1(n12007), .A2(n12673), .ZN(n12008) );
  AND2_X1 U11627 ( .A1(n12007), .A2(n13584), .ZN(n11988) );
  NAND2_X1 U11628 ( .A1(n12350), .A2(n12417), .ZN(n12168) );
  AND2_X1 U11629 ( .A1(n11653), .A2(n15752), .ZN(n9855) );
  NOR2_X1 U11630 ( .A1(n12672), .A2(n19098), .ZN(n12007) );
  AND3_X1 U11631 ( .A1(n12672), .A2(n10161), .A3(n12673), .ZN(n12020) );
  OAI211_X2 U11632 ( .C1(n11978), .C2(n11977), .A(n11976), .B(n11975), .ZN(
        n12672) );
  NAND2_X2 U11633 ( .A1(n11162), .A2(n20168), .ZN(n12536) );
  AND2_X2 U11634 ( .A1(n10428), .A2(n10411), .ZN(n11162) );
  INV_X1 U11635 ( .A(n11400), .ZN(n9856) );
  INV_X1 U11636 ( .A(n11400), .ZN(n9857) );
  NAND2_X2 U11637 ( .A1(n15758), .A2(n15737), .ZN(n11400) );
  NOR2_X4 U11638 ( .A1(n14199), .A2(n10281), .ZN(n14254) );
  NAND2_X2 U11639 ( .A1(n14071), .A2(n10705), .ZN(n14199) );
  OAI21_X2 U11640 ( .B1(n14891), .B2(n10273), .A(n12646), .ZN(n16049) );
  NOR2_X4 U11641 ( .A1(n14567), .A2(n14568), .ZN(n12655) );
  NAND4_X1 U11642 ( .A1(n10408), .A2(n10407), .A3(n10406), .A4(n10405), .ZN(
        n9859) );
  NAND2_X2 U11643 ( .A1(n14367), .A2(n10803), .ZN(n14721) );
  AND2_X2 U11644 ( .A1(n14254), .A2(n10203), .ZN(n14367) );
  NOR2_X2 U11645 ( .A1(n14606), .A2(n14705), .ZN(n14694) );
  NAND2_X2 U11646 ( .A1(n10578), .A2(n10537), .ZN(n13917) );
  XNOR2_X1 U11647 ( .A(n10434), .B(n10452), .ZN(n20264) );
  NAND2_X2 U11648 ( .A1(n10141), .A2(n10140), .ZN(n14934) );
  NAND3_X2 U11649 ( .A1(n10433), .A2(n10431), .A3(n10430), .ZN(n10454) );
  AND2_X1 U11650 ( .A1(n10284), .A2(n10293), .ZN(n9861) );
  AND2_X2 U11651 ( .A1(n10284), .A2(n10293), .ZN(n9862) );
  NOR2_X2 U11652 ( .A1(n14691), .A2(n14692), .ZN(n14680) );
  AND2_X1 U11653 ( .A1(n10284), .A2(n10290), .ZN(n9865) );
  AND2_X1 U11654 ( .A1(n10284), .A2(n10290), .ZN(n10510) );
  XNOR2_X1 U11655 ( .A(n10544), .B(n10543), .ZN(n13911) );
  AND2_X1 U11656 ( .A1(n13743), .A2(n10292), .ZN(n10498) );
  XNOR2_X2 U11657 ( .A(n13758), .B(n20292), .ZN(n10003) );
  XNOR2_X2 U11658 ( .A(n10497), .B(n10496), .ZN(n10551) );
  CLKBUF_X1 U11659 ( .A(n19083), .Z(n9868) );
  NOR4_X1 U11660 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(P2_STATEBS16_REG_SCAN_IN), .A4(n19802), .ZN(n19083) );
  NAND2_X1 U11661 ( .A1(n20182), .A2(n12633), .ZN(n10523) );
  AND2_X1 U11662 ( .A1(n9854), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11106) );
  OAI211_X1 U11663 ( .C1(n11106), .C2(n10525), .A(n10524), .B(n10523), .ZN(
        n10549) );
  INV_X1 U11664 ( .A(n14210), .ZN(n10107) );
  NAND2_X1 U11665 ( .A1(n13123), .A2(n13299), .ZN(n13126) );
  NAND2_X1 U11666 ( .A1(n10155), .A2(n12432), .ZN(n10154) );
  AND2_X1 U11667 ( .A1(n11788), .A2(n19290), .ZN(n11442) );
  NAND2_X2 U11668 ( .A1(n11442), .A2(n12432), .ZN(n11456) );
  OAI22_X1 U11669 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18727), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n13170), .ZN(n13176) );
  AOI21_X1 U11670 ( .B1(n18718), .B2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n13168), .ZN(n13174) );
  OAI22_X1 U11671 ( .A1(n18854), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B1(
        n18723), .B2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13173) );
  NAND2_X1 U11672 ( .A1(n14674), .A2(n9928), .ZN(n14567) );
  NAND2_X1 U11673 ( .A1(n20190), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n10801) );
  INV_X1 U11674 ( .A(n20093), .ZN(n10131) );
  OR2_X1 U11675 ( .A1(n13808), .A2(n11197), .ZN(n11243) );
  NAND2_X1 U11676 ( .A1(n10449), .A2(n10448), .ZN(n10495) );
  INV_X1 U11677 ( .A(n10439), .ZN(n10449) );
  AND3_X1 U11678 ( .A1(n10530), .A2(n10529), .A3(n10528), .ZN(n10531) );
  AOI21_X1 U11679 ( .B1(n10191), .B2(n10521), .A(n12631), .ZN(n10189) );
  NOR2_X1 U11680 ( .A1(n10476), .A2(n9869), .ZN(n10023) );
  NOR2_X1 U11681 ( .A1(n19286), .A2(n10078), .ZN(n10077) );
  NAND2_X1 U11682 ( .A1(n11662), .A2(n10267), .ZN(n12119) );
  INV_X1 U11683 ( .A(n12358), .ZN(n12165) );
  NAND2_X1 U11684 ( .A1(n11981), .A2(n11982), .ZN(n10101) );
  INV_X1 U11685 ( .A(n13360), .ZN(n10120) );
  INV_X1 U11686 ( .A(n11610), .ZN(n11602) );
  INV_X1 U11687 ( .A(n12363), .ZN(n12366) );
  OAI21_X2 U11688 ( .B1(n9992), .B2(n15712), .A(n9987), .ZN(n15674) );
  NAND2_X1 U11689 ( .A1(n9988), .A2(n9903), .ZN(n9987) );
  AND4_X1 U11690 ( .A1(n11737), .A2(n11736), .A3(n11735), .A4(n11734), .ZN(
        n11744) );
  OR2_X1 U11691 ( .A1(n11712), .A2(n11711), .ZN(n12096) );
  CLKBUF_X1 U11692 ( .A(n11543), .Z(n11606) );
  AND2_X1 U11694 ( .A1(n12897), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n12679) );
  INV_X1 U11695 ( .A(n11412), .ZN(n9979) );
  NOR3_X1 U11696 ( .A1(n13273), .A2(n15830), .A3(n13274), .ZN(n13257) );
  NOR2_X1 U11697 ( .A1(n13009), .A2(n13010), .ZN(n13027) );
  NAND2_X1 U11698 ( .A1(n10139), .A2(n12573), .ZN(n13383) );
  AND2_X1 U11699 ( .A1(n9912), .A2(n12637), .ZN(n10140) );
  INV_X1 U11700 ( .A(n14352), .ZN(n10106) );
  AND2_X1 U11701 ( .A1(n13839), .A2(n12696), .ZN(n12697) );
  AND2_X1 U11702 ( .A1(n9996), .A2(n9995), .ZN(n9994) );
  INV_X1 U11703 ( .A(n16288), .ZN(n9995) );
  XNOR2_X1 U11704 ( .A(n12678), .B(n12679), .ZN(n13582) );
  XNOR2_X1 U11705 ( .A(n13835), .B(n13623), .ZN(n13624) );
  NAND2_X1 U11706 ( .A1(n17818), .A2(n18043), .ZN(n13136) );
  INV_X1 U11707 ( .A(n18262), .ZN(n15830) );
  NAND2_X1 U11708 ( .A1(n14550), .A2(n14548), .ZN(n20808) );
  OR2_X1 U11709 ( .A1(n10573), .A2(n10572), .ZN(n12603) );
  NAND2_X1 U11710 ( .A1(n9886), .A2(n15351), .ZN(n10233) );
  NAND2_X1 U11711 ( .A1(n11448), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11491) );
  AND2_X1 U11712 ( .A1(n10214), .A2(n11765), .ZN(n11470) );
  NOR2_X1 U11713 ( .A1(n14035), .A2(n10215), .ZN(n10214) );
  NAND2_X1 U11714 ( .A1(n12380), .A2(n16370), .ZN(n10215) );
  INV_X1 U11715 ( .A(n11437), .ZN(n11438) );
  NOR2_X1 U11716 ( .A1(n14035), .A2(n19275), .ZN(n12431) );
  INV_X1 U11717 ( .A(n11371), .ZN(n11372) );
  AND2_X1 U11718 ( .A1(n13284), .A2(n13114), .ZN(n13116) );
  NOR2_X1 U11719 ( .A1(n9916), .A2(n10195), .ZN(n10194) );
  INV_X1 U11720 ( .A(n14608), .ZN(n10195) );
  INV_X1 U11721 ( .A(n11099), .ZN(n11074) );
  NAND2_X1 U11722 ( .A1(n15072), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11099) );
  AND2_X1 U11723 ( .A1(n10205), .A2(n10204), .ZN(n10203) );
  INV_X1 U11724 ( .A(n14369), .ZN(n10204) );
  AND2_X1 U11725 ( .A1(n10632), .A2(n10666), .ZN(n12601) );
  NOR2_X1 U11726 ( .A1(n14519), .A2(n20802), .ZN(n10552) );
  AND2_X1 U11727 ( .A1(n10136), .A2(n12630), .ZN(n10133) );
  AND3_X1 U11728 ( .A1(n14907), .A2(n14892), .A3(n12645), .ZN(n12646) );
  NAND2_X1 U11729 ( .A1(n10146), .A2(n16050), .ZN(n10145) );
  INV_X1 U11730 ( .A(n12646), .ZN(n10146) );
  NAND2_X1 U11731 ( .A1(n10004), .A2(n12641), .ZN(n14893) );
  NAND2_X1 U11732 ( .A1(n14906), .A2(n14892), .ZN(n10004) );
  NOR2_X1 U11733 ( .A1(n14740), .A2(n14739), .ZN(n14641) );
  NAND2_X1 U11734 ( .A1(n10037), .A2(n14160), .ZN(n10036) );
  INV_X1 U11735 ( .A(n14161), .ZN(n10037) );
  INV_X1 U11736 ( .A(n16090), .ZN(n10033) );
  NAND2_X1 U11737 ( .A1(n20264), .A2(n10477), .ZN(n9997) );
  NAND2_X1 U11738 ( .A1(n10479), .A2(n10478), .ZN(n20205) );
  INV_X1 U11739 ( .A(n20198), .ZN(n20297) );
  OR2_X1 U11740 ( .A1(n9854), .A2(n20806), .ZN(n10562) );
  NAND2_X1 U11741 ( .A1(n20182), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10563) );
  AOI21_X1 U11742 ( .B1(n11142), .B2(n11141), .A(n11140), .ZN(n11154) );
  NAND2_X1 U11743 ( .A1(n11626), .A2(n11625), .ZN(n12314) );
  NOR2_X1 U11744 ( .A1(n11459), .A2(n11441), .ZN(n10253) );
  AND2_X1 U11745 ( .A1(n11633), .A2(n11701), .ZN(n12313) );
  INV_X1 U11746 ( .A(n12314), .ZN(n12318) );
  NOR2_X1 U11747 ( .A1(n11799), .A2(n11798), .ZN(n11805) );
  OR2_X1 U11748 ( .A1(n11494), .A2(n15754), .ZN(n11486) );
  NOR2_X1 U11749 ( .A1(n15752), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12799) );
  NOR2_X1 U11750 ( .A1(n13336), .A2(n13337), .ZN(n10187) );
  NAND2_X1 U11751 ( .A1(n14138), .A2(n10174), .ZN(n12817) );
  AND2_X1 U11752 ( .A1(n9920), .A2(n12780), .ZN(n10174) );
  AND2_X1 U11753 ( .A1(n14035), .A2(n19297), .ZN(n10153) );
  NOR2_X1 U11754 ( .A1(n12486), .A2(n10110), .ZN(n10109) );
  INV_X1 U11755 ( .A(n12297), .ZN(n10110) );
  INV_X1 U11756 ( .A(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n10042) );
  NAND2_X1 U11757 ( .A1(n10117), .A2(n13927), .ZN(n10116) );
  INV_X1 U11758 ( .A(n13888), .ZN(n10117) );
  AND2_X1 U11759 ( .A1(n11514), .A2(n11521), .ZN(n10104) );
  INV_X1 U11760 ( .A(n12408), .ZN(n9965) );
  INV_X1 U11761 ( .A(n15200), .ZN(n10121) );
  NOR2_X1 U11762 ( .A1(n13348), .A2(n12417), .ZN(n12236) );
  INV_X1 U11763 ( .A(n15847), .ZN(n10182) );
  INV_X1 U11764 ( .A(n11613), .ZN(n11608) );
  NOR2_X1 U11765 ( .A1(n10116), .A2(n10115), .ZN(n10114) );
  NOR2_X1 U11766 ( .A1(n11722), .A2(n11721), .ZN(n12162) );
  NAND2_X1 U11767 ( .A1(n12341), .A2(n12101), .ZN(n9961) );
  NOR2_X1 U11768 ( .A1(n11806), .A2(n10181), .ZN(n10180) );
  INV_X1 U11769 ( .A(n14003), .ZN(n10181) );
  NOR2_X1 U11770 ( .A1(n11508), .A2(n14095), .ZN(n11501) );
  INV_X1 U11771 ( .A(n13828), .ZN(n11514) );
  INV_X1 U11772 ( .A(n13829), .ZN(n11515) );
  NAND2_X1 U11773 ( .A1(n12061), .A2(n12060), .ZN(n12105) );
  NAND2_X1 U11774 ( .A1(n12059), .A2(n12058), .ZN(n12060) );
  OAI211_X1 U11775 ( .C1(n11508), .C2(n11481), .A(n11480), .B(n11494), .ZN(
        n11979) );
  NOR2_X1 U11776 ( .A1(n10271), .A2(n11479), .ZN(n11480) );
  OAI21_X1 U11777 ( .B1(n11543), .B2(n12115), .A(n11478), .ZN(n11479) );
  OAI21_X1 U11778 ( .B1(n12672), .B2(n12683), .A(n12671), .ZN(n12693) );
  NOR2_X1 U11779 ( .A1(n11441), .A2(n11418), .ZN(n11421) );
  AND2_X1 U11780 ( .A1(n12672), .A2(n10161), .ZN(n10087) );
  NOR2_X1 U11781 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18870), .ZN(
        n13267) );
  OR3_X1 U11782 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18844), .A3(
        n18700), .ZN(n17215) );
  OAI21_X1 U11783 ( .B1(n15815), .B2(n15816), .A(n15804), .ZN(n16584) );
  NAND2_X1 U11784 ( .A1(n18862), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13015) );
  NAND2_X1 U11785 ( .A1(n10224), .A2(n10223), .ZN(n10222) );
  NOR2_X1 U11786 ( .A1(n10225), .A2(n20983), .ZN(n10223) );
  INV_X1 U11787 ( .A(n17687), .ZN(n10224) );
  NAND2_X1 U11788 ( .A1(n17835), .A2(n13125), .ZN(n13128) );
  OAI22_X1 U11789 ( .A1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n18691), .B1(
        n13177), .B2(n13176), .ZN(n13269) );
  AND2_X1 U11790 ( .A1(n13175), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n13177) );
  AOI21_X1 U11791 ( .B1(n13174), .B2(n13173), .A(n13172), .ZN(n13272) );
  OR2_X1 U11792 ( .A1(n13016), .A2(n13015), .ZN(n10259) );
  AND2_X1 U11793 ( .A1(n18694), .A2(n13277), .ZN(n14391) );
  AOI211_X1 U11794 ( .C1(n17200), .C2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A(
        n13225), .B(n13224), .ZN(n13226) );
  AOI211_X1 U11795 ( .C1(n17098), .C2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A(
        n13246), .B(n13245), .ZN(n13247) );
  NAND2_X1 U11796 ( .A1(n20022), .A2(n11269), .ZN(n11282) );
  NOR2_X1 U11797 ( .A1(n14558), .A2(n10208), .ZN(n10207) );
  INV_X1 U11798 ( .A(n12656), .ZN(n10208) );
  NAND2_X1 U11799 ( .A1(n11077), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n11172) );
  INV_X1 U11800 ( .A(n11054), .ZN(n11077) );
  INV_X1 U11801 ( .A(n10634), .ZN(n10635) );
  INV_X1 U11802 ( .A(n13886), .ZN(n10614) );
  NAND2_X1 U11803 ( .A1(n10608), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10634) );
  OAI21_X1 U11804 ( .B1(n13917), .B2(n10801), .A(n10269), .ZN(n10541) );
  NAND2_X1 U11805 ( .A1(n10548), .A2(n10547), .ZN(n10188) );
  INV_X1 U11806 ( .A(n15015), .ZN(n10008) );
  NAND2_X1 U11807 ( .A1(n12650), .A2(n15015), .ZN(n14869) );
  NAND2_X1 U11808 ( .A1(n14641), .A2(n11220), .ZN(n14642) );
  INV_X1 U11809 ( .A(n14644), .ZN(n11220) );
  NAND2_X1 U11810 ( .A1(n9957), .A2(n9956), .ZN(n14740) );
  NOR2_X1 U11811 ( .A1(n14256), .A2(n14308), .ZN(n9956) );
  NAND2_X1 U11812 ( .A1(n14246), .A2(n12636), .ZN(n10141) );
  NOR2_X1 U11813 ( .A1(n13944), .A2(n13943), .ZN(n11196) );
  INV_X1 U11814 ( .A(n13945), .ZN(n9955) );
  NAND2_X1 U11815 ( .A1(n20094), .A2(n10127), .ZN(n10126) );
  INV_X1 U11816 ( .A(n10129), .ZN(n10128) );
  AOI21_X1 U11817 ( .B1(n12600), .B2(n10131), .A(n10130), .ZN(n10124) );
  INV_X1 U11818 ( .A(n12600), .ZN(n10125) );
  NAND2_X1 U11819 ( .A1(n20094), .A2(n20093), .ZN(n20092) );
  AND2_X1 U11820 ( .A1(n14167), .A2(n14166), .ZN(n15054) );
  OR2_X1 U11821 ( .A1(n10551), .A2(n10138), .ZN(n10134) );
  OR2_X1 U11822 ( .A1(n10521), .A2(n10549), .ZN(n10138) );
  AND2_X1 U11823 ( .A1(n10549), .A2(n20806), .ZN(n10135) );
  NOR2_X1 U11824 ( .A1(n10533), .A2(n10532), .ZN(n10534) );
  NAND2_X1 U11825 ( .A1(n10476), .A2(n9869), .ZN(n10024) );
  INV_X1 U11826 ( .A(n10476), .ZN(n10025) );
  NAND2_X1 U11827 ( .A1(n10027), .A2(n10023), .ZN(n10022) );
  INV_X1 U11828 ( .A(n15901), .ZN(n13723) );
  OR2_X1 U11829 ( .A1(n20263), .A2(n9866), .ZN(n20204) );
  NOR2_X1 U11830 ( .A1(n13917), .A2(n10576), .ZN(n20383) );
  INV_X1 U11831 ( .A(n9866), .ZN(n20496) );
  AND2_X1 U11832 ( .A1(n20297), .A2(n20469), .ZN(n20598) );
  INV_X1 U11833 ( .A(n10421), .ZN(n20168) );
  NAND2_X1 U11834 ( .A1(n10563), .A2(n10562), .ZN(n11155) );
  AND2_X1 U11836 ( .A1(n13782), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n15897) );
  OR2_X1 U11837 ( .A1(n15119), .A2(n10053), .ZN(n10054) );
  NAND2_X1 U11838 ( .A1(n12266), .A2(n12265), .ZN(n16211) );
  INV_X1 U11839 ( .A(n15345), .ZN(n10070) );
  NAND2_X1 U11840 ( .A1(n11752), .A2(n12248), .ZN(n12253) );
  NAND2_X1 U11841 ( .A1(n12250), .A2(n12269), .ZN(n11752) );
  OR2_X1 U11842 ( .A1(n10075), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n10074) );
  OR2_X1 U11843 ( .A1(n10077), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n10075) );
  INV_X1 U11844 ( .A(n12119), .ZN(n10056) );
  NOR2_X1 U11845 ( .A1(n12119), .A2(n12118), .ZN(n12107) );
  INV_X1 U11846 ( .A(n10187), .ZN(n15095) );
  NOR2_X1 U11847 ( .A1(n19290), .A2(n13537), .ZN(n13559) );
  AND2_X1 U11848 ( .A1(n10062), .A2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n10061) );
  AND2_X1 U11849 ( .A1(n9881), .A2(n14323), .ZN(n10105) );
  NAND2_X1 U11850 ( .A1(n12366), .A2(n12102), .ZN(n12365) );
  OR2_X1 U11851 ( .A1(n12361), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n9996) );
  AND2_X1 U11852 ( .A1(n11527), .A2(n11526), .ZN(n13850) );
  AND2_X1 U11853 ( .A1(n13335), .A2(n9940), .ZN(n11615) );
  NAND2_X1 U11854 ( .A1(n12409), .A2(n12408), .ZN(n12495) );
  NOR2_X1 U11855 ( .A1(n15175), .A2(n13333), .ZN(n13335) );
  OR2_X1 U11856 ( .A1(n13332), .A2(n12417), .ZN(n12403) );
  NAND2_X1 U11857 ( .A1(n12402), .A2(n12408), .ZN(n12277) );
  AND2_X1 U11858 ( .A1(n12244), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15385) );
  NAND2_X1 U11859 ( .A1(n15410), .A2(n15368), .ZN(n15382) );
  NAND2_X1 U11860 ( .A1(n15398), .A2(n9984), .ZN(n15615) );
  INV_X1 U11861 ( .A(n15434), .ZN(n9984) );
  NAND2_X1 U11862 ( .A1(n10092), .A2(n15676), .ZN(n10089) );
  NOR2_X1 U11863 ( .A1(n15698), .A2(n15696), .ZN(n10212) );
  NAND2_X1 U11864 ( .A1(n9991), .A2(n9989), .ZN(n9992) );
  NAND2_X1 U11865 ( .A1(n9990), .A2(n12367), .ZN(n9989) );
  INV_X1 U11866 ( .A(n12360), .ZN(n10252) );
  NAND2_X1 U11867 ( .A1(n12357), .A2(n12356), .ZN(n12360) );
  AND2_X1 U11868 ( .A1(n12347), .A2(n14226), .ZN(n14218) );
  AND2_X1 U11869 ( .A1(n12400), .A2(n19808), .ZN(n12459) );
  INV_X1 U11870 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10211) );
  NAND2_X1 U11871 ( .A1(n13580), .A2(n12682), .ZN(n13625) );
  NAND2_X1 U11872 ( .A1(n13622), .A2(n13624), .ZN(n13837) );
  OR2_X1 U11873 ( .A1(n12693), .A2(n12692), .ZN(n13838) );
  NAND2_X1 U11874 ( .A1(n12690), .A2(n12689), .ZN(n13835) );
  OR2_X1 U11875 ( .A1(n12684), .A2(n12683), .ZN(n12690) );
  NAND2_X1 U11876 ( .A1(n19539), .A2(n14119), .ZN(n19447) );
  NAND2_X1 U11877 ( .A1(n19901), .A2(n14023), .ZN(n19889) );
  OR2_X1 U11878 ( .A1(n19539), .A2(n14119), .ZN(n19659) );
  OR2_X1 U11879 ( .A1(n19901), .A2(n19910), .ZN(n19688) );
  AOI21_X2 U11880 ( .B1(n13537), .B2(n16397), .A(n12321), .ZN(n19389) );
  AND2_X1 U11881 ( .A1(n16365), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n16397) );
  INV_X1 U11882 ( .A(n13106), .ZN(n10218) );
  INV_X1 U11883 ( .A(n17898), .ZN(n17908) );
  AND2_X1 U11884 ( .A1(n15906), .A2(n10274), .ZN(n13155) );
  NAND2_X1 U11885 ( .A1(n9890), .A2(n10241), .ZN(n17695) );
  INV_X1 U11886 ( .A(n10243), .ZN(n10242) );
  AOI21_X1 U11887 ( .B1(n18024), .B2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n10243) );
  INV_X1 U11888 ( .A(n18024), .ZN(n10239) );
  INV_X1 U11889 ( .A(n17754), .ZN(n10240) );
  INV_X1 U11890 ( .A(n18886), .ZN(n16589) );
  AND2_X1 U11891 ( .A1(n17898), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n17907) );
  NAND2_X1 U11892 ( .A1(n17907), .A2(n17901), .ZN(n17900) );
  NOR2_X1 U11893 ( .A1(n13238), .A2(n13237), .ZN(n18262) );
  NOR2_X1 U11894 ( .A1(n14504), .A2(n13782), .ZN(n11174) );
  AND2_X1 U11895 ( .A1(n20022), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20026) );
  AND2_X1 U11896 ( .A1(n14504), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13965) );
  INV_X1 U11897 ( .A(n14613), .ZN(n16020) );
  OR2_X1 U11898 ( .A1(n20098), .A2(n12661), .ZN(n14900) );
  INV_X1 U11899 ( .A(n20145), .ZN(n20114) );
  CLKBUF_X1 U11900 ( .A(n13910), .Z(n20529) );
  INV_X1 U11901 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20783) );
  OAI21_X1 U11902 ( .B1(n13909), .B2(n13908), .A(n20198), .ZN(n20791) );
  NOR2_X1 U11903 ( .A1(n18958), .A2(n11335), .ZN(n18942) );
  NAND2_X2 U11904 ( .A1(n11301), .A2(n11300), .ZN(n19079) );
  NAND2_X1 U11905 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n11300) );
  XNOR2_X1 U11906 ( .A(n12508), .B(n12507), .ZN(n14470) );
  XNOR2_X1 U11907 ( .A(n12521), .B(n11962), .ZN(n12453) );
  XNOR2_X1 U11908 ( .A(n12373), .B(n20998), .ZN(n12995) );
  NOR2_X1 U11909 ( .A1(n10257), .A2(n12528), .ZN(n10256) );
  XNOR2_X1 U11910 ( .A(n9968), .B(n9891), .ZN(n12988) );
  OAI21_X1 U11911 ( .B1(n12409), .B2(n9966), .A(n9962), .ZN(n9968) );
  NAND2_X1 U11912 ( .A1(n12453), .A2(n16344), .ZN(n10176) );
  NOR2_X1 U11913 ( .A1(n12452), .A2(n12480), .ZN(n10177) );
  NOR2_X1 U11914 ( .A1(n12479), .A2(n20998), .ZN(n12480) );
  OR2_X1 U11915 ( .A1(n12451), .A2(n12989), .ZN(n12452) );
  OR2_X1 U11916 ( .A1(n12454), .A2(n16326), .ZN(n10178) );
  AND2_X1 U11917 ( .A1(n12459), .A2(n19929), .ZN(n16338) );
  INV_X1 U11918 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19898) );
  NOR2_X1 U11919 ( .A1(n19476), .A2(n19889), .ZN(n19410) );
  NOR2_X1 U11920 ( .A1(n18747), .A2(n18901), .ZN(n18884) );
  NOR2_X1 U11921 ( .A1(n17291), .A2(n17434), .ZN(n17286) );
  NOR2_X1 U11922 ( .A1(n17540), .A2(n17357), .ZN(n17352) );
  NOR2_X1 U11923 ( .A1(n13304), .A2(n17913), .ZN(n17598) );
  NOR2_X1 U11924 ( .A1(n18236), .A2(n17905), .ZN(n17767) );
  NAND2_X1 U11925 ( .A1(n14393), .A2(n13314), .ZN(n17913) );
  INV_X1 U11926 ( .A(n17894), .ZN(n17914) );
  NOR2_X1 U11927 ( .A1(n18231), .A2(n18227), .ZN(n18220) );
  INV_X1 U11928 ( .A(n10444), .ZN(n10420) );
  AOI21_X1 U11929 ( .B1(n11155), .B2(n9858), .A(n11113), .ZN(n11115) );
  AOI22_X1 U11930 ( .A1(n11427), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n9857), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11409) );
  NAND2_X1 U11931 ( .A1(n11768), .A2(n11767), .ZN(n11769) );
  NAND2_X1 U11932 ( .A1(n12782), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n11767) );
  OAI21_X1 U11933 ( .B1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n18854), .A(
        n13169), .ZN(n13170) );
  OR2_X1 U11934 ( .A1(n13173), .A2(n13174), .ZN(n13169) );
  CLKBUF_X2 U11935 ( .A(n10596), .Z(n10481) );
  AND2_X1 U11936 ( .A1(n10626), .A2(n10625), .ZN(n10629) );
  XNOR2_X1 U11937 ( .A(n12612), .B(n10670), .ZN(n12621) );
  OR2_X1 U11938 ( .A1(n10652), .A2(n10651), .ZN(n12622) );
  NAND2_X1 U11939 ( .A1(n10522), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10192) );
  INV_X1 U11940 ( .A(n10562), .ZN(n10527) );
  NAND2_X1 U11941 ( .A1(n11646), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n11402) );
  INV_X1 U11942 ( .A(n11456), .ZN(n10151) );
  AOI21_X1 U11943 ( .B1(n14130), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A(
        n12006), .ZN(n12011) );
  NOR2_X1 U11944 ( .A1(n12684), .A2(n11990), .ZN(n12019) );
  AOI22_X1 U11945 ( .A1(n11427), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n9856), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11354) );
  NOR2_X1 U11946 ( .A1(n19290), .A2(n11451), .ZN(n11437) );
  NAND2_X1 U11947 ( .A1(n18870), .A2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13010) );
  NOR2_X1 U11948 ( .A1(n17401), .A2(n13096), .ZN(n13123) );
  NAND2_X1 U11949 ( .A1(n9958), .A2(n21089), .ZN(n11255) );
  NAND2_X1 U11950 ( .A1(n10467), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n10375) );
  AND2_X1 U11951 ( .A1(n10200), .A2(n10201), .ZN(n10199) );
  INV_X1 U11952 ( .A(n14595), .ZN(n10200) );
  AND2_X1 U11953 ( .A1(n10202), .A2(n14675), .ZN(n10201) );
  INV_X1 U11954 ( .A(n14668), .ZN(n10202) );
  INV_X1 U11955 ( .A(n10197), .ZN(n10196) );
  NOR2_X1 U11956 ( .A1(n10198), .A2(n14722), .ZN(n10197) );
  INV_X1 U11957 ( .A(n14626), .ZN(n10198) );
  AND2_X1 U11958 ( .A1(n10770), .A2(n10206), .ZN(n10205) );
  AND2_X1 U11959 ( .A1(n14640), .A2(n14743), .ZN(n10770) );
  INV_X1 U11960 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n21024) );
  INV_X1 U11961 ( .A(n11105), .ZN(n10414) );
  AND2_X1 U11962 ( .A1(n12562), .A2(n13400), .ZN(n13369) );
  OR2_X1 U11963 ( .A1(n14713), .A2(n14712), .ZN(n9951) );
  AND2_X1 U11964 ( .A1(n14911), .A2(n12640), .ZN(n14892) );
  NAND2_X1 U11965 ( .A1(n16064), .A2(n12639), .ZN(n14906) );
  AND2_X1 U11966 ( .A1(n14923), .A2(n14921), .ZN(n14907) );
  OAI21_X1 U11967 ( .B1(n12600), .B2(n10130), .A(n12611), .ZN(n10129) );
  OR2_X1 U11968 ( .A1(n10603), .A2(n10602), .ZN(n12602) );
  NAND2_X1 U11969 ( .A1(n20126), .A2(n12583), .ZN(n12591) );
  NAND2_X1 U11970 ( .A1(n9901), .A2(n20182), .ZN(n13409) );
  NAND2_X1 U11971 ( .A1(n9958), .A2(n11250), .ZN(n11175) );
  OR2_X1 U11972 ( .A1(n10491), .A2(n10490), .ZN(n12564) );
  INV_X1 U11973 ( .A(n10563), .ZN(n10026) );
  AOI21_X1 U11974 ( .B1(n10454), .B2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n10432), .ZN(n10434) );
  NOR2_X1 U11975 ( .A1(n15110), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n12263) );
  OR3_X1 U11976 ( .A1(n11632), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A3(
        n15918), .ZN(n11701) );
  AND2_X1 U11977 ( .A1(n11443), .A2(n19917), .ZN(n11789) );
  CLKBUF_X1 U11978 ( .A(n12945), .Z(n12955) );
  NAND2_X1 U11979 ( .A1(n9936), .A2(n15189), .ZN(n10171) );
  INV_X1 U11980 ( .A(n14350), .ZN(n10175) );
  AND2_X1 U11981 ( .A1(n9924), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n10062) );
  INV_X1 U11982 ( .A(n14142), .ZN(n11557) );
  INV_X1 U11983 ( .A(n12507), .ZN(n10108) );
  INV_X1 U11984 ( .A(n10233), .ZN(n10228) );
  NAND2_X1 U11985 ( .A1(n10232), .A2(n9886), .ZN(n10231) );
  INV_X1 U11986 ( .A(n15341), .ZN(n10232) );
  AND2_X1 U11987 ( .A1(n12368), .A2(n12455), .ZN(n10254) );
  INV_X1 U11988 ( .A(n11606), .ZN(n11609) );
  NAND2_X1 U11989 ( .A1(n10093), .A2(n10091), .ZN(n10090) );
  NAND2_X1 U11990 ( .A1(n10212), .A2(n15676), .ZN(n10091) );
  INV_X1 U11991 ( .A(n9994), .ZN(n9990) );
  INV_X1 U11992 ( .A(n15725), .ZN(n10183) );
  NOR2_X1 U11993 ( .A1(n10249), .A2(n12355), .ZN(n10248) );
  INV_X1 U11994 ( .A(n12350), .ZN(n12355) );
  NAND2_X1 U11995 ( .A1(n12164), .A2(n12163), .ZN(n12358) );
  NAND2_X1 U11996 ( .A1(n11451), .A2(n11789), .ZN(n11934) );
  NAND2_X1 U11997 ( .A1(n12379), .A2(n19297), .ZN(n10157) );
  CLKBUF_X1 U11998 ( .A(n12290), .Z(n12291) );
  INV_X1 U11999 ( .A(n12013), .ZN(n12012) );
  NOR2_X1 U12000 ( .A1(n12684), .A2(n12013), .ZN(n12014) );
  AND2_X1 U12001 ( .A1(n19098), .A2(n11989), .ZN(n11998) );
  OAI21_X1 U12002 ( .B1(n11343), .B2(n11342), .A(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11350) );
  NAND2_X1 U12003 ( .A1(n11348), .A2(n11651), .ZN(n11349) );
  NAND2_X1 U12004 ( .A1(n11367), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11375) );
  OAI21_X1 U12005 ( .B1(n11373), .B2(n11372), .A(n11651), .ZN(n11374) );
  NOR2_X1 U12006 ( .A1(n18705), .A2(n13014), .ZN(n13077) );
  NOR2_X1 U12007 ( .A1(n13016), .A2(n16947), .ZN(n13066) );
  INV_X1 U12008 ( .A(n13013), .ZN(n13240) );
  NOR2_X1 U12009 ( .A1(n18705), .A2(n13012), .ZN(n13088) );
  NAND2_X1 U12010 ( .A1(n17098), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n13067) );
  OR2_X1 U12011 ( .A1(n18705), .A2(n13009), .ZN(n9888) );
  INV_X1 U12012 ( .A(n16436), .ZN(n10238) );
  NAND2_X1 U12013 ( .A1(n17859), .A2(n13118), .ZN(n13121) );
  NAND2_X1 U12014 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13016) );
  NOR4_X1 U12015 ( .A1(n13262), .A2(n15830), .A3(n13253), .A4(n13256), .ZN(
        n13263) );
  AOI21_X1 U12016 ( .B1(n13262), .B2(n13261), .A(n15806), .ZN(n13266) );
  NAND2_X1 U12017 ( .A1(n10787), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n10818) );
  OR2_X1 U12018 ( .A1(n10690), .A2(n14080), .ZN(n10706) );
  NOR2_X2 U12019 ( .A1(n9951), .A2(n9950), .ZN(n14703) );
  INV_X1 U12020 ( .A(n14617), .ZN(n9950) );
  AOI21_X1 U12021 ( .B1(n11096), .B2(n14513), .A(n11076), .ZN(n12656) );
  NAND2_X1 U12022 ( .A1(n12655), .A2(n12656), .ZN(n14557) );
  OR2_X1 U12023 ( .A1(n11035), .A2(n14569), .ZN(n11054) );
  AOI21_X1 U12024 ( .B1(n11096), .B2(n14845), .A(n11033), .ZN(n14582) );
  NOR2_X1 U12025 ( .A1(n11011), .A2(n11010), .ZN(n11015) );
  NAND2_X1 U12026 ( .A1(n10970), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n11011) );
  AND2_X1 U12027 ( .A1(n10951), .A2(n10950), .ZN(n14682) );
  AND2_X1 U12028 ( .A1(n10906), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n10907) );
  NOR2_X1 U12029 ( .A1(n10871), .A2(n14616), .ZN(n10872) );
  AND2_X1 U12030 ( .A1(n10872), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n10906) );
  AND2_X1 U12031 ( .A1(n10870), .A2(n10869), .ZN(n14608) );
  CLKBUF_X1 U12032 ( .A(n14606), .Z(n14607) );
  NOR2_X1 U12033 ( .A1(n10837), .A2(n14633), .ZN(n10838) );
  NOR2_X1 U12034 ( .A1(n10818), .A2(n15999), .ZN(n10819) );
  NAND2_X1 U12035 ( .A1(n10819), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n10837) );
  NOR2_X1 U12036 ( .A1(n10771), .A2(n14648), .ZN(n10787) );
  INV_X1 U12037 ( .A(n14367), .ZN(n14730) );
  NAND2_X1 U12038 ( .A1(n10750), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n10771) );
  INV_X1 U12039 ( .A(n10764), .ZN(n10750) );
  OR2_X1 U12040 ( .A1(n14638), .A2(n14637), .ZN(n14639) );
  AND2_X1 U12041 ( .A1(n14744), .A2(n14743), .ZN(n14746) );
  NAND2_X1 U12042 ( .A1(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n10726), .ZN(
        n10764) );
  OR2_X1 U12043 ( .A1(n10706), .A2(n19967), .ZN(n10707) );
  NOR2_X1 U12044 ( .A1(n21019), .A2(n10707), .ZN(n10726) );
  INV_X1 U12045 ( .A(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n21019) );
  CLKBUF_X1 U12046 ( .A(n14254), .Z(n14255) );
  AND3_X1 U12047 ( .A1(n10689), .A2(n10688), .A3(n10687), .ZN(n14073) );
  CLKBUF_X1 U12048 ( .A(n14071), .Z(n14072) );
  NAND2_X1 U12049 ( .A1(n10664), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n10690) );
  INV_X1 U12050 ( .A(n10663), .ZN(n10664) );
  INV_X1 U12051 ( .A(n10655), .ZN(n10656) );
  NAND2_X1 U12052 ( .A1(n10656), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10663) );
  AOI21_X1 U12053 ( .B1(n12601), .B2(n10671), .A(n10640), .ZN(n13942) );
  AOI21_X1 U12054 ( .B1(n12594), .B2(n10671), .A(n10613), .ZN(n13886) );
  NAND2_X1 U12055 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n10582) );
  NOR2_X1 U12056 ( .A1(n21024), .A2(n10582), .ZN(n10608) );
  AND2_X1 U12057 ( .A1(n13369), .A2(n10414), .ZN(n15880) );
  INV_X1 U12058 ( .A(n14475), .ZN(n10000) );
  NOR2_X1 U12059 ( .A1(n14474), .A2(n10123), .ZN(n10122) );
  INV_X1 U12060 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n10123) );
  NOR2_X2 U12061 ( .A1(n14571), .A2(n14510), .ZN(n14552) );
  INV_X1 U12062 ( .A(n14839), .ZN(n10040) );
  INV_X1 U12063 ( .A(n14869), .ZN(n12652) );
  NAND2_X1 U12064 ( .A1(n12651), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14855) );
  NAND2_X1 U12065 ( .A1(n9960), .A2(n9959), .ZN(n14690) );
  INV_X1 U12066 ( .A(n14688), .ZN(n9959) );
  NAND2_X1 U12067 ( .A1(n10149), .A2(n9913), .ZN(n15014) );
  OAI211_X1 U12068 ( .C1(n10144), .C2(n10147), .A(n10143), .B(n12647), .ZN(
        n10149) );
  INV_X1 U12069 ( .A(n10145), .ZN(n10144) );
  INV_X1 U12070 ( .A(n9960), .ZN(n14700) );
  NOR2_X1 U12071 ( .A1(n16049), .A2(n12648), .ZN(n14873) );
  INV_X1 U12072 ( .A(n10147), .ZN(n10142) );
  NAND2_X1 U12073 ( .A1(n14735), .A2(n9948), .ZN(n14713) );
  NOR2_X1 U12074 ( .A1(n14630), .A2(n9949), .ZN(n9948) );
  INV_X1 U12075 ( .A(n14723), .ZN(n9949) );
  NAND2_X1 U12076 ( .A1(n14735), .A2(n14723), .ZN(n14725) );
  AND2_X1 U12077 ( .A1(n15054), .A2(n20121), .ZN(n16115) );
  AND2_X1 U12078 ( .A1(n11224), .A2(n11223), .ZN(n14375) );
  AND3_X1 U12079 ( .A1(n11218), .A2(n11243), .A3(n11217), .ZN(n14739) );
  AND2_X1 U12080 ( .A1(n11215), .A2(n11214), .ZN(n14256) );
  NOR2_X1 U12081 ( .A1(n14257), .A2(n14256), .ZN(n14305) );
  OR2_X1 U12082 ( .A1(n16081), .A2(n12635), .ZN(n14247) );
  INV_X1 U12083 ( .A(n14160), .ZN(n10038) );
  NAND2_X1 U12084 ( .A1(n14076), .A2(n14075), .ZN(n14204) );
  AND3_X1 U12085 ( .A1(n11199), .A2(n11243), .A3(n11198), .ZN(n13996) );
  INV_X1 U12086 ( .A(n13814), .ZN(n9954) );
  INV_X1 U12087 ( .A(n10265), .ZN(n9953) );
  OR2_X1 U12088 ( .A1(n20772), .A2(n12620), .ZN(n12590) );
  OR2_X1 U12089 ( .A1(n14165), .A2(n13726), .ZN(n20121) );
  INV_X1 U12090 ( .A(n13808), .ZN(n13820) );
  OAI21_X1 U12091 ( .B1(n10549), .B2(n9905), .A(n10137), .ZN(n10136) );
  NAND2_X1 U12092 ( .A1(n10549), .A2(n10522), .ZN(n10137) );
  INV_X1 U12093 ( .A(n10495), .ZN(n10496) );
  NAND2_X1 U12094 ( .A1(n13707), .A2(n10002), .ZN(n20234) );
  AND2_X1 U12095 ( .A1(n20383), .A2(n20496), .ZN(n20320) );
  AND2_X1 U12096 ( .A1(n20776), .A2(n20496), .ZN(n20439) );
  INV_X1 U12097 ( .A(n12574), .ZN(n20562) );
  NOR2_X1 U12098 ( .A1(n20569), .A2(n20496), .ZN(n20637) );
  INV_X1 U12099 ( .A(n20266), .ZN(n20638) );
  NAND2_X1 U12100 ( .A1(n12393), .A2(n12320), .ZN(n16365) );
  AND2_X1 U12101 ( .A1(n12314), .A2(n11635), .ZN(n16373) );
  NOR2_X1 U12102 ( .A1(n12280), .A2(n12279), .ZN(n12411) );
  OR2_X1 U12103 ( .A1(n10053), .A2(n15313), .ZN(n10052) );
  OR2_X1 U12104 ( .A1(n15119), .A2(n10053), .ZN(n10051) );
  NAND2_X1 U12106 ( .A1(n12263), .A2(n12262), .ZN(n12273) );
  NAND2_X1 U12107 ( .A1(n12264), .A2(n12272), .ZN(n12280) );
  NOR2_X1 U12108 ( .A1(n12253), .A2(n12252), .ZN(n10048) );
  INV_X1 U12109 ( .A(n10048), .ZN(n12256) );
  OR2_X1 U12110 ( .A1(n13345), .A2(n10053), .ZN(n10071) );
  NAND2_X1 U12111 ( .A1(n12206), .A2(n9929), .ZN(n12250) );
  NAND2_X1 U12112 ( .A1(n12206), .A2(n9880), .ZN(n12234) );
  NAND2_X1 U12113 ( .A1(n12191), .A2(n15144), .ZN(n12194) );
  AND2_X1 U12114 ( .A1(n12107), .A2(n12108), .ZN(n12126) );
  NOR2_X1 U12115 ( .A1(n10053), .A2(n14234), .ZN(n14356) );
  AND2_X1 U12116 ( .A1(n10279), .A2(n13951), .ZN(n10169) );
  NOR2_X1 U12117 ( .A1(n10164), .A2(n11835), .ZN(n10163) );
  NAND2_X1 U12118 ( .A1(n10187), .A2(n10186), .ZN(n15097) );
  INV_X1 U12119 ( .A(n15094), .ZN(n10186) );
  NOR2_X2 U12120 ( .A1(n15097), .A2(n12488), .ZN(n12516) );
  XNOR2_X1 U12121 ( .A(n12881), .B(n10278), .ZN(n15179) );
  NAND2_X1 U12122 ( .A1(n15183), .A2(n15185), .ZN(n15184) );
  NOR2_X1 U12123 ( .A1(n10173), .A2(n15230), .ZN(n15229) );
  INV_X1 U12124 ( .A(n12980), .ZN(n14030) );
  NAND2_X1 U12125 ( .A1(n10258), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n10257) );
  NOR2_X1 U12126 ( .A1(n12371), .A2(n15300), .ZN(n10258) );
  NAND2_X1 U12127 ( .A1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n12371) );
  NAND2_X1 U12128 ( .A1(n15219), .A2(n9937), .ZN(n15125) );
  OR2_X1 U12129 ( .A1(n15615), .A2(n12221), .ZN(n16240) );
  NAND2_X1 U12130 ( .A1(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n10041) );
  NOR2_X1 U12131 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n13431) );
  AND2_X1 U12132 ( .A1(n11540), .A2(n11539), .ZN(n13888) );
  AND2_X1 U12133 ( .A1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n10044) );
  INV_X1 U12134 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n15459) );
  AND2_X1 U12135 ( .A1(n10104), .A2(n10103), .ZN(n10102) );
  INV_X1 U12136 ( .A(n13850), .ZN(n10103) );
  NOR2_X1 U12137 ( .A1(n16300), .A2(n10045), .ZN(n10043) );
  AND2_X1 U12138 ( .A1(n11971), .A2(n11974), .ZN(n11978) );
  INV_X1 U12139 ( .A(n11981), .ZN(n11989) );
  INV_X1 U12140 ( .A(n9963), .ZN(n9962) );
  OAI21_X1 U12141 ( .B1(n12502), .B2(n9964), .A(n10280), .ZN(n9963) );
  NAND2_X1 U12142 ( .A1(n12493), .A2(n9965), .ZN(n9964) );
  NAND2_X1 U12143 ( .A1(n9967), .A2(n12493), .ZN(n9966) );
  XNOR2_X1 U12144 ( .A(n12277), .B(n12276), .ZN(n15298) );
  NOR2_X1 U12145 ( .A1(n12271), .A2(n12268), .ZN(n15310) );
  AND2_X1 U12146 ( .A1(n9937), .A2(n10119), .ZN(n10118) );
  INV_X1 U12147 ( .A(n15126), .ZN(n10119) );
  OR2_X1 U12148 ( .A1(n15587), .A2(n12449), .ZN(n15533) );
  CLKBUF_X1 U12149 ( .A(n15331), .Z(n15332) );
  NAND2_X1 U12150 ( .A1(n15219), .A2(n9935), .ZN(n15203) );
  NOR3_X1 U12151 ( .A1(n15573), .A2(n10185), .A3(n15572), .ZN(n15547) );
  NOR2_X1 U12152 ( .A1(n15573), .A2(n15572), .ZN(n15575) );
  NAND2_X1 U12153 ( .A1(n15219), .A2(n13349), .ZN(n15201) );
  OR2_X1 U12154 ( .A1(n12237), .A2(n15376), .ZN(n15371) );
  AND2_X1 U12155 ( .A1(n15216), .A2(n15217), .ZN(n15219) );
  AND2_X1 U12156 ( .A1(n11936), .A2(n11935), .ZN(n15847) );
  AND2_X1 U12157 ( .A1(n15632), .A2(n9921), .ZN(n14314) );
  NAND2_X1 U12158 ( .A1(n11558), .A2(n9878), .ZN(n14353) );
  AND2_X1 U12159 ( .A1(n12241), .A2(n15638), .ZN(n15626) );
  INV_X1 U12160 ( .A(n10099), .ZN(n15629) );
  OAI21_X1 U12161 ( .B1(n15445), .B2(n15362), .A(n15444), .ZN(n10099) );
  NAND2_X1 U12162 ( .A1(n15361), .A2(n15660), .ZN(n15445) );
  NAND2_X1 U12163 ( .A1(n10111), .A2(n10114), .ZN(n14016) );
  INV_X1 U12164 ( .A(n13879), .ZN(n10111) );
  NAND2_X1 U12165 ( .A1(n10114), .A2(n10113), .ZN(n10112) );
  INV_X1 U12166 ( .A(n14015), .ZN(n10113) );
  AND2_X1 U12167 ( .A1(n15726), .A2(n9873), .ZN(n14039) );
  INV_X1 U12168 ( .A(n14218), .ZN(n12348) );
  NAND2_X1 U12169 ( .A1(n10180), .A2(n14008), .ZN(n10179) );
  AND2_X1 U12170 ( .A1(n11513), .A2(n11512), .ZN(n13828) );
  NAND2_X1 U12171 ( .A1(n9982), .A2(n9981), .ZN(n9983) );
  INV_X1 U12172 ( .A(n12105), .ZN(n9981) );
  NAND2_X1 U12173 ( .A1(n12443), .A2(n9896), .ZN(n9975) );
  NAND2_X1 U12174 ( .A1(n11616), .A2(n19271), .ZN(n9974) );
  NOR2_X1 U12175 ( .A1(n13863), .A2(n11806), .ZN(n14004) );
  NAND2_X1 U12176 ( .A1(n10160), .A2(n10159), .ZN(n10162) );
  NAND2_X1 U12177 ( .A1(n12694), .A2(n19917), .ZN(n12688) );
  NAND2_X1 U12178 ( .A1(n12443), .A2(n9904), .ZN(n9972) );
  INV_X1 U12179 ( .A(n11616), .ZN(n9973) );
  OAI21_X1 U12180 ( .B1(n9980), .B2(n9979), .A(n11651), .ZN(n9978) );
  NAND2_X1 U12181 ( .A1(n9977), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9976) );
  INV_X1 U12182 ( .A(n19659), .ZN(n19537) );
  INV_X1 U12183 ( .A(n19688), .ZN(n19742) );
  INV_X1 U12184 ( .A(n19270), .ZN(n19296) );
  NOR2_X2 U12185 ( .A1(n14029), .A2(n16305), .ZN(n19295) );
  INV_X1 U12186 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n19735) );
  NOR2_X1 U12187 ( .A1(n16585), .A2(n16584), .ZN(n18684) );
  AOI21_X1 U12188 ( .B1(n13270), .B2(n13272), .A(n13269), .ZN(n18685) );
  NOR2_X1 U12189 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n16813), .ZN(n16799) );
  NOR2_X1 U12190 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n16824), .ZN(n16823) );
  NAND2_X1 U12191 ( .A1(n18904), .A2(n17428), .ZN(n16587) );
  NOR2_X1 U12192 ( .A1(n17230), .A2(n17247), .ZN(n17238) );
  INV_X1 U12193 ( .A(n17266), .ZN(n14395) );
  NOR2_X1 U12194 ( .A1(n17438), .A2(n10012), .ZN(n10011) );
  NOR2_X1 U12195 ( .A1(n17351), .A2(n10018), .ZN(n17315) );
  INV_X1 U12196 ( .A(n17327), .ZN(n10019) );
  OAI21_X1 U12197 ( .B1(n15812), .B2(n15813), .A(n14392), .ZN(n15919) );
  NOR2_X1 U12198 ( .A1(n16589), .A2(n17428), .ZN(n15920) );
  AND3_X1 U12199 ( .A1(n18685), .A2(n18880), .A3(n16584), .ZN(n15921) );
  INV_X1 U12200 ( .A(n17487), .ZN(n17429) );
  INV_X1 U12201 ( .A(n17491), .ZN(n17489) );
  INV_X1 U12202 ( .A(n16581), .ZN(n16580) );
  INV_X1 U12203 ( .A(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n17693) );
  NOR4_X1 U12204 ( .A1(n17810), .A2(n16836), .A3(n17789), .A4(n16816), .ZN(
        n17745) );
  INV_X1 U12205 ( .A(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n17789) );
  INV_X1 U12206 ( .A(n18690), .ZN(n13314) );
  OR2_X1 U12207 ( .A1(n17592), .A2(n13144), .ZN(n13145) );
  NAND2_X1 U12208 ( .A1(n10226), .A2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n10225) );
  INV_X1 U12209 ( .A(n13141), .ZN(n10226) );
  NOR2_X1 U12210 ( .A1(n17775), .A2(n18144), .ZN(n18022) );
  NOR2_X1 U12211 ( .A1(n13312), .A2(n17815), .ZN(n18103) );
  XNOR2_X1 U12212 ( .A(n13128), .B(n13127), .ZN(n17824) );
  INV_X1 U12213 ( .A(n13129), .ZN(n13127) );
  NOR2_X1 U12214 ( .A1(n17849), .A2(n17848), .ZN(n17847) );
  XNOR2_X1 U12215 ( .A(n13121), .B(n13120), .ZN(n17846) );
  INV_X1 U12216 ( .A(n13119), .ZN(n13120) );
  NAND2_X1 U12217 ( .A1(n17846), .A2(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n17845) );
  NOR2_X1 U12218 ( .A1(n17414), .A2(n13108), .ZN(n13114) );
  OR2_X1 U12219 ( .A1(n13287), .A2(n13110), .ZN(n13111) );
  INV_X1 U12220 ( .A(n15816), .ZN(n15803) );
  NAND2_X1 U12221 ( .A1(n10221), .A2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n10220) );
  INV_X1 U12222 ( .A(n10272), .ZN(n10221) );
  NOR2_X1 U12223 ( .A1(n15822), .A2(n15807), .ZN(n16454) );
  NAND2_X1 U12224 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n18700) );
  NAND2_X1 U12225 ( .A1(n15802), .A2(n10020), .ZN(n15816) );
  AOI21_X1 U12226 ( .B1(n14391), .B2(n13251), .A(n10021), .ZN(n10020) );
  AND2_X1 U12227 ( .A1(n15920), .A2(n17356), .ZN(n13251) );
  INV_X1 U12228 ( .A(n15804), .ZN(n10021) );
  NOR2_X1 U12229 ( .A1(n13189), .A2(n13188), .ZN(n18248) );
  NOR2_X1 U12230 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18245), .ZN(n18532) );
  NOR2_X1 U12231 ( .A1(n13217), .A2(n13216), .ZN(n18267) );
  INV_X1 U12232 ( .A(n13274), .ZN(n18271) );
  INV_X1 U12233 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n18901) );
  INV_X2 U12234 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n20802) );
  AND2_X1 U12235 ( .A1(n15935), .A2(n11286), .ZN(n14592) );
  INV_X1 U12236 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n15999) );
  INV_X1 U12237 ( .A(n20038), .ZN(n20010) );
  INV_X1 U12238 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n19967) );
  OR2_X1 U12239 ( .A1(n20023), .A2(n19980), .ZN(n19999) );
  OR2_X1 U12240 ( .A1(n11282), .A2(n11279), .ZN(n20023) );
  OR3_X1 U12241 ( .A1(n20808), .A2(n20103), .A3(n11171), .ZN(n20022) );
  OR2_X1 U12242 ( .A1(n13806), .A2(n19943), .ZN(n13812) );
  INV_X2 U12243 ( .A(n14718), .ZN(n14748) );
  NAND2_X1 U12244 ( .A1(n10209), .A2(n10210), .ZN(n14753) );
  NAND2_X1 U12245 ( .A1(n14557), .A2(n14558), .ZN(n10209) );
  INV_X1 U12246 ( .A(n14803), .ZN(n14798) );
  INV_X1 U12247 ( .A(n14802), .ZN(n14796) );
  NAND2_X1 U12248 ( .A1(n12540), .A2(n12539), .ZN(n20043) );
  OR2_X1 U12249 ( .A1(n14816), .A2(n13619), .ZN(n14814) );
  AND2_X1 U12250 ( .A1(n13418), .A2(n13417), .ZN(n20047) );
  BUF_X1 U12251 ( .A(n20071), .Z(n20064) );
  OR2_X1 U12252 ( .A1(n11172), .A2(n14560), .ZN(n11173) );
  INV_X1 U12253 ( .A(n14753), .ZN(n14824) );
  NAND2_X1 U12254 ( .A1(n14557), .A2(n12657), .ZN(n14509) );
  OR2_X1 U12255 ( .A1(n12656), .A2(n12655), .ZN(n12657) );
  AND2_X1 U12256 ( .A1(n14900), .A2(n12663), .ZN(n16077) );
  INV_X1 U12257 ( .A(n20097), .ZN(n20159) );
  INV_X1 U12258 ( .A(n14900), .ZN(n20091) );
  AND2_X1 U12259 ( .A1(n13418), .A2(n15880), .ZN(n20098) );
  AND2_X1 U12260 ( .A1(n20775), .A2(n12659), .ZN(n20097) );
  INV_X1 U12261 ( .A(n20098), .ZN(n19949) );
  AND2_X1 U12262 ( .A1(n14586), .A2(n14585), .ZN(n14972) );
  MUX2_X1 U12263 ( .A(n14839), .B(n14838), .S(n9913), .Z(n14841) );
  NAND2_X1 U12264 ( .A1(n14163), .A2(n14161), .ZN(n10034) );
  OAI21_X1 U12265 ( .B1(n20094), .B2(n10125), .A(n10124), .ZN(n16098) );
  NAND2_X1 U12266 ( .A1(n20092), .A2(n12600), .ZN(n16100) );
  OR2_X1 U12267 ( .A1(n14168), .A2(n15054), .ZN(n20120) );
  OR2_X1 U12268 ( .A1(n14165), .A2(n13395), .ZN(n20145) );
  OR2_X1 U12269 ( .A1(n14165), .A2(n13785), .ZN(n14167) );
  INV_X1 U12270 ( .A(n12563), .ZN(n10543) );
  INV_X1 U12271 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20461) );
  INV_X1 U12272 ( .A(n10536), .ZN(n10030) );
  NOR2_X1 U12273 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n15073) );
  OAI21_X1 U12274 ( .B1(n20315), .B2(n20298), .A(n20598), .ZN(n20316) );
  INV_X1 U12275 ( .A(n20369), .ZN(n20378) );
  NOR2_X1 U12276 ( .A1(n20790), .A2(n20380), .ZN(n20401) );
  AND2_X1 U12277 ( .A1(n20383), .A2(n20462), .ZN(n20402) );
  AND2_X1 U12278 ( .A1(n20439), .A2(n20562), .ZN(n20484) );
  NAND2_X1 U12279 ( .A1(n20776), .A2(n20462), .ZN(n20513) );
  OAI211_X1 U12280 ( .C1(n20623), .C2(n20599), .A(n20598), .B(n20597), .ZN(
        n20626) );
  INV_X1 U12281 ( .A(n20681), .ZN(n20688) );
  AND2_X1 U12282 ( .A1(n11160), .A2(n11159), .ZN(n15901) );
  OAI21_X1 U12283 ( .B1(n11158), .B2(n11157), .A(n11156), .ZN(n11160) );
  AND2_X1 U12284 ( .A1(n11155), .A2(n13492), .ZN(n11157) );
  INV_X1 U12285 ( .A(n15897), .ZN(n20695) );
  INV_X1 U12286 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n20413) );
  AOI221_X1 U12287 ( .B1(n20806), .B2(n13782), .C1(n15896), .C2(n13782), .A(
        n16203), .ZN(n16207) );
  AND2_X1 U12288 ( .A1(n10051), .A2(n10049), .ZN(n13329) );
  AND2_X1 U12289 ( .A1(n10052), .A2(n10050), .ZN(n10049) );
  INV_X1 U12290 ( .A(n15302), .ZN(n10050) );
  NAND2_X1 U12291 ( .A1(n10051), .A2(n10052), .ZN(n13330) );
  AND2_X1 U12292 ( .A1(n10054), .A2(n15313), .ZN(n16216) );
  NOR2_X1 U12293 ( .A1(n15324), .A2(n15120), .ZN(n15119) );
  NOR2_X1 U12294 ( .A1(n10053), .A2(n15135), .ZN(n15120) );
  NAND2_X1 U12295 ( .A1(n10048), .A2(n10047), .ZN(n15110) );
  NAND2_X1 U12296 ( .A1(n10053), .A2(n10070), .ZN(n10068) );
  NAND2_X1 U12297 ( .A1(n10067), .A2(n10065), .ZN(n10063) );
  NOR2_X1 U12298 ( .A1(n18943), .A2(n18959), .ZN(n10065) );
  AND2_X1 U12299 ( .A1(n10067), .A2(n10066), .ZN(n18958) );
  NOR2_X1 U12300 ( .A1(n12175), .A2(n10075), .ZN(n12178) );
  INV_X1 U12301 ( .A(n19101), .ZN(n19057) );
  INV_X1 U12302 ( .A(n19090), .ZN(n19072) );
  AND2_X1 U12303 ( .A1(n12107), .A2(n10058), .ZN(n12104) );
  NOR2_X1 U12304 ( .A1(n10060), .A2(n10059), .ZN(n10058) );
  INV_X1 U12305 ( .A(n12125), .ZN(n10059) );
  INV_X1 U12306 ( .A(n19088), .ZN(n19087) );
  INV_X1 U12307 ( .A(n19049), .ZN(n19095) );
  AND2_X1 U12308 ( .A1(n19074), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19101) );
  AND2_X1 U12309 ( .A1(n11558), .A2(n9881), .ZN(n14324) );
  OR2_X1 U12310 ( .A1(n11903), .A2(n11902), .ZN(n14064) );
  OR2_X1 U12311 ( .A1(n11888), .A2(n11887), .ZN(n14020) );
  OR2_X1 U12312 ( .A1(n11848), .A2(n11847), .ZN(n13921) );
  NAND2_X1 U12313 ( .A1(n9879), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n10164) );
  INV_X1 U12314 ( .A(n15215), .ZN(n15231) );
  INV_X1 U12315 ( .A(n13827), .ZN(n10165) );
  OR2_X1 U12316 ( .A1(n15192), .A2(n10156), .ZN(n15215) );
  AND2_X1 U12317 ( .A1(n15095), .A2(n13338), .ZN(n15486) );
  AND2_X1 U12318 ( .A1(n13574), .A2(n14030), .ZN(n19110) );
  NOR2_X1 U12319 ( .A1(n19116), .A2(n19156), .ZN(n19147) );
  INV_X1 U12320 ( .A(n19140), .ZN(n19155) );
  INV_X1 U12321 ( .A(n19160), .ZN(n19116) );
  OR2_X1 U12322 ( .A1(n19108), .A2(n13574), .ZN(n19129) );
  OR2_X1 U12323 ( .A1(n12678), .A2(n13562), .ZN(n14119) );
  NOR2_X1 U12324 ( .A1(n13335), .A2(n13334), .ZN(n15485) );
  NAND2_X1 U12325 ( .A1(n9906), .A2(n12357), .ZN(n9993) );
  INV_X1 U12326 ( .A(n16302), .ZN(n19256) );
  NAND2_X1 U12327 ( .A1(n19907), .A2(n19747), .ZN(n16305) );
  INV_X1 U12328 ( .A(n16295), .ZN(n19251) );
  INV_X1 U12329 ( .A(n16310), .ZN(n19246) );
  NAND2_X1 U12330 ( .A1(n12495), .A2(n12493), .ZN(n12501) );
  AOI21_X1 U12331 ( .B1(n12527), .B2(n16340), .A(n12526), .ZN(n12530) );
  INV_X1 U12332 ( .A(n10235), .ZN(n10234) );
  AOI21_X1 U12333 ( .B1(n15361), .B2(n12247), .A(n12246), .ZN(n15353) );
  XNOR2_X1 U12334 ( .A(n10094), .B(n9923), .ZN(n15585) );
  NAND2_X1 U12335 ( .A1(n15382), .A2(n10095), .ZN(n10094) );
  INV_X1 U12336 ( .A(n15383), .ZN(n10095) );
  INV_X1 U12337 ( .A(n15615), .ZN(n15624) );
  AND2_X1 U12338 ( .A1(n12465), .A2(n15665), .ZN(n16311) );
  AND2_X1 U12339 ( .A1(n9985), .A2(n15615), .ZN(n16247) );
  NAND2_X1 U12340 ( .A1(n15625), .A2(n15638), .ZN(n9985) );
  NAND2_X1 U12341 ( .A1(n10213), .A2(n10212), .ZN(n15673) );
  NAND2_X1 U12342 ( .A1(n9986), .A2(n9992), .ZN(n15708) );
  NAND2_X1 U12343 ( .A1(n9988), .A2(n9994), .ZN(n9986) );
  NAND2_X1 U12344 ( .A1(n12360), .A2(n12361), .ZN(n15453) );
  NAND2_X1 U12345 ( .A1(n10252), .A2(n12362), .ZN(n15454) );
  INV_X1 U12346 ( .A(n12673), .ZN(n13584) );
  INV_X1 U12347 ( .A(n15613), .ZN(n16351) );
  INV_X1 U12348 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19924) );
  INV_X1 U12349 ( .A(n14119), .ZN(n19921) );
  INV_X1 U12350 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19905) );
  INV_X1 U12351 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n15918) );
  AND2_X1 U12352 ( .A1(n13580), .A2(n13583), .ZN(n19910) );
  NAND2_X1 U12353 ( .A1(n13837), .A2(n13627), .ZN(n19901) );
  XNOR2_X1 U12354 ( .A(n13841), .B(n13840), .ZN(n19539) );
  NAND2_X1 U12355 ( .A1(n13837), .A2(n13836), .ZN(n13841) );
  NAND2_X1 U12356 ( .A1(n14128), .A2(n14127), .ZN(n19350) );
  OAI21_X1 U12357 ( .B1(n19393), .B2(n19392), .A(n19391), .ZN(n19411) );
  NOR2_X1 U12358 ( .A1(n19447), .A2(n19658), .ZN(n19439) );
  OAI21_X1 U12359 ( .B1(n19530), .B2(n19509), .A(n19747), .ZN(n19533) );
  NOR2_X1 U12360 ( .A1(n19476), .A2(n19688), .ZN(n19531) );
  INV_X1 U12361 ( .A(n19604), .ZN(n19595) );
  OAI21_X1 U12362 ( .B1(n19582), .B2(n19581), .A(n19580), .ZN(n19600) );
  INV_X1 U12363 ( .A(n19635), .ZN(n19599) );
  AOI211_X2 U12364 ( .C1(n14028), .C2(n14027), .A(n14026), .B(n19389), .ZN(
        n19657) );
  NOR2_X1 U12365 ( .A1(n19665), .A2(n19662), .ZN(n19683) );
  INV_X1 U12366 ( .A(n19784), .ZN(n19719) );
  OAI21_X1 U12367 ( .B1(n19700), .B2(n19699), .A(n19698), .ZN(n19729) );
  INV_X1 U12368 ( .A(n19703), .ZN(n19749) );
  INV_X1 U12369 ( .A(n19257), .ZN(n19740) );
  INV_X1 U12370 ( .A(n19707), .ZN(n19755) );
  INV_X1 U12371 ( .A(n19711), .ZN(n19761) );
  AND2_X1 U12372 ( .A1(n19275), .A2(n19296), .ZN(n19759) );
  INV_X1 U12373 ( .A(n19623), .ZN(n19767) );
  INV_X1 U12374 ( .A(n19717), .ZN(n19773) );
  AND2_X1 U12375 ( .A1(n19281), .A2(n19296), .ZN(n19771) );
  INV_X1 U12376 ( .A(n19800), .ZN(n19780) );
  AND2_X1 U12377 ( .A1(n19286), .A2(n19296), .ZN(n19777) );
  INV_X1 U12378 ( .A(n19726), .ZN(n19787) );
  NOR2_X2 U12379 ( .A1(n19689), .A2(n19688), .ZN(n19796) );
  NOR2_X1 U12380 ( .A1(n19744), .A2(n19739), .ZN(n19794) );
  AND2_X1 U12381 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n11636), .ZN(n19808) );
  NAND2_X1 U12382 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n21058), .ZN(n19937) );
  XOR2_X1 U12383 ( .A(n18886), .B(n18248), .Z(n18903) );
  NOR2_X1 U12384 ( .A1(n18684), .A2(n17491), .ZN(n18904) );
  NAND2_X1 U12385 ( .A1(n18884), .A2(n18685), .ZN(n17491) );
  NAND2_X1 U12386 ( .A1(n13314), .A2(n18884), .ZN(n16560) );
  NOR2_X1 U12387 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n16679), .ZN(n16660) );
  NOR2_X1 U12388 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n16745), .ZN(n16728) );
  NOR2_X1 U12389 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n16790), .ZN(n16775) );
  NOR2_X1 U12390 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n16894), .ZN(n16875) );
  INV_X1 U12391 ( .A(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n16924) );
  NAND2_X1 U12392 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n16958), .ZN(n16925) );
  INV_X1 U12393 ( .A(n16925), .ZN(n16944) );
  INV_X1 U12394 ( .A(n16930), .ZN(n16958) );
  INV_X1 U12395 ( .A(n16936), .ZN(n16954) );
  NOR2_X1 U12396 ( .A1(n17093), .A2(n17090), .ZN(n17077) );
  NAND2_X1 U12397 ( .A1(P3_EBX_REG_19__SCAN_IN), .A2(n17077), .ZN(n17076) );
  INV_X1 U12398 ( .A(n17131), .ZN(n17107) );
  NAND2_X1 U12399 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(n15796), .ZN(n17134) );
  NOR2_X1 U12400 ( .A1(n17189), .A2(n17207), .ZN(n17174) );
  NAND2_X1 U12401 ( .A1(P3_EBX_REG_11__SCAN_IN), .A2(n17174), .ZN(n17173) );
  NOR2_X1 U12402 ( .A1(n17233), .A2(n17210), .ZN(n17208) );
  NAND2_X1 U12403 ( .A1(P3_EBX_REG_9__SCAN_IN), .A2(n17208), .ZN(n17207) );
  INV_X1 U12404 ( .A(n17282), .ZN(n17277) );
  NAND2_X1 U12405 ( .A1(n17300), .A2(n9885), .ZN(n17291) );
  INV_X1 U12406 ( .A(n17304), .ZN(n17300) );
  NAND2_X1 U12407 ( .A1(n17300), .A2(P3_EAX_REG_25__SCAN_IN), .ZN(n17299) );
  NOR2_X1 U12408 ( .A1(n17356), .A2(n17309), .ZN(n17305) );
  NOR2_X1 U12409 ( .A1(n17314), .A2(n17444), .ZN(n17310) );
  NAND2_X1 U12410 ( .A1(n17310), .A2(P3_EAX_REG_23__SCAN_IN), .ZN(n17309) );
  NAND2_X1 U12411 ( .A1(n17315), .A2(P3_EAX_REG_21__SCAN_IN), .ZN(n17314) );
  NAND2_X1 U12412 ( .A1(P3_EAX_REG_16__SCAN_IN), .A2(n17352), .ZN(n17351) );
  NOR2_X1 U12413 ( .A1(n17388), .A2(n10013), .ZN(n17271) );
  INV_X1 U12414 ( .A(n17363), .ZN(n10014) );
  AND2_X1 U12415 ( .A1(n17272), .A2(n17356), .ZN(n17375) );
  NAND2_X1 U12416 ( .A1(n17399), .A2(P3_EAX_REG_7__SCAN_IN), .ZN(n17388) );
  NOR2_X1 U12417 ( .A1(n13094), .A2(n13093), .ZN(n17397) );
  NOR2_X1 U12418 ( .A1(n17420), .A2(n10015), .ZN(n17399) );
  NAND2_X1 U12419 ( .A1(n10016), .A2(P3_EAX_REG_6__SCAN_IN), .ZN(n10015) );
  INV_X1 U12420 ( .A(n17396), .ZN(n10016) );
  INV_X1 U12421 ( .A(n13281), .ZN(n17401) );
  NAND2_X1 U12422 ( .A1(n18713), .A2(n17272), .ZN(n17415) );
  INV_X1 U12423 ( .A(n17423), .ZN(n17418) );
  OAI21_X1 U12424 ( .B1(n15921), .B2(n10017), .A(n18884), .ZN(n17420) );
  AND2_X1 U12425 ( .A1(n15919), .A2(n15920), .ZN(n10017) );
  NOR2_X1 U12426 ( .A1(n10218), .A2(n10217), .ZN(n10216) );
  INV_X1 U12427 ( .A(n13105), .ZN(n10217) );
  CLKBUF_X1 U12428 ( .A(n17470), .Z(n17484) );
  CLKBUF_X1 U12430 ( .A(n17536), .Z(n17529) );
  INV_X1 U12431 ( .A(n17539), .ZN(n17530) );
  OR2_X1 U12432 ( .A1(n17491), .A2(n18735), .ZN(n17539) );
  NOR2_X1 U12433 ( .A1(n17529), .A2(n18886), .ZN(n17537) );
  INV_X1 U12434 ( .A(n17598), .ZN(n17822) );
  NAND2_X1 U12435 ( .A1(n18532), .A2(n18593), .ZN(n18343) );
  NAND2_X1 U12436 ( .A1(n17867), .A2(n17910), .ZN(n17905) );
  INV_X1 U12437 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n17904) );
  INV_X1 U12438 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n18236) );
  INV_X1 U12439 ( .A(n16447), .ZN(n15819) );
  OR2_X1 U12440 ( .A1(n17687), .A2(n10225), .ZN(n17612) );
  NOR2_X1 U12441 ( .A1(n17687), .A2(n13141), .ZN(n17637) );
  AND2_X1 U12442 ( .A1(n9890), .A2(n10244), .ZN(n17696) );
  NAND2_X1 U12443 ( .A1(n17705), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n10244) );
  CLKBUF_X1 U12444 ( .A(n17879), .Z(n18189) );
  AOI21_X2 U12445 ( .B1(n15833), .B2(n15832), .A(n18743), .ZN(n18227) );
  INV_X1 U12446 ( .A(n18224), .ZN(n18230) );
  INV_X1 U12447 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18723) );
  INV_X1 U12448 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n18727) );
  OAI21_X1 U12450 ( .B1(n14663), .B2(n20038), .A(n9900), .ZN(P1_U2809) );
  AOI21_X1 U12451 ( .B1(n10580), .B2(n20774), .A(n9938), .ZN(n20779) );
  AND2_X1 U12452 ( .A1(n11764), .A2(n11763), .ZN(n11966) );
  AND3_X1 U12453 ( .A1(n10178), .A2(n10177), .A3(n10176), .ZN(n12481) );
  INV_X1 U12454 ( .A(n12492), .ZN(n12499) );
  AOI21_X1 U12455 ( .B1(n16443), .B2(n17598), .A(n13321), .ZN(n13322) );
  OAI21_X1 U12456 ( .B1(n16446), .B2(n17914), .A(n13320), .ZN(n13321) );
  NAND2_X1 U12457 ( .A1(n11317), .A2(n10062), .ZN(n11312) );
  NAND2_X2 U12458 ( .A1(n12970), .A2(n11789), .ZN(n11817) );
  CLKBUF_X3 U12459 ( .A(n13088), .Z(n17213) );
  NAND2_X1 U12460 ( .A1(n15674), .A2(n10254), .ZN(n15386) );
  NAND2_X1 U12461 ( .A1(n15112), .A2(n15113), .ZN(n15111) );
  AND2_X1 U12462 ( .A1(n10475), .A2(n10026), .ZN(n9869) );
  NOR2_X1 U12463 ( .A1(n14721), .A2(n9916), .ZN(n14605) );
  NAND2_X1 U12464 ( .A1(n10193), .A2(n10197), .ZN(n14625) );
  AND2_X1 U12465 ( .A1(n13279), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n9870) );
  AND4_X1 U12466 ( .A1(n13193), .A2(n13192), .A3(n13191), .A4(n13190), .ZN(
        n9871) );
  OR2_X1 U12467 ( .A1(n12347), .A2(n14226), .ZN(n12351) );
  INV_X1 U12468 ( .A(n12351), .ZN(n10249) );
  NAND2_X1 U12469 ( .A1(n12206), .A2(n9922), .ZN(n9872) );
  NOR2_X1 U12470 ( .A1(n11838), .A2(n10183), .ZN(n9873) );
  AND2_X1 U12471 ( .A1(n11439), .A2(n11458), .ZN(n9874) );
  INV_X1 U12472 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n16300) );
  AND2_X1 U12473 ( .A1(n14138), .A2(n9917), .ZN(n9875) );
  NAND2_X1 U12474 ( .A1(n15632), .A2(n16312), .ZN(n15846) );
  OR2_X1 U12475 ( .A1(n11321), .A2(n9914), .ZN(n9876) );
  AND3_X1 U12476 ( .A1(n10046), .A2(n10043), .A3(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n9877) );
  AND2_X1 U12477 ( .A1(n11557), .A2(n10107), .ZN(n9878) );
  NAND2_X1 U12478 ( .A1(n14138), .A2(n14209), .ZN(n14208) );
  NAND2_X1 U12479 ( .A1(n11558), .A2(n11557), .ZN(n14141) );
  AND2_X1 U12480 ( .A1(n13827), .A2(n12700), .ZN(n9879) );
  NOR2_X1 U12481 ( .A1(n11751), .A2(n10080), .ZN(n9880) );
  AND2_X1 U12482 ( .A1(n11317), .A2(n9924), .ZN(n11313) );
  NOR2_X1 U12483 ( .A1(n15196), .A2(n12819), .ZN(n15188) );
  AND2_X1 U12484 ( .A1(n9878), .A2(n10106), .ZN(n9881) );
  INV_X1 U12485 ( .A(n10173), .ZN(n14382) );
  AND2_X1 U12486 ( .A1(n9921), .A2(n14315), .ZN(n9882) );
  NAND2_X1 U12487 ( .A1(n10628), .A2(n10579), .ZN(n20772) );
  INV_X1 U12488 ( .A(n10168), .ZN(n13950) );
  INV_X1 U12489 ( .A(n10167), .ZN(n14019) );
  AND2_X1 U12490 ( .A1(n10254), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n9883) );
  AND2_X1 U12491 ( .A1(n9883), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n9884) );
  AND2_X1 U12492 ( .A1(n10011), .A2(P3_EAX_REG_27__SCAN_IN), .ZN(n9885) );
  AND2_X2 U12493 ( .A1(n15743), .A2(n12799), .ZN(n11667) );
  OR3_X1 U12494 ( .A1(n13359), .A2(n12417), .A3(n15532), .ZN(n9886) );
  OR2_X1 U12495 ( .A1(n12362), .A2(n15730), .ZN(n9889) );
  NAND2_X1 U12496 ( .A1(n10162), .A2(n11982), .ZN(n10161) );
  AND2_X1 U12497 ( .A1(n13137), .A2(n13136), .ZN(n9890) );
  XNOR2_X1 U12498 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n12419), .ZN(
        n9891) );
  NAND2_X1 U12499 ( .A1(n14683), .A2(n14676), .ZN(n14670) );
  NAND2_X1 U12500 ( .A1(n9859), .A2(n12571), .ZN(n11250) );
  INV_X1 U12501 ( .A(n12502), .ZN(n9967) );
  AND2_X1 U12502 ( .A1(n15674), .A2(n9884), .ZN(n15340) );
  AND2_X1 U12503 ( .A1(n15674), .A2(n9883), .ZN(n15375) );
  NOR2_X1 U12504 ( .A1(n15331), .A2(n15333), .ZN(n15317) );
  NAND2_X1 U12505 ( .A1(n14674), .A2(n14675), .ZN(n14667) );
  NOR2_X1 U12506 ( .A1(n17605), .A2(n10222), .ZN(n9892) );
  NAND2_X1 U12507 ( .A1(n15398), .A2(n15399), .ZN(n9893) );
  OR2_X1 U12508 ( .A1(n13618), .A2(n10409), .ZN(n9894) );
  INV_X2 U12509 ( .A(n12412), .ZN(n19286) );
  INV_X1 U12510 ( .A(n11180), .ZN(n9958) );
  OR2_X2 U12511 ( .A1(n10329), .A2(n10328), .ZN(n10417) );
  NAND2_X1 U12512 ( .A1(n10088), .A2(n10089), .ZN(n15662) );
  NAND2_X1 U12513 ( .A1(n9993), .A2(n9996), .ZN(n16287) );
  NAND2_X1 U12514 ( .A1(n10158), .A2(n12677), .ZN(n12678) );
  AND2_X1 U12515 ( .A1(n14674), .A2(n10199), .ZN(n14580) );
  OR3_X1 U12516 ( .A1(n12524), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n12523), .ZN(n9895) );
  AND3_X1 U12517 ( .A1(n11419), .A2(n19297), .A3(n19271), .ZN(n9896) );
  OR2_X1 U12518 ( .A1(n12862), .A2(n12861), .ZN(n9897) );
  AND3_X1 U12519 ( .A1(n13196), .A2(n13194), .A3(n13197), .ZN(n9898) );
  AND2_X1 U12520 ( .A1(n15310), .A2(n15319), .ZN(n9899) );
  AND2_X1 U12521 ( .A1(n11291), .A2(n11290), .ZN(n9900) );
  AND3_X1 U12522 ( .A1(n9858), .A2(n11112), .A3(n12571), .ZN(n9901) );
  OR2_X1 U12523 ( .A1(n14509), .A2(n20159), .ZN(n9902) );
  AND2_X1 U12524 ( .A1(n9994), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n9903) );
  AND2_X1 U12525 ( .A1(n11419), .A2(n19297), .ZN(n9904) );
  INV_X1 U12526 ( .A(n15802), .ZN(n16585) );
  NAND2_X1 U12527 ( .A1(n16559), .A2(n18903), .ZN(n15802) );
  INV_X1 U12528 ( .A(n11459), .ZN(n12380) );
  BUF_X1 U12529 ( .A(n11459), .Z(n19275) );
  AND2_X1 U12530 ( .A1(n10522), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n9905) );
  INV_X1 U12531 ( .A(n13625), .ZN(n13622) );
  AND2_X1 U12532 ( .A1(n12356), .A2(n9889), .ZN(n9906) );
  NAND2_X1 U12533 ( .A1(n15252), .A2(n15251), .ZN(n13336) );
  OR2_X1 U12534 ( .A1(n10473), .A2(n10472), .ZN(n10475) );
  AND2_X1 U12535 ( .A1(n15161), .A2(n15160), .ZN(n15159) );
  OR2_X1 U12536 ( .A1(n10233), .A2(n12246), .ZN(n9907) );
  AND2_X1 U12537 ( .A1(n10272), .A2(n13107), .ZN(n9908) );
  OR2_X1 U12538 ( .A1(n12497), .A2(n12523), .ZN(n9909) );
  NAND2_X1 U12539 ( .A1(n17823), .A2(n13130), .ZN(n13279) );
  INV_X1 U12540 ( .A(n10521), .ZN(n10522) );
  AND2_X1 U12541 ( .A1(n9873), .A2(n14040), .ZN(n9910) );
  AND2_X1 U12542 ( .A1(n11462), .A2(n12392), .ZN(n9911) );
  NAND2_X1 U12543 ( .A1(n16081), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n9912) );
  INV_X2 U12544 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n15754) );
  NAND2_X1 U12545 ( .A1(n15184), .A2(n9897), .ZN(n12881) );
  NOR2_X1 U12546 ( .A1(n11319), .A2(n11332), .ZN(n11317) );
  NAND2_X1 U12547 ( .A1(n12305), .A2(n11637), .ZN(n12434) );
  NAND2_X1 U12548 ( .A1(n14138), .A2(n9920), .ZN(n10173) );
  OR2_X1 U12549 ( .A1(n16266), .A2(n10042), .ZN(n9914) );
  NAND2_X1 U12550 ( .A1(n11823), .A2(n11822), .ZN(n15726) );
  AND3_X1 U12551 ( .A1(n11440), .A2(n12434), .A3(n9874), .ZN(n12421) );
  NAND2_X1 U12552 ( .A1(n15726), .A2(n15725), .ZN(n14184) );
  NOR2_X1 U12553 ( .A1(n12175), .A2(n10077), .ZN(n12169) );
  NOR2_X1 U12554 ( .A1(n14322), .A2(n14381), .ZN(n14380) );
  INV_X1 U12555 ( .A(n16050), .ZN(n10148) );
  NOR3_X1 U12556 ( .A1(n11321), .A2(n9914), .A3(n10041), .ZN(n11318) );
  NOR2_X1 U12557 ( .A1(n14721), .A2(n14722), .ZN(n14624) );
  NAND2_X1 U12558 ( .A1(n15632), .A2(n9882), .ZN(n14313) );
  NAND2_X1 U12559 ( .A1(n14254), .A2(n10205), .ZN(n14368) );
  NOR3_X1 U12560 ( .A1(n11321), .A2(n9914), .A3(n15448), .ZN(n11320) );
  NOR2_X1 U12561 ( .A1(n11325), .A2(n15459), .ZN(n11326) );
  NOR2_X1 U12562 ( .A1(n11323), .A2(n16278), .ZN(n11324) );
  NOR2_X1 U12563 ( .A1(n11321), .A2(n16266), .ZN(n11322) );
  NOR2_X1 U12564 ( .A1(n11329), .A2(n11328), .ZN(n11330) );
  INV_X1 U12565 ( .A(n11329), .ZN(n10046) );
  AND2_X1 U12566 ( .A1(n17300), .A2(n10011), .ZN(n9915) );
  OR2_X1 U12567 ( .A1(n13581), .A2(n13582), .ZN(n13580) );
  OR2_X1 U12568 ( .A1(n10196), .A2(n14710), .ZN(n9916) );
  AND2_X1 U12569 ( .A1(n10175), .A2(n14209), .ZN(n9917) );
  AND2_X1 U12570 ( .A1(n10169), .A2(n14020), .ZN(n9918) );
  AND2_X1 U12571 ( .A1(n11317), .A2(n11292), .ZN(n11315) );
  OR2_X1 U12572 ( .A1(n14818), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n9919) );
  NOR2_X1 U12573 ( .A1(n13879), .A2(n10112), .ZN(n14017) );
  INV_X1 U12574 ( .A(n15350), .ZN(n10236) );
  AND2_X1 U12575 ( .A1(n9917), .A2(n12737), .ZN(n9920) );
  NAND2_X1 U12576 ( .A1(n10141), .A2(n12637), .ZN(n14280) );
  AND2_X1 U12577 ( .A1(n10182), .A2(n16312), .ZN(n9921) );
  NAND2_X1 U12578 ( .A1(n10034), .A2(n14160), .ZN(n16089) );
  NAND2_X1 U12579 ( .A1(n10081), .A2(n12131), .ZN(n14329) );
  AND2_X1 U12580 ( .A1(n9880), .A2(n10079), .ZN(n9922) );
  OR2_X1 U12581 ( .A1(n15385), .A2(n15384), .ZN(n9923) );
  INV_X1 U12582 ( .A(n12108), .ZN(n10060) );
  NAND2_X1 U12583 ( .A1(n11456), .A2(n10154), .ZN(n12374) );
  NAND2_X1 U12584 ( .A1(n20182), .A2(n11112), .ZN(n11105) );
  XNOR2_X1 U12585 ( .A(n12862), .B(n12858), .ZN(n15183) );
  INV_X1 U12586 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n11328) );
  XNOR2_X1 U12587 ( .A(n12817), .B(n12841), .ZN(n15195) );
  AND2_X1 U12588 ( .A1(n11292), .A2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n9924) );
  OR2_X1 U12589 ( .A1(n11700), .A2(n11699), .ZN(n11813) );
  NOR2_X1 U12590 ( .A1(n15188), .A2(n15189), .ZN(n9925) );
  NAND2_X1 U12591 ( .A1(n12327), .A2(n12328), .ZN(n9926) );
  AND2_X1 U12592 ( .A1(n10428), .A2(n10427), .ZN(n13399) );
  NAND2_X1 U12593 ( .A1(n11794), .A2(n19281), .ZN(n12379) );
  NOR2_X1 U12594 ( .A1(n14818), .A2(n14961), .ZN(n9927) );
  INV_X1 U12595 ( .A(n10076), .ZN(n12269) );
  NOR2_X1 U12596 ( .A1(n12175), .A2(n12412), .ZN(n10076) );
  AND2_X1 U12597 ( .A1(n10199), .A2(n14582), .ZN(n9928) );
  AND2_X1 U12598 ( .A1(n14380), .A2(n11573), .ZN(n15216) );
  AND2_X1 U12599 ( .A1(n9922), .A2(n15213), .ZN(n9929) );
  INV_X1 U12600 ( .A(n11593), .ZN(n15175) );
  NOR2_X1 U12601 ( .A1(n15111), .A2(n15176), .ZN(n11593) );
  AND2_X1 U12602 ( .A1(n15219), .A2(n10118), .ZN(n15112) );
  NAND2_X1 U12603 ( .A1(n10631), .A2(n10630), .ZN(n9930) );
  NAND2_X1 U12604 ( .A1(n10028), .A2(n13758), .ZN(n13707) );
  INV_X1 U12605 ( .A(n10093), .ZN(n10092) );
  OAI21_X1 U12606 ( .B1(n10212), .B2(n15676), .A(n15671), .ZN(n10093) );
  AND3_X1 U12607 ( .A1(n15699), .A2(n15694), .A3(n15717), .ZN(n9931) );
  INV_X1 U12608 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n15448) );
  OR2_X1 U12609 ( .A1(n11834), .A2(n11833), .ZN(n13883) );
  NOR2_X1 U12610 ( .A1(n11501), .A2(n11500), .ZN(n11504) );
  AND2_X1 U12611 ( .A1(n9858), .A2(n11112), .ZN(n12630) );
  AND2_X1 U12612 ( .A1(n9918), .A2(n14064), .ZN(n9932) );
  AND2_X1 U12613 ( .A1(n9882), .A2(n11939), .ZN(n9933) );
  OR2_X1 U12614 ( .A1(n11014), .A2(n11013), .ZN(n14595) );
  INV_X1 U12615 ( .A(n15212), .ZN(n15234) );
  INV_X1 U12616 ( .A(n16326), .ZN(n16340) );
  NAND2_X1 U12617 ( .A1(n13876), .A2(n13875), .ZN(n13874) );
  NOR2_X1 U12618 ( .A1(n10166), .A2(n10165), .ZN(n13766) );
  NAND2_X1 U12619 ( .A1(n13864), .A2(n10180), .ZN(n14005) );
  NOR2_X1 U12620 ( .A1(n13879), .A2(n10116), .ZN(n13926) );
  NAND2_X1 U12621 ( .A1(n19079), .A2(n11334), .ZN(n10067) );
  NOR2_X1 U12622 ( .A1(n11306), .A2(n15304), .ZN(n11302) );
  NOR2_X1 U12623 ( .A1(n13879), .A2(n13888), .ZN(n13889) );
  NAND2_X1 U12624 ( .A1(n12702), .A2(n10279), .ZN(n13924) );
  AND2_X1 U12625 ( .A1(n14062), .A2(n14140), .ZN(n14138) );
  NOR2_X1 U12626 ( .A1(n11310), .A2(n15343), .ZN(n11309) );
  AND2_X1 U12627 ( .A1(n11317), .A2(n10061), .ZN(n11311) );
  AND2_X1 U12628 ( .A1(n12702), .A2(n9932), .ZN(n14062) );
  AND2_X1 U12629 ( .A1(n13707), .A2(n10003), .ZN(n9934) );
  AND2_X1 U12630 ( .A1(n12459), .A2(n12424), .ZN(n16344) );
  INV_X1 U12631 ( .A(n16344), .ZN(n16313) );
  NOR3_X1 U12632 ( .A1(n11306), .A2(n15304), .A3(n10073), .ZN(n11294) );
  AND2_X1 U12633 ( .A1(n10121), .A2(n13349), .ZN(n9935) );
  NAND2_X1 U12634 ( .A1(n13855), .A2(n13878), .ZN(n13879) );
  AND2_X1 U12635 ( .A1(n13851), .A2(n13857), .ZN(n13855) );
  AND2_X1 U12636 ( .A1(n11515), .A2(n10102), .ZN(n13851) );
  OR3_X1 U12637 ( .A1(n12841), .A2(n12840), .A3(n15191), .ZN(n9936) );
  NAND2_X1 U12638 ( .A1(n11515), .A2(n11514), .ZN(n13768) );
  INV_X1 U12639 ( .A(n13953), .ZN(n10115) );
  AND2_X1 U12640 ( .A1(n9935), .A2(n10120), .ZN(n9937) );
  INV_X1 U12641 ( .A(n16342), .ZN(n16327) );
  AND2_X1 U12642 ( .A1(n12459), .A2(n19930), .ZN(n16342) );
  NAND2_X1 U12643 ( .A1(n14221), .A2(n11820), .ZN(n14336) );
  INV_X1 U12644 ( .A(n12207), .ZN(n10080) );
  NAND2_X1 U12645 ( .A1(n11515), .A2(n10104), .ZN(n13767) );
  INV_X1 U12646 ( .A(n13826), .ZN(n10166) );
  NOR2_X1 U12647 ( .A1(n10166), .A2(n10164), .ZN(n13881) );
  OR2_X1 U12648 ( .A1(n14204), .A2(n14205), .ZN(n14257) );
  INV_X1 U12649 ( .A(n14257), .ZN(n9957) );
  INV_X2 U12650 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n20806) );
  NOR2_X1 U12651 ( .A1(n11307), .A2(n15322), .ZN(n11304) );
  AND2_X1 U12652 ( .A1(n10003), .A2(n20773), .ZN(n9938) );
  NAND2_X1 U12653 ( .A1(n12702), .A2(n10169), .ZN(n10168) );
  NAND2_X1 U12654 ( .A1(n12702), .A2(n9918), .ZN(n10167) );
  OR2_X1 U12655 ( .A1(n19256), .A2(n19015), .ZN(n9939) );
  AND2_X1 U12656 ( .A1(n10109), .A2(n10108), .ZN(n9940) );
  AND2_X1 U12657 ( .A1(n10070), .A2(n15357), .ZN(n9941) );
  AND2_X1 U12658 ( .A1(n10071), .A2(n15357), .ZN(n9942) );
  INV_X1 U12659 ( .A(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n10073) );
  INV_X1 U12660 ( .A(n16293), .ZN(n19248) );
  NOR2_X1 U12661 ( .A1(n11306), .A2(n10072), .ZN(n11296) );
  INV_X1 U12662 ( .A(P2_EBX_REG_8__SCAN_IN), .ZN(n10078) );
  NOR2_X1 U12663 ( .A1(n13814), .A2(n13813), .ZN(n9943) );
  INV_X1 U12664 ( .A(n12458), .ZN(n19038) );
  INV_X1 U12665 ( .A(n19297), .ZN(n10156) );
  NAND2_X1 U12666 ( .A1(n14495), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n9944) );
  INV_X1 U12667 ( .A(P2_EBX_REG_24__SCAN_IN), .ZN(n10047) );
  OR2_X1 U12668 ( .A1(n9944), .A2(n10009), .ZN(n9945) );
  OR2_X1 U12669 ( .A1(n15501), .A2(n15300), .ZN(n9946) );
  INV_X1 U12670 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n10012) );
  INV_X1 U12671 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n10009) );
  INV_X1 U12672 ( .A(P2_EBX_REG_20__SCAN_IN), .ZN(n10079) );
  INV_X1 U12673 ( .A(n19389), .ZN(n19747) );
  AOI22_X2 U12674 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n19295), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n19294), .ZN(n19790) );
  AOI22_X2 U12675 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n19295), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n19294), .ZN(n19722) );
  NOR2_X2 U12676 ( .A1(n14030), .A2(n16305), .ZN(n19294) );
  AOI22_X2 U12677 ( .A1(DATAI_22_), .A2(n20161), .B1(BUF1_REG_22__SCAN_IN), 
        .B2(n20196), .ZN(n20682) );
  NOR2_X2 U12678 ( .A1(n18254), .A2(n18276), .ZN(n18569) );
  NOR3_X2 U12679 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18745), .A3(
        n18459), .ZN(n18429) );
  NOR2_X2 U12680 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n18864), .ZN(n18745) );
  AND2_X2 U12681 ( .A1(n13744), .A2(n10292), .ZN(n10335) );
  AND2_X2 U12682 ( .A1(n10581), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13744) );
  INV_X1 U12683 ( .A(n9951), .ZN(n14714) );
  NAND2_X1 U12684 ( .A1(n9954), .A2(n9952), .ZN(n13945) );
  NAND2_X1 U12685 ( .A1(n9955), .A2(n11196), .ZN(n13997) );
  XNOR2_X2 U12686 ( .A(n11268), .B(n11267), .ZN(n14663) );
  NOR2_X2 U12687 ( .A1(n14690), .A2(n14684), .ZN(n14683) );
  NAND2_X1 U12688 ( .A1(n12062), .A2(n11813), .ZN(n12341) );
  NAND2_X1 U12689 ( .A1(n9961), .A2(n12359), .ZN(n12347) );
  OR2_X2 U12690 ( .A1(n15361), .A2(n9907), .ZN(n10229) );
  NAND2_X2 U12691 ( .A1(n15662), .A2(n15661), .ZN(n15361) );
  INV_X1 U12692 ( .A(n14330), .ZN(n9970) );
  NAND3_X1 U12693 ( .A1(n9971), .A2(n9969), .A3(n9931), .ZN(n10213) );
  NAND2_X1 U12694 ( .A1(n12187), .A2(n9970), .ZN(n9969) );
  NAND3_X1 U12695 ( .A1(n12187), .A2(n10081), .A3(n12131), .ZN(n9971) );
  NAND2_X1 U12696 ( .A1(n14329), .A2(n14330), .ZN(n15457) );
  NAND2_X2 U12697 ( .A1(n9973), .A2(n9972), .ZN(n15774) );
  NAND2_X2 U12698 ( .A1(n11638), .A2(n13542), .ZN(n11616) );
  NAND3_X1 U12699 ( .A1(n16249), .A2(n16250), .A3(n9939), .ZN(P2_U3000) );
  NAND3_X1 U12700 ( .A1(n11472), .A2(n9975), .A3(n9974), .ZN(n12420) );
  INV_X2 U12701 ( .A(n11765), .ZN(n11443) );
  INV_X1 U12702 ( .A(n11637), .ZN(n12114) );
  NAND2_X1 U12703 ( .A1(n11765), .A2(n16370), .ZN(n11637) );
  NAND2_X2 U12704 ( .A1(n9978), .A2(n9976), .ZN(n16370) );
  NAND4_X1 U12705 ( .A1(n11416), .A2(n11414), .A3(n11417), .A4(n11415), .ZN(
        n9977) );
  NAND3_X1 U12706 ( .A1(n11413), .A2(n11410), .A3(n11411), .ZN(n9980) );
  AND2_X2 U12707 ( .A1(n11434), .A2(n11433), .ZN(n11765) );
  INV_X1 U12708 ( .A(n12106), .ZN(n9982) );
  NAND3_X1 U12709 ( .A1(n9983), .A2(n12338), .A3(n14100), .ZN(n14102) );
  NAND2_X2 U12710 ( .A1(n12106), .A2(n12105), .ZN(n12338) );
  NAND3_X1 U12711 ( .A1(n9889), .A2(n12356), .A3(n12367), .ZN(n9991) );
  NAND2_X1 U12712 ( .A1(n20205), .A2(n9997), .ZN(n13910) );
  XNOR2_X1 U12713 ( .A(n9998), .B(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14508) );
  NAND2_X1 U12714 ( .A1(n10000), .A2(n10122), .ZN(n9999) );
  NAND2_X1 U12715 ( .A1(n10001), .A2(n14475), .ZN(n14476) );
  OAI21_X1 U12716 ( .B1(n14839), .B2(n14961), .A(n16081), .ZN(n10001) );
  NAND2_X1 U12717 ( .A1(n10003), .A2(n20806), .ZN(n10575) );
  AOI21_X1 U12718 ( .B1(n10003), .B2(n13753), .A(n13752), .ZN(n13895) );
  INV_X1 U12719 ( .A(n10003), .ZN(n10002) );
  AOI22_X1 U12720 ( .A1(n13983), .A2(P1_REIP_REG_3__SCAN_IN), .B1(n20027), 
        .B2(n10003), .ZN(n13984) );
  OAI21_X1 U12721 ( .B1(n10008), .B2(n10007), .A(n9945), .ZN(n10006) );
  NAND2_X1 U12722 ( .A1(n12650), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n10007) );
  NAND2_X1 U12723 ( .A1(n10577), .A2(n10010), .ZN(n10666) );
  NAND3_X1 U12724 ( .A1(n10014), .A2(P3_EAX_REG_9__SCAN_IN), .A3(
        P3_EAX_REG_8__SCAN_IN), .ZN(n10013) );
  INV_X2 U12725 ( .A(n17356), .ZN(n18277) );
  NAND3_X2 U12726 ( .A1(n9898), .A2(n13195), .A3(n9871), .ZN(n17356) );
  NAND2_X1 U12727 ( .A1(n18248), .A2(n17356), .ZN(n13253) );
  NAND3_X1 U12728 ( .A1(n10019), .A2(P3_EAX_REG_19__SCAN_IN), .A3(
        P3_EAX_REG_20__SCAN_IN), .ZN(n10018) );
  INV_X2 U12729 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n18870) );
  OR2_X2 U12731 ( .A1(n10462), .A2(n10461), .ZN(n10028) );
  INV_X1 U12732 ( .A(n10535), .ZN(n10029) );
  OAI211_X2 U12733 ( .C1(n10027), .C2(n10025), .A(n10024), .B(n10022), .ZN(
        n10536) );
  NAND2_X1 U12734 ( .A1(n14163), .A2(n10035), .ZN(n10031) );
  NAND2_X1 U12735 ( .A1(n10031), .A2(n10032), .ZN(n14246) );
  NAND2_X2 U12736 ( .A1(n12649), .A2(n16081), .ZN(n15015) );
  NAND3_X1 U12737 ( .A1(n12650), .A2(n15015), .A3(n10009), .ZN(n14856) );
  INV_X1 U12738 ( .A(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n10045) );
  NAND4_X1 U12739 ( .A1(n10046), .A2(n10044), .A3(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A4(
        P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n11325) );
  NAND3_X1 U12740 ( .A1(n10046), .A2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A3(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n11327) );
  INV_X1 U12741 ( .A(n10054), .ZN(n16217) );
  INV_X1 U12742 ( .A(n12118), .ZN(n10057) );
  NAND3_X1 U12743 ( .A1(n10055), .A2(n12125), .A3(n12108), .ZN(n12167) );
  NAND2_X1 U12744 ( .A1(n11335), .A2(n11314), .ZN(n10064) );
  NAND2_X1 U12745 ( .A1(n10064), .A2(n10063), .ZN(n18941) );
  INV_X1 U12746 ( .A(n10067), .ZN(n18960) );
  INV_X1 U12747 ( .A(n18959), .ZN(n10066) );
  AOI21_X1 U12748 ( .B1(n13345), .B2(n15357), .A(n10053), .ZN(n13358) );
  NAND2_X1 U12749 ( .A1(n10069), .A2(n10068), .ZN(n13357) );
  NAND2_X1 U12750 ( .A1(n13345), .A2(n9941), .ZN(n10069) );
  INV_X1 U12751 ( .A(n10071), .ZN(n15857) );
  NAND3_X1 U12752 ( .A1(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_29__SCAN_IN), .A3(
        P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n10072) );
  NAND2_X1 U12753 ( .A1(n11296), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11298) );
  NAND2_X1 U12754 ( .A1(n12206), .A2(n12207), .ZN(n12225) );
  NAND2_X1 U12755 ( .A1(n14216), .A2(n14215), .ZN(n10081) );
  OR2_X2 U12756 ( .A1(n10082), .A2(n11972), .ZN(n11976) );
  NAND2_X1 U12757 ( .A1(n10082), .A2(n11969), .ZN(n11492) );
  NAND3_X1 U12758 ( .A1(n10082), .A2(n11973), .A3(n11974), .ZN(n11975) );
  OAI21_X1 U12759 ( .B1(n10082), .B2(n11969), .A(n11968), .ZN(n11493) );
  XNOR2_X2 U12760 ( .A(n11986), .B(n10082), .ZN(n12684) );
  NAND2_X2 U12761 ( .A1(n10101), .A2(n10100), .ZN(n10082) );
  NAND2_X4 U12762 ( .A1(n10084), .A2(n10083), .ZN(n11451) );
  NAND2_X1 U12763 ( .A1(n10086), .A2(n11651), .ZN(n10083) );
  NAND2_X1 U12764 ( .A1(n10085), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10084) );
  NAND4_X1 U12765 ( .A1(n11405), .A2(n10277), .A3(n11403), .A4(n11404), .ZN(
        n10085) );
  NAND4_X1 U12766 ( .A1(n11409), .A2(n11408), .A3(n11406), .A4(n11407), .ZN(
        n10086) );
  AND2_X2 U12767 ( .A1(n10087), .A2(n13584), .ZN(n12021) );
  NAND2_X1 U12768 ( .A1(n10213), .A2(n10090), .ZN(n10088) );
  NAND2_X1 U12769 ( .A1(n10096), .A2(n11460), .ZN(n11463) );
  NAND2_X1 U12770 ( .A1(n10097), .A2(n11456), .ZN(n10096) );
  NAND2_X1 U12771 ( .A1(n11458), .A2(n10098), .ZN(n10097) );
  INV_X1 U12772 ( .A(n11457), .ZN(n10098) );
  NOR2_X2 U12773 ( .A1(n11456), .A2(n19297), .ZN(n12439) );
  NAND2_X2 U12774 ( .A1(n11398), .A2(n11399), .ZN(n19290) );
  NAND2_X1 U12775 ( .A1(n11484), .A2(n11483), .ZN(n10100) );
  XNOR2_X2 U12776 ( .A(n11483), .B(n11482), .ZN(n11981) );
  NAND2_X1 U12777 ( .A1(n11558), .A2(n10105), .ZN(n14322) );
  NAND2_X1 U12778 ( .A1(n13335), .A2(n10109), .ZN(n12508) );
  NAND2_X1 U12779 ( .A1(n13335), .A2(n12297), .ZN(n12296) );
  NAND2_X1 U12780 ( .A1(n10551), .A2(n10135), .ZN(n10132) );
  NAND3_X1 U12781 ( .A1(n10134), .A2(n10136), .A3(n10132), .ZN(n12574) );
  NAND3_X1 U12782 ( .A1(n10134), .A2(n10133), .A3(n10132), .ZN(n10139) );
  OAI21_X1 U12783 ( .B1(n10142), .B2(n14891), .A(n10145), .ZN(n16051) );
  NAND2_X1 U12784 ( .A1(n14891), .A2(n10145), .ZN(n10143) );
  NAND2_X1 U12785 ( .A1(n10152), .A2(n10150), .ZN(n12442) );
  NAND3_X1 U12786 ( .A1(n10151), .A2(n11419), .A3(n10156), .ZN(n10150) );
  NAND4_X1 U12787 ( .A1(n10154), .A2(n11456), .A3(n12379), .A4(n10153), .ZN(
        n10152) );
  INV_X1 U12788 ( .A(n11794), .ZN(n10155) );
  NOR2_X1 U12789 ( .A1(n10157), .A2(n12374), .ZN(n12428) );
  INV_X1 U12790 ( .A(n11979), .ZN(n10159) );
  INV_X1 U12791 ( .A(n11980), .ZN(n10160) );
  NAND3_X1 U12792 ( .A1(n10162), .A2(n11982), .A3(n12676), .ZN(n10158) );
  NAND2_X1 U12793 ( .A1(n13826), .A2(n10163), .ZN(n13882) );
  NAND2_X1 U12794 ( .A1(n13826), .A2(n9879), .ZN(n13848) );
  INV_X1 U12795 ( .A(n12819), .ZN(n10170) );
  NAND2_X1 U12796 ( .A1(n10170), .A2(n9936), .ZN(n10172) );
  NOR2_X1 U12797 ( .A1(n13862), .A2(n13861), .ZN(n13863) );
  NAND2_X1 U12798 ( .A1(n15632), .A2(n9933), .ZN(n15596) );
  NAND2_X1 U12799 ( .A1(n15726), .A2(n9910), .ZN(n15689) );
  NOR2_X2 U12800 ( .A1(n15573), .A2(n10184), .ZN(n15550) );
  NAND3_X1 U12801 ( .A1(n13350), .A2(n15548), .A3(n11943), .ZN(n10184) );
  NAND2_X1 U12802 ( .A1(n15550), .A2(n13363), .ZN(n13362) );
  INV_X1 U12803 ( .A(n13350), .ZN(n10185) );
  NOR2_X2 U12804 ( .A1(n15129), .A2(n15115), .ZN(n15252) );
  NAND2_X1 U12805 ( .A1(n10188), .A2(n13700), .ZN(n13699) );
  OAI21_X1 U12806 ( .B1(n13700), .B2(n10188), .A(n13699), .ZN(n13958) );
  NAND3_X1 U12807 ( .A1(n13876), .A2(n10614), .A3(n13875), .ZN(n13941) );
  INV_X1 U12808 ( .A(n13941), .ZN(n10642) );
  NAND2_X1 U12809 ( .A1(n10551), .A2(n10191), .ZN(n10190) );
  AND2_X2 U12810 ( .A1(n10290), .A2(n10291), .ZN(n11078) );
  INV_X1 U12811 ( .A(n14721), .ZN(n10193) );
  NAND2_X1 U12812 ( .A1(n10193), .A2(n10194), .ZN(n14606) );
  NAND2_X1 U12813 ( .A1(n14254), .A2(n14300), .ZN(n14299) );
  OR2_X1 U12814 ( .A1(n14300), .A2(n14304), .ZN(n10206) );
  OR2_X2 U12815 ( .A1(n10351), .A2(n10352), .ZN(n12571) );
  NAND2_X1 U12816 ( .A1(n12655), .A2(n10207), .ZN(n10210) );
  AND2_X4 U12817 ( .A1(n15743), .A2(n15754), .ZN(n12797) );
  NAND2_X1 U12818 ( .A1(n17878), .A2(n18190), .ZN(n17879) );
  NAND2_X2 U12819 ( .A1(n17889), .A2(n13111), .ZN(n13113) );
  NAND2_X1 U12820 ( .A1(n17890), .A2(n17891), .ZN(n17889) );
  NOR2_X2 U12821 ( .A1(n13133), .A2(n9870), .ZN(n17809) );
  NOR2_X2 U12822 ( .A1(n13279), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13133) );
  NAND2_X1 U12823 ( .A1(n13104), .A2(n10216), .ZN(n17898) );
  INV_X1 U12824 ( .A(n17421), .ZN(n13108) );
  NAND2_X1 U12825 ( .A1(n13072), .A2(n9908), .ZN(n10219) );
  NOR2_X2 U12826 ( .A1(n13140), .A2(n17650), .ZN(n17687) );
  NAND3_X1 U12827 ( .A1(n10229), .A2(n10231), .A3(n10227), .ZN(n15330) );
  NAND4_X1 U12828 ( .A1(n10229), .A2(n10231), .A3(n10227), .A4(
        P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n10237) );
  NAND2_X1 U12829 ( .A1(n10230), .A2(n15351), .ZN(n15342) );
  OAI21_X1 U12830 ( .B1(n15361), .B2(n12246), .A(n10234), .ZN(n10230) );
  NAND2_X1 U12831 ( .A1(n10237), .A2(n12259), .ZN(n12261) );
  NOR2_X2 U12832 ( .A1(n17561), .A2(n17757), .ZN(n16447) );
  AOI21_X1 U12833 ( .B1(n17754), .B2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n10242), .ZN(n10241) );
  INV_X1 U12834 ( .A(n17705), .ZN(n13138) );
  NAND2_X1 U12835 ( .A1(n11981), .A2(n19098), .ZN(n12013) );
  NAND2_X2 U12836 ( .A1(n12062), .A2(n10245), .ZN(n12359) );
  XNOR2_X2 U12837 ( .A(n12359), .B(n12165), .ZN(n12350) );
  NAND2_X1 U12838 ( .A1(n12442), .A2(n16370), .ZN(n11450) );
  INV_X1 U12839 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10246) );
  NOR2_X2 U12840 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n15758) );
  NAND2_X1 U12841 ( .A1(n14220), .A2(n10248), .ZN(n10250) );
  NAND3_X1 U12842 ( .A1(n12353), .A2(n12354), .A3(n10250), .ZN(n14328) );
  NAND2_X1 U12843 ( .A1(n14220), .A2(n12351), .ZN(n10251) );
  NAND2_X1 U12844 ( .A1(n10251), .A2(n12350), .ZN(n12356) );
  AND2_X1 U12845 ( .A1(n15674), .A2(n12455), .ZN(n15398) );
  INV_X1 U12846 ( .A(n15311), .ZN(n10255) );
  NOR2_X1 U12847 ( .A1(n15311), .A2(n10257), .ZN(n12506) );
  NAND2_X1 U12848 ( .A1(n10255), .A2(n10256), .ZN(n12373) );
  NOR2_X1 U12849 ( .A1(n15311), .A2(n15501), .ZN(n15299) );
  OR2_X2 U12850 ( .A1(n15311), .A2(n9946), .ZN(n12372) );
  NAND2_X1 U12851 ( .A1(n15295), .A2(n16338), .ZN(n12498) );
  AOI21_X1 U12852 ( .B1(n15156), .B2(n19250), .A(n12992), .ZN(n12993) );
  NAND2_X1 U12853 ( .A1(n15156), .A2(n19097), .ZN(n11764) );
  NOR2_X1 U12854 ( .A1(n20772), .A2(n20408), .ZN(n20776) );
  NAND2_X1 U12855 ( .A1(n20772), .A2(n13917), .ZN(n20263) );
  NAND2_X1 U12856 ( .A1(n12650), .A2(n9913), .ZN(n12651) );
  INV_X1 U12857 ( .A(n12454), .ZN(n15156) );
  NAND2_X1 U12858 ( .A1(n12531), .A2(n19248), .ZN(n12515) );
  NOR3_X1 U12859 ( .A1(n10474), .A2(n11112), .A3(n10417), .ZN(n10354) );
  NAND2_X1 U12860 ( .A1(n15172), .A2(n15171), .ZN(n15170) );
  CLKBUF_X1 U12861 ( .A(n11963), .Z(n16390) );
  AOI22_X1 U12862 ( .A1(n11427), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n9856), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11370) );
  NAND2_X1 U12863 ( .A1(n14102), .A2(n12337), .ZN(n12342) );
  AND2_X1 U12864 ( .A1(n12901), .A2(n12900), .ZN(n12902) );
  INV_X1 U12865 ( .A(n19290), .ZN(n11452) );
  INV_X1 U12866 ( .A(n11985), .ZN(n11969) );
  OR2_X1 U12867 ( .A1(n12359), .A2(n12358), .ZN(n12363) );
  AOI22_X1 U12868 ( .A1(n12797), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11427), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11417) );
  AOI22_X1 U12869 ( .A1(n9845), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12828), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11403) );
  AOI22_X1 U12870 ( .A1(n11646), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11645), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11369) );
  AOI22_X1 U12871 ( .A1(n11646), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n11645), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11351) );
  NAND2_X1 U12872 ( .A1(n14506), .A2(n12541), .ZN(n12559) );
  NOR2_X1 U12873 ( .A1(n15179), .A2(n15178), .ZN(n15177) );
  OAI22_X1 U12874 ( .A1(n19452), .A2(n12033), .B1(n14124), .B2(n12032), .ZN(
        n12034) );
  INV_X1 U12875 ( .A(n10542), .ZN(n10544) );
  INV_X1 U12876 ( .A(n19067), .ZN(n19097) );
  AND2_X1 U12877 ( .A1(n20043), .A2(n13619), .ZN(n20040) );
  OR2_X1 U12879 ( .A1(n19415), .A2(n11991), .ZN(n10260) );
  INV_X1 U12880 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n13107) );
  AND3_X1 U12881 ( .A1(n12499), .A2(n12498), .A3(n9909), .ZN(n10261) );
  AND3_X1 U12882 ( .A1(n12011), .A2(n12010), .A3(n12009), .ZN(n10262) );
  NOR2_X1 U12883 ( .A1(n20493), .A2(n20783), .ZN(n10263) );
  AND2_X1 U12884 ( .A1(n11190), .A2(n11189), .ZN(n10265) );
  AND2_X1 U12885 ( .A1(n12987), .A2(n12986), .ZN(n10266) );
  OR2_X1 U12886 ( .A1(n11451), .A2(n13629), .ZN(n10267) );
  AND2_X1 U12887 ( .A1(n12881), .A2(n10278), .ZN(n10268) );
  INV_X1 U12888 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n14633) );
  AND2_X1 U12889 ( .A1(n10540), .A2(n10539), .ZN(n10269) );
  AND3_X1 U12890 ( .A1(n14499), .A2(n14503), .A3(n14498), .ZN(n10270) );
  INV_X1 U12891 ( .A(n14394), .ZN(n17267) );
  INV_X1 U12892 ( .A(n17267), .ZN(n17260) );
  INV_X1 U12893 ( .A(n14749), .ZN(n14719) );
  AND2_X1 U12894 ( .A1(n11610), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n10271) );
  AND2_X1 U12895 ( .A1(n14748), .A2(n14519), .ZN(n14378) );
  AND4_X1 U12896 ( .A1(n13062), .A2(n13061), .A3(n13060), .A4(n13059), .ZN(
        n10272) );
  INV_X1 U12897 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n13112) );
  OR2_X1 U12898 ( .A1(n14893), .A2(n12642), .ZN(n10273) );
  NOR2_X1 U12899 ( .A1(n13150), .A2(n13146), .ZN(n10274) );
  NOR2_X1 U12900 ( .A1(n20493), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n10275) );
  INV_X1 U12901 ( .A(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n20152) );
  OR2_X1 U12902 ( .A1(n12529), .A2(n12528), .ZN(n10276) );
  AND2_X1 U12903 ( .A1(n11402), .A2(n11401), .ZN(n10277) );
  NAND2_X1 U12904 ( .A1(n17630), .A2(n17910), .ZN(n17697) );
  AND3_X1 U12905 ( .A1(n12896), .A2(n12897), .A3(n12878), .ZN(n10278) );
  INV_X1 U12906 ( .A(n13427), .ZN(n12058) );
  INV_X1 U12907 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n13132) );
  AND2_X1 U12908 ( .A1(n12701), .A2(n13921), .ZN(n10279) );
  INV_X1 U12909 ( .A(n14209), .ZN(n12705) );
  OR2_X1 U12910 ( .A1(n11930), .A2(n11929), .ZN(n14209) );
  AND2_X1 U12911 ( .A1(n12503), .A2(n12500), .ZN(n10280) );
  AND2_X1 U12912 ( .A1(n10725), .A2(n10724), .ZN(n10281) );
  INV_X1 U12913 ( .A(n14072), .ZN(n14202) );
  INV_X1 U12914 ( .A(n10552), .ZN(n10639) );
  INV_X2 U12915 ( .A(n10639), .ZN(n11049) );
  INV_X1 U12916 ( .A(n14380), .ZN(n15227) );
  AND2_X1 U12917 ( .A1(n11998), .A2(n12684), .ZN(n10282) );
  INV_X1 U12918 ( .A(n15375), .ZN(n15387) );
  OAI22_X1 U12919 ( .A1(n12085), .A2(n11996), .B1(n19304), .B2(n11995), .ZN(
        n11997) );
  INV_X1 U12920 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10283) );
  INV_X1 U12921 ( .A(n10629), .ZN(n10630) );
  AND3_X1 U12922 ( .A1(n10447), .A2(n10446), .A3(n10445), .ZN(n10448) );
  NAND2_X1 U12923 ( .A1(n10429), .A2(n10527), .ZN(n10430) );
  AND2_X1 U12924 ( .A1(n19297), .A2(n19281), .ZN(n11458) );
  INV_X1 U12925 ( .A(n11114), .ZN(n11119) );
  OR2_X1 U12926 ( .A1(n10624), .A2(n10623), .ZN(n12614) );
  INV_X1 U12927 ( .A(n10667), .ZN(n10668) );
  INV_X1 U12928 ( .A(n10666), .ZN(n10669) );
  AND2_X1 U12929 ( .A1(n11147), .A2(n11166), .ZN(n11148) );
  AOI22_X1 U12930 ( .A1(n11646), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n9850), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11406) );
  INV_X1 U12931 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11339) );
  AOI22_X1 U12932 ( .A1(n11427), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__2__SCAN_IN), .B2(n12798), .ZN(n11347) );
  AOI22_X1 U12933 ( .A1(n11427), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n12929), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11359) );
  AOI22_X1 U12934 ( .A1(n12797), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n11427), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11379) );
  AND2_X1 U12935 ( .A1(n11154), .A2(n11152), .ZN(n11166) );
  INV_X1 U12936 ( .A(n14696), .ZN(n10905) );
  INV_X1 U12937 ( .A(n14729), .ZN(n10803) );
  INV_X1 U12938 ( .A(n14201), .ZN(n10705) );
  INV_X1 U12939 ( .A(n13942), .ZN(n10641) );
  INV_X1 U12940 ( .A(n10475), .ZN(n12585) );
  NOR2_X1 U12941 ( .A1(n10523), .A2(n20806), .ZN(n12631) );
  AOI22_X1 U12942 ( .A1(n10335), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n10597), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10294) );
  INV_X1 U12943 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n11293) );
  AND2_X1 U12944 ( .A1(n15205), .A2(n12818), .ZN(n12819) );
  OR2_X1 U12945 ( .A1(n12489), .A2(n15291), .ZN(n12490) );
  AND4_X1 U12946 ( .A1(n11741), .A2(n11740), .A3(n11739), .A4(n11738), .ZN(
        n11743) );
  INV_X1 U12947 ( .A(n11441), .ZN(n12432) );
  AND2_X1 U12948 ( .A1(n12684), .A2(n11998), .ZN(n11994) );
  AOI21_X1 U12949 ( .B1(n11154), .B2(n11153), .A(n11152), .ZN(n13492) );
  INV_X1 U12950 ( .A(n11034), .ZN(n11035) );
  INV_X1 U12951 ( .A(n10968), .ZN(n10969) );
  AND2_X1 U12952 ( .A1(n10654), .A2(n10653), .ZN(n10667) );
  NAND2_X1 U12953 ( .A1(n10605), .A2(n10604), .ZN(n10631) );
  OR2_X1 U12954 ( .A1(n16081), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n12638) );
  NAND2_X1 U12955 ( .A1(n11147), .A2(n12630), .ZN(n11156) );
  OR2_X1 U12956 ( .A1(n11632), .A2(n11624), .ZN(n11626) );
  INV_X1 U12957 ( .A(n13951), .ZN(n12703) );
  INV_X1 U12958 ( .A(n13769), .ZN(n11521) );
  AOI21_X1 U12959 ( .B1(n15237), .B2(n16344), .A(n12490), .ZN(n12491) );
  OR2_X1 U12960 ( .A1(n15599), .A2(n15414), .ZN(n15587) );
  NOR2_X1 U12961 ( .A1(n11674), .A2(n11673), .ZN(n12330) );
  AND2_X1 U12962 ( .A1(n12684), .A2(n12012), .ZN(n12004) );
  NAND2_X1 U12963 ( .A1(n12319), .A2(n12318), .ZN(n12320) );
  AND2_X1 U12964 ( .A1(n13268), .A2(n13267), .ZN(n13168) );
  INV_X1 U12965 ( .A(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n21055) );
  INV_X1 U12966 ( .A(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n21120) );
  NAND2_X1 U12967 ( .A1(n13116), .A2(n13293), .ZN(n13096) );
  NOR2_X1 U12968 ( .A1(n17275), .A2(n18271), .ZN(n13277) );
  INV_X1 U12969 ( .A(n18258), .ZN(n13262) );
  AND2_X1 U12970 ( .A1(n11204), .A2(n11203), .ZN(n13991) );
  OR2_X1 U12971 ( .A1(n15901), .A2(n13726), .ZN(n13806) );
  INV_X1 U12972 ( .A(n13392), .ZN(n13373) );
  AND2_X1 U12973 ( .A1(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n10969), .ZN(
        n10970) );
  OAI211_X1 U12974 ( .C1(n10675), .C2(n10609), .A(n10674), .B(n10673), .ZN(
        n13988) );
  AND2_X1 U12975 ( .A1(n20802), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n12658) );
  OR3_X1 U12976 ( .A1(n13735), .A2(n13734), .A3(n13733), .ZN(n13901) );
  OR2_X1 U12977 ( .A1(n11861), .A2(n11860), .ZN(n12701) );
  INV_X1 U12978 ( .A(n12861), .ZN(n12858) );
  AND2_X1 U12979 ( .A1(n13529), .A2(n13528), .ZN(n19165) );
  AND2_X1 U12980 ( .A1(n11520), .A2(n11519), .ZN(n13769) );
  AND2_X1 U12981 ( .A1(n15510), .A2(n12474), .ZN(n15474) );
  NAND2_X1 U12982 ( .A1(n17490), .A2(n16589), .ZN(n15804) );
  NOR2_X1 U12983 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n16867), .ZN(n16840) );
  INV_X1 U12984 ( .A(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n21007) );
  INV_X1 U12985 ( .A(n17670), .ZN(n16730) );
  NOR2_X1 U12986 ( .A1(n18018), .A2(n17705), .ZN(n17650) );
  NAND2_X1 U12987 ( .A1(n13134), .A2(n17757), .ZN(n17756) );
  NOR2_X1 U12988 ( .A1(n17818), .A2(n13279), .ZN(n17775) );
  NOR2_X1 U12989 ( .A1(n13298), .A2(n17847), .ZN(n13301) );
  INV_X1 U12990 ( .A(n17405), .ZN(n13293) );
  NAND3_X1 U12991 ( .A1(n13228), .A2(n13227), .A3(n13226), .ZN(n13273) );
  AND2_X1 U12992 ( .A1(n15950), .A2(P1_REIP_REG_23__SCAN_IN), .ZN(n15935) );
  AND2_X1 U12993 ( .A1(n11235), .A2(n11234), .ZN(n14712) );
  INV_X1 U12994 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n14648) );
  INV_X1 U12995 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n14080) );
  NAND2_X1 U12996 ( .A1(n10561), .A2(n10560), .ZN(n20292) );
  OR3_X1 U12997 ( .A1(n11282), .A2(n11281), .A3(n11280), .ZN(n19997) );
  NOR2_X2 U12998 ( .A1(n14642), .A2(n14375), .ZN(n14733) );
  XNOR2_X1 U12999 ( .A(n11173), .B(n11283), .ZN(n14504) );
  AND2_X1 U13000 ( .A1(n11015), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n11034) );
  INV_X1 U13001 ( .A(n14694), .ZN(n14707) );
  AOI21_X1 U13002 ( .B1(n12613), .B2(n10671), .A(n10661), .ZN(n14000) );
  AND2_X1 U13003 ( .A1(n12658), .A2(n20413), .ZN(n20775) );
  AND3_X1 U13004 ( .A1(n11192), .A2(n11243), .A3(n11191), .ZN(n13944) );
  INV_X1 U13005 ( .A(n20232), .ZN(n20467) );
  NAND2_X1 U13006 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n20297), .ZN(n20195) );
  INV_X1 U13007 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n13782) );
  INV_X1 U13008 ( .A(n11760), .ZN(n11761) );
  INV_X1 U13009 ( .A(n11644), .ZN(n11762) );
  XNOR2_X1 U13010 ( .A(n11298), .B(n11297), .ZN(n12991) );
  INV_X1 U13011 ( .A(n12403), .ZN(n12276) );
  OR3_X1 U13012 ( .A1(n18953), .A2(n12417), .A3(n15401), .ZN(n15393) );
  XNOR2_X1 U13013 ( .A(n12365), .B(n12364), .ZN(n16288) );
  INV_X1 U13014 ( .A(n12684), .ZN(n11987) );
  INV_X1 U13015 ( .A(n19910), .ZN(n14023) );
  NAND2_X1 U13016 ( .A1(n19539), .A2(n19921), .ZN(n19476) );
  AND2_X1 U13017 ( .A1(n16399), .A2(n19915), .ZN(n12321) );
  OR2_X1 U13018 ( .A1(n19901), .A2(n14023), .ZN(n19658) );
  OR2_X1 U13019 ( .A1(n19539), .A2(n19921), .ZN(n19689) );
  INV_X1 U13020 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n19802) );
  OR2_X1 U13021 ( .A1(n16687), .A2(n16765), .ZN(n16724) );
  INV_X1 U13022 ( .A(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n16816) );
  INV_X1 U13023 ( .A(n16939), .ZN(n16946) );
  INV_X1 U13024 ( .A(n18267), .ZN(n17275) );
  OAI21_X1 U13025 ( .B1(n17904), .B2(n17697), .A(n18343), .ZN(n17712) );
  INV_X1 U13026 ( .A(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n17751) );
  INV_X1 U13027 ( .A(n17805), .ZN(n17783) );
  OAI21_X1 U13028 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n18883), .A(n16560), 
        .ZN(n17910) );
  INV_X1 U13029 ( .A(n17818), .ZN(n17757) );
  NOR2_X1 U13030 ( .A1(n18059), .A2(n17738), .ZN(n18048) );
  NOR2_X1 U13031 ( .A1(n18710), .A2(n18699), .ZN(n18118) );
  NOR2_X1 U13032 ( .A1(n18163), .A2(n17839), .ZN(n17838) );
  NOR2_X1 U13033 ( .A1(n13207), .A2(n13206), .ZN(n18258) );
  AOI22_X1 U13034 ( .A1(n18682), .A2(n18681), .B1(n18686), .B2(n16454), .ZN(
        n18690) );
  AND2_X1 U13035 ( .A1(n15901), .A2(n13736), .ZN(n13418) );
  AND2_X1 U13036 ( .A1(n15897), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n13736) );
  NOR2_X1 U13037 ( .A1(n19999), .A2(n11284), .ZN(n19970) );
  INV_X1 U13038 ( .A(n19997), .ZN(n20025) );
  AND2_X1 U13039 ( .A1(n13812), .A2(n13811), .ZN(n14718) );
  NAND2_X1 U13040 ( .A1(n13734), .A2(n13736), .ZN(n12540) );
  INV_X1 U13041 ( .A(n20043), .ZN(n14816) );
  INV_X1 U13042 ( .A(n13603), .ZN(n20082) );
  NAND2_X1 U13043 ( .A1(n10907), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n10968) );
  NAND2_X1 U13044 ( .A1(n10838), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n10871) );
  NAND2_X1 U13045 ( .A1(n10635), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10655) );
  INV_X1 U13046 ( .A(n13699), .ZN(n13764) );
  NOR2_X1 U13047 ( .A1(n16152), .A2(n14490), .ZN(n16140) );
  NAND2_X1 U13048 ( .A1(n13381), .A2(n13736), .ZN(n14165) );
  INV_X1 U13049 ( .A(n20119), .ZN(n20107) );
  INV_X1 U13050 ( .A(n16177), .ZN(n20137) );
  INV_X1 U13051 ( .A(n20121), .ZN(n15051) );
  OAI221_X2 U13052 ( .B1(n20807), .B2(n15078), .C1(n16208), .C2(n15078), .A(
        n20806), .ZN(n20198) );
  NOR2_X1 U13053 ( .A1(n13723), .A2(n20413), .ZN(n15078) );
  OAI22_X1 U13054 ( .A1(n20165), .A2(n20164), .B1(n20469), .B2(n20293), .ZN(
        n20200) );
  INV_X1 U13055 ( .A(n20231), .ZN(n20221) );
  INV_X1 U13056 ( .A(n20260), .ZN(n20252) );
  INV_X1 U13057 ( .A(n20286), .ZN(n20287) );
  INV_X1 U13058 ( .A(n20319), .ZN(n20311) );
  INV_X1 U13059 ( .A(n20335), .ZN(n20344) );
  AND2_X1 U13060 ( .A1(n20320), .A2(n20562), .ZN(n20369) );
  OAI211_X1 U13061 ( .C1(n20429), .C2(n20413), .A(n20467), .B(n20412), .ZN(
        n20430) );
  INV_X1 U13062 ( .A(n20460), .ZN(n20446) );
  OAI22_X1 U13063 ( .A1(n20471), .A2(n20470), .B1(n20469), .B2(n20592), .ZN(
        n20488) );
  INV_X1 U13064 ( .A(n20513), .ZN(n20519) );
  AND2_X1 U13065 ( .A1(n9866), .A2(n20562), .ZN(n20501) );
  AND2_X1 U13066 ( .A1(n20563), .A2(n12574), .ZN(n20587) );
  INV_X1 U13067 ( .A(n20594), .ZN(n20625) );
  AND2_X1 U13068 ( .A1(n16373), .A2(n19808), .ZN(n11964) );
  NOR2_X1 U13069 ( .A1(n11762), .A2(n11761), .ZN(n11763) );
  NAND2_X1 U13070 ( .A1(n12527), .A2(n19097), .ZN(n13004) );
  NAND2_X1 U13071 ( .A1(n13433), .A2(n11643), .ZN(n19074) );
  INV_X1 U13072 ( .A(n19074), .ZN(n19091) );
  AND2_X1 U13073 ( .A1(n13437), .A2(n11640), .ZN(n19090) );
  AND2_X1 U13074 ( .A1(n19241), .A2(n16388), .ZN(n19088) );
  OR2_X1 U13075 ( .A1(n11916), .A2(n11915), .ZN(n14140) );
  OR2_X1 U13076 ( .A1(n11875), .A2(n11874), .ZN(n13951) );
  AND2_X1 U13077 ( .A1(n13838), .A2(n13839), .ZN(n13840) );
  AND2_X1 U13078 ( .A1(n13574), .A2(n14029), .ZN(n19109) );
  INV_X1 U13079 ( .A(n15285), .ZN(n19156) );
  INV_X1 U13080 ( .A(n13500), .ZN(n19242) );
  AND2_X1 U13081 ( .A1(n13438), .A2(n19166), .ZN(n19237) );
  AND2_X1 U13082 ( .A1(n16310), .A2(n15464), .ZN(n16302) );
  INV_X1 U13083 ( .A(n16305), .ZN(n19250) );
  AND2_X1 U13084 ( .A1(n14188), .A2(n14187), .ZN(n19135) );
  AND2_X1 U13085 ( .A1(n12459), .A2(n16366), .ZN(n15610) );
  OAI21_X1 U13086 ( .B1(n19267), .B2(n19266), .A(n19265), .ZN(n19300) );
  NAND2_X1 U13087 ( .A1(n19901), .A2(n19910), .ZN(n19540) );
  NOR2_X2 U13088 ( .A1(n19540), .A2(n19476), .ZN(n19349) );
  INV_X1 U13089 ( .A(n19373), .ZN(n19379) );
  NOR2_X1 U13090 ( .A1(n19388), .A2(n19386), .ZN(n19409) );
  NOR2_X1 U13091 ( .A1(n19476), .A2(n19658), .ZN(n19472) );
  NOR2_X1 U13092 ( .A1(n19688), .A2(n19447), .ZN(n19498) );
  OAI21_X1 U13093 ( .B1(n19514), .B2(n19513), .A(n19512), .ZN(n19532) );
  NOR2_X1 U13094 ( .A1(n19689), .A2(n19540), .ZN(n19553) );
  AND2_X1 U13095 ( .A1(n19611), .A2(n19609), .ZN(n19631) );
  INV_X1 U13096 ( .A(n19758), .ZN(n19704) );
  NOR2_X1 U13097 ( .A1(n19659), .A2(n19658), .ZN(n19718) );
  INV_X1 U13098 ( .A(n19734), .ZN(n19795) );
  AND3_X1 U13099 ( .A1(n21058), .A2(n19873), .A3(n19824), .ZN(n19818) );
  NOR2_X1 U13100 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n16650), .ZN(n16640) );
  NOR2_X1 U13101 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n16702), .ZN(n16688) );
  NOR2_X1 U13102 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n16719), .ZN(n16707) );
  NOR2_X1 U13103 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n16766), .ZN(n16754) );
  NAND2_X1 U13104 ( .A1(n17710), .A2(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n16762) );
  INV_X1 U13105 ( .A(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n16836) );
  INV_X1 U13106 ( .A(n18750), .ZN(n16882) );
  INV_X1 U13107 ( .A(P3_EBX_REG_3__SCAN_IN), .ZN(n17252) );
  NOR2_X1 U13108 ( .A1(n17356), .A2(n17076), .ZN(n17064) );
  NAND2_X1 U13109 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n17120), .ZN(n17090) );
  INV_X1 U13110 ( .A(n17173), .ZN(n17161) );
  NAND4_X1 U13111 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(P3_EBX_REG_3__SCAN_IN), 
        .A3(n14395), .A4(n17248), .ZN(n17247) );
  NAND3_X1 U13112 ( .A1(n14393), .A2(n17428), .A3(n15919), .ZN(n17266) );
  INV_X1 U13113 ( .A(n17415), .ZN(n17422) );
  INV_X1 U13114 ( .A(n18248), .ZN(n17428) );
  NOR2_X1 U13115 ( .A1(n18103), .A2(n18024), .ZN(n18058) );
  OAI22_X1 U13116 ( .A1(n18103), .A2(n17914), .B1(n17822), .B2(n18101), .ZN(
        n17805) );
  NAND2_X1 U13117 ( .A1(n17750), .A2(n17697), .ZN(n17903) );
  NAND2_X1 U13118 ( .A1(n17836), .A2(n17837), .ZN(n17835) );
  INV_X1 U13119 ( .A(n18532), .ZN(n18342) );
  NOR2_X1 U13120 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18864), .ZN(
        n18866) );
  INV_X1 U13121 ( .A(n18517), .ZN(n18523) );
  INV_X1 U13122 ( .A(P3_STATE_REG_1__SCAN_IN), .ZN(n18759) );
  NAND2_X1 U13123 ( .A1(n13418), .A2(n10386), .ZN(n14550) );
  INV_X1 U13124 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n20208) );
  INV_X1 U13125 ( .A(n20026), .ZN(n20014) );
  NAND2_X1 U13126 ( .A1(n20022), .A2(n11174), .ZN(n16023) );
  OR3_X1 U13127 ( .A1(n11282), .A2(n15890), .A3(n11278), .ZN(n20038) );
  NOR2_X1 U13128 ( .A1(n12557), .A2(n12556), .ZN(n12558) );
  INV_X1 U13129 ( .A(n16001), .ZN(n14811) );
  INV_X1 U13130 ( .A(n20047), .ZN(n20073) );
  NOR2_X1 U13131 ( .A1(n14550), .A2(n13587), .ZN(n13657) );
  INV_X1 U13132 ( .A(n16077), .ZN(n20102) );
  OR2_X1 U13133 ( .A1(n12660), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20128) );
  OR2_X1 U13134 ( .A1(n14165), .A2(n13388), .ZN(n16177) );
  INV_X1 U13135 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20790) );
  INV_X1 U13136 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20523) );
  AOI211_X1 U13137 ( .C1(P1_STATE2_REG_2__SCAN_IN), .C2(n20293), .A(n20232), 
        .B(n20156), .ZN(n20183) );
  OR2_X1 U13138 ( .A1(n20204), .A2(n20562), .ZN(n20231) );
  OR2_X1 U13139 ( .A1(n20204), .A2(n12574), .ZN(n20260) );
  OR2_X1 U13140 ( .A1(n20263), .A2(n20348), .ZN(n20286) );
  OR2_X1 U13141 ( .A1(n20263), .A2(n20261), .ZN(n20319) );
  INV_X1 U13142 ( .A(n20402), .ZN(n20372) );
  NAND2_X1 U13143 ( .A1(n20383), .A2(n20501), .ZN(n20433) );
  INV_X1 U13144 ( .A(n20484), .ZN(n20492) );
  NAND2_X1 U13145 ( .A1(n20776), .A2(n20501), .ZN(n20561) );
  NAND2_X1 U13146 ( .A1(n20637), .A2(n12574), .ZN(n20692) );
  INV_X1 U13147 ( .A(n20770), .ZN(n20766) );
  INV_X1 U13148 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n21058) );
  NAND2_X1 U13149 ( .A1(n12453), .A2(n19088), .ZN(n11965) );
  OR2_X1 U13150 ( .A1(n11758), .A2(n11756), .ZN(n19067) );
  AND2_X1 U13151 ( .A1(n12969), .A2(n19808), .ZN(n19140) );
  NAND2_X1 U13152 ( .A1(n19140), .A2(n10155), .ZN(n19160) );
  OR2_X1 U13153 ( .A1(n19236), .A2(n19170), .ZN(n19202) );
  NAND2_X1 U13154 ( .A1(n19168), .A2(n19818), .ZN(n19236) );
  INV_X1 U13155 ( .A(n19241), .ZN(n19166) );
  OR2_X1 U13156 ( .A1(n18916), .A2(n12058), .ZN(n16293) );
  INV_X1 U13157 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n16266) );
  INV_X1 U13158 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n16278) );
  NAND2_X1 U13159 ( .A1(n18916), .A2(n12322), .ZN(n16310) );
  AND2_X1 U13160 ( .A1(n12530), .A2(n10276), .ZN(n12533) );
  INV_X1 U13161 ( .A(n16338), .ZN(n16321) );
  INV_X1 U13162 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19914) );
  OR2_X1 U13163 ( .A1(n19540), .A2(n19447), .ZN(n19332) );
  INV_X1 U13164 ( .A(n19350), .ZN(n19338) );
  OR2_X1 U13165 ( .A1(n19447), .A2(n19889), .ZN(n19373) );
  INV_X1 U13166 ( .A(n19410), .ZN(n19387) );
  INV_X1 U13167 ( .A(n19439), .ZN(n19433) );
  INV_X1 U13168 ( .A(n19472), .ZN(n19461) );
  INV_X1 U13169 ( .A(n19498), .ZN(n19505) );
  INV_X1 U13170 ( .A(n19531), .ZN(n19525) );
  INV_X1 U13171 ( .A(n19553), .ZN(n19569) );
  NAND2_X1 U13172 ( .A1(n19537), .A2(n19536), .ZN(n19604) );
  NAND2_X1 U13173 ( .A1(n19571), .A2(n19570), .ZN(n19635) );
  INV_X1 U13174 ( .A(n19718), .ZN(n19733) );
  NAND2_X1 U13175 ( .A1(n19537), .A2(n19742), .ZN(n19800) );
  INV_X1 U13176 ( .A(n19885), .ZN(n19811) );
  INV_X1 U13177 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n18887) );
  INV_X1 U13178 ( .A(n16950), .ZN(n16955) );
  INV_X1 U13179 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n17852) );
  NOR2_X1 U13180 ( .A1(n16651), .A2(n17012), .ZN(n17015) );
  NAND2_X1 U13181 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n17064), .ZN(n17052) );
  INV_X1 U13182 ( .A(n13304), .ZN(n17393) );
  NOR2_X1 U13183 ( .A1(n13083), .A2(n13082), .ZN(n17405) );
  NOR2_X1 U13184 ( .A1(n18881), .A2(n17429), .ZN(n17470) );
  NAND2_X1 U13185 ( .A1(n17489), .A2(n17427), .ZN(n17487) );
  INV_X1 U13186 ( .A(n17537), .ZN(n17532) );
  INV_X1 U13187 ( .A(n17690), .ZN(n17721) );
  INV_X1 U13188 ( .A(n17819), .ZN(n17808) );
  INV_X1 U13189 ( .A(n17903), .ZN(n17897) );
  INV_X1 U13190 ( .A(n18220), .ZN(n18195) );
  INV_X1 U13191 ( .A(n18227), .ZN(n18214) );
  NOR2_X1 U13192 ( .A1(n18247), .A2(n15814), .ZN(n18869) );
  INV_X1 U13193 ( .A(n18884), .ZN(n18743) );
  INV_X1 U13194 ( .A(n18835), .ZN(n18832) );
  OR2_X1 U13195 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n18759), .ZN(n18899) );
  CLKBUF_X1 U13196 ( .A(n16551), .Z(n16552) );
  NAND2_X1 U13197 ( .A1(n12559), .A2(n12558), .ZN(P1_U2873) );
  OAI211_X1 U13198 ( .C1(n19949), .C2(n14959), .A(n9902), .B(n12666), .ZN(
        P1_U2970) );
  OAI211_X1 U13199 ( .C1(n15483), .C2(n16293), .A(n12370), .B(n12369), .ZN(
        P2_U2986) );
  OAI21_X1 U13200 ( .B1(n15297), .B2(n16327), .A(n10261), .ZN(P2_U3017) );
  AND2_X4 U13201 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13716) );
  AND2_X4 U13202 ( .A1(n10289), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10284) );
  AOI22_X1 U13203 ( .A1(n10400), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n9842), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10288) );
  AOI22_X1 U13204 ( .A1(n10710), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n10595), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10287) );
  AND2_X4 U13205 ( .A1(n10284), .A2(n13744), .ZN(n11079) );
  AOI22_X1 U13206 ( .A1(n11079), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n10510), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10286) );
  AOI22_X1 U13207 ( .A1(n10342), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n10330), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10285) );
  NAND4_X1 U13208 ( .A1(n10288), .A2(n10287), .A3(n10286), .A4(n10285), .ZN(
        n10299) );
  AND2_X4 U13209 ( .A1(n10292), .A2(n10293), .ZN(n10499) );
  AOI22_X1 U13210 ( .A1(n10498), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n10499), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10297) );
  AOI22_X1 U13211 ( .A1(n10387), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n10596), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10296) );
  AOI22_X1 U13212 ( .A1(n10467), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n11064), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10295) );
  AND2_X4 U13213 ( .A1(n10293), .A2(n13716), .ZN(n10597) );
  NAND4_X1 U13214 ( .A1(n10297), .A2(n10296), .A3(n10295), .A4(n10294), .ZN(
        n10298) );
  NAND2_X1 U13215 ( .A1(n10400), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n10303) );
  NAND2_X1 U13216 ( .A1(n9842), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n10302) );
  NAND2_X1 U13217 ( .A1(n10930), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n10301) );
  NAND2_X1 U13218 ( .A1(n10330), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n10300) );
  NAND2_X1 U13219 ( .A1(n10387), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n10307) );
  NAND2_X1 U13220 ( .A1(n10710), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n10306) );
  NAND2_X1 U13221 ( .A1(n11079), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n10305) );
  NAND2_X1 U13222 ( .A1(n9864), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n10304) );
  NAND2_X1 U13223 ( .A1(n10342), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n10311) );
  NAND2_X1 U13224 ( .A1(n10467), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n10310) );
  NAND2_X1 U13225 ( .A1(n10498), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n10309) );
  NAND2_X1 U13226 ( .A1(n10499), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n10308) );
  NAND2_X1 U13227 ( .A1(n10335), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n10315) );
  NAND2_X1 U13228 ( .A1(n10595), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n10314) );
  NAND2_X1 U13229 ( .A1(n10596), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n10313) );
  NAND2_X1 U13230 ( .A1(n10597), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n10312) );
  NAND4_X4 U13231 ( .A1(n10319), .A2(n10318), .A3(n10317), .A4(n10316), .ZN(
        n11112) );
  AOI22_X1 U13232 ( .A1(n10498), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n9841), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10323) );
  AOI22_X1 U13233 ( .A1(n10400), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10499), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10322) );
  AOI22_X1 U13234 ( .A1(n9867), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n10330), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10321) );
  BUF_X4 U13235 ( .A(n11078), .Z(n10908) );
  AOI22_X1 U13236 ( .A1(n10342), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n10908), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10320) );
  NAND4_X1 U13237 ( .A1(n10323), .A2(n10322), .A3(n10321), .A4(n10320), .ZN(
        n10329) );
  AOI22_X1 U13238 ( .A1(n10467), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n10597), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10327) );
  AOI22_X1 U13239 ( .A1(n9861), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n10596), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10326) );
  AOI22_X1 U13240 ( .A1(n10335), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n9864), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10325) );
  AOI22_X1 U13241 ( .A1(n10710), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n10387), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10324) );
  NAND4_X1 U13242 ( .A1(n10327), .A2(n10326), .A3(n10325), .A4(n10324), .ZN(
        n10328) );
  AOI22_X1 U13243 ( .A1(n10498), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n9842), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10334) );
  AOI22_X1 U13244 ( .A1(n10400), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n10499), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10333) );
  AOI22_X1 U13245 ( .A1(n11079), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n10330), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10332) );
  AOI22_X1 U13246 ( .A1(n10342), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n10908), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10331) );
  NAND4_X1 U13247 ( .A1(n10334), .A2(n10333), .A3(n10332), .A4(n10331), .ZN(
        n10341) );
  AOI22_X1 U13248 ( .A1(n10710), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n10387), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10339) );
  AOI22_X1 U13249 ( .A1(n10335), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n9865), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10338) );
  AOI22_X1 U13250 ( .A1(n9862), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n10596), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10337) );
  AOI22_X1 U13251 ( .A1(n10467), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n10597), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10336) );
  NAND4_X1 U13252 ( .A1(n10339), .A2(n10338), .A3(n10337), .A4(n10336), .ZN(
        n10340) );
  OR2_X2 U13253 ( .A1(n10341), .A2(n10340), .ZN(n10415) );
  INV_X2 U13254 ( .A(n10415), .ZN(n13376) );
  AOI22_X1 U13255 ( .A1(n10498), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n10980), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10346) );
  AOI22_X1 U13256 ( .A1(n10400), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10499), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10345) );
  AOI22_X1 U13257 ( .A1(n10342), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n10510), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10344) );
  AOI22_X1 U13258 ( .A1(n10387), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n10596), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10343) );
  NAND4_X1 U13259 ( .A1(n10346), .A2(n10345), .A3(n10344), .A4(n10343), .ZN(
        n10352) );
  AOI22_X1 U13260 ( .A1(n10710), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n10595), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10350) );
  AOI22_X1 U13261 ( .A1(n11079), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n10467), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10349) );
  AOI22_X1 U13262 ( .A1(n10335), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n10597), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10348) );
  AOI22_X1 U13263 ( .A1(n10930), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n10330), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10347) );
  NAND4_X1 U13264 ( .A1(n10350), .A2(n10349), .A3(n10348), .A4(n10347), .ZN(
        n10351) );
  NAND2_X1 U13265 ( .A1(n13376), .A2(n12571), .ZN(n10416) );
  INV_X1 U13266 ( .A(n10416), .ZN(n10353) );
  NAND2_X1 U13267 ( .A1(n10354), .A2(n10353), .ZN(n13487) );
  AOI22_X1 U13268 ( .A1(n10498), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n10980), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n10358) );
  AOI22_X1 U13269 ( .A1(n10400), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n10499), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10357) );
  AOI22_X1 U13270 ( .A1(n11079), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n10330), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10356) );
  AOI22_X1 U13271 ( .A1(n10342), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n10908), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10355) );
  NAND4_X1 U13272 ( .A1(n10358), .A2(n10357), .A3(n10356), .A4(n10355), .ZN(
        n10364) );
  AOI22_X1 U13273 ( .A1(n10710), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n10387), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10362) );
  AOI22_X1 U13274 ( .A1(n10335), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n10510), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10361) );
  AOI22_X1 U13275 ( .A1(n10595), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n10596), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n10360) );
  AOI22_X1 U13276 ( .A1(n10467), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n10597), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10359) );
  NAND4_X1 U13277 ( .A1(n10362), .A2(n10361), .A3(n10360), .A4(n10359), .ZN(
        n10363) );
  NAND2_X1 U13278 ( .A1(n10387), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n10368) );
  NAND2_X1 U13279 ( .A1(n10710), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n10367) );
  NAND2_X1 U13280 ( .A1(n10595), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n10366) );
  NAND2_X1 U13281 ( .A1(n10596), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n10365) );
  NAND2_X1 U13282 ( .A1(n10498), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n10372) );
  NAND2_X1 U13283 ( .A1(n10980), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n10371) );
  NAND2_X1 U13284 ( .A1(n10499), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n10370) );
  NAND2_X1 U13285 ( .A1(n10400), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n10369) );
  NAND2_X1 U13286 ( .A1(n10335), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n10376) );
  NAND2_X1 U13287 ( .A1(n9864), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n10374) );
  NAND2_X1 U13288 ( .A1(n10597), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n10373) );
  NAND2_X1 U13289 ( .A1(n11079), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n10380) );
  NAND2_X1 U13290 ( .A1(n10342), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n10379) );
  NAND2_X1 U13291 ( .A1(n10330), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n10378) );
  NAND2_X1 U13292 ( .A1(n10930), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n10377) );
  NAND2_X1 U13293 ( .A1(n13371), .A2(n9854), .ZN(n11161) );
  INV_X1 U13294 ( .A(n11161), .ZN(n10386) );
  NAND2_X1 U13295 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n20702) );
  OAI21_X1 U13296 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(P1_STATE_REG_2__SCAN_IN), 
        .A(n20702), .ZN(n11270) );
  INV_X1 U13297 ( .A(n11270), .ZN(n10385) );
  NAND2_X1 U13298 ( .A1(n10386), .A2(n10385), .ZN(n10412) );
  NAND2_X1 U13299 ( .A1(n10387), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n10391) );
  NAND2_X1 U13300 ( .A1(n10335), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n10390) );
  NAND2_X1 U13301 ( .A1(n10710), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n10389) );
  NAND2_X1 U13302 ( .A1(n10597), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n10388) );
  NAND2_X1 U13303 ( .A1(n10342), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n10395) );
  NAND2_X1 U13304 ( .A1(n10467), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n10394) );
  NAND2_X1 U13305 ( .A1(n10498), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n10393) );
  NAND2_X1 U13306 ( .A1(n9842), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n10392) );
  NAND2_X1 U13307 ( .A1(n10595), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n10399) );
  NAND2_X1 U13308 ( .A1(n11079), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n10398) );
  NAND2_X1 U13309 ( .A1(n10510), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n10397) );
  NAND2_X1 U13310 ( .A1(n10596), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n10396) );
  NAND2_X1 U13311 ( .A1(n10499), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n10404) );
  NAND2_X1 U13312 ( .A1(n10400), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n10403) );
  NAND2_X1 U13313 ( .A1(n10930), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n10402) );
  NAND2_X1 U13314 ( .A1(n10330), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n10401) );
  NAND3_X1 U13315 ( .A1(n13959), .A2(n10418), .A3(n13809), .ZN(n13709) );
  NAND2_X2 U13316 ( .A1(n10422), .A2(n11112), .ZN(n13618) );
  NAND2_X1 U13317 ( .A1(n10474), .A2(n14519), .ZN(n10409) );
  NAND2_X1 U13318 ( .A1(n13376), .A2(n11112), .ZN(n12566) );
  NAND3_X1 U13319 ( .A1(n12566), .A2(n20177), .A3(n13392), .ZN(n10410) );
  NAND2_X1 U13320 ( .A1(n9894), .A2(n10410), .ZN(n10428) );
  NOR2_X1 U13321 ( .A1(n11105), .A2(n9854), .ZN(n10411) );
  NAND2_X1 U13322 ( .A1(n13371), .A2(n13808), .ZN(n13385) );
  NAND4_X1 U13323 ( .A1(n10412), .A2(n13386), .A3(n12536), .A4(n13385), .ZN(
        n10413) );
  NAND2_X1 U13324 ( .A1(n10415), .A2(n9854), .ZN(n13405) );
  NAND2_X1 U13325 ( .A1(n11175), .A2(n10416), .ZN(n13390) );
  NAND2_X1 U13326 ( .A1(n10418), .A2(n10417), .ZN(n10419) );
  NAND2_X1 U13327 ( .A1(n12560), .A2(n20182), .ZN(n10444) );
  NAND2_X1 U13328 ( .A1(n10440), .A2(n13781), .ZN(n10425) );
  INV_X1 U13329 ( .A(n9854), .ZN(n20157) );
  AOI21_X1 U13330 ( .B1(n12630), .B2(n20190), .A(n20157), .ZN(n10424) );
  NAND3_X1 U13331 ( .A1(n13711), .A2(n10425), .A3(n13403), .ZN(n10426) );
  NAND2_X1 U13332 ( .A1(n10426), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10431) );
  NAND2_X1 U13333 ( .A1(n11105), .A2(n10415), .ZN(n10427) );
  NAND3_X1 U13334 ( .A1(n13399), .A2(n20168), .A3(n13718), .ZN(n10429) );
  NAND2_X1 U13335 ( .A1(n15073), .A2(n20806), .ZN(n12660) );
  NAND2_X1 U13336 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n10456) );
  OAI21_X1 U13337 ( .B1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n10456), .ZN(n20465) );
  NAND2_X1 U13338 ( .A1(n20695), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n10450) );
  OAI21_X1 U13339 ( .B1(n12660), .B2(n20465), .A(n10450), .ZN(n10432) );
  NAND2_X1 U13340 ( .A1(n10454), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10436) );
  MUX2_X1 U13341 ( .A(n12660), .B(n15897), .S(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .Z(n10435) );
  AOI21_X1 U13342 ( .B1(n13618), .B2(n12571), .A(n13477), .ZN(n10438) );
  INV_X1 U13343 ( .A(n13399), .ZN(n10437) );
  MUX2_X1 U13344 ( .A(n10438), .B(n10437), .S(n13959), .Z(n10439) );
  NAND3_X1 U13345 ( .A1(n10440), .A2(n9858), .A3(n13781), .ZN(n10447) );
  INV_X1 U13346 ( .A(n10441), .ZN(n10443) );
  NAND2_X1 U13347 ( .A1(n20157), .A2(n9858), .ZN(n13961) );
  NAND3_X1 U13348 ( .A1(n13961), .A2(n15073), .A3(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n10442) );
  NOR2_X1 U13349 ( .A1(n10443), .A2(n10442), .ZN(n10446) );
  NAND2_X1 U13350 ( .A1(n10444), .A2(n15891), .ZN(n10445) );
  AND2_X2 U13351 ( .A1(n10497), .A2(n10495), .ZN(n10477) );
  NAND2_X1 U13352 ( .A1(n10450), .A2(n10289), .ZN(n10451) );
  NAND2_X1 U13353 ( .A1(n10452), .A2(n10451), .ZN(n10453) );
  NAND2_X1 U13354 ( .A1(n10454), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10460) );
  INV_X1 U13355 ( .A(n12660), .ZN(n10458) );
  INV_X1 U13356 ( .A(n10456), .ZN(n10455) );
  NAND2_X1 U13357 ( .A1(n10455), .A2(n20461), .ZN(n20493) );
  NAND2_X1 U13358 ( .A1(n10456), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n10457) );
  NAND2_X1 U13359 ( .A1(n20493), .A2(n10457), .ZN(n20163) );
  AOI22_X1 U13360 ( .A1(n10458), .A2(n20163), .B1(n20695), .B2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n10459) );
  NAND2_X2 U13361 ( .A1(n10462), .A2(n10461), .ZN(n13758) );
  AOI22_X1 U13362 ( .A1(n11023), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n9863), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n10466) );
  AOI22_X1 U13363 ( .A1(n11057), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n10499), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10465) );
  AOI22_X1 U13364 ( .A1(n9867), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n11058), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10464) );
  AOI22_X1 U13365 ( .A1(n11065), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n10908), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10463) );
  NAND4_X1 U13366 ( .A1(n10466), .A2(n10465), .A3(n10464), .A4(n10463), .ZN(
        n10473) );
  AOI22_X1 U13367 ( .A1(n10925), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11085), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10471) );
  AOI22_X1 U13368 ( .A1(n11059), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n9864), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10470) );
  AOI22_X1 U13369 ( .A1(n10595), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n10481), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10469) );
  AOI22_X1 U13370 ( .A1(n11080), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n10597), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10468) );
  NAND4_X1 U13371 ( .A1(n10471), .A2(n10470), .A3(n10469), .A4(n10468), .ZN(
        n10472) );
  AOI22_X1 U13372 ( .A1(n11147), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n10527), .B2(n10475), .ZN(n10476) );
  INV_X1 U13373 ( .A(n20264), .ZN(n10479) );
  INV_X1 U13374 ( .A(n10477), .ZN(n10478) );
  INV_X1 U13375 ( .A(n13910), .ZN(n10480) );
  NAND2_X1 U13376 ( .A1(n10480), .A2(n20806), .ZN(n10494) );
  AOI22_X1 U13377 ( .A1(n10925), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n11085), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10485) );
  AOI22_X1 U13378 ( .A1(n11065), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11057), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10484) );
  AOI22_X1 U13379 ( .A1(n11079), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n9864), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10483) );
  AOI22_X1 U13380 ( .A1(n9862), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n10481), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10482) );
  NAND4_X1 U13381 ( .A1(n10485), .A2(n10484), .A3(n10483), .A4(n10482), .ZN(
        n10491) );
  AOI22_X1 U13382 ( .A1(n11023), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n10499), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10489) );
  AOI22_X1 U13383 ( .A1(n11080), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n11058), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10488) );
  AOI22_X1 U13384 ( .A1(n9863), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n11064), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10487) );
  AOI22_X1 U13385 ( .A1(n11059), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n10597), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10486) );
  NAND4_X1 U13386 ( .A1(n10489), .A2(n10488), .A3(n10487), .A4(n10486), .ZN(
        n10490) );
  INV_X1 U13387 ( .A(n12564), .ZN(n10492) );
  OR2_X1 U13388 ( .A1(n10563), .A2(n10492), .ZN(n10493) );
  AND2_X2 U13389 ( .A1(n10494), .A2(n10493), .ZN(n12563) );
  AOI22_X1 U13390 ( .A1(n11023), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n9863), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n10503) );
  AOI22_X1 U13391 ( .A1(n11057), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n10499), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10502) );
  AOI22_X1 U13392 ( .A1(n11079), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n11058), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10501) );
  AOI22_X1 U13393 ( .A1(n9831), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n10908), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10500) );
  NAND4_X1 U13394 ( .A1(n10503), .A2(n10502), .A3(n10501), .A4(n10500), .ZN(
        n10509) );
  AOI22_X1 U13395 ( .A1(n10925), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n10387), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10507) );
  AOI22_X1 U13396 ( .A1(n10335), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n9864), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10506) );
  AOI22_X1 U13397 ( .A1(n9862), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n10481), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10505) );
  AOI22_X1 U13398 ( .A1(n11080), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n10597), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10504) );
  NAND4_X1 U13399 ( .A1(n10507), .A2(n10506), .A3(n10505), .A4(n10504), .ZN(
        n10508) );
  NOR2_X1 U13400 ( .A1(n10563), .A2(n12633), .ZN(n10526) );
  AOI22_X1 U13401 ( .A1(n11065), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n9863), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10514) );
  AOI22_X1 U13402 ( .A1(n11057), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10499), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10513) );
  AOI22_X1 U13403 ( .A1(n10925), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10595), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10512) );
  AOI22_X1 U13404 ( .A1(n9864), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n11058), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10511) );
  NAND4_X1 U13405 ( .A1(n10514), .A2(n10513), .A3(n10512), .A4(n10511), .ZN(
        n10520) );
  AOI22_X1 U13406 ( .A1(n11079), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n11080), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10518) );
  AOI22_X1 U13407 ( .A1(n11085), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n10481), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10517) );
  AOI22_X1 U13408 ( .A1(n11023), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11064), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10516) );
  AOI22_X1 U13409 ( .A1(n11059), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n10597), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10515) );
  NAND4_X1 U13410 ( .A1(n10518), .A2(n10517), .A3(n10516), .A4(n10515), .ZN(
        n10519) );
  MUX2_X1 U13411 ( .A(n12631), .B(n10526), .S(n12570), .Z(n10521) );
  NOR2_X1 U13412 ( .A1(n12570), .A2(n20806), .ZN(n10525) );
  NAND2_X1 U13413 ( .A1(n11147), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n10524) );
  NAND2_X1 U13414 ( .A1(n11147), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n10530) );
  INV_X1 U13415 ( .A(n10526), .ZN(n10529) );
  NAND2_X1 U13416 ( .A1(n10527), .A2(n12564), .ZN(n10528) );
  INV_X1 U13417 ( .A(n10531), .ZN(n10532) );
  AOI21_X2 U13418 ( .B1(n12563), .B2(n10542), .A(n10534), .ZN(n10535) );
  NAND2_X2 U13419 ( .A1(n10536), .A2(n10535), .ZN(n10578) );
  INV_X1 U13420 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n13775) );
  XNOR2_X1 U13421 ( .A(n13775), .B(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n20035) );
  INV_X1 U13422 ( .A(n12658), .ZN(n10660) );
  OAI21_X1 U13423 ( .B1(n20035), .B2(n10609), .A(n10660), .ZN(n10538) );
  AOI21_X1 U13424 ( .B1(n11049), .B2(P1_EAX_REG_2__SCAN_IN), .A(n10538), .ZN(
        n10540) );
  AND2_X1 U13425 ( .A1(n13392), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n10606) );
  NAND2_X1 U13426 ( .A1(n10606), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10539) );
  NAND2_X1 U13427 ( .A1(n12658), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10558) );
  NAND2_X1 U13428 ( .A1(n13911), .A2(n10671), .ZN(n10548) );
  AOI22_X1 U13429 ( .A1(n11049), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n20802), .ZN(n10546) );
  NAND2_X1 U13430 ( .A1(n10606), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10545) );
  AND2_X1 U13431 ( .A1(n10546), .A2(n10545), .ZN(n10547) );
  NAND2_X1 U13432 ( .A1(n12574), .A2(n20190), .ZN(n10550) );
  NAND2_X1 U13433 ( .A1(n10550), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13609) );
  INV_X1 U13434 ( .A(n10606), .ZN(n10587) );
  NAND2_X1 U13435 ( .A1(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n20802), .ZN(
        n10554) );
  NAND2_X1 U13436 ( .A1(n10552), .A2(P1_EAX_REG_0__SCAN_IN), .ZN(n10553) );
  OAI211_X1 U13437 ( .C1(n10587), .C2(n9947), .A(n10554), .B(n10553), .ZN(
        n10555) );
  AOI21_X1 U13438 ( .B1(n10551), .B2(n10671), .A(n10555), .ZN(n13610) );
  OR2_X1 U13439 ( .A1(n13609), .A2(n13610), .ZN(n13607) );
  INV_X1 U13440 ( .A(n13610), .ZN(n10556) );
  OR2_X1 U13441 ( .A1(n10556), .A2(n10609), .ZN(n10557) );
  NAND2_X1 U13442 ( .A1(n13607), .A2(n10557), .ZN(n13700) );
  NAND2_X1 U13443 ( .A1(n13765), .A2(n13764), .ZN(n13763) );
  NAND2_X2 U13444 ( .A1(n13763), .A2(n10558), .ZN(n13876) );
  INV_X1 U13445 ( .A(n10578), .ZN(n10577) );
  NAND2_X1 U13446 ( .A1(n10454), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10561) );
  NOR3_X1 U13447 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n20461), .A3(
        n20523), .ZN(n20384) );
  INV_X1 U13448 ( .A(n20384), .ZN(n20380) );
  NAND3_X1 U13449 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20633) );
  INV_X1 U13450 ( .A(n20633), .ZN(n20640) );
  NAND2_X1 U13451 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20640), .ZN(
        n20630) );
  OAI21_X1 U13452 ( .B1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n20401), .A(
        n20630), .ZN(n20406) );
  OAI22_X1 U13453 ( .A1(n12660), .A2(n20406), .B1(n15897), .B2(n20783), .ZN(
        n10559) );
  INV_X1 U13454 ( .A(n10559), .ZN(n10560) );
  AOI22_X1 U13455 ( .A1(n11059), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n11085), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10567) );
  AOI22_X1 U13456 ( .A1(n11023), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10499), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10566) );
  AOI22_X1 U13457 ( .A1(n11080), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n10597), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10565) );
  AOI22_X1 U13458 ( .A1(n9863), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n10908), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10564) );
  NAND4_X1 U13459 ( .A1(n10567), .A2(n10566), .A3(n10565), .A4(n10564), .ZN(
        n10573) );
  AOI22_X1 U13460 ( .A1(n11065), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11057), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10571) );
  AOI22_X1 U13461 ( .A1(n10595), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n9864), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10570) );
  AOI22_X1 U13462 ( .A1(n10925), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n10481), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10569) );
  AOI22_X1 U13463 ( .A1(n11079), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11058), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10568) );
  NAND4_X1 U13464 ( .A1(n10571), .A2(n10570), .A3(n10569), .A4(n10568), .ZN(
        n10572) );
  AOI22_X1 U13465 ( .A1(n11155), .A2(n12603), .B1(n11147), .B2(
        P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10574) );
  NAND2_X1 U13466 ( .A1(n10578), .A2(n20294), .ZN(n10579) );
  INV_X1 U13467 ( .A(n20772), .ZN(n10580) );
  NAND2_X1 U13468 ( .A1(n10580), .A2(n10671), .ZN(n10590) );
  INV_X1 U13469 ( .A(n10582), .ZN(n10584) );
  INV_X1 U13470 ( .A(n10608), .ZN(n10583) );
  OAI21_X1 U13471 ( .B1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n10584), .A(
        n10583), .ZN(n13975) );
  AOI22_X1 U13472 ( .A1(n11096), .A2(n13975), .B1(n12658), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n10586) );
  NAND2_X1 U13473 ( .A1(n11049), .A2(P1_EAX_REG_3__SCAN_IN), .ZN(n10585) );
  OAI211_X1 U13474 ( .C1(n10587), .C2(n10581), .A(n10586), .B(n10585), .ZN(
        n10588) );
  INV_X1 U13475 ( .A(n10588), .ZN(n10589) );
  AOI22_X1 U13476 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n11023), .B1(
        n9863), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n10594) );
  AOI22_X1 U13477 ( .A1(n11057), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n10499), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10593) );
  AOI22_X1 U13478 ( .A1(n11079), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n11058), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10592) );
  INV_X1 U13479 ( .A(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n21135) );
  AOI22_X1 U13480 ( .A1(n11065), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n10908), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10591) );
  NAND4_X1 U13481 ( .A1(n10594), .A2(n10593), .A3(n10592), .A4(n10591), .ZN(
        n10603) );
  AOI22_X1 U13482 ( .A1(n10925), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n11085), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10601) );
  AOI22_X1 U13483 ( .A1(n11059), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n9865), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10600) );
  AOI22_X1 U13484 ( .A1(n10595), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n10481), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10599) );
  AOI22_X1 U13485 ( .A1(n11080), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n10597), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10598) );
  NAND4_X1 U13486 ( .A1(n10601), .A2(n10600), .A3(n10599), .A4(n10598), .ZN(
        n10602) );
  NAND2_X1 U13487 ( .A1(n11155), .A2(n12602), .ZN(n10605) );
  NAND2_X1 U13488 ( .A1(n11147), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n10604) );
  XNOR2_X1 U13489 ( .A(n10628), .B(n10631), .ZN(n12594) );
  NAND2_X1 U13490 ( .A1(n10606), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n10612) );
  INV_X1 U13491 ( .A(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n20013) );
  AOI21_X1 U13492 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n20013), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n10607) );
  AOI21_X1 U13493 ( .B1(n11049), .B2(P1_EAX_REG_4__SCAN_IN), .A(n10607), .ZN(
        n10611) );
  OAI21_X1 U13494 ( .B1(n10608), .B2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n10634), .ZN(n20101) );
  NOR2_X1 U13495 ( .A1(n20101), .A2(n10609), .ZN(n10610) );
  AOI21_X1 U13496 ( .B1(n10612), .B2(n10611), .A(n10610), .ZN(n10613) );
  INV_X1 U13497 ( .A(n10631), .ZN(n10627) );
  AOI22_X1 U13498 ( .A1(n11023), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n9863), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10618) );
  AOI22_X1 U13499 ( .A1(n11057), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n10499), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10617) );
  AOI22_X1 U13500 ( .A1(n9867), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11058), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10616) );
  AOI22_X1 U13501 ( .A1(n11065), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10908), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10615) );
  NAND4_X1 U13502 ( .A1(n10618), .A2(n10617), .A3(n10616), .A4(n10615), .ZN(
        n10624) );
  AOI22_X1 U13503 ( .A1(n10925), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11085), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10622) );
  AOI22_X1 U13504 ( .A1(n10335), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n9865), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10621) );
  AOI22_X1 U13505 ( .A1(n10595), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n10481), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10620) );
  AOI22_X1 U13506 ( .A1(n11080), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10597), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10619) );
  NAND4_X1 U13507 ( .A1(n10622), .A2(n10621), .A3(n10620), .A4(n10619), .ZN(
        n10623) );
  NAND2_X1 U13508 ( .A1(n11155), .A2(n12614), .ZN(n10626) );
  NAND2_X1 U13509 ( .A1(n11147), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n10625) );
  OAI21_X1 U13510 ( .B1(n10628), .B2(n10627), .A(n10629), .ZN(n10632) );
  INV_X1 U13511 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n10638) );
  INV_X1 U13512 ( .A(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n10633) );
  NAND2_X1 U13513 ( .A1(n10634), .A2(n10633), .ZN(n10636) );
  NAND2_X1 U13514 ( .A1(n10636), .A2(n10655), .ZN(n20007) );
  AOI22_X1 U13515 ( .A1(n20007), .A2(n11096), .B1(n12658), .B2(
        P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n10637) );
  OAI21_X1 U13516 ( .B1(n10639), .B2(n10638), .A(n10637), .ZN(n10640) );
  NAND2_X1 U13517 ( .A1(n10642), .A2(n10641), .ZN(n13939) );
  AOI22_X1 U13518 ( .A1(n11023), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n9863), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10646) );
  AOI22_X1 U13519 ( .A1(n11057), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n10499), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10645) );
  AOI22_X1 U13520 ( .A1(n9867), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11058), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10644) );
  AOI22_X1 U13521 ( .A1(n11065), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n10908), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10643) );
  NAND4_X1 U13522 ( .A1(n10646), .A2(n10645), .A3(n10644), .A4(n10643), .ZN(
        n10652) );
  AOI22_X1 U13523 ( .A1(n10925), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11085), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10650) );
  AOI22_X1 U13524 ( .A1(n10335), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n9865), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10649) );
  AOI22_X1 U13525 ( .A1(n9861), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n10481), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10648) );
  AOI22_X1 U13526 ( .A1(n11080), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n10597), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10647) );
  NAND4_X1 U13527 ( .A1(n10650), .A2(n10649), .A3(n10648), .A4(n10647), .ZN(
        n10651) );
  NAND2_X1 U13528 ( .A1(n11155), .A2(n12622), .ZN(n10654) );
  NAND2_X1 U13529 ( .A1(n11147), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n10653) );
  NAND2_X1 U13530 ( .A1(n10666), .A2(n10667), .ZN(n12613) );
  INV_X1 U13531 ( .A(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n10659) );
  OAI21_X1 U13532 ( .B1(n10656), .B2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n10663), .ZN(n19996) );
  NAND2_X1 U13533 ( .A1(n19996), .A2(n11096), .ZN(n10658) );
  NAND2_X1 U13534 ( .A1(n11049), .A2(P1_EAX_REG_6__SCAN_IN), .ZN(n10657) );
  OAI211_X1 U13535 ( .C1(n10660), .C2(n10659), .A(n10658), .B(n10657), .ZN(
        n10661) );
  NOR2_X2 U13536 ( .A1(n13939), .A2(n14000), .ZN(n13989) );
  INV_X1 U13537 ( .A(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n10662) );
  NAND2_X1 U13538 ( .A1(n10663), .A2(n10662), .ZN(n10665) );
  NAND2_X1 U13539 ( .A1(n10665), .A2(n10690), .ZN(n19985) );
  INV_X1 U13540 ( .A(n19985), .ZN(n10675) );
  AOI22_X1 U13541 ( .A1(n11155), .A2(n12633), .B1(n11147), .B2(
        P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10670) );
  INV_X1 U13542 ( .A(n12621), .ZN(n10672) );
  INV_X1 U13543 ( .A(n10801), .ZN(n10671) );
  NAND2_X1 U13544 ( .A1(n10672), .A2(n10671), .ZN(n10674) );
  AOI22_X1 U13545 ( .A1(n11049), .A2(P1_EAX_REG_7__SCAN_IN), .B1(n12658), .B2(
        P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n10673) );
  NAND2_X1 U13546 ( .A1(n13989), .A2(n13988), .ZN(n13987) );
  AOI22_X1 U13547 ( .A1(n10925), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n11085), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10679) );
  AOI22_X1 U13548 ( .A1(n11023), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10499), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10678) );
  AOI22_X1 U13549 ( .A1(n9865), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n10481), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10677) );
  AOI22_X1 U13550 ( .A1(n10930), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n11058), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10676) );
  NAND4_X1 U13551 ( .A1(n10679), .A2(n10678), .A3(n10677), .A4(n10676), .ZN(
        n10685) );
  AOI22_X1 U13552 ( .A1(n9867), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n11065), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10683) );
  AOI22_X1 U13553 ( .A1(n11057), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n9863), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10682) );
  AOI22_X1 U13554 ( .A1(n10335), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n9862), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10681) );
  AOI22_X1 U13555 ( .A1(n11080), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10597), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10680) );
  NAND4_X1 U13556 ( .A1(n10683), .A2(n10682), .A3(n10681), .A4(n10680), .ZN(
        n10684) );
  OAI21_X1 U13557 ( .B1(n10685), .B2(n10684), .A(n10671), .ZN(n10689) );
  INV_X1 U13558 ( .A(n10690), .ZN(n10686) );
  XNOR2_X1 U13559 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B(n10686), .ZN(
        n14250) );
  AOI22_X1 U13560 ( .A1(n11096), .A2(n14250), .B1(n12658), .B2(
        P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n10688) );
  NAND2_X1 U13561 ( .A1(n11049), .A2(P1_EAX_REG_8__SCAN_IN), .ZN(n10687) );
  NOR2_X2 U13562 ( .A1(n13987), .A2(n14073), .ZN(n14071) );
  XNOR2_X1 U13563 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .B(n10706), .ZN(
        n19971) );
  INV_X1 U13564 ( .A(n19971), .ZN(n14283) );
  AOI22_X1 U13565 ( .A1(n9831), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n9863), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10694) );
  AOI22_X1 U13566 ( .A1(n11023), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n10499), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10693) );
  AOI22_X1 U13567 ( .A1(n10925), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n10481), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10692) );
  AOI22_X1 U13568 ( .A1(n9861), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n11058), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10691) );
  NAND4_X1 U13569 ( .A1(n10694), .A2(n10693), .A3(n10692), .A4(n10691), .ZN(
        n10700) );
  AOI22_X1 U13570 ( .A1(n9867), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n11080), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10698) );
  AOI22_X1 U13571 ( .A1(n11085), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n9865), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10697) );
  AOI22_X1 U13572 ( .A1(n11057), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n10908), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10696) );
  AOI22_X1 U13573 ( .A1(n10335), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n10597), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10695) );
  NAND4_X1 U13574 ( .A1(n10698), .A2(n10697), .A3(n10696), .A4(n10695), .ZN(
        n10699) );
  OAI21_X1 U13575 ( .B1(n10700), .B2(n10699), .A(n10671), .ZN(n10703) );
  NAND2_X1 U13576 ( .A1(n11049), .A2(P1_EAX_REG_9__SCAN_IN), .ZN(n10702) );
  NAND2_X1 U13577 ( .A1(n12658), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n10701) );
  NAND3_X1 U13578 ( .A1(n10703), .A2(n10702), .A3(n10701), .ZN(n10704) );
  AOI21_X1 U13579 ( .B1(n14283), .B2(n11096), .A(n10704), .ZN(n14201) );
  NAND2_X1 U13580 ( .A1(n10707), .A2(n21019), .ZN(n10709) );
  INV_X1 U13581 ( .A(n10726), .ZN(n10708) );
  NAND2_X1 U13582 ( .A1(n10709), .A2(n10708), .ZN(n16033) );
  NAND2_X1 U13583 ( .A1(n16033), .A2(n11096), .ZN(n10725) );
  AOI22_X1 U13584 ( .A1(n10925), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n11085), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10714) );
  AOI22_X1 U13585 ( .A1(n11065), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n9863), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10713) );
  AOI22_X1 U13586 ( .A1(n11057), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n10499), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10712) );
  AOI22_X1 U13587 ( .A1(n10595), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n9833), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10711) );
  NAND4_X1 U13588 ( .A1(n10714), .A2(n10713), .A3(n10712), .A4(n10711), .ZN(
        n10720) );
  AOI22_X1 U13589 ( .A1(n10335), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n10481), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10718) );
  AOI22_X1 U13590 ( .A1(n11023), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n10930), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10717) );
  AOI22_X1 U13591 ( .A1(n9867), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11058), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10716) );
  AOI22_X1 U13592 ( .A1(n11080), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n10597), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10715) );
  NAND4_X1 U13593 ( .A1(n10718), .A2(n10717), .A3(n10716), .A4(n10715), .ZN(
        n10719) );
  OAI21_X1 U13594 ( .B1(n10720), .B2(n10719), .A(n10671), .ZN(n10723) );
  NAND2_X1 U13595 ( .A1(n11049), .A2(P1_EAX_REG_10__SCAN_IN), .ZN(n10722) );
  NAND2_X1 U13596 ( .A1(n12658), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n10721) );
  AND3_X1 U13597 ( .A1(n10723), .A2(n10722), .A3(n10721), .ZN(n10724) );
  NAND2_X1 U13598 ( .A1(n11049), .A2(P1_EAX_REG_11__SCAN_IN), .ZN(n10728) );
  OAI21_X1 U13599 ( .B1(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n10726), .A(
        n10764), .ZN(n16088) );
  AOI22_X1 U13600 ( .A1(n11096), .A2(n16088), .B1(n12658), .B2(
        P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n10727) );
  NAND2_X1 U13601 ( .A1(n10728), .A2(n10727), .ZN(n14300) );
  AOI22_X1 U13602 ( .A1(n11023), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n9863), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10732) );
  AOI22_X1 U13603 ( .A1(n11057), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n10499), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10731) );
  AOI22_X1 U13604 ( .A1(n11059), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n10481), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10730) );
  AOI22_X1 U13605 ( .A1(n11080), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n10597), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10729) );
  NAND4_X1 U13606 ( .A1(n10732), .A2(n10731), .A3(n10730), .A4(n10729), .ZN(
        n10738) );
  AOI22_X1 U13607 ( .A1(n10925), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11085), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10736) );
  AOI22_X1 U13608 ( .A1(n10595), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n9865), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10735) );
  AOI22_X1 U13609 ( .A1(n11065), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n10908), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10734) );
  AOI22_X1 U13610 ( .A1(n11079), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n11058), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10733) );
  NAND4_X1 U13611 ( .A1(n10736), .A2(n10735), .A3(n10734), .A4(n10733), .ZN(
        n10737) );
  OR2_X1 U13612 ( .A1(n10738), .A2(n10737), .ZN(n10739) );
  NAND2_X1 U13613 ( .A1(n10671), .A2(n10739), .ZN(n14637) );
  INV_X1 U13614 ( .A(n14637), .ZN(n14304) );
  AOI22_X1 U13615 ( .A1(n11065), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n9863), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10743) );
  AOI22_X1 U13616 ( .A1(n11057), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n10499), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10742) );
  AOI22_X1 U13617 ( .A1(n9867), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(n9865), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10741) );
  AOI22_X1 U13618 ( .A1(n9862), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n10481), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10740) );
  NAND4_X1 U13619 ( .A1(n10743), .A2(n10742), .A3(n10741), .A4(n10740), .ZN(
        n10749) );
  AOI22_X1 U13620 ( .A1(n10925), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11085), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10747) );
  AOI22_X1 U13621 ( .A1(n11080), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11058), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10746) );
  AOI22_X1 U13622 ( .A1(n11023), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n10908), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10745) );
  AOI22_X1 U13623 ( .A1(n11059), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10597), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10744) );
  NAND4_X1 U13624 ( .A1(n10747), .A2(n10746), .A3(n10745), .A4(n10744), .ZN(
        n10748) );
  NOR2_X1 U13625 ( .A1(n10749), .A2(n10748), .ZN(n10753) );
  XNOR2_X1 U13626 ( .A(n10771), .B(n14648), .ZN(n14929) );
  NAND2_X1 U13627 ( .A1(n14929), .A2(n11096), .ZN(n10752) );
  AOI22_X1 U13628 ( .A1(n11049), .A2(P1_EAX_REG_13__SCAN_IN), .B1(n12658), 
        .B2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n10751) );
  OAI211_X1 U13629 ( .C1(n10753), .C2(n10801), .A(n10752), .B(n10751), .ZN(
        n14640) );
  AOI22_X1 U13630 ( .A1(n10925), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n11085), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10757) );
  AOI22_X1 U13631 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n11057), .B1(
        n9863), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n10756) );
  AOI22_X1 U13632 ( .A1(n9862), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n9865), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10755) );
  AOI22_X1 U13633 ( .A1(n9831), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n10930), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10754) );
  NAND4_X1 U13634 ( .A1(n10757), .A2(n10756), .A3(n10755), .A4(n10754), .ZN(
        n10763) );
  AOI22_X1 U13635 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n11023), .B1(
        n10499), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10761) );
  AOI22_X1 U13636 ( .A1(n11059), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n10481), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10760) );
  AOI22_X1 U13637 ( .A1(n9867), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n11058), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10759) );
  AOI22_X1 U13638 ( .A1(n11080), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n10597), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10758) );
  NAND4_X1 U13639 ( .A1(n10761), .A2(n10760), .A3(n10759), .A4(n10758), .ZN(
        n10762) );
  OAI21_X1 U13640 ( .B1(n10763), .B2(n10762), .A(n10671), .ZN(n10769) );
  NAND2_X1 U13641 ( .A1(n11049), .A2(P1_EAX_REG_12__SCAN_IN), .ZN(n10768) );
  XNOR2_X1 U13642 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B(n10764), .ZN(
        n16076) );
  NAND2_X1 U13643 ( .A1(n12658), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n10765) );
  OAI21_X1 U13644 ( .B1(n16076), .B2(n10609), .A(n10765), .ZN(n10766) );
  INV_X1 U13645 ( .A(n10766), .ZN(n10767) );
  NAND3_X1 U13646 ( .A1(n10769), .A2(n10768), .A3(n10767), .ZN(n14743) );
  XOR2_X1 U13647 ( .A(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B(n10787), .Z(
        n16068) );
  INV_X1 U13648 ( .A(n16068), .ZN(n10786) );
  AOI22_X1 U13649 ( .A1(n11065), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n9863), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10775) );
  AOI22_X1 U13650 ( .A1(n11057), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n10499), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10774) );
  AOI22_X1 U13651 ( .A1(n10925), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n10481), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10773) );
  AOI22_X1 U13652 ( .A1(n9867), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n11058), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10772) );
  NAND4_X1 U13653 ( .A1(n10775), .A2(n10774), .A3(n10773), .A4(n10772), .ZN(
        n10781) );
  AOI22_X1 U13654 ( .A1(n11085), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n9861), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10779) );
  AOI22_X1 U13655 ( .A1(n11059), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n9865), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10778) );
  AOI22_X1 U13656 ( .A1(n11023), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n10908), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10777) );
  AOI22_X1 U13657 ( .A1(n11080), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n10597), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10776) );
  NAND4_X1 U13658 ( .A1(n10779), .A2(n10778), .A3(n10777), .A4(n10776), .ZN(
        n10780) );
  NOR2_X1 U13659 ( .A1(n10781), .A2(n10780), .ZN(n10784) );
  NAND2_X1 U13660 ( .A1(n11049), .A2(P1_EAX_REG_14__SCAN_IN), .ZN(n10783) );
  NAND2_X1 U13661 ( .A1(n12658), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n10782) );
  OAI211_X1 U13662 ( .C1(n10801), .C2(n10784), .A(n10783), .B(n10782), .ZN(
        n10785) );
  AOI21_X1 U13663 ( .B1(n10786), .B2(n11096), .A(n10785), .ZN(n14369) );
  XNOR2_X1 U13664 ( .A(n10818), .B(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15997) );
  INV_X1 U13665 ( .A(n15997), .ZN(n14917) );
  AOI22_X1 U13666 ( .A1(n10925), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n11085), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10791) );
  AOI22_X1 U13667 ( .A1(n11023), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n9831), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n10790) );
  AOI22_X1 U13668 ( .A1(n9862), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n9833), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10789) );
  AOI22_X1 U13669 ( .A1(n11079), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n11058), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n10788) );
  NAND4_X1 U13670 ( .A1(n10791), .A2(n10790), .A3(n10789), .A4(n10788), .ZN(
        n10797) );
  AOI22_X1 U13671 ( .A1(n11057), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n10499), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10795) );
  AOI22_X1 U13672 ( .A1(n11059), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n10481), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10794) );
  AOI22_X1 U13673 ( .A1(n9863), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n10930), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10793) );
  AOI22_X1 U13674 ( .A1(n11080), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n10597), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10792) );
  NAND4_X1 U13675 ( .A1(n10795), .A2(n10794), .A3(n10793), .A4(n10792), .ZN(
        n10796) );
  NOR2_X1 U13676 ( .A1(n10797), .A2(n10796), .ZN(n10800) );
  NAND2_X1 U13677 ( .A1(n11049), .A2(P1_EAX_REG_15__SCAN_IN), .ZN(n10799) );
  NAND2_X1 U13678 ( .A1(n12658), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n10798) );
  OAI211_X1 U13679 ( .C1(n10801), .C2(n10800), .A(n10799), .B(n10798), .ZN(
        n10802) );
  AOI21_X1 U13680 ( .B1(n14917), .B2(n11096), .A(n10802), .ZN(n14729) );
  INV_X1 U13681 ( .A(n13781), .ZN(n15072) );
  AOI22_X1 U13682 ( .A1(n11059), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10925), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10807) );
  AOI22_X1 U13683 ( .A1(n9831), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n9863), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10806) );
  AOI22_X1 U13684 ( .A1(n11023), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11057), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10805) );
  AOI22_X1 U13685 ( .A1(n11080), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n10597), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10804) );
  NAND4_X1 U13686 ( .A1(n10807), .A2(n10806), .A3(n10805), .A4(n10804), .ZN(
        n10813) );
  AOI22_X1 U13687 ( .A1(n9861), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(n9865), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10811) );
  AOI22_X1 U13688 ( .A1(n11085), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10481), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10810) );
  AOI22_X1 U13689 ( .A1(n10499), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n10908), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10809) );
  AOI22_X1 U13690 ( .A1(n11079), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11058), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10808) );
  NAND4_X1 U13691 ( .A1(n10811), .A2(n10810), .A3(n10809), .A4(n10808), .ZN(
        n10812) );
  NOR2_X1 U13692 ( .A1(n10813), .A2(n10812), .ZN(n10817) );
  NAND2_X1 U13693 ( .A1(n20802), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n10814) );
  NAND2_X1 U13694 ( .A1(n10609), .A2(n10814), .ZN(n10815) );
  AOI21_X1 U13695 ( .B1(n11049), .B2(P1_EAX_REG_16__SCAN_IN), .A(n10815), .ZN(
        n10816) );
  OAI21_X1 U13696 ( .B1(n11099), .B2(n10817), .A(n10816), .ZN(n10821) );
  OAI21_X1 U13697 ( .B1(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n10819), .A(
        n10837), .ZN(n16061) );
  OR2_X1 U13698 ( .A1(n10609), .A2(n16061), .ZN(n10820) );
  NAND2_X1 U13699 ( .A1(n10821), .A2(n10820), .ZN(n14722) );
  AOI22_X1 U13700 ( .A1(n10925), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n11085), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10825) );
  AOI22_X1 U13701 ( .A1(n11023), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n10499), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10824) );
  AOI22_X1 U13702 ( .A1(n9862), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n10481), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10823) );
  AOI22_X1 U13703 ( .A1(n9833), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n11064), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10822) );
  NAND4_X1 U13704 ( .A1(n10825), .A2(n10824), .A3(n10823), .A4(n10822), .ZN(
        n10831) );
  AOI22_X1 U13705 ( .A1(n9867), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n11080), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10829) );
  AOI22_X1 U13706 ( .A1(n11057), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n9863), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10828) );
  AOI22_X1 U13707 ( .A1(n11059), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n10597), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10827) );
  AOI22_X1 U13708 ( .A1(n9831), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n11058), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10826) );
  NAND4_X1 U13709 ( .A1(n10829), .A2(n10828), .A3(n10827), .A4(n10826), .ZN(
        n10830) );
  OR2_X1 U13710 ( .A1(n10831), .A2(n10830), .ZN(n10832) );
  NAND2_X1 U13711 ( .A1(n11074), .A2(n10832), .ZN(n10836) );
  XNOR2_X1 U13712 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B(n10837), .ZN(
        n14902) );
  NAND2_X1 U13713 ( .A1(n12658), .A2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n10833) );
  OAI21_X1 U13714 ( .B1(n14902), .B2(n10609), .A(n10833), .ZN(n10834) );
  AOI21_X1 U13715 ( .B1(n11049), .B2(P1_EAX_REG_17__SCAN_IN), .A(n10834), .ZN(
        n10835) );
  NAND2_X1 U13716 ( .A1(n10836), .A2(n10835), .ZN(n14626) );
  OR2_X1 U13717 ( .A1(n10838), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n10839) );
  NAND2_X1 U13718 ( .A1(n10839), .A2(n10871), .ZN(n16056) );
  AOI22_X1 U13719 ( .A1(n11023), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11065), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10843) );
  AOI22_X1 U13720 ( .A1(n11057), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n10499), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10842) );
  AOI22_X1 U13721 ( .A1(n11079), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n9861), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10841) );
  AOI22_X1 U13722 ( .A1(n10930), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n11058), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10840) );
  NAND4_X1 U13723 ( .A1(n10843), .A2(n10842), .A3(n10841), .A4(n10840), .ZN(
        n10849) );
  AOI22_X1 U13724 ( .A1(n10925), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11085), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10847) );
  AOI22_X1 U13725 ( .A1(n9863), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11080), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n10846) );
  AOI22_X1 U13726 ( .A1(n9833), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n10481), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10845) );
  AOI22_X1 U13727 ( .A1(n11059), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n10597), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10844) );
  NAND4_X1 U13728 ( .A1(n10847), .A2(n10846), .A3(n10845), .A4(n10844), .ZN(
        n10848) );
  NOR2_X1 U13729 ( .A1(n10849), .A2(n10848), .ZN(n10850) );
  NOR2_X1 U13730 ( .A1(n11099), .A2(n10850), .ZN(n10854) );
  INV_X1 U13731 ( .A(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n10852) );
  NAND2_X1 U13732 ( .A1(n11049), .A2(P1_EAX_REG_18__SCAN_IN), .ZN(n10851) );
  OAI211_X1 U13733 ( .C1(P1_STATE2_REG_2__SCAN_IN), .C2(n10852), .A(n10851), 
        .B(n10609), .ZN(n10853) );
  OAI22_X1 U13734 ( .A1(n16056), .A2(n10609), .B1(n10854), .B2(n10853), .ZN(
        n14710) );
  AOI22_X1 U13735 ( .A1(n11085), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n9862), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10858) );
  AOI22_X1 U13736 ( .A1(n11057), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n10499), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10857) );
  AOI22_X1 U13737 ( .A1(n11059), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n9833), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10856) );
  AOI22_X1 U13738 ( .A1(n11080), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n10597), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10855) );
  NAND4_X1 U13739 ( .A1(n10858), .A2(n10857), .A3(n10856), .A4(n10855), .ZN(
        n10864) );
  AOI22_X1 U13740 ( .A1(n11023), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n9863), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10862) );
  AOI22_X1 U13741 ( .A1(n10925), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n10481), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10861) );
  AOI22_X1 U13742 ( .A1(n9831), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10930), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10860) );
  AOI22_X1 U13743 ( .A1(n9867), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11058), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10859) );
  NAND4_X1 U13744 ( .A1(n10862), .A2(n10861), .A3(n10860), .A4(n10859), .ZN(
        n10863) );
  NOR2_X1 U13745 ( .A1(n10864), .A2(n10863), .ZN(n10868) );
  NAND2_X1 U13746 ( .A1(n20802), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n10865) );
  NAND2_X1 U13747 ( .A1(n10609), .A2(n10865), .ZN(n10866) );
  AOI21_X1 U13748 ( .B1(n11049), .B2(P1_EAX_REG_19__SCAN_IN), .A(n10866), .ZN(
        n10867) );
  OAI21_X1 U13749 ( .B1(n11099), .B2(n10868), .A(n10867), .ZN(n10870) );
  XNOR2_X1 U13750 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B(n10871), .ZN(
        n14619) );
  NAND2_X1 U13751 ( .A1(n11096), .A2(n14619), .ZN(n10869) );
  INV_X1 U13752 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n14616) );
  INV_X1 U13753 ( .A(n10906), .ZN(n10874) );
  OR2_X1 U13754 ( .A1(n10872), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n10873) );
  NAND2_X1 U13755 ( .A1(n10874), .A2(n10873), .ZN(n16048) );
  AOI22_X1 U13756 ( .A1(n9863), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11080), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n10878) );
  AOI22_X1 U13757 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n11023), .B1(
        n11057), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10877) );
  AOI22_X1 U13758 ( .A1(n10925), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n9833), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10876) );
  AOI22_X1 U13759 ( .A1(n11059), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n10597), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10875) );
  NAND4_X1 U13760 ( .A1(n10878), .A2(n10877), .A3(n10876), .A4(n10875), .ZN(
        n10884) );
  AOI22_X1 U13761 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n10499), .B1(
        n9831), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n10882) );
  AOI22_X1 U13762 ( .A1(n11079), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n9861), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10881) );
  AOI22_X1 U13763 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n11085), .B1(
        n10481), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10880) );
  AOI22_X1 U13764 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n10930), .B1(
        n11058), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10879) );
  NAND4_X1 U13765 ( .A1(n10882), .A2(n10881), .A3(n10880), .A4(n10879), .ZN(
        n10883) );
  NOR2_X1 U13766 ( .A1(n10884), .A2(n10883), .ZN(n10888) );
  NAND2_X1 U13767 ( .A1(n20802), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n10885) );
  NAND2_X1 U13768 ( .A1(n10609), .A2(n10885), .ZN(n10886) );
  AOI21_X1 U13769 ( .B1(n11049), .B2(P1_EAX_REG_20__SCAN_IN), .A(n10886), .ZN(
        n10887) );
  OAI21_X1 U13770 ( .B1(n11099), .B2(n10888), .A(n10887), .ZN(n10889) );
  OAI21_X1 U13771 ( .B1(n16048), .B2(n10609), .A(n10889), .ZN(n14705) );
  INV_X1 U13772 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n15972) );
  XNOR2_X1 U13773 ( .A(n10906), .B(n15972), .ZN(n15965) );
  NAND2_X1 U13774 ( .A1(n15965), .A2(n11096), .ZN(n10904) );
  AOI22_X1 U13775 ( .A1(n10925), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n9867), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10893) );
  AOI22_X1 U13776 ( .A1(n11023), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n9863), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10892) );
  AOI22_X1 U13777 ( .A1(n11057), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n10499), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10891) );
  AOI22_X1 U13778 ( .A1(n11065), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11058), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10890) );
  NAND4_X1 U13779 ( .A1(n10893), .A2(n10892), .A3(n10891), .A4(n10890), .ZN(
        n10899) );
  AOI22_X1 U13780 ( .A1(n9861), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(n9833), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10897) );
  AOI22_X1 U13781 ( .A1(n11080), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n10930), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10896) );
  AOI22_X1 U13782 ( .A1(n11085), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10481), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10895) );
  AOI22_X1 U13783 ( .A1(n11059), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10597), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10894) );
  NAND4_X1 U13784 ( .A1(n10897), .A2(n10896), .A3(n10895), .A4(n10894), .ZN(
        n10898) );
  NOR2_X1 U13785 ( .A1(n10899), .A2(n10898), .ZN(n10902) );
  AOI21_X1 U13786 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n15972), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n10900) );
  AOI21_X1 U13787 ( .B1(n11049), .B2(P1_EAX_REG_21__SCAN_IN), .A(n10900), .ZN(
        n10901) );
  OAI21_X1 U13788 ( .B1(n11099), .B2(n10902), .A(n10901), .ZN(n10903) );
  NAND2_X1 U13789 ( .A1(n10904), .A2(n10903), .ZN(n14696) );
  NAND2_X1 U13790 ( .A1(n14694), .A2(n10905), .ZN(n14691) );
  OAI21_X1 U13791 ( .B1(n10907), .B2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n10968), .ZN(n16043) );
  OR2_X1 U13792 ( .A1(n16043), .A2(n10609), .ZN(n10924) );
  AOI22_X1 U13793 ( .A1(n10925), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n11085), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10912) );
  AOI22_X1 U13794 ( .A1(n11023), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n9831), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10911) );
  AOI22_X1 U13795 ( .A1(n10335), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n10597), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10910) );
  AOI22_X1 U13796 ( .A1(n11080), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n10908), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10909) );
  NAND4_X1 U13797 ( .A1(n10912), .A2(n10911), .A3(n10910), .A4(n10909), .ZN(
        n10918) );
  AOI22_X1 U13798 ( .A1(n11057), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n10499), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10916) );
  AOI22_X1 U13799 ( .A1(n9867), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(n9833), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10915) );
  AOI22_X1 U13800 ( .A1(n9861), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n10481), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10914) );
  AOI22_X1 U13801 ( .A1(n9863), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11058), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10913) );
  NAND4_X1 U13802 ( .A1(n10916), .A2(n10915), .A3(n10914), .A4(n10913), .ZN(
        n10917) );
  NOR2_X1 U13803 ( .A1(n10918), .A2(n10917), .ZN(n10922) );
  NAND2_X1 U13804 ( .A1(n20802), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n10919) );
  NAND2_X1 U13805 ( .A1(n10609), .A2(n10919), .ZN(n10920) );
  AOI21_X1 U13806 ( .B1(n11049), .B2(P1_EAX_REG_22__SCAN_IN), .A(n10920), .ZN(
        n10921) );
  OAI21_X1 U13807 ( .B1(n11099), .B2(n10922), .A(n10921), .ZN(n10923) );
  NAND2_X1 U13808 ( .A1(n10924), .A2(n10923), .ZN(n14692) );
  AOI22_X1 U13809 ( .A1(n10925), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11085), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10929) );
  AOI22_X1 U13810 ( .A1(n11059), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n9833), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10928) );
  AOI22_X1 U13811 ( .A1(n10595), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n10481), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10927) );
  AOI22_X1 U13812 ( .A1(n11080), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n10597), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10926) );
  NAND4_X1 U13813 ( .A1(n10929), .A2(n10928), .A3(n10927), .A4(n10926), .ZN(
        n10936) );
  AOI22_X1 U13814 ( .A1(n11023), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n9863), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10934) );
  AOI22_X1 U13815 ( .A1(n11057), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n10499), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10933) );
  AOI22_X1 U13816 ( .A1(n9867), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11058), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10932) );
  AOI22_X1 U13817 ( .A1(n9831), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10930), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10931) );
  NAND4_X1 U13818 ( .A1(n10934), .A2(n10933), .A3(n10932), .A4(n10931), .ZN(
        n10935) );
  NOR2_X1 U13819 ( .A1(n10936), .A2(n10935), .ZN(n10952) );
  AOI22_X1 U13820 ( .A1(n11023), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11057), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10940) );
  AOI22_X1 U13821 ( .A1(n11059), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n9833), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10939) );
  AOI22_X1 U13822 ( .A1(n10925), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n10481), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10938) );
  AOI22_X1 U13823 ( .A1(n11080), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n10597), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10937) );
  NAND4_X1 U13824 ( .A1(n10940), .A2(n10939), .A3(n10938), .A4(n10937), .ZN(
        n10946) );
  AOI22_X1 U13825 ( .A1(n9863), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n10499), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10944) );
  AOI22_X1 U13826 ( .A1(n11085), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n9862), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10943) );
  AOI22_X1 U13827 ( .A1(n11065), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11064), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10942) );
  AOI22_X1 U13828 ( .A1(n9867), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11058), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n10941) );
  NAND4_X1 U13829 ( .A1(n10944), .A2(n10943), .A3(n10942), .A4(n10941), .ZN(
        n10945) );
  NOR2_X1 U13830 ( .A1(n10946), .A2(n10945), .ZN(n10953) );
  XNOR2_X1 U13831 ( .A(n10952), .B(n10953), .ZN(n10949) );
  INV_X1 U13832 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n15954) );
  OAI21_X1 U13833 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n15954), .A(n10609), 
        .ZN(n10947) );
  AOI21_X1 U13834 ( .B1(n11049), .B2(P1_EAX_REG_23__SCAN_IN), .A(n10947), .ZN(
        n10948) );
  OAI21_X1 U13835 ( .B1(n10949), .B2(n11099), .A(n10948), .ZN(n10951) );
  XNOR2_X1 U13836 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .B(n10968), .ZN(
        n15945) );
  NAND2_X1 U13837 ( .A1(n11096), .A2(n15945), .ZN(n10950) );
  AND2_X2 U13838 ( .A1(n14680), .A2(n14682), .ZN(n14674) );
  NOR2_X1 U13839 ( .A1(n10953), .A2(n10952), .ZN(n10975) );
  AOI22_X1 U13840 ( .A1(n11023), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n9863), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10957) );
  AOI22_X1 U13841 ( .A1(n11057), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n10499), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10956) );
  AOI22_X1 U13842 ( .A1(n9867), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11058), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10955) );
  AOI22_X1 U13843 ( .A1(n9831), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11064), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10954) );
  NAND4_X1 U13844 ( .A1(n10957), .A2(n10956), .A3(n10955), .A4(n10954), .ZN(
        n10963) );
  AOI22_X1 U13845 ( .A1(n10925), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n11085), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10961) );
  AOI22_X1 U13846 ( .A1(n11059), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n9833), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10960) );
  INV_X1 U13847 ( .A(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n20172) );
  AOI22_X1 U13848 ( .A1(n9862), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n10481), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10959) );
  AOI22_X1 U13849 ( .A1(n11080), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n10597), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10958) );
  NAND4_X1 U13850 ( .A1(n10961), .A2(n10960), .A3(n10959), .A4(n10958), .ZN(
        n10962) );
  OR2_X1 U13851 ( .A1(n10963), .A2(n10962), .ZN(n10974) );
  INV_X1 U13852 ( .A(n10974), .ZN(n10964) );
  XNOR2_X1 U13853 ( .A(n10975), .B(n10964), .ZN(n10965) );
  NAND2_X1 U13854 ( .A1(n10965), .A2(n11074), .ZN(n10973) );
  NAND2_X1 U13855 ( .A1(n20802), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n10966) );
  NAND2_X1 U13856 ( .A1(n10609), .A2(n10966), .ZN(n10967) );
  AOI21_X1 U13857 ( .B1(n11049), .B2(P1_EAX_REG_24__SCAN_IN), .A(n10967), .ZN(
        n10972) );
  OAI21_X1 U13858 ( .B1(n10970), .B2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n11011), .ZN(n15937) );
  NOR2_X1 U13859 ( .A1(n15937), .A2(n10609), .ZN(n10971) );
  AOI21_X1 U13860 ( .B1(n10973), .B2(n10972), .A(n10971), .ZN(n14675) );
  NAND2_X1 U13861 ( .A1(n10975), .A2(n10974), .ZN(n10993) );
  AOI22_X1 U13862 ( .A1(n11059), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n10925), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10979) );
  AOI22_X1 U13863 ( .A1(n11057), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n10499), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10978) );
  AOI22_X1 U13864 ( .A1(n11080), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n10597), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10977) );
  AOI22_X1 U13865 ( .A1(n11023), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11064), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10976) );
  NAND4_X1 U13866 ( .A1(n10979), .A2(n10978), .A3(n10977), .A4(n10976), .ZN(
        n10986) );
  AOI22_X1 U13867 ( .A1(n11065), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n9863), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10984) );
  AOI22_X1 U13868 ( .A1(n9861), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(n9833), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10983) );
  AOI22_X1 U13869 ( .A1(n11085), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n10481), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10982) );
  AOI22_X1 U13870 ( .A1(n11079), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11058), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10981) );
  NAND4_X1 U13871 ( .A1(n10984), .A2(n10983), .A3(n10982), .A4(n10981), .ZN(
        n10985) );
  NOR2_X1 U13872 ( .A1(n10986), .A2(n10985), .ZN(n10994) );
  XOR2_X1 U13873 ( .A(n10993), .B(n10994), .Z(n10987) );
  NAND2_X1 U13874 ( .A1(n10987), .A2(n11074), .ZN(n10990) );
  INV_X1 U13875 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n15924) );
  OAI21_X1 U13876 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n15924), .A(n10609), 
        .ZN(n10988) );
  AOI21_X1 U13877 ( .B1(n11049), .B2(P1_EAX_REG_25__SCAN_IN), .A(n10988), .ZN(
        n10989) );
  NAND2_X1 U13878 ( .A1(n10990), .A2(n10989), .ZN(n10992) );
  XNOR2_X1 U13879 ( .A(n11011), .B(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15927) );
  NAND2_X1 U13880 ( .A1(n15927), .A2(n11096), .ZN(n10991) );
  NAND2_X1 U13881 ( .A1(n10992), .A2(n10991), .ZN(n14668) );
  NOR2_X1 U13882 ( .A1(n10994), .A2(n10993), .ZN(n11018) );
  AOI22_X1 U13883 ( .A1(n11023), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n9863), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10998) );
  AOI22_X1 U13884 ( .A1(n11057), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n10499), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10997) );
  AOI22_X1 U13885 ( .A1(n9867), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11058), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10996) );
  AOI22_X1 U13886 ( .A1(n11065), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11064), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10995) );
  NAND4_X1 U13887 ( .A1(n10998), .A2(n10997), .A3(n10996), .A4(n10995), .ZN(
        n11004) );
  AOI22_X1 U13888 ( .A1(n10925), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11085), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11002) );
  AOI22_X1 U13889 ( .A1(n11059), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n9833), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11001) );
  AOI22_X1 U13890 ( .A1(n10595), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n10481), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11000) );
  INV_X1 U13891 ( .A(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n21145) );
  AOI22_X1 U13892 ( .A1(n11080), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10597), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10999) );
  NAND4_X1 U13893 ( .A1(n11002), .A2(n11001), .A3(n11000), .A4(n10999), .ZN(
        n11003) );
  OR2_X1 U13894 ( .A1(n11004), .A2(n11003), .ZN(n11017) );
  INV_X1 U13895 ( .A(n11017), .ZN(n11005) );
  XNOR2_X1 U13896 ( .A(n11018), .B(n11005), .ZN(n11008) );
  INV_X1 U13897 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n14596) );
  NAND2_X1 U13898 ( .A1(n11049), .A2(P1_EAX_REG_26__SCAN_IN), .ZN(n11006) );
  OAI211_X1 U13899 ( .C1(P1_STATE2_REG_2__SCAN_IN), .C2(n14596), .A(n11006), 
        .B(n10609), .ZN(n11007) );
  AOI21_X1 U13900 ( .B1(n11008), .B2(n11074), .A(n11007), .ZN(n11014) );
  INV_X1 U13901 ( .A(n11011), .ZN(n11009) );
  AOI21_X1 U13902 ( .B1(n11009), .B2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n11012) );
  NAND2_X1 U13903 ( .A1(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n11010) );
  OR2_X1 U13904 ( .A1(n11012), .A2(n11015), .ZN(n14851) );
  NOR2_X1 U13905 ( .A1(n14851), .A2(n10609), .ZN(n11013) );
  INV_X1 U13906 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n21108) );
  INV_X1 U13907 ( .A(n11015), .ZN(n11016) );
  AOI21_X1 U13908 ( .B1(n21108), .B2(n11016), .A(n11034), .ZN(n14845) );
  NAND2_X1 U13909 ( .A1(n11018), .A2(n11017), .ZN(n11037) );
  AOI22_X1 U13910 ( .A1(n10925), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n11085), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11022) );
  AOI22_X1 U13911 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n9833), .B1(
        n10481), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11021) );
  AOI22_X1 U13912 ( .A1(n11080), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11058), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11020) );
  AOI22_X1 U13913 ( .A1(n11059), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n10597), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11019) );
  NAND4_X1 U13914 ( .A1(n11022), .A2(n11021), .A3(n11020), .A4(n11019), .ZN(
        n11029) );
  AOI22_X1 U13915 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n11023), .B1(
        n9863), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11027) );
  AOI22_X1 U13916 ( .A1(n11057), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n10499), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11026) );
  AOI22_X1 U13917 ( .A1(n9867), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(n9862), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11025) );
  AOI22_X1 U13918 ( .A1(n9831), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11064), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11024) );
  NAND4_X1 U13919 ( .A1(n11027), .A2(n11026), .A3(n11025), .A4(n11024), .ZN(
        n11028) );
  NOR2_X1 U13920 ( .A1(n11029), .A2(n11028), .ZN(n11038) );
  XOR2_X1 U13921 ( .A(n11037), .B(n11038), .Z(n11032) );
  NAND2_X1 U13922 ( .A1(n11049), .A2(P1_EAX_REG_27__SCAN_IN), .ZN(n11030) );
  OAI211_X1 U13923 ( .C1(P1_STATE2_REG_2__SCAN_IN), .C2(n21108), .A(n11030), 
        .B(n10609), .ZN(n11031) );
  AOI21_X1 U13924 ( .B1(n11032), .B2(n11074), .A(n11031), .ZN(n11033) );
  INV_X1 U13925 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n14569) );
  NAND2_X1 U13926 ( .A1(n11035), .A2(n14569), .ZN(n11036) );
  NAND2_X1 U13927 ( .A1(n11054), .A2(n11036), .ZN(n14834) );
  NOR2_X1 U13928 ( .A1(n11038), .A2(n11037), .ZN(n11056) );
  AOI22_X1 U13929 ( .A1(n11023), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n9863), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11042) );
  AOI22_X1 U13930 ( .A1(n11057), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n10499), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11041) );
  AOI22_X1 U13931 ( .A1(n9867), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11058), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11040) );
  AOI22_X1 U13932 ( .A1(n11065), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11064), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11039) );
  NAND4_X1 U13933 ( .A1(n11042), .A2(n11041), .A3(n11040), .A4(n11039), .ZN(
        n11048) );
  AOI22_X1 U13934 ( .A1(n10925), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11085), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11046) );
  AOI22_X1 U13935 ( .A1(n11059), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n9833), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11045) );
  AOI22_X1 U13936 ( .A1(n9862), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n10481), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11044) );
  AOI22_X1 U13937 ( .A1(n11080), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n10597), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11043) );
  NAND4_X1 U13938 ( .A1(n11046), .A2(n11045), .A3(n11044), .A4(n11043), .ZN(
        n11047) );
  OR2_X1 U13939 ( .A1(n11048), .A2(n11047), .ZN(n11055) );
  XNOR2_X1 U13940 ( .A(n11056), .B(n11055), .ZN(n11052) );
  AOI21_X1 U13941 ( .B1(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n20802), .A(
        n11096), .ZN(n11051) );
  NAND2_X1 U13942 ( .A1(n11049), .A2(P1_EAX_REG_28__SCAN_IN), .ZN(n11050) );
  OAI211_X1 U13943 ( .C1(n11052), .C2(n11099), .A(n11051), .B(n11050), .ZN(
        n11053) );
  OAI21_X1 U13944 ( .B1(n10609), .B2(n14834), .A(n11053), .ZN(n14568) );
  XOR2_X1 U13945 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .B(n11077), .Z(
        n14513) );
  NAND2_X1 U13946 ( .A1(n11056), .A2(n11055), .ZN(n11092) );
  AOI22_X1 U13947 ( .A1(n11057), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n10499), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11063) );
  AOI22_X1 U13948 ( .A1(n11085), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n10481), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11062) );
  AOI22_X1 U13949 ( .A1(n11080), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11058), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11061) );
  AOI22_X1 U13950 ( .A1(n11059), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n10597), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11060) );
  NAND4_X1 U13951 ( .A1(n11063), .A2(n11062), .A3(n11061), .A4(n11060), .ZN(
        n11071) );
  AOI22_X1 U13952 ( .A1(n10925), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n9861), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11069) );
  AOI22_X1 U13953 ( .A1(n11023), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n9863), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11068) );
  AOI22_X1 U13954 ( .A1(n11079), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n9833), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11067) );
  AOI22_X1 U13955 ( .A1(n9831), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11064), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11066) );
  NAND4_X1 U13956 ( .A1(n11069), .A2(n11068), .A3(n11067), .A4(n11066), .ZN(
        n11070) );
  NOR2_X1 U13957 ( .A1(n11071), .A2(n11070), .ZN(n11093) );
  XOR2_X1 U13958 ( .A(n11092), .B(n11093), .Z(n11075) );
  INV_X1 U13959 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n12664) );
  NAND2_X1 U13960 ( .A1(n11049), .A2(P1_EAX_REG_29__SCAN_IN), .ZN(n11072) );
  OAI211_X1 U13961 ( .C1(P1_STATE2_REG_2__SCAN_IN), .C2(n12664), .A(n11072), 
        .B(n10609), .ZN(n11073) );
  AOI21_X1 U13962 ( .B1(n11075), .B2(n11074), .A(n11073), .ZN(n11076) );
  XOR2_X1 U13963 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .B(n11172), .Z(
        n14822) );
  AOI22_X1 U13964 ( .A1(n11057), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n10499), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11084) );
  AOI22_X1 U13965 ( .A1(n10335), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n9833), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11083) );
  AOI22_X1 U13966 ( .A1(n11079), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11078), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11082) );
  AOI22_X1 U13967 ( .A1(n11080), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n10597), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11081) );
  NAND4_X1 U13968 ( .A1(n11084), .A2(n11083), .A3(n11082), .A4(n11081), .ZN(
        n11091) );
  AOI22_X1 U13969 ( .A1(n10925), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11085), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11089) );
  AOI22_X1 U13970 ( .A1(n11023), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n9863), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11088) );
  AOI22_X1 U13971 ( .A1(n10595), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n10481), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11087) );
  AOI22_X1 U13972 ( .A1(n11065), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11058), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11086) );
  NAND4_X1 U13973 ( .A1(n11089), .A2(n11088), .A3(n11087), .A4(n11086), .ZN(
        n11090) );
  NOR2_X1 U13974 ( .A1(n11091), .A2(n11090), .ZN(n11095) );
  NOR2_X1 U13975 ( .A1(n11093), .A2(n11092), .ZN(n11094) );
  XOR2_X1 U13976 ( .A(n11095), .B(n11094), .Z(n11100) );
  AOI21_X1 U13977 ( .B1(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n20802), .A(
        n11096), .ZN(n11098) );
  NAND2_X1 U13978 ( .A1(n11049), .A2(P1_EAX_REG_30__SCAN_IN), .ZN(n11097) );
  OAI211_X1 U13979 ( .C1(n11100), .C2(n11099), .A(n11098), .B(n11097), .ZN(
        n11101) );
  OAI21_X1 U13980 ( .B1(n10609), .B2(n14822), .A(n11101), .ZN(n14558) );
  AOI22_X1 U13981 ( .A1(n11049), .A2(P1_EAX_REG_31__SCAN_IN), .B1(n12658), 
        .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n11102) );
  XNOR2_X2 U13982 ( .A(n14556), .B(n11102), .ZN(n14506) );
  NAND2_X1 U13983 ( .A1(n20790), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11114) );
  OAI21_X1 U13984 ( .B1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n20790), .A(
        n11114), .ZN(n11103) );
  INV_X1 U13985 ( .A(n11103), .ZN(n11108) );
  NAND2_X1 U13986 ( .A1(n11155), .A2(n11108), .ZN(n11104) );
  NAND2_X1 U13987 ( .A1(n11156), .A2(n11104), .ZN(n11111) );
  INV_X1 U13988 ( .A(n11106), .ZN(n11109) );
  NAND2_X1 U13989 ( .A1(n10418), .A2(n9854), .ZN(n11107) );
  NAND2_X1 U13990 ( .A1(n11107), .A2(n20168), .ZN(n11129) );
  OAI211_X1 U13991 ( .C1(n11105), .C2(n11109), .A(n11129), .B(n11108), .ZN(
        n11110) );
  NAND2_X1 U13992 ( .A1(n11111), .A2(n11110), .ZN(n11117) );
  NOR2_X1 U13993 ( .A1(n11112), .A2(n20806), .ZN(n11113) );
  MUX2_X1 U13994 ( .A(n20523), .B(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .S(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .Z(n11120) );
  XNOR2_X1 U13995 ( .A(n11120), .B(n11119), .ZN(n11164) );
  NAND2_X1 U13996 ( .A1(n11115), .A2(n9858), .ZN(n11146) );
  OAI211_X1 U13997 ( .C1(n11117), .C2(n11115), .A(n11164), .B(n11146), .ZN(
        n11127) );
  INV_X1 U13998 ( .A(n11115), .ZN(n11116) );
  NOR2_X1 U13999 ( .A1(n11164), .A2(n11116), .ZN(n11118) );
  NAND2_X1 U14000 ( .A1(n11118), .A2(n11117), .ZN(n11126) );
  NAND2_X1 U14001 ( .A1(n11120), .A2(n11119), .ZN(n11122) );
  NAND2_X1 U14002 ( .A1(n20523), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11121) );
  NAND2_X1 U14003 ( .A1(n11122), .A2(n11121), .ZN(n11133) );
  XNOR2_X1 U14004 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n11132) );
  XNOR2_X1 U14005 ( .A(n11133), .B(n11132), .ZN(n11163) );
  INV_X1 U14006 ( .A(n11163), .ZN(n11123) );
  NAND2_X1 U14007 ( .A1(n11155), .A2(n11123), .ZN(n11128) );
  NAND2_X1 U14008 ( .A1(n11147), .A2(n11163), .ZN(n11124) );
  NAND3_X1 U14009 ( .A1(n11128), .A2(n11129), .A3(n11124), .ZN(n11125) );
  NAND3_X1 U14010 ( .A1(n11127), .A2(n11126), .A3(n11125), .ZN(n11138) );
  INV_X1 U14011 ( .A(n11128), .ZN(n11131) );
  INV_X1 U14012 ( .A(n11129), .ZN(n11130) );
  NAND2_X1 U14013 ( .A1(n11131), .A2(n11130), .ZN(n11137) );
  INV_X1 U14014 ( .A(n11147), .ZN(n11136) );
  NAND2_X1 U14015 ( .A1(n11133), .A2(n11132), .ZN(n11135) );
  NAND2_X1 U14016 ( .A1(n20461), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11134) );
  NAND2_X1 U14017 ( .A1(n11135), .A2(n11134), .ZN(n11142) );
  XNOR2_X1 U14018 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n11141) );
  XNOR2_X1 U14019 ( .A(n11142), .B(n11141), .ZN(n11165) );
  AOI22_X1 U14020 ( .A1(n11138), .A2(n11137), .B1(n11136), .B2(n11165), .ZN(
        n11145) );
  INV_X1 U14021 ( .A(n11165), .ZN(n11139) );
  NOR2_X1 U14022 ( .A1(n11156), .A2(n11139), .ZN(n11144) );
  NOR2_X1 U14023 ( .A1(n10581), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n11140) );
  NOR2_X1 U14024 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n20152), .ZN(
        n11152) );
  INV_X1 U14025 ( .A(n11166), .ZN(n11143) );
  OAI22_X1 U14026 ( .A1(n11145), .A2(n11144), .B1(n11147), .B2(n11143), .ZN(
        n11151) );
  INV_X1 U14027 ( .A(n11146), .ZN(n11149) );
  AOI22_X1 U14028 ( .A1(n11149), .A2(n11148), .B1(
        P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n20806), .ZN(n11150) );
  NAND2_X1 U14029 ( .A1(n11151), .A2(n11150), .ZN(n11158) );
  NAND2_X1 U14030 ( .A1(n20152), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n11153) );
  INV_X1 U14031 ( .A(n13492), .ZN(n11168) );
  NAND2_X1 U14032 ( .A1(n11158), .A2(n11168), .ZN(n11159) );
  NOR4_X1 U14033 ( .A1(n11166), .A2(n11165), .A3(n11164), .A4(n11163), .ZN(
        n13491) );
  INV_X1 U14034 ( .A(n13491), .ZN(n11167) );
  AND3_X1 U14035 ( .A1(n11162), .A2(n11168), .A3(n11167), .ZN(n13480) );
  NAND2_X1 U14036 ( .A1(n13480), .A2(n13736), .ZN(n14548) );
  INV_X2 U14037 ( .A(n20128), .ZN(n20103) );
  NAND2_X1 U14038 ( .A1(n20802), .A2(n13782), .ZN(n20807) );
  NOR2_X1 U14039 ( .A1(n20413), .A2(n20807), .ZN(n15902) );
  INV_X1 U14040 ( .A(n15902), .ZN(n15898) );
  OR2_X1 U14041 ( .A1(n10609), .A2(n13782), .ZN(n11169) );
  MUX2_X1 U14042 ( .A(n15898), .B(n11169), .S(n20806), .Z(n11170) );
  INV_X1 U14043 ( .A(n11170), .ZN(n11171) );
  INV_X1 U14044 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n14560) );
  INV_X1 U14045 ( .A(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n11283) );
  NAND2_X1 U14046 ( .A1(n14506), .A2(n19992), .ZN(n11291) );
  AOI22_X1 U14047 ( .A1(n13396), .A2(P1_EBX_REG_30__SCAN_IN), .B1(n13820), 
        .B2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14553) );
  INV_X1 U14048 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n20151) );
  NAND2_X1 U14049 ( .A1(n11197), .A2(n20151), .ZN(n11177) );
  INV_X1 U14050 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n13963) );
  NAND2_X1 U14051 ( .A1(n13808), .A2(n13963), .ZN(n11176) );
  NAND3_X1 U14052 ( .A1(n11177), .A2(n11250), .A3(n11176), .ZN(n11178) );
  NAND2_X1 U14053 ( .A1(n11197), .A2(P1_EBX_REG_0__SCAN_IN), .ZN(n11182) );
  INV_X1 U14054 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n14656) );
  NAND2_X1 U14055 ( .A1(n9835), .A2(n14656), .ZN(n11181) );
  NAND2_X1 U14056 ( .A1(n11182), .A2(n11181), .ZN(n13397) );
  XNOR2_X1 U14057 ( .A(n11183), .B(n13397), .ZN(n13819) );
  NAND2_X1 U14058 ( .A1(n13819), .A2(n13808), .ZN(n13822) );
  NAND2_X1 U14059 ( .A1(n13822), .A2(n11183), .ZN(n13814) );
  OR2_X1 U14060 ( .A1(n9860), .A2(P1_EBX_REG_2__SCAN_IN), .ZN(n11188) );
  INV_X1 U14061 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n20135) );
  NAND2_X1 U14062 ( .A1(n11197), .A2(n20135), .ZN(n11186) );
  INV_X1 U14063 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n13816) );
  NAND2_X1 U14064 ( .A1(n13808), .A2(n13816), .ZN(n11185) );
  NAND3_X1 U14065 ( .A1(n11186), .A2(n9835), .A3(n11185), .ZN(n11187) );
  AND2_X1 U14066 ( .A1(n11188), .A2(n11187), .ZN(n13813) );
  NAND2_X2 U14067 ( .A1(n13808), .A2(n9835), .ZN(n11258) );
  MUX2_X1 U14068 ( .A(n11258), .B(n9835), .S(P1_EBX_REG_3__SCAN_IN), .Z(n11190) );
  OR2_X1 U14069 ( .A1(n13396), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11189) );
  MUX2_X1 U14070 ( .A(n9860), .B(n11197), .S(P1_EBX_REG_4__SCAN_IN), .Z(n11192) );
  NAND2_X1 U14071 ( .A1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n13820), .ZN(
        n11191) );
  INV_X1 U14072 ( .A(P1_EBX_REG_5__SCAN_IN), .ZN(n19998) );
  NAND2_X1 U14073 ( .A1(n13808), .A2(n19998), .ZN(n11194) );
  NAND2_X1 U14074 ( .A1(n9835), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11193) );
  NAND3_X1 U14075 ( .A1(n11194), .A2(n11197), .A3(n11193), .ZN(n11195) );
  OAI21_X1 U14076 ( .B1(n11258), .B2(P1_EBX_REG_5__SCAN_IN), .A(n11195), .ZN(
        n13943) );
  MUX2_X1 U14077 ( .A(n9860), .B(n11197), .S(P1_EBX_REG_6__SCAN_IN), .Z(n11199) );
  NAND2_X1 U14078 ( .A1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n13820), .ZN(
        n11198) );
  NOR2_X2 U14079 ( .A1(n13997), .A2(n13996), .ZN(n13998) );
  INV_X1 U14080 ( .A(n11258), .ZN(n11200) );
  INV_X1 U14081 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n13993) );
  NAND2_X1 U14082 ( .A1(n11200), .A2(n13993), .ZN(n11204) );
  NAND2_X1 U14083 ( .A1(n13808), .A2(n13993), .ZN(n11202) );
  NAND2_X1 U14084 ( .A1(n9835), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11201) );
  NAND3_X1 U14085 ( .A1(n11202), .A2(n11197), .A3(n11201), .ZN(n11203) );
  MUX2_X1 U14086 ( .A(n9860), .B(n11197), .S(P1_EBX_REG_8__SCAN_IN), .Z(n11207) );
  NAND2_X1 U14087 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n13820), .ZN(
        n11205) );
  AND2_X1 U14088 ( .A1(n11243), .A2(n11205), .ZN(n11206) );
  NAND2_X1 U14089 ( .A1(n11207), .A2(n11206), .ZN(n14075) );
  INV_X1 U14090 ( .A(P1_EBX_REG_9__SCAN_IN), .ZN(n11208) );
  NAND2_X1 U14091 ( .A1(n13808), .A2(n11208), .ZN(n11210) );
  NAND2_X1 U14092 ( .A1(n9835), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n11209) );
  NAND3_X1 U14093 ( .A1(n11210), .A2(n11197), .A3(n11209), .ZN(n11211) );
  OAI21_X1 U14094 ( .B1(n11258), .B2(P1_EBX_REG_9__SCAN_IN), .A(n11211), .ZN(
        n14205) );
  OR2_X1 U14095 ( .A1(n9860), .A2(P1_EBX_REG_10__SCAN_IN), .ZN(n11215) );
  NAND2_X1 U14096 ( .A1(n11197), .A2(n16080), .ZN(n11213) );
  INV_X1 U14097 ( .A(P1_EBX_REG_10__SCAN_IN), .ZN(n16029) );
  NAND2_X1 U14098 ( .A1(n13808), .A2(n16029), .ZN(n11212) );
  NAND3_X1 U14099 ( .A1(n11213), .A2(n9835), .A3(n11212), .ZN(n11214) );
  MUX2_X1 U14100 ( .A(n11258), .B(n9835), .S(P1_EBX_REG_11__SCAN_IN), .Z(
        n11216) );
  OAI21_X1 U14101 ( .B1(n13396), .B2(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n11216), .ZN(n14308) );
  MUX2_X1 U14102 ( .A(n9860), .B(n11197), .S(P1_EBX_REG_12__SCAN_IN), .Z(
        n11218) );
  NAND2_X1 U14103 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n13820), .ZN(
        n11217) );
  MUX2_X1 U14104 ( .A(n11258), .B(n9835), .S(P1_EBX_REG_13__SCAN_IN), .Z(
        n11219) );
  OAI21_X1 U14105 ( .B1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n13396), .A(
        n11219), .ZN(n14644) );
  OR2_X1 U14106 ( .A1(n9860), .A2(P1_EBX_REG_14__SCAN_IN), .ZN(n11224) );
  INV_X1 U14107 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n16143) );
  NAND2_X1 U14108 ( .A1(n11197), .A2(n16143), .ZN(n11222) );
  INV_X1 U14109 ( .A(P1_EBX_REG_14__SCAN_IN), .ZN(n16005) );
  NAND2_X1 U14110 ( .A1(n13808), .A2(n16005), .ZN(n11221) );
  NAND3_X1 U14111 ( .A1(n11222), .A2(n9835), .A3(n11221), .ZN(n11223) );
  MUX2_X1 U14112 ( .A(n11258), .B(n11250), .S(P1_EBX_REG_15__SCAN_IN), .Z(
        n11225) );
  OAI21_X1 U14113 ( .B1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n13396), .A(
        n11225), .ZN(n11226) );
  INV_X1 U14114 ( .A(n11226), .ZN(n14732) );
  OR2_X1 U14115 ( .A1(n9860), .A2(P1_EBX_REG_16__SCAN_IN), .ZN(n11230) );
  INV_X1 U14116 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15047) );
  NAND2_X1 U14117 ( .A1(n11197), .A2(n15047), .ZN(n11228) );
  INV_X1 U14118 ( .A(P1_EBX_REG_16__SCAN_IN), .ZN(n14726) );
  NAND2_X1 U14119 ( .A1(n13808), .A2(n14726), .ZN(n11227) );
  NAND3_X1 U14120 ( .A1(n11228), .A2(n9835), .A3(n11227), .ZN(n11229) );
  NAND2_X1 U14121 ( .A1(n11230), .A2(n11229), .ZN(n14723) );
  MUX2_X1 U14122 ( .A(n11258), .B(n9835), .S(P1_EBX_REG_17__SCAN_IN), .Z(
        n11231) );
  OAI21_X1 U14123 ( .B1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n13396), .A(
        n11231), .ZN(n14630) );
  OR2_X1 U14124 ( .A1(n9860), .A2(P1_EBX_REG_18__SCAN_IN), .ZN(n11235) );
  INV_X1 U14125 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n16123) );
  NAND2_X1 U14126 ( .A1(n11197), .A2(n16123), .ZN(n11233) );
  INV_X1 U14127 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n15981) );
  NAND2_X1 U14128 ( .A1(n13808), .A2(n15981), .ZN(n11232) );
  NAND3_X1 U14129 ( .A1(n11233), .A2(n9835), .A3(n11232), .ZN(n11234) );
  MUX2_X1 U14130 ( .A(n11258), .B(n9835), .S(P1_EBX_REG_19__SCAN_IN), .Z(
        n11237) );
  OR2_X1 U14131 ( .A1(n13396), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n11236) );
  AND2_X1 U14132 ( .A1(n11237), .A2(n11236), .ZN(n14617) );
  MUX2_X1 U14133 ( .A(n9860), .B(n11197), .S(P1_EBX_REG_20__SCAN_IN), .Z(
        n11240) );
  NAND2_X1 U14134 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n13820), .ZN(
        n11238) );
  AND2_X1 U14135 ( .A1(n11243), .A2(n11238), .ZN(n11239) );
  NAND2_X1 U14136 ( .A1(n11240), .A2(n11239), .ZN(n14702) );
  NAND2_X1 U14137 ( .A1(n14703), .A2(n14702), .ZN(n14697) );
  MUX2_X1 U14138 ( .A(n11258), .B(n9835), .S(P1_EBX_REG_21__SCAN_IN), .Z(
        n11241) );
  OAI21_X1 U14139 ( .B1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .B2(n13396), .A(
        n11241), .ZN(n14698) );
  MUX2_X1 U14140 ( .A(n9860), .B(n11197), .S(P1_EBX_REG_22__SCAN_IN), .Z(
        n11244) );
  NAND2_X1 U14141 ( .A1(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n13820), .ZN(
        n11242) );
  AND3_X1 U14142 ( .A1(n11244), .A2(n11243), .A3(n11242), .ZN(n14688) );
  MUX2_X1 U14143 ( .A(n11258), .B(n11250), .S(P1_EBX_REG_23__SCAN_IN), .Z(
        n11245) );
  OAI21_X1 U14144 ( .B1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n13396), .A(
        n11245), .ZN(n14684) );
  OR2_X1 U14145 ( .A1(n9860), .A2(P1_EBX_REG_24__SCAN_IN), .ZN(n11249) );
  INV_X1 U14146 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14999) );
  NAND2_X1 U14147 ( .A1(n11197), .A2(n14999), .ZN(n11247) );
  INV_X1 U14148 ( .A(P1_EBX_REG_24__SCAN_IN), .ZN(n15936) );
  NAND2_X1 U14149 ( .A1(n13808), .A2(n15936), .ZN(n11246) );
  NAND3_X1 U14150 ( .A1(n11247), .A2(n9835), .A3(n11246), .ZN(n11248) );
  NAND2_X1 U14151 ( .A1(n11249), .A2(n11248), .ZN(n14676) );
  INV_X1 U14152 ( .A(P1_EBX_REG_25__SCAN_IN), .ZN(n20935) );
  NAND2_X1 U14153 ( .A1(n13808), .A2(n20935), .ZN(n11252) );
  NAND2_X1 U14154 ( .A1(n9835), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n11251) );
  NAND3_X1 U14155 ( .A1(n11252), .A2(n9958), .A3(n11251), .ZN(n11253) );
  OAI21_X1 U14156 ( .B1(n11258), .B2(P1_EBX_REG_25__SCAN_IN), .A(n11253), .ZN(
        n14671) );
  NOR2_X2 U14157 ( .A1(n14670), .A2(n14671), .ZN(n14598) );
  OR2_X1 U14158 ( .A1(n9860), .A2(P1_EBX_REG_26__SCAN_IN), .ZN(n11257) );
  INV_X1 U14159 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n21089) );
  INV_X1 U14160 ( .A(P1_EBX_REG_26__SCAN_IN), .ZN(n14666) );
  NAND2_X1 U14161 ( .A1(n13808), .A2(n14666), .ZN(n11254) );
  NAND3_X1 U14162 ( .A1(n11255), .A2(n9835), .A3(n11254), .ZN(n11256) );
  NAND2_X1 U14163 ( .A1(n11257), .A2(n11256), .ZN(n14597) );
  NAND2_X1 U14164 ( .A1(n14598), .A2(n14597), .ZN(n14583) );
  MUX2_X1 U14165 ( .A(n11258), .B(n9835), .S(P1_EBX_REG_27__SCAN_IN), .Z(
        n11259) );
  OAI21_X1 U14166 ( .B1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n13396), .A(
        n11259), .ZN(n14584) );
  OR2_X2 U14167 ( .A1(n14583), .A2(n14584), .ZN(n14586) );
  OR2_X1 U14168 ( .A1(n9860), .A2(P1_EBX_REG_28__SCAN_IN), .ZN(n11263) );
  INV_X1 U14169 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n14831) );
  NAND2_X1 U14170 ( .A1(n11197), .A2(n14831), .ZN(n11261) );
  INV_X1 U14171 ( .A(P1_EBX_REG_28__SCAN_IN), .ZN(n14664) );
  NAND2_X1 U14172 ( .A1(n13808), .A2(n14664), .ZN(n11260) );
  NAND3_X1 U14173 ( .A1(n11261), .A2(n9835), .A3(n11260), .ZN(n11262) );
  AND2_X1 U14174 ( .A1(n11263), .A2(n11262), .ZN(n14570) );
  OR2_X2 U14175 ( .A1(n14586), .A2(n14570), .ZN(n14571) );
  OR2_X1 U14176 ( .A1(n13396), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n11265) );
  INV_X1 U14177 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n11264) );
  NAND2_X1 U14178 ( .A1(n9846), .A2(n11264), .ZN(n11266) );
  NAND2_X1 U14179 ( .A1(n11265), .A2(n11266), .ZN(n14551) );
  MUX2_X1 U14180 ( .A(n14551), .B(n11266), .S(n13477), .Z(n14510) );
  MUX2_X1 U14181 ( .A(n9835), .B(n14553), .S(n14552), .Z(n11268) );
  AOI22_X1 U14182 ( .A1(n13396), .A2(P1_EBX_REG_31__SCAN_IN), .B1(n13820), 
        .B2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n11267) );
  AND2_X1 U14183 ( .A1(n9854), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n11269) );
  NAND2_X1 U14184 ( .A1(READY1), .A2(READY11_REG_SCAN_IN), .ZN(n20810) );
  AND2_X1 U14185 ( .A1(n20810), .A2(n20208), .ZN(n15890) );
  NAND2_X1 U14186 ( .A1(n10421), .A2(P1_EBX_REG_31__SCAN_IN), .ZN(n11278) );
  AND2_X1 U14187 ( .A1(P1_REIP_REG_29__SCAN_IN), .A2(P1_REIP_REG_30__SCAN_IN), 
        .ZN(n11277) );
  OR2_X1 U14188 ( .A1(n11270), .A2(P1_STATE_REG_0__SCAN_IN), .ZN(n13727) );
  INV_X1 U14189 ( .A(n20810), .ZN(n20701) );
  AOI21_X1 U14190 ( .B1(n20168), .B2(n13727), .A(n20701), .ZN(n13372) );
  NAND2_X1 U14191 ( .A1(n13372), .A2(n20208), .ZN(n11279) );
  NAND2_X1 U14192 ( .A1(n20023), .A2(n20022), .ZN(n14613) );
  AND2_X1 U14193 ( .A1(P1_REIP_REG_27__SCAN_IN), .A2(P1_REIP_REG_28__SCAN_IN), 
        .ZN(n11287) );
  INV_X1 U14194 ( .A(n11287), .ZN(n11276) );
  INV_X1 U14195 ( .A(n20022), .ZN(n19979) );
  NAND4_X1 U14196 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(P1_REIP_REG_1__SCAN_IN), 
        .A3(P1_REIP_REG_3__SCAN_IN), .A4(P1_REIP_REG_2__SCAN_IN), .ZN(n19980)
         );
  NAND4_X1 U14197 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(P1_REIP_REG_7__SCAN_IN), 
        .A3(P1_REIP_REG_6__SCAN_IN), .A4(P1_REIP_REG_5__SCAN_IN), .ZN(n11284)
         );
  NOR3_X1 U14198 ( .A1(n19979), .A2(n19980), .A3(n11284), .ZN(n14611) );
  NAND4_X1 U14199 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(P1_REIP_REG_13__SCAN_IN), 
        .A3(P1_REIP_REG_12__SCAN_IN), .A4(P1_REIP_REG_11__SCAN_IN), .ZN(n14610) );
  NAND3_X1 U14200 ( .A1(P1_REIP_REG_17__SCAN_IN), .A2(P1_REIP_REG_16__SCAN_IN), 
        .A3(P1_REIP_REG_15__SCAN_IN), .ZN(n14614) );
  NAND2_X1 U14201 ( .A1(P1_REIP_REG_19__SCAN_IN), .A2(P1_REIP_REG_18__SCAN_IN), 
        .ZN(n15975) );
  NAND3_X1 U14202 ( .A1(P1_REIP_REG_20__SCAN_IN), .A2(P1_REIP_REG_9__SCAN_IN), 
        .A3(P1_REIP_REG_10__SCAN_IN), .ZN(n11271) );
  NOR4_X1 U14203 ( .A1(n14610), .A2(n14614), .A3(n15975), .A4(n11271), .ZN(
        n15961) );
  AND4_X1 U14204 ( .A1(P1_REIP_REG_23__SCAN_IN), .A2(n15961), .A3(
        P1_REIP_REG_22__SCAN_IN), .A4(P1_REIP_REG_21__SCAN_IN), .ZN(n11272) );
  NAND2_X1 U14205 ( .A1(n14611), .A2(n11272), .ZN(n11273) );
  NAND2_X1 U14206 ( .A1(n11273), .A2(n14613), .ZN(n15946) );
  AND3_X1 U14207 ( .A1(P1_REIP_REG_24__SCAN_IN), .A2(P1_REIP_REG_25__SCAN_IN), 
        .A3(P1_REIP_REG_26__SCAN_IN), .ZN(n11286) );
  INV_X1 U14208 ( .A(n11286), .ZN(n11274) );
  NAND2_X1 U14209 ( .A1(n14613), .A2(n11274), .ZN(n11275) );
  NAND2_X1 U14210 ( .A1(n15946), .A2(n11275), .ZN(n14601) );
  AOI21_X1 U14211 ( .B1(n11276), .B2(n14613), .A(n14601), .ZN(n14579) );
  OAI21_X1 U14212 ( .B1(n11277), .B2(n16020), .A(n14579), .ZN(n14563) );
  INV_X1 U14213 ( .A(n11278), .ZN(n11281) );
  INV_X1 U14214 ( .A(n11279), .ZN(n11280) );
  INV_X1 U14215 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n14662) );
  OAI22_X1 U14216 ( .A1(n20014), .A2(n11283), .B1(n19997), .B2(n14662), .ZN(
        n11289) );
  NAND2_X1 U14217 ( .A1(n19970), .A2(n15961), .ZN(n15959) );
  NAND2_X1 U14218 ( .A1(P1_REIP_REG_22__SCAN_IN), .A2(P1_REIP_REG_21__SCAN_IN), 
        .ZN(n11285) );
  NOR2_X1 U14219 ( .A1(n15959), .A2(n11285), .ZN(n15950) );
  NAND2_X1 U14220 ( .A1(n14592), .A2(n11287), .ZN(n14559) );
  INV_X1 U14221 ( .A(P1_REIP_REG_30__SCAN_IN), .ZN(n14820) );
  INV_X1 U14222 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n20751) );
  NOR4_X1 U14223 ( .A1(n14559), .A2(P1_REIP_REG_31__SCAN_IN), .A3(n14820), 
        .A4(n20751), .ZN(n11288) );
  AOI211_X1 U14224 ( .C1(P1_REIP_REG_31__SCAN_IN), .C2(n14563), .A(n11289), 
        .B(n11288), .ZN(n11290) );
  NAND2_X1 U14225 ( .A1(n11326), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11323) );
  NAND2_X1 U14226 ( .A1(n11324), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n11321) );
  NAND2_X1 U14227 ( .A1(n11318), .A2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n11319) );
  INV_X1 U14228 ( .A(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n11332) );
  AND2_X1 U14229 ( .A1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n11292) );
  NAND2_X1 U14230 ( .A1(n11311), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n11310) );
  INV_X1 U14231 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n15343) );
  NAND2_X1 U14232 ( .A1(n11309), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n11307) );
  INV_X1 U14233 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n15322) );
  INV_X1 U14234 ( .A(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n16210) );
  NAND2_X1 U14235 ( .A1(n11304), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11306) );
  INV_X1 U14236 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n15304) );
  NOR2_X1 U14237 ( .A1(n11294), .A2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n11295) );
  OR2_X1 U14238 ( .A1(n11296), .A2(n11295), .ZN(n15289) );
  INV_X1 U14239 ( .A(n15289), .ZN(n11336) );
  INV_X1 U14240 ( .A(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n11297) );
  INV_X1 U14241 ( .A(n12991), .ZN(n11299) );
  NAND2_X1 U14242 ( .A1(n11299), .A2(n13537), .ZN(n11301) );
  INV_X1 U14243 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n20998) );
  NOR2_X1 U14244 ( .A1(n11302), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n11303) );
  OR2_X1 U14245 ( .A1(n11294), .A2(n11303), .ZN(n12325) );
  INV_X1 U14246 ( .A(n12325), .ZN(n15105) );
  AOI21_X1 U14247 ( .B1(n15304), .B2(n11306), .A(n11302), .ZN(n15302) );
  INV_X1 U14248 ( .A(n11304), .ZN(n11308) );
  NAND2_X1 U14249 ( .A1(n11308), .A2(n16210), .ZN(n11305) );
  NAND2_X1 U14250 ( .A1(n11306), .A2(n11305), .ZN(n15313) );
  INV_X1 U14251 ( .A(n15313), .ZN(n16218) );
  AOI21_X1 U14252 ( .B1(n15322), .B2(n11307), .A(n11304), .ZN(n15324) );
  OAI21_X1 U14253 ( .B1(n11309), .B2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n11307), .ZN(n15335) );
  INV_X1 U14254 ( .A(n15335), .ZN(n15137) );
  AOI21_X1 U14255 ( .B1(n15343), .B2(n11310), .A(n11309), .ZN(n15345) );
  OAI21_X1 U14256 ( .B1(n11311), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n11310), .ZN(n15357) );
  INV_X1 U14257 ( .A(n15357), .ZN(n15858) );
  AOI21_X1 U14258 ( .B1(n11312), .B2(n11293), .A(n11311), .ZN(n15378) );
  OAI21_X1 U14259 ( .B1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n11313), .A(
        n11312), .ZN(n11314) );
  INV_X1 U14260 ( .A(n11314), .ZN(n18943) );
  NOR2_X1 U14261 ( .A1(n11315), .A2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n11316) );
  NOR2_X1 U14262 ( .A1(n11313), .A2(n11316), .ZN(n18959) );
  XNOR2_X1 U14263 ( .A(n11317), .B(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n18984) );
  OAI21_X1 U14264 ( .B1(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n11318), .A(
        n11319), .ZN(n19009) );
  AOI21_X1 U14265 ( .B1(n15448), .B2(n9876), .A(n11320), .ZN(n19025) );
  AOI21_X1 U14266 ( .B1(n16266), .B2(n11321), .A(n11322), .ZN(n16259) );
  AOI21_X1 U14267 ( .B1(n16278), .B2(n11323), .A(n11324), .ZN(n16271) );
  AOI21_X1 U14268 ( .B1(n15459), .B2(n11325), .A(n11326), .ZN(n19047) );
  AOI21_X1 U14269 ( .B1(n16300), .B2(n11327), .A(n9877), .ZN(n19081) );
  AOI21_X1 U14270 ( .B1(n11328), .B2(n11329), .A(n11330), .ZN(n16301) );
  OAI22_X1 U14271 ( .A1(n13537), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(P2_STATE2_REG_0__SCAN_IN), .ZN(
        n15739) );
  INV_X1 U14272 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n13537) );
  INV_X1 U14273 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13691) );
  OAI22_X1 U14274 ( .A1(n13537), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(
        n13691), .B2(P2_STATE2_REG_0__SCAN_IN), .ZN(n14357) );
  AND2_X1 U14275 ( .A1(n15739), .A2(n14357), .ZN(n14234) );
  OAI21_X1 U14276 ( .B1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n11329), .ZN(n14236) );
  NAND2_X1 U14277 ( .A1(n14234), .A2(n14236), .ZN(n14050) );
  NOR2_X1 U14278 ( .A1(n16301), .A2(n14050), .ZN(n14147) );
  OAI21_X1 U14279 ( .B1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n11330), .A(
        n11327), .ZN(n19255) );
  NAND2_X1 U14280 ( .A1(n14147), .A2(n19255), .ZN(n19078) );
  NOR2_X1 U14281 ( .A1(n19081), .A2(n19078), .ZN(n19063) );
  OAI21_X1 U14282 ( .B1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n9877), .A(
        n11325), .ZN(n19065) );
  NAND2_X1 U14283 ( .A1(n19063), .A2(n19065), .ZN(n19046) );
  NOR2_X1 U14284 ( .A1(n19047), .A2(n19046), .ZN(n14180) );
  OAI21_X1 U14285 ( .B1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n11326), .A(
        n11323), .ZN(n16292) );
  NAND2_X1 U14286 ( .A1(n14180), .A2(n16292), .ZN(n14041) );
  NOR2_X1 U14287 ( .A1(n16271), .A2(n14041), .ZN(n19039) );
  OAI21_X1 U14288 ( .B1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n11324), .A(
        n11321), .ZN(n19040) );
  NAND2_X1 U14289 ( .A1(n19039), .A2(n19040), .ZN(n15141) );
  NOR2_X1 U14290 ( .A1(n16259), .A2(n15141), .ZN(n14262) );
  OAI21_X1 U14291 ( .B1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n11322), .A(
        n9876), .ZN(n16258) );
  NAND2_X1 U14292 ( .A1(n14262), .A2(n16258), .ZN(n19024) );
  NOR2_X1 U14293 ( .A1(n19025), .A2(n19024), .ZN(n19013) );
  INV_X1 U14294 ( .A(n11318), .ZN(n11331) );
  OAI21_X1 U14295 ( .B1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n11320), .A(
        n11331), .ZN(n19015) );
  AND2_X1 U14296 ( .A1(n19013), .A2(n19015), .ZN(n19010) );
  NAND2_X1 U14297 ( .A1(n19009), .A2(n19010), .ZN(n18990) );
  AOI21_X1 U14298 ( .B1(n11332), .B2(n11319), .A(n11317), .ZN(n18991) );
  NOR2_X1 U14299 ( .A1(n18990), .A2(n18991), .ZN(n18985) );
  AND2_X1 U14300 ( .A1(n18984), .A2(n18985), .ZN(n18966) );
  AOI21_X1 U14301 ( .B1(n11317), .B2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .A(
        P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n11333) );
  OR2_X1 U14302 ( .A1(n11315), .A2(n11333), .ZN(n18967) );
  NAND2_X1 U14303 ( .A1(n18966), .A2(n18967), .ZN(n11334) );
  NOR2_X1 U14304 ( .A1(n11335), .A2(n18941), .ZN(n13346) );
  NOR2_X1 U14305 ( .A1(n15378), .A2(n13346), .ZN(n13345) );
  NOR2_X1 U14306 ( .A1(n10053), .A2(n13357), .ZN(n15136) );
  NOR2_X1 U14307 ( .A1(n15137), .A2(n15136), .ZN(n15135) );
  NOR2_X1 U14308 ( .A1(n10053), .A2(n13329), .ZN(n15104) );
  NOR2_X1 U14309 ( .A1(n15105), .A2(n15104), .ZN(n15103) );
  NOR2_X1 U14310 ( .A1(n10053), .A2(n15103), .ZN(n15083) );
  NOR2_X1 U14311 ( .A1(n11336), .A2(n15083), .ZN(n15084) );
  XNOR2_X1 U14312 ( .A(n11296), .B(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12996) );
  NAND4_X1 U14313 ( .A1(n9868), .A2(n15084), .A3(n12996), .A4(n19079), .ZN(
        n11967) );
  AND2_X4 U14314 ( .A1(n11655), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12945) );
  AOI22_X1 U14315 ( .A1(n11427), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12945), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11338) );
  AOI22_X1 U14316 ( .A1(n12797), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n9857), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11337) );
  NAND2_X1 U14317 ( .A1(n11338), .A2(n11337), .ZN(n11343) );
  AND2_X4 U14318 ( .A1(n11653), .A2(n15752), .ZN(n12949) );
  AND2_X2 U14319 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11654) );
  AOI22_X1 U14320 ( .A1(n12949), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12828), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11341) );
  AND2_X2 U14321 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n12290) );
  AND2_X4 U14322 ( .A1(n12290), .A2(n15737), .ZN(n11646) );
  AND2_X4 U14323 ( .A1(n12290), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11645) );
  AOI22_X1 U14324 ( .A1(n11646), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11645), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11340) );
  NAND2_X1 U14325 ( .A1(n11341), .A2(n11340), .ZN(n11342) );
  INV_X2 U14326 ( .A(n11400), .ZN(n12798) );
  AOI22_X1 U14327 ( .A1(n9855), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12945), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11346) );
  AOI22_X1 U14328 ( .A1(n12797), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n9852), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11345) );
  AOI22_X1 U14329 ( .A1(n11646), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n11645), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11344) );
  NAND4_X1 U14330 ( .A1(n11347), .A2(n11346), .A3(n11345), .A4(n11344), .ZN(
        n11348) );
  AOI22_X1 U14331 ( .A1(n12949), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12945), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11353) );
  AOI22_X1 U14332 ( .A1(n12797), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12828), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11352) );
  NAND4_X1 U14333 ( .A1(n11354), .A2(n11353), .A3(n11352), .A4(n11351), .ZN(
        n11355) );
  NAND2_X1 U14334 ( .A1(n11355), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11362) );
  INV_X2 U14335 ( .A(n11400), .ZN(n12929) );
  AOI22_X1 U14336 ( .A1(n12949), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n12945), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11358) );
  AOI22_X1 U14337 ( .A1(n12797), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n9830), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11357) );
  AOI22_X1 U14338 ( .A1(n11646), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n11645), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11356) );
  NAND4_X1 U14339 ( .A1(n11359), .A2(n11358), .A3(n11357), .A4(n11356), .ZN(
        n11360) );
  NAND2_X1 U14340 ( .A1(n11360), .A2(n11651), .ZN(n11361) );
  AOI22_X1 U14341 ( .A1(n11427), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12798), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11366) );
  AOI22_X1 U14342 ( .A1(n12949), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12945), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11365) );
  AOI22_X1 U14343 ( .A1(n12797), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12828), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11364) );
  AOI22_X1 U14344 ( .A1(n11646), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11645), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11363) );
  NAND4_X1 U14345 ( .A1(n11366), .A2(n11365), .A3(n11364), .A4(n11363), .ZN(
        n11367) );
  AOI22_X1 U14346 ( .A1(n12797), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n9855), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11368) );
  NAND3_X1 U14347 ( .A1(n11370), .A2(n11369), .A3(n11368), .ZN(n11373) );
  AOI22_X1 U14348 ( .A1(n12945), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n12828), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11371) );
  NAND2_X1 U14349 ( .A1(n11375), .A2(n11374), .ZN(n11435) );
  AOI22_X1 U14350 ( .A1(n12798), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n12945), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11378) );
  AOI22_X1 U14351 ( .A1(n12949), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n9852), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11377) );
  AOI22_X1 U14352 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n11645), .B1(
        n11646), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11376) );
  NAND4_X1 U14353 ( .A1(n11379), .A2(n11378), .A3(n11377), .A4(n11376), .ZN(
        n11380) );
  NAND2_X1 U14354 ( .A1(n11380), .A2(n11651), .ZN(n11387) );
  AOI22_X1 U14355 ( .A1(n12949), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11427), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11384) );
  AOI22_X1 U14356 ( .A1(n12945), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n9830), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11383) );
  AOI22_X1 U14357 ( .A1(n12797), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12798), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11382) );
  AOI22_X1 U14358 ( .A1(n11646), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11645), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11381) );
  NAND4_X1 U14359 ( .A1(n11384), .A2(n11383), .A3(n11382), .A4(n11381), .ZN(
        n11385) );
  NAND2_X1 U14360 ( .A1(n11385), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11386) );
  AOI22_X1 U14361 ( .A1(n9857), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11427), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11391) );
  AOI22_X1 U14362 ( .A1(n12949), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12945), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11390) );
  AOI22_X1 U14363 ( .A1(n12797), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n9853), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11389) );
  AOI22_X1 U14364 ( .A1(n11646), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11645), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11388) );
  NAND4_X1 U14365 ( .A1(n11391), .A2(n11390), .A3(n11389), .A4(n11388), .ZN(
        n11392) );
  NAND2_X1 U14366 ( .A1(n11392), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11399) );
  AOI22_X1 U14367 ( .A1(n11427), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__6__SCAN_IN), .B2(n12929), .ZN(n11396) );
  AOI22_X1 U14368 ( .A1(n12949), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12945), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11395) );
  AOI22_X1 U14369 ( .A1(n12797), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n9830), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11394) );
  AOI22_X1 U14370 ( .A1(n11646), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11645), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11393) );
  NAND4_X1 U14371 ( .A1(n11396), .A2(n11395), .A3(n11394), .A4(n11393), .ZN(
        n11397) );
  NAND2_X1 U14372 ( .A1(n11397), .A2(n11651), .ZN(n11398) );
  AOI22_X1 U14373 ( .A1(n11427), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12929), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11405) );
  AOI22_X1 U14374 ( .A1(n9848), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12945), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11404) );
  NAND2_X1 U14375 ( .A1(n11645), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n11401) );
  AOI22_X1 U14376 ( .A1(n9847), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12945), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11408) );
  AOI22_X1 U14377 ( .A1(n9844), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(n9830), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11407) );
  AOI22_X1 U14378 ( .A1(n12949), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12945), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11413) );
  AOI22_X1 U14379 ( .A1(n12797), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n12929), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11412) );
  AOI22_X1 U14380 ( .A1(n11427), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n9853), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11411) );
  AOI22_X1 U14381 ( .A1(n11646), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n11645), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11410) );
  AOI22_X1 U14382 ( .A1(n12949), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12798), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11416) );
  AOI22_X1 U14383 ( .A1(n12945), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n9830), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11415) );
  AOI22_X1 U14384 ( .A1(n11646), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11645), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11414) );
  NAND2_X2 U14385 ( .A1(n11963), .A2(n16370), .ZN(n11638) );
  INV_X1 U14386 ( .A(n11451), .ZN(n11418) );
  INV_X1 U14387 ( .A(n11435), .ZN(n11419) );
  AND2_X1 U14388 ( .A1(n11436), .A2(n19290), .ZN(n12985) );
  NAND2_X2 U14389 ( .A1(n11461), .A2(n12392), .ZN(n13542) );
  AOI22_X1 U14390 ( .A1(n12797), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n11427), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11425) );
  AOI22_X1 U14391 ( .A1(n12949), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n12945), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11424) );
  AOI22_X1 U14392 ( .A1(n12798), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n9852), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11423) );
  AOI22_X1 U14393 ( .A1(n11646), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n11645), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11422) );
  AND4_X1 U14394 ( .A1(n11425), .A2(n11424), .A3(n11423), .A4(n11422), .ZN(
        n11426) );
  NAND2_X1 U14395 ( .A1(n11426), .A2(n11651), .ZN(n11434) );
  AOI22_X1 U14396 ( .A1(n12949), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12945), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11431) );
  AOI22_X1 U14397 ( .A1(n12797), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n9853), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11430) );
  AOI22_X1 U14398 ( .A1(n11646), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11645), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11429) );
  AOI22_X1 U14399 ( .A1(n12798), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n11427), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11428) );
  NAND2_X1 U14400 ( .A1(n11432), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11433) );
  AND2_X1 U14401 ( .A1(n11443), .A2(n12380), .ZN(n12426) );
  OAI21_X1 U14402 ( .B1(n12114), .B2(n11438), .A(n11419), .ZN(n11440) );
  NAND2_X1 U14403 ( .A1(n14035), .A2(n11794), .ZN(n11439) );
  NAND2_X1 U14404 ( .A1(n12392), .A2(n11443), .ZN(n12305) );
  INV_X1 U14405 ( .A(n11508), .ZN(n11448) );
  INV_X1 U14406 ( .A(P2_EBX_REG_1__SCAN_IN), .ZN(n13585) );
  NAND2_X1 U14407 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n11446) );
  INV_X1 U14408 ( .A(n11638), .ZN(n11444) );
  AND2_X4 U14409 ( .A1(n13559), .A2(n13427), .ZN(n12897) );
  AND2_X4 U14410 ( .A1(n11444), .A2(n12897), .ZN(n11610) );
  NAND2_X1 U14411 ( .A1(n11610), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n11445) );
  OAI211_X1 U14412 ( .C1(n11543), .C2(n13585), .A(n11446), .B(n11445), .ZN(
        n11447) );
  AOI21_X2 U14413 ( .B1(n11448), .B2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n11447), .ZN(n11483) );
  NAND2_X1 U14414 ( .A1(n11794), .A2(n19271), .ZN(n12430) );
  OR2_X1 U14415 ( .A1(n12439), .A2(n12430), .ZN(n11449) );
  NAND2_X1 U14416 ( .A1(n11450), .A2(n11449), .ZN(n11466) );
  INV_X1 U14417 ( .A(n11963), .ZN(n11455) );
  NOR2_X2 U14418 ( .A1(n11452), .A2(n11788), .ZN(n11457) );
  NAND2_X1 U14419 ( .A1(n11453), .A2(n11457), .ZN(n12387) );
  NAND3_X1 U14420 ( .A1(n12387), .A2(n12380), .A3(n13427), .ZN(n11454) );
  NAND2_X1 U14421 ( .A1(n11455), .A2(n11454), .ZN(n12422) );
  AOI21_X1 U14422 ( .B1(n11794), .B2(n14035), .A(n19275), .ZN(n11460) );
  INV_X1 U14423 ( .A(n11461), .ZN(n11462) );
  NAND2_X1 U14424 ( .A1(n11463), .A2(n9911), .ZN(n12437) );
  OAI21_X1 U14425 ( .B1(n12422), .B2(n12392), .A(n12437), .ZN(n11464) );
  INV_X1 U14426 ( .A(n11464), .ZN(n11465) );
  AOI22_X1 U14427 ( .A1(n15774), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(n13431), 
        .B2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n11467) );
  OAI21_X2 U14428 ( .B1(n11494), .B2(n10246), .A(n11467), .ZN(n11482) );
  NAND2_X1 U14429 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_STATE2_REG_0__SCAN_IN), .ZN(n11468) );
  NAND2_X1 U14430 ( .A1(n11543), .A2(n11468), .ZN(n11469) );
  OAI21_X1 U14431 ( .B1(n11471), .B2(n11470), .A(n11469), .ZN(n11476) );
  INV_X1 U14432 ( .A(n13431), .ZN(n11473) );
  OAI22_X1 U14433 ( .A1(n11472), .A2(n13537), .B1(n11473), .B2(n19924), .ZN(
        n11474) );
  INV_X1 U14434 ( .A(n11474), .ZN(n11475) );
  NAND2_X1 U14435 ( .A1(n11476), .A2(n11475), .ZN(n11980) );
  INV_X1 U14436 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n11481) );
  INV_X1 U14437 ( .A(P2_EBX_REG_0__SCAN_IN), .ZN(n12115) );
  AND2_X1 U14438 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n11477) );
  NOR2_X1 U14439 ( .A1(n13431), .A2(n11477), .ZN(n11478) );
  INV_X1 U14440 ( .A(n11482), .ZN(n11484) );
  AOI21_X1 U14441 ( .B1(n13537), .B2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n11485) );
  INV_X1 U14442 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n13629) );
  NAND2_X1 U14443 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n11488) );
  NAND2_X1 U14444 ( .A1(n11610), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n11487) );
  OAI211_X1 U14445 ( .C1(n11543), .C2(n13629), .A(n11488), .B(n11487), .ZN(
        n11489) );
  INV_X1 U14446 ( .A(n11489), .ZN(n11490) );
  NAND2_X1 U14447 ( .A1(n11493), .A2(n11492), .ZN(n11502) );
  INV_X1 U14448 ( .A(n11494), .ZN(n11495) );
  NAND2_X1 U14449 ( .A1(n11495), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11497) );
  NAND2_X1 U14450 ( .A1(n13431), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n11496) );
  NAND2_X1 U14451 ( .A1(n11497), .A2(n11496), .ZN(n11503) );
  INV_X1 U14452 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n14095) );
  INV_X1 U14453 ( .A(P2_EBX_REG_3__SCAN_IN), .ZN(n14054) );
  NAND2_X1 U14454 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n11499) );
  NAND2_X1 U14455 ( .A1(n11610), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n11498) );
  OAI211_X1 U14456 ( .C1(n11543), .C2(n14054), .A(n11499), .B(n11498), .ZN(
        n11500) );
  XNOR2_X2 U14457 ( .A(n11503), .B(n11504), .ZN(n11971) );
  NAND2_X1 U14458 ( .A1(n11502), .A2(n11971), .ZN(n11507) );
  INV_X1 U14459 ( .A(n11503), .ZN(n11505) );
  NAND2_X1 U14460 ( .A1(n11505), .A2(n11504), .ZN(n11506) );
  NAND2_X1 U14461 ( .A1(n11507), .A2(n11506), .ZN(n13829) );
  INV_X1 U14462 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n21161) );
  OR2_X1 U14463 ( .A1(n11613), .A2(n21161), .ZN(n11513) );
  INV_X1 U14464 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n13831) );
  NAND2_X1 U14465 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n11510) );
  NAND2_X1 U14466 ( .A1(n11610), .A2(P2_REIP_REG_4__SCAN_IN), .ZN(n11509) );
  OAI211_X1 U14467 ( .C1(n11606), .C2(n13831), .A(n11510), .B(n11509), .ZN(
        n11511) );
  INV_X1 U14468 ( .A(n11511), .ZN(n11512) );
  INV_X1 U14469 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n14226) );
  OR2_X1 U14470 ( .A1(n11613), .A2(n14226), .ZN(n11520) );
  INV_X1 U14471 ( .A(P2_EBX_REG_5__SCAN_IN), .ZN(n19073) );
  NAND2_X1 U14472 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n11517) );
  NAND2_X1 U14473 ( .A1(n11610), .A2(P2_REIP_REG_5__SCAN_IN), .ZN(n11516) );
  OAI211_X1 U14474 ( .C1(n11606), .C2(n19073), .A(n11517), .B(n11516), .ZN(
        n11518) );
  INV_X1 U14475 ( .A(n11518), .ZN(n11519) );
  INV_X1 U14476 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n12425) );
  OR2_X1 U14477 ( .A1(n11613), .A2(n12425), .ZN(n11527) );
  INV_X1 U14478 ( .A(P2_EBX_REG_6__SCAN_IN), .ZN(n11524) );
  NAND2_X1 U14479 ( .A1(n11610), .A2(P2_REIP_REG_6__SCAN_IN), .ZN(n11523) );
  NAND2_X1 U14480 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n11522) );
  OAI211_X1 U14481 ( .C1(n11606), .C2(n11524), .A(n11523), .B(n11522), .ZN(
        n11525) );
  INV_X1 U14482 ( .A(n11525), .ZN(n11526) );
  INV_X1 U14483 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n11530) );
  INV_X1 U14484 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n15730) );
  OR2_X1 U14485 ( .A1(n11613), .A2(n15730), .ZN(n11529) );
  AOI22_X1 U14486 ( .A1(n11609), .A2(P2_EBX_REG_7__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11528) );
  OAI211_X1 U14487 ( .C1(n11602), .C2(n11530), .A(n11529), .B(n11528), .ZN(
        n13857) );
  INV_X1 U14488 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n12364) );
  OR2_X1 U14489 ( .A1(n11613), .A2(n12364), .ZN(n11535) );
  NAND2_X1 U14490 ( .A1(n11610), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n11532) );
  NAND2_X1 U14491 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n11531) );
  OAI211_X1 U14492 ( .C1(n11606), .C2(n10078), .A(n11532), .B(n11531), .ZN(
        n11533) );
  INV_X1 U14493 ( .A(n11533), .ZN(n11534) );
  NAND2_X1 U14494 ( .A1(n11535), .A2(n11534), .ZN(n13878) );
  INV_X1 U14495 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15712) );
  OR2_X1 U14496 ( .A1(n11613), .A2(n15712), .ZN(n11540) );
  INV_X1 U14497 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n12184) );
  NAND2_X1 U14498 ( .A1(n11610), .A2(P2_REIP_REG_9__SCAN_IN), .ZN(n11537) );
  NAND2_X1 U14499 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n11536) );
  OAI211_X1 U14500 ( .C1(n11606), .C2(n12184), .A(n11537), .B(n11536), .ZN(
        n11538) );
  INV_X1 U14501 ( .A(n11538), .ZN(n11539) );
  INV_X1 U14502 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n12180) );
  OR2_X1 U14503 ( .A1(n11613), .A2(n12180), .ZN(n11546) );
  INV_X1 U14504 ( .A(P2_EBX_REG_10__SCAN_IN), .ZN(n19034) );
  NAND2_X1 U14505 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n11542) );
  NAND2_X1 U14506 ( .A1(n11610), .A2(P2_REIP_REG_10__SCAN_IN), .ZN(n11541) );
  OAI211_X1 U14507 ( .C1(n11543), .C2(n19034), .A(n11542), .B(n11541), .ZN(
        n11544) );
  INV_X1 U14508 ( .A(n11544), .ZN(n11545) );
  NAND2_X1 U14509 ( .A1(n11546), .A2(n11545), .ZN(n13927) );
  INV_X1 U14510 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n11878) );
  INV_X1 U14511 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15676) );
  OR2_X1 U14512 ( .A1(n11613), .A2(n15676), .ZN(n11548) );
  AOI22_X1 U14513 ( .A1(n11609), .A2(P2_EBX_REG_11__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), 
        .ZN(n11547) );
  OAI211_X1 U14514 ( .C1(n11602), .C2(n11878), .A(n11548), .B(n11547), .ZN(
        n13953) );
  INV_X1 U14515 ( .A(P2_EBX_REG_12__SCAN_IN), .ZN(n14270) );
  NAND2_X1 U14516 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n11550) );
  NAND2_X1 U14517 ( .A1(n11610), .A2(P2_REIP_REG_12__SCAN_IN), .ZN(n11549) );
  OAI211_X1 U14518 ( .C1(n11606), .C2(n14270), .A(n11550), .B(n11549), .ZN(
        n11551) );
  AOI21_X1 U14519 ( .B1(n11608), .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n11551), .ZN(n14015) );
  INV_X1 U14520 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n15449) );
  INV_X1 U14521 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n21086) );
  OR2_X1 U14522 ( .A1(n11613), .A2(n21086), .ZN(n11553) );
  AOI22_X1 U14523 ( .A1(n11609), .A2(P2_EBX_REG_13__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), 
        .ZN(n11552) );
  OAI211_X1 U14524 ( .C1(n11602), .C2(n15449), .A(n11553), .B(n11552), .ZN(
        n14066) );
  NAND2_X1 U14525 ( .A1(n14017), .A2(n14066), .ZN(n14065) );
  INV_X1 U14526 ( .A(n14065), .ZN(n11558) );
  INV_X1 U14527 ( .A(P2_EBX_REG_14__SCAN_IN), .ZN(n14146) );
  NAND2_X1 U14528 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n11555) );
  NAND2_X1 U14529 ( .A1(n11610), .A2(P2_REIP_REG_14__SCAN_IN), .ZN(n11554) );
  OAI211_X1 U14530 ( .C1(n11606), .C2(n14146), .A(n11555), .B(n11554), .ZN(
        n11556) );
  AOI21_X1 U14531 ( .B1(n11608), .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n11556), .ZN(n14142) );
  INV_X1 U14532 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n12216) );
  NAND2_X1 U14533 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n11560) );
  NAND2_X1 U14534 ( .A1(n11610), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n11559) );
  OAI211_X1 U14535 ( .C1(n11606), .C2(n12216), .A(n11560), .B(n11559), .ZN(
        n11561) );
  AOI21_X1 U14536 ( .B1(n11608), .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n11561), .ZN(n14210) );
  INV_X1 U14537 ( .A(P2_EBX_REG_16__SCAN_IN), .ZN(n18992) );
  NAND2_X1 U14538 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n11563) );
  NAND2_X1 U14539 ( .A1(n11610), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n11562) );
  OAI211_X1 U14540 ( .C1(n11606), .C2(n18992), .A(n11563), .B(n11562), .ZN(
        n11564) );
  AOI21_X1 U14541 ( .B1(n11608), .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n11564), .ZN(n14352) );
  INV_X1 U14542 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n21095) );
  INV_X1 U14543 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15622) );
  OR2_X1 U14544 ( .A1(n11613), .A2(n15622), .ZN(n11566) );
  AOI22_X1 U14545 ( .A1(n11609), .A2(P2_EBX_REG_17__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), 
        .ZN(n11565) );
  OAI211_X1 U14546 ( .C1(n21095), .C2(n11602), .A(n11566), .B(n11565), .ZN(
        n14323) );
  INV_X1 U14547 ( .A(P2_EBX_REG_18__SCAN_IN), .ZN(n18968) );
  NAND2_X1 U14548 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n11568) );
  NAND2_X1 U14549 ( .A1(n11610), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n11567) );
  OAI211_X1 U14550 ( .C1(n11606), .C2(n18968), .A(n11568), .B(n11567), .ZN(
        n11569) );
  AOI21_X1 U14551 ( .B1(n11608), .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n11569), .ZN(n14381) );
  INV_X1 U14552 ( .A(P2_EBX_REG_19__SCAN_IN), .ZN(n12228) );
  NAND2_X1 U14553 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n11571) );
  INV_X1 U14554 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n19854) );
  OR2_X1 U14555 ( .A1(n11602), .A2(n19854), .ZN(n11570) );
  OAI211_X1 U14556 ( .C1(n11606), .C2(n12228), .A(n11571), .B(n11570), .ZN(
        n11572) );
  AOI21_X1 U14557 ( .B1(n11608), .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n11572), .ZN(n15226) );
  INV_X1 U14558 ( .A(n15226), .ZN(n11573) );
  INV_X1 U14559 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n19856) );
  INV_X1 U14560 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15388) );
  OR2_X1 U14561 ( .A1(n11613), .A2(n15388), .ZN(n11575) );
  AOI22_X1 U14562 ( .A1(n11609), .A2(P2_EBX_REG_20__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), 
        .ZN(n11574) );
  OAI211_X1 U14563 ( .C1(n11602), .C2(n19856), .A(n11575), .B(n11574), .ZN(
        n15217) );
  INV_X1 U14564 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n21126) );
  INV_X1 U14565 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n15376) );
  OR2_X1 U14566 ( .A1(n11613), .A2(n15376), .ZN(n11577) );
  AOI22_X1 U14567 ( .A1(n11609), .A2(P2_EBX_REG_21__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), 
        .ZN(n11576) );
  OAI211_X1 U14568 ( .C1(n11602), .C2(n21126), .A(n11577), .B(n11576), .ZN(
        n13349) );
  INV_X1 U14569 ( .A(P2_EBX_REG_22__SCAN_IN), .ZN(n11580) );
  NAND2_X1 U14570 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n11579) );
  INV_X1 U14571 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n15861) );
  OR2_X1 U14572 ( .A1(n11602), .A2(n15861), .ZN(n11578) );
  OAI211_X1 U14573 ( .C1(n11606), .C2(n11580), .A(n11579), .B(n11578), .ZN(
        n11581) );
  AOI21_X1 U14574 ( .B1(n11608), .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n11581), .ZN(n15200) );
  INV_X1 U14575 ( .A(P2_EBX_REG_23__SCAN_IN), .ZN(n11753) );
  NAND2_X1 U14576 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n11583) );
  INV_X1 U14577 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n19860) );
  OR2_X1 U14578 ( .A1(n11602), .A2(n19860), .ZN(n11582) );
  OAI211_X1 U14579 ( .C1(n11606), .C2(n11753), .A(n11583), .B(n11582), .ZN(
        n11584) );
  AOI21_X1 U14580 ( .B1(n11608), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n11584), .ZN(n13360) );
  NAND2_X1 U14581 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n11586) );
  NAND2_X1 U14582 ( .A1(n11610), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n11585) );
  OAI211_X1 U14583 ( .C1(n11606), .C2(n10047), .A(n11586), .B(n11585), .ZN(
        n11587) );
  AOI21_X1 U14584 ( .B1(n11608), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n11587), .ZN(n15126) );
  INV_X1 U14585 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n19864) );
  INV_X1 U14586 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15509) );
  OR2_X1 U14587 ( .A1(n11613), .A2(n15509), .ZN(n11589) );
  AOI22_X1 U14588 ( .A1(n11609), .A2(P2_EBX_REG_25__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), 
        .ZN(n11588) );
  OAI211_X1 U14589 ( .C1(n11602), .C2(n19864), .A(n11589), .B(n11588), .ZN(
        n15113) );
  INV_X1 U14590 ( .A(P2_EBX_REG_26__SCAN_IN), .ZN(n12262) );
  NAND2_X1 U14591 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n11591) );
  INV_X1 U14592 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n19866) );
  OR2_X1 U14593 ( .A1(n11602), .A2(n19866), .ZN(n11590) );
  OAI211_X1 U14594 ( .C1(n11606), .C2(n12262), .A(n11591), .B(n11590), .ZN(
        n11592) );
  AOI21_X1 U14595 ( .B1(n11608), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n11592), .ZN(n15176) );
  INV_X1 U14596 ( .A(P2_EBX_REG_27__SCAN_IN), .ZN(n13331) );
  NAND2_X1 U14597 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n11595) );
  INV_X1 U14598 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n21193) );
  OR2_X1 U14599 ( .A1(n11602), .A2(n21193), .ZN(n11594) );
  OAI211_X1 U14600 ( .C1(n11606), .C2(n13331), .A(n11595), .B(n11594), .ZN(
        n11596) );
  AOI21_X1 U14601 ( .B1(n11608), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n11596), .ZN(n13333) );
  INV_X1 U14602 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n19869) );
  INV_X1 U14603 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15473) );
  OR2_X1 U14604 ( .A1(n11613), .A2(n15473), .ZN(n11598) );
  AOI22_X1 U14605 ( .A1(n11609), .A2(P2_EBX_REG_28__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), 
        .ZN(n11597) );
  OAI211_X1 U14606 ( .C1(n11602), .C2(n19869), .A(n11598), .B(n11597), .ZN(
        n12297) );
  INV_X1 U14607 ( .A(P2_EBX_REG_29__SCAN_IN), .ZN(n15089) );
  NAND2_X1 U14608 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n11600) );
  INV_X1 U14609 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n19871) );
  OR2_X1 U14610 ( .A1(n11602), .A2(n19871), .ZN(n11599) );
  OAI211_X1 U14611 ( .C1(n11606), .C2(n15089), .A(n11600), .B(n11599), .ZN(
        n11601) );
  AOI21_X1 U14612 ( .B1(n11608), .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n11601), .ZN(n12486) );
  INV_X1 U14613 ( .A(P2_EBX_REG_30__SCAN_IN), .ZN(n11605) );
  NAND2_X1 U14614 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n11604) );
  INV_X1 U14615 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n12509) );
  OR2_X1 U14616 ( .A1(n11602), .A2(n12509), .ZN(n11603) );
  OAI211_X1 U14617 ( .C1(n11606), .C2(n11605), .A(n11604), .B(n11603), .ZN(
        n11607) );
  AOI21_X1 U14618 ( .B1(n11608), .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n11607), .ZN(n12507) );
  AOI22_X1 U14619 ( .A1(n11609), .A2(P2_EBX_REG_31__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n11612) );
  NAND2_X1 U14620 ( .A1(n11610), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n11611) );
  OAI211_X1 U14621 ( .C1(n11613), .C2(n20998), .A(n11612), .B(n11611), .ZN(
        n11614) );
  XNOR2_X1 U14622 ( .A(n11615), .B(n11614), .ZN(n12454) );
  XNOR2_X1 U14623 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n12298) );
  NAND2_X1 U14624 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n19924), .ZN(
        n12113) );
  INV_X1 U14625 ( .A(n12113), .ZN(n11617) );
  NAND2_X1 U14626 ( .A1(n12298), .A2(n11617), .ZN(n11619) );
  NAND2_X1 U14627 ( .A1(n19914), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11618) );
  NAND2_X1 U14628 ( .A1(n11619), .A2(n11618), .ZN(n11629) );
  XNOR2_X1 U14629 ( .A(n15752), .B(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n11627) );
  NAND2_X1 U14630 ( .A1(n11629), .A2(n11627), .ZN(n11621) );
  NAND2_X1 U14631 ( .A1(n19905), .A2(n15752), .ZN(n11620) );
  NAND2_X1 U14632 ( .A1(n11621), .A2(n11620), .ZN(n11631) );
  XNOR2_X1 U14633 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n11630) );
  NAND2_X1 U14634 ( .A1(n11631), .A2(n11630), .ZN(n11623) );
  NAND2_X1 U14635 ( .A1(n19898), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11622) );
  NAND2_X1 U14636 ( .A1(n11623), .A2(n11622), .ZN(n11632) );
  AND2_X1 U14637 ( .A1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n15918), .ZN(
        n11624) );
  INV_X1 U14638 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n13545) );
  NAND2_X1 U14639 ( .A1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n13545), .ZN(
        n11625) );
  XNOR2_X1 U14640 ( .A(n12298), .B(n12113), .ZN(n12301) );
  INV_X1 U14641 ( .A(n11627), .ZN(n11628) );
  XNOR2_X1 U14642 ( .A(n11629), .B(n11628), .ZN(n12307) );
  XNOR2_X1 U14643 ( .A(n11631), .B(n11630), .ZN(n11687) );
  INV_X1 U14644 ( .A(n11687), .ZN(n11633) );
  NAND2_X1 U14645 ( .A1(n12307), .A2(n12313), .ZN(n12289) );
  INV_X1 U14646 ( .A(n12289), .ZN(n11634) );
  NAND2_X1 U14647 ( .A1(n12301), .A2(n11634), .ZN(n11635) );
  NAND2_X1 U14648 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19802), .ZN(n11641) );
  INV_X1 U14649 ( .A(n11641), .ZN(n11636) );
  NAND2_X1 U14650 ( .A1(n11616), .A2(n11964), .ZN(n13433) );
  OR2_X1 U14651 ( .A1(n13433), .A2(n12308), .ZN(n11758) );
  INV_X1 U14652 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n19573) );
  NAND2_X1 U14653 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n19803) );
  NAND2_X1 U14654 ( .A1(n19573), .A2(n19803), .ZN(n11756) );
  INV_X1 U14655 ( .A(n11964), .ZN(n13419) );
  NOR2_X1 U14656 ( .A1(n11638), .A2(n13419), .ZN(n13437) );
  INV_X1 U14657 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n15158) );
  NAND2_X1 U14658 ( .A1(n11756), .A2(n15158), .ZN(n11639) );
  NAND2_X2 U14659 ( .A1(n19940), .A2(P2_STATE_REG_2__SCAN_IN), .ZN(n19873) );
  NOR2_X1 U14660 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(P2_STATE_REG_2__SCAN_IN), 
        .ZN(n18913) );
  INV_X1 U14661 ( .A(n18913), .ZN(n19824) );
  NAND2_X1 U14662 ( .A1(n19818), .A2(n19803), .ZN(n16372) );
  INV_X1 U14663 ( .A(n16372), .ZN(n13530) );
  AOI22_X1 U14664 ( .A1(n13427), .A2(n11639), .B1(n19573), .B2(n13530), .ZN(
        n11640) );
  NOR2_X2 U14665 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19691) );
  NAND2_X1 U14666 ( .A1(n13431), .A2(n19691), .ZN(n12458) );
  INV_X1 U14667 ( .A(n19038), .ZN(n15684) );
  NOR3_X1 U14668 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n11641), .A3(n19917), 
        .ZN(n16395) );
  NOR2_X1 U14669 ( .A1(n9868), .A2(n16395), .ZN(n11642) );
  AND2_X1 U14670 ( .A1(n15684), .A2(n11642), .ZN(n11643) );
  AOI22_X1 U14671 ( .A1(P2_EBX_REG_31__SCAN_IN), .A2(n19090), .B1(
        P2_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n19101), .ZN(n11644) );
  AND2_X1 U14672 ( .A1(n12944), .A2(n11651), .ZN(n11766) );
  AOI22_X1 U14673 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n11723), .B1(
        n12781), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11650) );
  AOI22_X1 U14674 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n12782), .B1(
        n11727), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11649) );
  AND2_X2 U14675 ( .A1(n11427), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11772) );
  AOI22_X1 U14676 ( .A1(n11772), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11771), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11648) );
  INV_X1 U14677 ( .A(n11645), .ZN(n12801) );
  AND2_X2 U14678 ( .A1(n12953), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11770) );
  AOI22_X1 U14679 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n11777), .B1(
        n11770), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11647) );
  NAND4_X1 U14680 ( .A1(n11650), .A2(n11649), .A3(n11648), .A4(n11647), .ZN(
        n11661) );
  AND2_X2 U14681 ( .A1(n12945), .A2(n11651), .ZN(n11778) );
  AOI22_X1 U14682 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n11778), .B1(
        n11680), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11659) );
  INV_X2 U14683 ( .A(n10264), .ZN(n12788) );
  AOI22_X1 U14684 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n12783), .B1(
        n12788), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11658) );
  AOI22_X1 U14686 ( .A1(n11776), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n12789), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11657) );
  AOI22_X1 U14687 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n11667), .B1(
        n11668), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11656) );
  NAND4_X1 U14688 ( .A1(n11659), .A2(n11658), .A3(n11657), .A4(n11656), .ZN(
        n11660) );
  NOR2_X1 U14689 ( .A1(n11661), .A2(n11660), .ZN(n12328) );
  INV_X1 U14690 ( .A(n12307), .ZN(n12306) );
  NAND2_X1 U14691 ( .A1(n12285), .A2(n11451), .ZN(n11662) );
  AOI22_X1 U14692 ( .A1(n12781), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n11777), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11666) );
  AOI22_X1 U14693 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n12783), .B1(
        n12788), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11665) );
  AOI22_X1 U14694 ( .A1(n11723), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n11770), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11664) );
  AOI22_X1 U14695 ( .A1(n11778), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n11771), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11663) );
  NAND4_X1 U14696 ( .A1(n11666), .A2(n11665), .A3(n11664), .A4(n11663), .ZN(
        n11674) );
  AOI22_X1 U14697 ( .A1(n11667), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n11668), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11672) );
  AOI22_X1 U14698 ( .A1(n11776), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n12789), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11671) );
  AOI22_X1 U14699 ( .A1(n12782), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11680), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11670) );
  AOI22_X1 U14700 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n11727), .B1(
        n11772), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11669) );
  NAND4_X1 U14701 ( .A1(n11672), .A2(n11671), .A3(n11670), .A4(n11669), .ZN(
        n11673) );
  NAND2_X1 U14702 ( .A1(n13585), .A2(n12115), .ZN(n11675) );
  MUX2_X1 U14703 ( .A(n12330), .B(n11675), .S(n12412), .Z(n12118) );
  AOI22_X1 U14704 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n11723), .B1(
        n12781), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11679) );
  AOI22_X1 U14705 ( .A1(n11727), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12783), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11678) );
  AOI22_X1 U14706 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n11668), .B1(
        n12789), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11677) );
  AOI22_X1 U14707 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n11667), .B1(
        n11776), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11676) );
  NAND4_X1 U14708 ( .A1(n11679), .A2(n11678), .A3(n11677), .A4(n11676), .ZN(
        n11686) );
  AOI22_X1 U14709 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n11778), .B1(
        n11680), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11684) );
  AOI22_X1 U14710 ( .A1(n12782), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11771), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11683) );
  AOI22_X1 U14711 ( .A1(n11772), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11770), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11682) );
  AOI22_X1 U14712 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n11777), .B1(
        n12788), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11681) );
  NAND4_X1 U14713 ( .A1(n11684), .A2(n11683), .A3(n11682), .A4(n11681), .ZN(
        n11685) );
  NAND2_X1 U14714 ( .A1(n12308), .A2(n11687), .ZN(n11688) );
  OAI21_X1 U14715 ( .B1(n12308), .B2(n12059), .A(n11688), .ZN(n11689) );
  INV_X1 U14716 ( .A(n11689), .ZN(n11690) );
  MUX2_X1 U14717 ( .A(n11690), .B(n14054), .S(n11788), .Z(n12108) );
  AOI22_X1 U14718 ( .A1(n11723), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11772), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11694) );
  AOI22_X1 U14719 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n12781), .B1(
        n11727), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11693) );
  AOI22_X1 U14720 ( .A1(n12782), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n11771), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11692) );
  AOI22_X1 U14721 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n12783), .B1(
        n11770), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11691) );
  NAND4_X1 U14722 ( .A1(n11694), .A2(n11693), .A3(n11692), .A4(n11691), .ZN(
        n11700) );
  AOI22_X1 U14723 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n11778), .B1(
        n11680), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11698) );
  AOI22_X1 U14724 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n11777), .B1(
        n12788), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11697) );
  AOI22_X1 U14725 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n11668), .B1(
        n12789), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11696) );
  AOI22_X1 U14726 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n11667), .B1(
        n11776), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11695) );
  NAND4_X1 U14727 ( .A1(n11698), .A2(n11697), .A3(n11696), .A4(n11695), .ZN(
        n11699) );
  MUX2_X1 U14728 ( .A(n11813), .B(n11701), .S(n12308), .Z(n11702) );
  MUX2_X1 U14729 ( .A(n13831), .B(n11702), .S(n19286), .Z(n12125) );
  AOI22_X1 U14730 ( .A1(n12781), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11772), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11706) );
  AOI22_X1 U14731 ( .A1(n11723), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11727), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11705) );
  AOI22_X1 U14732 ( .A1(n12782), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11771), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11704) );
  AOI22_X1 U14733 ( .A1(n11770), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12783), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11703) );
  NAND4_X1 U14734 ( .A1(n11706), .A2(n11705), .A3(n11704), .A4(n11703), .ZN(
        n11712) );
  AOI22_X1 U14735 ( .A1(n11778), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11680), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11710) );
  AOI22_X1 U14736 ( .A1(n12788), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11777), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11709) );
  AOI22_X1 U14737 ( .A1(n11776), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n12789), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11708) );
  AOI22_X1 U14738 ( .A1(n11667), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n11668), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11707) );
  NAND4_X1 U14739 ( .A1(n11710), .A2(n11709), .A3(n11708), .A4(n11707), .ZN(
        n11711) );
  MUX2_X1 U14740 ( .A(n19073), .B(n12096), .S(n19286), .Z(n12103) );
  AOI22_X1 U14741 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n12781), .B1(
        n11772), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11716) );
  AOI22_X1 U14742 ( .A1(n11723), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11727), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11715) );
  AOI22_X1 U14743 ( .A1(n12782), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11771), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11714) );
  AOI22_X1 U14744 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n11777), .B1(
        n11770), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11713) );
  NAND4_X1 U14745 ( .A1(n11716), .A2(n11715), .A3(n11714), .A4(n11713), .ZN(
        n11722) );
  AOI22_X1 U14746 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n11778), .B1(
        n11680), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11720) );
  AOI22_X1 U14747 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n12783), .B1(
        n12788), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11719) );
  AOI22_X1 U14748 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n11776), .B1(
        n12789), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11718) );
  AOI22_X1 U14749 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n11667), .B1(
        n11668), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11717) );
  NAND4_X1 U14750 ( .A1(n11720), .A2(n11719), .A3(n11718), .A4(n11717), .ZN(
        n11721) );
  MUX2_X1 U14751 ( .A(n12162), .B(P2_EBX_REG_6__SCAN_IN), .S(n12412), .Z(
        n12166) );
  INV_X1 U14752 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n13858) );
  INV_X1 U14753 ( .A(n11723), .ZN(n11726) );
  INV_X1 U14754 ( .A(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12948) );
  INV_X1 U14755 ( .A(n11772), .ZN(n11725) );
  INV_X1 U14756 ( .A(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11724) );
  OAI22_X1 U14757 ( .A1(n11726), .A2(n12948), .B1(n11725), .B2(n11724), .ZN(
        n11733) );
  INV_X1 U14758 ( .A(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11731) );
  INV_X1 U14759 ( .A(n11727), .ZN(n11730) );
  INV_X1 U14760 ( .A(n11771), .ZN(n11729) );
  INV_X1 U14761 ( .A(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11728) );
  OAI22_X1 U14762 ( .A1(n11731), .A2(n11730), .B1(n11729), .B2(n11728), .ZN(
        n11732) );
  NOR2_X1 U14763 ( .A1(n11733), .A2(n11732), .ZN(n11745) );
  NAND2_X1 U14764 ( .A1(n12782), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n11737) );
  NAND2_X1 U14765 ( .A1(n12781), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n11736) );
  NAND2_X1 U14766 ( .A1(n11777), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n11735) );
  NAND2_X1 U14767 ( .A1(n11770), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n11734) );
  AOI22_X1 U14768 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n11776), .B1(
        n12789), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11741) );
  AOI22_X1 U14769 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n11667), .B1(
        n11668), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11740) );
  NAND2_X1 U14770 ( .A1(n11778), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n11739) );
  NAND2_X1 U14771 ( .A1(n11680), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n11738) );
  AOI22_X1 U14772 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n12783), .B1(
        n12788), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11742) );
  MUX2_X1 U14773 ( .A(n13858), .B(n12102), .S(n19286), .Z(n12172) );
  NAND2_X1 U14774 ( .A1(n12173), .A2(n12172), .ZN(n12175) );
  INV_X1 U14775 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n15144) );
  NAND2_X1 U14776 ( .A1(n12412), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n11746) );
  NAND2_X1 U14777 ( .A1(n12412), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n12211) );
  AND2_X2 U14778 ( .A1(n12213), .A2(n12211), .ZN(n12200) );
  NAND2_X1 U14779 ( .A1(n14146), .A2(n12216), .ZN(n11747) );
  NAND2_X1 U14780 ( .A1(n12412), .A2(n11747), .ZN(n11748) );
  NOR2_X1 U14781 ( .A1(n19286), .A2(n18992), .ZN(n11749) );
  NOR2_X2 U14782 ( .A1(n12219), .A2(n11749), .ZN(n12206) );
  NAND2_X1 U14783 ( .A1(n12412), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n12207) );
  NOR2_X1 U14784 ( .A1(P2_EBX_REG_18__SCAN_IN), .A2(P2_EBX_REG_19__SCAN_IN), 
        .ZN(n11750) );
  NOR2_X1 U14785 ( .A1(n19286), .A2(n11750), .ZN(n11751) );
  INV_X1 U14786 ( .A(P2_EBX_REG_21__SCAN_IN), .ZN(n15213) );
  NAND2_X1 U14787 ( .A1(n12412), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n12248) );
  NOR2_X1 U14788 ( .A1(n19286), .A2(n11753), .ZN(n12252) );
  NAND2_X1 U14789 ( .A1(n12273), .A2(n12269), .ZN(n12264) );
  NAND2_X1 U14790 ( .A1(n12412), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n12272) );
  INV_X1 U14791 ( .A(P2_EBX_REG_28__SCAN_IN), .ZN(n11754) );
  NOR2_X1 U14792 ( .A1(n19286), .A2(n11754), .ZN(n12279) );
  NAND2_X1 U14793 ( .A1(n12412), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n12410) );
  NAND2_X1 U14794 ( .A1(n12411), .A2(n12410), .ZN(n12414) );
  OAI21_X1 U14795 ( .B1(n12414), .B2(P2_EBX_REG_30__SCAN_IN), .A(n12412), .ZN(
        n11755) );
  NAND2_X1 U14796 ( .A1(n11755), .A2(n12269), .ZN(n12418) );
  INV_X1 U14797 ( .A(n12418), .ZN(n11759) );
  NAND2_X1 U14798 ( .A1(P2_EBX_REG_31__SCAN_IN), .A2(n11756), .ZN(n11757) );
  NOR2_X2 U14799 ( .A1(n11758), .A2(n11757), .ZN(n19049) );
  AOI22_X1 U14800 ( .A1(n11759), .A2(n19049), .B1(P2_REIP_REG_31__SCAN_IN), 
        .B2(n19091), .ZN(n11760) );
  AOI22_X1 U14801 ( .A1(n11723), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11766), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11768) );
  AOI21_X1 U14802 ( .B1(n12783), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A(
        n11769), .ZN(n11775) );
  AOI22_X1 U14803 ( .A1(n11770), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n11771), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11774) );
  AOI22_X1 U14804 ( .A1(n11772), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12788), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11773) );
  NAND3_X1 U14805 ( .A1(n11775), .A2(n11774), .A3(n11773), .ZN(n11784) );
  AOI22_X1 U14806 ( .A1(n11776), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n12789), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11782) );
  AOI22_X1 U14807 ( .A1(n11667), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n11668), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11781) );
  AOI22_X1 U14808 ( .A1(n11727), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11777), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11780) );
  AOI22_X1 U14809 ( .A1(n11778), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11680), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11779) );
  NAND4_X1 U14810 ( .A1(n11782), .A2(n11781), .A3(n11780), .A4(n11779), .ZN(
        n11783) );
  NOR2_X1 U14811 ( .A1(n11784), .A2(n11783), .ZN(n12331) );
  NAND2_X1 U14812 ( .A1(n10155), .A2(n11792), .ZN(n11800) );
  OAI22_X1 U14813 ( .A1(n19297), .A2(P2_STATE2_REG_3__SCAN_IN), .B1(n19924), 
        .B2(n19917), .ZN(n11785) );
  INV_X1 U14814 ( .A(n11785), .ZN(n11786) );
  AND2_X1 U14815 ( .A1(n11788), .A2(n19297), .ZN(n12970) );
  INV_X1 U14816 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n18929) );
  INV_X1 U14817 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n13576) );
  OAI21_X1 U14818 ( .B1(n19297), .B2(n13576), .A(n19917), .ZN(n11790) );
  AOI21_X1 U14819 ( .B1(n11792), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n11790), .ZN(n11791) );
  OAI21_X1 U14820 ( .B1(n11817), .B2(n18929), .A(n11791), .ZN(n13569) );
  INV_X1 U14821 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n19831) );
  NOR2_X1 U14822 ( .A1(n19297), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n11802) );
  AOI22_X1 U14823 ( .A1(n11802), .A2(P2_EAX_REG_1__SCAN_IN), .B1(n11792), .B2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n11793) );
  OAI21_X1 U14824 ( .B1(n11817), .B2(n19831), .A(n11793), .ZN(n11797) );
  OR2_X1 U14825 ( .A1(n12330), .A2(n11934), .ZN(n11796) );
  NAND2_X1 U14826 ( .A1(n11794), .A2(n19297), .ZN(n12382) );
  MUX2_X1 U14827 ( .A(n12382), .B(n19914), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n11795) );
  NAND2_X1 U14828 ( .A1(n11796), .A2(n11795), .ZN(n13550) );
  NOR2_X1 U14829 ( .A1(n13551), .A2(n13550), .ZN(n11799) );
  NOR2_X1 U14830 ( .A1(n13567), .A2(n11797), .ZN(n11798) );
  NAND2_X1 U14831 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n11801) );
  OAI211_X1 U14832 ( .C1(n11934), .C2(n12328), .A(n11801), .B(n11800), .ZN(
        n11804) );
  XNOR2_X1 U14833 ( .A(n11805), .B(n11804), .ZN(n13862) );
  INV_X1 U14834 ( .A(n11817), .ZN(n11931) );
  INV_X1 U14835 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n21092) );
  INV_X1 U14836 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n21090) );
  AOI22_X1 U14837 ( .A1(n11960), .A2(P2_EAX_REG_2__SCAN_IN), .B1(n11958), .B2(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n11803) );
  OAI21_X1 U14838 ( .B1(n11817), .B2(n21092), .A(n11803), .ZN(n13861) );
  NOR2_X1 U14839 ( .A1(n11805), .A2(n11804), .ZN(n11806) );
  INV_X1 U14840 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n11812) );
  AOI22_X1 U14841 ( .A1(n11958), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B1(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n11808) );
  NAND2_X1 U14842 ( .A1(n11960), .A2(P2_EAX_REG_3__SCAN_IN), .ZN(n11807) );
  AND2_X1 U14843 ( .A1(n11808), .A2(n11807), .ZN(n11811) );
  INV_X1 U14844 ( .A(n12059), .ZN(n11809) );
  OR2_X1 U14845 ( .A1(n11934), .A2(n11809), .ZN(n11810) );
  OAI211_X1 U14846 ( .C1(n11817), .C2(n11812), .A(n11811), .B(n11810), .ZN(
        n14003) );
  INV_X1 U14847 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n11816) );
  AOI22_X1 U14848 ( .A1(n11960), .A2(P2_EAX_REG_4__SCAN_IN), .B1(n11792), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n11815) );
  INV_X1 U14849 ( .A(n11813), .ZN(n12339) );
  OR2_X1 U14850 ( .A1(n11934), .A2(n12339), .ZN(n11814) );
  OAI211_X1 U14851 ( .C1(n11817), .C2(n11816), .A(n11815), .B(n11814), .ZN(
        n14008) );
  AOI22_X1 U14852 ( .A1(n11931), .A2(P2_REIP_REG_5__SCAN_IN), .B1(n11792), 
        .B2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n11819) );
  INV_X1 U14853 ( .A(n11934), .ZN(n11849) );
  AOI22_X1 U14854 ( .A1(n11849), .A2(n12096), .B1(n11960), .B2(
        P2_EAX_REG_5__SCAN_IN), .ZN(n11818) );
  NAND2_X1 U14855 ( .A1(n11819), .A2(n11818), .ZN(n14222) );
  NAND2_X1 U14856 ( .A1(n14223), .A2(n14222), .ZN(n14221) );
  OR2_X1 U14857 ( .A1(n11934), .A2(n12162), .ZN(n11820) );
  INV_X1 U14858 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n19838) );
  AOI22_X1 U14859 ( .A1(n11960), .A2(P2_EAX_REG_6__SCAN_IN), .B1(n11792), .B2(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n11821) );
  OAI21_X1 U14860 ( .B1(n11817), .B2(n19838), .A(n11821), .ZN(n14337) );
  NAND2_X1 U14861 ( .A1(n14336), .A2(n14337), .ZN(n11823) );
  OR2_X1 U14862 ( .A1(n11934), .A2(n12417), .ZN(n11822) );
  AOI22_X1 U14863 ( .A1(n11960), .A2(P2_EAX_REG_7__SCAN_IN), .B1(n11792), .B2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n11824) );
  OAI21_X1 U14864 ( .B1(n11817), .B2(n11530), .A(n11824), .ZN(n15725) );
  INV_X1 U14865 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n14190) );
  AOI22_X1 U14866 ( .A1(n11960), .A2(P2_EAX_REG_8__SCAN_IN), .B1(n11958), .B2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n11837) );
  AOI22_X1 U14867 ( .A1(n11723), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12781), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11828) );
  AOI22_X1 U14868 ( .A1(n12782), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n11771), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11827) );
  AOI22_X1 U14869 ( .A1(n11772), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11727), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11826) );
  AOI22_X1 U14870 ( .A1(n12788), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12783), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11825) );
  NAND4_X1 U14871 ( .A1(n11828), .A2(n11827), .A3(n11826), .A4(n11825), .ZN(
        n11834) );
  AOI22_X1 U14872 ( .A1(n11778), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n11680), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11832) );
  AOI22_X1 U14873 ( .A1(n11777), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n11770), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11831) );
  AOI22_X1 U14874 ( .A1(n11776), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n12789), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11830) );
  AOI22_X1 U14875 ( .A1(n11667), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n11668), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11829) );
  NAND4_X1 U14876 ( .A1(n11832), .A2(n11831), .A3(n11830), .A4(n11829), .ZN(
        n11833) );
  INV_X1 U14877 ( .A(n13883), .ZN(n11835) );
  OR2_X1 U14878 ( .A1(n11934), .A2(n11835), .ZN(n11836) );
  OAI211_X1 U14879 ( .C1(n11817), .C2(n14190), .A(n11837), .B(n11836), .ZN(
        n14186) );
  INV_X1 U14880 ( .A(n14186), .ZN(n11838) );
  AOI22_X1 U14881 ( .A1(n11931), .A2(P2_REIP_REG_9__SCAN_IN), .B1(n11960), 
        .B2(P2_EAX_REG_9__SCAN_IN), .ZN(n11851) );
  AOI22_X1 U14882 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n12781), .B1(
        n11772), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11842) );
  AOI22_X1 U14883 ( .A1(n11723), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11727), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11841) );
  AOI22_X1 U14884 ( .A1(n12782), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n11771), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11840) );
  AOI22_X1 U14885 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n11770), .B1(
        n12783), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11839) );
  NAND4_X1 U14886 ( .A1(n11842), .A2(n11841), .A3(n11840), .A4(n11839), .ZN(
        n11848) );
  AOI22_X1 U14887 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n11680), .B1(
        n11778), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11846) );
  AOI22_X1 U14888 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n11777), .B1(
        n12788), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11845) );
  AOI22_X1 U14889 ( .A1(n11776), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n12789), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11844) );
  AOI22_X1 U14890 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n11667), .B1(
        n11668), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11843) );
  NAND4_X1 U14891 ( .A1(n11846), .A2(n11845), .A3(n11844), .A4(n11843), .ZN(
        n11847) );
  AOI22_X1 U14892 ( .A1(n11849), .A2(n13921), .B1(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n11958), .ZN(n11850) );
  NAND2_X1 U14893 ( .A1(n11851), .A2(n11850), .ZN(n14040) );
  INV_X1 U14894 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n11864) );
  AOI22_X1 U14895 ( .A1(n11960), .A2(P2_EAX_REG_10__SCAN_IN), .B1(n11958), 
        .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n11863) );
  AOI22_X1 U14896 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n12781), .B1(
        n12782), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11855) );
  AOI22_X1 U14897 ( .A1(n11772), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11771), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11854) );
  AOI22_X1 U14898 ( .A1(n11723), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11727), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11853) );
  AOI22_X1 U14899 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n12788), .B1(
        n12783), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11852) );
  NAND4_X1 U14900 ( .A1(n11855), .A2(n11854), .A3(n11853), .A4(n11852), .ZN(
        n11861) );
  AOI22_X1 U14901 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n11778), .B1(
        n11680), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11859) );
  AOI22_X1 U14902 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n11777), .B1(
        n11770), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11858) );
  AOI22_X1 U14903 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n11776), .B1(
        n12789), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11857) );
  AOI22_X1 U14904 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n11667), .B1(
        n11668), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11856) );
  NAND4_X1 U14905 ( .A1(n11859), .A2(n11858), .A3(n11857), .A4(n11856), .ZN(
        n11860) );
  INV_X1 U14906 ( .A(n12701), .ZN(n13922) );
  OR2_X1 U14907 ( .A1(n11934), .A2(n13922), .ZN(n11862) );
  OAI211_X1 U14908 ( .C1(n11817), .C2(n11864), .A(n11863), .B(n11862), .ZN(
        n11865) );
  INV_X1 U14909 ( .A(n11865), .ZN(n15688) );
  NOR2_X2 U14910 ( .A1(n15689), .A2(n15688), .ZN(n15146) );
  AOI22_X1 U14911 ( .A1(n11960), .A2(P2_EAX_REG_11__SCAN_IN), .B1(n11958), 
        .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n11877) );
  AOI22_X1 U14912 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n12781), .B1(
        n11772), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11869) );
  AOI22_X1 U14913 ( .A1(n11723), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11727), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11868) );
  AOI22_X1 U14914 ( .A1(n12782), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n11771), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11867) );
  AOI22_X1 U14915 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n11770), .B1(
        n12783), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11866) );
  NAND4_X1 U14916 ( .A1(n11869), .A2(n11868), .A3(n11867), .A4(n11866), .ZN(
        n11875) );
  AOI22_X1 U14917 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n11778), .B1(
        n11680), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11873) );
  AOI22_X1 U14918 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n11777), .B1(
        n12788), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11872) );
  AOI22_X1 U14919 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n11776), .B1(
        n12789), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11871) );
  AOI22_X1 U14920 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n11667), .B1(
        n11668), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11870) );
  NAND4_X1 U14921 ( .A1(n11873), .A2(n11872), .A3(n11871), .A4(n11870), .ZN(
        n11874) );
  OR2_X1 U14922 ( .A1(n11934), .A2(n12703), .ZN(n11876) );
  OAI211_X1 U14923 ( .C1(n11817), .C2(n11878), .A(n11877), .B(n11876), .ZN(
        n15147) );
  NAND2_X1 U14924 ( .A1(n15146), .A2(n15147), .ZN(n14263) );
  INV_X1 U14925 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n11892) );
  AOI22_X1 U14926 ( .A1(n11960), .A2(P2_EAX_REG_12__SCAN_IN), .B1(n11958), 
        .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n11891) );
  AOI22_X1 U14927 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n11723), .B1(
        n12782), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11882) );
  AOI22_X1 U14928 ( .A1(n12781), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n11771), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11881) );
  AOI22_X1 U14929 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n11772), .B1(
        n11727), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11880) );
  AOI22_X1 U14930 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n11770), .B1(
        n12788), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11879) );
  NAND4_X1 U14931 ( .A1(n11882), .A2(n11881), .A3(n11880), .A4(n11879), .ZN(
        n11888) );
  AOI22_X1 U14932 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n11778), .B1(
        n11680), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11886) );
  AOI22_X1 U14933 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n11777), .B1(
        n12783), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11885) );
  AOI22_X1 U14934 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n11776), .B1(
        n12789), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11884) );
  AOI22_X1 U14935 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n11667), .B1(
        n11668), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11883) );
  NAND4_X1 U14936 ( .A1(n11886), .A2(n11885), .A3(n11884), .A4(n11883), .ZN(
        n11887) );
  INV_X1 U14937 ( .A(n14020), .ZN(n11889) );
  OR2_X1 U14938 ( .A1(n11934), .A2(n11889), .ZN(n11890) );
  OAI211_X1 U14939 ( .C1(n11817), .C2(n11892), .A(n11891), .B(n11890), .ZN(
        n14265) );
  INV_X1 U14940 ( .A(n14265), .ZN(n11893) );
  AOI22_X1 U14941 ( .A1(n11960), .A2(P2_EAX_REG_13__SCAN_IN), .B1(n11958), 
        .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n11906) );
  AOI22_X1 U14942 ( .A1(n12781), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11772), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11897) );
  AOI22_X1 U14943 ( .A1(n11723), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11727), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11896) );
  AOI22_X1 U14944 ( .A1(n12782), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n11771), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11895) );
  AOI22_X1 U14945 ( .A1(n11770), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n12783), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11894) );
  NAND4_X1 U14946 ( .A1(n11897), .A2(n11896), .A3(n11895), .A4(n11894), .ZN(
        n11903) );
  AOI22_X1 U14947 ( .A1(n11778), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11680), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11901) );
  AOI22_X1 U14948 ( .A1(n12788), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11777), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11900) );
  AOI22_X1 U14949 ( .A1(n11776), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n12789), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11899) );
  AOI22_X1 U14950 ( .A1(n11667), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11668), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11898) );
  NAND4_X1 U14951 ( .A1(n11901), .A2(n11900), .A3(n11899), .A4(n11898), .ZN(
        n11902) );
  INV_X1 U14952 ( .A(n14064), .ZN(n11904) );
  OR2_X1 U14953 ( .A1(n11934), .A2(n11904), .ZN(n11905) );
  OAI211_X1 U14954 ( .C1(n11817), .C2(n15449), .A(n11906), .B(n11905), .ZN(
        n15647) );
  NAND2_X1 U14955 ( .A1(n14266), .A2(n15647), .ZN(n15648) );
  INV_X1 U14956 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n11919) );
  AOI22_X1 U14957 ( .A1(n11960), .A2(P2_EAX_REG_14__SCAN_IN), .B1(n11958), 
        .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n11918) );
  AOI22_X1 U14958 ( .A1(n11723), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11727), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11910) );
  AOI22_X1 U14959 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n12781), .B1(
        n11772), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11909) );
  AOI22_X1 U14960 ( .A1(n12782), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n11771), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11908) );
  AOI22_X1 U14961 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n11770), .B1(
        n12783), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11907) );
  NAND4_X1 U14962 ( .A1(n11910), .A2(n11909), .A3(n11908), .A4(n11907), .ZN(
        n11916) );
  AOI22_X1 U14963 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n11778), .B1(
        n11680), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11914) );
  AOI22_X1 U14964 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n11777), .B1(
        n12788), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11913) );
  AOI22_X1 U14965 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n12789), .B1(
        n11668), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11912) );
  AOI22_X1 U14966 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n11667), .B1(
        n11776), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11911) );
  NAND4_X1 U14967 ( .A1(n11914), .A2(n11913), .A3(n11912), .A4(n11911), .ZN(
        n11915) );
  INV_X1 U14968 ( .A(n14140), .ZN(n12704) );
  OR2_X1 U14969 ( .A1(n11934), .A2(n12704), .ZN(n11917) );
  OAI211_X1 U14970 ( .C1(n11817), .C2(n11919), .A(n11918), .B(n11917), .ZN(
        n15631) );
  INV_X1 U14971 ( .A(n15631), .ZN(n11920) );
  AOI22_X1 U14972 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n12781), .B1(
        n11772), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11924) );
  AOI22_X1 U14973 ( .A1(n11723), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11727), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11923) );
  AOI22_X1 U14974 ( .A1(n12782), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n11771), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11922) );
  AOI22_X1 U14975 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n11770), .B1(
        n12783), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11921) );
  NAND4_X1 U14976 ( .A1(n11924), .A2(n11923), .A3(n11922), .A4(n11921), .ZN(
        n11930) );
  AOI22_X1 U14977 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n11778), .B1(
        n11680), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11928) );
  AOI22_X1 U14978 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n11777), .B1(
        n12788), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11927) );
  AOI22_X1 U14979 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n11776), .B1(
        n12789), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11926) );
  AOI22_X1 U14980 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n11667), .B1(
        n11668), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11925) );
  NAND4_X1 U14981 ( .A1(n11928), .A2(n11927), .A3(n11926), .A4(n11925), .ZN(
        n11929) );
  NAND2_X1 U14982 ( .A1(n11931), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n11933) );
  AOI22_X1 U14983 ( .A1(n11960), .A2(P2_EAX_REG_15__SCAN_IN), .B1(n11958), 
        .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n11932) );
  OAI211_X1 U14984 ( .C1(n12705), .C2(n11934), .A(n11933), .B(n11932), .ZN(
        n16312) );
  NAND2_X1 U14985 ( .A1(n11931), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n11936) );
  AOI22_X1 U14986 ( .A1(n11960), .A2(P2_EAX_REG_16__SCAN_IN), .B1(n11958), 
        .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n11935) );
  AOI22_X1 U14987 ( .A1(n11960), .A2(P2_EAX_REG_17__SCAN_IN), .B1(n11792), 
        .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n11937) );
  OAI21_X1 U14988 ( .B1(n11817), .B2(n21095), .A(n11937), .ZN(n14315) );
  INV_X1 U14989 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n15411) );
  AOI22_X1 U14990 ( .A1(n11960), .A2(P2_EAX_REG_18__SCAN_IN), .B1(n11792), 
        .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n11938) );
  OAI21_X1 U14991 ( .B1(n11817), .B2(n15411), .A(n11938), .ZN(n11939) );
  INV_X1 U14992 ( .A(n11939), .ZN(n15598) );
  AOI22_X1 U14993 ( .A1(n11960), .A2(P2_EAX_REG_19__SCAN_IN), .B1(n11792), 
        .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n11940) );
  OAI21_X1 U14994 ( .B1(n11817), .B2(n19854), .A(n11940), .ZN(n11941) );
  INV_X1 U14995 ( .A(n11941), .ZN(n15280) );
  AOI22_X1 U14996 ( .A1(n11960), .A2(P2_EAX_REG_20__SCAN_IN), .B1(n11792), 
        .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n11942) );
  OAI21_X1 U14997 ( .B1(n11817), .B2(n19856), .A(n11942), .ZN(n11943) );
  INV_X1 U14998 ( .A(n11943), .ZN(n15572) );
  AOI22_X1 U14999 ( .A1(n11960), .A2(P2_EAX_REG_21__SCAN_IN), .B1(n11958), 
        .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n11944) );
  OAI21_X1 U15000 ( .B1(n11817), .B2(n21126), .A(n11944), .ZN(n13350) );
  AOI22_X1 U15001 ( .A1(n11960), .A2(P2_EAX_REG_22__SCAN_IN), .B1(n11958), 
        .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n11945) );
  OAI21_X1 U15002 ( .B1(n11817), .B2(n15861), .A(n11945), .ZN(n15548) );
  AOI22_X1 U15003 ( .A1(n11960), .A2(P2_EAX_REG_23__SCAN_IN), .B1(n11958), 
        .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n11946) );
  OAI21_X1 U15004 ( .B1(n11817), .B2(n19860), .A(n11946), .ZN(n13363) );
  NAND2_X1 U15005 ( .A1(n11931), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n11948) );
  AOI22_X1 U15006 ( .A1(n11960), .A2(P2_EAX_REG_24__SCAN_IN), .B1(n11958), 
        .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n11947) );
  AND2_X1 U15007 ( .A1(n11948), .A2(n11947), .ZN(n15127) );
  OR2_X2 U15008 ( .A1(n13362), .A2(n15127), .ZN(n15129) );
  NAND2_X1 U15009 ( .A1(n11931), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n11950) );
  AOI22_X1 U15010 ( .A1(n11960), .A2(P2_EAX_REG_25__SCAN_IN), .B1(n11958), 
        .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n11949) );
  AND2_X1 U15011 ( .A1(n11950), .A2(n11949), .ZN(n15115) );
  AOI22_X1 U15012 ( .A1(n11960), .A2(P2_EAX_REG_26__SCAN_IN), .B1(n11958), 
        .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n11951) );
  OAI21_X1 U15013 ( .B1(n11817), .B2(n19866), .A(n11951), .ZN(n15251) );
  NAND2_X1 U15014 ( .A1(n11931), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n11953) );
  AOI22_X1 U15015 ( .A1(n11960), .A2(P2_EAX_REG_27__SCAN_IN), .B1(n11958), 
        .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n11952) );
  AND2_X1 U15016 ( .A1(n11953), .A2(n11952), .ZN(n13337) );
  NAND2_X1 U15017 ( .A1(n11931), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n11955) );
  AOI22_X1 U15018 ( .A1(n11960), .A2(P2_EAX_REG_28__SCAN_IN), .B1(n11958), 
        .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n11954) );
  AND2_X1 U15019 ( .A1(n11955), .A2(n11954), .ZN(n15094) );
  NAND2_X1 U15020 ( .A1(n11931), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n11957) );
  AOI22_X1 U15021 ( .A1(n11960), .A2(P2_EAX_REG_29__SCAN_IN), .B1(n11958), 
        .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n11956) );
  AND2_X1 U15022 ( .A1(n11957), .A2(n11956), .ZN(n12488) );
  AOI22_X1 U15023 ( .A1(n11960), .A2(P2_EAX_REG_30__SCAN_IN), .B1(n11958), 
        .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n11959) );
  OAI21_X1 U15024 ( .B1(n11817), .B2(n12509), .A(n11959), .ZN(n12517) );
  NAND2_X1 U15025 ( .A1(n12516), .A2(n12517), .ZN(n12521) );
  INV_X1 U15026 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n19874) );
  AOI22_X1 U15027 ( .A1(n11960), .A2(P2_EAX_REG_31__SCAN_IN), .B1(n11792), 
        .B2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n11961) );
  OAI21_X1 U15028 ( .B1(n11817), .B2(n19874), .A(n11961), .ZN(n11962) );
  AND2_X1 U15029 ( .A1(n19271), .A2(n16370), .ZN(n16389) );
  AND3_X2 U15030 ( .A1(n16390), .A2(n16389), .A3(n11964), .ZN(n19241) );
  NOR2_X1 U15031 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n16372), .ZN(n16388) );
  NAND3_X1 U15032 ( .A1(n11967), .A2(n11966), .A3(n11965), .ZN(P2_U2824) );
  NAND2_X1 U15033 ( .A1(n11985), .A2(n11984), .ZN(n11974) );
  INV_X1 U15034 ( .A(n11971), .ZN(n11973) );
  NAND2_X1 U15035 ( .A1(n11969), .A2(n11968), .ZN(n11970) );
  AND2_X1 U15036 ( .A1(n11973), .A2(n11970), .ZN(n11977) );
  NAND2_X1 U15037 ( .A1(n11971), .A2(n11970), .ZN(n11972) );
  INV_X1 U15038 ( .A(n11982), .ZN(n11983) );
  XNOR2_X2 U15039 ( .A(n11989), .B(n11983), .ZN(n12673) );
  XNOR2_X1 U15040 ( .A(n11985), .B(n11984), .ZN(n11986) );
  INV_X1 U15041 ( .A(n12071), .ZN(n14031) );
  NAND2_X1 U15042 ( .A1(n14031), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n11993) );
  INV_X2 U15043 ( .A(n11987), .ZN(n13628) );
  INV_X1 U15044 ( .A(n19508), .ZN(n19511) );
  NAND2_X1 U15045 ( .A1(n19511), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n11992) );
  BUF_X4 U15046 ( .A(n12672), .Z(n13842) );
  INV_X1 U15047 ( .A(n11998), .ZN(n11990) );
  NAND2_X1 U15048 ( .A1(n13842), .A2(n12019), .ZN(n19415) );
  INV_X1 U15049 ( .A(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11991) );
  NAND3_X1 U15050 ( .A1(n11993), .A2(n11992), .A3(n10260), .ZN(n12003) );
  NAND2_X2 U15051 ( .A1(n12021), .A2(n13628), .ZN(n12072) );
  INV_X1 U15052 ( .A(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12001) );
  INV_X1 U15053 ( .A(n12672), .ZN(n14053) );
  NAND3_X2 U15054 ( .A1(n13628), .A2(n12012), .A3(n14053), .ZN(n12085) );
  INV_X1 U15055 ( .A(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11996) );
  INV_X1 U15056 ( .A(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11995) );
  INV_X1 U15057 ( .A(n11997), .ZN(n12000) );
  INV_X1 U15058 ( .A(n19542), .ZN(n19545) );
  NAND2_X1 U15059 ( .A1(n19545), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n11999) );
  OAI211_X1 U15060 ( .C1(n12072), .C2(n12001), .A(n12000), .B(n11999), .ZN(
        n12002) );
  NOR2_X1 U15061 ( .A1(n12003), .A2(n12002), .ZN(n12027) );
  INV_X1 U15062 ( .A(n14124), .ZN(n14130) );
  INV_X1 U15063 ( .A(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12005) );
  OAI21_X1 U15064 ( .B1(n19358), .B2(n12005), .A(n13427), .ZN(n12006) );
  INV_X1 U15065 ( .A(n12064), .ZN(n19579) );
  NAND2_X1 U15066 ( .A1(n19579), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n12010) );
  INV_X1 U15067 ( .A(n12063), .ZN(n19697) );
  NAND2_X1 U15068 ( .A1(n19697), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n12009) );
  INV_X1 U15069 ( .A(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12017) );
  INV_X1 U15070 ( .A(n12014), .ZN(n12015) );
  OR2_X2 U15071 ( .A1(n12015), .A2(n13842), .ZN(n12080) );
  INV_X1 U15072 ( .A(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12016) );
  INV_X1 U15073 ( .A(n12018), .ZN(n12025) );
  NAND2_X1 U15074 ( .A1(n14053), .A2(n12019), .ZN(n12148) );
  INV_X1 U15075 ( .A(n12148), .ZN(n19660) );
  NAND2_X1 U15076 ( .A1(n19660), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n12024) );
  INV_X1 U15077 ( .A(n19452), .ZN(n19444) );
  NAND2_X1 U15078 ( .A1(n19444), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n12023) );
  INV_X1 U15079 ( .A(n12141), .ZN(n19384) );
  NAND2_X1 U15080 ( .A1(n19384), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n12022) );
  NAND3_X1 U15081 ( .A1(n12027), .A2(n10262), .A3(n12026), .ZN(n12029) );
  OR2_X1 U15082 ( .A1(n12331), .A2(n13427), .ZN(n12329) );
  INV_X1 U15083 ( .A(n12329), .ZN(n15465) );
  INV_X1 U15084 ( .A(n12330), .ZN(n12028) );
  NAND2_X1 U15085 ( .A1(n15465), .A2(n12028), .ZN(n12327) );
  AND2_X2 U15086 ( .A1(n12029), .A2(n9926), .ZN(n12106) );
  INV_X1 U15087 ( .A(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12031) );
  INV_X1 U15088 ( .A(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12030) );
  OAI22_X1 U15089 ( .A1(n12031), .A2(n12063), .B1(n12064), .B2(n12030), .ZN(
        n12035) );
  INV_X1 U15090 ( .A(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12033) );
  INV_X1 U15091 ( .A(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12032) );
  NOR2_X1 U15092 ( .A1(n12035), .A2(n12034), .ZN(n12056) );
  INV_X1 U15093 ( .A(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n14038) );
  INV_X1 U15094 ( .A(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12036) );
  OAI22_X1 U15095 ( .A1(n14038), .A2(n12071), .B1(n19508), .B2(n12036), .ZN(
        n12040) );
  INV_X1 U15096 ( .A(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12038) );
  INV_X1 U15097 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12037) );
  OAI22_X1 U15098 ( .A1(n12038), .A2(n12141), .B1(n12072), .B2(n12037), .ZN(
        n12039) );
  NOR2_X1 U15099 ( .A1(n12040), .A2(n12039), .ZN(n12055) );
  INV_X1 U15100 ( .A(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12042) );
  INV_X1 U15101 ( .A(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12041) );
  OAI22_X1 U15102 ( .A1(n12042), .A2(n19482), .B1(n12080), .B2(n12041), .ZN(
        n12046) );
  INV_X1 U15103 ( .A(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12044) );
  INV_X1 U15104 ( .A(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12043) );
  OAI22_X1 U15105 ( .A1(n12044), .A2(n19415), .B1(n12148), .B2(n12043), .ZN(
        n12045) );
  NOR2_X1 U15106 ( .A1(n12046), .A2(n12045), .ZN(n12054) );
  INV_X1 U15107 ( .A(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12048) );
  INV_X1 U15108 ( .A(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12047) );
  OAI22_X1 U15109 ( .A1(n19304), .A2(n12048), .B1(n12085), .B2(n12047), .ZN(
        n12052) );
  INV_X1 U15110 ( .A(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12050) );
  INV_X1 U15111 ( .A(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12049) );
  OAI22_X1 U15112 ( .A1(n19542), .A2(n12050), .B1(n19358), .B2(n12049), .ZN(
        n12051) );
  NOR2_X1 U15113 ( .A1(n12052), .A2(n12051), .ZN(n12053) );
  NAND4_X1 U15114 ( .A1(n12056), .A2(n12055), .A3(n12054), .A4(n12053), .ZN(
        n12057) );
  NAND2_X1 U15115 ( .A1(n12057), .A2(n13427), .ZN(n12061) );
  INV_X1 U15116 ( .A(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12066) );
  INV_X1 U15117 ( .A(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12065) );
  OAI22_X1 U15118 ( .A1(n12066), .A2(n12063), .B1(n12064), .B2(n12065), .ZN(
        n12070) );
  INV_X1 U15119 ( .A(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12068) );
  INV_X1 U15120 ( .A(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12067) );
  OAI22_X1 U15121 ( .A1(n12068), .A2(n19452), .B1(n14124), .B2(n12067), .ZN(
        n12069) );
  NOR2_X1 U15122 ( .A1(n12070), .A2(n12069), .ZN(n12095) );
  INV_X1 U15123 ( .A(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12073) );
  INV_X1 U15124 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13846) );
  OAI22_X1 U15125 ( .A1(n12073), .A2(n12071), .B1(n12072), .B2(n13846), .ZN(
        n12077) );
  INV_X1 U15126 ( .A(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12075) );
  INV_X1 U15127 ( .A(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12074) );
  OAI22_X1 U15128 ( .A1(n12075), .A2(n19508), .B1(n12141), .B2(n12074), .ZN(
        n12076) );
  NOR2_X1 U15129 ( .A1(n12077), .A2(n12076), .ZN(n12094) );
  INV_X1 U15130 ( .A(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12079) );
  INV_X1 U15131 ( .A(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12078) );
  OAI22_X1 U15132 ( .A1(n12079), .A2(n19415), .B1(n12148), .B2(n12078), .ZN(
        n12084) );
  INV_X1 U15133 ( .A(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12082) );
  INV_X1 U15134 ( .A(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12081) );
  OAI22_X1 U15135 ( .A1(n12082), .A2(n19482), .B1(n12080), .B2(n12081), .ZN(
        n12083) );
  NOR2_X1 U15136 ( .A1(n12084), .A2(n12083), .ZN(n12093) );
  INV_X1 U15137 ( .A(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12087) );
  INV_X1 U15138 ( .A(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12086) );
  OAI22_X1 U15139 ( .A1(n12087), .A2(n19542), .B1(n12085), .B2(n12086), .ZN(
        n12091) );
  INV_X1 U15140 ( .A(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12089) );
  INV_X1 U15141 ( .A(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12088) );
  OAI22_X1 U15142 ( .A1(n12089), .A2(n19304), .B1(n19358), .B2(n12088), .ZN(
        n12090) );
  NOR2_X1 U15143 ( .A1(n12091), .A2(n12090), .ZN(n12092) );
  NAND4_X1 U15144 ( .A1(n12095), .A2(n12094), .A3(n12093), .A4(n12092), .ZN(
        n12099) );
  INV_X1 U15145 ( .A(n12096), .ZN(n12097) );
  NAND2_X1 U15146 ( .A1(n12097), .A2(n19271), .ZN(n12098) );
  INV_X1 U15147 ( .A(n12100), .ZN(n12101) );
  OAI21_X1 U15148 ( .B1(n12104), .B2(n12103), .A(n12167), .ZN(n19075) );
  OAI21_X2 U15149 ( .B1(n12347), .B2(n12102), .A(n19075), .ZN(n12130) );
  XNOR2_X1 U15150 ( .A(n12130), .B(n14226), .ZN(n14215) );
  INV_X1 U15151 ( .A(n12126), .ZN(n12111) );
  INV_X1 U15152 ( .A(n12107), .ZN(n12109) );
  NAND2_X1 U15153 ( .A1(n12109), .A2(n10060), .ZN(n12110) );
  NAND2_X1 U15154 ( .A1(n12111), .A2(n12110), .ZN(n14057) );
  AND2_X1 U15155 ( .A1(n14057), .A2(n14095), .ZN(n12112) );
  NAND2_X1 U15156 ( .A1(n12123), .A2(n12112), .ZN(n14086) );
  INV_X1 U15157 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n15749) );
  OAI21_X1 U15158 ( .B1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n19924), .A(
        n12113), .ZN(n12300) );
  MUX2_X1 U15159 ( .A(n12300), .B(n12331), .S(n12114), .Z(n12286) );
  MUX2_X1 U15160 ( .A(n12286), .B(n12115), .S(n12412), .Z(n19094) );
  NOR2_X1 U15161 ( .A1(n19094), .A2(n11481), .ZN(n13548) );
  NAND3_X1 U15162 ( .A1(n12412), .A2(P2_EBX_REG_1__SCAN_IN), .A3(
        P2_EBX_REG_0__SCAN_IN), .ZN(n12116) );
  NAND2_X1 U15163 ( .A1(n12118), .A2(n12116), .ZN(n14362) );
  INV_X1 U15164 ( .A(n14362), .ZN(n13547) );
  NAND2_X1 U15165 ( .A1(n13548), .A2(n13547), .ZN(n12117) );
  NOR2_X1 U15166 ( .A1(n13548), .A2(n13547), .ZN(n13546) );
  AOI21_X1 U15167 ( .B1(n15749), .B2(n12117), .A(n13546), .ZN(n14527) );
  XNOR2_X1 U15168 ( .A(n12119), .B(n12118), .ZN(n14240) );
  XNOR2_X1 U15169 ( .A(n14240), .B(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n14528) );
  NAND2_X1 U15170 ( .A1(n14527), .A2(n14528), .ZN(n12122) );
  INV_X1 U15171 ( .A(n14240), .ZN(n12120) );
  NAND2_X1 U15172 ( .A1(n12120), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12121) );
  NAND2_X1 U15173 ( .A1(n12122), .A2(n12121), .ZN(n14087) );
  NAND2_X1 U15174 ( .A1(n14086), .A2(n14087), .ZN(n14085) );
  NAND2_X1 U15175 ( .A1(n12123), .A2(n14057), .ZN(n12124) );
  NAND2_X1 U15176 ( .A1(n14085), .A2(n14089), .ZN(n14109) );
  XNOR2_X1 U15177 ( .A(n12126), .B(n12125), .ZN(n14156) );
  XNOR2_X1 U15178 ( .A(n14156), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n14108) );
  NAND2_X1 U15179 ( .A1(n14109), .A2(n14108), .ZN(n12129) );
  INV_X1 U15180 ( .A(n14156), .ZN(n12127) );
  NAND2_X1 U15181 ( .A1(n12127), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12128) );
  NAND2_X1 U15182 ( .A1(n12129), .A2(n12128), .ZN(n14216) );
  NAND2_X1 U15183 ( .A1(n12130), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12131) );
  INV_X1 U15184 ( .A(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12133) );
  INV_X1 U15185 ( .A(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12132) );
  OAI22_X1 U15186 ( .A1(n12133), .A2(n12063), .B1(n19452), .B2(n12132), .ZN(
        n12137) );
  INV_X1 U15187 ( .A(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12135) );
  INV_X1 U15188 ( .A(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12134) );
  OAI22_X1 U15189 ( .A1(n12135), .A2(n12064), .B1(n14124), .B2(n12134), .ZN(
        n12136) );
  NOR2_X1 U15190 ( .A1(n12137), .A2(n12136), .ZN(n12161) );
  INV_X1 U15191 ( .A(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12139) );
  INV_X1 U15192 ( .A(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12138) );
  OAI22_X1 U15193 ( .A1(n12139), .A2(n12071), .B1(n12072), .B2(n12138), .ZN(
        n12144) );
  INV_X1 U15194 ( .A(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12142) );
  INV_X1 U15195 ( .A(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12140) );
  OAI22_X1 U15196 ( .A1(n12142), .A2(n19508), .B1(n12141), .B2(n12140), .ZN(
        n12143) );
  NOR2_X1 U15197 ( .A1(n12144), .A2(n12143), .ZN(n12160) );
  INV_X1 U15198 ( .A(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12146) );
  INV_X1 U15199 ( .A(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12145) );
  OAI22_X1 U15200 ( .A1(n12146), .A2(n19415), .B1(n19482), .B2(n12145), .ZN(
        n12151) );
  INV_X1 U15201 ( .A(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12149) );
  INV_X1 U15202 ( .A(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12147) );
  OAI22_X1 U15203 ( .A1(n12149), .A2(n12080), .B1(n12148), .B2(n12147), .ZN(
        n12150) );
  NOR2_X1 U15204 ( .A1(n12151), .A2(n12150), .ZN(n12159) );
  INV_X1 U15205 ( .A(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12153) );
  INV_X1 U15206 ( .A(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12152) );
  OAI22_X1 U15207 ( .A1(n12153), .A2(n19542), .B1(n12085), .B2(n12152), .ZN(
        n12157) );
  INV_X1 U15208 ( .A(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12155) );
  INV_X1 U15209 ( .A(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12154) );
  OAI22_X1 U15210 ( .A1(n12155), .A2(n19304), .B1(n19358), .B2(n12154), .ZN(
        n12156) );
  NOR2_X1 U15211 ( .A1(n12157), .A2(n12156), .ZN(n12158) );
  NAND4_X1 U15212 ( .A1(n12161), .A2(n12160), .A3(n12159), .A4(n12158), .ZN(
        n12164) );
  NAND2_X1 U15213 ( .A1(n12162), .A2(n12058), .ZN(n12163) );
  XNOR2_X1 U15214 ( .A(n12167), .B(n12166), .ZN(n19059) );
  NOR2_X1 U15215 ( .A1(n19286), .A2(n10078), .ZN(n12170) );
  AND2_X1 U15216 ( .A1(n12175), .A2(n12170), .ZN(n12171) );
  OR2_X1 U15217 ( .A1(n12169), .A2(n12171), .ZN(n14183) );
  NOR2_X1 U15218 ( .A1(n14183), .A2(n12417), .ZN(n12181) );
  NAND2_X1 U15219 ( .A1(n12181), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n16280) );
  OR2_X1 U15220 ( .A1(n12173), .A2(n12172), .ZN(n12174) );
  AND2_X1 U15221 ( .A1(n12175), .A2(n12174), .ZN(n19050) );
  NAND2_X1 U15222 ( .A1(n19050), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16281) );
  AND2_X1 U15223 ( .A1(n16280), .A2(n16281), .ZN(n15692) );
  NAND2_X1 U15224 ( .A1(n12176), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n15456) );
  AND2_X1 U15225 ( .A1(n15692), .A2(n15456), .ZN(n12187) );
  NAND2_X1 U15226 ( .A1(n12412), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n12177) );
  OAI21_X1 U15227 ( .B1(n12178), .B2(n12177), .A(n12269), .ZN(n12179) );
  OR2_X1 U15228 ( .A1(n12191), .A2(n12179), .ZN(n19036) );
  OAI21_X1 U15229 ( .B1(n19036), .B2(n12417), .A(n12180), .ZN(n15699) );
  INV_X1 U15230 ( .A(n12181), .ZN(n12182) );
  NAND2_X1 U15231 ( .A1(n12182), .A2(n12364), .ZN(n16279) );
  INV_X1 U15232 ( .A(n19050), .ZN(n12183) );
  NAND2_X1 U15233 ( .A1(n12183), .A2(n15730), .ZN(n16283) );
  AND2_X1 U15234 ( .A1(n16279), .A2(n16283), .ZN(n15694) );
  NOR2_X1 U15235 ( .A1(n19286), .A2(n12184), .ZN(n12185) );
  XNOR2_X1 U15236 ( .A(n12169), .B(n12185), .ZN(n14044) );
  NAND2_X1 U15237 ( .A1(n14044), .A2(n12102), .ZN(n12186) );
  NAND2_X1 U15238 ( .A1(n12186), .A2(n15712), .ZN(n15717) );
  AND2_X1 U15239 ( .A1(n12102), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n12188) );
  AND2_X1 U15240 ( .A1(n14044), .A2(n12188), .ZN(n15696) );
  NAND2_X1 U15241 ( .A1(n12102), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n12189) );
  NOR2_X1 U15242 ( .A1(n19036), .A2(n12189), .ZN(n15698) );
  NAND2_X1 U15243 ( .A1(n12412), .A2(P2_EBX_REG_11__SCAN_IN), .ZN(n12190) );
  OR2_X1 U15244 ( .A1(n12191), .A2(n12190), .ZN(n15151) );
  NOR2_X1 U15245 ( .A1(n12192), .A2(n12417), .ZN(n12193) );
  NAND2_X1 U15246 ( .A1(n15151), .A2(n12193), .ZN(n15671) );
  NAND2_X1 U15247 ( .A1(P2_EBX_REG_12__SCAN_IN), .A2(n12194), .ZN(n12195) );
  NOR2_X1 U15248 ( .A1(n19286), .A2(n12195), .ZN(n12196) );
  OR2_X1 U15249 ( .A1(n12213), .A2(n12196), .ZN(n14275) );
  NOR2_X1 U15250 ( .A1(n14275), .A2(n12417), .ZN(n12214) );
  NAND2_X1 U15251 ( .A1(n12214), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n15661) );
  NOR2_X1 U15252 ( .A1(n19286), .A2(n15213), .ZN(n12197) );
  AOI21_X1 U15253 ( .B1(n9872), .B2(n12197), .A(n10076), .ZN(n12198) );
  NAND2_X1 U15254 ( .A1(n12250), .A2(n12198), .ZN(n13348) );
  NOR2_X1 U15255 ( .A1(n12236), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15370) );
  NOR2_X1 U15256 ( .A1(n12200), .A2(n14146), .ZN(n12199) );
  MUX2_X1 U15257 ( .A(n12200), .B(n12199), .S(n12412), .Z(n12202) );
  NAND2_X1 U15258 ( .A1(n12200), .A2(n14146), .ZN(n12218) );
  INV_X1 U15259 ( .A(n12218), .ZN(n12201) );
  NOR2_X1 U15260 ( .A1(n12202), .A2(n12201), .ZN(n19017) );
  NAND2_X1 U15261 ( .A1(n19017), .A2(n12102), .ZN(n12241) );
  INV_X1 U15262 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n15638) );
  NAND3_X1 U15263 ( .A1(n12219), .A2(P2_EBX_REG_16__SCAN_IN), .A3(n12412), 
        .ZN(n12203) );
  OAI211_X1 U15264 ( .C1(n12219), .C2(P2_EBX_REG_16__SCAN_IN), .A(n12203), .B(
        n12269), .ZN(n18993) );
  INV_X1 U15265 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15614) );
  OAI21_X1 U15266 ( .B1(n18993), .B2(n12417), .A(n15614), .ZN(n12205) );
  NAND2_X1 U15267 ( .A1(n12102), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12204) );
  OR2_X1 U15268 ( .A1(n18993), .A2(n12204), .ZN(n15364) );
  NAND2_X1 U15269 ( .A1(n12205), .A2(n15364), .ZN(n15849) );
  INV_X1 U15270 ( .A(n12206), .ZN(n12208) );
  NAND2_X1 U15271 ( .A1(n12208), .A2(n10080), .ZN(n12209) );
  NAND2_X1 U15272 ( .A1(n12225), .A2(n12209), .ZN(n18978) );
  OR2_X1 U15273 ( .A1(n18978), .A2(n12417), .ZN(n12210) );
  NAND2_X1 U15274 ( .A1(n12210), .A2(n15622), .ZN(n15366) );
  INV_X1 U15275 ( .A(n12211), .ZN(n12212) );
  XNOR2_X1 U15276 ( .A(n12213), .B(n12212), .ZN(n19027) );
  NAND2_X1 U15277 ( .A1(n19027), .A2(n12102), .ZN(n12240) );
  NAND2_X1 U15278 ( .A1(n12240), .A2(n21086), .ZN(n15443) );
  INV_X1 U15279 ( .A(n12214), .ZN(n12215) );
  INV_X1 U15280 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n15659) );
  NAND2_X1 U15281 ( .A1(n12215), .A2(n15659), .ZN(n15660) );
  NOR2_X1 U15282 ( .A1(n19286), .A2(n12216), .ZN(n12217) );
  NAND2_X1 U15283 ( .A1(n12218), .A2(n12217), .ZN(n12220) );
  NAND2_X1 U15284 ( .A1(n12220), .A2(n12219), .ZN(n18999) );
  OR2_X1 U15285 ( .A1(n18999), .A2(n12417), .ZN(n12222) );
  INV_X1 U15286 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n12221) );
  NAND2_X1 U15287 ( .A1(n12222), .A2(n12221), .ZN(n15431) );
  NAND4_X1 U15288 ( .A1(n15366), .A2(n15443), .A3(n15660), .A4(n15431), .ZN(
        n12223) );
  NOR4_X1 U15289 ( .A1(n15370), .A2(n15626), .A3(n15849), .A4(n12223), .ZN(
        n12235) );
  NAND2_X1 U15290 ( .A1(n12225), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n12224) );
  MUX2_X1 U15291 ( .A(n12225), .B(n12224), .S(n12412), .Z(n12226) );
  OR2_X1 U15292 ( .A1(n12225), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n12230) );
  NAND2_X1 U15293 ( .A1(n12226), .A2(n12230), .ZN(n18970) );
  OR2_X1 U15294 ( .A1(n18970), .A2(n12417), .ZN(n12227) );
  INV_X1 U15295 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n15414) );
  NAND2_X1 U15296 ( .A1(n12227), .A2(n15414), .ZN(n15408) );
  NOR2_X1 U15297 ( .A1(n19286), .A2(n12228), .ZN(n12229) );
  NAND2_X1 U15298 ( .A1(n12230), .A2(n12229), .ZN(n12231) );
  NAND2_X1 U15299 ( .A1(n12231), .A2(n12234), .ZN(n18953) );
  OR2_X1 U15300 ( .A1(n18953), .A2(n12417), .ZN(n12232) );
  INV_X1 U15301 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15401) );
  NAND2_X1 U15302 ( .A1(n12232), .A2(n15401), .ZN(n15394) );
  NAND2_X1 U15303 ( .A1(n15408), .A2(n15394), .ZN(n15383) );
  NAND2_X1 U15304 ( .A1(n12412), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n12233) );
  XNOR2_X1 U15305 ( .A(n12234), .B(n12233), .ZN(n18945) );
  NAND2_X1 U15306 ( .A1(n18945), .A2(n12102), .ZN(n12243) );
  AND2_X1 U15307 ( .A1(n12243), .A2(n15388), .ZN(n15384) );
  NOR2_X1 U15308 ( .A1(n15383), .A2(n15384), .ZN(n15369) );
  AND2_X1 U15309 ( .A1(n12235), .A2(n15369), .ZN(n12247) );
  INV_X1 U15310 ( .A(n12236), .ZN(n12237) );
  NAND2_X1 U15311 ( .A1(n12102), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n12238) );
  OR2_X1 U15312 ( .A1(n18978), .A2(n12238), .ZN(n15365) );
  NAND2_X1 U15313 ( .A1(n12102), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n12239) );
  OR2_X1 U15314 ( .A1(n18999), .A2(n12239), .ZN(n15430) );
  OR2_X1 U15315 ( .A1(n12240), .A2(n21086), .ZN(n15444) );
  AND4_X1 U15316 ( .A1(n15365), .A2(n15364), .A3(n15430), .A4(n15444), .ZN(
        n12242) );
  OR2_X1 U15317 ( .A1(n12241), .A2(n15638), .ZN(n15428) );
  NAND3_X1 U15318 ( .A1(n15371), .A2(n12242), .A3(n15428), .ZN(n12245) );
  INV_X1 U15319 ( .A(n12243), .ZN(n12244) );
  OR3_X2 U15320 ( .A1(n18970), .A2(n12417), .A3(n15414), .ZN(n15407) );
  NAND2_X1 U15321 ( .A1(n15407), .A2(n15393), .ZN(n15367) );
  INV_X1 U15322 ( .A(n12248), .ZN(n12251) );
  INV_X1 U15323 ( .A(n12253), .ZN(n12249) );
  AOI21_X1 U15324 ( .B1(n12251), .B2(n12250), .A(n12249), .ZN(n15859) );
  AOI21_X1 U15325 ( .B1(n15859), .B2(n12102), .A(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15350) );
  NAND3_X1 U15326 ( .A1(n15859), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A3(
        n12102), .ZN(n15351) );
  NAND2_X1 U15327 ( .A1(n12253), .A2(n12252), .ZN(n12254) );
  NAND2_X1 U15328 ( .A1(n12256), .A2(n12254), .ZN(n13359) );
  OR2_X1 U15329 ( .A1(n13359), .A2(n12417), .ZN(n12255) );
  XNOR2_X1 U15330 ( .A(n12255), .B(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15341) );
  INV_X1 U15331 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15532) );
  NAND2_X1 U15332 ( .A1(n12412), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n12257) );
  MUX2_X1 U15333 ( .A(P2_EBX_REG_24__SCAN_IN), .B(n12257), .S(n12256), .Z(
        n12258) );
  NAND2_X1 U15334 ( .A1(n12258), .A2(n12269), .ZN(n15131) );
  NOR2_X1 U15335 ( .A1(n15131), .A2(n12417), .ZN(n15328) );
  INV_X1 U15336 ( .A(n15328), .ZN(n12259) );
  INV_X1 U15337 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15333) );
  NAND2_X1 U15338 ( .A1(n15330), .A2(n15333), .ZN(n12260) );
  AND2_X2 U15339 ( .A1(n12261), .A2(n12260), .ZN(n15308) );
  OR3_X1 U15340 ( .A1(n12263), .A2(n12262), .A3(n19286), .ZN(n12266) );
  INV_X1 U15341 ( .A(n12264), .ZN(n12265) );
  INV_X1 U15342 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15501) );
  NOR3_X1 U15343 ( .A1(n16211), .A2(n12417), .A3(n15501), .ZN(n12271) );
  INV_X1 U15344 ( .A(n16211), .ZN(n12267) );
  AOI21_X1 U15345 ( .B1(n12267), .B2(n12102), .A(
        P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n12268) );
  NAND2_X1 U15346 ( .A1(n12269), .A2(n12102), .ZN(n12270) );
  NAND2_X1 U15347 ( .A1(n12270), .A2(n15509), .ZN(n15319) );
  NOR2_X1 U15348 ( .A1(n12270), .A2(n15509), .ZN(n15318) );
  NOR2_X1 U15349 ( .A1(n12271), .A2(n15318), .ZN(n12408) );
  INV_X1 U15350 ( .A(n12272), .ZN(n12274) );
  NAND2_X1 U15351 ( .A1(n12274), .A2(n12273), .ZN(n12275) );
  NAND2_X1 U15352 ( .A1(n12280), .A2(n12275), .ZN(n13332) );
  INV_X1 U15353 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15300) );
  INV_X1 U15354 ( .A(n12277), .ZN(n12278) );
  OAI22_X1 U15355 ( .A1(n15298), .A2(n15300), .B1(n12278), .B2(n12403), .ZN(
        n12284) );
  AND2_X1 U15356 ( .A1(n12280), .A2(n12279), .ZN(n12281) );
  OR2_X1 U15357 ( .A1(n12281), .A2(n12411), .ZN(n15102) );
  INV_X1 U15358 ( .A(n15102), .ZN(n12282) );
  NAND2_X1 U15359 ( .A1(n12282), .A2(n12102), .ZN(n12404) );
  XNOR2_X1 U15360 ( .A(n12404), .B(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12283) );
  XNOR2_X1 U15361 ( .A(n12284), .B(n12283), .ZN(n15483) );
  OAI21_X1 U15362 ( .B1(n12286), .B2(n12299), .A(n12285), .ZN(n12287) );
  AOI21_X1 U15363 ( .B1(n12287), .B2(n12313), .A(n12318), .ZN(n19927) );
  INV_X1 U15364 ( .A(n16389), .ZN(n12288) );
  NOR2_X1 U15365 ( .A1(n12387), .A2(n12288), .ZN(n19930) );
  NAND2_X1 U15366 ( .A1(n19927), .A2(n19930), .ZN(n12397) );
  NOR2_X1 U15367 ( .A1(n12387), .A2(n12308), .ZN(n19929) );
  OAI21_X1 U15368 ( .B1(n12300), .B2(n12289), .A(n16373), .ZN(n12293) );
  INV_X1 U15369 ( .A(n12782), .ZN(n12292) );
  AOI21_X1 U15370 ( .B1(n12291), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n13539) );
  AOI21_X1 U15371 ( .B1(n12292), .B2(n13539), .A(P2_FLUSH_REG_SCAN_IN), .ZN(
        n19916) );
  MUX2_X1 U15372 ( .A(n12293), .B(n19916), .S(P2_STATE2_REG_1__SCAN_IN), .Z(
        n19928) );
  INV_X1 U15373 ( .A(n19928), .ZN(n12388) );
  NAND2_X1 U15374 ( .A1(n19929), .A2(n12388), .ZN(n12294) );
  NAND2_X1 U15375 ( .A1(n12397), .A2(n12294), .ZN(n12295) );
  NAND2_X1 U15376 ( .A1(n12295), .A2(n19808), .ZN(n18916) );
  OAI21_X1 U15377 ( .B1(n13335), .B2(n12297), .A(n12296), .ZN(n15472) );
  INV_X1 U15378 ( .A(n15472), .ZN(n15108) );
  AND2_X1 U15379 ( .A1(n19691), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19907) );
  INV_X1 U15380 ( .A(n12298), .ZN(n12299) );
  OAI21_X1 U15381 ( .B1(n12299), .B2(n12300), .A(n12114), .ZN(n12304) );
  NAND2_X1 U15382 ( .A1(n19271), .A2(n12300), .ZN(n12302) );
  NAND3_X1 U15383 ( .A1(n12302), .A2(n12392), .A3(n12301), .ZN(n12303) );
  OAI211_X1 U15384 ( .C1(n12306), .C2(n12305), .A(n12304), .B(n12303), .ZN(
        n12312) );
  NAND2_X1 U15385 ( .A1(n16370), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n19170) );
  NAND2_X1 U15386 ( .A1(n13427), .A2(n19170), .ZN(n12309) );
  MUX2_X1 U15387 ( .A(n12309), .B(n12308), .S(n12307), .Z(n12311) );
  INV_X1 U15388 ( .A(n12313), .ZN(n12310) );
  AOI21_X1 U15389 ( .B1(n12312), .B2(n12311), .A(n12310), .ZN(n12316) );
  NOR2_X1 U15390 ( .A1(n12114), .A2(n12313), .ZN(n12315) );
  OAI21_X1 U15391 ( .B1(n12316), .B2(n12315), .A(n12314), .ZN(n12317) );
  MUX2_X1 U15392 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B(n12317), .S(
        P2_STATE2_REG_0__SCAN_IN), .Z(n12393) );
  INV_X1 U15393 ( .A(n19170), .ZN(n12319) );
  AOI21_X1 U15394 ( .B1(n19735), .B2(n19802), .A(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n16399) );
  NAND2_X1 U15395 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n19915) );
  NOR2_X1 U15396 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n15767) );
  OR2_X1 U15397 ( .A1(n19691), .A2(n15767), .ZN(n19920) );
  NAND2_X1 U15398 ( .A1(n19920), .A2(n13537), .ZN(n12322) );
  NAND2_X1 U15399 ( .A1(n13537), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n12683) );
  NAND2_X1 U15400 ( .A1(n19573), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n12323) );
  NAND2_X1 U15401 ( .A1(n12683), .A2(n12323), .ZN(n15464) );
  NAND2_X1 U15402 ( .A1(n19038), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n15476) );
  NAND2_X1 U15403 ( .A1(n19246), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12324) );
  OAI211_X1 U15404 ( .C1(n19256), .C2(n12325), .A(n15476), .B(n12324), .ZN(
        n12326) );
  AOI21_X1 U15405 ( .B1(n15108), .B2(n19250), .A(n12326), .ZN(n12370) );
  XOR2_X1 U15406 ( .A(n12328), .B(n12327), .Z(n14524) );
  NAND2_X1 U15407 ( .A1(n12329), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n15466) );
  XNOR2_X1 U15408 ( .A(n12331), .B(n12330), .ZN(n12332) );
  NOR2_X1 U15409 ( .A1(n15466), .A2(n12332), .ZN(n12333) );
  XNOR2_X1 U15410 ( .A(n15466), .B(n12332), .ZN(n13553) );
  NOR2_X1 U15411 ( .A1(n15749), .A2(n13553), .ZN(n13552) );
  NOR2_X1 U15412 ( .A1(n12333), .A2(n13552), .ZN(n12334) );
  XNOR2_X1 U15413 ( .A(n21090), .B(n12334), .ZN(n14523) );
  NOR2_X1 U15414 ( .A1(n14524), .A2(n14523), .ZN(n14522) );
  NOR2_X1 U15415 ( .A1(n12334), .A2(n21090), .ZN(n12335) );
  OR2_X1 U15416 ( .A1(n14522), .A2(n12335), .ZN(n12336) );
  XNOR2_X1 U15417 ( .A(n12336), .B(n14095), .ZN(n14100) );
  NAND2_X1 U15418 ( .A1(n12336), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12337) );
  NAND2_X1 U15419 ( .A1(n12338), .A2(n12339), .ZN(n12340) );
  NAND2_X1 U15420 ( .A1(n12341), .A2(n12340), .ZN(n12343) );
  XNOR2_X1 U15421 ( .A(n12342), .B(n12343), .ZN(n14107) );
  NAND2_X1 U15422 ( .A1(n14107), .A2(n21161), .ZN(n12346) );
  INV_X1 U15423 ( .A(n12342), .ZN(n12344) );
  NAND2_X1 U15424 ( .A1(n12344), .A2(n12343), .ZN(n12345) );
  NAND2_X1 U15425 ( .A1(n12346), .A2(n12345), .ZN(n14217) );
  INV_X1 U15426 ( .A(n14217), .ZN(n12349) );
  NAND2_X1 U15427 ( .A1(n10249), .A2(n12358), .ZN(n12354) );
  INV_X1 U15428 ( .A(n14220), .ZN(n12352) );
  NAND2_X1 U15429 ( .A1(n12352), .A2(n12355), .ZN(n12353) );
  NAND2_X1 U15430 ( .A1(n14328), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12357) );
  XNOR2_X1 U15431 ( .A(n12363), .B(n12102), .ZN(n12361) );
  INV_X1 U15432 ( .A(n12361), .ZN(n12362) );
  NAND3_X1 U15433 ( .A1(n12366), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A3(
        n12102), .ZN(n12367) );
  AND2_X1 U15434 ( .A1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n12455) );
  NAND2_X1 U15435 ( .A1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n12466) );
  NAND2_X1 U15436 ( .A1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15616) );
  AND2_X1 U15437 ( .A1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n15636) );
  NAND2_X1 U15438 ( .A1(n15636), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n15434) );
  OR2_X1 U15439 ( .A1(n15616), .A2(n15434), .ZN(n15413) );
  NOR2_X1 U15440 ( .A1(n12466), .A2(n15413), .ZN(n15399) );
  AND2_X1 U15441 ( .A1(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n15399), .ZN(
        n12368) );
  AND2_X1 U15442 ( .A1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15521) );
  NAND2_X1 U15443 ( .A1(n15340), .A2(n15521), .ZN(n15331) );
  NAND2_X1 U15444 ( .A1(n15317), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15311) );
  XNOR2_X1 U15445 ( .A(n12372), .B(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n15471) );
  OR2_X1 U15446 ( .A1(n18916), .A2(n13427), .ZN(n16295) );
  NAND2_X1 U15447 ( .A1(n15471), .A2(n19251), .ZN(n12369) );
  INV_X1 U15448 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n12523) );
  INV_X1 U15449 ( .A(n12995), .ZN(n12401) );
  AND2_X1 U15450 ( .A1(n16365), .A2(n13427), .ZN(n13529) );
  NAND3_X1 U15451 ( .A1(n13529), .A2(n19275), .A3(n13530), .ZN(n12399) );
  NAND2_X1 U15452 ( .A1(n19271), .A2(n19281), .ZN(n12375) );
  NAND2_X1 U15453 ( .A1(n12375), .A2(n12392), .ZN(n12377) );
  AOI21_X1 U15454 ( .B1(n12377), .B2(n12376), .A(n19275), .ZN(n12378) );
  NOR2_X1 U15455 ( .A1(n12374), .A2(n12378), .ZN(n12385) );
  NAND2_X1 U15456 ( .A1(n12379), .A2(n12380), .ZN(n12381) );
  NAND2_X1 U15457 ( .A1(n13542), .A2(n12381), .ZN(n12384) );
  NAND3_X1 U15458 ( .A1(n16390), .A2(n16373), .A3(n13530), .ZN(n12383) );
  OAI21_X1 U15459 ( .B1(n12382), .B2(n11442), .A(n16389), .ZN(n12429) );
  NAND4_X1 U15460 ( .A1(n12385), .A2(n12384), .A3(n12383), .A4(n12429), .ZN(
        n13532) );
  INV_X1 U15461 ( .A(n19803), .ZN(n19812) );
  NOR2_X1 U15462 ( .A1(n12426), .A2(n19812), .ZN(n12386) );
  OAI211_X1 U15463 ( .C1(n16390), .C2(n19271), .A(n16373), .B(n12386), .ZN(
        n12390) );
  INV_X1 U15464 ( .A(n12387), .ZN(n16371) );
  NAND3_X1 U15465 ( .A1(n16371), .A2(n13427), .A3(n12388), .ZN(n12389) );
  NAND2_X1 U15466 ( .A1(n12390), .A2(n12389), .ZN(n12391) );
  NOR2_X1 U15467 ( .A1(n13532), .A2(n12391), .ZN(n12398) );
  INV_X1 U15468 ( .A(n13529), .ZN(n12395) );
  AOI21_X1 U15469 ( .B1(n12393), .B2(n12392), .A(n12432), .ZN(n12394) );
  NAND2_X1 U15470 ( .A1(n12395), .A2(n12394), .ZN(n12396) );
  NAND4_X1 U15471 ( .A1(n12399), .A2(n12398), .A3(n12397), .A4(n12396), .ZN(
        n12400) );
  NAND2_X1 U15472 ( .A1(n12401), .A2(n16342), .ZN(n12483) );
  AOI21_X1 U15473 ( .B1(n15473), .B2(n15300), .A(n12404), .ZN(n12406) );
  INV_X1 U15474 ( .A(n12404), .ZN(n12405) );
  OAI22_X1 U15475 ( .A1(n12407), .A2(n12406), .B1(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n12405), .ZN(n12409) );
  XNOR2_X1 U15476 ( .A(n12411), .B(n12410), .ZN(n12416) );
  OAI21_X1 U15477 ( .B1(n12416), .B2(n12417), .A(n12523), .ZN(n12493) );
  NAND2_X1 U15478 ( .A1(n12412), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n12413) );
  XNOR2_X1 U15479 ( .A(n12414), .B(n12413), .ZN(n13003) );
  AOI21_X1 U15480 ( .B1(n13003), .B2(n12102), .A(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n12502) );
  AND2_X1 U15481 ( .A1(n12102), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12415) );
  NAND2_X1 U15482 ( .A1(n13003), .A2(n12415), .ZN(n12503) );
  INV_X1 U15483 ( .A(n12416), .ZN(n15091) );
  NAND3_X1 U15484 ( .A1(n15091), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n12102), .ZN(n12500) );
  NOR2_X1 U15485 ( .A1(n12418), .A2(n12417), .ZN(n12419) );
  NAND2_X1 U15486 ( .A1(n12988), .A2(n16338), .ZN(n12482) );
  NAND2_X1 U15487 ( .A1(n12459), .A2(n12420), .ZN(n16326) );
  NAND2_X1 U15488 ( .A1(n12421), .A2(n12422), .ZN(n13531) );
  NAND2_X1 U15489 ( .A1(n11616), .A2(n13427), .ZN(n12423) );
  NAND2_X1 U15490 ( .A1(n13531), .A2(n12423), .ZN(n12424) );
  NAND2_X1 U15491 ( .A1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n14339) );
  OR2_X1 U15492 ( .A1(n12425), .A2(n14339), .ZN(n12456) );
  AND2_X1 U15493 ( .A1(n12426), .A2(n19286), .ZN(n12427) );
  AND2_X1 U15494 ( .A1(n12421), .A2(n12427), .ZN(n16366) );
  INV_X1 U15495 ( .A(n15610), .ZN(n12446) );
  OR2_X1 U15496 ( .A1(n12428), .A2(n19271), .ZN(n15735) );
  NAND2_X1 U15497 ( .A1(n15735), .A2(n12429), .ZN(n12441) );
  NAND2_X1 U15498 ( .A1(n12430), .A2(n12431), .ZN(n12438) );
  INV_X1 U15499 ( .A(n12431), .ZN(n12433) );
  NAND2_X1 U15500 ( .A1(n12433), .A2(n12432), .ZN(n12435) );
  INV_X1 U15501 ( .A(n12434), .ZN(n13426) );
  AOI22_X1 U15502 ( .A1(n12435), .A2(n13426), .B1(n19275), .B2(n16370), .ZN(
        n12436) );
  OAI211_X1 U15503 ( .C1(n12439), .C2(n12438), .A(n12437), .B(n12436), .ZN(
        n12440) );
  AOI21_X1 U15504 ( .B1(n12441), .B2(n14035), .A(n12440), .ZN(n12444) );
  NAND2_X1 U15505 ( .A1(n12442), .A2(n12443), .ZN(n12968) );
  NAND2_X1 U15506 ( .A1(n12444), .A2(n12968), .ZN(n15781) );
  OR2_X1 U15507 ( .A1(n15781), .A2(n13563), .ZN(n12445) );
  NAND2_X1 U15508 ( .A1(n12459), .A2(n12445), .ZN(n15612) );
  NAND2_X1 U15509 ( .A1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n14529) );
  NAND2_X1 U15510 ( .A1(n21090), .A2(n14529), .ZN(n14525) );
  INV_X1 U15511 ( .A(n14529), .ZN(n12457) );
  AOI22_X1 U15512 ( .A1(n15610), .A2(n14525), .B1(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n12457), .ZN(n14094) );
  NOR2_X1 U15513 ( .A1(n14094), .A2(n14095), .ZN(n14224) );
  NAND2_X1 U15514 ( .A1(n15613), .A2(n14224), .ZN(n14114) );
  NOR2_X1 U15515 ( .A1(n12456), .A2(n14114), .ZN(n16332) );
  NAND3_X1 U15516 ( .A1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A3(n16332), .ZN(n15713) );
  NOR2_X1 U15517 ( .A1(n15712), .A2(n15713), .ZN(n15687) );
  NAND2_X1 U15518 ( .A1(n12455), .A2(n15687), .ZN(n15666) );
  NOR2_X1 U15519 ( .A1(n15434), .A2(n15666), .ZN(n16316) );
  INV_X1 U15520 ( .A(n15616), .ZN(n12447) );
  AND2_X1 U15521 ( .A1(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n12447), .ZN(
        n12448) );
  NAND2_X1 U15522 ( .A1(n16316), .A2(n12448), .ZN(n15599) );
  NOR2_X1 U15523 ( .A1(n15401), .A2(n15388), .ZN(n12468) );
  NAND2_X1 U15524 ( .A1(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n12468), .ZN(
        n12449) );
  NAND2_X1 U15525 ( .A1(n15521), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n12450) );
  NOR2_X1 U15526 ( .A1(n15533), .A2(n12450), .ZN(n15510) );
  NOR2_X1 U15527 ( .A1(n15509), .A2(n15501), .ZN(n12474) );
  NOR2_X1 U15528 ( .A1(n15473), .A2(n15300), .ZN(n12476) );
  NAND2_X1 U15529 ( .A1(n15474), .A2(n12476), .ZN(n12524) );
  INV_X1 U15530 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n12528) );
  NOR4_X1 U15531 ( .A1(n12524), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n12523), .A4(n12528), .ZN(n12451) );
  NOR2_X1 U15532 ( .A1(n15684), .A2(n19874), .ZN(n12989) );
  NAND2_X1 U15533 ( .A1(n15613), .A2(n15434), .ZN(n12465) );
  INV_X1 U15534 ( .A(n12455), .ZN(n12464) );
  NAND2_X1 U15535 ( .A1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n16331) );
  INV_X1 U15536 ( .A(n14525), .ZN(n14093) );
  OR4_X1 U15537 ( .A1(n14095), .A2(n12456), .A3(n16331), .A4(n14093), .ZN(
        n12463) );
  NOR2_X1 U15538 ( .A1(n15612), .A2(n12457), .ZN(n12460) );
  INV_X1 U15539 ( .A(n12458), .ZN(n19245) );
  NOR2_X1 U15540 ( .A1(n12459), .A2(n19245), .ZN(n16339) );
  OR2_X1 U15541 ( .A1(n12460), .A2(n16339), .ZN(n14532) );
  INV_X1 U15542 ( .A(n14532), .ZN(n12462) );
  INV_X1 U15543 ( .A(n15612), .ZN(n12461) );
  NAND2_X1 U15544 ( .A1(n12461), .A2(n21090), .ZN(n14530) );
  NAND2_X1 U15545 ( .A1(n12462), .A2(n14530), .ZN(n14092) );
  AOI21_X1 U15546 ( .B1(n15613), .B2(n12463), .A(n14092), .ZN(n15711) );
  OAI21_X1 U15547 ( .B1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n16351), .A(
        n15711), .ZN(n15686) );
  AOI21_X1 U15548 ( .B1(n12464), .B2(n15613), .A(n15686), .ZN(n15665) );
  NAND2_X1 U15549 ( .A1(n16351), .A2(n16311), .ZN(n12471) );
  INV_X1 U15550 ( .A(n12471), .ZN(n12472) );
  OAI21_X1 U15551 ( .B1(n15616), .B2(n12466), .A(n15613), .ZN(n12467) );
  NAND2_X1 U15552 ( .A1(n16311), .A2(n12467), .ZN(n15607) );
  INV_X1 U15553 ( .A(n12468), .ZN(n15571) );
  NAND2_X1 U15554 ( .A1(n15613), .A2(n15571), .ZN(n12469) );
  NAND2_X1 U15555 ( .A1(n12469), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12470) );
  OR2_X1 U15556 ( .A1(n15607), .A2(n12470), .ZN(n15561) );
  NAND2_X1 U15557 ( .A1(n15561), .A2(n12471), .ZN(n15546) );
  OAI21_X1 U15558 ( .B1(n15521), .B2(n12472), .A(n15546), .ZN(n15528) );
  AND2_X1 U15559 ( .A1(n15613), .A2(n15333), .ZN(n12473) );
  NOR2_X1 U15560 ( .A1(n15528), .A2(n12473), .ZN(n15507) );
  INV_X1 U15561 ( .A(n12474), .ZN(n15498) );
  NAND2_X1 U15562 ( .A1(n15613), .A2(n15498), .ZN(n12475) );
  NAND2_X1 U15563 ( .A1(n15507), .A2(n12475), .ZN(n15492) );
  AOI21_X1 U15564 ( .B1(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n12476), .A(
        n16351), .ZN(n12477) );
  NOR2_X1 U15565 ( .A1(n15492), .A2(n12477), .ZN(n12529) );
  OAI21_X1 U15566 ( .B1(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n16351), .A(
        n12529), .ZN(n12478) );
  INV_X1 U15567 ( .A(n12478), .ZN(n12479) );
  NAND3_X1 U15568 ( .A1(n12483), .A2(n12482), .A3(n12481), .ZN(P2_U3015) );
  INV_X1 U15569 ( .A(n12506), .ZN(n12485) );
  OAI21_X1 U15570 ( .B1(n12372), .B2(n15473), .A(n12523), .ZN(n12484) );
  NAND2_X1 U15571 ( .A1(n12485), .A2(n12484), .ZN(n15297) );
  NAND2_X1 U15572 ( .A1(n12296), .A2(n12486), .ZN(n12487) );
  NAND2_X1 U15573 ( .A1(n12508), .A2(n12487), .ZN(n15293) );
  AOI21_X1 U15574 ( .B1(n12488), .B2(n15097), .A(n12516), .ZN(n15237) );
  NOR2_X1 U15575 ( .A1(n12524), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12489) );
  NOR2_X1 U15576 ( .A1(n15684), .A2(n19871), .ZN(n15291) );
  OAI21_X1 U15577 ( .B1(n15293), .B2(n16326), .A(n12491), .ZN(n12492) );
  NAND2_X1 U15578 ( .A1(n12500), .A2(n12493), .ZN(n12494) );
  XNOR2_X1 U15579 ( .A(n12495), .B(n12494), .ZN(n15295) );
  INV_X1 U15580 ( .A(n15492), .ZN(n12496) );
  NAND2_X1 U15581 ( .A1(n15474), .A2(n15300), .ZN(n15489) );
  NAND2_X1 U15582 ( .A1(n12496), .A2(n15489), .ZN(n15480) );
  AOI21_X1 U15583 ( .B1(n15474), .B2(n15473), .A(n15480), .ZN(n12497) );
  NAND2_X1 U15584 ( .A1(n12501), .A2(n12500), .ZN(n12505) );
  NAND2_X1 U15585 ( .A1(n9967), .A2(n12503), .ZN(n12504) );
  XNOR2_X1 U15586 ( .A(n12506), .B(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12534) );
  NOR2_X1 U15587 ( .A1(n15684), .A2(n12509), .ZN(n12522) );
  NOR2_X1 U15588 ( .A1(n19256), .A2(n12996), .ZN(n12510) );
  AOI211_X1 U15589 ( .C1(n19246), .C2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n12522), .B(n12510), .ZN(n12511) );
  OAI21_X1 U15590 ( .B1(n14470), .B2(n16305), .A(n12511), .ZN(n12512) );
  INV_X1 U15591 ( .A(n12512), .ZN(n12513) );
  NAND3_X1 U15592 ( .A1(n12515), .A2(n12514), .A3(n12513), .ZN(P2_U2984) );
  INV_X1 U15593 ( .A(n14470), .ZN(n12527) );
  INV_X1 U15594 ( .A(n12516), .ZN(n12519) );
  INV_X1 U15595 ( .A(n12517), .ZN(n12518) );
  NAND2_X1 U15596 ( .A1(n12519), .A2(n12518), .ZN(n12520) );
  NAND2_X1 U15597 ( .A1(n12521), .A2(n12520), .ZN(n13001) );
  INV_X1 U15598 ( .A(n12522), .ZN(n12525) );
  OAI211_X1 U15599 ( .C1(n13001), .C2(n16313), .A(n12525), .B(n9895), .ZN(
        n12526) );
  NAND2_X1 U15600 ( .A1(n12531), .A2(n16338), .ZN(n12532) );
  OAI211_X1 U15601 ( .C1(n12534), .C2(n16327), .A(n12533), .B(n12532), .ZN(
        P2_U3016) );
  AOI21_X1 U15602 ( .B1(n13781), .B2(n20157), .A(n10416), .ZN(n12562) );
  AND2_X1 U15603 ( .A1(n12562), .A2(n13959), .ZN(n13384) );
  INV_X1 U15604 ( .A(n13384), .ZN(n13715) );
  OAI21_X1 U15605 ( .B1(n20701), .B2(n13385), .A(n13715), .ZN(n12535) );
  NAND2_X1 U15606 ( .A1(n15901), .A2(n12535), .ZN(n12538) );
  INV_X1 U15607 ( .A(n12536), .ZN(n13899) );
  NOR3_X1 U15608 ( .A1(n13492), .A2(n20701), .A3(n13491), .ZN(n13370) );
  NAND2_X1 U15609 ( .A1(n13899), .A2(n13370), .ZN(n12537) );
  NAND2_X1 U15610 ( .A1(n12538), .A2(n12537), .ZN(n13734) );
  NAND4_X1 U15611 ( .A1(n20182), .A2(n20194), .A3(n13736), .A4(n10417), .ZN(
        n13807) );
  OR2_X1 U15612 ( .A1(n13709), .A2(n13807), .ZN(n12539) );
  AND2_X1 U15613 ( .A1(n20043), .A2(n20194), .ZN(n12541) );
  NOR4_X1 U15614 ( .A1(P1_ADDRESS_REG_16__SCAN_IN), .A2(
        P1_ADDRESS_REG_15__SCAN_IN), .A3(P1_ADDRESS_REG_14__SCAN_IN), .A4(
        P1_ADDRESS_REG_13__SCAN_IN), .ZN(n12545) );
  NOR4_X1 U15615 ( .A1(P1_ADDRESS_REG_20__SCAN_IN), .A2(
        P1_ADDRESS_REG_19__SCAN_IN), .A3(P1_ADDRESS_REG_18__SCAN_IN), .A4(
        P1_ADDRESS_REG_17__SCAN_IN), .ZN(n12544) );
  NOR4_X1 U15616 ( .A1(P1_ADDRESS_REG_7__SCAN_IN), .A2(
        P1_ADDRESS_REG_6__SCAN_IN), .A3(P1_ADDRESS_REG_5__SCAN_IN), .A4(
        P1_ADDRESS_REG_4__SCAN_IN), .ZN(n12543) );
  NOR4_X1 U15617 ( .A1(P1_ADDRESS_REG_12__SCAN_IN), .A2(
        P1_ADDRESS_REG_11__SCAN_IN), .A3(P1_ADDRESS_REG_9__SCAN_IN), .A4(
        P1_ADDRESS_REG_8__SCAN_IN), .ZN(n12542) );
  AND4_X1 U15618 ( .A1(n12545), .A2(n12544), .A3(n12543), .A4(n12542), .ZN(
        n12550) );
  NOR4_X1 U15619 ( .A1(P1_ADDRESS_REG_1__SCAN_IN), .A2(
        P1_ADDRESS_REG_0__SCAN_IN), .A3(P1_ADDRESS_REG_10__SCAN_IN), .A4(
        P1_ADDRESS_REG_3__SCAN_IN), .ZN(n12548) );
  NOR4_X1 U15620 ( .A1(P1_ADDRESS_REG_24__SCAN_IN), .A2(
        P1_ADDRESS_REG_23__SCAN_IN), .A3(P1_ADDRESS_REG_22__SCAN_IN), .A4(
        P1_ADDRESS_REG_21__SCAN_IN), .ZN(n12547) );
  NOR4_X1 U15621 ( .A1(P1_ADDRESS_REG_28__SCAN_IN), .A2(
        P1_ADDRESS_REG_27__SCAN_IN), .A3(P1_ADDRESS_REG_26__SCAN_IN), .A4(
        P1_ADDRESS_REG_25__SCAN_IN), .ZN(n12546) );
  INV_X1 U15622 ( .A(P1_ADDRESS_REG_2__SCAN_IN), .ZN(n20715) );
  AND4_X1 U15623 ( .A1(n12548), .A2(n12547), .A3(n12546), .A4(n20715), .ZN(
        n12549) );
  NAND2_X1 U15624 ( .A1(n12550), .A2(n12549), .ZN(n12551) );
  AND2_X2 U15625 ( .A1(n12551), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n20160)
         );
  AND2_X1 U15626 ( .A1(n13392), .A2(n20160), .ZN(n12552) );
  NAND2_X1 U15627 ( .A1(n20043), .A2(n12552), .ZN(n14802) );
  INV_X1 U15628 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n12553) );
  NOR2_X1 U15629 ( .A1(n14802), .A2(n12553), .ZN(n12557) );
  NOR3_X1 U15630 ( .A1(n14816), .A2(n20160), .A3(n13373), .ZN(n12554) );
  AOI22_X1 U15631 ( .A1(n14806), .A2(DATAI_31_), .B1(P1_EAX_REG_31__SCAN_IN), 
        .B2(n14816), .ZN(n12555) );
  INV_X1 U15632 ( .A(n12555), .ZN(n12556) );
  NAND2_X1 U15633 ( .A1(n10414), .A2(n20190), .ZN(n12561) );
  AND2_X1 U15634 ( .A1(n12561), .A2(n12560), .ZN(n13400) );
  NAND2_X1 U15635 ( .A1(n12563), .A2(n9858), .ZN(n12569) );
  NAND2_X1 U15636 ( .A1(n12570), .A2(n12564), .ZN(n12586) );
  OAI21_X1 U15637 ( .B1(n12564), .B2(n12570), .A(n12586), .ZN(n12565) );
  INV_X1 U15638 ( .A(n12565), .ZN(n12567) );
  AOI21_X1 U15639 ( .B1(n12567), .B2(n15891), .A(n12566), .ZN(n12568) );
  INV_X1 U15640 ( .A(n12630), .ZN(n12620) );
  INV_X1 U15641 ( .A(n12570), .ZN(n12572) );
  AND2_X1 U15642 ( .A1(n12571), .A2(n20157), .ZN(n12578) );
  AOI21_X1 U15643 ( .B1(n12572), .B2(n15891), .A(n12578), .ZN(n12573) );
  NAND2_X1 U15644 ( .A1(n13383), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13382) );
  INV_X1 U15645 ( .A(n12575), .ZN(n12576) );
  OR2_X1 U15646 ( .A1(n13382), .A2(n12576), .ZN(n12577) );
  OR2_X1 U15647 ( .A1(n13917), .A2(n12620), .ZN(n12581) );
  XNOR2_X1 U15648 ( .A(n12586), .B(n12585), .ZN(n12579) );
  AOI21_X1 U15649 ( .B1(n12579), .B2(n15891), .A(n12578), .ZN(n12580) );
  NAND2_X1 U15650 ( .A1(n12581), .A2(n12580), .ZN(n13778) );
  NAND2_X1 U15651 ( .A1(n13777), .A2(n13778), .ZN(n20126) );
  NAND2_X1 U15652 ( .A1(n12582), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12583) );
  INV_X1 U15653 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n12584) );
  NAND2_X1 U15654 ( .A1(n12586), .A2(n12585), .ZN(n12605) );
  INV_X1 U15655 ( .A(n12603), .ZN(n12587) );
  XNOR2_X1 U15656 ( .A(n12605), .B(n12587), .ZN(n12588) );
  NAND2_X1 U15657 ( .A1(n12588), .A2(n15891), .ZN(n12589) );
  NAND2_X1 U15658 ( .A1(n12590), .A2(n12589), .ZN(n13932) );
  NAND2_X1 U15659 ( .A1(n12591), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12592) );
  INV_X1 U15660 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n12593) );
  NAND2_X1 U15661 ( .A1(n12594), .A2(n12630), .ZN(n12598) );
  NAND2_X1 U15662 ( .A1(n12605), .A2(n12603), .ZN(n12595) );
  XNOR2_X1 U15663 ( .A(n12595), .B(n12602), .ZN(n12596) );
  NAND2_X1 U15664 ( .A1(n12596), .A2(n15891), .ZN(n12597) );
  NAND2_X1 U15665 ( .A1(n12598), .A2(n12597), .ZN(n20093) );
  NAND2_X1 U15666 ( .A1(n12601), .A2(n12630), .ZN(n12609) );
  AND2_X1 U15667 ( .A1(n12603), .A2(n12602), .ZN(n12604) );
  AND2_X1 U15668 ( .A1(n12605), .A2(n12604), .ZN(n12615) );
  INV_X1 U15669 ( .A(n12614), .ZN(n12606) );
  XNOR2_X1 U15670 ( .A(n12615), .B(n12606), .ZN(n12607) );
  NAND2_X1 U15671 ( .A1(n12607), .A2(n15891), .ZN(n12608) );
  NAND2_X1 U15672 ( .A1(n12609), .A2(n12608), .ZN(n12610) );
  INV_X1 U15673 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n16199) );
  XNOR2_X1 U15674 ( .A(n12610), .B(n16199), .ZN(n16099) );
  NAND2_X1 U15675 ( .A1(n12610), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12611) );
  NAND3_X1 U15676 ( .A1(n12612), .A2(n12630), .A3(n12613), .ZN(n12618) );
  NAND2_X1 U15677 ( .A1(n12615), .A2(n12614), .ZN(n12623) );
  XNOR2_X1 U15678 ( .A(n12622), .B(n12623), .ZN(n12616) );
  NAND2_X1 U15679 ( .A1(n15891), .A2(n12616), .ZN(n12617) );
  NAND2_X1 U15680 ( .A1(n12618), .A2(n12617), .ZN(n12619) );
  OR2_X1 U15681 ( .A1(n12619), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n14161) );
  NAND2_X1 U15682 ( .A1(n12619), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n14160) );
  OR2_X1 U15683 ( .A1(n12621), .A2(n12620), .ZN(n12628) );
  INV_X1 U15684 ( .A(n12622), .ZN(n12624) );
  NOR2_X1 U15685 ( .A1(n12624), .A2(n12623), .ZN(n12634) );
  INV_X1 U15686 ( .A(n12634), .ZN(n12625) );
  XNOR2_X1 U15687 ( .A(n12633), .B(n12625), .ZN(n12626) );
  NAND2_X1 U15688 ( .A1(n15891), .A2(n12626), .ZN(n12627) );
  NAND2_X1 U15689 ( .A1(n12628), .A2(n12627), .ZN(n12629) );
  NAND2_X1 U15690 ( .A1(n12629), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16090) );
  AND2_X1 U15691 ( .A1(n12631), .A2(n12630), .ZN(n12632) );
  AND3_X1 U15692 ( .A1(n15891), .A2(n12634), .A3(n12633), .ZN(n12635) );
  NAND2_X1 U15693 ( .A1(n14247), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12637) );
  AOI21_X1 U15694 ( .B1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A(n16081), .ZN(n14922) );
  NOR2_X1 U15695 ( .A1(n16081), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n14925) );
  NAND2_X1 U15696 ( .A1(n16081), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n16062) );
  OAI21_X1 U15697 ( .B1(n16081), .B2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n16062), .ZN(n14926) );
  OR2_X1 U15698 ( .A1(n16081), .A2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12639) );
  NAND2_X1 U15699 ( .A1(n16081), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n14911) );
  OAI21_X1 U15700 ( .B1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A(n16081), .ZN(n12640) );
  NOR2_X1 U15701 ( .A1(n16081), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15043) );
  XNOR2_X1 U15702 ( .A(n16081), .B(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15046) );
  NOR2_X1 U15703 ( .A1(n15043), .A2(n15046), .ZN(n12641) );
  NOR2_X1 U15704 ( .A1(n16081), .A2(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n12642) );
  NAND2_X1 U15705 ( .A1(n16081), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n14923) );
  INV_X1 U15706 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n12643) );
  NAND2_X1 U15707 ( .A1(n16080), .A2(n12643), .ZN(n12644) );
  NAND2_X1 U15708 ( .A1(n16081), .A2(n12644), .ZN(n14921) );
  OAI21_X1 U15709 ( .B1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A(n16081), .ZN(n12645) );
  XNOR2_X1 U15710 ( .A(n16081), .B(n16123), .ZN(n16050) );
  NAND2_X1 U15711 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n14492) );
  INV_X1 U15712 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n15025) );
  NOR2_X1 U15713 ( .A1(n14492), .A2(n15025), .ZN(n12647) );
  NAND2_X1 U15714 ( .A1(n15014), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n12650) );
  AND2_X1 U15715 ( .A1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n14495) );
  INV_X1 U15716 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15034) );
  NAND3_X1 U15717 ( .A1(n16109), .A2(n15034), .A3(n16123), .ZN(n12648) );
  NAND2_X1 U15718 ( .A1(n14873), .A2(n15025), .ZN(n12649) );
  INV_X1 U15719 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n14985) );
  NAND2_X1 U15720 ( .A1(n14999), .A2(n14985), .ZN(n14826) );
  OAI21_X2 U15721 ( .B1(n14856), .B2(n14826), .A(n16081), .ZN(n14848) );
  INV_X1 U15722 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14840) );
  NAND2_X1 U15723 ( .A1(n14840), .A2(n14831), .ZN(n14961) );
  AND2_X1 U15724 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n14963) );
  INV_X1 U15725 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n12653) );
  OR2_X1 U15726 ( .A1(n16081), .A2(n12653), .ZN(n14474) );
  NAND2_X1 U15727 ( .A1(n16081), .A2(n12653), .ZN(n14818) );
  NAND2_X1 U15728 ( .A1(n14474), .A2(n14818), .ZN(n12654) );
  XNOR2_X1 U15729 ( .A(n14476), .B(n12654), .ZN(n14959) );
  NAND2_X1 U15730 ( .A1(n20806), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n16202) );
  INV_X1 U15731 ( .A(n16202), .ZN(n12659) );
  NAND2_X1 U15732 ( .A1(n20802), .A2(n20413), .ZN(n20786) );
  NAND2_X1 U15733 ( .A1(n12660), .A2(n20786), .ZN(n20809) );
  AND2_X1 U15734 ( .A1(n20809), .A2(n20806), .ZN(n12661) );
  NAND2_X1 U15735 ( .A1(n20806), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n15889) );
  NAND2_X1 U15736 ( .A1(n20208), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n12662) );
  AND2_X1 U15737 ( .A1(n15889), .A2(n12662), .ZN(n13611) );
  INV_X1 U15738 ( .A(n13611), .ZN(n12663) );
  NAND2_X1 U15739 ( .A1(n20103), .A2(P1_REIP_REG_29__SCAN_IN), .ZN(n14953) );
  OAI21_X1 U15740 ( .B1(n14900), .B2(n12664), .A(n14953), .ZN(n12665) );
  AOI21_X1 U15741 ( .B1(n14513), .B2(n16077), .A(n12665), .ZN(n12666) );
  NAND2_X1 U15742 ( .A1(n19290), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12694) );
  AND2_X1 U15743 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19606) );
  NAND2_X1 U15744 ( .A1(n19898), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n19449) );
  INV_X1 U15745 ( .A(n19449), .ZN(n12667) );
  NAND2_X1 U15746 ( .A1(n19606), .A2(n12667), .ZN(n19481) );
  NAND2_X1 U15747 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19737) );
  INV_X1 U15748 ( .A(n19737), .ZN(n12668) );
  NAND2_X1 U15749 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n12668), .ZN(
        n19260) );
  NAND2_X1 U15750 ( .A1(n19260), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n12669) );
  NAND2_X1 U15751 ( .A1(n19481), .A2(n12669), .ZN(n12670) );
  AND2_X1 U15752 ( .A1(n12670), .A2(n19691), .ZN(n14032) );
  AOI21_X1 U15753 ( .B1(n12688), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n14032), .ZN(n12671) );
  AND2_X1 U15754 ( .A1(n12897), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n12692) );
  NAND2_X1 U15755 ( .A1(n12897), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n13623) );
  INV_X1 U15756 ( .A(n13623), .ZN(n13834) );
  INV_X1 U15757 ( .A(n12683), .ZN(n12676) );
  NAND2_X1 U15758 ( .A1(n12673), .A2(n12676), .ZN(n12675) );
  NAND2_X1 U15759 ( .A1(n19924), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19572) );
  NAND2_X1 U15760 ( .A1(n19914), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n19538) );
  NAND2_X1 U15761 ( .A1(n19572), .A2(n19538), .ZN(n19575) );
  AND2_X1 U15762 ( .A1(n19691), .A2(n19575), .ZN(n14129) );
  AOI21_X1 U15763 ( .B1(n12688), .B2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n14129), .ZN(n12674) );
  NAND2_X1 U15764 ( .A1(n12675), .A2(n12674), .ZN(n13581) );
  AOI22_X1 U15765 ( .A1(n12688), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n19691), .B2(n19924), .ZN(n12677) );
  INV_X1 U15766 ( .A(n12678), .ZN(n12681) );
  INV_X1 U15767 ( .A(n12679), .ZN(n12680) );
  NAND2_X1 U15768 ( .A1(n12681), .A2(n12680), .ZN(n12682) );
  NAND3_X1 U15769 ( .A1(n13838), .A2(n13834), .A3(n13622), .ZN(n12699) );
  NAND2_X1 U15770 ( .A1(n13625), .A2(n13623), .ZN(n12691) );
  INV_X1 U15771 ( .A(n19691), .ZN(n19886) );
  INV_X1 U15772 ( .A(n19606), .ZN(n12685) );
  NAND2_X1 U15773 ( .A1(n12685), .A2(n19905), .ZN(n12686) );
  NAND2_X1 U15774 ( .A1(n12686), .A2(n19260), .ZN(n14024) );
  NOR2_X1 U15775 ( .A1(n19886), .A2(n14024), .ZN(n12687) );
  AOI21_X1 U15776 ( .B1(n12688), .B2(n15752), .A(n12687), .ZN(n12689) );
  NAND3_X1 U15777 ( .A1(n13838), .A2(n12691), .A3(n13835), .ZN(n12698) );
  NAND2_X1 U15778 ( .A1(n12693), .A2(n12692), .ZN(n13839) );
  INV_X1 U15779 ( .A(n12694), .ZN(n12695) );
  NAND2_X1 U15780 ( .A1(n12695), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n12696) );
  NAND3_X1 U15781 ( .A1(n12699), .A2(n12698), .A3(n12697), .ZN(n13826) );
  AND2_X1 U15782 ( .A1(n12897), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n13827) );
  AND2_X1 U15783 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12700) );
  INV_X1 U15784 ( .A(n13882), .ZN(n12702) );
  AOI22_X1 U15785 ( .A1(n12781), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11772), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12709) );
  AOI22_X1 U15786 ( .A1(n11723), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11727), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12708) );
  AOI22_X1 U15787 ( .A1(n12782), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n11771), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12707) );
  AOI22_X1 U15788 ( .A1(n11770), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n12783), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12706) );
  NAND4_X1 U15789 ( .A1(n12709), .A2(n12708), .A3(n12707), .A4(n12706), .ZN(
        n12715) );
  AOI22_X1 U15790 ( .A1(n11778), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n11680), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12713) );
  AOI22_X1 U15791 ( .A1(n12788), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11777), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12712) );
  AOI22_X1 U15792 ( .A1(n11776), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n12789), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12711) );
  AOI22_X1 U15793 ( .A1(n11667), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11668), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12710) );
  NAND4_X1 U15794 ( .A1(n12713), .A2(n12712), .A3(n12711), .A4(n12710), .ZN(
        n12714) );
  NOR2_X1 U15795 ( .A1(n12715), .A2(n12714), .ZN(n14350) );
  AOI22_X1 U15796 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n12781), .B1(
        n11772), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12719) );
  AOI22_X1 U15797 ( .A1(n11723), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11727), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12718) );
  AOI22_X1 U15798 ( .A1(n12782), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n11771), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12717) );
  AOI22_X1 U15799 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n11770), .B1(
        n12783), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12716) );
  NAND4_X1 U15800 ( .A1(n12719), .A2(n12718), .A3(n12717), .A4(n12716), .ZN(
        n12725) );
  AOI22_X1 U15801 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n11778), .B1(
        n11680), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12723) );
  AOI22_X1 U15802 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n12788), .B1(
        n11777), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12722) );
  AOI22_X1 U15803 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n11776), .B1(
        n12789), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12721) );
  AOI22_X1 U15804 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n11667), .B1(
        n11668), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12720) );
  NAND4_X1 U15805 ( .A1(n12723), .A2(n12722), .A3(n12721), .A4(n12720), .ZN(
        n12724) );
  NOR2_X1 U15806 ( .A1(n12725), .A2(n12724), .ZN(n14384) );
  INV_X1 U15807 ( .A(n14384), .ZN(n12736) );
  AOI22_X1 U15808 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n12781), .B1(
        n11772), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12729) );
  AOI22_X1 U15809 ( .A1(n11723), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11727), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12728) );
  AOI22_X1 U15810 ( .A1(n12782), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n11771), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12727) );
  AOI22_X1 U15811 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n11770), .B1(
        n12783), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12726) );
  NAND4_X1 U15812 ( .A1(n12729), .A2(n12728), .A3(n12727), .A4(n12726), .ZN(
        n12735) );
  AOI22_X1 U15813 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n11778), .B1(
        n11680), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12733) );
  AOI22_X1 U15814 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n12788), .B1(
        n11777), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12732) );
  AOI22_X1 U15815 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n11776), .B1(
        n12789), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12731) );
  AOI22_X1 U15816 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n11667), .B1(
        n11668), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12730) );
  NAND4_X1 U15817 ( .A1(n12733), .A2(n12732), .A3(n12731), .A4(n12730), .ZN(
        n12734) );
  OR2_X1 U15818 ( .A1(n12735), .A2(n12734), .ZN(n14312) );
  AND2_X1 U15819 ( .A1(n12736), .A2(n14312), .ZN(n12737) );
  AOI22_X1 U15820 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n12781), .B1(
        n11772), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12741) );
  AOI22_X1 U15821 ( .A1(n11723), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11727), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12740) );
  AOI22_X1 U15822 ( .A1(n12782), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n11771), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12739) );
  AOI22_X1 U15823 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n11770), .B1(
        n12783), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12738) );
  NAND4_X1 U15824 ( .A1(n12741), .A2(n12740), .A3(n12739), .A4(n12738), .ZN(
        n12747) );
  AOI22_X1 U15825 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n11778), .B1(
        n11680), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12745) );
  AOI22_X1 U15826 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n11777), .B1(
        n12788), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12744) );
  AOI22_X1 U15827 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n11776), .B1(
        n12789), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12743) );
  AOI22_X1 U15828 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n11667), .B1(
        n11668), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12742) );
  NAND4_X1 U15829 ( .A1(n12745), .A2(n12744), .A3(n12743), .A4(n12742), .ZN(
        n12746) );
  NOR2_X1 U15830 ( .A1(n12747), .A2(n12746), .ZN(n15230) );
  AOI22_X1 U15831 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n12781), .B1(
        n11772), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12751) );
  AOI22_X1 U15832 ( .A1(n11723), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11727), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12750) );
  AOI22_X1 U15833 ( .A1(n12782), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n11771), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12749) );
  AOI22_X1 U15834 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n11770), .B1(
        n12783), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12748) );
  NAND4_X1 U15835 ( .A1(n12751), .A2(n12750), .A3(n12749), .A4(n12748), .ZN(
        n12757) );
  AOI22_X1 U15836 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n11778), .B1(
        n11680), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12755) );
  AOI22_X1 U15837 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n11777), .B1(
        n12788), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12754) );
  AOI22_X1 U15838 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n11776), .B1(
        n12789), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12753) );
  AOI22_X1 U15839 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n11667), .B1(
        n11668), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12752) );
  NAND4_X1 U15840 ( .A1(n12755), .A2(n12754), .A3(n12753), .A4(n12752), .ZN(
        n12756) );
  NOR2_X1 U15841 ( .A1(n12757), .A2(n12756), .ZN(n15206) );
  INV_X1 U15842 ( .A(n15206), .ZN(n12778) );
  AOI22_X1 U15843 ( .A1(n12781), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11772), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12761) );
  AOI22_X1 U15844 ( .A1(n11723), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11727), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12760) );
  AOI22_X1 U15845 ( .A1(n12782), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n11771), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12759) );
  AOI22_X1 U15846 ( .A1(n11770), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n12783), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12758) );
  NAND4_X1 U15847 ( .A1(n12761), .A2(n12760), .A3(n12759), .A4(n12758), .ZN(
        n12767) );
  AOI22_X1 U15848 ( .A1(n11778), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11680), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12765) );
  AOI22_X1 U15849 ( .A1(n12788), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11777), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12764) );
  AOI22_X1 U15850 ( .A1(n11776), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n12789), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12763) );
  AOI22_X1 U15851 ( .A1(n11667), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11668), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12762) );
  NAND4_X1 U15852 ( .A1(n12765), .A2(n12764), .A3(n12763), .A4(n12762), .ZN(
        n12766) );
  OR2_X1 U15853 ( .A1(n12767), .A2(n12766), .ZN(n15211) );
  AOI22_X1 U15854 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n12781), .B1(
        n11772), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12771) );
  AOI22_X1 U15855 ( .A1(n11723), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n11727), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12770) );
  AOI22_X1 U15856 ( .A1(n12782), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n11771), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12769) );
  AOI22_X1 U15857 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n11770), .B1(
        n12783), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12768) );
  NAND4_X1 U15858 ( .A1(n12771), .A2(n12770), .A3(n12769), .A4(n12768), .ZN(
        n12777) );
  AOI22_X1 U15859 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n11778), .B1(
        n11680), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12775) );
  AOI22_X1 U15860 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n11777), .B1(
        n12788), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12774) );
  AOI22_X1 U15861 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n11776), .B1(
        n12789), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12773) );
  AOI22_X1 U15862 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n11667), .B1(
        n11668), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12772) );
  NAND4_X1 U15863 ( .A1(n12775), .A2(n12774), .A3(n12773), .A4(n12772), .ZN(
        n12776) );
  OR2_X1 U15864 ( .A1(n12777), .A2(n12776), .ZN(n15220) );
  AND2_X1 U15865 ( .A1(n15211), .A2(n15220), .ZN(n15204) );
  NAND2_X1 U15866 ( .A1(n12778), .A2(n15204), .ZN(n12779) );
  NOR2_X1 U15867 ( .A1(n15230), .A2(n12779), .ZN(n12780) );
  AOI22_X1 U15868 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n12781), .B1(
        n11772), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12787) );
  AOI22_X1 U15869 ( .A1(n11723), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11727), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12786) );
  AOI22_X1 U15870 ( .A1(n12782), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n11771), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12785) );
  AOI22_X1 U15871 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n11770), .B1(
        n12783), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12784) );
  NAND4_X1 U15872 ( .A1(n12787), .A2(n12786), .A3(n12785), .A4(n12784), .ZN(
        n12796) );
  AOI22_X1 U15873 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n11778), .B1(
        n11680), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12794) );
  AOI22_X1 U15874 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n11777), .B1(
        n12788), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12793) );
  AOI22_X1 U15875 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n11776), .B1(
        n12789), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12792) );
  AOI22_X1 U15876 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n11667), .B1(
        n11668), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12791) );
  NAND4_X1 U15877 ( .A1(n12794), .A2(n12793), .A3(n12792), .A4(n12791), .ZN(
        n12795) );
  NOR2_X1 U15878 ( .A1(n12796), .A2(n12795), .ZN(n12835) );
  AOI22_X1 U15879 ( .A1(n12944), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n12941), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12807) );
  AOI22_X1 U15880 ( .A1(n12954), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12798), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12806) );
  AOI22_X1 U15881 ( .A1(n12953), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n9852), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12805) );
  NAND2_X1 U15882 ( .A1(n12955), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n12803) );
  AND2_X1 U15883 ( .A1(n15752), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12800) );
  OR2_X1 U15884 ( .A1(n12800), .A2(n12799), .ZN(n12956) );
  NAND2_X1 U15885 ( .A1(n11652), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n12802) );
  AND3_X1 U15886 ( .A1(n12803), .A2(n12956), .A3(n12802), .ZN(n12804) );
  NAND4_X1 U15887 ( .A1(n12807), .A2(n12806), .A3(n12805), .A4(n12804), .ZN(
        n12815) );
  AOI22_X1 U15888 ( .A1(n12954), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n9856), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12813) );
  INV_X1 U15889 ( .A(n12956), .ZN(n12922) );
  NAND2_X1 U15890 ( .A1(n12945), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n12809) );
  NAND2_X1 U15891 ( .A1(n12953), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n12808) );
  AND3_X1 U15892 ( .A1(n12922), .A2(n12809), .A3(n12808), .ZN(n12812) );
  AOI22_X1 U15893 ( .A1(n12944), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n9830), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12811) );
  AOI22_X1 U15894 ( .A1(n12941), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11652), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12810) );
  NAND4_X1 U15895 ( .A1(n12813), .A2(n12812), .A3(n12811), .A4(n12810), .ZN(
        n12814) );
  NAND2_X1 U15896 ( .A1(n12815), .A2(n12814), .ZN(n12840) );
  NOR2_X1 U15897 ( .A1(n19271), .A2(n12840), .ZN(n12816) );
  XOR2_X1 U15898 ( .A(n12835), .B(n12816), .Z(n12841) );
  INV_X1 U15899 ( .A(n12840), .ZN(n12836) );
  NAND2_X1 U15900 ( .A1(n12058), .A2(n12836), .ZN(n15197) );
  INV_X1 U15901 ( .A(n12817), .ZN(n15205) );
  INV_X1 U15902 ( .A(n12841), .ZN(n12818) );
  AOI22_X1 U15903 ( .A1(n12954), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12941), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12825) );
  NAND2_X1 U15904 ( .A1(n12945), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n12821) );
  NAND2_X1 U15905 ( .A1(n12953), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n12820) );
  AND3_X1 U15906 ( .A1(n12922), .A2(n12821), .A3(n12820), .ZN(n12824) );
  AOI22_X1 U15907 ( .A1(n12944), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12950), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12823) );
  AOI22_X1 U15908 ( .A1(n12929), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11652), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12822) );
  NAND4_X1 U15909 ( .A1(n12825), .A2(n12824), .A3(n12823), .A4(n12822), .ZN(
        n12834) );
  INV_X1 U15910 ( .A(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n21142) );
  AOI22_X1 U15911 ( .A1(n12954), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12941), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12832) );
  NAND2_X1 U15912 ( .A1(n12955), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n12827) );
  INV_X1 U15913 ( .A(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n19335) );
  NAND2_X1 U15914 ( .A1(n12953), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n12826) );
  AND3_X1 U15915 ( .A1(n12827), .A2(n12956), .A3(n12826), .ZN(n12831) );
  AOI22_X1 U15916 ( .A1(n12944), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n12950), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12830) );
  AOI22_X1 U15917 ( .A1(n9857), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n11652), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12829) );
  NAND4_X1 U15918 ( .A1(n12832), .A2(n12831), .A3(n12830), .A4(n12829), .ZN(
        n12833) );
  AND2_X1 U15919 ( .A1(n12834), .A2(n12833), .ZN(n12839) );
  INV_X1 U15920 ( .A(n12835), .ZN(n12837) );
  AND2_X1 U15921 ( .A1(n12837), .A2(n12836), .ZN(n12838) );
  NAND2_X1 U15922 ( .A1(n12838), .A2(n12839), .ZN(n12842) );
  OAI211_X1 U15923 ( .C1(n12839), .C2(n12838), .A(n12897), .B(n12842), .ZN(
        n15189) );
  NAND2_X1 U15924 ( .A1(n19271), .A2(n12839), .ZN(n15191) );
  INV_X1 U15925 ( .A(n12842), .ZN(n12857) );
  AOI22_X1 U15926 ( .A1(n12954), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12941), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12848) );
  NAND2_X1 U15927 ( .A1(n12945), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n12844) );
  NAND2_X1 U15928 ( .A1(n12953), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n12843) );
  AND3_X1 U15929 ( .A1(n12922), .A2(n12844), .A3(n12843), .ZN(n12847) );
  AOI22_X1 U15930 ( .A1(n12944), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12950), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12846) );
  AOI22_X1 U15931 ( .A1(n9856), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11652), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12845) );
  NAND4_X1 U15932 ( .A1(n12848), .A2(n12847), .A3(n12846), .A4(n12845), .ZN(
        n12856) );
  AOI22_X1 U15933 ( .A1(n12798), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n12941), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12854) );
  NAND2_X1 U15934 ( .A1(n12955), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n12850) );
  INV_X1 U15935 ( .A(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n21044) );
  NAND2_X1 U15936 ( .A1(n12953), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n12849) );
  AND3_X1 U15937 ( .A1(n12850), .A2(n12956), .A3(n12849), .ZN(n12853) );
  AOI22_X1 U15938 ( .A1(n12954), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12950), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12852) );
  AOI22_X1 U15939 ( .A1(n12944), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n11652), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12851) );
  NAND4_X1 U15940 ( .A1(n12854), .A2(n12853), .A3(n12852), .A4(n12851), .ZN(
        n12855) );
  AND2_X1 U15941 ( .A1(n12856), .A2(n12855), .ZN(n12859) );
  NAND2_X1 U15942 ( .A1(n12857), .A2(n12859), .ZN(n12877) );
  OAI211_X1 U15943 ( .C1(n12857), .C2(n12859), .A(n12897), .B(n12877), .ZN(
        n12861) );
  INV_X1 U15944 ( .A(n12859), .ZN(n12860) );
  NOR2_X1 U15945 ( .A1(n13427), .A2(n12860), .ZN(n15185) );
  NAND2_X1 U15946 ( .A1(n12955), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(
        n12864) );
  NAND2_X1 U15947 ( .A1(n12953), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n12863) );
  AND3_X1 U15948 ( .A1(n12922), .A2(n12864), .A3(n12863), .ZN(n12868) );
  AOI22_X1 U15949 ( .A1(n12954), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12941), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12867) );
  AOI22_X1 U15950 ( .A1(n12944), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12950), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12866) );
  AOI22_X1 U15951 ( .A1(n12929), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11652), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12865) );
  NAND4_X1 U15952 ( .A1(n12868), .A2(n12867), .A3(n12866), .A4(n12865), .ZN(
        n12876) );
  AOI22_X1 U15953 ( .A1(n12954), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12941), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12874) );
  NAND2_X1 U15954 ( .A1(n12955), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n12870) );
  NAND2_X1 U15955 ( .A1(n12953), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n12869) );
  AND3_X1 U15956 ( .A1(n12870), .A2(n12956), .A3(n12869), .ZN(n12873) );
  AOI22_X1 U15957 ( .A1(n12944), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n12950), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12872) );
  AOI22_X1 U15958 ( .A1(n9857), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n11652), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12871) );
  NAND4_X1 U15959 ( .A1(n12874), .A2(n12873), .A3(n12872), .A4(n12871), .ZN(
        n12875) );
  NAND2_X1 U15960 ( .A1(n12876), .A2(n12875), .ZN(n12879) );
  OR2_X1 U15961 ( .A1(n12877), .A2(n12879), .ZN(n12896) );
  NAND2_X1 U15962 ( .A1(n12877), .A2(n12879), .ZN(n12878) );
  INV_X1 U15963 ( .A(n12879), .ZN(n12880) );
  NAND2_X1 U15964 ( .A1(n19271), .A2(n12880), .ZN(n15178) );
  NAND2_X1 U15965 ( .A1(n12955), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n12883) );
  NAND2_X1 U15966 ( .A1(n12953), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n12882) );
  AND3_X1 U15967 ( .A1(n12922), .A2(n12883), .A3(n12882), .ZN(n12887) );
  AOI22_X1 U15968 ( .A1(n12954), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n12941), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12886) );
  AOI22_X1 U15969 ( .A1(n12944), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n12950), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12885) );
  AOI22_X1 U15970 ( .A1(n9856), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11652), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12884) );
  NAND4_X1 U15971 ( .A1(n12887), .A2(n12886), .A3(n12885), .A4(n12884), .ZN(
        n12895) );
  AOI22_X1 U15972 ( .A1(n12954), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n12941), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12893) );
  NAND2_X1 U15973 ( .A1(n12955), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n12889) );
  NAND2_X1 U15974 ( .A1(n12953), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n12888) );
  AND3_X1 U15975 ( .A1(n12889), .A2(n12956), .A3(n12888), .ZN(n12892) );
  AOI22_X1 U15976 ( .A1(n12944), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n12950), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12891) );
  AOI22_X1 U15977 ( .A1(n12798), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n11652), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12890) );
  NAND4_X1 U15978 ( .A1(n12893), .A2(n12892), .A3(n12891), .A4(n12890), .ZN(
        n12894) );
  NAND2_X1 U15979 ( .A1(n12895), .A2(n12894), .ZN(n12903) );
  INV_X1 U15980 ( .A(n12903), .ZN(n12899) );
  INV_X1 U15981 ( .A(n12896), .ZN(n12898) );
  OR2_X1 U15982 ( .A1(n12896), .A2(n12903), .ZN(n12936) );
  OAI211_X1 U15983 ( .C1(n12899), .C2(n12898), .A(n12936), .B(n12897), .ZN(
        n12900) );
  NOR2_X1 U15984 ( .A1(n13427), .A2(n12903), .ZN(n15171) );
  INV_X1 U15985 ( .A(n12904), .ZN(n12919) );
  NAND2_X1 U15986 ( .A1(n12955), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n12906) );
  NAND2_X1 U15987 ( .A1(n12953), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n12905) );
  AND3_X1 U15988 ( .A1(n12922), .A2(n12906), .A3(n12905), .ZN(n12910) );
  AOI22_X1 U15989 ( .A1(n12954), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12941), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12909) );
  AOI22_X1 U15990 ( .A1(n12944), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12950), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12908) );
  AOI22_X1 U15991 ( .A1(n9857), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11652), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12907) );
  NAND4_X1 U15992 ( .A1(n12910), .A2(n12909), .A3(n12908), .A4(n12907), .ZN(
        n12918) );
  AOI22_X1 U15993 ( .A1(n12954), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12941), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12916) );
  NAND2_X1 U15994 ( .A1(n12955), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n12912) );
  NAND2_X1 U15995 ( .A1(n12953), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n12911) );
  AND3_X1 U15996 ( .A1(n12912), .A2(n12956), .A3(n12911), .ZN(n12915) );
  AOI22_X1 U15997 ( .A1(n12944), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n12950), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12914) );
  AOI22_X1 U15998 ( .A1(n12929), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11652), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12913) );
  NAND4_X1 U15999 ( .A1(n12916), .A2(n12915), .A3(n12914), .A4(n12913), .ZN(
        n12917) );
  NAND2_X1 U16000 ( .A1(n12918), .A2(n12917), .ZN(n15166) );
  AOI22_X1 U16001 ( .A1(n12929), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12941), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12926) );
  NAND2_X1 U16002 ( .A1(n12955), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n12921) );
  NAND2_X1 U16003 ( .A1(n11652), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n12920) );
  AND3_X1 U16004 ( .A1(n12922), .A2(n12921), .A3(n12920), .ZN(n12925) );
  AOI22_X1 U16005 ( .A1(n12944), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12950), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12924) );
  AOI22_X1 U16006 ( .A1(n12954), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12953), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12923) );
  NAND4_X1 U16007 ( .A1(n12926), .A2(n12925), .A3(n12924), .A4(n12923), .ZN(
        n12935) );
  AOI22_X1 U16008 ( .A1(n12944), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n12941), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12933) );
  NAND2_X1 U16009 ( .A1(n12955), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n12928) );
  NAND2_X1 U16010 ( .A1(n11652), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(
        n12927) );
  AND3_X1 U16011 ( .A1(n12928), .A2(n12956), .A3(n12927), .ZN(n12932) );
  AOI22_X1 U16012 ( .A1(n12954), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12950), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12931) );
  AOI22_X1 U16013 ( .A1(n12929), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n12953), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12930) );
  NAND4_X1 U16014 ( .A1(n12933), .A2(n12932), .A3(n12931), .A4(n12930), .ZN(
        n12934) );
  NAND2_X1 U16015 ( .A1(n12935), .A2(n12934), .ZN(n12939) );
  INV_X1 U16016 ( .A(n12936), .ZN(n15165) );
  NOR2_X1 U16017 ( .A1(n12058), .A2(n15166), .ZN(n12937) );
  NAND2_X1 U16018 ( .A1(n15165), .A2(n12937), .ZN(n12938) );
  NOR2_X1 U16019 ( .A1(n12938), .A2(n12939), .ZN(n12940) );
  AOI21_X1 U16020 ( .B1(n12939), .B2(n12938), .A(n12940), .ZN(n15160) );
  NOR2_X1 U16021 ( .A1(n15159), .A2(n12940), .ZN(n12965) );
  AOI22_X1 U16022 ( .A1(n12929), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12941), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12943) );
  AOI22_X1 U16023 ( .A1(n12797), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12950), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12942) );
  NAND2_X1 U16024 ( .A1(n12943), .A2(n12942), .ZN(n12963) );
  AOI22_X1 U16025 ( .A1(n12944), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12953), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12947) );
  AOI21_X1 U16026 ( .B1(n12945), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A(
        n12956), .ZN(n12946) );
  OAI211_X1 U16027 ( .C1(n12801), .C2(n12948), .A(n12947), .B(n12946), .ZN(
        n12962) );
  AOI22_X1 U16028 ( .A1(n12944), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n12941), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12952) );
  AOI22_X1 U16029 ( .A1(n12798), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n12950), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12951) );
  NAND2_X1 U16030 ( .A1(n12952), .A2(n12951), .ZN(n12961) );
  AOI22_X1 U16031 ( .A1(n12797), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12953), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12959) );
  NAND2_X1 U16032 ( .A1(n12955), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n12958) );
  NAND2_X1 U16033 ( .A1(n11652), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n12957) );
  NAND4_X1 U16034 ( .A1(n12959), .A2(n12958), .A3(n12957), .A4(n12956), .ZN(
        n12960) );
  OAI22_X1 U16035 ( .A1(n12963), .A2(n12962), .B1(n12961), .B2(n12960), .ZN(
        n12964) );
  XNOR2_X1 U16036 ( .A(n12965), .B(n12964), .ZN(n14473) );
  NAND2_X1 U16037 ( .A1(n12434), .A2(n19803), .ZN(n16374) );
  INV_X1 U16038 ( .A(n16373), .ZN(n16363) );
  NOR2_X1 U16039 ( .A1(n16374), .A2(n16363), .ZN(n12966) );
  AND2_X1 U16040 ( .A1(n11616), .A2(n12966), .ZN(n12967) );
  AOI21_X1 U16041 ( .B1(n16365), .B2(n16366), .A(n12967), .ZN(n13534) );
  NAND2_X1 U16042 ( .A1(n13534), .A2(n12968), .ZN(n12969) );
  NAND2_X1 U16043 ( .A1(n19140), .A2(n10156), .ZN(n15285) );
  AND2_X1 U16044 ( .A1(n19140), .A2(n12970), .ZN(n19108) );
  NOR4_X1 U16045 ( .A1(P2_ADDRESS_REG_14__SCAN_IN), .A2(
        P2_ADDRESS_REG_13__SCAN_IN), .A3(P2_ADDRESS_REG_12__SCAN_IN), .A4(
        P2_ADDRESS_REG_11__SCAN_IN), .ZN(n12974) );
  NOR4_X1 U16046 ( .A1(P2_ADDRESS_REG_18__SCAN_IN), .A2(
        P2_ADDRESS_REG_17__SCAN_IN), .A3(P2_ADDRESS_REG_16__SCAN_IN), .A4(
        P2_ADDRESS_REG_15__SCAN_IN), .ZN(n12973) );
  NOR4_X1 U16047 ( .A1(P2_ADDRESS_REG_6__SCAN_IN), .A2(
        P2_ADDRESS_REG_5__SCAN_IN), .A3(P2_ADDRESS_REG_4__SCAN_IN), .A4(
        P2_ADDRESS_REG_3__SCAN_IN), .ZN(n12972) );
  NOR4_X1 U16048 ( .A1(P2_ADDRESS_REG_10__SCAN_IN), .A2(
        P2_ADDRESS_REG_9__SCAN_IN), .A3(P2_ADDRESS_REG_8__SCAN_IN), .A4(
        P2_ADDRESS_REG_7__SCAN_IN), .ZN(n12971) );
  NAND4_X1 U16049 ( .A1(n12974), .A2(n12973), .A3(n12972), .A4(n12971), .ZN(
        n12979) );
  NOR4_X1 U16050 ( .A1(P2_ADDRESS_REG_1__SCAN_IN), .A2(
        P2_ADDRESS_REG_0__SCAN_IN), .A3(P2_ADDRESS_REG_28__SCAN_IN), .A4(
        P2_ADDRESS_REG_27__SCAN_IN), .ZN(n12977) );
  NOR4_X1 U16051 ( .A1(P2_ADDRESS_REG_22__SCAN_IN), .A2(
        P2_ADDRESS_REG_21__SCAN_IN), .A3(P2_ADDRESS_REG_20__SCAN_IN), .A4(
        P2_ADDRESS_REG_19__SCAN_IN), .ZN(n12976) );
  NOR4_X1 U16052 ( .A1(P2_ADDRESS_REG_26__SCAN_IN), .A2(
        P2_ADDRESS_REG_25__SCAN_IN), .A3(P2_ADDRESS_REG_24__SCAN_IN), .A4(
        P2_ADDRESS_REG_23__SCAN_IN), .ZN(n12975) );
  INV_X1 U16053 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n19834) );
  NAND4_X1 U16054 ( .A1(n12977), .A2(n12976), .A3(n12975), .A4(n19834), .ZN(
        n12978) );
  OAI21_X1 U16055 ( .B1(n12979), .B2(n12978), .A(P2_ADDRESS_REG_29__SCAN_IN), 
        .ZN(n12980) );
  NAND2_X1 U16056 ( .A1(n14029), .A2(BUF2_REG_14__SCAN_IN), .ZN(n12982) );
  INV_X1 U16057 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n14371) );
  OR2_X1 U16058 ( .A1(n14029), .A2(n14371), .ZN(n12981) );
  NAND2_X1 U16059 ( .A1(n12982), .A2(n12981), .ZN(n19238) );
  AOI22_X1 U16060 ( .A1(n19108), .A2(n19238), .B1(n19155), .B2(
        P2_EAX_REG_30__SCAN_IN), .ZN(n12983) );
  OAI21_X1 U16061 ( .B1(n13001), .B2(n15285), .A(n12983), .ZN(n12984) );
  INV_X1 U16062 ( .A(n12984), .ZN(n12987) );
  AND2_X1 U16063 ( .A1(n19140), .A2(n12985), .ZN(n13574) );
  AOI22_X1 U16064 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n19110), .B1(n19109), .B2(
        BUF2_REG_30__SCAN_IN), .ZN(n12986) );
  OAI21_X1 U16065 ( .B1(n14473), .B2(n19160), .A(n10266), .ZN(P2_U2889) );
  NAND2_X1 U16066 ( .A1(n12988), .A2(n19248), .ZN(n12994) );
  AOI21_X1 U16067 ( .B1(n19246), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n12989), .ZN(n12990) );
  OAI21_X1 U16068 ( .B1(n19256), .B2(n12991), .A(n12990), .ZN(n12992) );
  OAI211_X1 U16069 ( .C1(n12995), .C2(n16295), .A(n12994), .B(n12993), .ZN(
        P2_U2983) );
  NOR2_X1 U16070 ( .A1(n10053), .A2(n15084), .ZN(n12997) );
  XNOR2_X1 U16071 ( .A(n12997), .B(n12996), .ZN(n12998) );
  NAND2_X1 U16072 ( .A1(n12998), .A2(n9868), .ZN(n13007) );
  AOI22_X1 U16073 ( .A1(n19091), .A2(P2_REIP_REG_30__SCAN_IN), .B1(n19090), 
        .B2(P2_EBX_REG_30__SCAN_IN), .ZN(n13000) );
  NAND2_X1 U16074 ( .A1(n19101), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12999) );
  OAI211_X1 U16075 ( .C1(n13001), .C2(n19087), .A(n13000), .B(n12999), .ZN(
        n13002) );
  AOI21_X1 U16076 ( .B1(n13003), .B2(n19049), .A(n13002), .ZN(n13005) );
  AND2_X1 U16077 ( .A1(n13005), .A2(n13004), .ZN(n13006) );
  NAND2_X1 U16078 ( .A1(n13007), .A2(n13006), .ZN(P2_U2825) );
  AOI22_X1 U16079 ( .A1(n17211), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n9839), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n13025) );
  AOI22_X1 U16080 ( .A1(n9849), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(n9838), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n13024) );
  INV_X1 U16081 ( .A(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n21192) );
  AOI22_X1 U16082 ( .A1(n17112), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n17213), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n13008) );
  OAI21_X1 U16083 ( .B1(n13161), .B2(n21192), .A(n13008), .ZN(n13022) );
  AOI22_X1 U16084 ( .A1(n9832), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(n9837), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n13020) );
  NOR2_X1 U16085 ( .A1(n13014), .A2(n13010), .ZN(n13011) );
  AOI22_X1 U16086 ( .A1(n17199), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n17194), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n13019) );
  NOR2_X2 U16087 ( .A1(n16947), .A2(n13012), .ZN(n13013) );
  NOR2_X1 U16088 ( .A1(n16947), .A2(n13014), .ZN(n13063) );
  AOI22_X1 U16089 ( .A1(n17193), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n17216), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n13018) );
  INV_X2 U16090 ( .A(n10259), .ZN(n17153) );
  INV_X2 U16091 ( .A(n17215), .ZN(n15785) );
  AOI22_X1 U16092 ( .A1(n17153), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n15785), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n13017) );
  NAND4_X1 U16093 ( .A1(n13020), .A2(n13019), .A3(n13018), .A4(n13017), .ZN(
        n13021) );
  AOI211_X1 U16094 ( .C1(n17219), .C2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A(
        n13022), .B(n13021), .ZN(n13023) );
  NAND3_X1 U16095 ( .A1(n13025), .A2(n13024), .A3(n13023), .ZN(n13304) );
  AOI22_X1 U16096 ( .A1(n9832), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(n9839), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n13036) );
  AOI22_X1 U16097 ( .A1(n17220), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n9837), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n13035) );
  INV_X1 U16098 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n17246) );
  AOI22_X1 U16099 ( .A1(n17112), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17213), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n13026) );
  OAI21_X1 U16100 ( .B1(n9887), .B2(n17246), .A(n13026), .ZN(n13033) );
  CLKBUF_X3 U16101 ( .A(n13065), .Z(n17211) );
  AOI22_X1 U16102 ( .A1(n17153), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17211), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n13031) );
  INV_X2 U16103 ( .A(n17136), .ZN(n17194) );
  AOI22_X1 U16104 ( .A1(n17194), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17216), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n13030) );
  INV_X2 U16105 ( .A(n17215), .ZN(n17148) );
  AOI22_X1 U16106 ( .A1(n9838), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n17148), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n13029) );
  INV_X2 U16107 ( .A(n13240), .ZN(n17193) );
  AOI22_X1 U16108 ( .A1(n9849), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n17193), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n13028) );
  NAND4_X1 U16109 ( .A1(n13031), .A2(n13030), .A3(n13029), .A4(n13028), .ZN(
        n13032) );
  AOI211_X1 U16110 ( .C1(n17098), .C2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A(
        n13033), .B(n13032), .ZN(n13034) );
  NAND3_X1 U16111 ( .A1(n13036), .A2(n13035), .A3(n13034), .ZN(n13281) );
  AOI22_X1 U16112 ( .A1(n9849), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(n9837), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n13046) );
  AOI22_X1 U16113 ( .A1(n17193), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n9839), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n13045) );
  AOI22_X1 U16114 ( .A1(n17211), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17213), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n13037) );
  OAI21_X1 U16115 ( .B1(n13161), .B2(n21055), .A(n13037), .ZN(n13043) );
  AOI22_X1 U16116 ( .A1(n17199), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17216), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n13041) );
  INV_X2 U16117 ( .A(n9887), .ZN(n17219) );
  INV_X2 U16118 ( .A(n9888), .ZN(n17112) );
  AOI22_X1 U16119 ( .A1(n17219), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n17112), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n13040) );
  AOI22_X1 U16120 ( .A1(n17153), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n17148), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n13039) );
  AOI22_X1 U16121 ( .A1(n17194), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n9838), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n13038) );
  NAND4_X1 U16122 ( .A1(n13041), .A2(n13040), .A3(n13039), .A4(n13038), .ZN(
        n13042) );
  AOI211_X1 U16123 ( .C1(n17200), .C2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A(
        n13043), .B(n13042), .ZN(n13044) );
  NAND3_X1 U16124 ( .A1(n13046), .A2(n13045), .A3(n13044), .ZN(n13284) );
  AOI22_X1 U16125 ( .A1(n9851), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n13065), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n13051) );
  INV_X2 U16126 ( .A(n13161), .ZN(n17177) );
  AOI22_X1 U16127 ( .A1(n17199), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17177), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n13050) );
  AOI22_X1 U16128 ( .A1(n9832), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n17148), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n13049) );
  AOI22_X1 U16129 ( .A1(n13013), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n9837), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n13048) );
  NAND4_X1 U16130 ( .A1(n13051), .A2(n13050), .A3(n13049), .A4(n13048), .ZN(
        n13057) );
  AOI22_X1 U16131 ( .A1(n17153), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n13088), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n13055) );
  AOI22_X1 U16132 ( .A1(n17217), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n9838), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n13054) );
  INV_X1 U16133 ( .A(n9888), .ZN(n17176) );
  AOI22_X1 U16134 ( .A1(n17176), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n13058), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n13053) );
  AOI22_X1 U16135 ( .A1(n13160), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n17216), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n13052) );
  NAND4_X1 U16136 ( .A1(n13055), .A2(n13054), .A3(n13053), .A4(n13052), .ZN(
        n13056) );
  NOR2_X2 U16137 ( .A1(n13057), .A2(n13056), .ZN(n17414) );
  AOI22_X1 U16138 ( .A1(n17219), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n13011), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n13062) );
  AOI22_X1 U16139 ( .A1(n9832), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n13160), .ZN(n13061) );
  AOI22_X1 U16140 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n17148), .B1(
        P3_INSTQUEUE_REG_12__1__SCAN_IN), .B2(n17192), .ZN(n13060) );
  AOI22_X1 U16141 ( .A1(n13013), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_6__1__SCAN_IN), .B2(n13058), .ZN(n13059) );
  AOI22_X1 U16142 ( .A1(n13047), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n13063), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n13064) );
  OAI21_X1 U16143 ( .B1(n9888), .B2(n21120), .A(n13064), .ZN(n13071) );
  INV_X2 U16144 ( .A(n10259), .ZN(n17212) );
  AOI22_X1 U16145 ( .A1(n17212), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_3__1__SCAN_IN), .B2(n9838), .ZN(n13069) );
  AOI22_X1 U16146 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n9837), .B1(
        n13065), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n13068) );
  NAND3_X1 U16147 ( .A1(n13069), .A2(n13068), .A3(n13067), .ZN(n13070) );
  AOI22_X1 U16148 ( .A1(n9849), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n17177), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n13076) );
  AOI22_X1 U16149 ( .A1(n9832), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17112), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n13075) );
  AOI22_X1 U16150 ( .A1(n9838), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17213), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n13074) );
  AOI22_X1 U16151 ( .A1(n17212), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n17148), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n13073) );
  NAND4_X1 U16152 ( .A1(n13076), .A2(n13075), .A3(n13074), .A4(n13073), .ZN(
        n13083) );
  INV_X2 U16153 ( .A(n13219), .ZN(n17147) );
  AOI22_X1 U16154 ( .A1(n17147), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n9839), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n13081) );
  AOI22_X1 U16155 ( .A1(n17199), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17193), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n13080) );
  AOI22_X1 U16156 ( .A1(n9837), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17211), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n13079) );
  AOI22_X1 U16157 ( .A1(n17219), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n17194), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n13078) );
  NAND4_X1 U16158 ( .A1(n13081), .A2(n13080), .A3(n13079), .A4(n13078), .ZN(
        n13082) );
  AOI22_X1 U16159 ( .A1(n17176), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n9838), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n13087) );
  AOI22_X1 U16160 ( .A1(n17199), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17177), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n13086) );
  AOI22_X1 U16161 ( .A1(n9832), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17148), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13085) );
  AOI22_X1 U16162 ( .A1(n9851), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(n9849), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n13084) );
  NAND4_X1 U16163 ( .A1(n13087), .A2(n13086), .A3(n13085), .A4(n13084), .ZN(
        n13094) );
  AOI22_X1 U16164 ( .A1(n9837), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(n9839), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n13092) );
  AOI22_X1 U16165 ( .A1(n17147), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17213), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n13091) );
  AOI22_X1 U16166 ( .A1(n17193), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17194), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n13090) );
  AOI22_X1 U16167 ( .A1(n17212), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17211), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n13089) );
  NAND4_X1 U16168 ( .A1(n13092), .A2(n13091), .A3(n13090), .A4(n13089), .ZN(
        n13093) );
  INV_X1 U16169 ( .A(n17397), .ZN(n13299) );
  INV_X1 U16170 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n17594) );
  NOR2_X1 U16171 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17818), .ZN(
        n17685) );
  INV_X1 U16172 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n18015) );
  NAND2_X1 U16173 ( .A1(n17685), .A2(n18015), .ZN(n13095) );
  NOR2_X1 U16174 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n13095), .ZN(
        n17651) );
  INV_X1 U16175 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n17989) );
  NAND2_X1 U16176 ( .A1(n17651), .A2(n17989), .ZN(n17635) );
  NOR3_X1 U16177 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(n17635), .ZN(n13139) );
  INV_X1 U16178 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n18127) );
  INV_X1 U16179 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18116) );
  NOR2_X1 U16180 ( .A1(n18127), .A2(n18116), .ZN(n17784) );
  NAND2_X1 U16181 ( .A1(n17784), .A2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n18108) );
  INV_X1 U16182 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n18100) );
  NOR2_X1 U16183 ( .A1(n18108), .A2(n18100), .ZN(n18070) );
  NAND2_X1 U16184 ( .A1(n18070), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n18068) );
  INV_X1 U16185 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n18074) );
  NOR2_X1 U16186 ( .A1(n18068), .A2(n18074), .ZN(n18041) );
  NAND2_X1 U16187 ( .A1(n18041), .A2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n18024) );
  XOR2_X1 U16188 ( .A(n17401), .B(n13096), .Z(n13119) );
  NAND2_X1 U16189 ( .A1(n13108), .A2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13109) );
  AOI22_X1 U16190 ( .A1(n17176), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17213), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n13106) );
  AOI22_X1 U16191 ( .A1(n17212), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n17216), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n13105) );
  INV_X1 U16192 ( .A(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n21111) );
  AOI22_X1 U16193 ( .A1(n13065), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n9838), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n13097) );
  OAI21_X1 U16194 ( .B1(n9887), .B2(n21111), .A(n13097), .ZN(n13103) );
  AOI22_X1 U16195 ( .A1(n13013), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n13011), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n13101) );
  AOI22_X1 U16196 ( .A1(n9837), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n13058), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n13100) );
  AOI22_X1 U16197 ( .A1(n13066), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n13160), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n13099) );
  AOI22_X1 U16198 ( .A1(n13047), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n17148), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n13098) );
  NAND4_X1 U16199 ( .A1(n13101), .A2(n13100), .A3(n13099), .A4(n13098), .ZN(
        n13102) );
  AOI211_X1 U16200 ( .C1(n9832), .C2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A(
        n13103), .B(n13102), .ZN(n13104) );
  INV_X1 U16201 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n18226) );
  NAND2_X1 U16202 ( .A1(n13109), .A2(n17900), .ZN(n17890) );
  XOR2_X1 U16203 ( .A(n17414), .B(n17421), .Z(n13110) );
  XNOR2_X1 U16204 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n13110), .ZN(
        n17891) );
  INV_X1 U16205 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n13287) );
  NAND2_X1 U16206 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n13113), .ZN(
        n13115) );
  INV_X1 U16207 ( .A(n13284), .ZN(n17409) );
  XNOR2_X1 U16208 ( .A(n17409), .B(n13114), .ZN(n18190) );
  NAND2_X1 U16209 ( .A1(n13115), .A2(n17879), .ZN(n17860) );
  INV_X1 U16210 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n18187) );
  XNOR2_X1 U16211 ( .A(n17405), .B(n13116), .ZN(n13117) );
  XNOR2_X1 U16212 ( .A(n18187), .B(n13117), .ZN(n17861) );
  NAND2_X1 U16213 ( .A1(n17860), .A2(n17861), .ZN(n17859) );
  NAND2_X1 U16214 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n13117), .ZN(
        n13118) );
  NAND2_X1 U16215 ( .A1(n13119), .A2(n13121), .ZN(n13122) );
  NAND2_X1 U16216 ( .A1(n13122), .A2(n17845), .ZN(n17836) );
  INV_X1 U16217 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n18163) );
  XNOR2_X1 U16218 ( .A(n17397), .B(n13123), .ZN(n13124) );
  XNOR2_X1 U16219 ( .A(n18163), .B(n13124), .ZN(n17837) );
  NAND2_X1 U16220 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n13124), .ZN(
        n13125) );
  AOI21_X1 U16221 ( .B1(n17393), .B2(n13126), .A(n17818), .ZN(n13129) );
  NAND2_X1 U16222 ( .A1(n17824), .A2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n17823) );
  NAND2_X1 U16223 ( .A1(n13129), .A2(n13128), .ZN(n13130) );
  INV_X1 U16224 ( .A(n13133), .ZN(n13131) );
  INV_X1 U16225 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n20983) );
  NAND2_X1 U16226 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n18018) );
  NAND2_X1 U16227 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n17988) );
  INV_X1 U16228 ( .A(n17988), .ZN(n17653) );
  NAND3_X1 U16229 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(n17653), .ZN(n13141) );
  NOR2_X1 U16230 ( .A1(n18018), .A2(n13141), .ZN(n17976) );
  NAND2_X1 U16231 ( .A1(n17976), .A2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n17964) );
  NOR2_X1 U16232 ( .A1(n20983), .A2(n17964), .ZN(n17608) );
  NOR4_X1 U16233 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A4(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n13135) );
  NOR2_X1 U16234 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n17774) );
  NAND3_X1 U16235 ( .A1(n13133), .A2(n17774), .A3(n13132), .ZN(n13134) );
  OAI21_X1 U16236 ( .B1(n17818), .B2(n13135), .A(n17756), .ZN(n17704) );
  INV_X1 U16237 ( .A(n17704), .ZN(n13137) );
  INV_X1 U16238 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n18043) );
  INV_X1 U16239 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n21008) );
  NAND2_X2 U16240 ( .A1(n17695), .A2(n17757), .ZN(n17659) );
  OAI221_X1 U16241 ( .B1(n13139), .B2(n13138), .C1(n13139), .C2(n17608), .A(
        n17659), .ZN(n17606) );
  NOR2_X2 U16242 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17606), .ZN(
        n17605) );
  INV_X1 U16243 ( .A(n17659), .ZN(n13140) );
  INV_X1 U16244 ( .A(n17605), .ZN(n17593) );
  NAND2_X1 U16245 ( .A1(n17757), .A2(n17593), .ZN(n13142) );
  OAI221_X1 U16246 ( .B1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n17757), 
        .C1(n17594), .C2(n9892), .A(n13142), .ZN(n17571) );
  NOR2_X1 U16247 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n17571), .ZN(
        n17570) );
  NOR2_X1 U16248 ( .A1(n9892), .A2(n17757), .ZN(n17592) );
  INV_X1 U16249 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n13143) );
  NOR2_X1 U16250 ( .A1(n17594), .A2(n13143), .ZN(n15836) );
  INV_X1 U16251 ( .A(n15836), .ZN(n17923) );
  AND2_X1 U16252 ( .A1(n17818), .A2(n17923), .ZN(n13144) );
  NOR2_X2 U16253 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n13147), .ZN(
        n17559) );
  INV_X1 U16254 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n17553) );
  NAND2_X1 U16255 ( .A1(n17559), .A2(n17553), .ZN(n15820) );
  OAI21_X1 U16256 ( .B1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n15820), .A(
        n17757), .ZN(n15906) );
  INV_X1 U16257 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n18848) );
  NOR2_X1 U16258 ( .A1(n18848), .A2(n17757), .ZN(n13150) );
  NOR2_X1 U16259 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n17818), .ZN(
        n13146) );
  INV_X1 U16260 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15837) );
  NOR2_X1 U16261 ( .A1(n15837), .A2(n17553), .ZN(n16426) );
  NAND2_X1 U16262 ( .A1(n16426), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16436) );
  NAND2_X1 U16263 ( .A1(n15907), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n13154) );
  AOI21_X1 U16264 ( .B1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n18848), .A(
        n13148), .ZN(n13149) );
  NAND2_X1 U16265 ( .A1(n13149), .A2(n15906), .ZN(n13153) );
  AOI22_X1 U16266 ( .A1(n18848), .A2(n17757), .B1(n13150), .B2(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n13151) );
  INV_X1 U16267 ( .A(n13151), .ZN(n13152) );
  AOI22_X2 U16268 ( .A1(n13155), .A2(n13154), .B1(n13153), .B2(n13152), .ZN(
        n16442) );
  AOI22_X1 U16269 ( .A1(n9837), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n17211), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n13159) );
  AOI22_X1 U16270 ( .A1(n17112), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_4__1__SCAN_IN), .B2(n17147), .ZN(n13158) );
  AOI22_X1 U16271 ( .A1(n17192), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n15785), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n13157) );
  AOI22_X1 U16272 ( .A1(n9838), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(n9839), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n13156) );
  NAND4_X1 U16273 ( .A1(n13159), .A2(n13158), .A3(n13157), .A4(n13156), .ZN(
        n13167) );
  AOI22_X1 U16274 ( .A1(n17098), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n9849), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n13165) );
  INV_X2 U16275 ( .A(n17080), .ZN(n17200) );
  AOI22_X1 U16276 ( .A1(n9851), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n17200), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n13164) );
  INV_X2 U16277 ( .A(n13161), .ZN(n17220) );
  AOI22_X1 U16278 ( .A1(n17220), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n17194), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n13163) );
  AOI22_X1 U16279 ( .A1(n17193), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n17153), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n13162) );
  NAND4_X1 U16280 ( .A1(n13165), .A2(n13164), .A3(n13163), .A4(n13162), .ZN(
        n13166) );
  NAND2_X1 U16281 ( .A1(n18236), .A2(P3_STATE2_REG_0__SCAN_IN), .ZN(n18747) );
  NOR2_X1 U16282 ( .A1(n18886), .A2(n18743), .ZN(n14393) );
  AOI22_X1 U16283 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n18718), .B1(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n18862), .ZN(n13268) );
  NOR2_X1 U16284 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18727), .ZN(
        n13171) );
  NAND2_X1 U16285 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n13170), .ZN(
        n13175) );
  AOI22_X1 U16286 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n13176), .B1(
        n13171), .B2(n13175), .ZN(n13179) );
  AOI21_X1 U16287 ( .B1(n18870), .B2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(
        n13267), .ZN(n13271) );
  AND2_X1 U16288 ( .A1(n13268), .A2(n13271), .ZN(n13178) );
  OAI21_X1 U16289 ( .B1(n13174), .B2(n13173), .A(n13179), .ZN(n13172) );
  INV_X1 U16290 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n18691) );
  AOI211_X2 U16291 ( .C1(n13179), .C2(n13178), .A(n13272), .B(n13269), .ZN(
        n18682) );
  AOI22_X1 U16292 ( .A1(n17200), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n9837), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n13183) );
  AOI22_X1 U16293 ( .A1(n9851), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17153), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n13182) );
  AOI22_X1 U16294 ( .A1(n17217), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n9838), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n13181) );
  AOI22_X1 U16295 ( .A1(n13160), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n17148), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n13180) );
  NAND4_X1 U16296 ( .A1(n13183), .A2(n13182), .A3(n13181), .A4(n13180), .ZN(
        n13189) );
  AOI22_X1 U16297 ( .A1(n17112), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17213), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n13187) );
  AOI22_X1 U16298 ( .A1(n17098), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17177), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n13186) );
  AOI22_X1 U16299 ( .A1(n17193), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17211), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n13185) );
  AOI22_X1 U16300 ( .A1(n17147), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n9839), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n13184) );
  NAND4_X1 U16301 ( .A1(n13187), .A2(n13186), .A3(n13185), .A4(n13184), .ZN(
        n13188) );
  AOI22_X1 U16302 ( .A1(n17112), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n13058), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n13193) );
  AOI22_X1 U16303 ( .A1(n17212), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n17220), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n13192) );
  AOI22_X1 U16304 ( .A1(n17219), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n9837), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n13191) );
  AOI22_X1 U16305 ( .A1(n17199), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n15785), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n13190) );
  AOI22_X1 U16306 ( .A1(n9849), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(n9838), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n13197) );
  AOI22_X1 U16307 ( .A1(n17200), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n17194), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n13196) );
  AOI22_X1 U16308 ( .A1(n17193), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n17147), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n13195) );
  AOI22_X1 U16309 ( .A1(n17211), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n17192), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n13194) );
  AOI22_X1 U16310 ( .A1(n17112), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n9837), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n13201) );
  AOI22_X1 U16311 ( .A1(n17193), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17153), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n13200) );
  AOI22_X1 U16312 ( .A1(n17220), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17211), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n13199) );
  AOI22_X1 U16313 ( .A1(n9839), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n15785), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n13198) );
  NAND4_X1 U16314 ( .A1(n13201), .A2(n13200), .A3(n13199), .A4(n13198), .ZN(
        n13207) );
  AOI22_X1 U16315 ( .A1(n9851), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17213), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n13205) );
  AOI22_X1 U16316 ( .A1(n17098), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17147), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n13204) );
  AOI22_X1 U16317 ( .A1(n9849), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n17194), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n13203) );
  AOI22_X1 U16318 ( .A1(n17200), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n9838), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n13202) );
  NAND4_X1 U16319 ( .A1(n13205), .A2(n13204), .A3(n13203), .A4(n13202), .ZN(
        n13206) );
  NOR2_X2 U16320 ( .A1(n18277), .A2(n18258), .ZN(n13264) );
  AOI22_X1 U16321 ( .A1(n17193), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n9839), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n13211) );
  AOI22_X1 U16322 ( .A1(n17098), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17147), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13210) );
  AOI22_X1 U16323 ( .A1(n17220), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n13065), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n13209) );
  AOI22_X1 U16324 ( .A1(n9849), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n15785), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n13208) );
  NAND4_X1 U16325 ( .A1(n13211), .A2(n13210), .A3(n13209), .A4(n13208), .ZN(
        n13217) );
  AOI22_X1 U16326 ( .A1(n17217), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n9838), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n13215) );
  AOI22_X1 U16327 ( .A1(n17112), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n9837), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n13214) );
  AOI22_X1 U16328 ( .A1(n17153), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17213), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n13213) );
  AOI22_X1 U16329 ( .A1(n9851), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17200), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n13212) );
  NAND4_X1 U16330 ( .A1(n13215), .A2(n13214), .A3(n13213), .A4(n13212), .ZN(
        n13216) );
  AOI22_X1 U16331 ( .A1(n17193), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17112), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n13228) );
  AOI22_X1 U16332 ( .A1(n17220), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n17194), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n13227) );
  INV_X1 U16333 ( .A(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n21013) );
  AOI22_X1 U16334 ( .A1(n9837), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n13058), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n13218) );
  OAI21_X1 U16335 ( .B1(n13219), .B2(n21013), .A(n13218), .ZN(n13225) );
  AOI22_X1 U16336 ( .A1(n17098), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n9838), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n13223) );
  AOI22_X1 U16337 ( .A1(n17219), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n17153), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n13222) );
  AOI22_X1 U16338 ( .A1(n13160), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n17211), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n13221) );
  AOI22_X1 U16339 ( .A1(n17192), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n15785), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n13220) );
  NAND4_X1 U16340 ( .A1(n13223), .A2(n13222), .A3(n13221), .A4(n13220), .ZN(
        n13224) );
  NOR2_X1 U16341 ( .A1(n18267), .A2(n13273), .ZN(n15826) );
  AOI22_X1 U16342 ( .A1(n17200), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n9837), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n13232) );
  AOI22_X1 U16343 ( .A1(n17098), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17112), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n13231) );
  AOI22_X1 U16344 ( .A1(n17193), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n9838), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n13230) );
  AOI22_X1 U16345 ( .A1(n17211), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n15785), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n13229) );
  NAND4_X1 U16346 ( .A1(n13232), .A2(n13231), .A3(n13230), .A4(n13229), .ZN(
        n13238) );
  AOI22_X1 U16347 ( .A1(n9849), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n17147), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n13236) );
  AOI22_X1 U16348 ( .A1(n17220), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17213), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n13235) );
  AOI22_X1 U16349 ( .A1(n17217), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n9839), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n13234) );
  AOI22_X1 U16350 ( .A1(n17219), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n17153), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n13233) );
  NAND4_X1 U16351 ( .A1(n13236), .A2(n13235), .A3(n13234), .A4(n13233), .ZN(
        n13237) );
  AOI22_X1 U16352 ( .A1(n9838), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(n9839), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n13249) );
  AOI22_X1 U16353 ( .A1(n9849), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n17211), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n13248) );
  AOI22_X1 U16354 ( .A1(n17217), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17112), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n13239) );
  OAI21_X1 U16355 ( .B1(n13240), .B2(n21007), .A(n13239), .ZN(n13246) );
  AOI22_X1 U16356 ( .A1(n17219), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n17200), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n13244) );
  AOI22_X1 U16357 ( .A1(n17153), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17216), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n13243) );
  AOI22_X1 U16358 ( .A1(n17220), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17213), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n13242) );
  AOI22_X1 U16359 ( .A1(n9837), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n15785), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n13241) );
  NAND4_X1 U16360 ( .A1(n13244), .A2(n13243), .A3(n13242), .A4(n13241), .ZN(
        n13245) );
  NOR2_X1 U16361 ( .A1(n18262), .A2(n13274), .ZN(n18695) );
  NAND3_X1 U16362 ( .A1(n13264), .A2(n15826), .A3(n18695), .ZN(n15812) );
  NOR2_X2 U16363 ( .A1(n18903), .A2(n15812), .ZN(n18710) );
  NOR2_X2 U16364 ( .A1(n13262), .A2(n13273), .ZN(n18694) );
  NAND4_X1 U16365 ( .A1(n13264), .A2(n18267), .A3(n13257), .A4(n17428), .ZN(
        n13250) );
  NAND2_X1 U16366 ( .A1(n17275), .A2(n13274), .ZN(n13256) );
  NAND2_X1 U16367 ( .A1(n13263), .A2(n13273), .ZN(n15805) );
  NAND2_X1 U16368 ( .A1(n13250), .A2(n15805), .ZN(n16559) );
  INV_X1 U16369 ( .A(n13250), .ZN(n17490) );
  NOR2_X1 U16370 ( .A1(n18248), .A2(n16589), .ZN(n13252) );
  NOR2_X1 U16371 ( .A1(n13274), .A2(n18267), .ZN(n18713) );
  OR2_X1 U16372 ( .A1(n18277), .A2(n18713), .ZN(n15922) );
  NAND2_X1 U16373 ( .A1(n13252), .A2(n15922), .ZN(n15808) );
  OAI21_X1 U16374 ( .B1(n15826), .B2(n13257), .A(n15808), .ZN(n13261) );
  AOI22_X1 U16375 ( .A1(n18258), .A2(n13253), .B1(n18262), .B2(n18713), .ZN(
        n13260) );
  INV_X1 U16376 ( .A(n13273), .ZN(n18254) );
  NAND2_X1 U16377 ( .A1(n18248), .A2(n16589), .ZN(n13254) );
  NAND2_X1 U16378 ( .A1(n18254), .A2(n13254), .ZN(n13276) );
  AOI21_X1 U16379 ( .B1(n17356), .B2(n13256), .A(n18262), .ZN(n13255) );
  AOI21_X1 U16380 ( .B1(n13256), .B2(n13276), .A(n13255), .ZN(n13259) );
  NOR2_X1 U16381 ( .A1(n13273), .A2(n13256), .ZN(n15831) );
  OAI21_X1 U16382 ( .B1(n13257), .B2(n15831), .A(n18248), .ZN(n13258) );
  NAND3_X1 U16383 ( .A1(n13260), .A2(n13259), .A3(n13258), .ZN(n15806) );
  NAND2_X1 U16384 ( .A1(n13263), .A2(n13266), .ZN(n15815) );
  INV_X1 U16385 ( .A(n13264), .ZN(n13275) );
  NAND3_X1 U16386 ( .A1(n13275), .A2(n16589), .A3(n15802), .ZN(n13265) );
  NAND2_X1 U16387 ( .A1(n13266), .A2(n13265), .ZN(n18693) );
  AOI21_X4 U16388 ( .B1(n18694), .B2(n15803), .A(n18693), .ZN(n18692) );
  XOR2_X1 U16389 ( .A(n13268), .B(n13267), .Z(n13270) );
  INV_X1 U16390 ( .A(n18685), .ZN(n15825) );
  AOI21_X1 U16391 ( .B1(n13272), .B2(n13271), .A(n15825), .ZN(n18686) );
  NOR2_X1 U16392 ( .A1(n18886), .A2(n13273), .ZN(n15824) );
  NAND2_X1 U16393 ( .A1(n15824), .A2(n13274), .ZN(n15822) );
  NOR3_X1 U16394 ( .A1(n13277), .A2(n13276), .A3(n13275), .ZN(n13278) );
  OAI21_X1 U16395 ( .B1(n18262), .B2(n18713), .A(n13278), .ZN(n15807) );
  NOR2_X2 U16396 ( .A1(n17393), .A2(n17913), .ZN(n17819) );
  NAND2_X1 U16397 ( .A1(n16442), .A2(n17819), .ZN(n13323) );
  INV_X1 U16398 ( .A(n17976), .ZN(n17639) );
  NAND4_X1 U16399 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A4(n15836), .ZN(n15840) );
  NOR2_X1 U16400 ( .A1(n17639), .A2(n15840), .ZN(n17925) );
  INV_X1 U16401 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n18059) );
  INV_X1 U16402 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n18144) );
  NAND2_X1 U16403 ( .A1(n18041), .A2(n18022), .ZN(n17738) );
  NAND2_X1 U16404 ( .A1(n17925), .A2(n18048), .ZN(n17916) );
  NOR2_X1 U16405 ( .A1(n16436), .A2(n17916), .ZN(n16425) );
  NAND2_X1 U16406 ( .A1(n16425), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n13280) );
  XNOR2_X1 U16407 ( .A(n13280), .B(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n16443) );
  NAND2_X1 U16408 ( .A1(n17898), .A2(n17421), .ZN(n13285) );
  NAND2_X1 U16409 ( .A1(n17414), .A2(n13285), .ZN(n13283) );
  NAND2_X1 U16410 ( .A1(n13283), .A2(n13284), .ZN(n13294) );
  NOR2_X1 U16411 ( .A1(n17405), .A2(n13294), .ZN(n13282) );
  NAND2_X1 U16412 ( .A1(n13282), .A2(n13281), .ZN(n13300) );
  NOR2_X1 U16413 ( .A1(n17397), .A2(n13300), .ZN(n13305) );
  NAND2_X1 U16414 ( .A1(n13305), .A2(n13304), .ZN(n13306) );
  XNOR2_X1 U16415 ( .A(n13282), .B(n17401), .ZN(n13297) );
  AND2_X1 U16416 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n13297), .ZN(
        n13298) );
  XNOR2_X1 U16417 ( .A(n13284), .B(n13283), .ZN(n13291) );
  NOR2_X1 U16418 ( .A1(n13291), .A2(n13112), .ZN(n13292) );
  XOR2_X1 U16419 ( .A(n17414), .B(n13285), .Z(n13286) );
  NOR2_X1 U16420 ( .A1(n13286), .A2(n13287), .ZN(n13290) );
  XNOR2_X1 U16421 ( .A(n13287), .B(n13286), .ZN(n17886) );
  NOR2_X1 U16422 ( .A1(n13108), .A2(n18226), .ZN(n13289) );
  NAND3_X1 U16423 ( .A1(n17908), .A2(n13108), .A3(n18226), .ZN(n13288) );
  OAI221_X1 U16424 ( .B1(n13289), .B2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .C1(
        n17908), .C2(n13108), .A(n13288), .ZN(n17885) );
  NOR2_X1 U16425 ( .A1(n17886), .A2(n17885), .ZN(n17884) );
  NOR2_X1 U16426 ( .A1(n13290), .A2(n17884), .ZN(n17874) );
  XNOR2_X1 U16427 ( .A(n13291), .B(n13112), .ZN(n17873) );
  NOR2_X1 U16428 ( .A1(n17874), .A2(n17873), .ZN(n17872) );
  NOR2_X1 U16429 ( .A1(n13292), .A2(n17872), .ZN(n13295) );
  NOR2_X1 U16430 ( .A1(n13295), .A2(n18187), .ZN(n13296) );
  XOR2_X1 U16431 ( .A(n13294), .B(n13293), .Z(n17866) );
  XNOR2_X1 U16432 ( .A(n18187), .B(n13295), .ZN(n17865) );
  NOR2_X1 U16433 ( .A1(n17866), .A2(n17865), .ZN(n17864) );
  NOR2_X1 U16434 ( .A1(n13296), .A2(n17864), .ZN(n17849) );
  XNOR2_X1 U16435 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B(n13297), .ZN(
        n17848) );
  XOR2_X1 U16436 ( .A(n13300), .B(n13299), .Z(n13302) );
  NOR2_X1 U16437 ( .A1(n13301), .A2(n13302), .ZN(n13303) );
  XNOR2_X1 U16438 ( .A(n13302), .B(n13301), .ZN(n17839) );
  NOR2_X1 U16439 ( .A1(n13303), .A2(n17838), .ZN(n13307) );
  XNOR2_X1 U16440 ( .A(n13305), .B(n13304), .ZN(n13308) );
  NAND2_X1 U16441 ( .A1(n13307), .A2(n13308), .ZN(n17828) );
  NAND2_X1 U16442 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n17828), .ZN(
        n13310) );
  NOR2_X1 U16443 ( .A1(n13306), .A2(n13310), .ZN(n13312) );
  INV_X1 U16444 ( .A(n13306), .ZN(n13311) );
  OR2_X1 U16445 ( .A1(n13308), .A2(n13307), .ZN(n17829) );
  OAI21_X1 U16446 ( .B1(n13311), .B2(n13310), .A(n17829), .ZN(n13309) );
  AOI21_X1 U16447 ( .B1(n13311), .B2(n13310), .A(n13309), .ZN(n17816) );
  NAND2_X1 U16448 ( .A1(n18058), .A2(n17925), .ZN(n17917) );
  NOR2_X1 U16449 ( .A1(n17917), .A2(n16436), .ZN(n16427) );
  NAND2_X1 U16450 ( .A1(n16427), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n13313) );
  XOR2_X1 U16451 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n13313), .Z(
        n16446) );
  NOR2_X2 U16452 ( .A1(n16589), .A2(n16560), .ZN(n17894) );
  NAND2_X1 U16453 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n17867) );
  NOR2_X1 U16454 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n18902) );
  INV_X1 U16455 ( .A(n18902), .ZN(n18849) );
  INV_X1 U16456 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n18864) );
  NAND2_X1 U16457 ( .A1(n18901), .A2(n18864), .ZN(n16556) );
  AND2_X1 U16458 ( .A1(n18849), .A2(n16556), .ZN(n18883) );
  NOR2_X2 U16459 ( .A1(n17888), .A2(n16924), .ZN(n17868) );
  NAND2_X1 U16460 ( .A1(n17868), .A2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n17851) );
  NOR2_X2 U16461 ( .A1(n17851), .A2(n17852), .ZN(n17853) );
  NAND2_X1 U16462 ( .A1(n17853), .A2(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n16854) );
  NOR2_X2 U16463 ( .A1(n17904), .A2(n16854), .ZN(n16779) );
  NAND2_X1 U16464 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n17810) );
  NAND2_X2 U16465 ( .A1(n16779), .A2(n17745), .ZN(n17748) );
  INV_X1 U16466 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n17763) );
  NOR2_X1 U16467 ( .A1(n17763), .A2(n17751), .ZN(n17744) );
  NAND2_X1 U16468 ( .A1(n17744), .A2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n17714) );
  NOR2_X4 U16469 ( .A1(n17748), .A2(n17714), .ZN(n17710) );
  INV_X2 U16470 ( .A(n16762), .ZN(n16751) );
  NOR2_X4 U16471 ( .A1(n16750), .A2(n17693), .ZN(n17670) );
  NAND2_X1 U16472 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n17672) );
  OR2_X2 U16473 ( .A1(n16730), .A2(n17672), .ZN(n17629) );
  INV_X1 U16474 ( .A(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n17663) );
  NOR2_X2 U16475 ( .A1(n17629), .A2(n17663), .ZN(n16582) );
  NAND2_X1 U16476 ( .A1(n16582), .A2(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n16581) );
  INV_X1 U16477 ( .A(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n17618) );
  NOR2_X2 U16478 ( .A1(n17586), .A2(n17618), .ZN(n16579) );
  NAND3_X2 U16479 ( .A1(n16579), .A2(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n17542) );
  INV_X1 U16480 ( .A(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n17574) );
  NOR2_X2 U16481 ( .A1(n17542), .A2(n17574), .ZN(n16572) );
  NAND3_X1 U16482 ( .A1(n16572), .A2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n16573) );
  INV_X1 U16483 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n16610) );
  NOR2_X2 U16484 ( .A1(n16573), .A2(n16610), .ZN(n16417) );
  NAND2_X1 U16485 ( .A1(n16417), .A2(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n13315) );
  INV_X4 U16486 ( .A(n9843), .ZN(n16789) );
  INV_X1 U16487 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n18823) );
  INV_X1 U16488 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n18891) );
  NOR2_X1 U16489 ( .A1(n18823), .A2(n18218), .ZN(n16440) );
  INV_X1 U16490 ( .A(n16854), .ZN(n17746) );
  NAND2_X1 U16491 ( .A1(n17746), .A2(n17745), .ZN(n17733) );
  NOR2_X1 U16492 ( .A1(n17714), .A2(n17733), .ZN(n17707) );
  NAND3_X1 U16493 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A3(n17707), .ZN(n17692) );
  NOR2_X1 U16494 ( .A1(n17693), .A2(n17692), .ZN(n17671) );
  NAND3_X1 U16495 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A3(n17671), .ZN(n17662) );
  NOR2_X1 U16496 ( .A1(n17663), .A2(n17662), .ZN(n17631) );
  NAND3_X1 U16497 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A3(n17631), .ZN(n17615) );
  NOR2_X1 U16498 ( .A1(n17618), .A2(n17615), .ZN(n17599) );
  NAND3_X1 U16499 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A3(n17599), .ZN(n17573) );
  NOR2_X1 U16500 ( .A1(n17574), .A2(n17573), .ZN(n17546) );
  NAND3_X1 U16501 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A3(n17546), .ZN(n16415) );
  NOR2_X1 U16502 ( .A1(n16610), .A2(n16415), .ZN(n13316) );
  NOR2_X1 U16503 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18901), .ZN(n17630) );
  AOI221_X1 U16504 ( .B1(P3_STATE2_REG_2__SCAN_IN), .B2(n18236), .C1(n18901), 
        .C2(P3_STATE2_REG_1__SCAN_IN), .A(n18866), .ZN(n18245) );
  NOR3_X2 U16505 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(P3_STATE2_REG_3__SCAN_IN), .A3(n18887), .ZN(n18593) );
  NAND2_X1 U16506 ( .A1(n13316), .A2(n17712), .ZN(n16407) );
  INV_X1 U16507 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n20969) );
  XOR2_X1 U16508 ( .A(n20969), .B(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .Z(
        n13318) );
  NOR2_X1 U16509 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n17697), .ZN(
        n16416) );
  INV_X1 U16510 ( .A(n16573), .ZN(n16419) );
  INV_X1 U16511 ( .A(n17630), .ZN(n17909) );
  OR2_X1 U16512 ( .A1(n18343), .A2(n13316), .ZN(n13317) );
  OAI211_X1 U16513 ( .C1(n16419), .C2(n17909), .A(n17910), .B(n13317), .ZN(
        n16424) );
  NOR2_X1 U16514 ( .A1(n16416), .A2(n16424), .ZN(n16406) );
  OAI22_X1 U16515 ( .A1(n16407), .A2(n13318), .B1(n16406), .B2(n20969), .ZN(
        n13319) );
  AOI211_X1 U16516 ( .C1(n17767), .C2(n16789), .A(n16440), .B(n13319), .ZN(
        n13320) );
  NAND2_X1 U16517 ( .A1(n13323), .A2(n13322), .ZN(P3_U2799) );
  INV_X1 U16518 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n19926) );
  NOR2_X1 U16519 ( .A1(P2_BE_N_REG_0__SCAN_IN), .A2(n19926), .ZN(n13325) );
  NOR4_X1 U16520 ( .A1(P2_BE_N_REG_1__SCAN_IN), .A2(P2_BE_N_REG_2__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n13324) );
  INV_X1 U16521 ( .A(P2_BE_N_REG_3__SCAN_IN), .ZN(n20943) );
  NAND4_X1 U16522 ( .A1(P2_M_IO_N_REG_SCAN_IN), .A2(n13325), .A3(n13324), .A4(
        n20943), .ZN(n13328) );
  NOR2_X1 U16523 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n13328), .ZN(n16536)
         );
  INV_X1 U16524 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n20799) );
  NOR3_X1 U16525 ( .A1(P1_D_C_N_REG_SCAN_IN), .A2(P1_BE_N_REG_0__SCAN_IN), 
        .A3(n20799), .ZN(n13327) );
  NOR4_X1 U16526 ( .A1(P1_BE_N_REG_1__SCAN_IN), .A2(P1_BE_N_REG_2__SCAN_IN), 
        .A3(P1_BE_N_REG_3__SCAN_IN), .A4(P1_ADS_N_REG_SCAN_IN), .ZN(n13326) );
  NAND4_X1 U16527 ( .A1(n20160), .A2(P1_M_IO_N_REG_SCAN_IN), .A3(n13327), .A4(
        n13326), .ZN(U214) );
  NOR2_X1 U16528 ( .A1(n14029), .A2(n13328), .ZN(n16465) );
  NAND2_X1 U16529 ( .A1(n16465), .A2(U214), .ZN(U212) );
  INV_X1 U16530 ( .A(n9868), .ZN(n19809) );
  AOI211_X1 U16531 ( .C1(n15302), .C2(n13330), .A(n13329), .B(n19809), .ZN(
        n13344) );
  OAI22_X1 U16532 ( .A1(n13331), .A2(n19072), .B1(n21193), .B2(n19074), .ZN(
        n13343) );
  OAI22_X1 U16533 ( .A1(n13332), .A2(n19095), .B1(n15304), .B2(n19057), .ZN(
        n13342) );
  AND2_X1 U16534 ( .A1(n15175), .A2(n13333), .ZN(n13334) );
  INV_X1 U16535 ( .A(n15485), .ZN(n13340) );
  NAND2_X1 U16536 ( .A1(n13336), .A2(n13337), .ZN(n13338) );
  INV_X1 U16537 ( .A(n15486), .ZN(n13339) );
  OAI22_X1 U16538 ( .A1(n13340), .A2(n19067), .B1(n13339), .B2(n19087), .ZN(
        n13341) );
  OR4_X1 U16539 ( .A1(n13344), .A2(n13343), .A3(n13342), .A4(n13341), .ZN(
        P2_U2828) );
  AOI211_X1 U16540 ( .C1(n15378), .C2(n13346), .A(n13345), .B(n19809), .ZN(
        n13356) );
  AOI22_X1 U16541 ( .A1(P2_EBX_REG_21__SCAN_IN), .A2(n19090), .B1(
        P2_REIP_REG_21__SCAN_IN), .B2(n19091), .ZN(n13347) );
  INV_X1 U16542 ( .A(n13347), .ZN(n13355) );
  OAI22_X1 U16543 ( .A1(n13348), .A2(n19095), .B1(n11293), .B2(n19057), .ZN(
        n13354) );
  OAI21_X1 U16544 ( .B1(n15219), .B2(n13349), .A(n15201), .ZN(n15560) );
  OR2_X1 U16545 ( .A1(n15575), .A2(n13350), .ZN(n13352) );
  INV_X1 U16546 ( .A(n15547), .ZN(n13351) );
  NAND2_X1 U16547 ( .A1(n13352), .A2(n13351), .ZN(n15565) );
  OAI22_X1 U16548 ( .A1(n15560), .A2(n19067), .B1(n15565), .B2(n19087), .ZN(
        n13353) );
  OR4_X1 U16549 ( .A1(n13356), .A2(n13355), .A3(n13354), .A4(n13353), .ZN(
        P2_U2834) );
  AOI211_X1 U16550 ( .C1(n15345), .C2(n13358), .A(n13357), .B(n19809), .ZN(
        n13368) );
  OAI22_X1 U16551 ( .A1(n11753), .A2(n19072), .B1(n19860), .B2(n19074), .ZN(
        n13367) );
  OAI22_X1 U16552 ( .A1(n13359), .A2(n19095), .B1(n15343), .B2(n19057), .ZN(
        n13366) );
  NAND2_X1 U16553 ( .A1(n15203), .A2(n13360), .ZN(n13361) );
  NAND2_X1 U16554 ( .A1(n15125), .A2(n13361), .ZN(n15347) );
  OR2_X1 U16555 ( .A1(n15550), .A2(n13363), .ZN(n13364) );
  NAND2_X1 U16556 ( .A1(n13362), .A2(n13364), .ZN(n15537) );
  OAI22_X1 U16557 ( .A1(n15347), .A2(n19067), .B1(n19087), .B2(n15537), .ZN(
        n13365) );
  OR4_X1 U16558 ( .A1(n13368), .A2(n13367), .A3(n13366), .A4(n13365), .ZN(
        P2_U2832) );
  NOR2_X1 U16559 ( .A1(n13781), .A2(n20168), .ZN(n13391) );
  OAI21_X1 U16560 ( .B1(n13369), .B2(n11162), .A(n13403), .ZN(n13730) );
  AOI21_X1 U16561 ( .B1(n13723), .B2(n13391), .A(n13730), .ZN(n13380) );
  NAND2_X1 U16562 ( .A1(n9858), .A2(n13727), .ZN(n13484) );
  NAND2_X1 U16563 ( .A1(n13370), .A2(n13484), .ZN(n13378) );
  NAND2_X1 U16564 ( .A1(n15892), .A2(n13372), .ZN(n13374) );
  NAND3_X1 U16565 ( .A1(n13374), .A2(n9854), .A3(n13373), .ZN(n13375) );
  NAND2_X1 U16566 ( .A1(n15901), .A2(n13375), .ZN(n13377) );
  MUX2_X1 U16567 ( .A(n13378), .B(n13377), .S(n13376), .Z(n13379) );
  NAND2_X1 U16568 ( .A1(n13380), .A2(n13379), .ZN(n13381) );
  NAND2_X1 U16569 ( .A1(n14165), .A2(n20128), .ZN(n14170) );
  NAND2_X1 U16570 ( .A1(n11162), .A2(n9858), .ZN(n13785) );
  INV_X1 U16571 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n20122) );
  AOI21_X1 U16572 ( .B1(n14170), .B2(n14167), .A(n20122), .ZN(n13414) );
  OAI21_X1 U16573 ( .B1(n13383), .B2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n13382), .ZN(n13617) );
  OR2_X1 U16574 ( .A1(n15880), .A2(n13384), .ZN(n13489) );
  OAI211_X1 U16575 ( .C1(n20182), .C2(n13386), .A(n12536), .B(n13385), .ZN(
        n13387) );
  NOR2_X1 U16576 ( .A1(n13489), .A2(n13387), .ZN(n13388) );
  NOR2_X1 U16577 ( .A1(n13617), .A2(n16177), .ZN(n13413) );
  INV_X1 U16578 ( .A(n13961), .ZN(n13389) );
  NAND2_X1 U16579 ( .A1(n13389), .A2(n11105), .ZN(n13708) );
  AND2_X1 U16580 ( .A1(n13390), .A2(n13708), .ZN(n13408) );
  NAND2_X1 U16581 ( .A1(n13408), .A2(n13391), .ZN(n13726) );
  NAND2_X1 U16582 ( .A1(n15051), .A2(n20122), .ZN(n20149) );
  INV_X1 U16583 ( .A(n20149), .ZN(n13412) );
  INV_X1 U16584 ( .A(n13709), .ZN(n13394) );
  AND2_X1 U16585 ( .A1(n13392), .A2(n20182), .ZN(n13393) );
  AOI22_X1 U16586 ( .A1(n15892), .A2(n15891), .B1(n13394), .B2(n13393), .ZN(
        n13395) );
  OR2_X1 U16587 ( .A1(n13396), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13398) );
  NAND2_X1 U16588 ( .A1(n13398), .A2(n13397), .ZN(n14655) );
  INV_X1 U16589 ( .A(n13959), .ZN(n13404) );
  NAND2_X1 U16590 ( .A1(n13400), .A2(n13718), .ZN(n13401) );
  NAND2_X1 U16591 ( .A1(n13401), .A2(n9858), .ZN(n13402) );
  OAI211_X1 U16592 ( .C1(n13399), .C2(n13404), .A(n13403), .B(n13402), .ZN(
        n13714) );
  OAI21_X1 U16593 ( .B1(n13718), .B2(n10417), .A(n13405), .ZN(n13406) );
  INV_X1 U16594 ( .A(n13406), .ZN(n13407) );
  OAI211_X1 U16595 ( .C1(n9854), .C2(n13409), .A(n13408), .B(n13407), .ZN(
        n13410) );
  NOR2_X1 U16596 ( .A1(n13714), .A2(n13410), .ZN(n14164) );
  OR3_X1 U16597 ( .A1(n14165), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A3(
        n14164), .ZN(n14169) );
  OR2_X1 U16598 ( .A1(n20128), .A2(n14657), .ZN(n13612) );
  OAI211_X1 U16599 ( .C1(n20145), .C2(n14655), .A(n14169), .B(n13612), .ZN(
        n13411) );
  OR4_X1 U16600 ( .A1(n13414), .A2(n13413), .A3(n13412), .A4(n13411), .ZN(
        P1_U3031) );
  INV_X1 U16601 ( .A(n15891), .ZN(n20800) );
  AOI21_X1 U16602 ( .B1(n13785), .B2(n20800), .A(n13727), .ZN(n13416) );
  INV_X1 U16603 ( .A(n15892), .ZN(n13415) );
  NAND2_X1 U16604 ( .A1(n13785), .A2(n13415), .ZN(n13728) );
  AND2_X1 U16605 ( .A1(n13416), .A2(n13728), .ZN(n13417) );
  NOR2_X1 U16606 ( .A1(n20802), .A2(n13782), .ZN(n16204) );
  INV_X1 U16607 ( .A(n16204), .ZN(n16208) );
  OR2_X1 U16608 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n16208), .ZN(n20045) );
  INV_X2 U16609 ( .A(n20045), .ZN(n20811) );
  AND2_X1 U16610 ( .A1(n20064), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(P1_U2905)
         );
  OR2_X1 U16611 ( .A1(n13542), .A2(n13419), .ZN(n14363) );
  INV_X1 U16612 ( .A(n14363), .ZN(n19100) );
  INV_X1 U16613 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .ZN(n19939) );
  INV_X1 U16614 ( .A(n13437), .ZN(n13421) );
  AND2_X1 U16615 ( .A1(n19691), .A2(n19802), .ZN(n13424) );
  INV_X1 U16616 ( .A(n13424), .ZN(n13420) );
  OAI211_X1 U16617 ( .C1(n19100), .C2(n19939), .A(n13421), .B(n13420), .ZN(
        P2_U2814) );
  INV_X1 U16618 ( .A(n13433), .ZN(n13423) );
  INV_X1 U16619 ( .A(P2_CODEFETCH_REG_SCAN_IN), .ZN(n13422) );
  INV_X1 U16620 ( .A(n15767), .ZN(n19890) );
  NAND2_X1 U16621 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19735), .ZN(n19804) );
  OAI22_X1 U16622 ( .A1(n13423), .A2(n13422), .B1(n19890), .B2(n19804), .ZN(
        P2_U2816) );
  OAI21_X1 U16623 ( .B1(n13424), .B2(P2_READREQUEST_REG_SCAN_IN), .A(n13433), 
        .ZN(n13425) );
  OAI21_X1 U16624 ( .B1(n13426), .B2(n13433), .A(n13425), .ZN(P2_U3612) );
  INV_X1 U16625 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n19813) );
  NOR2_X1 U16626 ( .A1(n12434), .A2(n13537), .ZN(n13430) );
  OAI21_X1 U16627 ( .B1(P2_STATEBS16_REG_SCAN_IN), .B2(n13427), .A(n19818), 
        .ZN(n13429) );
  AOI21_X1 U16628 ( .B1(P2_STATE2_REG_2__SCAN_IN), .B2(n19803), .A(n16399), 
        .ZN(n13428) );
  AOI21_X1 U16629 ( .B1(n13430), .B2(n13429), .A(n13428), .ZN(n13435) );
  NOR2_X1 U16630 ( .A1(n13431), .A2(n19735), .ZN(n16392) );
  NOR2_X1 U16631 ( .A1(n19915), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n19196) );
  INV_X1 U16632 ( .A(n19196), .ZN(n19169) );
  INV_X1 U16633 ( .A(n19169), .ZN(n19234) );
  NAND2_X1 U16634 ( .A1(n19803), .A2(n19234), .ZN(n13432) );
  OAI211_X1 U16635 ( .C1(P2_STATE2_REG_3__SCAN_IN), .C2(n16392), .A(n13433), 
        .B(n13432), .ZN(n13434) );
  MUX2_X1 U16636 ( .A(n19813), .B(n13435), .S(n13434), .Z(n13436) );
  INV_X1 U16637 ( .A(n13436), .ZN(P2_U3610) );
  NAND2_X1 U16638 ( .A1(n13437), .A2(n19803), .ZN(n13438) );
  AOI22_X1 U16639 ( .A1(n19237), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n19241), 
        .B2(P2_EAX_REG_2__SCAN_IN), .ZN(n13439) );
  NOR2_X2 U16640 ( .A1(n13438), .A2(n12058), .ZN(n19239) );
  OAI22_X1 U16641 ( .A1(n14029), .A2(BUF1_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n14030), .ZN(n19276) );
  INV_X1 U16642 ( .A(n19276), .ZN(n16234) );
  NAND2_X1 U16643 ( .A1(n19239), .A2(n16234), .ZN(n13501) );
  NAND2_X1 U16644 ( .A1(n13439), .A2(n13501), .ZN(P2_U2969) );
  AOI22_X1 U16645 ( .A1(n19237), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n19241), 
        .B2(P2_EAX_REG_9__SCAN_IN), .ZN(n13444) );
  INV_X1 U16646 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n13440) );
  OR2_X1 U16647 ( .A1(n14029), .A2(n13440), .ZN(n13442) );
  NAND2_X1 U16648 ( .A1(n14029), .A2(BUF2_REG_9__SCAN_IN), .ZN(n13441) );
  AND2_X1 U16649 ( .A1(n13442), .A2(n13441), .ZN(n19133) );
  INV_X1 U16650 ( .A(n19133), .ZN(n13443) );
  NAND2_X1 U16651 ( .A1(n19239), .A2(n13443), .ZN(n13518) );
  NAND2_X1 U16652 ( .A1(n13444), .A2(n13518), .ZN(P2_U2976) );
  AOI22_X1 U16653 ( .A1(n19237), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n19241), 
        .B2(P2_EAX_REG_1__SCAN_IN), .ZN(n13445) );
  AOI22_X1 U16654 ( .A1(n14030), .A2(BUF1_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n14029), .ZN(n19272) );
  INV_X1 U16655 ( .A(n19272), .ZN(n14317) );
  NAND2_X1 U16656 ( .A1(n19239), .A2(n14317), .ZN(n13526) );
  NAND2_X1 U16657 ( .A1(n13445), .A2(n13526), .ZN(P2_U2968) );
  AOI22_X1 U16658 ( .A1(n19237), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n19241), 
        .B2(P2_EAX_REG_0__SCAN_IN), .ZN(n13446) );
  INV_X1 U16659 ( .A(BUF1_REG_0__SCAN_IN), .ZN(n16516) );
  INV_X1 U16660 ( .A(BUF2_REG_0__SCAN_IN), .ZN(n21157) );
  AOI22_X1 U16661 ( .A1(n14030), .A2(n16516), .B1(n21157), .B2(n14029), .ZN(
        n19107) );
  NAND2_X1 U16662 ( .A1(n19239), .A2(n19107), .ZN(n13448) );
  NAND2_X1 U16663 ( .A1(n13446), .A2(n13448), .ZN(P2_U2967) );
  AOI22_X1 U16664 ( .A1(n19237), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n19241), 
        .B2(P2_EAX_REG_7__SCAN_IN), .ZN(n13447) );
  AOI22_X1 U16665 ( .A1(n14030), .A2(BUF1_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n14029), .ZN(n19299) );
  INV_X1 U16666 ( .A(n19299), .ZN(n15268) );
  NAND2_X1 U16667 ( .A1(n19239), .A2(n15268), .ZN(n13522) );
  NAND2_X1 U16668 ( .A1(n13447), .A2(n13522), .ZN(P2_U2974) );
  AOI22_X1 U16669 ( .A1(n19237), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(n19241), 
        .B2(P2_EAX_REG_16__SCAN_IN), .ZN(n13449) );
  NAND2_X1 U16670 ( .A1(n13449), .A2(n13448), .ZN(P2_U2952) );
  AOI22_X1 U16671 ( .A1(n19237), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n19241), 
        .B2(P2_EAX_REG_8__SCAN_IN), .ZN(n13454) );
  INV_X1 U16672 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n13450) );
  OR2_X1 U16673 ( .A1(n14029), .A2(n13450), .ZN(n13452) );
  NAND2_X1 U16674 ( .A1(n14029), .A2(BUF2_REG_8__SCAN_IN), .ZN(n13451) );
  AND2_X1 U16675 ( .A1(n13452), .A2(n13451), .ZN(n19136) );
  INV_X1 U16676 ( .A(n19136), .ZN(n13453) );
  NAND2_X1 U16677 ( .A1(n19239), .A2(n13453), .ZN(n13508) );
  NAND2_X1 U16678 ( .A1(n13454), .A2(n13508), .ZN(P2_U2975) );
  AOI22_X1 U16679 ( .A1(n19237), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n19241), 
        .B2(P2_EAX_REG_4__SCAN_IN), .ZN(n13455) );
  INV_X1 U16680 ( .A(BUF1_REG_4__SCAN_IN), .ZN(n16506) );
  INV_X1 U16681 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n18261) );
  AOI22_X1 U16682 ( .A1(n14030), .A2(n16506), .B1(n18261), .B2(n14029), .ZN(
        n19282) );
  NAND2_X1 U16683 ( .A1(n19239), .A2(n19282), .ZN(n13510) );
  NAND2_X1 U16684 ( .A1(n13455), .A2(n13510), .ZN(P2_U2971) );
  AOI22_X1 U16685 ( .A1(n19237), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n19241), 
        .B2(P2_EAX_REG_5__SCAN_IN), .ZN(n13456) );
  AOI22_X1 U16686 ( .A1(n14030), .A2(BUF1_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n14029), .ZN(n19287) );
  INV_X1 U16687 ( .A(n19287), .ZN(n15274) );
  NAND2_X1 U16688 ( .A1(n19239), .A2(n15274), .ZN(n13524) );
  NAND2_X1 U16689 ( .A1(n13456), .A2(n13524), .ZN(P2_U2972) );
  AOI22_X1 U16690 ( .A1(n19237), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n19241), 
        .B2(P2_EAX_REG_11__SCAN_IN), .ZN(n13461) );
  INV_X1 U16691 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n13457) );
  OR2_X1 U16692 ( .A1(n14029), .A2(n13457), .ZN(n13459) );
  NAND2_X1 U16693 ( .A1(n14029), .A2(BUF2_REG_11__SCAN_IN), .ZN(n13458) );
  AND2_X1 U16694 ( .A1(n13459), .A2(n13458), .ZN(n19127) );
  INV_X1 U16695 ( .A(n19127), .ZN(n13460) );
  NAND2_X1 U16696 ( .A1(n19239), .A2(n13460), .ZN(n13514) );
  NAND2_X1 U16697 ( .A1(n13461), .A2(n13514), .ZN(P2_U2978) );
  AOI22_X1 U16698 ( .A1(n19237), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n19241), 
        .B2(P2_EAX_REG_6__SCAN_IN), .ZN(n13462) );
  OAI22_X1 U16699 ( .A1(n14029), .A2(BUF1_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n14030), .ZN(n19291) );
  INV_X1 U16700 ( .A(n19291), .ZN(n16224) );
  NAND2_X1 U16701 ( .A1(n19239), .A2(n16224), .ZN(n13512) );
  NAND2_X1 U16702 ( .A1(n13462), .A2(n13512), .ZN(P2_U2973) );
  AOI22_X1 U16703 ( .A1(n19237), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n19241), 
        .B2(P2_EAX_REG_3__SCAN_IN), .ZN(n13463) );
  AOI22_X1 U16704 ( .A1(n14030), .A2(BUF1_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n14029), .ZN(n19154) );
  INV_X1 U16705 ( .A(n19154), .ZN(n15282) );
  NAND2_X1 U16706 ( .A1(n19239), .A2(n15282), .ZN(n13516) );
  NAND2_X1 U16707 ( .A1(n13463), .A2(n13516), .ZN(P2_U2970) );
  INV_X1 U16708 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n19214) );
  NAND2_X1 U16709 ( .A1(n14029), .A2(BUF2_REG_10__SCAN_IN), .ZN(n13465) );
  INV_X1 U16710 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n21071) );
  OR2_X1 U16711 ( .A1(n14029), .A2(n21071), .ZN(n13464) );
  NAND2_X1 U16712 ( .A1(n13465), .A2(n13464), .ZN(n19130) );
  NAND2_X1 U16713 ( .A1(n19239), .A2(n19130), .ZN(n13471) );
  NAND2_X1 U16714 ( .A1(n19237), .A2(P2_LWORD_REG_10__SCAN_IN), .ZN(n13466) );
  OAI211_X1 U16715 ( .C1(n19214), .C2(n19166), .A(n13471), .B(n13466), .ZN(
        P2_U2977) );
  INV_X1 U16716 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n19178) );
  NAND2_X1 U16717 ( .A1(n14029), .A2(BUF2_REG_12__SCAN_IN), .ZN(n13468) );
  INV_X1 U16718 ( .A(BUF1_REG_12__SCAN_IN), .ZN(n16495) );
  OR2_X1 U16719 ( .A1(n14029), .A2(n16495), .ZN(n13467) );
  NAND2_X1 U16720 ( .A1(n13468), .A2(n13467), .ZN(n19124) );
  NAND2_X1 U16721 ( .A1(n19239), .A2(n19124), .ZN(n13473) );
  NAND2_X1 U16722 ( .A1(n19237), .A2(P2_UWORD_REG_12__SCAN_IN), .ZN(n13469) );
  OAI211_X1 U16723 ( .C1(n19178), .C2(n19166), .A(n13473), .B(n13469), .ZN(
        P2_U2964) );
  INV_X1 U16724 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n19182) );
  NAND2_X1 U16725 ( .A1(n19237), .A2(P2_UWORD_REG_10__SCAN_IN), .ZN(n13470) );
  OAI211_X1 U16726 ( .C1(n19182), .C2(n19166), .A(n13471), .B(n13470), .ZN(
        P2_U2962) );
  INV_X1 U16727 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n19210) );
  NAND2_X1 U16728 ( .A1(n19237), .A2(P2_LWORD_REG_12__SCAN_IN), .ZN(n13472) );
  OAI211_X1 U16729 ( .C1(n19210), .C2(n19166), .A(n13473), .B(n13472), .ZN(
        P2_U2979) );
  INV_X1 U16730 ( .A(P2_LWORD_REG_15__SCAN_IN), .ZN(n13476) );
  INV_X1 U16731 ( .A(n19237), .ZN(n13500) );
  INV_X1 U16732 ( .A(n19239), .ZN(n13475) );
  AOI22_X1 U16733 ( .A1(n14030), .A2(BUF1_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n14029), .ZN(n19117) );
  INV_X1 U16734 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n13474) );
  OAI222_X1 U16735 ( .A1(n13476), .A2(n13500), .B1(n13475), .B2(n19117), .C1(
        n19166), .C2(n13474), .ZN(P2_U2982) );
  NOR2_X1 U16736 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n20786), .ZN(n14547) );
  NOR2_X1 U16737 ( .A1(P1_READREQUEST_REG_SCAN_IN), .A2(n14547), .ZN(n13479)
         );
  OAI21_X1 U16738 ( .B1(n13959), .B2(n13477), .A(n20808), .ZN(n13478) );
  OAI21_X1 U16739 ( .B1(n13479), .B2(n20808), .A(n13478), .ZN(P1_U3487) );
  OR2_X1 U16740 ( .A1(n15901), .A2(n13959), .ZN(n13483) );
  INV_X1 U16741 ( .A(n13480), .ZN(n13481) );
  NAND2_X1 U16742 ( .A1(n13481), .A2(n11161), .ZN(n13482) );
  NAND2_X1 U16743 ( .A1(n13483), .A2(n13482), .ZN(n19944) );
  OR2_X1 U16744 ( .A1(n13484), .A2(n9854), .ZN(n13485) );
  NAND2_X1 U16745 ( .A1(n13485), .A2(n20810), .ZN(n20803) );
  AOI21_X1 U16746 ( .B1(n15891), .B2(n13727), .A(n20803), .ZN(n13486) );
  OR2_X1 U16747 ( .A1(n19944), .A2(n13486), .ZN(n15884) );
  AND2_X1 U16748 ( .A1(n15884), .A2(n13736), .ZN(n19951) );
  INV_X1 U16749 ( .A(P1_MORE_REG_SCAN_IN), .ZN(n13499) );
  NOR2_X1 U16750 ( .A1(n13487), .A2(n20157), .ZN(n13488) );
  NOR2_X1 U16751 ( .A1(n13489), .A2(n13488), .ZN(n13495) );
  INV_X1 U16752 ( .A(n13726), .ZN(n13490) );
  NAND2_X1 U16753 ( .A1(n15901), .A2(n13490), .ZN(n13494) );
  OAI21_X1 U16754 ( .B1(n13492), .B2(n13491), .A(n11162), .ZN(n13493) );
  OAI211_X1 U16755 ( .C1(n15901), .C2(n13495), .A(n13494), .B(n13493), .ZN(
        n13496) );
  NAND2_X1 U16756 ( .A1(n13496), .A2(n14519), .ZN(n15881) );
  INV_X1 U16757 ( .A(n15881), .ZN(n13497) );
  NAND2_X1 U16758 ( .A1(n19951), .A2(n13497), .ZN(n13498) );
  OAI21_X1 U16759 ( .B1(n19951), .B2(n13499), .A(n13498), .ZN(P1_U3484) );
  AOI22_X1 U16760 ( .A1(n19242), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(
        P2_EAX_REG_18__SCAN_IN), .B2(n19241), .ZN(n13502) );
  NAND2_X1 U16761 ( .A1(n13502), .A2(n13501), .ZN(P2_U2954) );
  AOI22_X1 U16762 ( .A1(n19242), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(
        P2_EAX_REG_29__SCAN_IN), .B2(n19241), .ZN(n13507) );
  INV_X1 U16763 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n13503) );
  OR2_X1 U16764 ( .A1(n14029), .A2(n13503), .ZN(n13505) );
  NAND2_X1 U16765 ( .A1(n14029), .A2(BUF2_REG_13__SCAN_IN), .ZN(n13504) );
  AND2_X1 U16766 ( .A1(n13505), .A2(n13504), .ZN(n19122) );
  INV_X1 U16767 ( .A(n19122), .ZN(n13506) );
  NAND2_X1 U16768 ( .A1(n19239), .A2(n13506), .ZN(n13520) );
  NAND2_X1 U16769 ( .A1(n13507), .A2(n13520), .ZN(P2_U2965) );
  AOI22_X1 U16770 ( .A1(n19242), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(
        P2_EAX_REG_24__SCAN_IN), .B2(n19241), .ZN(n13509) );
  NAND2_X1 U16771 ( .A1(n13509), .A2(n13508), .ZN(P2_U2960) );
  AOI22_X1 U16772 ( .A1(n19242), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(
        P2_EAX_REG_20__SCAN_IN), .B2(n19241), .ZN(n13511) );
  NAND2_X1 U16773 ( .A1(n13511), .A2(n13510), .ZN(P2_U2956) );
  AOI22_X1 U16774 ( .A1(n19242), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(
        P2_EAX_REG_22__SCAN_IN), .B2(n19241), .ZN(n13513) );
  NAND2_X1 U16775 ( .A1(n13513), .A2(n13512), .ZN(P2_U2958) );
  AOI22_X1 U16776 ( .A1(n19242), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(
        P2_EAX_REG_27__SCAN_IN), .B2(n19241), .ZN(n13515) );
  NAND2_X1 U16777 ( .A1(n13515), .A2(n13514), .ZN(P2_U2963) );
  AOI22_X1 U16778 ( .A1(n19242), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n19241), 
        .B2(P2_EAX_REG_19__SCAN_IN), .ZN(n13517) );
  NAND2_X1 U16779 ( .A1(n13517), .A2(n13516), .ZN(P2_U2955) );
  AOI22_X1 U16780 ( .A1(n19242), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(
        P2_EAX_REG_25__SCAN_IN), .B2(n19241), .ZN(n13519) );
  NAND2_X1 U16781 ( .A1(n13519), .A2(n13518), .ZN(P2_U2961) );
  AOI22_X1 U16782 ( .A1(n19242), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n19241), 
        .B2(P2_EAX_REG_13__SCAN_IN), .ZN(n13521) );
  NAND2_X1 U16783 ( .A1(n13521), .A2(n13520), .ZN(P2_U2980) );
  AOI22_X1 U16784 ( .A1(n19242), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n19241), 
        .B2(P2_EAX_REG_23__SCAN_IN), .ZN(n13523) );
  NAND2_X1 U16785 ( .A1(n13523), .A2(n13522), .ZN(P2_U2959) );
  AOI22_X1 U16786 ( .A1(n19242), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n19241), 
        .B2(P2_EAX_REG_21__SCAN_IN), .ZN(n13525) );
  NAND2_X1 U16787 ( .A1(n13525), .A2(n13524), .ZN(P2_U2957) );
  AOI22_X1 U16788 ( .A1(n19242), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n19241), 
        .B2(P2_EAX_REG_17__SCAN_IN), .ZN(n13527) );
  NAND2_X1 U16789 ( .A1(n13527), .A2(n13526), .ZN(P2_U2953) );
  INV_X1 U16790 ( .A(n13542), .ZN(n13528) );
  NAND2_X1 U16791 ( .A1(n19165), .A2(n13530), .ZN(n13536) );
  INV_X1 U16792 ( .A(n16365), .ZN(n16367) );
  INV_X1 U16793 ( .A(n13531), .ZN(n16364) );
  NAND2_X1 U16794 ( .A1(n16367), .A2(n16364), .ZN(n13564) );
  INV_X1 U16795 ( .A(n13532), .ZN(n13533) );
  AND3_X1 U16796 ( .A1(n13534), .A2(n13564), .A3(n13533), .ZN(n13535) );
  NAND2_X1 U16797 ( .A1(n13536), .A2(n13535), .ZN(n16354) );
  INV_X1 U16798 ( .A(n16354), .ZN(n16380) );
  INV_X1 U16799 ( .A(n19808), .ZN(n18914) );
  NOR2_X1 U16800 ( .A1(n13537), .A2(n19915), .ZN(n16403) );
  AOI22_X1 U16801 ( .A1(n13537), .A2(P2_STATE2_REG_3__SCAN_IN), .B1(n16403), 
        .B2(P2_FLUSH_REG_SCAN_IN), .ZN(n13538) );
  OAI21_X1 U16802 ( .B1(n16380), .B2(n18914), .A(n13538), .ZN(n15783) );
  INV_X1 U16803 ( .A(n15783), .ZN(n13543) );
  INV_X1 U16804 ( .A(n13539), .ZN(n13540) );
  NAND2_X1 U16805 ( .A1(n19271), .A2(n13540), .ZN(n13541) );
  OR2_X1 U16806 ( .A1(n13542), .A2(n13541), .ZN(n16376) );
  OR3_X1 U16807 ( .A1(n13543), .A2(n19890), .A3(n16376), .ZN(n13544) );
  OAI21_X1 U16808 ( .B1(n13545), .B2(n15783), .A(n13544), .ZN(P2_U3595) );
  AOI21_X1 U16809 ( .B1(n13548), .B2(n13547), .A(n13546), .ZN(n13549) );
  XNOR2_X1 U16810 ( .A(n13549), .B(n15749), .ZN(n13692) );
  AOI22_X1 U16811 ( .A1(n13692), .A2(n16338), .B1(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n16339), .ZN(n13557) );
  XNOR2_X1 U16812 ( .A(n13551), .B(n13550), .ZN(n19906) );
  NOR2_X1 U16813 ( .A1(n15684), .A2(n19831), .ZN(n13693) );
  AOI21_X1 U16814 ( .B1(n16344), .B2(n19906), .A(n13693), .ZN(n13556) );
  AOI21_X1 U16815 ( .B1(n15749), .B2(n13553), .A(n13552), .ZN(n13694) );
  NAND2_X1 U16816 ( .A1(n16342), .A2(n13694), .ZN(n13555) );
  OAI211_X1 U16817 ( .C1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(n15613), .B(n14529), .ZN(n13554) );
  AND4_X1 U16818 ( .A1(n13557), .A2(n13556), .A3(n13555), .A4(n13554), .ZN(
        n13558) );
  OAI21_X1 U16819 ( .B1(n13584), .B2(n16326), .A(n13558), .ZN(P2_U3045) );
  INV_X1 U16820 ( .A(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n13560) );
  OAI211_X1 U16821 ( .C1(n12058), .C2(n13560), .A(n13559), .B(n19917), .ZN(
        n13561) );
  INV_X1 U16822 ( .A(n13561), .ZN(n13562) );
  INV_X1 U16823 ( .A(n13563), .ZN(n15756) );
  NAND2_X1 U16824 ( .A1(n13564), .A2(n15756), .ZN(n13565) );
  AND2_X2 U16825 ( .A1(n13565), .A2(n19808), .ZN(n15212) );
  MUX2_X1 U16826 ( .A(n10161), .B(n12115), .S(n15234), .Z(n13566) );
  OAI21_X1 U16827 ( .B1(n14119), .B2(n15215), .A(n13566), .ZN(P2_U2887) );
  AOI21_X1 U16828 ( .B1(n14119), .B2(n19116), .A(n19156), .ZN(n13579) );
  INV_X1 U16829 ( .A(n13567), .ZN(n13573) );
  INV_X1 U16830 ( .A(n13568), .ZN(n13571) );
  INV_X1 U16831 ( .A(n13569), .ZN(n13570) );
  NAND2_X1 U16832 ( .A1(n13571), .A2(n13570), .ZN(n13572) );
  NAND2_X1 U16833 ( .A1(n13573), .A2(n13572), .ZN(n16343) );
  NAND3_X1 U16834 ( .A1(n19921), .A2(n19116), .A3(n16343), .ZN(n13575) );
  OAI21_X1 U16835 ( .B1(n19140), .B2(n13576), .A(n13575), .ZN(n13577) );
  AOI21_X1 U16836 ( .B1(n19107), .B2(n19129), .A(n13577), .ZN(n13578) );
  OAI21_X1 U16837 ( .B1(n13579), .B2(n16343), .A(n13578), .ZN(P2_U2919) );
  NAND2_X1 U16838 ( .A1(n13581), .A2(n13582), .ZN(n13583) );
  MUX2_X1 U16839 ( .A(n13585), .B(n13584), .S(n15212), .Z(n13586) );
  OAI21_X1 U16840 ( .B1(n19910), .B2(n15215), .A(n13586), .ZN(P2_U2886) );
  NOR2_X1 U16841 ( .A1(n15891), .A2(n20810), .ZN(n13587) );
  INV_X1 U16842 ( .A(n13657), .ZN(n20075) );
  OR2_X1 U16843 ( .A1(n20075), .A2(n10421), .ZN(n13631) );
  INV_X1 U16844 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n14809) );
  NAND2_X1 U16845 ( .A1(n13657), .A2(n9859), .ZN(n13603) );
  INV_X1 U16846 ( .A(DATAI_15_), .ZN(n13589) );
  INV_X1 U16847 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n13588) );
  MUX2_X1 U16848 ( .A(n13589), .B(n13588), .S(n20160), .Z(n14810) );
  INV_X1 U16849 ( .A(P1_LWORD_REG_15__SCAN_IN), .ZN(n20046) );
  OAI222_X1 U16850 ( .A1(n13631), .A2(n14809), .B1(n13603), .B2(n14810), .C1(
        n13657), .C2(n20046), .ZN(P1_U2967) );
  INV_X1 U16851 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n21045) );
  NAND2_X1 U16852 ( .A1(n20047), .A2(n9854), .ZN(n13804) );
  AOI22_X1 U16853 ( .A1(P1_UWORD_REG_8__SCAN_IN), .A2(n20811), .B1(n20071), 
        .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n13590) );
  OAI21_X1 U16854 ( .B1(n21045), .B2(n13804), .A(n13590), .ZN(P1_U2912) );
  INV_X1 U16855 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n13592) );
  AOI22_X1 U16856 ( .A1(P1_UWORD_REG_12__SCAN_IN), .A2(n20811), .B1(n20071), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n13591) );
  OAI21_X1 U16857 ( .B1(n13592), .B2(n13804), .A(n13591), .ZN(P1_U2908) );
  INV_X1 U16858 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n13594) );
  AOI22_X1 U16859 ( .A1(P1_UWORD_REG_14__SCAN_IN), .A2(n20811), .B1(n20071), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .ZN(n13593) );
  OAI21_X1 U16860 ( .B1(n13594), .B2(n13804), .A(n13593), .ZN(P1_U2906) );
  INV_X1 U16861 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n13596) );
  AOI22_X1 U16862 ( .A1(P1_UWORD_REG_10__SCAN_IN), .A2(n20811), .B1(n20071), 
        .B2(P1_DATAO_REG_26__SCAN_IN), .ZN(n13595) );
  OAI21_X1 U16863 ( .B1(n13596), .B2(n13804), .A(n13595), .ZN(P1_U2910) );
  INV_X1 U16864 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n13598) );
  AOI22_X1 U16865 ( .A1(P1_UWORD_REG_13__SCAN_IN), .A2(n20811), .B1(n20071), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n13597) );
  OAI21_X1 U16866 ( .B1(n13598), .B2(n13804), .A(n13597), .ZN(P1_U2907) );
  INV_X1 U16867 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n13600) );
  AOI22_X1 U16868 ( .A1(P1_UWORD_REG_11__SCAN_IN), .A2(n20811), .B1(n20071), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n13599) );
  OAI21_X1 U16869 ( .B1(n13600), .B2(n13804), .A(n13599), .ZN(P1_U2909) );
  INV_X1 U16870 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n13602) );
  AOI22_X1 U16871 ( .A1(P1_UWORD_REG_9__SCAN_IN), .A2(n20811), .B1(n20071), 
        .B2(P1_DATAO_REG_25__SCAN_IN), .ZN(n13601) );
  OAI21_X1 U16872 ( .B1(n13602), .B2(n13804), .A(n13601), .ZN(P1_U2911) );
  MUX2_X1 U16873 ( .A(DATAI_8_), .B(BUF1_REG_8__SCAN_IN), .S(n20160), .Z(
        n14770) );
  NAND2_X1 U16874 ( .A1(n20082), .A2(n14770), .ZN(n13606) );
  NAND2_X1 U16875 ( .A1(n20075), .A2(P1_UWORD_REG_8__SCAN_IN), .ZN(n13604) );
  OAI211_X1 U16876 ( .C1(n21045), .C2(n13631), .A(n13606), .B(n13604), .ZN(
        P1_U2945) );
  INV_X1 U16877 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n20057) );
  NAND2_X1 U16878 ( .A1(n20075), .A2(P1_LWORD_REG_8__SCAN_IN), .ZN(n13605) );
  OAI211_X1 U16879 ( .C1(n20057), .C2(n13631), .A(n13606), .B(n13605), .ZN(
        P1_U2960) );
  INV_X1 U16880 ( .A(n13607), .ZN(n13608) );
  AOI21_X1 U16881 ( .B1(n13610), .B2(n13609), .A(n13608), .ZN(n14660) );
  NAND2_X1 U16882 ( .A1(n14660), .A2(n20097), .ZN(n13616) );
  NAND2_X1 U16883 ( .A1(n13611), .A2(n14900), .ZN(n13614) );
  INV_X1 U16884 ( .A(n13612), .ZN(n13613) );
  AOI21_X1 U16885 ( .B1(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n13614), .A(
        n13613), .ZN(n13615) );
  OAI211_X1 U16886 ( .C1(n13617), .C2(n19949), .A(n13616), .B(n13615), .ZN(
        P1_U2999) );
  INV_X1 U16887 ( .A(n14660), .ZN(n13845) );
  NAND2_X1 U16888 ( .A1(n13618), .A2(n14519), .ZN(n13619) );
  INV_X2 U16889 ( .A(n20040), .ZN(n14815) );
  INV_X1 U16890 ( .A(n20160), .ZN(n20158) );
  NAND2_X1 U16891 ( .A1(n20158), .A2(DATAI_0_), .ZN(n13621) );
  NAND2_X1 U16892 ( .A1(n20160), .A2(BUF1_REG_0__SCAN_IN), .ZN(n13620) );
  AND2_X1 U16893 ( .A1(n13621), .A2(n13620), .ZN(n20162) );
  INV_X1 U16894 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n20074) );
  OAI222_X1 U16895 ( .A1(n13845), .A2(n14815), .B1(n14814), .B2(n20162), .C1(
        n20043), .C2(n20074), .ZN(P1_U2904) );
  INV_X1 U16896 ( .A(n13624), .ZN(n13626) );
  NAND2_X1 U16897 ( .A1(n13626), .A2(n13625), .ZN(n13627) );
  MUX2_X1 U16898 ( .A(n13629), .B(n13628), .S(n15212), .Z(n13630) );
  OAI21_X1 U16899 ( .B1(n19901), .B2(n15215), .A(n13630), .ZN(P2_U2885) );
  INV_X2 U16900 ( .A(n13631), .ZN(n20088) );
  AOI22_X1 U16901 ( .A1(n20088), .A2(P1_EAX_REG_2__SCAN_IN), .B1(
        P1_LWORD_REG_2__SCAN_IN), .B2(n13688), .ZN(n13635) );
  NAND2_X1 U16902 ( .A1(n20158), .A2(DATAI_2_), .ZN(n13633) );
  NAND2_X1 U16903 ( .A1(n20160), .A2(BUF1_REG_2__SCAN_IN), .ZN(n13632) );
  AND2_X1 U16904 ( .A1(n13633), .A2(n13632), .ZN(n20173) );
  INV_X1 U16905 ( .A(n20173), .ZN(n13634) );
  NAND2_X1 U16906 ( .A1(n20082), .A2(n13634), .ZN(n13646) );
  NAND2_X1 U16907 ( .A1(n13635), .A2(n13646), .ZN(P1_U2954) );
  AOI22_X1 U16908 ( .A1(n20088), .A2(P1_EAX_REG_10__SCAN_IN), .B1(
        P1_LWORD_REG_10__SCAN_IN), .B2(n13688), .ZN(n13638) );
  INV_X1 U16909 ( .A(DATAI_10_), .ZN(n13637) );
  NAND2_X1 U16910 ( .A1(n20160), .A2(BUF1_REG_10__SCAN_IN), .ZN(n13636) );
  OAI21_X1 U16911 ( .B1(n20160), .B2(n13637), .A(n13636), .ZN(n14762) );
  NAND2_X1 U16912 ( .A1(n20082), .A2(n14762), .ZN(n13677) );
  NAND2_X1 U16913 ( .A1(n13638), .A2(n13677), .ZN(P1_U2962) );
  AOI22_X1 U16914 ( .A1(n20088), .A2(P1_EAX_REG_6__SCAN_IN), .B1(
        P1_LWORD_REG_6__SCAN_IN), .B2(n13688), .ZN(n13642) );
  NAND2_X1 U16915 ( .A1(n20158), .A2(DATAI_6_), .ZN(n13640) );
  NAND2_X1 U16916 ( .A1(n20160), .A2(BUF1_REG_6__SCAN_IN), .ZN(n13639) );
  AND2_X1 U16917 ( .A1(n13640), .A2(n13639), .ZN(n20191) );
  INV_X1 U16918 ( .A(n20191), .ZN(n13641) );
  NAND2_X1 U16919 ( .A1(n20082), .A2(n13641), .ZN(n13666) );
  NAND2_X1 U16920 ( .A1(n13642), .A2(n13666), .ZN(P1_U2958) );
  AOI22_X1 U16921 ( .A1(n20088), .A2(P1_EAX_REG_19__SCAN_IN), .B1(
        P1_UWORD_REG_3__SCAN_IN), .B2(n13688), .ZN(n13645) );
  NAND2_X1 U16922 ( .A1(n20158), .A2(DATAI_3_), .ZN(n13644) );
  NAND2_X1 U16923 ( .A1(n20160), .A2(BUF1_REG_3__SCAN_IN), .ZN(n13643) );
  AND2_X1 U16924 ( .A1(n13644), .A2(n13643), .ZN(n20178) );
  INV_X1 U16925 ( .A(n20178), .ZN(n14787) );
  NAND2_X1 U16926 ( .A1(n20082), .A2(n14787), .ZN(n13689) );
  NAND2_X1 U16927 ( .A1(n13645), .A2(n13689), .ZN(P1_U2940) );
  AOI22_X1 U16928 ( .A1(n20088), .A2(P1_EAX_REG_18__SCAN_IN), .B1(
        P1_UWORD_REG_2__SCAN_IN), .B2(n13688), .ZN(n13647) );
  NAND2_X1 U16929 ( .A1(n13647), .A2(n13646), .ZN(P1_U2939) );
  AOI22_X1 U16930 ( .A1(n20088), .A2(P1_EAX_REG_17__SCAN_IN), .B1(
        P1_UWORD_REG_1__SCAN_IN), .B2(n13688), .ZN(n13650) );
  NAND2_X1 U16931 ( .A1(n20158), .A2(DATAI_1_), .ZN(n13649) );
  NAND2_X1 U16932 ( .A1(n20160), .A2(BUF1_REG_1__SCAN_IN), .ZN(n13648) );
  AND2_X1 U16933 ( .A1(n13649), .A2(n13648), .ZN(n20169) );
  INV_X1 U16934 ( .A(n20169), .ZN(n14797) );
  NAND2_X1 U16935 ( .A1(n20082), .A2(n14797), .ZN(n13675) );
  NAND2_X1 U16936 ( .A1(n13650), .A2(n13675), .ZN(P1_U2938) );
  AOI22_X1 U16937 ( .A1(n20088), .A2(P1_EAX_REG_16__SCAN_IN), .B1(
        P1_UWORD_REG_0__SCAN_IN), .B2(n13688), .ZN(n13652) );
  INV_X1 U16938 ( .A(n20162), .ZN(n13651) );
  NAND2_X1 U16939 ( .A1(n20082), .A2(n13651), .ZN(n13684) );
  NAND2_X1 U16940 ( .A1(n13652), .A2(n13684), .ZN(P1_U2937) );
  AOI22_X1 U16941 ( .A1(n20088), .A2(P1_EAX_REG_4__SCAN_IN), .B1(
        P1_LWORD_REG_4__SCAN_IN), .B2(n13688), .ZN(n13656) );
  NAND2_X1 U16942 ( .A1(n20158), .A2(DATAI_4_), .ZN(n13654) );
  NAND2_X1 U16943 ( .A1(n20160), .A2(BUF1_REG_4__SCAN_IN), .ZN(n13653) );
  AND2_X1 U16944 ( .A1(n13654), .A2(n13653), .ZN(n20184) );
  INV_X1 U16945 ( .A(n20184), .ZN(n13655) );
  NAND2_X1 U16946 ( .A1(n20082), .A2(n13655), .ZN(n13671) );
  NAND2_X1 U16947 ( .A1(n13656), .A2(n13671), .ZN(P1_U2956) );
  INV_X1 U16948 ( .A(n13657), .ZN(n13688) );
  AOI22_X1 U16949 ( .A1(n20088), .A2(P1_EAX_REG_27__SCAN_IN), .B1(
        P1_UWORD_REG_11__SCAN_IN), .B2(n13688), .ZN(n13660) );
  INV_X1 U16950 ( .A(DATAI_11_), .ZN(n13659) );
  NAND2_X1 U16951 ( .A1(n20160), .A2(BUF1_REG_11__SCAN_IN), .ZN(n13658) );
  OAI21_X1 U16952 ( .B1(n20160), .B2(n13659), .A(n13658), .ZN(n14759) );
  NAND2_X1 U16953 ( .A1(n20082), .A2(n14759), .ZN(n13686) );
  NAND2_X1 U16954 ( .A1(n13660), .A2(n13686), .ZN(P1_U2948) );
  AOI22_X1 U16955 ( .A1(n20088), .A2(P1_EAX_REG_5__SCAN_IN), .B1(
        P1_LWORD_REG_5__SCAN_IN), .B2(n13688), .ZN(n13663) );
  NAND2_X1 U16956 ( .A1(n20158), .A2(DATAI_5_), .ZN(n13662) );
  NAND2_X1 U16957 ( .A1(n20160), .A2(BUF1_REG_5__SCAN_IN), .ZN(n13661) );
  AND2_X1 U16958 ( .A1(n13662), .A2(n13661), .ZN(n20187) );
  INV_X1 U16959 ( .A(n20187), .ZN(n14780) );
  NAND2_X1 U16960 ( .A1(n20082), .A2(n14780), .ZN(n13664) );
  NAND2_X1 U16961 ( .A1(n13663), .A2(n13664), .ZN(P1_U2957) );
  AOI22_X1 U16962 ( .A1(n20088), .A2(P1_EAX_REG_21__SCAN_IN), .B1(
        P1_UWORD_REG_5__SCAN_IN), .B2(n13688), .ZN(n13665) );
  NAND2_X1 U16963 ( .A1(n13665), .A2(n13664), .ZN(P1_U2942) );
  AOI22_X1 U16964 ( .A1(n20088), .A2(P1_EAX_REG_22__SCAN_IN), .B1(
        P1_UWORD_REG_6__SCAN_IN), .B2(n13688), .ZN(n13667) );
  NAND2_X1 U16965 ( .A1(n13667), .A2(n13666), .ZN(P1_U2943) );
  AOI22_X1 U16966 ( .A1(n20088), .A2(P1_EAX_REG_13__SCAN_IN), .B1(
        P1_LWORD_REG_13__SCAN_IN), .B2(n13688), .ZN(n13670) );
  INV_X1 U16967 ( .A(DATAI_13_), .ZN(n13669) );
  NAND2_X1 U16968 ( .A1(n20160), .A2(BUF1_REG_13__SCAN_IN), .ZN(n13668) );
  OAI21_X1 U16969 ( .B1(n20160), .B2(n13669), .A(n13668), .ZN(n14812) );
  NAND2_X1 U16970 ( .A1(n20082), .A2(n14812), .ZN(n13673) );
  NAND2_X1 U16971 ( .A1(n13670), .A2(n13673), .ZN(P1_U2965) );
  AOI22_X1 U16972 ( .A1(n20088), .A2(P1_EAX_REG_20__SCAN_IN), .B1(
        P1_UWORD_REG_4__SCAN_IN), .B2(n13688), .ZN(n13672) );
  NAND2_X1 U16973 ( .A1(n13672), .A2(n13671), .ZN(P1_U2941) );
  AOI22_X1 U16974 ( .A1(n20088), .A2(P1_EAX_REG_29__SCAN_IN), .B1(
        P1_UWORD_REG_13__SCAN_IN), .B2(n13688), .ZN(n13674) );
  NAND2_X1 U16975 ( .A1(n13674), .A2(n13673), .ZN(P1_U2950) );
  AOI22_X1 U16976 ( .A1(n20088), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_LWORD_REG_1__SCAN_IN), .B2(n13688), .ZN(n13676) );
  NAND2_X1 U16977 ( .A1(n13676), .A2(n13675), .ZN(P1_U2953) );
  AOI22_X1 U16978 ( .A1(n20088), .A2(P1_EAX_REG_26__SCAN_IN), .B1(
        P1_UWORD_REG_10__SCAN_IN), .B2(n13688), .ZN(n13678) );
  NAND2_X1 U16979 ( .A1(n13678), .A2(n13677), .ZN(P1_U2947) );
  AOI22_X1 U16980 ( .A1(n20088), .A2(P1_EAX_REG_7__SCAN_IN), .B1(
        P1_LWORD_REG_7__SCAN_IN), .B2(n13688), .ZN(n13681) );
  NAND2_X1 U16981 ( .A1(n20158), .A2(DATAI_7_), .ZN(n13680) );
  NAND2_X1 U16982 ( .A1(n20160), .A2(BUF1_REG_7__SCAN_IN), .ZN(n13679) );
  AND2_X1 U16983 ( .A1(n13680), .A2(n13679), .ZN(n20199) );
  INV_X1 U16984 ( .A(n20199), .ZN(n14773) );
  NAND2_X1 U16985 ( .A1(n20082), .A2(n14773), .ZN(n13682) );
  NAND2_X1 U16986 ( .A1(n13681), .A2(n13682), .ZN(P1_U2959) );
  AOI22_X1 U16987 ( .A1(n20088), .A2(P1_EAX_REG_23__SCAN_IN), .B1(
        P1_UWORD_REG_7__SCAN_IN), .B2(n13688), .ZN(n13683) );
  NAND2_X1 U16988 ( .A1(n13683), .A2(n13682), .ZN(P1_U2944) );
  AOI22_X1 U16989 ( .A1(n20088), .A2(P1_EAX_REG_0__SCAN_IN), .B1(
        P1_LWORD_REG_0__SCAN_IN), .B2(n13688), .ZN(n13685) );
  NAND2_X1 U16990 ( .A1(n13685), .A2(n13684), .ZN(P1_U2952) );
  AOI22_X1 U16991 ( .A1(n20088), .A2(P1_EAX_REG_11__SCAN_IN), .B1(
        P1_LWORD_REG_11__SCAN_IN), .B2(n13688), .ZN(n13687) );
  NAND2_X1 U16992 ( .A1(n13687), .A2(n13686), .ZN(P1_U2963) );
  AOI22_X1 U16993 ( .A1(n20088), .A2(P1_EAX_REG_3__SCAN_IN), .B1(
        P1_LWORD_REG_3__SCAN_IN), .B2(n13688), .ZN(n13690) );
  NAND2_X1 U16994 ( .A1(n13690), .A2(n13689), .ZN(P1_U2955) );
  AOI22_X1 U16995 ( .A1(n13692), .A2(n19248), .B1(n16302), .B2(n13691), .ZN(
        n13696) );
  AOI21_X1 U16996 ( .B1(n19251), .B2(n13694), .A(n13693), .ZN(n13695) );
  OAI211_X1 U16997 ( .C1(n13691), .C2(n16310), .A(n13696), .B(n13695), .ZN(
        n13697) );
  AOI21_X1 U16998 ( .B1(n12673), .B2(n19250), .A(n13697), .ZN(n13698) );
  INV_X1 U16999 ( .A(n13698), .ZN(P2_U3013) );
  INV_X1 U17000 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n13701) );
  NOR2_X1 U17001 ( .A1(n20128), .A2(n13701), .ZN(n20141) );
  NOR2_X1 U17002 ( .A1(n20102), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13702) );
  AOI211_X1 U17003 ( .C1(n20091), .C2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n20141), .B(n13702), .ZN(n13706) );
  OR2_X1 U17004 ( .A1(n13703), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n20138) );
  NAND3_X1 U17005 ( .A1(n20138), .A2(n13704), .A3(n20098), .ZN(n13705) );
  OAI211_X1 U17006 ( .C1(n13958), .C2(n20159), .A(n13706), .B(n13705), .ZN(
        P1_U2998) );
  INV_X1 U17007 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n20070) );
  OAI222_X1 U17008 ( .A1(n13958), .A2(n14815), .B1(n14814), .B2(n20169), .C1(
        n20043), .C2(n20070), .ZN(P1_U2903) );
  NAND2_X1 U17009 ( .A1(n13709), .A2(n13708), .ZN(n13710) );
  NOR2_X1 U17010 ( .A1(n15892), .A2(n13710), .ZN(n13712) );
  NAND3_X1 U17011 ( .A1(n12536), .A2(n13712), .A3(n13711), .ZN(n13713) );
  NOR2_X1 U17012 ( .A1(n13714), .A2(n13713), .ZN(n15069) );
  NAND2_X1 U17013 ( .A1(n13715), .A2(n13726), .ZN(n13748) );
  XNOR2_X1 U17014 ( .A(n13716), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13724) );
  NOR2_X1 U17015 ( .A1(n13785), .A2(n10289), .ZN(n13717) );
  NOR2_X1 U17016 ( .A1(n13785), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n15071) );
  MUX2_X1 U17017 ( .A(n13717), .B(n15071), .S(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n13720) );
  INV_X1 U17018 ( .A(n15069), .ZN(n13753) );
  NOR3_X1 U17019 ( .A1(n13753), .A2(n13718), .A3(n13724), .ZN(n13719) );
  AOI211_X1 U17020 ( .C1(n13748), .C2(n13724), .A(n13720), .B(n13719), .ZN(
        n13721) );
  OAI21_X1 U17021 ( .B1(n13707), .B2(n15069), .A(n13721), .ZN(n13894) );
  INV_X1 U17022 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n13722) );
  AOI22_X1 U17023 ( .A1(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n20151), .B2(n13722), .ZN(
        n15074) );
  NOR2_X1 U17024 ( .A1(n13782), .A2(n20122), .ZN(n15076) );
  INV_X1 U17025 ( .A(n13724), .ZN(n13725) );
  AOI222_X1 U17026 ( .A1(n13894), .A2(n15073), .B1(n15074), .B2(n15076), .C1(
        n15078), .C2(n13725), .ZN(n13738) );
  INV_X1 U17027 ( .A(n13806), .ZN(n13735) );
  INV_X1 U17028 ( .A(n13727), .ZN(n20801) );
  NAND4_X1 U17029 ( .A1(n15901), .A2(n20801), .A3(n20810), .A4(n13728), .ZN(
        n13732) );
  NOR2_X1 U17030 ( .A1(n13961), .A2(n10415), .ZN(n13729) );
  NOR2_X1 U17031 ( .A1(n13730), .A2(n13729), .ZN(n13731) );
  NAND2_X1 U17032 ( .A1(n13732), .A2(n13731), .ZN(n13733) );
  INV_X1 U17033 ( .A(n13901), .ZN(n15870) );
  INV_X1 U17034 ( .A(n13736), .ZN(n19943) );
  NAND2_X1 U17035 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n16204), .ZN(n13908) );
  INV_X1 U17036 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n19950) );
  OAI22_X1 U17037 ( .A1(n15870), .A2(n19943), .B1(n13908), .B2(n19950), .ZN(
        n13760) );
  AOI21_X1 U17038 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n20806), .A(n13760), 
        .ZN(n13787) );
  NAND2_X1 U17039 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n13787), .ZN(
        n13737) );
  OAI21_X1 U17040 ( .B1(n13738), .B2(n13787), .A(n13737), .ZN(P1_U3472) );
  AOI21_X1 U17041 ( .B1(n13716), .B2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13739) );
  NOR2_X1 U17042 ( .A1(n10597), .A2(n13739), .ZN(n13754) );
  NAND3_X1 U17043 ( .A1(n15069), .A2(n13809), .A3(n13754), .ZN(n13751) );
  INV_X1 U17044 ( .A(n13743), .ZN(n13740) );
  MUX2_X1 U17045 ( .A(n13740), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n13716), .Z(n13742) );
  INV_X1 U17046 ( .A(n13744), .ZN(n13741) );
  NAND2_X1 U17047 ( .A1(n13742), .A2(n13741), .ZN(n13747) );
  AOI21_X1 U17048 ( .B1(n13744), .B2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n13743), .ZN(n13745) );
  NOR2_X1 U17049 ( .A1(n13785), .A2(n13745), .ZN(n13746) );
  AOI21_X1 U17050 ( .B1(n13748), .B2(n13747), .A(n13746), .ZN(n13750) );
  NAND2_X1 U17051 ( .A1(n15071), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13749) );
  NAND3_X1 U17052 ( .A1(n13751), .A2(n13750), .A3(n13749), .ZN(n13752) );
  INV_X1 U17053 ( .A(n13895), .ZN(n13755) );
  AOI22_X1 U17054 ( .A1(n13755), .A2(n15073), .B1(n13754), .B2(n15078), .ZN(
        n13757) );
  NAND2_X1 U17055 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n13787), .ZN(
        n13756) );
  OAI21_X1 U17056 ( .B1(n13757), .B2(n13787), .A(n13756), .ZN(P1_U3469) );
  INV_X1 U17057 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n13762) );
  INV_X1 U17058 ( .A(n13787), .ZN(n15081) );
  INV_X1 U17059 ( .A(n20292), .ZN(n20528) );
  OR2_X1 U17060 ( .A1(n13758), .A2(n20528), .ZN(n13759) );
  XNOR2_X1 U17061 ( .A(n13759), .B(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n20009) );
  NAND4_X1 U17062 ( .A1(n13760), .A2(n15073), .A3(n13899), .A4(n20009), .ZN(
        n13761) );
  OAI21_X1 U17063 ( .B1(n13762), .B2(n15081), .A(n13761), .ZN(P1_U3468) );
  OAI21_X1 U17064 ( .B1(n13765), .B2(n13764), .A(n13763), .ZN(n20032) );
  INV_X1 U17065 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n20068) );
  OAI222_X1 U17066 ( .A1(n20032), .A2(n14815), .B1(n14814), .B2(n20173), .C1(
        n20043), .C2(n20068), .ZN(P1_U2902) );
  XNOR2_X1 U17067 ( .A(n13766), .B(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13773) );
  NAND2_X1 U17068 ( .A1(n13768), .A2(n13769), .ZN(n13770) );
  AND2_X1 U17069 ( .A1(n13767), .A2(n13770), .ZN(n19082) );
  NOR2_X1 U17070 ( .A1(n15212), .A2(n19073), .ZN(n13771) );
  AOI21_X1 U17071 ( .B1(n19082), .B2(n15212), .A(n13771), .ZN(n13772) );
  OAI21_X1 U17072 ( .B1(n13773), .B2(n15215), .A(n13772), .ZN(P2_U2882) );
  INV_X1 U17073 ( .A(P1_REIP_REG_2__SCAN_IN), .ZN(n13774) );
  OAI22_X1 U17074 ( .A1(n14900), .A2(n13775), .B1(n20128), .B2(n13774), .ZN(
        n13776) );
  AOI21_X1 U17075 ( .B1(n20035), .B2(n16077), .A(n13776), .ZN(n13780) );
  OR2_X1 U17076 ( .A1(n13778), .A2(n13777), .ZN(n20127) );
  NAND3_X1 U17077 ( .A1(n20127), .A2(n20126), .A3(n20098), .ZN(n13779) );
  OAI211_X1 U17078 ( .C1(n20032), .C2(n20159), .A(n13780), .B(n13779), .ZN(
        P1_U2997) );
  INV_X1 U17079 ( .A(n10551), .ZN(n20784) );
  OAI22_X1 U17080 ( .A1(n20784), .A2(n15069), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n13781), .ZN(n15868) );
  INV_X1 U17081 ( .A(n15078), .ZN(n13783) );
  OAI22_X1 U17082 ( .A1(n13783), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n13782), .ZN(n13784) );
  AOI21_X1 U17083 ( .B1(n15073), .B2(n15868), .A(n13784), .ZN(n13788) );
  NOR2_X1 U17084 ( .A1(n13785), .A2(n9947), .ZN(n15867) );
  AOI22_X1 U17085 ( .A1(n15867), .A2(n15073), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n13787), .ZN(n13786) );
  OAI21_X1 U17086 ( .B1(n13788), .B2(n13787), .A(n13786), .ZN(P1_U3474) );
  INV_X1 U17087 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n13790) );
  AOI22_X1 U17088 ( .A1(P1_UWORD_REG_6__SCAN_IN), .A2(n20811), .B1(n20064), 
        .B2(P1_DATAO_REG_22__SCAN_IN), .ZN(n13789) );
  OAI21_X1 U17089 ( .B1(n13790), .B2(n13804), .A(n13789), .ZN(P1_U2914) );
  INV_X1 U17090 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n13792) );
  AOI22_X1 U17091 ( .A1(P1_UWORD_REG_0__SCAN_IN), .A2(n20811), .B1(n20064), 
        .B2(P1_DATAO_REG_16__SCAN_IN), .ZN(n13791) );
  OAI21_X1 U17092 ( .B1(n13792), .B2(n13804), .A(n13791), .ZN(P1_U2920) );
  INV_X1 U17093 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n13794) );
  AOI22_X1 U17094 ( .A1(P1_UWORD_REG_1__SCAN_IN), .A2(n20811), .B1(n20064), 
        .B2(P1_DATAO_REG_17__SCAN_IN), .ZN(n13793) );
  OAI21_X1 U17095 ( .B1(n13794), .B2(n13804), .A(n13793), .ZN(P1_U2919) );
  INV_X1 U17096 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n13796) );
  AOI22_X1 U17097 ( .A1(P1_UWORD_REG_2__SCAN_IN), .A2(n20811), .B1(n20064), 
        .B2(P1_DATAO_REG_18__SCAN_IN), .ZN(n13795) );
  OAI21_X1 U17098 ( .B1(n13796), .B2(n13804), .A(n13795), .ZN(P1_U2918) );
  INV_X1 U17099 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n13798) );
  AOI22_X1 U17100 ( .A1(P1_UWORD_REG_3__SCAN_IN), .A2(n20811), .B1(n20064), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n13797) );
  OAI21_X1 U17101 ( .B1(n13798), .B2(n13804), .A(n13797), .ZN(P1_U2917) );
  INV_X1 U17102 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n13800) );
  AOI22_X1 U17103 ( .A1(P1_UWORD_REG_7__SCAN_IN), .A2(n20811), .B1(n20064), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n13799) );
  OAI21_X1 U17104 ( .B1(n13800), .B2(n13804), .A(n13799), .ZN(P1_U2913) );
  INV_X1 U17105 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n13802) );
  AOI22_X1 U17106 ( .A1(P1_UWORD_REG_5__SCAN_IN), .A2(n20811), .B1(n20064), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n13801) );
  OAI21_X1 U17107 ( .B1(n13802), .B2(n13804), .A(n13801), .ZN(P1_U2915) );
  INV_X1 U17108 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n13805) );
  AOI22_X1 U17109 ( .A1(P1_UWORD_REG_4__SCAN_IN), .A2(n20811), .B1(n20064), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n13803) );
  OAI21_X1 U17110 ( .B1(n13805), .B2(n13804), .A(n13803), .ZN(P1_U2916) );
  INV_X1 U17111 ( .A(n13807), .ZN(n13810) );
  NAND4_X1 U17112 ( .A1(n13810), .A2(n10418), .A3(n13809), .A4(n13808), .ZN(
        n13811) );
  NAND2_X2 U17113 ( .A1(n14748), .A2(n20194), .ZN(n14749) );
  AND2_X1 U17114 ( .A1(n13814), .A2(n13813), .ZN(n13815) );
  OR2_X1 U17115 ( .A1(n9943), .A2(n13815), .ZN(n20129) );
  OAI22_X1 U17116 ( .A1(n14749), .A2(n20129), .B1(n13816), .B2(n14748), .ZN(
        n13817) );
  INV_X1 U17117 ( .A(n13817), .ZN(n13818) );
  OAI21_X1 U17118 ( .B1(n20032), .B2(n14747), .A(n13818), .ZN(P1_U2870) );
  INV_X2 U17119 ( .A(n14378), .ZN(n14747) );
  INV_X1 U17120 ( .A(n13819), .ZN(n13821) );
  NAND2_X1 U17121 ( .A1(n13821), .A2(n13820), .ZN(n13823) );
  AND2_X1 U17122 ( .A1(n13823), .A2(n13822), .ZN(n20144) );
  OAI22_X1 U17123 ( .A1(n14749), .A2(n20144), .B1(n13963), .B2(n14748), .ZN(
        n13824) );
  INV_X1 U17124 ( .A(n13824), .ZN(n13825) );
  OAI21_X1 U17125 ( .B1(n13958), .B2(n14747), .A(n13825), .ZN(P1_U2871) );
  INV_X1 U17126 ( .A(n13766), .ZN(n13847) );
  OAI21_X1 U17127 ( .B1(n13827), .B2(n13826), .A(n13847), .ZN(n19142) );
  NAND2_X1 U17128 ( .A1(n13829), .A2(n13828), .ZN(n13830) );
  AND2_X1 U17129 ( .A1(n13768), .A2(n13830), .ZN(n19249) );
  NOR2_X1 U17130 ( .A1(n15212), .A2(n13831), .ZN(n13832) );
  AOI21_X1 U17131 ( .B1(n19249), .B2(n15212), .A(n13832), .ZN(n13833) );
  OAI21_X1 U17132 ( .B1(n19142), .B2(n15215), .A(n13833), .ZN(P2_U2883) );
  NAND2_X1 U17133 ( .A1(n13835), .A2(n13834), .ZN(n13836) );
  INV_X1 U17134 ( .A(n15212), .ZN(n15192) );
  NOR2_X1 U17135 ( .A1(n13842), .A2(n15192), .ZN(n13843) );
  AOI21_X1 U17136 ( .B1(P2_EBX_REG_3__SCAN_IN), .B2(n15192), .A(n13843), .ZN(
        n13844) );
  OAI21_X1 U17137 ( .B1(n19539), .B2(n15215), .A(n13844), .ZN(P2_U2884) );
  OAI222_X1 U17138 ( .A1(n14655), .A2(n14749), .B1(n14748), .B2(n14656), .C1(
        n13845), .C2(n14747), .ZN(P1_U2872) );
  NOR2_X1 U17139 ( .A1(n13847), .A2(n13846), .ZN(n13849) );
  OAI211_X1 U17140 ( .C1(n13849), .C2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A(
        n15231), .B(n13848), .ZN(n13854) );
  AND2_X1 U17141 ( .A1(n13767), .A2(n13850), .ZN(n13852) );
  OR2_X1 U17142 ( .A1(n13852), .A2(n13851), .ZN(n19066) );
  INV_X1 U17143 ( .A(n19066), .ZN(n14342) );
  NAND2_X1 U17144 ( .A1(n14342), .A2(n15212), .ZN(n13853) );
  OAI211_X1 U17145 ( .C1(n15212), .C2(n11524), .A(n13854), .B(n13853), .ZN(
        P2_U2881) );
  XOR2_X1 U17146 ( .A(n13848), .B(P2_INSTQUEUE_REG_0__7__SCAN_IN), .Z(n13860)
         );
  INV_X1 U17147 ( .A(n13855), .ZN(n13856) );
  OAI21_X1 U17148 ( .B1(n13851), .B2(n13857), .A(n13856), .ZN(n19052) );
  MUX2_X1 U17149 ( .A(n13858), .B(n19052), .S(n15212), .Z(n13859) );
  OAI21_X1 U17150 ( .B1(n13860), .B2(n15215), .A(n13859), .ZN(P2_U2880) );
  NAND2_X1 U17151 ( .A1(n13862), .A2(n13861), .ZN(n13865) );
  INV_X1 U17152 ( .A(n13863), .ZN(n13864) );
  AND2_X1 U17153 ( .A1(n13865), .A2(n13864), .ZN(n14534) );
  XNOR2_X1 U17154 ( .A(n19901), .B(n14534), .ZN(n13870) );
  INV_X1 U17155 ( .A(n19906), .ZN(n13866) );
  NAND2_X1 U17156 ( .A1(n19910), .A2(n13866), .ZN(n13867) );
  OAI21_X1 U17157 ( .B1(n19910), .B2(n13866), .A(n13867), .ZN(n19158) );
  NOR2_X1 U17158 ( .A1(n14119), .A2(n16343), .ZN(n19159) );
  NOR2_X1 U17159 ( .A1(n19158), .A2(n19159), .ZN(n19157) );
  INV_X1 U17160 ( .A(n13867), .ZN(n13868) );
  NOR2_X1 U17161 ( .A1(n19157), .A2(n13868), .ZN(n13869) );
  NOR2_X1 U17162 ( .A1(n13869), .A2(n13870), .ZN(n14007) );
  AOI21_X1 U17163 ( .B1(n13870), .B2(n13869), .A(n14007), .ZN(n13873) );
  AOI22_X1 U17164 ( .A1(n19129), .A2(n16234), .B1(P2_EAX_REG_2__SCAN_IN), .B2(
        n19155), .ZN(n13872) );
  INV_X1 U17165 ( .A(n14534), .ZN(n19903) );
  NAND2_X1 U17166 ( .A1(n19903), .A2(n19156), .ZN(n13871) );
  OAI211_X1 U17167 ( .C1(n13873), .C2(n19160), .A(n13872), .B(n13871), .ZN(
        P2_U2917) );
  OAI21_X1 U17168 ( .B1(n13876), .B2(n13875), .A(n13874), .ZN(n13986) );
  INV_X1 U17169 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n20066) );
  OAI222_X1 U17170 ( .A1(n13986), .A2(n14815), .B1(n14814), .B2(n20178), .C1(
        n20043), .C2(n20066), .ZN(P1_U2901) );
  OR2_X1 U17171 ( .A1(n9943), .A2(n10265), .ZN(n13877) );
  NAND2_X1 U17172 ( .A1(n13945), .A2(n13877), .ZN(n20111) );
  INV_X1 U17173 ( .A(P1_EBX_REG_3__SCAN_IN), .ZN(n13974) );
  OAI222_X1 U17174 ( .A1(n20111), .A2(n14749), .B1(n13974), .B2(n14748), .C1(
        n14747), .C2(n13986), .ZN(P1_U2869) );
  OR2_X1 U17175 ( .A1(n13855), .A2(n13878), .ZN(n13880) );
  AND2_X1 U17176 ( .A1(n13880), .A2(n13879), .ZN(n16289) );
  INV_X1 U17177 ( .A(n16289), .ZN(n16325) );
  OAI211_X1 U17178 ( .C1(n13881), .C2(n13883), .A(n13882), .B(n15231), .ZN(
        n13885) );
  NAND2_X1 U17179 ( .A1(n15234), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n13884) );
  OAI211_X1 U17180 ( .C1(n16325), .C2(n15234), .A(n13885), .B(n13884), .ZN(
        P2_U2879) );
  XOR2_X1 U17181 ( .A(n13886), .B(n13874), .Z(n20096) );
  INV_X1 U17182 ( .A(n20096), .ZN(n13916) );
  XOR2_X1 U17183 ( .A(n13944), .B(n13945), .Z(n20104) );
  AOI22_X1 U17184 ( .A1(n14719), .A2(n20104), .B1(P1_EBX_REG_4__SCAN_IN), .B2(
        n14718), .ZN(n13887) );
  OAI21_X1 U17185 ( .B1(n13916), .B2(n14747), .A(n13887), .ZN(P1_U2868) );
  XOR2_X1 U17186 ( .A(n13882), .B(n13921), .Z(n13893) );
  NAND2_X1 U17187 ( .A1(n13888), .A2(n13879), .ZN(n13891) );
  INV_X1 U17188 ( .A(n13889), .ZN(n13890) );
  AND2_X1 U17189 ( .A1(n13891), .A2(n13890), .ZN(n16275) );
  INV_X1 U17190 ( .A(n16275), .ZN(n15709) );
  MUX2_X1 U17191 ( .A(n15709), .B(n12184), .S(n15234), .Z(n13892) );
  OAI21_X1 U17192 ( .B1(n13893), .B2(n15215), .A(n13892), .ZN(P2_U2878) );
  NOR2_X1 U17193 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(n13782), .ZN(n13903) );
  MUX2_X1 U17194 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n13894), .S(
        n13901), .Z(n15875) );
  AOI22_X1 U17195 ( .A1(n13903), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n15875), .B2(n13782), .ZN(n13898) );
  MUX2_X1 U17196 ( .A(n10581), .B(n13895), .S(n13901), .Z(n15877) );
  INV_X1 U17197 ( .A(n15877), .ZN(n13896) );
  AOI22_X1 U17198 ( .A1(n13903), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n13782), .B2(n13896), .ZN(n13897) );
  NOR2_X1 U17199 ( .A1(n13898), .A2(n13897), .ZN(n15878) );
  INV_X1 U17200 ( .A(n15878), .ZN(n13907) );
  NAND2_X1 U17201 ( .A1(n20009), .A2(n13899), .ZN(n13900) );
  NAND2_X1 U17202 ( .A1(n13900), .A2(n13901), .ZN(n13906) );
  OAI21_X1 U17203 ( .B1(n13901), .B2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(
        n13782), .ZN(n13902) );
  INV_X1 U17204 ( .A(n13902), .ZN(n13905) );
  AND2_X1 U17205 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n13903), .ZN(
        n13904) );
  AOI21_X1 U17206 ( .B1(n13906), .B2(n13905), .A(n13904), .ZN(n15887) );
  OAI21_X1 U17207 ( .B1(n13907), .B2(n10291), .A(n15887), .ZN(n15895) );
  NOR2_X1 U17208 ( .A1(n15895), .A2(P1_FLUSH_REG_SCAN_IN), .ZN(n13909) );
  NAND2_X1 U17209 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n20413), .ZN(n20773) );
  INV_X1 U17210 ( .A(n20773), .ZN(n20785) );
  OR2_X1 U17211 ( .A1(n9866), .A2(n20786), .ZN(n13912) );
  NOR2_X1 U17212 ( .A1(P1_STATEBS16_REG_SCAN_IN), .A2(n20786), .ZN(n20774) );
  INV_X1 U17213 ( .A(n20774), .ZN(n20526) );
  NAND2_X1 U17214 ( .A1(n13912), .A2(n20526), .ZN(n20262) );
  OAI21_X1 U17215 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n9866), .A(n20262), 
        .ZN(n13913) );
  OAI21_X1 U17216 ( .B1(n20529), .B2(n20785), .A(n13913), .ZN(n13914) );
  NAND2_X1 U17217 ( .A1(n20791), .A2(n13914), .ZN(n13915) );
  OAI21_X1 U17218 ( .B1(n20791), .B2(n20523), .A(n13915), .ZN(P1_U3477) );
  INV_X1 U17219 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n20063) );
  OAI222_X1 U17220 ( .A1(n14815), .A2(n13916), .B1(n14814), .B2(n20184), .C1(
        n20043), .C2(n20063), .ZN(P1_U2900) );
  NOR2_X1 U17221 ( .A1(n13707), .A2(n20785), .ZN(n13919) );
  AND2_X1 U17222 ( .A1(n9866), .A2(n20775), .ZN(n20382) );
  MUX2_X1 U17223 ( .A(n20262), .B(n20382), .S(n13917), .Z(n13918) );
  OAI21_X1 U17224 ( .B1(n13919), .B2(n13918), .A(n20791), .ZN(n13920) );
  OAI21_X1 U17225 ( .B1(n20791), .B2(n20461), .A(n13920), .ZN(P1_U3476) );
  INV_X1 U17226 ( .A(n13921), .ZN(n13923) );
  OAI21_X1 U17227 ( .B1(n13882), .B2(n13923), .A(n13922), .ZN(n13925) );
  NAND3_X1 U17228 ( .A1(n13925), .A2(n15231), .A3(n13924), .ZN(n13930) );
  NOR2_X1 U17229 ( .A1(n13927), .A2(n13889), .ZN(n13928) );
  NOR2_X1 U17230 ( .A1(n13926), .A2(n13928), .ZN(n19042) );
  NAND2_X1 U17231 ( .A1(n19042), .A2(n15212), .ZN(n13929) );
  OAI211_X1 U17232 ( .C1(n15212), .C2(n19034), .A(n13930), .B(n13929), .ZN(
        P2_U2877) );
  OAI21_X1 U17233 ( .B1(n13933), .B2(n13932), .A(n13931), .ZN(n13934) );
  INV_X1 U17234 ( .A(n13934), .ZN(n20115) );
  NAND2_X1 U17235 ( .A1(n20115), .A2(n20098), .ZN(n13938) );
  INV_X1 U17236 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n13935) );
  NOR2_X1 U17237 ( .A1(n20128), .A2(n13935), .ZN(n20112) );
  NOR2_X1 U17238 ( .A1(n20102), .A2(n13975), .ZN(n13936) );
  AOI211_X1 U17239 ( .C1(n20091), .C2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A(
        n20112), .B(n13936), .ZN(n13937) );
  OAI211_X1 U17240 ( .C1(n20159), .C2(n13986), .A(n13938), .B(n13937), .ZN(
        P1_U2996) );
  INV_X1 U17241 ( .A(n13939), .ZN(n13940) );
  AOI21_X1 U17242 ( .B1(n13942), .B2(n13941), .A(n13940), .ZN(n20004) );
  OAI21_X1 U17243 ( .B1(n13945), .B2(n13944), .A(n13943), .ZN(n13946) );
  AND2_X1 U17244 ( .A1(n13946), .A2(n13997), .ZN(n20000) );
  INV_X1 U17245 ( .A(n20000), .ZN(n16193) );
  OAI22_X1 U17246 ( .A1(n14749), .A2(n16193), .B1(n19998), .B2(n14748), .ZN(
        n13947) );
  AOI21_X1 U17247 ( .B1(n20004), .B2(n14378), .A(n13947), .ZN(n13948) );
  INV_X1 U17248 ( .A(n13948), .ZN(P1_U2867) );
  INV_X1 U17249 ( .A(n20004), .ZN(n13949) );
  OAI222_X1 U17250 ( .A1(n13949), .A2(n14815), .B1(n14814), .B2(n20187), .C1(
        n20043), .C2(n10638), .ZN(P1_U2899) );
  INV_X1 U17251 ( .A(n13924), .ZN(n13952) );
  OAI211_X1 U17252 ( .C1(n13952), .C2(n13951), .A(n10168), .B(n15231), .ZN(
        n13957) );
  INV_X1 U17253 ( .A(n13926), .ZN(n13954) );
  NAND2_X1 U17254 ( .A1(n13954), .A2(n10115), .ZN(n13955) );
  AND2_X1 U17255 ( .A1(n13955), .A2(n14016), .ZN(n16263) );
  NAND2_X1 U17256 ( .A1(n16263), .A2(n15212), .ZN(n13956) );
  OAI211_X1 U17257 ( .C1(n15212), .C2(n15144), .A(n13957), .B(n13956), .ZN(
        P2_U2876) );
  INV_X1 U17258 ( .A(n13958), .ZN(n13972) );
  NAND3_X1 U17259 ( .A1(n20022), .A2(P1_STATE2_REG_2__SCAN_IN), .A3(n13959), 
        .ZN(n13960) );
  NAND2_X1 U17260 ( .A1(n16023), .A2(n13960), .ZN(n20017) );
  INV_X1 U17261 ( .A(n20529), .ZN(n20591) );
  NOR2_X1 U17262 ( .A1(n13961), .A2(n20802), .ZN(n13962) );
  AND2_X1 U17263 ( .A1(n20022), .A2(n13962), .ZN(n20027) );
  AOI22_X1 U17264 ( .A1(n20591), .A2(n20027), .B1(n20026), .B2(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13970) );
  OAI22_X1 U17265 ( .A1(n20144), .A2(n20038), .B1(n13963), .B2(n19997), .ZN(
        n13964) );
  AOI21_X1 U17266 ( .B1(n19979), .B2(P1_REIP_REG_1__SCAN_IN), .A(n13964), .ZN(
        n13969) );
  OR2_X1 U17267 ( .A1(n20023), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n13968) );
  INV_X1 U17268 ( .A(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13966) );
  NAND2_X1 U17269 ( .A1(n20034), .A2(n13966), .ZN(n13967) );
  NAND4_X1 U17270 ( .A1(n13970), .A2(n13969), .A3(n13968), .A4(n13967), .ZN(
        n13971) );
  AOI21_X1 U17271 ( .B1(n13972), .B2(n20017), .A(n13971), .ZN(n13973) );
  INV_X1 U17272 ( .A(n13973), .ZN(P1_U2839) );
  INV_X1 U17273 ( .A(n20017), .ZN(n20031) );
  OAI22_X1 U17274 ( .A1(n20038), .A2(n20111), .B1(n19997), .B2(n13974), .ZN(
        n13981) );
  NAND3_X1 U17275 ( .A1(P1_REIP_REG_2__SCAN_IN), .A2(P1_REIP_REG_1__SCAN_IN), 
        .A3(n13935), .ZN(n13979) );
  NAND2_X1 U17276 ( .A1(n20026), .A2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13978) );
  INV_X1 U17277 ( .A(n13975), .ZN(n13976) );
  NAND2_X1 U17278 ( .A1(n20034), .A2(n13976), .ZN(n13977) );
  OAI211_X1 U17279 ( .C1(n20023), .C2(n13979), .A(n13978), .B(n13977), .ZN(
        n13980) );
  NOR2_X1 U17280 ( .A1(n13981), .A2(n13980), .ZN(n13985) );
  NOR2_X1 U17281 ( .A1(n13774), .A2(n13701), .ZN(n13982) );
  OAI21_X1 U17282 ( .B1(n20023), .B2(n13982), .A(n20022), .ZN(n13983) );
  OAI211_X1 U17283 ( .C1(n13986), .C2(n20031), .A(n13985), .B(n13984), .ZN(
        P1_U2837) );
  OR2_X1 U17284 ( .A1(n13989), .A2(n13988), .ZN(n13990) );
  AND2_X1 U17285 ( .A1(n13987), .A2(n13990), .ZN(n19982) );
  NOR2_X1 U17286 ( .A1(n13998), .A2(n13991), .ZN(n13992) );
  OR2_X1 U17287 ( .A1(n14076), .A2(n13992), .ZN(n16185) );
  OAI22_X1 U17288 ( .A1(n14749), .A2(n16185), .B1(n13993), .B2(n14748), .ZN(
        n13994) );
  AOI21_X1 U17289 ( .B1(n19982), .B2(n14378), .A(n13994), .ZN(n13995) );
  INV_X1 U17290 ( .A(n13995), .ZN(P1_U2865) );
  AND2_X1 U17291 ( .A1(n13997), .A2(n13996), .ZN(n13999) );
  OR2_X1 U17292 ( .A1(n13999), .A2(n13998), .ZN(n19988) );
  XOR2_X1 U17293 ( .A(n13939), .B(n14000), .Z(n19993) );
  INV_X1 U17294 ( .A(n19993), .ZN(n14013) );
  INV_X1 U17295 ( .A(P1_EBX_REG_6__SCAN_IN), .ZN(n14001) );
  OAI222_X1 U17296 ( .A1(n19988), .A2(n14749), .B1(n14747), .B2(n14013), .C1(
        n14001), .C2(n14748), .ZN(P1_U2866) );
  INV_X1 U17297 ( .A(n19982), .ZN(n14002) );
  INV_X1 U17298 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n20059) );
  OAI222_X1 U17299 ( .A1(n14002), .A2(n14815), .B1(n14814), .B2(n20199), .C1(
        n20043), .C2(n20059), .ZN(P1_U2897) );
  OR2_X1 U17300 ( .A1(n14004), .A2(n14003), .ZN(n14006) );
  NAND2_X1 U17301 ( .A1(n14006), .A2(n14005), .ZN(n14091) );
  AOI21_X1 U17302 ( .B1(n14534), .B2(n19901), .A(n14007), .ZN(n19150) );
  XNOR2_X1 U17303 ( .A(n19539), .B(n14091), .ZN(n19149) );
  NOR2_X1 U17304 ( .A1(n19150), .A2(n19149), .ZN(n19148) );
  AOI21_X1 U17305 ( .B1(n19539), .B2(n14091), .A(n19148), .ZN(n14009) );
  XNOR2_X1 U17306 ( .A(n14005), .B(n14008), .ZN(n14154) );
  NOR2_X1 U17307 ( .A1(n14009), .A2(n14154), .ZN(n19143) );
  XNOR2_X1 U17308 ( .A(n19143), .B(n19142), .ZN(n14012) );
  AOI22_X1 U17309 ( .A1(n19156), .A2(n14154), .B1(P2_EAX_REG_4__SCAN_IN), .B2(
        n19155), .ZN(n14011) );
  NAND2_X1 U17310 ( .A1(n19129), .A2(n19282), .ZN(n14010) );
  OAI211_X1 U17311 ( .C1(n14012), .C2(n19160), .A(n14011), .B(n14010), .ZN(
        P2_U2915) );
  INV_X1 U17312 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n14014) );
  OAI222_X1 U17313 ( .A1(n20043), .A2(n14014), .B1(n14814), .B2(n20191), .C1(
        n14815), .C2(n14013), .ZN(P1_U2898) );
  AND2_X1 U17314 ( .A1(n14016), .A2(n14015), .ZN(n14018) );
  OR2_X1 U17315 ( .A1(n14018), .A2(n14017), .ZN(n16252) );
  OAI211_X1 U17316 ( .C1(n13950), .C2(n14020), .A(n10167), .B(n15231), .ZN(
        n14022) );
  NAND2_X1 U17317 ( .A1(n15234), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n14021) );
  OAI211_X1 U17318 ( .C1(n16252), .C2(n15234), .A(n14022), .B(n14021), .ZN(
        P2_U2875) );
  NOR2_X2 U17319 ( .A1(n19689), .A2(n19658), .ZN(n19684) );
  NOR2_X2 U17320 ( .A1(n19659), .A2(n19889), .ZN(n19654) );
  OAI21_X1 U17321 ( .B1(n19684), .B2(n19654), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n14028) );
  INV_X1 U17322 ( .A(n14024), .ZN(n19385) );
  INV_X1 U17323 ( .A(n19575), .ZN(n19450) );
  NAND3_X1 U17324 ( .A1(n19385), .A2(n19450), .A3(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n14027) );
  AOI21_X1 U17325 ( .B1(n12071), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n14025) );
  NAND3_X1 U17326 ( .A1(n19914), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19666) );
  NOR2_X1 U17327 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19666), .ZN(
        n19652) );
  NOR2_X1 U17328 ( .A1(n14025), .A2(n19652), .ZN(n14026) );
  AOI22_X1 U17329 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n19295), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n19294), .ZN(n19623) );
  AOI22_X2 U17330 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n19295), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n19294), .ZN(n19770) );
  INV_X1 U17331 ( .A(n19770), .ZN(n19620) );
  AOI22_X1 U17332 ( .A1(n19654), .A2(n19767), .B1(n19684), .B2(n19620), .ZN(
        n14037) );
  OAI21_X1 U17333 ( .B1(n14031), .B2(n19652), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n14034) );
  NAND3_X1 U17334 ( .A1(n14032), .A2(n19450), .A3(n19385), .ZN(n14033) );
  NAND2_X1 U17335 ( .A1(n14034), .A2(n14033), .ZN(n19653) );
  NOR2_X2 U17336 ( .A1(n19154), .A2(n19389), .ZN(n19766) );
  NAND2_X1 U17337 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19747), .ZN(n19270) );
  AND2_X1 U17338 ( .A1(n14035), .A2(n19296), .ZN(n19765) );
  AOI22_X1 U17339 ( .A1(n19653), .A2(n19766), .B1(n19765), .B2(n19652), .ZN(
        n14036) );
  OAI211_X1 U17340 ( .C1(n19657), .C2(n14038), .A(n14037), .B(n14036), .ZN(
        P2_U3147) );
  XOR2_X1 U17341 ( .A(n14039), .B(n14040), .Z(n15716) );
  INV_X1 U17342 ( .A(n15716), .ZN(n19134) );
  NAND2_X1 U17343 ( .A1(n19079), .A2(n14041), .ZN(n14042) );
  XNOR2_X1 U17344 ( .A(n16271), .B(n14042), .ZN(n14043) );
  NAND2_X1 U17345 ( .A1(n14043), .A2(n9868), .ZN(n14049) );
  AOI22_X1 U17346 ( .A1(n14044), .A2(n19049), .B1(n19101), .B2(
        P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n14045) );
  OAI211_X1 U17347 ( .C1(n12184), .C2(n19072), .A(n14045), .B(n15684), .ZN(
        n14047) );
  NOR2_X1 U17348 ( .A1(n15709), .A2(n19067), .ZN(n14046) );
  AOI211_X1 U17349 ( .C1(P2_REIP_REG_9__SCAN_IN), .C2(n19091), .A(n14047), .B(
        n14046), .ZN(n14048) );
  OAI211_X1 U17350 ( .C1(n19134), .C2(n19087), .A(n14049), .B(n14048), .ZN(
        P2_U2846) );
  NAND2_X1 U17351 ( .A1(n19079), .A2(n14050), .ZN(n14051) );
  XNOR2_X1 U17352 ( .A(n16301), .B(n14051), .ZN(n14052) );
  NAND2_X1 U17353 ( .A1(n14052), .A2(n9868), .ZN(n14061) );
  OAI22_X1 U17354 ( .A1(n14054), .A2(n19072), .B1(n11812), .B2(n19074), .ZN(
        n14055) );
  AOI21_X1 U17355 ( .B1(n19101), .B2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A(
        n14055), .ZN(n14056) );
  OAI21_X1 U17356 ( .B1(n14057), .B2(n19095), .A(n14056), .ZN(n14059) );
  NOR2_X1 U17357 ( .A1(n14091), .A2(n19087), .ZN(n14058) );
  AOI211_X1 U17358 ( .C1(n19097), .C2(n14053), .A(n14059), .B(n14058), .ZN(
        n14060) );
  OAI211_X1 U17359 ( .C1(n19539), .C2(n14363), .A(n14061), .B(n14060), .ZN(
        P2_U2852) );
  INV_X1 U17360 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n14070) );
  INV_X1 U17361 ( .A(n14062), .ZN(n14063) );
  OAI211_X1 U17362 ( .C1(n14019), .C2(n14064), .A(n14063), .B(n15231), .ZN(
        n14069) );
  OAI21_X1 U17363 ( .B1(n14017), .B2(n14066), .A(n14065), .ZN(n19029) );
  INV_X1 U17364 ( .A(n19029), .ZN(n14067) );
  NAND2_X1 U17365 ( .A1(n14067), .A2(n15212), .ZN(n14068) );
  OAI211_X1 U17366 ( .C1(n15212), .C2(n14070), .A(n14069), .B(n14068), .ZN(
        P2_U2874) );
  AOI21_X1 U17367 ( .B1(n14073), .B2(n13987), .A(n14072), .ZN(n14252) );
  INV_X1 U17368 ( .A(n14252), .ZN(n14106) );
  INV_X1 U17369 ( .A(n14814), .ZN(n20039) );
  AOI22_X1 U17370 ( .A1(n20039), .A2(n14770), .B1(P1_EAX_REG_8__SCAN_IN), .B2(
        n14816), .ZN(n14074) );
  OAI21_X1 U17371 ( .B1(n14106), .B2(n14815), .A(n14074), .ZN(P1_U2896) );
  INV_X1 U17372 ( .A(n14250), .ZN(n14083) );
  OR2_X1 U17373 ( .A1(n14076), .A2(n14075), .ZN(n14077) );
  NAND2_X1 U17374 ( .A1(n14204), .A2(n14077), .ZN(n16178) );
  INV_X1 U17375 ( .A(P1_REIP_REG_8__SCAN_IN), .ZN(n20721) );
  NAND4_X1 U17376 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(P1_REIP_REG_6__SCAN_IN), 
        .A3(P1_REIP_REG_5__SCAN_IN), .A4(n20721), .ZN(n14078) );
  OAI22_X1 U17377 ( .A1(n20038), .A2(n16178), .B1(n19999), .B2(n14078), .ZN(
        n14082) );
  OR2_X1 U17378 ( .A1(n14611), .A2(n16020), .ZN(n15960) );
  INV_X1 U17379 ( .A(n15960), .ZN(n19969) );
  AOI22_X1 U17380 ( .A1(P1_EBX_REG_8__SCAN_IN), .A2(n20025), .B1(
        P1_REIP_REG_8__SCAN_IN), .B2(n19969), .ZN(n14079) );
  NAND2_X1 U17381 ( .A1(n14547), .A2(n20022), .ZN(n20011) );
  OAI211_X1 U17382 ( .C1(n20014), .C2(n14080), .A(n14079), .B(n20011), .ZN(
        n14081) );
  AOI211_X1 U17383 ( .C1(n20034), .C2(n14083), .A(n14082), .B(n14081), .ZN(
        n14084) );
  OAI21_X1 U17384 ( .B1(n16023), .B2(n14106), .A(n14084), .ZN(P1_U2832) );
  INV_X1 U17385 ( .A(n14085), .ZN(n14090) );
  AOI21_X1 U17386 ( .B1(n14089), .B2(n14086), .A(n14087), .ZN(n14088) );
  AOI21_X1 U17387 ( .B1(n14090), .B2(n14089), .A(n14088), .ZN(n16307) );
  INV_X1 U17388 ( .A(n16307), .ZN(n14105) );
  INV_X1 U17389 ( .A(n14091), .ZN(n19892) );
  AOI21_X1 U17390 ( .B1(n15610), .B2(n14093), .A(n14092), .ZN(n14110) );
  INV_X1 U17391 ( .A(n14110), .ZN(n14097) );
  NOR2_X1 U17392 ( .A1(n16351), .A2(n14094), .ZN(n14096) );
  MUX2_X1 U17393 ( .A(n14097), .B(n14096), .S(n14095), .Z(n14099) );
  OAI22_X1 U17394 ( .A1(n13842), .A2(n16326), .B1(n11812), .B2(n12458), .ZN(
        n14098) );
  AOI211_X1 U17395 ( .C1(n19892), .C2(n16344), .A(n14099), .B(n14098), .ZN(
        n14104) );
  OR2_X1 U17396 ( .A1(n14101), .A2(n14100), .ZN(n16303) );
  NAND3_X1 U17397 ( .A1(n16303), .A2(n16342), .A3(n14102), .ZN(n14103) );
  OAI211_X1 U17398 ( .C1(n14105), .C2(n16321), .A(n14104), .B(n14103), .ZN(
        P2_U3043) );
  INV_X1 U17399 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n21061) );
  OAI222_X1 U17400 ( .A1(n16178), .A2(n14749), .B1(n14748), .B2(n21061), .C1(
        n14747), .C2(n14106), .ZN(P1_U2864) );
  XNOR2_X1 U17401 ( .A(n14107), .B(n21161), .ZN(n19252) );
  INV_X1 U17402 ( .A(n19252), .ZN(n14118) );
  XOR2_X1 U17403 ( .A(n14109), .B(n14108), .Z(n19247) );
  NAND2_X1 U17404 ( .A1(n19247), .A2(n16338), .ZN(n14117) );
  OAI21_X1 U17405 ( .B1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n16351), .A(
        n14110), .ZN(n14338) );
  NOR2_X1 U17406 ( .A1(n11816), .A2(n15684), .ZN(n14111) );
  AOI21_X1 U17407 ( .B1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n14338), .A(
        n14111), .ZN(n14113) );
  NAND2_X1 U17408 ( .A1(n16344), .A2(n14154), .ZN(n14112) );
  OAI211_X1 U17409 ( .C1(n14114), .C2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A(
        n14113), .B(n14112), .ZN(n14115) );
  AOI21_X1 U17410 ( .B1(n19249), .B2(n16340), .A(n14115), .ZN(n14116) );
  OAI211_X1 U17411 ( .C1(n14118), .C2(n16327), .A(n14117), .B(n14116), .ZN(
        P2_U3042) );
  INV_X1 U17412 ( .A(n19349), .ZN(n14120) );
  NAND2_X1 U17413 ( .A1(n19373), .A2(n14120), .ZN(n14121) );
  NAND2_X1 U17414 ( .A1(n14121), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n14123) );
  NOR2_X1 U17415 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19354) );
  NAND2_X1 U17416 ( .A1(n19575), .A2(n19354), .ZN(n14122) );
  NAND2_X1 U17417 ( .A1(n14123), .A2(n14122), .ZN(n14128) );
  NAND2_X1 U17418 ( .A1(n14124), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n14125) );
  NAND2_X1 U17419 ( .A1(n14125), .A2(n19917), .ZN(n14126) );
  INV_X1 U17420 ( .A(n19354), .ZN(n19305) );
  NOR2_X1 U17421 ( .A1(n19572), .A2(n19305), .ZN(n19347) );
  INV_X1 U17422 ( .A(n19347), .ZN(n14134) );
  AOI21_X1 U17423 ( .B1(n14126), .B2(n14134), .A(n19389), .ZN(n14127) );
  INV_X1 U17424 ( .A(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n14137) );
  INV_X1 U17425 ( .A(n14129), .ZN(n19446) );
  OAI21_X1 U17426 ( .B1(n14130), .B2(n19347), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n14131) );
  OAI21_X1 U17427 ( .B1(n19305), .B2(n19446), .A(n14131), .ZN(n19348) );
  INV_X1 U17428 ( .A(n19107), .ZN(n14132) );
  NOR2_X2 U17429 ( .A1(n14132), .A2(n19389), .ZN(n19741) );
  NAND2_X1 U17430 ( .A1(n16370), .A2(n19296), .ZN(n19257) );
  AOI22_X1 U17431 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n19295), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n19294), .ZN(n19703) );
  AOI22_X1 U17432 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n19295), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n19294), .ZN(n19752) );
  INV_X1 U17433 ( .A(n19752), .ZN(n19690) );
  AOI22_X1 U17434 ( .A1(n19349), .A2(n19749), .B1(n19379), .B2(n19690), .ZN(
        n14133) );
  OAI21_X1 U17435 ( .B1(n19257), .B2(n14134), .A(n14133), .ZN(n14135) );
  AOI21_X1 U17436 ( .B1(n19348), .B2(n19741), .A(n14135), .ZN(n14136) );
  OAI21_X1 U17437 ( .B1(n19338), .B2(n14137), .A(n14136), .ZN(P2_U3064) );
  INV_X1 U17438 ( .A(n14138), .ZN(n14139) );
  OAI211_X1 U17439 ( .C1(n14062), .C2(n14140), .A(n15231), .B(n14139), .ZN(
        n14145) );
  NAND2_X1 U17440 ( .A1(n14065), .A2(n14142), .ZN(n14143) );
  AND2_X1 U17441 ( .A1(n14141), .A2(n14143), .ZN(n19020) );
  NAND2_X1 U17442 ( .A1(n19020), .A2(n15212), .ZN(n14144) );
  OAI211_X1 U17443 ( .C1(n15212), .C2(n14146), .A(n14145), .B(n14144), .ZN(
        P2_U2873) );
  INV_X1 U17444 ( .A(n19255), .ZN(n14150) );
  NOR2_X1 U17445 ( .A1(n10053), .A2(n14147), .ZN(n14149) );
  AOI21_X1 U17446 ( .B1(n14150), .B2(n14149), .A(n19809), .ZN(n14148) );
  OAI21_X1 U17447 ( .B1(n14150), .B2(n14149), .A(n14148), .ZN(n14159) );
  NOR2_X1 U17448 ( .A1(n19074), .A2(n11816), .ZN(n14151) );
  AOI211_X1 U17449 ( .C1(n19090), .C2(P2_EBX_REG_4__SCAN_IN), .A(n19245), .B(
        n14151), .ZN(n14152) );
  OAI21_X1 U17450 ( .B1(n10045), .B2(n19057), .A(n14152), .ZN(n14153) );
  AOI21_X1 U17451 ( .B1(n19088), .B2(n14154), .A(n14153), .ZN(n14155) );
  OAI21_X1 U17452 ( .B1(n14156), .B2(n19095), .A(n14155), .ZN(n14157) );
  AOI21_X1 U17453 ( .B1(n19249), .B2(n19097), .A(n14157), .ZN(n14158) );
  OAI211_X1 U17454 ( .C1(n19142), .C2(n14363), .A(n14159), .B(n14158), .ZN(
        P2_U2851) );
  NAND2_X1 U17455 ( .A1(n14161), .A2(n14160), .ZN(n14162) );
  XNOR2_X1 U17456 ( .A(n14163), .B(n14162), .ZN(n16095) );
  NAND2_X1 U17457 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n14288) );
  NAND2_X1 U17458 ( .A1(n14167), .A2(n20122), .ZN(n20139) );
  INV_X1 U17459 ( .A(n20139), .ZN(n14168) );
  OR2_X1 U17460 ( .A1(n14165), .A2(n14164), .ZN(n14166) );
  NOR2_X1 U17461 ( .A1(n14288), .A2(n20120), .ZN(n14173) );
  INV_X1 U17462 ( .A(n14173), .ZN(n14172) );
  NAND2_X1 U17463 ( .A1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n20106) );
  NOR2_X1 U17464 ( .A1(n20106), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n16195) );
  INV_X1 U17465 ( .A(n16195), .ZN(n14171) );
  INV_X1 U17466 ( .A(n15054), .ZN(n20125) );
  OR2_X1 U17467 ( .A1(n14288), .A2(n20106), .ZN(n14477) );
  NOR2_X1 U17468 ( .A1(n16199), .A2(n20106), .ZN(n14286) );
  OAI21_X1 U17469 ( .B1(n20122), .B2(n20151), .A(n20135), .ZN(n14289) );
  NAND2_X1 U17470 ( .A1(n14170), .A2(n14169), .ZN(n20123) );
  INV_X1 U17471 ( .A(n20123), .ZN(n20150) );
  OAI221_X1 U17472 ( .B1(n20121), .B2(n14286), .C1(n20121), .C2(n14289), .A(
        n20150), .ZN(n16156) );
  AOI21_X1 U17473 ( .B1(n20125), .B2(n14477), .A(n16156), .ZN(n16200) );
  OAI21_X1 U17474 ( .B1(n14172), .B2(n14171), .A(n16200), .ZN(n16175) );
  NOR2_X1 U17475 ( .A1(n15051), .A2(n14173), .ZN(n16168) );
  INV_X1 U17476 ( .A(n16168), .ZN(n14174) );
  NAND2_X1 U17477 ( .A1(n14289), .A2(n14174), .ZN(n20119) );
  NAND2_X1 U17478 ( .A1(n14286), .A2(n20107), .ZN(n16180) );
  INV_X1 U17479 ( .A(n16180), .ZN(n14175) );
  INV_X1 U17480 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n16181) );
  AOI22_X1 U17481 ( .A1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n16175), .B1(
        n14175), .B2(n16181), .ZN(n14177) );
  NAND2_X1 U17482 ( .A1(n20103), .A2(P1_REIP_REG_6__SCAN_IN), .ZN(n14176) );
  OAI211_X1 U17483 ( .C1(n20145), .C2(n19988), .A(n14177), .B(n14176), .ZN(
        n14178) );
  AOI21_X1 U17484 ( .B1(n20137), .B2(n16095), .A(n14178), .ZN(n14179) );
  INV_X1 U17485 ( .A(n14179), .ZN(P1_U3025) );
  NOR2_X1 U17486 ( .A1(n10053), .A2(n14180), .ZN(n14181) );
  XNOR2_X1 U17487 ( .A(n14181), .B(n16292), .ZN(n14182) );
  NAND2_X1 U17488 ( .A1(n14182), .A2(n9868), .ZN(n14198) );
  INV_X1 U17489 ( .A(n14183), .ZN(n14196) );
  NAND2_X1 U17490 ( .A1(n19101), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n14194) );
  INV_X1 U17491 ( .A(n14184), .ZN(n14185) );
  OR2_X1 U17492 ( .A1(n14186), .A2(n14185), .ZN(n14188) );
  INV_X1 U17493 ( .A(n14039), .ZN(n14187) );
  NAND2_X1 U17494 ( .A1(n19088), .A2(n19135), .ZN(n14189) );
  OAI21_X1 U17495 ( .B1(n19074), .B2(n14190), .A(n14189), .ZN(n14191) );
  INV_X1 U17496 ( .A(n14191), .ZN(n14193) );
  AOI21_X1 U17497 ( .B1(n19090), .B2(P2_EBX_REG_8__SCAN_IN), .A(n19038), .ZN(
        n14192) );
  NAND3_X1 U17498 ( .A1(n14194), .A2(n14193), .A3(n14192), .ZN(n14195) );
  AOI21_X1 U17499 ( .B1(n14196), .B2(n19049), .A(n14195), .ZN(n14197) );
  OAI211_X1 U17500 ( .C1(n16325), .C2(n19067), .A(n14198), .B(n14197), .ZN(
        P2_U2847) );
  INV_X1 U17501 ( .A(n14199), .ZN(n14200) );
  AND2_X1 U17502 ( .A1(n14202), .A2(n14201), .ZN(n14203) );
  NOR2_X1 U17503 ( .A1(n14200), .A2(n14203), .ZN(n20041) );
  INV_X1 U17504 ( .A(n20041), .ZN(n14207) );
  AOI21_X1 U17505 ( .B1(n14205), .B2(n14204), .A(n9957), .ZN(n19965) );
  AOI22_X1 U17506 ( .A1(n19965), .A2(n14719), .B1(n14718), .B2(
        P1_EBX_REG_9__SCAN_IN), .ZN(n14206) );
  OAI21_X1 U17507 ( .B1(n14207), .B2(n14747), .A(n14206), .ZN(P1_U2863) );
  OAI211_X1 U17508 ( .C1(n14138), .C2(n14209), .A(n15231), .B(n14208), .ZN(
        n14214) );
  NAND2_X1 U17509 ( .A1(n14141), .A2(n14210), .ZN(n14211) );
  NAND2_X1 U17510 ( .A1(n14353), .A2(n14211), .ZN(n19005) );
  INV_X1 U17511 ( .A(n19005), .ZN(n14212) );
  NAND2_X1 U17512 ( .A1(n14212), .A2(n15212), .ZN(n14213) );
  OAI211_X1 U17513 ( .C1(n15212), .C2(n12216), .A(n14214), .B(n14213), .ZN(
        P2_U2872) );
  XNOR2_X1 U17514 ( .A(n14215), .B(n14216), .ZN(n16294) );
  OAI21_X1 U17515 ( .B1(n10249), .B2(n14218), .A(n14217), .ZN(n14219) );
  OAI21_X1 U17516 ( .B1(n14220), .B2(n10249), .A(n14219), .ZN(n16296) );
  INV_X1 U17517 ( .A(n16296), .ZN(n14232) );
  OAI21_X1 U17518 ( .B1(n14223), .B2(n14222), .A(n14221), .ZN(n19146) );
  INV_X1 U17519 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n19836) );
  NOR2_X1 U17520 ( .A1(n19836), .A2(n15684), .ZN(n14228) );
  INV_X1 U17521 ( .A(n14224), .ZN(n14335) );
  NAND2_X1 U17522 ( .A1(n15613), .A2(n14339), .ZN(n14225) );
  AOI211_X1 U17523 ( .C1(n14226), .C2(n21161), .A(n14335), .B(n14225), .ZN(
        n14227) );
  AOI211_X1 U17524 ( .C1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .C2(n14338), .A(
        n14228), .B(n14227), .ZN(n14230) );
  NAND2_X1 U17525 ( .A1(n19082), .A2(n16340), .ZN(n14229) );
  OAI211_X1 U17526 ( .C1(n19146), .C2(n16313), .A(n14230), .B(n14229), .ZN(
        n14231) );
  AOI21_X1 U17527 ( .B1(n14232), .B2(n16342), .A(n14231), .ZN(n14233) );
  OAI21_X1 U17528 ( .B1(n16321), .B2(n16294), .A(n14233), .ZN(P2_U3041) );
  INV_X1 U17529 ( .A(n14236), .ZN(n14539) );
  INV_X1 U17530 ( .A(n14356), .ZN(n14235) );
  AOI221_X1 U17531 ( .B1(n14539), .B2(n14356), .C1(n14236), .C2(n14235), .A(
        n19809), .ZN(n14237) );
  INV_X1 U17532 ( .A(n14237), .ZN(n14245) );
  AOI22_X1 U17533 ( .A1(P2_EBX_REG_2__SCAN_IN), .A2(n19090), .B1(
        P2_REIP_REG_2__SCAN_IN), .B2(n19091), .ZN(n14239) );
  NAND2_X1 U17534 ( .A1(n19101), .A2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n14238) );
  OAI211_X1 U17535 ( .C1(n19095), .C2(n14240), .A(n14239), .B(n14238), .ZN(
        n14242) );
  NOR2_X1 U17536 ( .A1(n14534), .A2(n19087), .ZN(n14241) );
  AOI211_X1 U17537 ( .C1(n19097), .C2(n14243), .A(n14242), .B(n14241), .ZN(
        n14244) );
  OAI211_X1 U17538 ( .C1(n19901), .C2(n14363), .A(n14245), .B(n14244), .ZN(
        P2_U2853) );
  XOR2_X1 U17539 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B(n14247), .Z(
        n14248) );
  XNOR2_X1 U17540 ( .A(n14246), .B(n14248), .ZN(n16176) );
  AOI22_X1 U17541 ( .A1(n20091), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B1(
        n20103), .B2(P1_REIP_REG_8__SCAN_IN), .ZN(n14249) );
  OAI21_X1 U17542 ( .B1(n20102), .B2(n14250), .A(n14249), .ZN(n14251) );
  AOI21_X1 U17543 ( .B1(n14252), .B2(n20097), .A(n14251), .ZN(n14253) );
  OAI21_X1 U17544 ( .B1(n16176), .B2(n19949), .A(n14253), .ZN(P1_U2991) );
  AOI21_X1 U17545 ( .B1(n10281), .B2(n14199), .A(n14255), .ZN(n16035) );
  AND2_X1 U17546 ( .A1(n14257), .A2(n14256), .ZN(n14258) );
  OR2_X1 U17547 ( .A1(n14305), .A2(n14258), .ZN(n16028) );
  OAI22_X1 U17548 ( .A1(n16028), .A2(n14749), .B1(n16029), .B2(n14748), .ZN(
        n14259) );
  AOI21_X1 U17549 ( .B1(n16035), .B2(n14378), .A(n14259), .ZN(n14260) );
  INV_X1 U17550 ( .A(n14260), .ZN(P1_U2862) );
  NOR3_X1 U17551 ( .A1(n10053), .A2(n14262), .A3(n19809), .ZN(n15143) );
  INV_X1 U17552 ( .A(n16258), .ZN(n14261) );
  OAI211_X1 U17553 ( .C1(n10053), .C2(n14262), .A(n9868), .B(n14261), .ZN(
        n14274) );
  INV_X1 U17554 ( .A(n14263), .ZN(n14264) );
  OR2_X1 U17555 ( .A1(n14265), .A2(n14264), .ZN(n14268) );
  INV_X1 U17556 ( .A(n14266), .ZN(n14267) );
  AND2_X1 U17557 ( .A1(n14268), .A2(n14267), .ZN(n15667) );
  AOI22_X1 U17558 ( .A1(n19091), .A2(P2_REIP_REG_12__SCAN_IN), .B1(n19088), 
        .B2(n15667), .ZN(n14269) );
  OAI211_X1 U17559 ( .C1(n14270), .C2(n19072), .A(n14269), .B(n15684), .ZN(
        n14272) );
  NOR2_X1 U17560 ( .A1(n16252), .A2(n19067), .ZN(n14271) );
  AOI211_X1 U17561 ( .C1(n19101), .C2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n14272), .B(n14271), .ZN(n14273) );
  OAI211_X1 U17562 ( .C1(n14275), .C2(n19095), .A(n14274), .B(n14273), .ZN(
        n14276) );
  AOI21_X1 U17563 ( .B1(n15143), .B2(n16258), .A(n14276), .ZN(n14277) );
  INV_X1 U17564 ( .A(n14277), .ZN(P2_U2843) );
  INV_X1 U17565 ( .A(n16035), .ZN(n14279) );
  INV_X1 U17566 ( .A(n14762), .ZN(n14278) );
  INV_X1 U17567 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n21136) );
  OAI222_X1 U17568 ( .A1(n14815), .A2(n14279), .B1(n14814), .B2(n14278), .C1(
        n20043), .C2(n21136), .ZN(P1_U2894) );
  XNOR2_X1 U17569 ( .A(n9913), .B(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n14281) );
  XNOR2_X1 U17570 ( .A(n14280), .B(n14281), .ZN(n14298) );
  AOI22_X1 U17571 ( .A1(n20091), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .B1(
        n20103), .B2(P1_REIP_REG_9__SCAN_IN), .ZN(n14282) );
  OAI21_X1 U17572 ( .B1(n20102), .B2(n14283), .A(n14282), .ZN(n14284) );
  AOI21_X1 U17573 ( .B1(n20041), .B2(n20097), .A(n14284), .ZN(n14285) );
  OAI21_X1 U17574 ( .B1(n14298), .B2(n19949), .A(n14285), .ZN(P1_U2990) );
  INV_X1 U17575 ( .A(P1_REIP_REG_9__SCAN_IN), .ZN(n21039) );
  NOR2_X1 U17576 ( .A1(n20128), .A2(n21039), .ZN(n14296) );
  INV_X1 U17577 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n16184) );
  INV_X1 U17578 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16191) );
  NOR3_X1 U17579 ( .A1(n16184), .A2(n16191), .A3(n16181), .ZN(n15060) );
  NAND2_X1 U17580 ( .A1(n14286), .A2(n14289), .ZN(n14478) );
  INV_X1 U17581 ( .A(n14478), .ZN(n14287) );
  NAND2_X1 U17582 ( .A1(n15060), .A2(n14287), .ZN(n14292) );
  NOR2_X1 U17583 ( .A1(n16168), .A2(n14292), .ZN(n14294) );
  INV_X1 U17584 ( .A(n14288), .ZN(n14291) );
  NOR2_X1 U17585 ( .A1(n20121), .A2(n14289), .ZN(n20131) );
  NOR2_X1 U17586 ( .A1(n20131), .A2(n20123), .ZN(n14290) );
  OAI21_X1 U17587 ( .B1(n15054), .B2(n14291), .A(n14290), .ZN(n20116) );
  NAND2_X1 U17588 ( .A1(n16115), .A2(n20150), .ZN(n14482) );
  OAI21_X1 U17589 ( .B1(n20116), .B2(n14292), .A(n14482), .ZN(n15063) );
  INV_X1 U17590 ( .A(n15063), .ZN(n14293) );
  MUX2_X1 U17591 ( .A(n14294), .B(n14293), .S(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .Z(n14295) );
  AOI211_X1 U17592 ( .C1(n20114), .C2(n19965), .A(n14296), .B(n14295), .ZN(
        n14297) );
  OAI21_X1 U17593 ( .B1(n14298), .B2(n16177), .A(n14297), .ZN(P1_U3022) );
  INV_X1 U17594 ( .A(n14255), .ZN(n14302) );
  INV_X1 U17595 ( .A(n14300), .ZN(n14301) );
  NAND2_X1 U17596 ( .A1(n14302), .A2(n14301), .ZN(n14303) );
  NAND2_X1 U17597 ( .A1(n14299), .A2(n14303), .ZN(n14638) );
  XNOR2_X1 U17598 ( .A(n14638), .B(n14304), .ZN(n16085) );
  INV_X1 U17599 ( .A(n16085), .ZN(n16022) );
  INV_X1 U17600 ( .A(P1_EBX_REG_11__SCAN_IN), .ZN(n14310) );
  INV_X1 U17601 ( .A(n14305), .ZN(n14307) );
  INV_X1 U17602 ( .A(n14740), .ZN(n14306) );
  AOI21_X1 U17603 ( .B1(n14308), .B2(n14307), .A(n14306), .ZN(n16167) );
  INV_X1 U17604 ( .A(n16167), .ZN(n14309) );
  OAI222_X1 U17605 ( .A1(n16022), .A2(n14747), .B1(n14748), .B2(n14310), .C1(
        n14749), .C2(n14309), .ZN(P1_U2861) );
  INV_X1 U17606 ( .A(n14759), .ZN(n14311) );
  INV_X1 U17607 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n20053) );
  OAI222_X1 U17608 ( .A1(n16022), .A2(n14815), .B1(n14814), .B2(n14311), .C1(
        n20043), .C2(n20053), .ZN(P1_U2893) );
  NAND2_X1 U17609 ( .A1(n9875), .A2(n14312), .ZN(n14383) );
  OAI21_X1 U17610 ( .B1(n9875), .B2(n14312), .A(n14383), .ZN(n14327) );
  OR2_X1 U17611 ( .A1(n14315), .A2(n14314), .ZN(n14316) );
  NAND2_X1 U17612 ( .A1(n14313), .A2(n14316), .ZN(n18980) );
  AOI22_X1 U17613 ( .A1(n19110), .A2(BUF1_REG_17__SCAN_IN), .B1(n19109), .B2(
        BUF2_REG_17__SCAN_IN), .ZN(n14319) );
  AOI22_X1 U17614 ( .A1(n19108), .A2(n14317), .B1(n19155), .B2(
        P2_EAX_REG_17__SCAN_IN), .ZN(n14318) );
  OAI211_X1 U17615 ( .C1(n15285), .C2(n18980), .A(n14319), .B(n14318), .ZN(
        n14320) );
  INV_X1 U17616 ( .A(n14320), .ZN(n14321) );
  OAI21_X1 U17617 ( .B1(n14327), .B2(n19160), .A(n14321), .ZN(P2_U2902) );
  OAI21_X1 U17618 ( .B1(n14324), .B2(n14323), .A(n14322), .ZN(n15421) );
  NOR2_X1 U17619 ( .A1(n15421), .A2(n15192), .ZN(n14325) );
  AOI21_X1 U17620 ( .B1(P2_EBX_REG_17__SCAN_IN), .B2(n15234), .A(n14325), .ZN(
        n14326) );
  OAI21_X1 U17621 ( .B1(n14327), .B2(n15215), .A(n14326), .ZN(P2_U2870) );
  XNOR2_X1 U17622 ( .A(n14328), .B(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n14349) );
  XOR2_X1 U17623 ( .A(n14329), .B(n14330), .Z(n14347) );
  OAI22_X1 U17624 ( .A1(n19838), .A2(n15684), .B1(n19256), .B2(n19065), .ZN(
        n14331) );
  AOI21_X1 U17625 ( .B1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n19246), .A(
        n14331), .ZN(n14332) );
  OAI21_X1 U17626 ( .B1(n19066), .B2(n16305), .A(n14332), .ZN(n14333) );
  AOI21_X1 U17627 ( .B1(n14347), .B2(n19248), .A(n14333), .ZN(n14334) );
  OAI21_X1 U17628 ( .B1(n14349), .B2(n16295), .A(n14334), .ZN(P2_U3008) );
  NOR4_X1 U17629 ( .A1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n16351), .A3(
        n14339), .A4(n14335), .ZN(n14346) );
  XNOR2_X1 U17630 ( .A(n14336), .B(n14337), .ZN(n19139) );
  AOI21_X1 U17631 ( .B1(n15613), .B2(n14339), .A(n14338), .ZN(n15723) );
  INV_X1 U17632 ( .A(n15723), .ZN(n14341) );
  NOR2_X1 U17633 ( .A1(n19838), .A2(n15684), .ZN(n14340) );
  AOI21_X1 U17634 ( .B1(n14341), .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n14340), .ZN(n14344) );
  NAND2_X1 U17635 ( .A1(n14342), .A2(n16340), .ZN(n14343) );
  OAI211_X1 U17636 ( .C1(n19139), .C2(n16313), .A(n14344), .B(n14343), .ZN(
        n14345) );
  AOI211_X1 U17637 ( .C1(n14347), .C2(n16338), .A(n14346), .B(n14345), .ZN(
        n14348) );
  OAI21_X1 U17638 ( .B1(n14349), .B2(n16327), .A(n14348), .ZN(P2_U3040) );
  AND2_X1 U17639 ( .A1(n14208), .A2(n14350), .ZN(n14351) );
  NOR2_X1 U17640 ( .A1(n9875), .A2(n14351), .ZN(n19112) );
  NAND2_X1 U17641 ( .A1(n19112), .A2(n15231), .ZN(n14355) );
  XOR2_X1 U17642 ( .A(n14353), .B(n14352), .Z(n18995) );
  NAND2_X1 U17643 ( .A1(n18995), .A2(n15212), .ZN(n14354) );
  OAI211_X1 U17644 ( .C1(n15212), .C2(n18992), .A(n14355), .B(n14354), .ZN(
        P2_U2871) );
  OAI21_X1 U17645 ( .B1(n15739), .B2(n14357), .A(n14356), .ZN(n15748) );
  NAND2_X1 U17646 ( .A1(n19906), .A2(n19088), .ZN(n14361) );
  NAND2_X1 U17647 ( .A1(n9868), .A2(n10053), .ZN(n18977) );
  AOI22_X1 U17648 ( .A1(P2_EBX_REG_1__SCAN_IN), .A2(n19090), .B1(
        P2_REIP_REG_1__SCAN_IN), .B2(n19091), .ZN(n14358) );
  OAI21_X1 U17649 ( .B1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n18977), .A(
        n14358), .ZN(n14359) );
  AOI21_X1 U17650 ( .B1(n19101), .B2(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n14359), .ZN(n14360) );
  OAI211_X1 U17651 ( .C1(n19095), .C2(n14362), .A(n14361), .B(n14360), .ZN(
        n14365) );
  NOR2_X1 U17652 ( .A1(n19910), .A2(n14363), .ZN(n14364) );
  AOI211_X1 U17653 ( .C1(n19097), .C2(n12673), .A(n14365), .B(n14364), .ZN(
        n14366) );
  OAI21_X1 U17654 ( .B1(n15748), .B2(n19809), .A(n14366), .ZN(P2_U2854) );
  NAND2_X1 U17655 ( .A1(n14368), .A2(n14369), .ZN(n14370) );
  AND2_X1 U17656 ( .A1(n14730), .A2(n14370), .ZN(n16069) );
  INV_X1 U17657 ( .A(n16069), .ZN(n14374) );
  INV_X1 U17658 ( .A(DATAI_14_), .ZN(n14372) );
  MUX2_X1 U17659 ( .A(n14372), .B(n14371), .S(n20160), .Z(n20080) );
  INV_X1 U17660 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n14373) );
  OAI222_X1 U17661 ( .A1(n14374), .A2(n14815), .B1(n14814), .B2(n20080), .C1(
        n14373), .C2(n20043), .ZN(P1_U2890) );
  AND2_X1 U17662 ( .A1(n14642), .A2(n14375), .ZN(n14376) );
  OR2_X1 U17663 ( .A1(n14376), .A2(n14733), .ZN(n16137) );
  OAI22_X1 U17664 ( .A1(n16137), .A2(n14749), .B1(n16005), .B2(n14748), .ZN(
        n14377) );
  AOI21_X1 U17665 ( .B1(n16069), .B2(n14378), .A(n14377), .ZN(n14379) );
  INV_X1 U17666 ( .A(n14379), .ZN(P1_U2858) );
  AOI21_X1 U17667 ( .B1(n14381), .B2(n14322), .A(n14380), .ZN(n18973) );
  INV_X1 U17668 ( .A(n18973), .ZN(n15603) );
  AOI21_X1 U17669 ( .B1(n14384), .B2(n14383), .A(n14382), .ZN(n16235) );
  NAND2_X1 U17670 ( .A1(n16235), .A2(n15231), .ZN(n14386) );
  NAND2_X1 U17671 ( .A1(n15234), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n14385) );
  OAI211_X1 U17672 ( .C1(n15603), .C2(n15234), .A(n14386), .B(n14385), .ZN(
        P2_U2869) );
  OAI211_X1 U17673 ( .C1(n18844), .C2(n18700), .A(n10259), .B(n18691), .ZN(
        n18237) );
  NOR2_X1 U17674 ( .A1(P3_FLUSH_REG_SCAN_IN), .A2(n18237), .ZN(n14387) );
  NAND3_X1 U17675 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_0__SCAN_IN), .A3(P3_STATE2_REG_2__SCAN_IN), .ZN(n18836)
         );
  OAI21_X1 U17676 ( .B1(n14387), .B2(n18836), .A(n18342), .ZN(n18242) );
  INV_X1 U17677 ( .A(n18242), .ZN(n14388) );
  INV_X1 U17678 ( .A(n17867), .ZN(n17709) );
  NOR2_X1 U17679 ( .A1(n17709), .A2(n18883), .ZN(n15799) );
  AOI21_X1 U17680 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n15799), .ZN(n15800) );
  NOR2_X1 U17681 ( .A1(n14388), .A2(n15800), .ZN(n14390) );
  NOR2_X1 U17682 ( .A1(n18864), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n18281) );
  OR2_X1 U17683 ( .A1(n18281), .A2(n14388), .ZN(n15798) );
  OR2_X1 U17684 ( .A1(n18593), .A2(n15798), .ZN(n14389) );
  MUX2_X1 U17685 ( .A(n14390), .B(n14389), .S(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .Z(P3_U2864) );
  AND2_X1 U17686 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(P3_EBX_REG_27__SCAN_IN), 
        .ZN(n16993) );
  INV_X1 U17687 ( .A(n18682), .ZN(n15813) );
  NAND3_X1 U17688 ( .A1(n18277), .A2(n18262), .A3(n14391), .ZN(n14392) );
  NOR2_X1 U17689 ( .A1(n17356), .A2(n17266), .ZN(n17263) );
  INV_X1 U17690 ( .A(n17263), .ZN(n17269) );
  NAND2_X1 U17691 ( .A1(n14395), .A2(n17356), .ZN(n14394) );
  INV_X1 U17692 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n16651) );
  INV_X1 U17693 ( .A(P3_EBX_REG_18__SCAN_IN), .ZN(n17093) );
  INV_X1 U17694 ( .A(P3_EBX_REG_14__SCAN_IN), .ZN(n20937) );
  INV_X1 U17695 ( .A(P3_EBX_REG_10__SCAN_IN), .ZN(n17189) );
  INV_X1 U17696 ( .A(P3_EBX_REG_8__SCAN_IN), .ZN(n17233) );
  INV_X1 U17697 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n17230) );
  INV_X1 U17698 ( .A(P3_EBX_REG_2__SCAN_IN), .ZN(n17256) );
  NAND2_X1 U17699 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n17257) );
  NOR2_X1 U17700 ( .A1(n17256), .A2(n17257), .ZN(n17248) );
  NAND3_X1 U17701 ( .A1(P3_EBX_REG_7__SCAN_IN), .A2(P3_EBX_REG_6__SCAN_IN), 
        .A3(n17238), .ZN(n17210) );
  NOR2_X2 U17702 ( .A1(n20937), .A2(n17134), .ZN(n17133) );
  NAND2_X1 U17703 ( .A1(P3_EBX_REG_15__SCAN_IN), .A2(n17133), .ZN(n17131) );
  AND2_X2 U17704 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n17107), .ZN(n17120) );
  NAND3_X1 U17705 ( .A1(P3_EBX_REG_23__SCAN_IN), .A2(P3_EBX_REG_22__SCAN_IN), 
        .A3(P3_EBX_REG_21__SCAN_IN), .ZN(n16963) );
  NOR2_X2 U17706 ( .A1(n17052), .A2(n16963), .ZN(n17025) );
  NAND2_X1 U17707 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n17025), .ZN(n17012) );
  NAND2_X1 U17708 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n17015), .ZN(n17006) );
  NAND2_X1 U17709 ( .A1(n14394), .A2(n17006), .ZN(n17004) );
  OAI21_X1 U17710 ( .B1(n16993), .B2(n17269), .A(n17004), .ZN(n16998) );
  AOI22_X1 U17711 ( .A1(n17153), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n9837), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n14399) );
  AOI22_X1 U17712 ( .A1(n17219), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17098), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n14398) );
  AOI22_X1 U17713 ( .A1(n9849), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17213), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n14397) );
  AOI22_X1 U17714 ( .A1(n17112), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n15785), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n14396) );
  NAND4_X1 U17715 ( .A1(n14399), .A2(n14398), .A3(n14397), .A4(n14396), .ZN(
        n14405) );
  AOI22_X1 U17716 ( .A1(n17220), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17211), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n14403) );
  AOI22_X1 U17717 ( .A1(n17200), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n9839), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n14402) );
  AOI22_X1 U17718 ( .A1(n17147), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n9838), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n14401) );
  AOI22_X1 U17719 ( .A1(n17193), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17194), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n14400) );
  NAND4_X1 U17720 ( .A1(n14403), .A2(n14402), .A3(n14401), .A4(n14400), .ZN(
        n14404) );
  NOR2_X1 U17721 ( .A1(n14405), .A2(n14404), .ZN(n17002) );
  AOI22_X1 U17722 ( .A1(n17200), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n17112), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n14409) );
  AOI22_X1 U17723 ( .A1(n17193), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17194), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n14408) );
  AOI22_X1 U17724 ( .A1(n17147), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n9838), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n14407) );
  AOI22_X1 U17725 ( .A1(n17192), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n15785), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n14406) );
  NAND4_X1 U17726 ( .A1(n14409), .A2(n14408), .A3(n14407), .A4(n14406), .ZN(
        n14415) );
  AOI22_X1 U17727 ( .A1(n9851), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n17220), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n14413) );
  AOI22_X1 U17728 ( .A1(n17098), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n17153), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n14412) );
  AOI22_X1 U17729 ( .A1(n9837), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17211), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n14411) );
  AOI22_X1 U17730 ( .A1(n9849), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(n9839), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n14410) );
  NAND4_X1 U17731 ( .A1(n14413), .A2(n14412), .A3(n14411), .A4(n14410), .ZN(
        n14414) );
  NOR2_X1 U17732 ( .A1(n14415), .A2(n14414), .ZN(n17013) );
  AOI22_X1 U17733 ( .A1(n17200), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17194), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n14419) );
  AOI22_X1 U17734 ( .A1(n9849), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(n9837), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n14418) );
  AOI22_X1 U17735 ( .A1(n17098), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n17216), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n14417) );
  AOI22_X1 U17736 ( .A1(n17112), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n15785), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n14416) );
  NAND4_X1 U17737 ( .A1(n14419), .A2(n14418), .A3(n14417), .A4(n14416), .ZN(
        n14425) );
  AOI22_X1 U17738 ( .A1(n17153), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n9839), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n14423) );
  AOI22_X1 U17739 ( .A1(n17219), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17220), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n14422) );
  AOI22_X1 U17740 ( .A1(n9838), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17213), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n14421) );
  AOI22_X1 U17741 ( .A1(n17193), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17211), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n14420) );
  NAND4_X1 U17742 ( .A1(n14423), .A2(n14422), .A3(n14421), .A4(n14420), .ZN(
        n14424) );
  NOR2_X1 U17743 ( .A1(n14425), .A2(n14424), .ZN(n17023) );
  AOI22_X1 U17744 ( .A1(n17199), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n17177), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n14429) );
  AOI22_X1 U17745 ( .A1(n17193), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n17212), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n14428) );
  AOI22_X1 U17746 ( .A1(n9839), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n17213), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n14427) );
  AOI22_X1 U17747 ( .A1(n9837), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n15785), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n14426) );
  NAND4_X1 U17748 ( .A1(n14429), .A2(n14428), .A3(n14427), .A4(n14426), .ZN(
        n14435) );
  AOI22_X1 U17749 ( .A1(n9832), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n17112), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n14433) );
  AOI22_X1 U17750 ( .A1(n17217), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n9838), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n14432) );
  AOI22_X1 U17751 ( .A1(n9849), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n17216), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n14431) );
  AOI22_X1 U17752 ( .A1(n9851), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n17211), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n14430) );
  NAND4_X1 U17753 ( .A1(n14433), .A2(n14432), .A3(n14431), .A4(n14430), .ZN(
        n14434) );
  NOR2_X1 U17754 ( .A1(n14435), .A2(n14434), .ZN(n17022) );
  NOR2_X1 U17755 ( .A1(n17023), .A2(n17022), .ZN(n17018) );
  AOI22_X1 U17756 ( .A1(n17199), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n17211), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n14446) );
  AOI22_X1 U17757 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n9838), .B1(
        n17112), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n14445) );
  AOI22_X1 U17758 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n17192), .B1(
        P3_INSTQUEUE_REG_13__1__SCAN_IN), .B2(n17220), .ZN(n14436) );
  OAI21_X1 U17759 ( .B1(n14437), .B2(n21120), .A(n14436), .ZN(n14443) );
  AOI22_X1 U17760 ( .A1(n9832), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(n9837), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n14441) );
  AOI22_X1 U17761 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n17153), .B1(
        P3_INSTQUEUE_REG_12__1__SCAN_IN), .B2(n17193), .ZN(n14440) );
  AOI22_X1 U17762 ( .A1(n17217), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_2__1__SCAN_IN), .B2(n15785), .ZN(n14439) );
  AOI22_X1 U17763 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n17147), .B1(
        P3_INSTQUEUE_REG_9__1__SCAN_IN), .B2(n9839), .ZN(n14438) );
  NAND4_X1 U17764 ( .A1(n14441), .A2(n14440), .A3(n14439), .A4(n14438), .ZN(
        n14442) );
  AOI211_X1 U17765 ( .C1(n17219), .C2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A(
        n14443), .B(n14442), .ZN(n14444) );
  NAND3_X1 U17766 ( .A1(n14446), .A2(n14445), .A3(n14444), .ZN(n17017) );
  NAND2_X1 U17767 ( .A1(n17018), .A2(n17017), .ZN(n17016) );
  NOR2_X1 U17768 ( .A1(n17013), .A2(n17016), .ZN(n17009) );
  AOI22_X1 U17769 ( .A1(n9832), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17216), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n14456) );
  AOI22_X1 U17770 ( .A1(n9849), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17213), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n14455) );
  AOI22_X1 U17771 ( .A1(n17193), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17177), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n14447) );
  OAI21_X1 U17772 ( .B1(n17136), .B2(n21055), .A(n14447), .ZN(n14453) );
  AOI22_X1 U17773 ( .A1(n9838), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(n9839), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n14451) );
  AOI22_X1 U17774 ( .A1(n17153), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n17112), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n14450) );
  AOI22_X1 U17775 ( .A1(n17219), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n9837), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n14449) );
  AOI22_X1 U17776 ( .A1(n17211), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n15785), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n14448) );
  NAND4_X1 U17777 ( .A1(n14451), .A2(n14450), .A3(n14449), .A4(n14448), .ZN(
        n14452) );
  AOI211_X1 U17778 ( .C1(n17098), .C2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .A(
        n14453), .B(n14452), .ZN(n14454) );
  NAND3_X1 U17779 ( .A1(n14456), .A2(n14455), .A3(n14454), .ZN(n17008) );
  NAND2_X1 U17780 ( .A1(n17009), .A2(n17008), .ZN(n17007) );
  NOR2_X1 U17781 ( .A1(n17002), .A2(n17007), .ZN(n17001) );
  AOI22_X1 U17782 ( .A1(n9849), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17153), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n14460) );
  AOI22_X1 U17783 ( .A1(n9851), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n17194), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n14459) );
  AOI22_X1 U17784 ( .A1(n9832), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17211), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n14458) );
  AOI22_X1 U17785 ( .A1(n9837), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n15785), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n14457) );
  NAND4_X1 U17786 ( .A1(n14460), .A2(n14459), .A3(n14458), .A4(n14457), .ZN(
        n14466) );
  AOI22_X1 U17787 ( .A1(n17147), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n17213), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n14464) );
  AOI22_X1 U17788 ( .A1(n17220), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n9839), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n14463) );
  AOI22_X1 U17789 ( .A1(n17112), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n9838), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n14462) );
  AOI22_X1 U17790 ( .A1(n17199), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n17193), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n14461) );
  NAND4_X1 U17791 ( .A1(n14464), .A2(n14463), .A3(n14462), .A4(n14461), .ZN(
        n14465) );
  NOR2_X1 U17792 ( .A1(n14466), .A2(n14465), .ZN(n16994) );
  XNOR2_X1 U17793 ( .A(n17001), .B(n16994), .ZN(n17285) );
  AOI22_X1 U17794 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n16998), .B1(n17267), 
        .B2(n17285), .ZN(n14469) );
  INV_X1 U17795 ( .A(P3_EBX_REG_28__SCAN_IN), .ZN(n14467) );
  INV_X1 U17796 ( .A(n17006), .ZN(n17011) );
  NAND3_X1 U17797 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(n14467), .A3(n17011), 
        .ZN(n14468) );
  NAND2_X1 U17798 ( .A1(n14469), .A2(n14468), .ZN(P3_U2675) );
  NOR2_X1 U17799 ( .A1(n14470), .A2(n15192), .ZN(n14471) );
  AOI21_X1 U17800 ( .B1(P2_EBX_REG_30__SCAN_IN), .B2(n15192), .A(n14471), .ZN(
        n14472) );
  OAI21_X1 U17801 ( .B1(n14473), .B2(n15215), .A(n14472), .ZN(P2_U2857) );
  INV_X1 U17802 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n21070) );
  NOR2_X1 U17803 ( .A1(n15025), .A2(n21070), .ZN(n15017) );
  NAND3_X1 U17804 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A3(n15060), .ZN(n16154) );
  OR3_X1 U17805 ( .A1(n16199), .A2(n14477), .A3(n16154), .ZN(n16158) );
  NAND3_X1 U17806 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n14490) );
  NOR2_X1 U17807 ( .A1(n16158), .A2(n14490), .ZN(n15053) );
  INV_X1 U17808 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15048) );
  NOR3_X1 U17809 ( .A1(n15048), .A2(n16143), .A3(n15047), .ZN(n16124) );
  NAND2_X1 U17810 ( .A1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n16124), .ZN(
        n16117) );
  NOR2_X1 U17811 ( .A1(n16123), .A2(n16117), .ZN(n14491) );
  INV_X1 U17812 ( .A(n14491), .ZN(n14480) );
  INV_X1 U17813 ( .A(n14490), .ZN(n14479) );
  NOR2_X1 U17814 ( .A1(n16154), .A2(n14478), .ZN(n16171) );
  NAND2_X1 U17815 ( .A1(n14479), .A2(n16171), .ZN(n15050) );
  AOI221_X1 U17816 ( .B1(n14480), .B2(n15051), .C1(n15050), .C2(n15051), .A(
        n20123), .ZN(n14481) );
  OAI221_X1 U17817 ( .B1(n15054), .B2(n15053), .C1(n15054), .C2(n14491), .A(
        n14481), .ZN(n16111) );
  OAI21_X1 U17818 ( .B1(n14492), .B2(n16111), .A(n14482), .ZN(n15026) );
  OAI21_X1 U17819 ( .B1(n16115), .B2(n15017), .A(n15026), .ZN(n15011) );
  NOR2_X1 U17820 ( .A1(n20121), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14483) );
  NOR2_X1 U17821 ( .A1(n15011), .A2(n14483), .ZN(n14998) );
  NAND2_X1 U17822 ( .A1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n14485) );
  NOR2_X1 U17823 ( .A1(n20121), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14484) );
  AOI21_X1 U17824 ( .B1(n20125), .B2(n14485), .A(n14484), .ZN(n14486) );
  NAND2_X1 U17825 ( .A1(n14998), .A2(n14486), .ZN(n14995) );
  INV_X1 U17826 ( .A(n14495), .ZN(n14487) );
  OR2_X1 U17827 ( .A1(n14995), .A2(n14487), .ZN(n14968) );
  INV_X1 U17828 ( .A(n14963), .ZN(n14951) );
  NAND2_X1 U17829 ( .A1(n14998), .A2(n16115), .ZN(n14967) );
  OAI21_X1 U17830 ( .B1(n14968), .B2(n14951), .A(n14967), .ZN(n14950) );
  OAI21_X1 U17831 ( .B1(n16115), .B2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14488) );
  INV_X1 U17832 ( .A(n14488), .ZN(n14489) );
  NAND2_X1 U17833 ( .A1(n14950), .A2(n14489), .ZN(n14945) );
  NAND3_X1 U17834 ( .A1(n14945), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n14967), .ZN(n14499) );
  NAND2_X1 U17835 ( .A1(n20103), .A2(P1_REIP_REG_31__SCAN_IN), .ZN(n14503) );
  NOR2_X1 U17836 ( .A1(n16158), .A2(n20120), .ZN(n16153) );
  AOI21_X1 U17837 ( .B1(n16171), .B2(n15051), .A(n16153), .ZN(n16152) );
  NAND2_X1 U17838 ( .A1(n14491), .A2(n16140), .ZN(n16108) );
  INV_X1 U17839 ( .A(n14492), .ZN(n14493) );
  NAND3_X1 U17840 ( .A1(n14493), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n14494) );
  NOR2_X1 U17841 ( .A1(n16108), .A2(n14494), .ZN(n15000) );
  AND2_X1 U17842 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14986) );
  AND2_X1 U17843 ( .A1(n14495), .A2(n14986), .ZN(n14496) );
  NAND2_X1 U17844 ( .A1(n15000), .A2(n14496), .ZN(n14975) );
  NAND2_X1 U17845 ( .A1(n14963), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14497) );
  NOR2_X1 U17846 ( .A1(n14975), .A2(n14497), .ZN(n14946) );
  NAND3_X1 U17847 ( .A1(n14946), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n13722), .ZN(n14498) );
  INV_X1 U17848 ( .A(n14500), .ZN(n14501) );
  OAI21_X1 U17849 ( .B1(n14508), .B2(n16177), .A(n14501), .ZN(P1_U3000) );
  NAND2_X1 U17850 ( .A1(n20091), .A2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14502) );
  OAI211_X1 U17851 ( .C1(n20102), .C2(n14504), .A(n14503), .B(n14502), .ZN(
        n14505) );
  AOI21_X1 U17852 ( .B1(n14506), .B2(n20097), .A(n14505), .ZN(n14507) );
  OAI21_X1 U17853 ( .B1(n14508), .B2(n19949), .A(n14507), .ZN(P1_U2968) );
  AND2_X1 U17854 ( .A1(n14571), .A2(n14510), .ZN(n14511) );
  NOR2_X1 U17855 ( .A1(n14552), .A2(n14511), .ZN(n14952) );
  AOI22_X1 U17856 ( .A1(n14952), .A2(n14719), .B1(n14718), .B2(
        P1_EBX_REG_29__SCAN_IN), .ZN(n14512) );
  OAI21_X1 U17857 ( .B1(n14509), .B2(n14747), .A(n14512), .ZN(P1_U2843) );
  NOR2_X1 U17858 ( .A1(n14559), .A2(P1_REIP_REG_29__SCAN_IN), .ZN(n14517) );
  AOI22_X1 U17859 ( .A1(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n20026), .B1(
        n20034), .B2(n14513), .ZN(n14515) );
  NAND2_X1 U17860 ( .A1(n20025), .A2(P1_EBX_REG_29__SCAN_IN), .ZN(n14514) );
  OAI211_X1 U17861 ( .C1(n14579), .C2(n20751), .A(n14515), .B(n14514), .ZN(
        n14516) );
  AOI211_X1 U17862 ( .C1(n14952), .C2(n20010), .A(n14517), .B(n14516), .ZN(
        n14518) );
  OAI21_X1 U17863 ( .B1(n14509), .B2(n16023), .A(n14518), .ZN(P1_U2811) );
  AOI22_X1 U17864 ( .A1(n14796), .A2(BUF1_REG_29__SCAN_IN), .B1(
        P1_EAX_REG_29__SCAN_IN), .B2(n14816), .ZN(n14521) );
  NAND3_X1 U17865 ( .A1(n20043), .A2(n10418), .A3(n14519), .ZN(n14803) );
  AOI22_X1 U17866 ( .A1(n14806), .A2(DATAI_29_), .B1(n14798), .B2(n14812), 
        .ZN(n14520) );
  OAI211_X1 U17867 ( .C1(n14509), .C2(n14815), .A(n14521), .B(n14520), .ZN(
        P1_U2875) );
  AOI21_X1 U17868 ( .B1(n14524), .B2(n14523), .A(n14522), .ZN(n14544) );
  OAI21_X1 U17869 ( .B1(n14529), .B2(n21090), .A(n14525), .ZN(n14526) );
  AOI22_X1 U17870 ( .A1(n16342), .A2(n14544), .B1(n15610), .B2(n14526), .ZN(
        n14537) );
  XOR2_X1 U17871 ( .A(n14528), .B(n14527), .Z(n14538) );
  NAND2_X1 U17872 ( .A1(n19038), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n14540) );
  OAI21_X1 U17873 ( .B1(n14530), .B2(n14529), .A(n14540), .ZN(n14531) );
  AOI21_X1 U17874 ( .B1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n14532), .A(
        n14531), .ZN(n14533) );
  OAI21_X1 U17875 ( .B1(n14534), .B2(n16313), .A(n14533), .ZN(n14535) );
  AOI21_X1 U17876 ( .B1(n16338), .B2(n14538), .A(n14535), .ZN(n14536) );
  OAI211_X1 U17877 ( .C1(n13628), .C2(n16326), .A(n14537), .B(n14536), .ZN(
        P2_U3044) );
  NAND2_X1 U17878 ( .A1(n14538), .A2(n19248), .ZN(n14546) );
  INV_X1 U17879 ( .A(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n14542) );
  NAND2_X1 U17880 ( .A1(n16302), .A2(n14539), .ZN(n14541) );
  OAI211_X1 U17881 ( .C1(n16310), .C2(n14542), .A(n14541), .B(n14540), .ZN(
        n14543) );
  AOI21_X1 U17882 ( .B1(n14544), .B2(n19251), .A(n14543), .ZN(n14545) );
  OAI211_X1 U17883 ( .C1(n16305), .C2(n10247), .A(n14546), .B(n14545), .ZN(
        P2_U3012) );
  INV_X1 U17884 ( .A(n14547), .ZN(n19946) );
  NAND2_X1 U17885 ( .A1(n14548), .A2(P1_MEMORYFETCH_REG_SCAN_IN), .ZN(n14549)
         );
  NAND3_X1 U17886 ( .A1(n14550), .A2(n19946), .A3(n14549), .ZN(P1_U2801) );
  OAI22_X1 U17887 ( .A1(n14552), .A2(n9835), .B1(n14571), .B2(n14551), .ZN(
        n14555) );
  INV_X1 U17888 ( .A(n14553), .ZN(n14554) );
  XNOR2_X1 U17889 ( .A(n14555), .B(n14554), .ZN(n14942) );
  NAND2_X1 U17890 ( .A1(n14824), .A2(n19992), .ZN(n14566) );
  OAI21_X1 U17891 ( .B1(n14559), .B2(n20751), .A(n14820), .ZN(n14564) );
  INV_X1 U17892 ( .A(P1_EBX_REG_30__SCAN_IN), .ZN(n21110) );
  NOR2_X1 U17893 ( .A1(n19997), .A2(n21110), .ZN(n14562) );
  OAI22_X1 U17894 ( .A1(n14560), .A2(n20014), .B1(n20006), .B2(n14822), .ZN(
        n14561) );
  AOI211_X1 U17895 ( .C1(n14564), .C2(n14563), .A(n14562), .B(n14561), .ZN(
        n14565) );
  OAI211_X1 U17896 ( .C1(n20038), .C2(n14942), .A(n14566), .B(n14565), .ZN(
        P1_U2810) );
  AOI21_X1 U17897 ( .B1(n14592), .B2(P1_REIP_REG_27__SCAN_IN), .A(
        P1_REIP_REG_28__SCAN_IN), .ZN(n14578) );
  AOI21_X1 U17899 ( .B1(n14568), .B2(n14581), .A(n12655), .ZN(n14836) );
  NAND2_X1 U17900 ( .A1(n14836), .A2(n19992), .ZN(n14577) );
  OAI22_X1 U17901 ( .A1(n14569), .A2(n20014), .B1(n20006), .B2(n14834), .ZN(
        n14575) );
  INV_X1 U17902 ( .A(n14586), .ZN(n14573) );
  INV_X1 U17903 ( .A(n14570), .ZN(n14572) );
  OAI21_X1 U17904 ( .B1(n14573), .B2(n14572), .A(n14571), .ZN(n14960) );
  NOR2_X1 U17905 ( .A1(n14960), .A2(n20038), .ZN(n14574) );
  AOI211_X1 U17906 ( .C1(n20025), .C2(P1_EBX_REG_28__SCAN_IN), .A(n14575), .B(
        n14574), .ZN(n14576) );
  OAI211_X1 U17907 ( .C1(n14579), .C2(n14578), .A(n14577), .B(n14576), .ZN(
        P1_U2812) );
  NAND2_X1 U17908 ( .A1(n14583), .A2(n14584), .ZN(n14585) );
  AOI22_X1 U17909 ( .A1(n14845), .A2(n20034), .B1(P1_EBX_REG_27__SCAN_IN), 
        .B2(n20025), .ZN(n14587) );
  OAI21_X1 U17910 ( .B1(n21108), .B2(n20014), .A(n14587), .ZN(n14588) );
  INV_X1 U17911 ( .A(n14588), .ZN(n14590) );
  NAND2_X1 U17912 ( .A1(n14601), .A2(P1_REIP_REG_27__SCAN_IN), .ZN(n14589) );
  NAND2_X1 U17913 ( .A1(n14590), .A2(n14589), .ZN(n14591) );
  AOI21_X1 U17914 ( .B1(n14972), .B2(n20010), .A(n14591), .ZN(n14594) );
  INV_X1 U17915 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n20749) );
  NAND2_X1 U17916 ( .A1(n14592), .A2(n20749), .ZN(n14593) );
  OAI211_X1 U17917 ( .C1(n14842), .C2(n16023), .A(n14594), .B(n14593), .ZN(
        P1_U2813) );
  AOI21_X1 U17918 ( .B1(n14595), .B2(n9829), .A(n14580), .ZN(n14853) );
  INV_X1 U17919 ( .A(n14853), .ZN(n14765) );
  OAI22_X1 U17920 ( .A1(n14596), .A2(n20014), .B1(n20006), .B2(n14851), .ZN(
        n14600) );
  OAI21_X1 U17921 ( .B1(n14598), .B2(n14597), .A(n14583), .ZN(n14980) );
  NOR2_X1 U17922 ( .A1(n14980), .A2(n20038), .ZN(n14599) );
  AOI211_X1 U17923 ( .C1(P1_EBX_REG_26__SCAN_IN), .C2(n20025), .A(n14600), .B(
        n14599), .ZN(n14604) );
  AND3_X1 U17924 ( .A1(n15935), .A2(P1_REIP_REG_24__SCAN_IN), .A3(
        P1_REIP_REG_25__SCAN_IN), .ZN(n14602) );
  OAI21_X1 U17925 ( .B1(n14602), .B2(P1_REIP_REG_26__SCAN_IN), .A(n14601), 
        .ZN(n14603) );
  OAI211_X1 U17926 ( .C1(n14765), .C2(n16023), .A(n14604), .B(n14603), .ZN(
        P1_U2814) );
  OAI21_X1 U17927 ( .B1(n14605), .B2(n14608), .A(n14607), .ZN(n14885) );
  NAND2_X1 U17928 ( .A1(P1_REIP_REG_16__SCAN_IN), .A2(P1_REIP_REG_15__SCAN_IN), 
        .ZN(n15991) );
  NAND3_X1 U17929 ( .A1(P1_REIP_REG_13__SCAN_IN), .A2(P1_REIP_REG_12__SCAN_IN), 
        .A3(P1_REIP_REG_11__SCAN_IN), .ZN(n14609) );
  NAND3_X1 U17930 ( .A1(n19970), .A2(P1_REIP_REG_9__SCAN_IN), .A3(
        P1_REIP_REG_10__SCAN_IN), .ZN(n16027) );
  NOR2_X1 U17931 ( .A1(n14609), .A2(n16027), .ZN(n16008) );
  NAND2_X1 U17932 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(n16008), .ZN(n16004) );
  NOR2_X1 U17933 ( .A1(n15991), .A2(n16004), .ZN(n14629) );
  NAND2_X1 U17934 ( .A1(P1_REIP_REG_17__SCAN_IN), .A2(n14629), .ZN(n15984) );
  NOR2_X1 U17935 ( .A1(P1_REIP_REG_19__SCAN_IN), .A2(n15984), .ZN(n14622) );
  INV_X1 U17936 ( .A(n14610), .ZN(n14612) );
  AND3_X1 U17937 ( .A1(P1_REIP_REG_9__SCAN_IN), .A2(P1_REIP_REG_10__SCAN_IN), 
        .A3(n14611), .ZN(n16019) );
  AOI21_X1 U17938 ( .B1(n14612), .B2(n16019), .A(n16020), .ZN(n16007) );
  AOI21_X1 U17939 ( .B1(n14614), .B2(n14613), .A(n16007), .ZN(n14627) );
  OAI21_X1 U17940 ( .B1(n16020), .B2(P1_REIP_REG_18__SCAN_IN), .A(n14627), 
        .ZN(n15985) );
  AOI22_X1 U17941 ( .A1(P1_EBX_REG_19__SCAN_IN), .A2(n20025), .B1(
        P1_REIP_REG_19__SCAN_IN), .B2(n15985), .ZN(n14615) );
  OAI211_X1 U17942 ( .C1(n20014), .C2(n14616), .A(n14615), .B(n20011), .ZN(
        n14621) );
  NOR2_X1 U17943 ( .A1(n14714), .A2(n14617), .ZN(n14618) );
  OR2_X1 U17944 ( .A1(n14703), .A2(n14618), .ZN(n16105) );
  INV_X1 U17945 ( .A(n14619), .ZN(n14887) );
  OAI22_X1 U17946 ( .A1(n16105), .A2(n20038), .B1(n14887), .B2(n20006), .ZN(
        n14620) );
  AOI211_X1 U17947 ( .C1(n14622), .C2(P1_REIP_REG_18__SCAN_IN), .A(n14621), 
        .B(n14620), .ZN(n14623) );
  OAI21_X1 U17948 ( .B1(n14885), .B2(n16023), .A(n14623), .ZN(P1_U2821) );
  OAI21_X1 U17949 ( .B1(n14624), .B2(n14626), .A(n14625), .ZN(n14905) );
  INV_X1 U17950 ( .A(n14627), .ZN(n14628) );
  OAI21_X1 U17951 ( .B1(P1_REIP_REG_17__SCAN_IN), .B2(n14629), .A(n14628), 
        .ZN(n14636) );
  NAND2_X1 U17952 ( .A1(n14725), .A2(n14630), .ZN(n14631) );
  AND2_X1 U17953 ( .A1(n14713), .A2(n14631), .ZN(n16125) );
  AOI22_X1 U17954 ( .A1(n14902), .A2(n20034), .B1(P1_EBX_REG_17__SCAN_IN), 
        .B2(n20025), .ZN(n14632) );
  OAI211_X1 U17955 ( .C1(n20014), .C2(n14633), .A(n14632), .B(n20011), .ZN(
        n14634) );
  AOI21_X1 U17956 ( .B1(n20010), .B2(n16125), .A(n14634), .ZN(n14635) );
  OAI211_X1 U17957 ( .C1(n14905), .C2(n16023), .A(n14636), .B(n14635), .ZN(
        P1_U2823) );
  NAND2_X1 U17958 ( .A1(n14639), .A2(n14299), .ZN(n14744) );
  OAI21_X1 U17959 ( .B1(n14746), .B2(n14640), .A(n14368), .ZN(n14933) );
  NAND2_X1 U17960 ( .A1(P1_REIP_REG_12__SCAN_IN), .A2(P1_REIP_REG_11__SCAN_IN), 
        .ZN(n14645) );
  NOR3_X1 U17961 ( .A1(P1_REIP_REG_13__SCAN_IN), .A2(n14645), .A3(n16027), 
        .ZN(n14651) );
  INV_X1 U17962 ( .A(n14641), .ZN(n14742) );
  INV_X1 U17963 ( .A(n14642), .ZN(n14643) );
  AOI21_X1 U17964 ( .B1(n14644), .B2(n14742), .A(n14643), .ZN(n16146) );
  INV_X1 U17965 ( .A(n14645), .ZN(n14646) );
  AOI21_X1 U17966 ( .B1(n14646), .B2(n16019), .A(n16020), .ZN(n16015) );
  AOI22_X1 U17967 ( .A1(n20010), .A2(n16146), .B1(P1_REIP_REG_13__SCAN_IN), 
        .B2(n16015), .ZN(n14647) );
  OAI211_X1 U17968 ( .C1(n20014), .C2(n14648), .A(n14647), .B(n20011), .ZN(
        n14650) );
  INV_X1 U17969 ( .A(P1_EBX_REG_13__SCAN_IN), .ZN(n14738) );
  OAI22_X1 U17970 ( .A1(n20006), .A2(n14929), .B1(n19997), .B2(n14738), .ZN(
        n14649) );
  NOR3_X1 U17971 ( .A1(n14651), .A2(n14650), .A3(n14649), .ZN(n14652) );
  OAI21_X1 U17972 ( .B1(n14933), .B2(n16023), .A(n14652), .ZN(P1_U2827) );
  NAND2_X1 U17973 ( .A1(n20014), .A2(n20006), .ZN(n14653) );
  AOI22_X1 U17974 ( .A1(n14653), .A2(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .B1(
        n10551), .B2(n20027), .ZN(n14654) );
  OAI21_X1 U17975 ( .B1(n20038), .B2(n14655), .A(n14654), .ZN(n14659) );
  INV_X1 U17976 ( .A(P1_REIP_REG_0__SCAN_IN), .ZN(n14657) );
  OAI22_X1 U17977 ( .A1(n16020), .A2(n14657), .B1(n14656), .B2(n19997), .ZN(
        n14658) );
  AOI211_X1 U17978 ( .C1(n14660), .C2(n20017), .A(n14659), .B(n14658), .ZN(
        n14661) );
  INV_X1 U17979 ( .A(n14661), .ZN(P1_U2840) );
  OAI22_X1 U17980 ( .A1(n14663), .A2(n14749), .B1(n14662), .B2(n14748), .ZN(
        P1_U2841) );
  OAI222_X1 U17981 ( .A1(n14747), .A2(n14753), .B1(n14748), .B2(n21110), .C1(
        n14942), .C2(n14749), .ZN(P1_U2842) );
  INV_X1 U17982 ( .A(n14836), .ZN(n14758) );
  OAI222_X1 U17983 ( .A1(n14664), .A2(n14748), .B1(n14749), .B2(n14960), .C1(
        n14758), .C2(n14747), .ZN(P1_U2844) );
  AOI22_X1 U17984 ( .A1(n14972), .A2(n14719), .B1(P1_EBX_REG_27__SCAN_IN), 
        .B2(n14718), .ZN(n14665) );
  OAI21_X1 U17985 ( .B1(n14842), .B2(n14747), .A(n14665), .ZN(P1_U2845) );
  OAI222_X1 U17986 ( .A1(n14666), .A2(n14748), .B1(n14749), .B2(n14980), .C1(
        n14765), .C2(n14747), .ZN(P1_U2846) );
  NAND2_X1 U17987 ( .A1(n14667), .A2(n14668), .ZN(n14669) );
  NAND2_X1 U17988 ( .A1(n9829), .A2(n14669), .ZN(n15928) );
  XNOR2_X1 U17989 ( .A(n14670), .B(n14671), .ZN(n15934) );
  OAI22_X1 U17990 ( .A1(n15934), .A2(n14749), .B1(n20935), .B2(n14748), .ZN(
        n14672) );
  INV_X1 U17991 ( .A(n14672), .ZN(n14673) );
  OAI21_X1 U17992 ( .B1(n15928), .B2(n14747), .A(n14673), .ZN(P1_U2847) );
  OAI21_X1 U17993 ( .B1(n14674), .B2(n14675), .A(n14667), .ZN(n14864) );
  OR2_X1 U17994 ( .A1(n14683), .A2(n14676), .ZN(n14677) );
  NAND2_X1 U17995 ( .A1(n14670), .A2(n14677), .ZN(n15944) );
  OAI22_X1 U17996 ( .A1(n15944), .A2(n14749), .B1(n15936), .B2(n14748), .ZN(
        n14678) );
  INV_X1 U17997 ( .A(n14678), .ZN(n14679) );
  OAI21_X1 U17998 ( .B1(n14864), .B2(n14747), .A(n14679), .ZN(P1_U2848) );
  INV_X1 U17999 ( .A(n14674), .ZN(n14681) );
  INV_X1 U18000 ( .A(P1_EBX_REG_23__SCAN_IN), .ZN(n14687) );
  INV_X1 U18001 ( .A(n14683), .ZN(n14686) );
  NAND2_X1 U18002 ( .A1(n14690), .A2(n14684), .ZN(n14685) );
  NAND2_X1 U18003 ( .A1(n14686), .A2(n14685), .ZN(n15947) );
  OAI222_X1 U18004 ( .A1(n14747), .A2(n15948), .B1(n14748), .B2(n14687), .C1(
        n15947), .C2(n14749), .ZN(P1_U2849) );
  NAND2_X1 U18005 ( .A1(n14700), .A2(n14688), .ZN(n14689) );
  NAND2_X1 U18006 ( .A1(n14690), .A2(n14689), .ZN(n15964) );
  INV_X1 U18007 ( .A(P1_EBX_REG_22__SCAN_IN), .ZN(n21060) );
  AND2_X1 U18008 ( .A1(n14691), .A2(n14692), .ZN(n14693) );
  OR2_X1 U18009 ( .A1(n14693), .A2(n14680), .ZN(n15955) );
  OAI222_X1 U18010 ( .A1(n14749), .A2(n15964), .B1(n14748), .B2(n21060), .C1(
        n15955), .C2(n14747), .ZN(P1_U2850) );
  INV_X1 U18011 ( .A(n14691), .ZN(n14695) );
  AOI21_X1 U18012 ( .B1(n14696), .B2(n14707), .A(n14695), .ZN(n14878) );
  INV_X1 U18013 ( .A(n14878), .ZN(n15967) );
  INV_X1 U18014 ( .A(P1_EBX_REG_21__SCAN_IN), .ZN(n14701) );
  NAND2_X1 U18015 ( .A1(n14697), .A2(n14698), .ZN(n14699) );
  AND2_X1 U18016 ( .A1(n14700), .A2(n14699), .ZN(n15029) );
  INV_X1 U18017 ( .A(n15029), .ZN(n15966) );
  OAI222_X1 U18018 ( .A1(n14747), .A2(n15967), .B1(n14748), .B2(n14701), .C1(
        n15966), .C2(n14749), .ZN(P1_U2851) );
  OR2_X1 U18019 ( .A1(n14703), .A2(n14702), .ZN(n14704) );
  NAND2_X1 U18020 ( .A1(n14697), .A2(n14704), .ZN(n15980) );
  INV_X1 U18021 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n14708) );
  NAND2_X1 U18022 ( .A1(n14607), .A2(n14705), .ZN(n14706) );
  AND2_X1 U18023 ( .A1(n14707), .A2(n14706), .ZN(n16044) );
  INV_X1 U18024 ( .A(n16044), .ZN(n14786) );
  OAI222_X1 U18025 ( .A1(n14749), .A2(n15980), .B1(n14748), .B2(n14708), .C1(
        n14747), .C2(n14786), .ZN(P1_U2852) );
  INV_X1 U18026 ( .A(P1_EBX_REG_19__SCAN_IN), .ZN(n14709) );
  OAI222_X1 U18027 ( .A1(n14747), .A2(n14885), .B1(n14748), .B2(n14709), .C1(
        n16105), .C2(n14749), .ZN(P1_U2853) );
  AND2_X1 U18028 ( .A1(n14625), .A2(n14710), .ZN(n14711) );
  OR2_X1 U18029 ( .A1(n14605), .A2(n14711), .ZN(n15983) );
  AND2_X1 U18030 ( .A1(n14713), .A2(n14712), .ZN(n14715) );
  OR2_X1 U18031 ( .A1(n14715), .A2(n14714), .ZN(n16116) );
  OAI22_X1 U18032 ( .A1(n16116), .A2(n14749), .B1(n15981), .B2(n14748), .ZN(
        n14716) );
  INV_X1 U18033 ( .A(n14716), .ZN(n14717) );
  OAI21_X1 U18034 ( .B1(n15983), .B2(n14747), .A(n14717), .ZN(P1_U2854) );
  AOI22_X1 U18035 ( .A1(n16125), .A2(n14719), .B1(P1_EBX_REG_17__SCAN_IN), 
        .B2(n14718), .ZN(n14720) );
  OAI21_X1 U18036 ( .B1(n14905), .B2(n14747), .A(n14720), .ZN(P1_U2855) );
  AOI21_X1 U18037 ( .B1(n14722), .B2(n14721), .A(n14624), .ZN(n16058) );
  INV_X1 U18038 ( .A(n16058), .ZN(n14808) );
  OR2_X1 U18039 ( .A1(n14735), .A2(n14723), .ZN(n14724) );
  NAND2_X1 U18040 ( .A1(n14725), .A2(n14724), .ZN(n15995) );
  OAI22_X1 U18041 ( .A1(n15995), .A2(n14749), .B1(n14726), .B2(n14748), .ZN(
        n14727) );
  INV_X1 U18042 ( .A(n14727), .ZN(n14728) );
  OAI21_X1 U18043 ( .B1(n14808), .B2(n14747), .A(n14728), .ZN(P1_U2856) );
  NAND2_X1 U18044 ( .A1(n14730), .A2(n14729), .ZN(n14731) );
  AND2_X1 U18045 ( .A1(n14721), .A2(n14731), .ZN(n16001) );
  INV_X1 U18046 ( .A(P1_EBX_REG_15__SCAN_IN), .ZN(n14736) );
  NOR2_X1 U18047 ( .A1(n14733), .A2(n14732), .ZN(n14734) );
  OR2_X1 U18048 ( .A1(n14735), .A2(n14734), .ZN(n15996) );
  OAI222_X1 U18049 ( .A1(n14747), .A2(n14811), .B1(n14748), .B2(n14736), .C1(
        n15996), .C2(n14749), .ZN(P1_U2857) );
  INV_X1 U18050 ( .A(n16146), .ZN(n14737) );
  OAI222_X1 U18051 ( .A1(n14738), .A2(n14748), .B1(n14747), .B2(n14933), .C1(
        n14749), .C2(n14737), .ZN(P1_U2859) );
  NAND2_X1 U18052 ( .A1(n14740), .A2(n14739), .ZN(n14741) );
  NAND2_X1 U18053 ( .A1(n14742), .A2(n14741), .ZN(n16160) );
  INV_X1 U18054 ( .A(P1_EBX_REG_12__SCAN_IN), .ZN(n16012) );
  NOR2_X1 U18055 ( .A1(n14744), .A2(n14743), .ZN(n14745) );
  NOR2_X1 U18056 ( .A1(n14746), .A2(n14745), .ZN(n16075) );
  INV_X1 U18057 ( .A(n16075), .ZN(n16018) );
  OAI222_X1 U18058 ( .A1(n16160), .A2(n14749), .B1(n14748), .B2(n16012), .C1(
        n14747), .C2(n16018), .ZN(P1_U2860) );
  INV_X1 U18059 ( .A(BUF1_REG_30__SCAN_IN), .ZN(n16467) );
  OAI22_X1 U18060 ( .A1(n14802), .A2(n16467), .B1(n13594), .B2(n20043), .ZN(
        n14751) );
  NOR2_X1 U18061 ( .A1(n14803), .A2(n20080), .ZN(n14750) );
  AOI211_X1 U18062 ( .C1(n14806), .C2(DATAI_30_), .A(n14751), .B(n14750), .ZN(
        n14752) );
  OAI21_X1 U18063 ( .B1(n14753), .B2(n14815), .A(n14752), .ZN(P1_U2874) );
  AOI22_X1 U18064 ( .A1(n14796), .A2(BUF1_REG_28__SCAN_IN), .B1(
        P1_EAX_REG_28__SCAN_IN), .B2(n14816), .ZN(n14757) );
  INV_X1 U18065 ( .A(DATAI_12_), .ZN(n14755) );
  NAND2_X1 U18066 ( .A1(n20160), .A2(BUF1_REG_12__SCAN_IN), .ZN(n14754) );
  OAI21_X1 U18067 ( .B1(n20160), .B2(n14755), .A(n14754), .ZN(n20078) );
  AOI22_X1 U18068 ( .A1(n14806), .A2(DATAI_28_), .B1(n14798), .B2(n20078), 
        .ZN(n14756) );
  OAI211_X1 U18069 ( .C1(n14758), .C2(n14815), .A(n14757), .B(n14756), .ZN(
        P1_U2876) );
  AOI22_X1 U18070 ( .A1(n14796), .A2(BUF1_REG_27__SCAN_IN), .B1(
        P1_EAX_REG_27__SCAN_IN), .B2(n14816), .ZN(n14761) );
  AOI22_X1 U18071 ( .A1(n14806), .A2(DATAI_27_), .B1(n14798), .B2(n14759), 
        .ZN(n14760) );
  OAI211_X1 U18072 ( .C1(n14842), .C2(n14815), .A(n14761), .B(n14760), .ZN(
        P1_U2877) );
  AOI22_X1 U18073 ( .A1(n14796), .A2(BUF1_REG_26__SCAN_IN), .B1(
        P1_EAX_REG_26__SCAN_IN), .B2(n14816), .ZN(n14764) );
  AOI22_X1 U18074 ( .A1(n14806), .A2(DATAI_26_), .B1(n14798), .B2(n14762), 
        .ZN(n14763) );
  OAI211_X1 U18075 ( .C1(n14765), .C2(n14815), .A(n14764), .B(n14763), .ZN(
        P1_U2878) );
  AOI22_X1 U18076 ( .A1(n14796), .A2(BUF1_REG_25__SCAN_IN), .B1(
        P1_EAX_REG_25__SCAN_IN), .B2(n14816), .ZN(n14769) );
  INV_X1 U18077 ( .A(DATAI_9_), .ZN(n14767) );
  NAND2_X1 U18078 ( .A1(n20160), .A2(BUF1_REG_9__SCAN_IN), .ZN(n14766) );
  OAI21_X1 U18079 ( .B1(n20160), .B2(n14767), .A(n14766), .ZN(n20076) );
  AOI22_X1 U18080 ( .A1(n14806), .A2(DATAI_25_), .B1(n14798), .B2(n20076), 
        .ZN(n14768) );
  OAI211_X1 U18081 ( .C1(n15928), .C2(n14815), .A(n14769), .B(n14768), .ZN(
        P1_U2879) );
  AOI22_X1 U18082 ( .A1(n14796), .A2(BUF1_REG_24__SCAN_IN), .B1(
        P1_EAX_REG_24__SCAN_IN), .B2(n14816), .ZN(n14772) );
  AOI22_X1 U18083 ( .A1(n14806), .A2(DATAI_24_), .B1(n14798), .B2(n14770), 
        .ZN(n14771) );
  OAI211_X1 U18084 ( .C1(n14864), .C2(n14815), .A(n14772), .B(n14771), .ZN(
        P1_U2880) );
  AOI22_X1 U18085 ( .A1(n14796), .A2(BUF1_REG_23__SCAN_IN), .B1(
        P1_EAX_REG_23__SCAN_IN), .B2(n14816), .ZN(n14775) );
  AOI22_X1 U18086 ( .A1(n14806), .A2(DATAI_23_), .B1(n14798), .B2(n14773), 
        .ZN(n14774) );
  OAI211_X1 U18087 ( .C1(n15948), .C2(n14815), .A(n14775), .B(n14774), .ZN(
        P1_U2881) );
  INV_X1 U18088 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n14776) );
  OAI22_X1 U18089 ( .A1(n14802), .A2(n14776), .B1(n13790), .B2(n20043), .ZN(
        n14778) );
  NOR2_X1 U18090 ( .A1(n14803), .A2(n20191), .ZN(n14777) );
  AOI211_X1 U18091 ( .C1(n14806), .C2(DATAI_22_), .A(n14778), .B(n14777), .ZN(
        n14779) );
  OAI21_X1 U18092 ( .B1(n15955), .B2(n14815), .A(n14779), .ZN(P1_U2882) );
  AOI22_X1 U18093 ( .A1(n14796), .A2(BUF1_REG_21__SCAN_IN), .B1(
        P1_EAX_REG_21__SCAN_IN), .B2(n14816), .ZN(n14782) );
  AOI22_X1 U18094 ( .A1(n14806), .A2(DATAI_21_), .B1(n14798), .B2(n14780), 
        .ZN(n14781) );
  OAI211_X1 U18095 ( .C1(n15967), .C2(n14815), .A(n14782), .B(n14781), .ZN(
        P1_U2883) );
  INV_X1 U18096 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n16484) );
  OAI22_X1 U18097 ( .A1(n14802), .A2(n16484), .B1(n13805), .B2(n20043), .ZN(
        n14784) );
  NOR2_X1 U18098 ( .A1(n14803), .A2(n20184), .ZN(n14783) );
  AOI211_X1 U18099 ( .C1(n14806), .C2(DATAI_20_), .A(n14784), .B(n14783), .ZN(
        n14785) );
  OAI21_X1 U18100 ( .B1(n14786), .B2(n14815), .A(n14785), .ZN(P1_U2884) );
  AOI22_X1 U18101 ( .A1(n14796), .A2(BUF1_REG_19__SCAN_IN), .B1(
        P1_EAX_REG_19__SCAN_IN), .B2(n14816), .ZN(n14789) );
  AOI22_X1 U18102 ( .A1(n14806), .A2(DATAI_19_), .B1(n14798), .B2(n14787), 
        .ZN(n14788) );
  OAI211_X1 U18103 ( .C1(n14885), .C2(n14815), .A(n14789), .B(n14788), .ZN(
        P1_U2885) );
  INV_X1 U18104 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n14790) );
  NOR2_X1 U18105 ( .A1(n14802), .A2(n14790), .ZN(n14794) );
  INV_X1 U18106 ( .A(n14806), .ZN(n14792) );
  INV_X1 U18107 ( .A(DATAI_18_), .ZN(n14791) );
  OAI22_X1 U18108 ( .A1(n14792), .A2(n14791), .B1(n20173), .B2(n14803), .ZN(
        n14793) );
  AOI211_X1 U18109 ( .C1(n14816), .C2(P1_EAX_REG_18__SCAN_IN), .A(n14794), .B(
        n14793), .ZN(n14795) );
  OAI21_X1 U18110 ( .B1(n15983), .B2(n14815), .A(n14795), .ZN(P1_U2886) );
  AOI22_X1 U18111 ( .A1(n14796), .A2(BUF1_REG_17__SCAN_IN), .B1(
        P1_EAX_REG_17__SCAN_IN), .B2(n14816), .ZN(n14800) );
  AOI22_X1 U18112 ( .A1(n14806), .A2(DATAI_17_), .B1(n14798), .B2(n14797), 
        .ZN(n14799) );
  OAI211_X1 U18113 ( .C1(n14905), .C2(n14815), .A(n14800), .B(n14799), .ZN(
        P1_U2887) );
  INV_X1 U18114 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n14801) );
  OAI22_X1 U18115 ( .A1(n14802), .A2(n14801), .B1(n13792), .B2(n20043), .ZN(
        n14805) );
  NOR2_X1 U18116 ( .A1(n14803), .A2(n20162), .ZN(n14804) );
  AOI211_X1 U18117 ( .C1(n14806), .C2(DATAI_16_), .A(n14805), .B(n14804), .ZN(
        n14807) );
  OAI21_X1 U18118 ( .B1(n14808), .B2(n14815), .A(n14807), .ZN(P1_U2888) );
  OAI222_X1 U18119 ( .A1(n14815), .A2(n14811), .B1(n14814), .B2(n14810), .C1(
        n20043), .C2(n14809), .ZN(P1_U2889) );
  INV_X1 U18120 ( .A(n14812), .ZN(n14813) );
  INV_X1 U18121 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n20971) );
  OAI222_X1 U18122 ( .A1(n14815), .A2(n14933), .B1(n14814), .B2(n14813), .C1(
        n20043), .C2(n20971), .ZN(P1_U2891) );
  AOI22_X1 U18123 ( .A1(n20039), .A2(n20078), .B1(P1_EAX_REG_12__SCAN_IN), 
        .B2(n14816), .ZN(n14817) );
  OAI21_X1 U18124 ( .B1(n16018), .B2(n14815), .A(n14817), .ZN(P1_U2892) );
  XNOR2_X1 U18125 ( .A(n14819), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14949) );
  NOR2_X1 U18126 ( .A1(n20128), .A2(n14820), .ZN(n14943) );
  AOI21_X1 U18127 ( .B1(n20091), .B2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n14943), .ZN(n14821) );
  OAI21_X1 U18128 ( .B1(n20102), .B2(n14822), .A(n14821), .ZN(n14823) );
  AOI21_X1 U18129 ( .B1(n14824), .B2(n20097), .A(n14823), .ZN(n14825) );
  OAI21_X1 U18130 ( .B1(n14949), .B2(n19949), .A(n14825), .ZN(P1_U2969) );
  NOR4_X1 U18131 ( .A1(n14826), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A4(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14827) );
  NAND2_X1 U18132 ( .A1(n16081), .A2(n14827), .ZN(n14830) );
  NAND3_X1 U18133 ( .A1(n9913), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14829) );
  NAND3_X1 U18134 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14981) );
  AOI21_X1 U18135 ( .B1(n9913), .B2(n14981), .A(n12652), .ZN(n14828) );
  MUX2_X1 U18136 ( .A(n14830), .B(n14829), .S(n14828), .Z(n14832) );
  XNOR2_X1 U18137 ( .A(n14832), .B(n14831), .ZN(n14971) );
  INV_X1 U18138 ( .A(P1_REIP_REG_28__SCAN_IN), .ZN(n20753) );
  NOR2_X1 U18139 ( .A1(n20128), .A2(n20753), .ZN(n14965) );
  AOI21_X1 U18140 ( .B1(n20091), .B2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n14965), .ZN(n14833) );
  OAI21_X1 U18141 ( .B1(n20102), .B2(n14834), .A(n14833), .ZN(n14835) );
  AOI21_X1 U18142 ( .B1(n14836), .B2(n20097), .A(n14835), .ZN(n14837) );
  OAI21_X1 U18143 ( .B1(n14971), .B2(n19949), .A(n14837), .ZN(P1_U2971) );
  XNOR2_X1 U18144 ( .A(n14841), .B(n14840), .ZN(n14979) );
  NAND2_X1 U18145 ( .A1(n20103), .A2(P1_REIP_REG_27__SCAN_IN), .ZN(n14973) );
  OAI21_X1 U18146 ( .B1(n14900), .B2(n21108), .A(n14973), .ZN(n14844) );
  NOR2_X1 U18147 ( .A1(n14842), .A2(n20159), .ZN(n14843) );
  AOI211_X1 U18148 ( .C1(n16077), .C2(n14845), .A(n14844), .B(n14843), .ZN(
        n14846) );
  OAI21_X1 U18149 ( .B1(n19949), .B2(n14979), .A(n14846), .ZN(P1_U2972) );
  OAI21_X1 U18150 ( .B1(n12652), .B2(n14981), .A(n9913), .ZN(n14847) );
  NAND2_X1 U18151 ( .A1(n14848), .A2(n14847), .ZN(n14849) );
  XNOR2_X1 U18152 ( .A(n14849), .B(n21089), .ZN(n14991) );
  INV_X1 U18153 ( .A(P1_REIP_REG_26__SCAN_IN), .ZN(n20747) );
  NOR2_X1 U18154 ( .A1(n20128), .A2(n20747), .ZN(n14983) );
  AOI21_X1 U18155 ( .B1(n20091), .B2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n14983), .ZN(n14850) );
  OAI21_X1 U18156 ( .B1(n20102), .B2(n14851), .A(n14850), .ZN(n14852) );
  AOI21_X1 U18157 ( .B1(n14853), .B2(n20097), .A(n14852), .ZN(n14854) );
  OAI21_X1 U18158 ( .B1(n19949), .B2(n14991), .A(n14854), .ZN(P1_U2973) );
  MUX2_X1 U18159 ( .A(n14999), .B(n14856), .S(n16081), .Z(n14857) );
  AOI21_X1 U18160 ( .B1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n14855), .A(
        n14857), .ZN(n14858) );
  XNOR2_X1 U18161 ( .A(n14858), .B(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14997) );
  INV_X1 U18162 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n15929) );
  OR2_X1 U18163 ( .A1(n20128), .A2(n15929), .ZN(n14993) );
  OAI21_X1 U18164 ( .B1(n14900), .B2(n15924), .A(n14993), .ZN(n14860) );
  NOR2_X1 U18165 ( .A1(n15928), .A2(n20159), .ZN(n14859) );
  AOI211_X1 U18166 ( .C1(n16077), .C2(n15927), .A(n14860), .B(n14859), .ZN(
        n14861) );
  OAI21_X1 U18167 ( .B1(n19949), .B2(n14997), .A(n14861), .ZN(P1_U2974) );
  NAND2_X1 U18168 ( .A1(n14855), .A2(n12652), .ZN(n14862) );
  MUX2_X1 U18169 ( .A(n14855), .B(n14862), .S(n16081), .Z(n14863) );
  XNOR2_X1 U18170 ( .A(n14863), .B(n14999), .ZN(n15006) );
  INV_X1 U18171 ( .A(n14864), .ZN(n15942) );
  NAND2_X1 U18172 ( .A1(n20103), .A2(P1_REIP_REG_24__SCAN_IN), .ZN(n15001) );
  NAND2_X1 U18173 ( .A1(n20091), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14865) );
  OAI211_X1 U18174 ( .C1(n20102), .C2(n15937), .A(n15001), .B(n14865), .ZN(
        n14866) );
  AOI21_X1 U18175 ( .B1(n15942), .B2(n20097), .A(n14866), .ZN(n14867) );
  OAI21_X1 U18176 ( .B1(n19949), .B2(n15006), .A(n14867), .ZN(P1_U2975) );
  XNOR2_X1 U18177 ( .A(n9913), .B(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14868) );
  XNOR2_X1 U18178 ( .A(n14869), .B(n14868), .ZN(n15013) );
  NAND2_X1 U18179 ( .A1(n20103), .A2(P1_REIP_REG_23__SCAN_IN), .ZN(n15007) );
  OAI21_X1 U18180 ( .B1(n14900), .B2(n15954), .A(n15007), .ZN(n14871) );
  NOR2_X1 U18181 ( .A1(n15948), .A2(n20159), .ZN(n14870) );
  AOI211_X1 U18182 ( .C1(n16077), .C2(n15945), .A(n14871), .B(n14870), .ZN(
        n14872) );
  OAI21_X1 U18183 ( .B1(n15013), .B2(n19949), .A(n14872), .ZN(P1_U2976) );
  AND2_X1 U18184 ( .A1(n9913), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n14883) );
  NAND2_X1 U18185 ( .A1(n16051), .A2(n14883), .ZN(n15032) );
  INV_X1 U18186 ( .A(n15032), .ZN(n14874) );
  AOI22_X1 U18187 ( .A1(n14874), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .B1(
        n16081), .B2(n14873), .ZN(n14875) );
  XNOR2_X1 U18188 ( .A(n14875), .B(n15025), .ZN(n15031) );
  NAND2_X1 U18189 ( .A1(n15965), .A2(n16077), .ZN(n14876) );
  NAND2_X1 U18190 ( .A1(n20103), .A2(P1_REIP_REG_21__SCAN_IN), .ZN(n15023) );
  OAI211_X1 U18191 ( .C1(n14900), .C2(n15972), .A(n14876), .B(n15023), .ZN(
        n14877) );
  AOI21_X1 U18192 ( .B1(n14878), .B2(n20097), .A(n14877), .ZN(n14879) );
  OAI21_X1 U18193 ( .B1(n15031), .B2(n19949), .A(n14879), .ZN(P1_U2978) );
  AOI21_X1 U18194 ( .B1(n16081), .B2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n16051), .ZN(n14884) );
  NOR2_X1 U18195 ( .A1(n9913), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n14880) );
  NAND2_X1 U18196 ( .A1(n14884), .A2(n14880), .ZN(n15033) );
  INV_X1 U18197 ( .A(n15033), .ZN(n14882) );
  NOR3_X1 U18198 ( .A1(n14884), .A2(n14883), .A3(n14880), .ZN(n14881) );
  AOI211_X1 U18199 ( .C1(n14884), .C2(n14883), .A(n14882), .B(n14881), .ZN(
        n16104) );
  INV_X1 U18200 ( .A(n14885), .ZN(n14889) );
  AOI22_X1 U18201 ( .A1(n20091), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B1(
        n20103), .B2(P1_REIP_REG_19__SCAN_IN), .ZN(n14886) );
  OAI21_X1 U18202 ( .B1(n20102), .B2(n14887), .A(n14886), .ZN(n14888) );
  AOI21_X1 U18203 ( .B1(n14889), .B2(n20097), .A(n14888), .ZN(n14890) );
  OAI21_X1 U18204 ( .B1(n16104), .B2(n19949), .A(n14890), .ZN(P1_U2980) );
  INV_X1 U18205 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n21021) );
  NAND2_X1 U18206 ( .A1(n14891), .A2(n14907), .ZN(n16065) );
  INV_X1 U18207 ( .A(n14892), .ZN(n14895) );
  INV_X1 U18208 ( .A(n14893), .ZN(n14894) );
  OAI21_X1 U18209 ( .B1(n16065), .B2(n14895), .A(n14894), .ZN(n14896) );
  NAND2_X1 U18210 ( .A1(n16081), .A2(n14896), .ZN(n14897) );
  OAI22_X1 U18211 ( .A1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n14897), .B1(
        n16081), .B2(n14896), .ZN(n14898) );
  XNOR2_X1 U18212 ( .A(n21021), .B(n14898), .ZN(n16126) );
  NAND2_X1 U18213 ( .A1(n16126), .A2(n20098), .ZN(n14904) );
  INV_X1 U18214 ( .A(P1_REIP_REG_17__SCAN_IN), .ZN(n14899) );
  OAI22_X1 U18215 ( .A1(n14900), .A2(n14633), .B1(n20128), .B2(n14899), .ZN(
        n14901) );
  AOI21_X1 U18216 ( .B1(n16077), .B2(n14902), .A(n14901), .ZN(n14903) );
  OAI211_X1 U18217 ( .C1(n20159), .C2(n14905), .A(n14904), .B(n14903), .ZN(
        P1_U2982) );
  INV_X1 U18218 ( .A(n14891), .ZN(n14910) );
  INV_X1 U18219 ( .A(n14906), .ZN(n14909) );
  OAI211_X1 U18220 ( .C1(n9913), .C2(n16143), .A(n14907), .B(n16062), .ZN(
        n14908) );
  AOI21_X1 U18221 ( .B1(n14910), .B2(n14909), .A(n14908), .ZN(n14914) );
  AND2_X1 U18222 ( .A1(n14914), .A2(n14911), .ZN(n15044) );
  INV_X1 U18223 ( .A(n15044), .ZN(n14915) );
  INV_X1 U18224 ( .A(n14911), .ZN(n14912) );
  NOR2_X1 U18225 ( .A1(n15043), .A2(n14912), .ZN(n14913) );
  OAI22_X1 U18226 ( .A1(n14915), .A2(n15043), .B1(n14914), .B2(n14913), .ZN(
        n16133) );
  INV_X1 U18227 ( .A(n16133), .ZN(n14920) );
  AOI22_X1 U18228 ( .A1(n20091), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B1(
        n20103), .B2(P1_REIP_REG_15__SCAN_IN), .ZN(n14916) );
  OAI21_X1 U18229 ( .B1(n20102), .B2(n14917), .A(n14916), .ZN(n14918) );
  AOI21_X1 U18230 ( .B1(n16001), .B2(n20097), .A(n14918), .ZN(n14919) );
  OAI21_X1 U18231 ( .B1(n14920), .B2(n19949), .A(n14919), .ZN(P1_U2984) );
  OAI21_X1 U18232 ( .B1(n14891), .B2(n14922), .A(n14921), .ZN(n16074) );
  INV_X1 U18233 ( .A(n14925), .ZN(n14924) );
  NAND2_X1 U18234 ( .A1(n14924), .A2(n14923), .ZN(n16073) );
  NOR2_X1 U18235 ( .A1(n16074), .A2(n16073), .ZN(n16072) );
  NOR2_X1 U18236 ( .A1(n16072), .A2(n14925), .ZN(n14927) );
  XNOR2_X1 U18237 ( .A(n14927), .B(n14926), .ZN(n16147) );
  NAND2_X1 U18238 ( .A1(n16147), .A2(n20098), .ZN(n14932) );
  INV_X1 U18239 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n14928) );
  NOR2_X1 U18240 ( .A1(n20128), .A2(n14928), .ZN(n16145) );
  NOR2_X1 U18241 ( .A1(n20102), .A2(n14929), .ZN(n14930) );
  AOI211_X1 U18242 ( .C1(n20091), .C2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .A(
        n16145), .B(n14930), .ZN(n14931) );
  OAI211_X1 U18243 ( .C1(n20159), .C2(n14933), .A(n14932), .B(n14931), .ZN(
        P1_U2986) );
  AND2_X1 U18244 ( .A1(n14934), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n14936) );
  XNOR2_X1 U18245 ( .A(n14891), .B(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n14935) );
  MUX2_X1 U18246 ( .A(n14936), .B(n14935), .S(n9913), .Z(n14937) );
  NOR3_X1 U18247 ( .A1(n14934), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(
        n9913), .ZN(n16082) );
  NOR2_X1 U18248 ( .A1(n14937), .A2(n16082), .ZN(n15068) );
  INV_X1 U18249 ( .A(P1_REIP_REG_10__SCAN_IN), .ZN(n14938) );
  NOR2_X1 U18250 ( .A1(n20128), .A2(n14938), .ZN(n15065) );
  AOI21_X1 U18251 ( .B1(n20091), .B2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n15065), .ZN(n14939) );
  OAI21_X1 U18252 ( .B1(n20102), .B2(n16033), .A(n14939), .ZN(n14940) );
  AOI21_X1 U18253 ( .B1(n16035), .B2(n20097), .A(n14940), .ZN(n14941) );
  OAI21_X1 U18254 ( .B1(n15068), .B2(n19949), .A(n14941), .ZN(P1_U2989) );
  INV_X1 U18255 ( .A(n14942), .ZN(n14944) );
  AOI21_X1 U18256 ( .B1(n14944), .B2(n20114), .A(n14943), .ZN(n14948) );
  OAI21_X1 U18257 ( .B1(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n14946), .A(
        n14945), .ZN(n14947) );
  OAI211_X1 U18258 ( .C1(n14949), .C2(n16177), .A(n14948), .B(n14947), .ZN(
        P1_U3001) );
  INV_X1 U18259 ( .A(n14950), .ZN(n14957) );
  NOR3_X1 U18260 ( .A1(n14975), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n14951), .ZN(n14956) );
  INV_X1 U18261 ( .A(n14952), .ZN(n14954) );
  OAI21_X1 U18262 ( .B1(n14954), .B2(n20145), .A(n14953), .ZN(n14955) );
  AOI211_X1 U18263 ( .C1(n14957), .C2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n14956), .B(n14955), .ZN(n14958) );
  OAI21_X1 U18264 ( .B1(n14959), .B2(n16177), .A(n14958), .ZN(P1_U3002) );
  INV_X1 U18265 ( .A(n14960), .ZN(n14966) );
  INV_X1 U18266 ( .A(n14961), .ZN(n14962) );
  NOR3_X1 U18267 ( .A1(n14975), .A2(n14963), .A3(n14962), .ZN(n14964) );
  AOI211_X1 U18268 ( .C1(n14966), .C2(n20114), .A(n14965), .B(n14964), .ZN(
        n14970) );
  AND2_X1 U18269 ( .A1(n14968), .A2(n14967), .ZN(n14977) );
  NAND2_X1 U18270 ( .A1(n14977), .A2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14969) );
  OAI211_X1 U18271 ( .C1(n14971), .C2(n16177), .A(n14970), .B(n14969), .ZN(
        P1_U3003) );
  NAND2_X1 U18272 ( .A1(n14972), .A2(n20114), .ZN(n14974) );
  OAI211_X1 U18273 ( .C1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n14975), .A(
        n14974), .B(n14973), .ZN(n14976) );
  AOI21_X1 U18274 ( .B1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n14977), .A(
        n14976), .ZN(n14978) );
  OAI21_X1 U18275 ( .B1(n14979), .B2(n16177), .A(n14978), .ZN(P1_U3004) );
  INV_X1 U18276 ( .A(n14980), .ZN(n14984) );
  INV_X1 U18277 ( .A(n15000), .ZN(n15008) );
  NOR3_X1 U18278 ( .A1(n15008), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        n14981), .ZN(n14982) );
  AOI211_X1 U18279 ( .C1(n20114), .C2(n14984), .A(n14983), .B(n14982), .ZN(
        n14990) );
  AND2_X1 U18280 ( .A1(n14986), .A2(n14985), .ZN(n14987) );
  NAND2_X1 U18281 ( .A1(n15000), .A2(n14987), .ZN(n14992) );
  INV_X1 U18282 ( .A(n14992), .ZN(n14988) );
  OAI21_X1 U18283 ( .B1(n14988), .B2(n14995), .A(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n14989) );
  OAI211_X1 U18284 ( .C1(n14991), .C2(n16177), .A(n14990), .B(n14989), .ZN(
        P1_U3005) );
  OAI211_X1 U18285 ( .C1(n15934), .C2(n20145), .A(n14993), .B(n14992), .ZN(
        n14994) );
  AOI21_X1 U18286 ( .B1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n14995), .A(
        n14994), .ZN(n14996) );
  OAI21_X1 U18287 ( .B1(n14997), .B2(n16177), .A(n14996), .ZN(P1_U3006) );
  OAI21_X1 U18288 ( .B1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n20120), .A(
        n14998), .ZN(n15004) );
  NAND3_X1 U18289 ( .A1(n15000), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        n14999), .ZN(n15002) );
  OAI211_X1 U18290 ( .C1(n20145), .C2(n15944), .A(n15002), .B(n15001), .ZN(
        n15003) );
  AOI21_X1 U18291 ( .B1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n15004), .A(
        n15003), .ZN(n15005) );
  OAI21_X1 U18292 ( .B1(n15006), .B2(n16177), .A(n15005), .ZN(P1_U3007) );
  OAI21_X1 U18293 ( .B1(n15947), .B2(n20145), .A(n15007), .ZN(n15010) );
  NOR2_X1 U18294 ( .A1(n15008), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15009) );
  AOI211_X1 U18295 ( .C1(n15011), .C2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n15010), .B(n15009), .ZN(n15012) );
  OAI21_X1 U18296 ( .B1(n15013), .B2(n16177), .A(n15012), .ZN(P1_U3008) );
  NAND2_X1 U18297 ( .A1(n15015), .A2(n15014), .ZN(n15016) );
  XNOR2_X1 U18298 ( .A(n15016), .B(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n16039) );
  INV_X1 U18299 ( .A(n16039), .ZN(n15022) );
  INV_X1 U18300 ( .A(n15964), .ZN(n15020) );
  INV_X1 U18301 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n20741) );
  OAI22_X1 U18302 ( .A1(n21070), .A2(n15026), .B1(n20128), .B2(n20741), .ZN(
        n15019) );
  INV_X1 U18303 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n16109) );
  NOR2_X1 U18304 ( .A1(n16109), .A2(n16108), .ZN(n15037) );
  NAND2_X1 U18305 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n15037), .ZN(
        n15024) );
  AOI211_X1 U18306 ( .C1(n15025), .C2(n21070), .A(n15017), .B(n15024), .ZN(
        n15018) );
  AOI211_X1 U18307 ( .C1(n20114), .C2(n15020), .A(n15019), .B(n15018), .ZN(
        n15021) );
  OAI21_X1 U18308 ( .B1(n15022), .B2(n16177), .A(n15021), .ZN(P1_U3009) );
  OAI21_X1 U18309 ( .B1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .B2(n15024), .A(
        n15023), .ZN(n15028) );
  NOR2_X1 U18310 ( .A1(n15026), .A2(n15025), .ZN(n15027) );
  AOI211_X1 U18311 ( .C1(n20114), .C2(n15029), .A(n15028), .B(n15027), .ZN(
        n15030) );
  OAI21_X1 U18312 ( .B1(n15031), .B2(n16177), .A(n15030), .ZN(P1_U3010) );
  NAND2_X1 U18313 ( .A1(n15033), .A2(n15032), .ZN(n15035) );
  XNOR2_X1 U18314 ( .A(n15035), .B(n15034), .ZN(n16045) );
  INV_X1 U18315 ( .A(n16045), .ZN(n15042) );
  INV_X1 U18316 ( .A(n16111), .ZN(n15036) );
  OAI21_X1 U18317 ( .B1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n16108), .A(
        n15036), .ZN(n15040) );
  AOI22_X1 U18318 ( .A1(n20103), .A2(P1_REIP_REG_20__SCAN_IN), .B1(n15034), 
        .B2(n15037), .ZN(n15038) );
  OAI21_X1 U18319 ( .B1(n15980), .B2(n20145), .A(n15038), .ZN(n15039) );
  AOI21_X1 U18320 ( .B1(n15040), .B2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n15039), .ZN(n15041) );
  OAI21_X1 U18321 ( .B1(n15042), .B2(n16177), .A(n15041), .ZN(P1_U3011) );
  NOR2_X1 U18322 ( .A1(n15044), .A2(n15043), .ZN(n15045) );
  XNOR2_X1 U18323 ( .A(n15046), .B(n15045), .ZN(n16057) );
  INV_X1 U18324 ( .A(n16057), .ZN(n15059) );
  NAND2_X1 U18325 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n16140), .ZN(
        n16136) );
  AOI221_X1 U18326 ( .B1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .C1(n15048), .C2(n15047), .A(
        n16136), .ZN(n15049) );
  INV_X1 U18327 ( .A(n15049), .ZN(n15058) );
  AOI21_X1 U18328 ( .B1(n15051), .B2(n15050), .A(n20123), .ZN(n15052) );
  OAI21_X1 U18329 ( .B1(n15054), .B2(n15053), .A(n15052), .ZN(n16148) );
  INV_X1 U18330 ( .A(n16148), .ZN(n16144) );
  OAI21_X1 U18331 ( .B1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n16115), .A(
        n16144), .ZN(n16131) );
  INV_X1 U18332 ( .A(P1_REIP_REG_16__SCAN_IN), .ZN(n15055) );
  OAI22_X1 U18333 ( .A1(n15995), .A2(n20145), .B1(n20128), .B2(n15055), .ZN(
        n15056) );
  AOI21_X1 U18334 ( .B1(n16131), .B2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n15056), .ZN(n15057) );
  OAI211_X1 U18335 ( .C1(n15059), .C2(n16177), .A(n15058), .B(n15057), .ZN(
        P1_U3015) );
  INV_X1 U18336 ( .A(n16028), .ZN(n15066) );
  INV_X1 U18337 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16080) );
  INV_X1 U18338 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15061) );
  OAI221_X1 U18339 ( .B1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .C1(n16080), .C2(n15061), .A(
        n15060), .ZN(n15062) );
  OAI22_X1 U18340 ( .A1(n16080), .A2(n15063), .B1(n16180), .B2(n15062), .ZN(
        n15064) );
  AOI211_X1 U18341 ( .C1(n20114), .C2(n15066), .A(n15065), .B(n15064), .ZN(
        n15067) );
  OAI21_X1 U18342 ( .B1(n15068), .B2(n16177), .A(n15067), .ZN(P1_U3021) );
  NOR2_X1 U18343 ( .A1(n10291), .A2(n13716), .ZN(n15077) );
  NOR2_X1 U18344 ( .A1(n20529), .A2(n15069), .ZN(n15070) );
  AOI211_X1 U18345 ( .C1(n15072), .C2(n15077), .A(n15071), .B(n15070), .ZN(
        n15869) );
  INV_X1 U18346 ( .A(n15073), .ZN(n15080) );
  INV_X1 U18347 ( .A(n15074), .ZN(n15075) );
  AOI22_X1 U18348 ( .A1(n15078), .A2(n15077), .B1(n15076), .B2(n15075), .ZN(
        n15079) );
  OAI21_X1 U18349 ( .B1(n15869), .B2(n15080), .A(n15079), .ZN(n15082) );
  MUX2_X1 U18350 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n15082), .S(
        n15081), .Z(P1_U3473) );
  INV_X1 U18351 ( .A(n15083), .ZN(n15086) );
  INV_X1 U18352 ( .A(n15084), .ZN(n15085) );
  OAI211_X1 U18353 ( .C1(n15086), .C2(n15289), .A(n15085), .B(n9868), .ZN(
        n15093) );
  NAND2_X1 U18354 ( .A1(n15237), .A2(n19088), .ZN(n15088) );
  AOI22_X1 U18355 ( .A1(P2_REIP_REG_29__SCAN_IN), .A2(n19091), .B1(
        P2_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n19101), .ZN(n15087) );
  OAI211_X1 U18356 ( .C1(n19072), .C2(n15089), .A(n15088), .B(n15087), .ZN(
        n15090) );
  AOI21_X1 U18357 ( .B1(n15091), .B2(n19049), .A(n15090), .ZN(n15092) );
  OAI211_X1 U18358 ( .C1(n19067), .C2(n15293), .A(n15093), .B(n15092), .ZN(
        P2_U2826) );
  NAND2_X1 U18359 ( .A1(n15095), .A2(n15094), .ZN(n15096) );
  NAND2_X1 U18360 ( .A1(n15097), .A2(n15096), .ZN(n15477) );
  INV_X1 U18361 ( .A(n15477), .ZN(n15243) );
  NAND2_X1 U18362 ( .A1(n19090), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n15099) );
  NAND2_X1 U18363 ( .A1(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n19101), .ZN(
        n15098) );
  OAI211_X1 U18364 ( .C1(n19074), .C2(n19869), .A(n15099), .B(n15098), .ZN(
        n15100) );
  AOI21_X1 U18365 ( .B1(n15243), .B2(n19088), .A(n15100), .ZN(n15101) );
  OAI21_X1 U18366 ( .B1(n15102), .B2(n19095), .A(n15101), .ZN(n15107) );
  AOI211_X1 U18367 ( .C1(n15105), .C2(n15104), .A(n15103), .B(n19809), .ZN(
        n15106) );
  AOI211_X1 U18368 ( .C1(n19097), .C2(n15108), .A(n15107), .B(n15106), .ZN(
        n15109) );
  INV_X1 U18369 ( .A(n15109), .ZN(P2_U2827) );
  XOR2_X1 U18370 ( .A(P2_EBX_REG_25__SCAN_IN), .B(n15110), .Z(n15123) );
  OR2_X1 U18371 ( .A1(n15112), .A2(n15113), .ZN(n15114) );
  NAND2_X1 U18372 ( .A1(n15111), .A2(n15114), .ZN(n15514) );
  AOI21_X1 U18373 ( .B1(n15115), .B2(n15129), .A(n15252), .ZN(n15511) );
  AOI22_X1 U18374 ( .A1(P2_EBX_REG_25__SCAN_IN), .A2(n19090), .B1(
        P2_REIP_REG_25__SCAN_IN), .B2(n19091), .ZN(n15116) );
  OAI21_X1 U18375 ( .B1(n19057), .B2(n15322), .A(n15116), .ZN(n15117) );
  AOI21_X1 U18376 ( .B1(n15511), .B2(n19088), .A(n15117), .ZN(n15118) );
  OAI21_X1 U18377 ( .B1(n15514), .B2(n19067), .A(n15118), .ZN(n15122) );
  AOI211_X1 U18378 ( .C1(n15120), .C2(n15324), .A(n19809), .B(n15119), .ZN(
        n15121) );
  AOI211_X1 U18379 ( .C1(n19049), .C2(n15123), .A(n15122), .B(n15121), .ZN(
        n15124) );
  INV_X1 U18380 ( .A(n15124), .ZN(P2_U2830) );
  AOI21_X1 U18381 ( .B1(n15126), .B2(n15125), .A(n15112), .ZN(n15337) );
  INV_X1 U18382 ( .A(n15337), .ZN(n15526) );
  NAND2_X1 U18383 ( .A1(n13362), .A2(n15127), .ZN(n15128) );
  NAND2_X1 U18384 ( .A1(n15129), .A2(n15128), .ZN(n15262) );
  AOI22_X1 U18385 ( .A1(P2_EBX_REG_24__SCAN_IN), .A2(n19090), .B1(
        P2_REIP_REG_24__SCAN_IN), .B2(n19091), .ZN(n15134) );
  INV_X1 U18386 ( .A(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n15130) );
  OAI22_X1 U18387 ( .A1(n15131), .A2(n19095), .B1(n15130), .B2(n19057), .ZN(
        n15132) );
  INV_X1 U18388 ( .A(n15132), .ZN(n15133) );
  OAI211_X1 U18389 ( .C1(n15262), .C2(n19087), .A(n15134), .B(n15133), .ZN(
        n15139) );
  AOI211_X1 U18390 ( .C1(n15137), .C2(n15136), .A(n15135), .B(n19809), .ZN(
        n15138) );
  NOR2_X1 U18391 ( .A1(n15139), .A2(n15138), .ZN(n15140) );
  OAI21_X1 U18392 ( .B1(n19067), .B2(n15526), .A(n15140), .ZN(P2_U2831) );
  INV_X1 U18393 ( .A(n18977), .ZN(n19002) );
  NAND2_X1 U18394 ( .A1(n16259), .A2(n15141), .ZN(n15142) );
  AOI22_X1 U18395 ( .A1(n16259), .A2(n19002), .B1(n15143), .B2(n15142), .ZN(
        n15155) );
  OAI22_X1 U18396 ( .A1(n15144), .A2(n19072), .B1(n16266), .B2(n19057), .ZN(
        n15145) );
  AOI211_X1 U18397 ( .C1(P2_REIP_REG_11__SCAN_IN), .C2(n19091), .A(n19038), 
        .B(n15145), .ZN(n15154) );
  OR2_X1 U18398 ( .A1(n15147), .A2(n15146), .ZN(n15148) );
  NAND2_X1 U18399 ( .A1(n15148), .A2(n14263), .ZN(n19128) );
  INV_X1 U18400 ( .A(n19128), .ZN(n15149) );
  AOI22_X1 U18401 ( .A1(n16263), .A2(n19097), .B1(n19088), .B2(n15149), .ZN(
        n15153) );
  INV_X1 U18402 ( .A(n12192), .ZN(n15150) );
  NAND3_X1 U18403 ( .A1(n15151), .A2(n15150), .A3(n19049), .ZN(n15152) );
  NAND4_X1 U18404 ( .A1(n15155), .A2(n15154), .A3(n15153), .A4(n15152), .ZN(
        P2_U2844) );
  NAND2_X1 U18405 ( .A1(n15156), .A2(n15212), .ZN(n15157) );
  OAI21_X1 U18406 ( .B1(n15212), .B2(n15158), .A(n15157), .ZN(P2_U2856) );
  INV_X1 U18407 ( .A(n15159), .ZN(n15162) );
  OR2_X1 U18408 ( .A1(n15161), .A2(n15160), .ZN(n15235) );
  NAND3_X1 U18409 ( .A1(n15162), .A2(n15231), .A3(n15235), .ZN(n15164) );
  NAND2_X1 U18410 ( .A1(n15234), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n15163) );
  OAI211_X1 U18411 ( .C1(n15234), .C2(n15293), .A(n15164), .B(n15163), .ZN(
        P2_U2858) );
  NOR2_X1 U18412 ( .A1(n12904), .A2(n15165), .ZN(n15167) );
  XNOR2_X1 U18413 ( .A(n15167), .B(n15166), .ZN(n15246) );
  NOR2_X1 U18414 ( .A1(n15472), .A2(n15192), .ZN(n15168) );
  AOI21_X1 U18415 ( .B1(P2_EBX_REG_28__SCAN_IN), .B2(n15192), .A(n15168), .ZN(
        n15169) );
  OAI21_X1 U18416 ( .B1(n15246), .B2(n15215), .A(n15169), .ZN(P2_U2859) );
  OAI21_X1 U18417 ( .B1(n15172), .B2(n15171), .A(n15170), .ZN(n15250) );
  NAND2_X1 U18418 ( .A1(n15234), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n15174) );
  NAND2_X1 U18419 ( .A1(n15485), .A2(n15212), .ZN(n15173) );
  OAI211_X1 U18420 ( .C1(n15250), .C2(n15215), .A(n15174), .B(n15173), .ZN(
        P2_U2860) );
  AOI21_X1 U18421 ( .B1(n15176), .B2(n15111), .A(n11593), .ZN(n16215) );
  INV_X1 U18422 ( .A(n16215), .ZN(n15182) );
  AOI21_X1 U18423 ( .B1(n15179), .B2(n15178), .A(n15177), .ZN(n15256) );
  NAND2_X1 U18424 ( .A1(n15256), .A2(n15231), .ZN(n15181) );
  NAND2_X1 U18425 ( .A1(n15234), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n15180) );
  OAI211_X1 U18426 ( .C1(n15182), .C2(n15234), .A(n15181), .B(n15180), .ZN(
        P2_U2861) );
  OAI21_X1 U18427 ( .B1(n15183), .B2(n15185), .A(n15184), .ZN(n15261) );
  NOR2_X1 U18428 ( .A1(n15514), .A2(n15192), .ZN(n15186) );
  AOI21_X1 U18429 ( .B1(P2_EBX_REG_25__SCAN_IN), .B2(n15234), .A(n15186), .ZN(
        n15187) );
  OAI21_X1 U18430 ( .B1(n15261), .B2(n15215), .A(n15187), .ZN(P2_U2862) );
  AOI21_X1 U18431 ( .B1(n15188), .B2(n15189), .A(n9925), .ZN(n15190) );
  XOR2_X1 U18432 ( .A(n15191), .B(n15190), .Z(n15267) );
  NOR2_X1 U18433 ( .A1(n15526), .A2(n15192), .ZN(n15193) );
  AOI21_X1 U18434 ( .B1(P2_EBX_REG_24__SCAN_IN), .B2(n15234), .A(n15193), .ZN(
        n15194) );
  OAI21_X1 U18435 ( .B1(n15267), .B2(n15215), .A(n15194), .ZN(P2_U2863) );
  AOI21_X1 U18436 ( .B1(n15195), .B2(n15197), .A(n15196), .ZN(n15272) );
  NAND2_X1 U18437 ( .A1(n15272), .A2(n15231), .ZN(n15199) );
  INV_X1 U18438 ( .A(n15347), .ZN(n15540) );
  NAND2_X1 U18439 ( .A1(n15540), .A2(n15212), .ZN(n15198) );
  OAI211_X1 U18440 ( .C1(n15212), .C2(n11753), .A(n15199), .B(n15198), .ZN(
        P2_U2864) );
  NAND2_X1 U18441 ( .A1(n15201), .A2(n15200), .ZN(n15202) );
  AND2_X1 U18442 ( .A1(n15203), .A2(n15202), .ZN(n15856) );
  INV_X1 U18443 ( .A(n15856), .ZN(n15209) );
  NAND2_X1 U18444 ( .A1(n15229), .A2(n15204), .ZN(n15210) );
  AOI21_X1 U18445 ( .B1(n15206), .B2(n15210), .A(n15205), .ZN(n16226) );
  NAND2_X1 U18446 ( .A1(n16226), .A2(n15231), .ZN(n15208) );
  NAND2_X1 U18447 ( .A1(n15234), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n15207) );
  OAI211_X1 U18448 ( .C1(n15209), .C2(n15234), .A(n15208), .B(n15207), .ZN(
        P2_U2865) );
  AND2_X1 U18449 ( .A1(n15229), .A2(n15220), .ZN(n15221) );
  OAI21_X1 U18450 ( .B1(n15221), .B2(n15211), .A(n15210), .ZN(n15279) );
  MUX2_X1 U18451 ( .A(n15213), .B(n15560), .S(n15212), .Z(n15214) );
  OAI21_X1 U18452 ( .B1(n15279), .B2(n15215), .A(n15214), .ZN(P2_U2866) );
  NOR2_X1 U18453 ( .A1(n15216), .A2(n15217), .ZN(n15218) );
  OR2_X1 U18454 ( .A1(n15219), .A2(n15218), .ZN(n18948) );
  INV_X1 U18455 ( .A(n15220), .ZN(n15223) );
  INV_X1 U18456 ( .A(n15229), .ZN(n15222) );
  AOI21_X1 U18457 ( .B1(n15223), .B2(n15222), .A(n15221), .ZN(n16230) );
  NAND2_X1 U18458 ( .A1(n16230), .A2(n15231), .ZN(n15225) );
  NAND2_X1 U18459 ( .A1(n15234), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n15224) );
  OAI211_X1 U18460 ( .C1(n18948), .C2(n15234), .A(n15225), .B(n15224), .ZN(
        P2_U2867) );
  AND2_X1 U18461 ( .A1(n15227), .A2(n15226), .ZN(n15228) );
  OR2_X1 U18462 ( .A1(n15228), .A2(n15216), .ZN(n18957) );
  AOI21_X1 U18463 ( .B1(n15230), .B2(n10173), .A(n15229), .ZN(n15287) );
  NAND2_X1 U18464 ( .A1(n15287), .A2(n15231), .ZN(n15233) );
  NAND2_X1 U18465 ( .A1(n15234), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n15232) );
  OAI211_X1 U18466 ( .C1(n18957), .C2(n15234), .A(n15233), .B(n15232), .ZN(
        P2_U2868) );
  NAND2_X1 U18467 ( .A1(n15235), .A2(n19116), .ZN(n15240) );
  INV_X1 U18468 ( .A(n19108), .ZN(n15263) );
  INV_X1 U18469 ( .A(P2_EAX_REG_29__SCAN_IN), .ZN(n19176) );
  OAI22_X1 U18470 ( .A1(n15263), .A2(n19122), .B1(n19140), .B2(n19176), .ZN(
        n15236) );
  AOI21_X1 U18471 ( .B1(n19156), .B2(n15237), .A(n15236), .ZN(n15239) );
  AOI22_X1 U18472 ( .A1(n19110), .A2(BUF1_REG_29__SCAN_IN), .B1(n19109), .B2(
        BUF2_REG_29__SCAN_IN), .ZN(n15238) );
  OAI211_X1 U18473 ( .C1(n15240), .C2(n15159), .A(n15239), .B(n15238), .ZN(
        P2_U2890) );
  INV_X1 U18474 ( .A(n19124), .ZN(n15241) );
  OAI22_X1 U18475 ( .A1(n15263), .A2(n15241), .B1(n19140), .B2(n19178), .ZN(
        n15242) );
  AOI21_X1 U18476 ( .B1(n19156), .B2(n15243), .A(n15242), .ZN(n15245) );
  AOI22_X1 U18477 ( .A1(n19110), .A2(BUF1_REG_28__SCAN_IN), .B1(n19109), .B2(
        BUF2_REG_28__SCAN_IN), .ZN(n15244) );
  OAI211_X1 U18478 ( .C1(n15246), .C2(n19160), .A(n15245), .B(n15244), .ZN(
        P2_U2891) );
  INV_X1 U18479 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n19180) );
  OAI22_X1 U18480 ( .A1(n15263), .A2(n19127), .B1(n19140), .B2(n19180), .ZN(
        n15247) );
  AOI21_X1 U18481 ( .B1(n19156), .B2(n15486), .A(n15247), .ZN(n15249) );
  AOI22_X1 U18482 ( .A1(n19110), .A2(BUF1_REG_27__SCAN_IN), .B1(n19109), .B2(
        BUF2_REG_27__SCAN_IN), .ZN(n15248) );
  OAI211_X1 U18483 ( .C1(n15250), .C2(n19160), .A(n15249), .B(n15248), .ZN(
        P2_U2892) );
  OAI21_X1 U18484 ( .B1(n15252), .B2(n15251), .A(n13336), .ZN(n16213) );
  AOI22_X1 U18485 ( .A1(n19110), .A2(BUF1_REG_26__SCAN_IN), .B1(n19109), .B2(
        BUF2_REG_26__SCAN_IN), .ZN(n15254) );
  AOI22_X1 U18486 ( .A1(n19108), .A2(n19130), .B1(n19155), .B2(
        P2_EAX_REG_26__SCAN_IN), .ZN(n15253) );
  OAI211_X1 U18487 ( .C1(n15285), .C2(n16213), .A(n15254), .B(n15253), .ZN(
        n15255) );
  AOI21_X1 U18488 ( .B1(n15256), .B2(n19116), .A(n15255), .ZN(n15257) );
  INV_X1 U18489 ( .A(n15257), .ZN(P2_U2893) );
  INV_X1 U18490 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n19184) );
  OAI22_X1 U18491 ( .A1(n15263), .A2(n19133), .B1(n19140), .B2(n19184), .ZN(
        n15258) );
  AOI21_X1 U18492 ( .B1(n19156), .B2(n15511), .A(n15258), .ZN(n15260) );
  AOI22_X1 U18493 ( .A1(n19110), .A2(BUF1_REG_25__SCAN_IN), .B1(n19109), .B2(
        BUF2_REG_25__SCAN_IN), .ZN(n15259) );
  OAI211_X1 U18494 ( .C1(n15261), .C2(n19160), .A(n15260), .B(n15259), .ZN(
        P2_U2894) );
  INV_X1 U18495 ( .A(n15262), .ZN(n15524) );
  INV_X1 U18496 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n19186) );
  OAI22_X1 U18497 ( .A1(n15263), .A2(n19136), .B1(n19140), .B2(n19186), .ZN(
        n15264) );
  AOI21_X1 U18498 ( .B1(n19156), .B2(n15524), .A(n15264), .ZN(n15266) );
  AOI22_X1 U18499 ( .A1(n19110), .A2(BUF1_REG_24__SCAN_IN), .B1(n19109), .B2(
        BUF2_REG_24__SCAN_IN), .ZN(n15265) );
  OAI211_X1 U18500 ( .C1(n15267), .C2(n19160), .A(n15266), .B(n15265), .ZN(
        P2_U2895) );
  AOI22_X1 U18501 ( .A1(n19110), .A2(BUF1_REG_23__SCAN_IN), .B1(n19109), .B2(
        BUF2_REG_23__SCAN_IN), .ZN(n15270) );
  AOI22_X1 U18502 ( .A1(n19108), .A2(n15268), .B1(n19155), .B2(
        P2_EAX_REG_23__SCAN_IN), .ZN(n15269) );
  OAI211_X1 U18503 ( .C1(n15285), .C2(n15537), .A(n15270), .B(n15269), .ZN(
        n15271) );
  AOI21_X1 U18504 ( .B1(n15272), .B2(n19116), .A(n15271), .ZN(n15273) );
  INV_X1 U18505 ( .A(n15273), .ZN(P2_U2896) );
  AOI22_X1 U18506 ( .A1(n19110), .A2(BUF1_REG_21__SCAN_IN), .B1(n19109), .B2(
        BUF2_REG_21__SCAN_IN), .ZN(n15276) );
  AOI22_X1 U18507 ( .A1(n19108), .A2(n15274), .B1(n19155), .B2(
        P2_EAX_REG_21__SCAN_IN), .ZN(n15275) );
  OAI211_X1 U18508 ( .C1(n15285), .C2(n15565), .A(n15276), .B(n15275), .ZN(
        n15277) );
  INV_X1 U18509 ( .A(n15277), .ZN(n15278) );
  OAI21_X1 U18510 ( .B1(n15279), .B2(n19160), .A(n15278), .ZN(P2_U2898) );
  NAND2_X1 U18511 ( .A1(n15596), .A2(n15280), .ZN(n15281) );
  NAND2_X1 U18512 ( .A1(n15573), .A2(n15281), .ZN(n18965) );
  AOI22_X1 U18513 ( .A1(n19110), .A2(BUF1_REG_19__SCAN_IN), .B1(n19109), .B2(
        BUF2_REG_19__SCAN_IN), .ZN(n15284) );
  AOI22_X1 U18514 ( .A1(n19108), .A2(n15282), .B1(n19155), .B2(
        P2_EAX_REG_19__SCAN_IN), .ZN(n15283) );
  OAI211_X1 U18515 ( .C1(n15285), .C2(n18965), .A(n15284), .B(n15283), .ZN(
        n15286) );
  AOI21_X1 U18516 ( .B1(n15287), .B2(n19116), .A(n15286), .ZN(n15288) );
  INV_X1 U18517 ( .A(n15288), .ZN(P2_U2900) );
  NOR2_X1 U18518 ( .A1(n19256), .A2(n15289), .ZN(n15290) );
  AOI211_X1 U18519 ( .C1(n19246), .C2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n15291), .B(n15290), .ZN(n15292) );
  OAI21_X1 U18520 ( .B1(n15293), .B2(n16305), .A(n15292), .ZN(n15294) );
  AOI21_X1 U18521 ( .B1(n15295), .B2(n19248), .A(n15294), .ZN(n15296) );
  OAI21_X1 U18522 ( .B1(n15297), .B2(n16295), .A(n15296), .ZN(P2_U2985) );
  XNOR2_X1 U18523 ( .A(n15298), .B(n15300), .ZN(n15495) );
  INV_X1 U18524 ( .A(n15299), .ZN(n15301) );
  NAND2_X1 U18525 ( .A1(n15301), .A2(n15300), .ZN(n15484) );
  NAND3_X1 U18526 ( .A1(n15484), .A2(n19251), .A3(n12372), .ZN(n15307) );
  NAND2_X1 U18527 ( .A1(n16302), .A2(n15302), .ZN(n15303) );
  OR2_X1 U18528 ( .A1(n15684), .A2(n21193), .ZN(n15488) );
  OAI211_X1 U18529 ( .C1(n16310), .C2(n15304), .A(n15303), .B(n15488), .ZN(
        n15305) );
  AOI21_X1 U18530 ( .B1(n15485), .B2(n19250), .A(n15305), .ZN(n15306) );
  OAI211_X1 U18531 ( .C1(n15495), .C2(n16293), .A(n15307), .B(n15306), .ZN(
        P2_U2987) );
  OAI21_X1 U18532 ( .B1(n15308), .B2(n15318), .A(n15319), .ZN(n15309) );
  XOR2_X1 U18533 ( .A(n15310), .B(n15309), .Z(n15506) );
  AOI21_X1 U18534 ( .B1(n15501), .B2(n15311), .A(n15299), .ZN(n15496) );
  NAND2_X1 U18535 ( .A1(n15496), .A2(n19251), .ZN(n15316) );
  NOR2_X1 U18536 ( .A1(n15684), .A2(n19866), .ZN(n15497) );
  AOI21_X1 U18537 ( .B1(n19246), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n15497), .ZN(n15312) );
  OAI21_X1 U18538 ( .B1(n19256), .B2(n15313), .A(n15312), .ZN(n15314) );
  AOI21_X1 U18539 ( .B1(n16215), .B2(n19250), .A(n15314), .ZN(n15315) );
  OAI211_X1 U18540 ( .C1(n16293), .C2(n15506), .A(n15316), .B(n15315), .ZN(
        P2_U2988) );
  OAI21_X1 U18541 ( .B1(n15317), .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n15311), .ZN(n15519) );
  INV_X1 U18542 ( .A(n15318), .ZN(n15320) );
  NAND2_X1 U18543 ( .A1(n15320), .A2(n15319), .ZN(n15321) );
  XNOR2_X1 U18544 ( .A(n15308), .B(n15321), .ZN(n15517) );
  NOR2_X1 U18545 ( .A1(n15684), .A2(n19864), .ZN(n15508) );
  NOR2_X1 U18546 ( .A1(n16310), .A2(n15322), .ZN(n15323) );
  AOI211_X1 U18547 ( .C1(n15324), .C2(n16302), .A(n15508), .B(n15323), .ZN(
        n15325) );
  OAI21_X1 U18548 ( .B1(n15514), .B2(n16305), .A(n15325), .ZN(n15326) );
  AOI21_X1 U18549 ( .B1(n15517), .B2(n19248), .A(n15326), .ZN(n15327) );
  OAI21_X1 U18550 ( .B1(n15519), .B2(n16295), .A(n15327), .ZN(P2_U2989) );
  XNOR2_X1 U18551 ( .A(n15328), .B(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15329) );
  XNOR2_X1 U18552 ( .A(n15330), .B(n15329), .ZN(n15531) );
  AOI21_X1 U18553 ( .B1(n15333), .B2(n15332), .A(n15317), .ZN(n15520) );
  NAND2_X1 U18554 ( .A1(n15520), .A2(n19251), .ZN(n15339) );
  AOI22_X1 U18555 ( .A1(n19246), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .B1(
        P2_REIP_REG_24__SCAN_IN), .B2(n19038), .ZN(n15334) );
  OAI21_X1 U18556 ( .B1(n19256), .B2(n15335), .A(n15334), .ZN(n15336) );
  AOI21_X1 U18557 ( .B1(n15337), .B2(n19250), .A(n15336), .ZN(n15338) );
  OAI211_X1 U18558 ( .C1(n15531), .C2(n16293), .A(n15339), .B(n15338), .ZN(
        P2_U2990) );
  INV_X1 U18559 ( .A(n15340), .ZN(n15355) );
  INV_X1 U18560 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15551) );
  NOR2_X1 U18561 ( .A1(n15355), .A2(n15551), .ZN(n15354) );
  OAI21_X1 U18562 ( .B1(n15354), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n15332), .ZN(n15544) );
  XOR2_X1 U18563 ( .A(n15342), .B(n15341), .Z(n15541) );
  NAND2_X1 U18564 ( .A1(n19038), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n15536) );
  OAI21_X1 U18565 ( .B1(n16310), .B2(n15343), .A(n15536), .ZN(n15344) );
  AOI21_X1 U18566 ( .B1(n16302), .B2(n15345), .A(n15344), .ZN(n15346) );
  OAI21_X1 U18567 ( .B1(n15347), .B2(n16305), .A(n15346), .ZN(n15348) );
  AOI21_X1 U18568 ( .B1(n15541), .B2(n19248), .A(n15348), .ZN(n15349) );
  OAI21_X1 U18569 ( .B1(n15544), .B2(n16295), .A(n15349), .ZN(P2_U2991) );
  NAND2_X1 U18570 ( .A1(n10236), .A2(n15351), .ZN(n15352) );
  XNOR2_X1 U18571 ( .A(n15353), .B(n15352), .ZN(n15559) );
  AOI21_X1 U18572 ( .B1(n15551), .B2(n15355), .A(n15354), .ZN(n15545) );
  NAND2_X1 U18573 ( .A1(n15545), .A2(n19251), .ZN(n15360) );
  AOI22_X1 U18574 ( .A1(n19246), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B1(
        P2_REIP_REG_22__SCAN_IN), .B2(n19038), .ZN(n15356) );
  OAI21_X1 U18575 ( .B1(n19256), .B2(n15357), .A(n15356), .ZN(n15358) );
  AOI21_X1 U18576 ( .B1(n15856), .B2(n19250), .A(n15358), .ZN(n15359) );
  OAI211_X1 U18577 ( .C1(n15559), .C2(n16293), .A(n15360), .B(n15359), .ZN(
        P2_U2992) );
  INV_X1 U18578 ( .A(n15443), .ZN(n15362) );
  NAND2_X1 U18579 ( .A1(n15428), .A2(n15430), .ZN(n15363) );
  OAI21_X1 U18580 ( .B1(n15429), .B2(n15363), .A(n15431), .ZN(n15848) );
  OAI21_X1 U18581 ( .B1(n15848), .B2(n15849), .A(n15364), .ZN(n15420) );
  NAND2_X1 U18582 ( .A1(n15366), .A2(n15365), .ZN(n15419) );
  INV_X1 U18583 ( .A(n15367), .ZN(n15368) );
  AOI21_X1 U18584 ( .B1(n15382), .B2(n15369), .A(n15385), .ZN(n15374) );
  INV_X1 U18585 ( .A(n15370), .ZN(n15372) );
  NAND2_X1 U18586 ( .A1(n15372), .A2(n15371), .ZN(n15373) );
  XNOR2_X1 U18587 ( .A(n15374), .B(n15373), .ZN(n15570) );
  AOI21_X1 U18588 ( .B1(n15376), .B2(n15387), .A(n15340), .ZN(n15568) );
  NAND2_X1 U18589 ( .A1(n19038), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n15563) );
  OAI21_X1 U18590 ( .B1(n16310), .B2(n11293), .A(n15563), .ZN(n15377) );
  AOI21_X1 U18591 ( .B1(n16302), .B2(n15378), .A(n15377), .ZN(n15379) );
  OAI21_X1 U18592 ( .B1(n15560), .B2(n16305), .A(n15379), .ZN(n15380) );
  AOI21_X1 U18593 ( .B1(n15568), .B2(n19251), .A(n15380), .ZN(n15381) );
  OAI21_X1 U18594 ( .B1(n15570), .B2(n16293), .A(n15381), .ZN(P2_U2993) );
  AOI21_X1 U18595 ( .B1(n15388), .B2(n15386), .A(n15375), .ZN(n15583) );
  NOR2_X1 U18596 ( .A1(n15684), .A2(n19856), .ZN(n15576) );
  AOI21_X1 U18597 ( .B1(n19246), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n15576), .ZN(n15390) );
  NAND2_X1 U18598 ( .A1(n16302), .A2(n18943), .ZN(n15389) );
  OAI211_X1 U18599 ( .C1(n18948), .C2(n16305), .A(n15390), .B(n15389), .ZN(
        n15391) );
  AOI21_X1 U18600 ( .B1(n15583), .B2(n19251), .A(n15391), .ZN(n15392) );
  OAI21_X1 U18601 ( .B1(n15585), .B2(n16293), .A(n15392), .ZN(P2_U2994) );
  NAND2_X1 U18602 ( .A1(n15394), .A2(n15393), .ZN(n15397) );
  INV_X1 U18603 ( .A(n15408), .ZN(n15395) );
  AOI21_X1 U18604 ( .B1(n15410), .B2(n15407), .A(n15395), .ZN(n15396) );
  XOR2_X1 U18605 ( .A(n15397), .B(n15396), .Z(n15595) );
  INV_X1 U18606 ( .A(n15386), .ZN(n15400) );
  AOI21_X1 U18607 ( .B1(n15401), .B2(n9893), .A(n15400), .ZN(n15593) );
  INV_X1 U18608 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n15402) );
  OR2_X1 U18609 ( .A1(n15684), .A2(n19854), .ZN(n15586) );
  OAI21_X1 U18610 ( .B1(n16310), .B2(n15402), .A(n15586), .ZN(n15403) );
  AOI21_X1 U18611 ( .B1(n18959), .B2(n16302), .A(n15403), .ZN(n15404) );
  OAI21_X1 U18612 ( .B1(n18957), .B2(n16305), .A(n15404), .ZN(n15405) );
  AOI21_X1 U18613 ( .B1(n15593), .B2(n19251), .A(n15405), .ZN(n15406) );
  OAI21_X1 U18614 ( .B1(n15595), .B2(n16293), .A(n15406), .ZN(P2_U2995) );
  NAND2_X1 U18615 ( .A1(n15408), .A2(n15407), .ZN(n15409) );
  XNOR2_X1 U18616 ( .A(n15410), .B(n15409), .ZN(n15609) );
  NOR2_X1 U18617 ( .A1(n15684), .A2(n15411), .ZN(n15601) );
  AOI21_X1 U18618 ( .B1(n19246), .B2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n15601), .ZN(n15412) );
  OAI21_X1 U18619 ( .B1(n18967), .B2(n19256), .A(n15412), .ZN(n15417) );
  OAI21_X1 U18620 ( .B1(n16241), .B2(n15622), .A(n15414), .ZN(n15415) );
  NAND2_X1 U18621 ( .A1(n9893), .A2(n15415), .ZN(n15604) );
  NOR2_X1 U18622 ( .A1(n15604), .A2(n16295), .ZN(n15416) );
  AOI211_X1 U18623 ( .C1(n19250), .C2(n18973), .A(n15417), .B(n15416), .ZN(
        n15418) );
  OAI21_X1 U18624 ( .B1(n16293), .B2(n15609), .A(n15418), .ZN(P2_U2996) );
  XNOR2_X1 U18625 ( .A(n16241), .B(n15622), .ZN(n15427) );
  XNOR2_X1 U18626 ( .A(n15420), .B(n15419), .ZN(n15619) );
  NAND2_X1 U18627 ( .A1(n15619), .A2(n19248), .ZN(n15426) );
  INV_X1 U18628 ( .A(n15421), .ZN(n18982) );
  NOR2_X1 U18629 ( .A1(n21095), .A2(n12458), .ZN(n15424) );
  INV_X1 U18630 ( .A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n15422) );
  OAI22_X1 U18631 ( .A1(n16310), .A2(n15422), .B1(n19256), .B2(n18984), .ZN(
        n15423) );
  AOI211_X1 U18632 ( .C1(n18982), .C2(n19250), .A(n15424), .B(n15423), .ZN(
        n15425) );
  OAI211_X1 U18633 ( .C1(n16295), .C2(n15427), .A(n15426), .B(n15425), .ZN(
        P2_U2997) );
  INV_X1 U18634 ( .A(n15428), .ZN(n15627) );
  NOR2_X1 U18635 ( .A1(n15429), .A2(n15627), .ZN(n15433) );
  NAND2_X1 U18636 ( .A1(n15431), .A2(n15430), .ZN(n15432) );
  XNOR2_X1 U18637 ( .A(n15433), .B(n15432), .ZN(n16322) );
  NAND2_X1 U18638 ( .A1(n15615), .A2(n12221), .ZN(n15435) );
  NAND2_X1 U18639 ( .A1(n16240), .A2(n15435), .ZN(n16317) );
  INV_X1 U18640 ( .A(n16317), .ZN(n15440) );
  INV_X1 U18641 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n15436) );
  OAI22_X1 U18642 ( .A1(n16310), .A2(n15436), .B1(n19256), .B2(n19009), .ZN(
        n15439) );
  INV_X1 U18643 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n15437) );
  OAI22_X1 U18644 ( .A1(n19005), .A2(n16305), .B1(n15437), .B2(n12458), .ZN(
        n15438) );
  AOI211_X1 U18645 ( .C1(n15440), .C2(n19251), .A(n15439), .B(n15438), .ZN(
        n15441) );
  OAI21_X1 U18646 ( .B1(n16322), .B2(n16293), .A(n15441), .ZN(P2_U2999) );
  NAND2_X1 U18647 ( .A1(n15398), .A2(n15636), .ZN(n15625) );
  OAI21_X1 U18648 ( .B1(n15675), .B2(n15659), .A(n21086), .ZN(n15442) );
  NAND2_X1 U18649 ( .A1(n15625), .A2(n15442), .ZN(n15658) );
  NAND2_X1 U18650 ( .A1(n15444), .A2(n15443), .ZN(n15446) );
  XOR2_X1 U18651 ( .A(n15446), .B(n15445), .Z(n15656) );
  INV_X1 U18652 ( .A(n19025), .ZN(n15447) );
  OAI22_X1 U18653 ( .A1(n16310), .A2(n15448), .B1(n19256), .B2(n15447), .ZN(
        n15451) );
  OAI22_X1 U18654 ( .A1(n19029), .A2(n16305), .B1(n15449), .B2(n12458), .ZN(
        n15450) );
  AOI211_X1 U18655 ( .C1(n15656), .C2(n19248), .A(n15451), .B(n15450), .ZN(
        n15452) );
  OAI21_X1 U18656 ( .B1(n15658), .B2(n16295), .A(n15452), .ZN(P2_U3001) );
  NAND2_X1 U18657 ( .A1(n15454), .A2(n15453), .ZN(n15455) );
  XNOR2_X1 U18658 ( .A(n15455), .B(n15730), .ZN(n15734) );
  NAND2_X1 U18659 ( .A1(n15457), .A2(n15456), .ZN(n16284) );
  NAND2_X1 U18660 ( .A1(n16281), .A2(n16283), .ZN(n15458) );
  XNOR2_X1 U18661 ( .A(n16284), .B(n15458), .ZN(n15731) );
  OAI22_X1 U18662 ( .A1(n16310), .A2(n15459), .B1(n11530), .B2(n15684), .ZN(
        n15460) );
  AOI21_X1 U18663 ( .B1(n16302), .B2(n19047), .A(n15460), .ZN(n15461) );
  OAI21_X1 U18664 ( .B1(n19052), .B2(n16305), .A(n15461), .ZN(n15462) );
  AOI21_X1 U18665 ( .B1(n15731), .B2(n19248), .A(n15462), .ZN(n15463) );
  OAI21_X1 U18666 ( .B1(n15734), .B2(n16295), .A(n15463), .ZN(P2_U3007) );
  XNOR2_X1 U18667 ( .A(n19094), .B(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n16337) );
  AOI22_X1 U18668 ( .A1(n19250), .A2(n19098), .B1(n19248), .B2(n16337), .ZN(
        n15470) );
  OR2_X1 U18669 ( .A1(n15684), .A2(n18929), .ZN(n16347) );
  OAI21_X1 U18670 ( .B1(n19246), .B2(n15464), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n15469) );
  NAND2_X1 U18671 ( .A1(n15465), .A2(n11481), .ZN(n15467) );
  AND2_X1 U18672 ( .A1(n15467), .A2(n15466), .ZN(n16341) );
  NAND2_X1 U18673 ( .A1(n19251), .A2(n16341), .ZN(n15468) );
  NAND4_X1 U18674 ( .A1(n15470), .A2(n16347), .A3(n15469), .A4(n15468), .ZN(
        P2_U3014) );
  NAND2_X1 U18675 ( .A1(n15471), .A2(n16342), .ZN(n15482) );
  NOR2_X1 U18676 ( .A1(n15472), .A2(n16326), .ZN(n15479) );
  NAND3_X1 U18677 ( .A1(n15474), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A3(
        n15473), .ZN(n15475) );
  OAI211_X1 U18678 ( .C1(n16313), .C2(n15477), .A(n15476), .B(n15475), .ZN(
        n15478) );
  AOI211_X1 U18679 ( .C1(n15480), .C2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n15479), .B(n15478), .ZN(n15481) );
  OAI211_X1 U18680 ( .C1(n15483), .C2(n16321), .A(n15482), .B(n15481), .ZN(
        P2_U3018) );
  NAND3_X1 U18681 ( .A1(n15484), .A2(n16342), .A3(n12372), .ZN(n15494) );
  NAND2_X1 U18682 ( .A1(n15485), .A2(n16340), .ZN(n15490) );
  NAND2_X1 U18683 ( .A1(n16344), .A2(n15486), .ZN(n15487) );
  NAND4_X1 U18684 ( .A1(n15490), .A2(n15489), .A3(n15488), .A4(n15487), .ZN(
        n15491) );
  AOI21_X1 U18685 ( .B1(n15492), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n15491), .ZN(n15493) );
  OAI211_X1 U18686 ( .C1(n15495), .C2(n16321), .A(n15494), .B(n15493), .ZN(
        P2_U3019) );
  NAND2_X1 U18687 ( .A1(n15496), .A2(n16342), .ZN(n15505) );
  INV_X1 U18688 ( .A(n15497), .ZN(n15500) );
  OAI211_X1 U18689 ( .C1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(n15510), .B(n15498), .ZN(
        n15499) );
  OAI211_X1 U18690 ( .C1(n16313), .C2(n16213), .A(n15500), .B(n15499), .ZN(
        n15503) );
  NOR2_X1 U18691 ( .A1(n15507), .A2(n15501), .ZN(n15502) );
  AOI211_X1 U18692 ( .C1(n16215), .C2(n16340), .A(n15503), .B(n15502), .ZN(
        n15504) );
  OAI211_X1 U18693 ( .C1(n15506), .C2(n16321), .A(n15505), .B(n15504), .ZN(
        P2_U3020) );
  NOR2_X1 U18694 ( .A1(n15507), .A2(n15509), .ZN(n15516) );
  AOI21_X1 U18695 ( .B1(n15510), .B2(n15509), .A(n15508), .ZN(n15513) );
  NAND2_X1 U18696 ( .A1(n16344), .A2(n15511), .ZN(n15512) );
  OAI211_X1 U18697 ( .C1(n15514), .C2(n16326), .A(n15513), .B(n15512), .ZN(
        n15515) );
  AOI211_X1 U18698 ( .C1(n15517), .C2(n16338), .A(n15516), .B(n15515), .ZN(
        n15518) );
  OAI21_X1 U18699 ( .B1(n15519), .B2(n16327), .A(n15518), .ZN(P2_U3021) );
  NAND2_X1 U18700 ( .A1(n15520), .A2(n16342), .ZN(n15530) );
  INV_X1 U18701 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n19862) );
  NOR2_X1 U18702 ( .A1(n19862), .A2(n15684), .ZN(n15523) );
  INV_X1 U18703 ( .A(n15521), .ZN(n15534) );
  NOR3_X1 U18704 ( .A1(n15533), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(
        n15534), .ZN(n15522) );
  AOI211_X1 U18705 ( .C1(n16344), .C2(n15524), .A(n15523), .B(n15522), .ZN(
        n15525) );
  OAI21_X1 U18706 ( .B1(n15526), .B2(n16326), .A(n15525), .ZN(n15527) );
  AOI21_X1 U18707 ( .B1(n15528), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n15527), .ZN(n15529) );
  OAI211_X1 U18708 ( .C1(n15531), .C2(n16321), .A(n15530), .B(n15529), .ZN(
        P2_U3022) );
  NOR2_X1 U18709 ( .A1(n15546), .A2(n15532), .ZN(n15539) );
  INV_X1 U18710 ( .A(n15533), .ZN(n15552) );
  OAI211_X1 U18711 ( .C1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(n15552), .B(n15534), .ZN(
        n15535) );
  OAI211_X1 U18712 ( .C1(n16313), .C2(n15537), .A(n15536), .B(n15535), .ZN(
        n15538) );
  AOI211_X1 U18713 ( .C1(n15540), .C2(n16340), .A(n15539), .B(n15538), .ZN(
        n15543) );
  NAND2_X1 U18714 ( .A1(n15541), .A2(n16338), .ZN(n15542) );
  OAI211_X1 U18715 ( .C1(n15544), .C2(n16327), .A(n15543), .B(n15542), .ZN(
        P2_U3023) );
  NAND2_X1 U18716 ( .A1(n15545), .A2(n16342), .ZN(n15558) );
  NOR2_X1 U18717 ( .A1(n15546), .A2(n15551), .ZN(n15556) );
  NOR2_X1 U18718 ( .A1(n15548), .A2(n15547), .ZN(n15549) );
  OR2_X1 U18719 ( .A1(n15550), .A2(n15549), .ZN(n15855) );
  NAND2_X1 U18720 ( .A1(P2_REIP_REG_22__SCAN_IN), .A2(n19038), .ZN(n15554) );
  NAND2_X1 U18721 ( .A1(n15552), .A2(n15551), .ZN(n15553) );
  OAI211_X1 U18722 ( .C1(n16313), .C2(n15855), .A(n15554), .B(n15553), .ZN(
        n15555) );
  AOI211_X1 U18723 ( .C1(n15856), .C2(n16340), .A(n15556), .B(n15555), .ZN(
        n15557) );
  OAI211_X1 U18724 ( .C1(n15559), .C2(n16321), .A(n15558), .B(n15557), .ZN(
        P2_U3024) );
  NOR2_X1 U18725 ( .A1(n15560), .A2(n16326), .ZN(n15567) );
  NOR2_X1 U18726 ( .A1(n15587), .A2(n15571), .ZN(n15562) );
  OAI21_X1 U18727 ( .B1(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .B2(n15562), .A(
        n15561), .ZN(n15564) );
  OAI211_X1 U18728 ( .C1(n16313), .C2(n15565), .A(n15564), .B(n15563), .ZN(
        n15566) );
  AOI211_X1 U18729 ( .C1(n15568), .C2(n16342), .A(n15567), .B(n15566), .ZN(
        n15569) );
  OAI21_X1 U18730 ( .B1(n15570), .B2(n16321), .A(n15569), .ZN(P2_U3025) );
  OAI21_X1 U18731 ( .B1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(n15571), .ZN(n15579) );
  AND2_X1 U18732 ( .A1(n15573), .A2(n15572), .ZN(n15574) );
  NOR2_X1 U18733 ( .A1(n15575), .A2(n15574), .ZN(n18951) );
  NAND2_X1 U18734 ( .A1(n16344), .A2(n18951), .ZN(n15578) );
  INV_X1 U18735 ( .A(n15576), .ZN(n15577) );
  OAI211_X1 U18736 ( .C1(n15587), .C2(n15579), .A(n15578), .B(n15577), .ZN(
        n15580) );
  AOI21_X1 U18737 ( .B1(n15607), .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n15580), .ZN(n15581) );
  OAI21_X1 U18738 ( .B1(n18948), .B2(n16326), .A(n15581), .ZN(n15582) );
  AOI21_X1 U18739 ( .B1(n15583), .B2(n16342), .A(n15582), .ZN(n15584) );
  OAI21_X1 U18740 ( .B1(n15585), .B2(n16321), .A(n15584), .ZN(P2_U3026) );
  INV_X1 U18741 ( .A(n18965), .ZN(n15589) );
  OAI21_X1 U18742 ( .B1(n15587), .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n15586), .ZN(n15588) );
  AOI21_X1 U18743 ( .B1(n16344), .B2(n15589), .A(n15588), .ZN(n15591) );
  NAND2_X1 U18744 ( .A1(n15607), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15590) );
  OAI211_X1 U18745 ( .C1(n18957), .C2(n16326), .A(n15591), .B(n15590), .ZN(
        n15592) );
  AOI21_X1 U18746 ( .B1(n15593), .B2(n16342), .A(n15592), .ZN(n15594) );
  OAI21_X1 U18747 ( .B1(n15595), .B2(n16321), .A(n15594), .ZN(P2_U3027) );
  INV_X1 U18748 ( .A(n15596), .ZN(n15597) );
  AOI21_X1 U18749 ( .B1(n15598), .B2(n14313), .A(n15597), .ZN(n18972) );
  NOR2_X1 U18750 ( .A1(n15599), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15600) );
  AOI211_X1 U18751 ( .C1(n16344), .C2(n18972), .A(n15601), .B(n15600), .ZN(
        n15602) );
  OAI21_X1 U18752 ( .B1(n15603), .B2(n16326), .A(n15602), .ZN(n15606) );
  NOR2_X1 U18753 ( .A1(n15604), .A2(n16327), .ZN(n15605) );
  AOI211_X1 U18754 ( .C1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .C2(n15607), .A(
        n15606), .B(n15605), .ZN(n15608) );
  OAI21_X1 U18755 ( .B1(n16321), .B2(n15609), .A(n15608), .ZN(P2_U3028) );
  OAI21_X1 U18756 ( .B1(n16342), .B2(n15610), .A(n16241), .ZN(n15611) );
  OAI211_X1 U18757 ( .C1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n15612), .A(
        n15611), .B(n16311), .ZN(n15850) );
  AOI21_X1 U18758 ( .B1(n15614), .B2(n15613), .A(n15850), .ZN(n15623) );
  OAI22_X1 U18759 ( .A1(n16313), .A2(n18980), .B1(n21095), .B2(n12458), .ZN(
        n15618) );
  AOI21_X1 U18760 ( .B1(n15624), .B2(n16342), .A(n16316), .ZN(n15851) );
  NOR3_X1 U18761 ( .A1(n15851), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A3(
        n15616), .ZN(n15617) );
  AOI211_X1 U18762 ( .C1(n18982), .C2(n16340), .A(n15618), .B(n15617), .ZN(
        n15621) );
  NAND2_X1 U18763 ( .A1(n15619), .A2(n16338), .ZN(n15620) );
  OAI211_X1 U18764 ( .C1(n15623), .C2(n15622), .A(n15621), .B(n15620), .ZN(
        P2_U3029) );
  INV_X1 U18765 ( .A(n16247), .ZN(n15646) );
  NOR2_X1 U18766 ( .A1(n15627), .A2(n15626), .ZN(n15628) );
  XNOR2_X1 U18767 ( .A(n15629), .B(n15628), .ZN(n16248) );
  INV_X1 U18768 ( .A(n19020), .ZN(n15643) );
  INV_X1 U18769 ( .A(n15648), .ZN(n15630) );
  OR2_X1 U18770 ( .A1(n15631), .A2(n15630), .ZN(n15634) );
  INV_X1 U18771 ( .A(n15632), .ZN(n15633) );
  AND2_X1 U18772 ( .A1(n15634), .A2(n15633), .ZN(n19119) );
  NOR2_X1 U18773 ( .A1(n15684), .A2(n11919), .ZN(n15641) );
  NOR2_X1 U18774 ( .A1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n15666), .ZN(
        n15650) );
  OAI21_X1 U18775 ( .B1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n15666), .A(
        n15665), .ZN(n15651) );
  NOR2_X1 U18776 ( .A1(n15650), .A2(n15651), .ZN(n15639) );
  INV_X1 U18777 ( .A(n15666), .ZN(n15635) );
  NAND3_X1 U18778 ( .A1(n15636), .A2(n15638), .A3(n15635), .ZN(n15637) );
  OAI21_X1 U18779 ( .B1(n15639), .B2(n15638), .A(n15637), .ZN(n15640) );
  AOI211_X1 U18780 ( .C1(n16344), .C2(n19119), .A(n15641), .B(n15640), .ZN(
        n15642) );
  OAI21_X1 U18781 ( .B1(n15643), .B2(n16326), .A(n15642), .ZN(n15644) );
  AOI21_X1 U18782 ( .B1(n16248), .B2(n16338), .A(n15644), .ZN(n15645) );
  OAI21_X1 U18783 ( .B1(n15646), .B2(n16327), .A(n15645), .ZN(P2_U3032) );
  OR2_X1 U18784 ( .A1(n15647), .A2(n14266), .ZN(n15649) );
  NAND2_X1 U18785 ( .A1(n15649), .A2(n15648), .ZN(n19123) );
  NOR2_X1 U18786 ( .A1(n16313), .A2(n19123), .ZN(n15655) );
  AOI22_X1 U18787 ( .A1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n15651), .B1(
        P2_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n15650), .ZN(n15653) );
  OR2_X1 U18788 ( .A1(n15449), .A2(n15684), .ZN(n15652) );
  OAI211_X1 U18789 ( .C1(n19029), .C2(n16326), .A(n15653), .B(n15652), .ZN(
        n15654) );
  AOI211_X1 U18790 ( .C1(n15656), .C2(n16338), .A(n15655), .B(n15654), .ZN(
        n15657) );
  OAI21_X1 U18791 ( .B1(n15658), .B2(n16327), .A(n15657), .ZN(P2_U3033) );
  XNOR2_X1 U18792 ( .A(n15675), .B(n15659), .ZN(n16251) );
  NAND2_X1 U18793 ( .A1(n15661), .A2(n15660), .ZN(n15663) );
  XOR2_X1 U18794 ( .A(n15663), .B(n15662), .Z(n16254) );
  NAND2_X1 U18795 ( .A1(P2_REIP_REG_12__SCAN_IN), .A2(n19038), .ZN(n15664) );
  OAI221_X1 U18796 ( .B1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n15666), 
        .C1(n15659), .C2(n15665), .A(n15664), .ZN(n15669) );
  INV_X1 U18797 ( .A(n15667), .ZN(n19126) );
  OAI22_X1 U18798 ( .A1(n16252), .A2(n16326), .B1(n16313), .B2(n19126), .ZN(
        n15668) );
  AOI211_X1 U18799 ( .C1(n16254), .C2(n16338), .A(n15669), .B(n15668), .ZN(
        n15670) );
  OAI21_X1 U18800 ( .B1(n16251), .B2(n16327), .A(n15670), .ZN(P2_U3034) );
  XNOR2_X1 U18801 ( .A(n15671), .B(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n15672) );
  XNOR2_X1 U18802 ( .A(n15673), .B(n15672), .ZN(n16260) );
  INV_X1 U18803 ( .A(n15674), .ZN(n15707) );
  NOR2_X1 U18804 ( .A1(n15707), .A2(n12180), .ZN(n15683) );
  OAI21_X1 U18805 ( .B1(n15683), .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n15675), .ZN(n16261) );
  OR2_X1 U18806 ( .A1(n16261), .A2(n16327), .ZN(n15682) );
  XNOR2_X1 U18807 ( .A(n15676), .B(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n15680) );
  NAND2_X1 U18808 ( .A1(n15686), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n15678) );
  AOI22_X1 U18809 ( .A1(n16263), .A2(n16340), .B1(P2_REIP_REG_11__SCAN_IN), 
        .B2(n19038), .ZN(n15677) );
  OAI211_X1 U18810 ( .C1(n16313), .C2(n19128), .A(n15678), .B(n15677), .ZN(
        n15679) );
  AOI21_X1 U18811 ( .B1(n15687), .B2(n15680), .A(n15679), .ZN(n15681) );
  OAI211_X1 U18812 ( .C1(n16260), .C2(n16321), .A(n15682), .B(n15681), .ZN(
        P2_U3035) );
  AOI21_X1 U18813 ( .B1(n12180), .B2(n15707), .A(n15683), .ZN(n16267) );
  NAND2_X1 U18814 ( .A1(n16267), .A2(n16342), .ZN(n15706) );
  NOR2_X1 U18815 ( .A1(n11864), .A2(n15684), .ZN(n15685) );
  AOI221_X1 U18816 ( .B1(n15687), .B2(n12180), .C1(n15686), .C2(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A(n15685), .ZN(n15705) );
  XNOR2_X1 U18817 ( .A(n15689), .B(n15688), .ZN(n19132) );
  INV_X1 U18818 ( .A(n19042), .ZN(n15690) );
  OAI22_X1 U18819 ( .A1(n19132), .A2(n16313), .B1(n16326), .B2(n15690), .ZN(
        n15691) );
  INV_X1 U18820 ( .A(n15691), .ZN(n15704) );
  INV_X1 U18821 ( .A(n15692), .ZN(n15693) );
  OR2_X1 U18822 ( .A1(n16284), .A2(n15693), .ZN(n15695) );
  NAND2_X1 U18823 ( .A1(n15695), .A2(n15694), .ZN(n15720) );
  INV_X1 U18824 ( .A(n15717), .ZN(n15697) );
  INV_X1 U18825 ( .A(n15696), .ZN(n15718) );
  OAI21_X1 U18826 ( .B1(n15720), .B2(n15697), .A(n15718), .ZN(n15702) );
  INV_X1 U18827 ( .A(n15698), .ZN(n15700) );
  NAND2_X1 U18828 ( .A1(n15700), .A2(n15699), .ZN(n15701) );
  XNOR2_X1 U18829 ( .A(n15702), .B(n15701), .ZN(n16268) );
  NAND2_X1 U18830 ( .A1(n16268), .A2(n16338), .ZN(n15703) );
  NAND4_X1 U18831 ( .A1(n15706), .A2(n15705), .A3(n15704), .A4(n15703), .ZN(
        P2_U3036) );
  OAI21_X1 U18832 ( .B1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n15708), .A(
        n15707), .ZN(n16273) );
  NOR2_X1 U18833 ( .A1(n15709), .A2(n16326), .ZN(n15715) );
  NAND2_X1 U18834 ( .A1(P2_REIP_REG_9__SCAN_IN), .A2(n19038), .ZN(n15710) );
  OAI221_X1 U18835 ( .B1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n15713), .C1(
        n15712), .C2(n15711), .A(n15710), .ZN(n15714) );
  AOI211_X1 U18836 ( .C1(n15716), .C2(n16344), .A(n15715), .B(n15714), .ZN(
        n15722) );
  NAND2_X1 U18837 ( .A1(n15718), .A2(n15717), .ZN(n15719) );
  XNOR2_X1 U18838 ( .A(n15720), .B(n15719), .ZN(n16272) );
  OR2_X1 U18839 ( .A1(n16272), .A2(n16321), .ZN(n15721) );
  OAI211_X1 U18840 ( .C1(n16273), .C2(n16327), .A(n15722), .B(n15721), .ZN(
        P2_U3037) );
  OAI21_X1 U18841 ( .B1(n16351), .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n15723), .ZN(n16323) );
  AOI22_X1 U18842 ( .A1(n16323), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .B1(
        n19038), .B2(P2_REIP_REG_7__SCAN_IN), .ZN(n15724) );
  OAI21_X1 U18843 ( .B1(n19052), .B2(n16326), .A(n15724), .ZN(n15729) );
  OR2_X1 U18844 ( .A1(n15726), .A2(n15725), .ZN(n15727) );
  NAND2_X1 U18845 ( .A1(n15727), .A2(n14184), .ZN(n19138) );
  NOR2_X1 U18846 ( .A1(n19138), .A2(n16313), .ZN(n15728) );
  AOI211_X1 U18847 ( .C1(n16332), .C2(n15730), .A(n15729), .B(n15728), .ZN(
        n15733) );
  NAND2_X1 U18848 ( .A1(n15731), .A2(n16338), .ZN(n15732) );
  OAI211_X1 U18849 ( .C1(n15734), .C2(n16327), .A(n15733), .B(n15732), .ZN(
        P2_U3039) );
  INV_X1 U18850 ( .A(n16397), .ZN(n15782) );
  INV_X1 U18851 ( .A(n12421), .ZN(n15736) );
  NAND2_X1 U18852 ( .A1(n15736), .A2(n15735), .ZN(n15742) );
  MUX2_X1 U18853 ( .A(n15774), .B(n15742), .S(n15737), .Z(n15738) );
  AOI21_X1 U18854 ( .B1(n19098), .B2(n15781), .A(n15738), .ZN(n16352) );
  INV_X1 U18855 ( .A(n15739), .ZN(n19099) );
  AOI22_X1 U18856 ( .A1(n10053), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        n19099), .B2(n19079), .ZN(n15747) );
  INV_X1 U18857 ( .A(n15747), .ZN(n15740) );
  OAI222_X1 U18858 ( .A1(n15782), .A2(n12678), .B1(n19890), .B2(n16352), .C1(
        n19802), .C2(n15740), .ZN(n15741) );
  MUX2_X1 U18859 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B(n15741), .S(
        n15783), .Z(P2_U3601) );
  INV_X1 U18860 ( .A(n15774), .ZN(n15745) );
  OAI21_X1 U18861 ( .B1(n11653), .B2(n15743), .A(n15742), .ZN(n15744) );
  OAI21_X1 U18862 ( .B1(n15745), .B2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n15744), .ZN(n15746) );
  AOI21_X1 U18863 ( .B1(n12673), .B2(n15781), .A(n15746), .ZN(n16353) );
  NOR2_X1 U18864 ( .A1(n15747), .A2(n19802), .ZN(n15766) );
  INV_X1 U18865 ( .A(n15766), .ZN(n15750) );
  OAI21_X1 U18866 ( .B1(n19079), .B2(n15749), .A(n15748), .ZN(n15765) );
  OAI222_X1 U18867 ( .A1(n19890), .A2(n16353), .B1(n15782), .B2(n19910), .C1(
        n15750), .C2(n15765), .ZN(n15751) );
  MUX2_X1 U18868 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n15751), .S(
        n15783), .Z(P2_U3600) );
  INV_X1 U18869 ( .A(n15781), .ZN(n15753) );
  OR2_X1 U18870 ( .A1(n13628), .A2(n15753), .ZN(n15764) );
  INV_X1 U18871 ( .A(n11654), .ZN(n15755) );
  NAND2_X1 U18872 ( .A1(n15755), .A2(n15754), .ZN(n15770) );
  INV_X1 U18873 ( .A(n15770), .ZN(n15772) );
  NAND2_X1 U18874 ( .A1(n11472), .A2(n15756), .ZN(n15757) );
  NAND2_X1 U18875 ( .A1(n15757), .A2(n12801), .ZN(n15775) );
  OR2_X1 U18876 ( .A1(n16364), .A2(n16366), .ZN(n15771) );
  OAI21_X1 U18877 ( .B1(n11652), .B2(n15772), .A(n15771), .ZN(n15761) );
  NOR2_X1 U18878 ( .A1(n15758), .A2(n12291), .ZN(n15759) );
  NAND2_X1 U18879 ( .A1(n15774), .A2(n15759), .ZN(n15760) );
  OAI211_X1 U18880 ( .C1(n15772), .C2(n15775), .A(n15761), .B(n15760), .ZN(
        n15762) );
  INV_X1 U18881 ( .A(n15762), .ZN(n15763) );
  NAND2_X1 U18882 ( .A1(n15764), .A2(n15763), .ZN(n16358) );
  AOI22_X1 U18883 ( .A1(n16358), .A2(n15767), .B1(n15766), .B2(n15765), .ZN(
        n15768) );
  OAI21_X1 U18884 ( .B1(n19901), .B2(n15782), .A(n15768), .ZN(n15769) );
  MUX2_X1 U18885 ( .A(n15752), .B(n15769), .S(n15783), .Z(P2_U3599) );
  AOI22_X1 U18886 ( .A1(n15771), .A2(n15770), .B1(n12291), .B2(n15774), .ZN(
        n15778) );
  INV_X1 U18887 ( .A(n12291), .ZN(n15773) );
  AOI21_X1 U18888 ( .B1(n15774), .B2(n15773), .A(n15772), .ZN(n15776) );
  AND2_X1 U18889 ( .A1(n15776), .A2(n15775), .ZN(n15777) );
  MUX2_X1 U18890 ( .A(n15778), .B(n15777), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n15779) );
  NAND2_X1 U18891 ( .A1(n15779), .A2(n10264), .ZN(n15780) );
  AOI21_X1 U18892 ( .B1(n14053), .B2(n15781), .A(n15780), .ZN(n16357) );
  OAI22_X1 U18893 ( .A1(n19539), .A2(n15782), .B1(n16357), .B2(n19890), .ZN(
        n15784) );
  MUX2_X1 U18894 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n15784), .S(
        n15783), .Z(P2_U3596) );
  AOI22_X1 U18895 ( .A1(n17199), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17211), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n15789) );
  AOI22_X1 U18896 ( .A1(n17147), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n9837), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n15788) );
  AOI22_X1 U18897 ( .A1(n9849), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n15785), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n15787) );
  AOI22_X1 U18898 ( .A1(n17220), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17194), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n15786) );
  NAND4_X1 U18899 ( .A1(n15789), .A2(n15788), .A3(n15787), .A4(n15786), .ZN(
        n15795) );
  AOI22_X1 U18900 ( .A1(n17112), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n9838), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n15793) );
  AOI22_X1 U18901 ( .A1(n9832), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n17153), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n15792) );
  AOI22_X1 U18902 ( .A1(n9851), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(n9839), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n15791) );
  AOI22_X1 U18903 ( .A1(n13013), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n17213), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n15790) );
  NAND4_X1 U18904 ( .A1(n15793), .A2(n15792), .A3(n15791), .A4(n15790), .ZN(
        n15794) );
  NOR2_X1 U18905 ( .A1(n15795), .A2(n15794), .ZN(n17368) );
  NOR2_X1 U18906 ( .A1(n17267), .A2(n15796), .ZN(n17160) );
  INV_X1 U18907 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n16792) );
  OAI222_X1 U18908 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(n18277), .B1(
        P3_EBX_REG_13__SCAN_IN), .B2(n15796), .C1(n17160), .C2(n16792), .ZN(
        n15797) );
  OAI21_X1 U18909 ( .B1(n17368), .B2(n17260), .A(n15797), .ZN(P3_U2690) );
  NAND2_X1 U18910 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18459) );
  AOI221_X1 U18911 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n18459), .C1(n15799), 
        .C2(n18459), .A(n15798), .ZN(n18241) );
  NOR2_X1 U18912 ( .A1(n15800), .A2(n18718), .ZN(n15801) );
  OAI21_X1 U18913 ( .B1(n15801), .B2(n18593), .A(n18242), .ZN(n18239) );
  AOI22_X1 U18914 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18241), .B1(
        n18239), .B2(n18723), .ZN(P3_U2865) );
  NOR2_X1 U18915 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18864), .ZN(n18247) );
  NAND2_X1 U18916 ( .A1(READY22_REG_SCAN_IN), .A2(READY2), .ZN(n18880) );
  INV_X1 U18917 ( .A(n18880), .ZN(n18889) );
  NOR2_X1 U18918 ( .A1(n18889), .A2(n15825), .ZN(n15810) );
  INV_X1 U18919 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n18767) );
  INV_X2 U18920 ( .A(n18899), .ZN(n18898) );
  NAND2_X2 U18921 ( .A1(n18898), .A2(P3_STATE_REG_2__SCAN_IN), .ZN(n18826) );
  OAI211_X1 U18922 ( .C1(P3_STATE_REG_1__SCAN_IN), .C2(P3_STATE_REG_2__SCAN_IN), .A(n18767), .B(n18826), .ZN(n18885) );
  NOR2_X1 U18923 ( .A1(n15802), .A2(n18885), .ZN(n17427) );
  OAI21_X1 U18924 ( .B1(n15807), .B2(n15806), .A(n15805), .ZN(n15809) );
  NAND2_X1 U18925 ( .A1(n15809), .A2(n15808), .ZN(n15827) );
  AOI211_X1 U18926 ( .C1(n15810), .C2(n17427), .A(n15921), .B(n15827), .ZN(
        n15811) );
  OAI21_X1 U18927 ( .B1(n15813), .B2(n15812), .A(n15811), .ZN(n18711) );
  INV_X1 U18928 ( .A(n18711), .ZN(n18721) );
  INV_X1 U18929 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n21087) );
  OAI22_X1 U18930 ( .A1(n18721), .A2(n18743), .B1(n21087), .B2(n18836), .ZN(
        n15814) );
  INV_X1 U18931 ( .A(n18869), .ZN(n18860) );
  INV_X1 U18932 ( .A(n18700), .ZN(n18704) );
  AOI21_X1 U18933 ( .B1(n18704), .B2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n15817) );
  NOR3_X1 U18934 ( .A1(n15817), .A2(n15816), .A3(n15815), .ZN(n18733) );
  NAND3_X1 U18935 ( .A1(n18860), .A2(n18902), .A3(n18733), .ZN(n15818) );
  OAI21_X1 U18936 ( .B1(n18860), .B2(n18691), .A(n15818), .ZN(P3_U3284) );
  AOI22_X1 U18937 ( .A1(n17818), .A2(n17553), .B1(n15820), .B2(n15819), .ZN(
        n15821) );
  XNOR2_X1 U18938 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B(n15821), .ZN(
        n16434) );
  INV_X1 U18939 ( .A(n16454), .ZN(n18687) );
  INV_X1 U18940 ( .A(n15822), .ZN(n15829) );
  OAI21_X1 U18941 ( .B1(n18254), .B2(n16589), .A(n18885), .ZN(n15823) );
  OAI21_X1 U18942 ( .B1(n15824), .B2(n15823), .A(n18880), .ZN(n16558) );
  NOR3_X1 U18943 ( .A1(n15826), .A2(n15825), .A3(n16558), .ZN(n15828) );
  AOI211_X1 U18944 ( .C1(n15829), .C2(n18686), .A(n15828), .B(n15827), .ZN(
        n15833) );
  OAI21_X1 U18945 ( .B1(n15831), .B2(n15830), .A(n18682), .ZN(n15832) );
  NOR3_X4 U18946 ( .A1(n17393), .A2(n18687), .A3(n18214), .ZN(n18147) );
  INV_X1 U18947 ( .A(n18147), .ZN(n18123) );
  NAND2_X1 U18948 ( .A1(n16454), .A2(n17393), .ZN(n18083) );
  NOR2_X1 U18949 ( .A1(n18214), .A2(n18083), .ZN(n18021) );
  INV_X1 U18950 ( .A(n18021), .ZN(n18151) );
  NAND2_X1 U18951 ( .A1(n18681), .A2(n18227), .ZN(n18224) );
  OAI22_X1 U18952 ( .A1(n16425), .A2(n18151), .B1(n16427), .B2(n18224), .ZN(
        n15911) );
  INV_X2 U18953 ( .A(n18218), .ZN(n18231) );
  INV_X1 U18954 ( .A(n18118), .ZN(n18109) );
  INV_X1 U18955 ( .A(n18710), .ZN(n18203) );
  NAND2_X1 U18956 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18179) );
  NAND3_X1 U18957 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n18049) );
  NOR2_X1 U18958 ( .A1(n18179), .A2(n18049), .ZN(n18137) );
  INV_X1 U18959 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n20916) );
  NOR3_X1 U18960 ( .A1(n20916), .A2(n18163), .A3(n18144), .ZN(n18050) );
  NAND2_X1 U18961 ( .A1(n18137), .A2(n18050), .ZN(n18066) );
  NOR2_X1 U18962 ( .A1(n18024), .A2(n18066), .ZN(n17919) );
  NAND2_X1 U18963 ( .A1(n17925), .A2(n17919), .ZN(n15841) );
  NAND2_X1 U18964 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n17919), .ZN(
        n18039) );
  NOR2_X1 U18965 ( .A1(n17639), .A2(n18039), .ZN(n17980) );
  NOR2_X1 U18966 ( .A1(n15840), .A2(n15837), .ZN(n16458) );
  AOI21_X1 U18967 ( .B1(n17980), .B2(n16458), .A(n18692), .ZN(n15834) );
  AOI211_X1 U18968 ( .C1(n18699), .C2(n15841), .A(n15834), .B(n18220), .ZN(
        n15835) );
  AOI21_X1 U18969 ( .B1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18201) );
  NOR2_X1 U18970 ( .A1(n18201), .A2(n18049), .ZN(n18136) );
  NAND2_X1 U18971 ( .A1(n18050), .A2(n18136), .ZN(n18038) );
  NOR2_X1 U18972 ( .A1(n18024), .A2(n18038), .ZN(n17974) );
  INV_X1 U18973 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n17611) );
  NOR3_X1 U18974 ( .A1(n20983), .A2(n17611), .A3(n17964), .ZN(n17918) );
  NAND2_X1 U18975 ( .A1(n17974), .A2(n17918), .ZN(n17942) );
  NAND2_X1 U18976 ( .A1(n18710), .A2(n17942), .ZN(n17940) );
  OAI211_X1 U18977 ( .C1(n15836), .C2(n18203), .A(n15835), .B(n17940), .ZN(
        n15910) );
  AOI21_X1 U18978 ( .B1(n18109), .B2(n15837), .A(n15910), .ZN(n16450) );
  NAND2_X1 U18979 ( .A1(n18227), .A2(n18139), .ZN(n18140) );
  OAI22_X1 U18980 ( .A1(n18231), .A2(n16450), .B1(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n18140), .ZN(n15838) );
  INV_X1 U18981 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n18819) );
  NOR2_X1 U18982 ( .A1(n18218), .A2(n18819), .ZN(n16421) );
  AOI221_X1 U18983 ( .B1(n15911), .B2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), 
        .C1(n15838), .C2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A(n16421), .ZN(
        n15845) );
  INV_X1 U18984 ( .A(n17974), .ZN(n18017) );
  NOR2_X1 U18985 ( .A1(n18203), .A2(n18017), .ZN(n16455) );
  INV_X1 U18986 ( .A(n17980), .ZN(n15839) );
  NOR3_X1 U18987 ( .A1(n18692), .A2(n15840), .A3(n15839), .ZN(n15843) );
  INV_X1 U18988 ( .A(n18699), .ZN(n18714) );
  NOR2_X1 U18989 ( .A1(n18714), .A2(n15841), .ZN(n15842) );
  AOI211_X1 U18990 ( .C1(n17925), .C2(n16455), .A(n15843), .B(n15842), .ZN(
        n16438) );
  INV_X1 U18991 ( .A(n18083), .ZN(n18102) );
  AOI22_X1 U18992 ( .A1(n18681), .A2(n18058), .B1(n18048), .B2(n18102), .ZN(
        n16457) );
  INV_X1 U18993 ( .A(n17925), .ZN(n16409) );
  AOI211_X1 U18994 ( .C1(n16438), .C2(n16457), .A(n18214), .B(n16409), .ZN(
        n15909) );
  INV_X1 U18995 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16429) );
  NAND3_X1 U18996 ( .A1(n16426), .A2(n15909), .A3(n16429), .ZN(n15844) );
  OAI211_X1 U18997 ( .C1(n16434), .C2(n18123), .A(n15845), .B(n15844), .ZN(
        P3_U2833) );
  AOI21_X1 U18998 ( .B1(n15847), .B2(n15846), .A(n14314), .ZN(n19111) );
  AOI22_X1 U18999 ( .A1(n18995), .A2(n16340), .B1(n16344), .B2(n19111), .ZN(
        n15854) );
  XOR2_X1 U19000 ( .A(n15849), .B(n15848), .Z(n16239) );
  AOI22_X1 U19001 ( .A1(n16239), .A2(n16338), .B1(
        P2_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n15850), .ZN(n15853) );
  OR3_X1 U19002 ( .A1(n15851), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        n12221), .ZN(n15852) );
  NAND2_X1 U19003 ( .A1(P2_REIP_REG_16__SCAN_IN), .A2(n19245), .ZN(n16244) );
  NAND4_X1 U19004 ( .A1(n15854), .A2(n15853), .A3(n15852), .A4(n16244), .ZN(
        P2_U3030) );
  INV_X1 U19005 ( .A(n15855), .ZN(n16225) );
  AOI22_X1 U19006 ( .A1(n15856), .A2(n19097), .B1(n19088), .B2(n16225), .ZN(
        n15866) );
  AOI211_X1 U19007 ( .C1(n15858), .C2(n15857), .A(n9942), .B(n19809), .ZN(
        n15864) );
  INV_X1 U19008 ( .A(n15859), .ZN(n15862) );
  INV_X1 U19009 ( .A(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n15860) );
  OAI222_X1 U19010 ( .A1(n19095), .A2(n15862), .B1(n19074), .B2(n15861), .C1(
        n15860), .C2(n19057), .ZN(n15863) );
  AOI211_X1 U19011 ( .C1(n19090), .C2(P2_EBX_REG_22__SCAN_IN), .A(n15864), .B(
        n15863), .ZN(n15865) );
  NAND2_X1 U19012 ( .A1(n15866), .A2(n15865), .ZN(P2_U2833) );
  NOR3_X1 U19013 ( .A1(n15868), .A2(n15867), .A3(n20790), .ZN(n15873) );
  AOI211_X1 U19014 ( .C1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .C2(n15873), .A(
        n15870), .B(n15869), .ZN(n15871) );
  INV_X1 U19015 ( .A(n15871), .ZN(n15872) );
  OAI21_X1 U19016 ( .B1(n15873), .B2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(
        n15872), .ZN(n15874) );
  AOI222_X1 U19017 ( .A1(n15875), .A2(n20461), .B1(n15875), .B2(n15874), .C1(
        n20461), .C2(n15874), .ZN(n15876) );
  AOI222_X1 U19018 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n15877), 
        .B1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n15876), .C1(n15877), 
        .C2(n15876), .ZN(n15879) );
  AOI21_X1 U19019 ( .B1(n15879), .B2(n20152), .A(n15878), .ZN(n15888) );
  NOR2_X1 U19020 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(P1_MORE_REG_SCAN_IN), .ZN(
        n15883) );
  INV_X1 U19021 ( .A(n15880), .ZN(n15882) );
  OAI211_X1 U19022 ( .C1(n15884), .C2(n15883), .A(n15882), .B(n15881), .ZN(
        n15885) );
  INV_X1 U19023 ( .A(n15885), .ZN(n15886) );
  NAND3_X1 U19024 ( .A1(n15888), .A2(n15887), .A3(n15886), .ZN(n15896) );
  OAI21_X1 U19025 ( .B1(n20810), .B2(n15889), .A(n20695), .ZN(n15894) );
  NAND4_X1 U19026 ( .A1(n15892), .A2(n15891), .A3(n20801), .A4(n15890), .ZN(
        n15893) );
  NAND2_X1 U19027 ( .A1(n15894), .A2(n15893), .ZN(n16203) );
  NOR2_X1 U19028 ( .A1(n15895), .A2(n16208), .ZN(n20788) );
  AOI21_X1 U19029 ( .B1(n15897), .B2(n15896), .A(n20788), .ZN(n15899) );
  OAI211_X1 U19030 ( .C1(P1_STATE2_REG_2__SCAN_IN), .C2(n20810), .A(n15899), 
        .B(n15898), .ZN(n15900) );
  NOR2_X1 U19031 ( .A1(n16207), .A2(n15900), .ZN(n15905) );
  NAND2_X1 U19032 ( .A1(n15902), .A2(n15901), .ZN(n15903) );
  NAND2_X1 U19033 ( .A1(n20806), .A2(n15903), .ZN(n15904) );
  OAI22_X1 U19034 ( .A1(n15905), .A2(n20806), .B1(n16207), .B2(n15904), .ZN(
        P1_U3161) );
  NAND2_X1 U19035 ( .A1(n15907), .A2(n15906), .ZN(n15908) );
  XOR2_X1 U19036 ( .A(n15908), .B(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .Z(
        n16414) );
  NOR2_X1 U19037 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16436), .ZN(
        n16410) );
  AOI22_X1 U19038 ( .A1(n18231), .A2(P3_REIP_REG_30__SCAN_IN), .B1(n16410), 
        .B2(n15909), .ZN(n15914) );
  INV_X1 U19039 ( .A(n18140), .ZN(n18221) );
  AOI22_X1 U19040 ( .A1(n18221), .A2(n16436), .B1(n18218), .B2(n15910), .ZN(
        n16435) );
  INV_X1 U19041 ( .A(n16435), .ZN(n15912) );
  OAI21_X1 U19042 ( .B1(n15912), .B2(n15911), .A(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15913) );
  OAI211_X1 U19043 ( .C1(n18123), .C2(n16414), .A(n15914), .B(n15913), .ZN(
        P3_U2832) );
  INV_X1 U19044 ( .A(HOLD), .ZN(n19822) );
  INV_X1 U19045 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n20712) );
  NAND2_X1 U19046 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(n20712), .ZN(n20700) );
  AOI21_X1 U19047 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n20701), .A(n20801), 
        .ZN(n15916) );
  OAI211_X1 U19048 ( .C1(n20712), .C2(n19822), .A(P1_STATE_REG_0__SCAN_IN), 
        .B(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n15915) );
  OAI211_X1 U19049 ( .C1(n19822), .C2(n20700), .A(n15916), .B(n15915), .ZN(
        P1_U3195) );
  NOR2_X1 U19050 ( .A1(n19803), .A2(n19804), .ZN(n16394) );
  AOI221_X1 U19051 ( .B1(P2_STATEBS16_REG_SCAN_IN), .B2(
        P2_STATE2_REG_1__SCAN_IN), .C1(P2_STATE2_REG_0__SCAN_IN), .C2(
        P2_STATE2_REG_1__SCAN_IN), .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n15917)
         );
  NOR3_X1 U19052 ( .A1(n16394), .A2(n16403), .A3(n15917), .ZN(P2_U3178) );
  INV_X1 U19053 ( .A(n19925), .ZN(n19922) );
  NOR2_X1 U19054 ( .A1(n15918), .A2(n19922), .ZN(P2_U3047) );
  INV_X1 U19055 ( .A(n17420), .ZN(n17272) );
  NAND2_X1 U19056 ( .A1(n18277), .A2(n17272), .ZN(n17404) );
  INV_X1 U19057 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n17488) );
  NOR2_X1 U19058 ( .A1(n15922), .A2(n17420), .ZN(n17423) );
  AOI22_X1 U19059 ( .A1(n17423), .A2(BUF2_REG_0__SCAN_IN), .B1(n17422), .B2(
        n17898), .ZN(n15923) );
  OAI221_X1 U19060 ( .B1(P3_EAX_REG_0__SCAN_IN), .B2(n17404), .C1(n17488), 
        .C2(n17272), .A(n15923), .ZN(P3_U2735) );
  AOI221_X1 U19061 ( .B1(P1_REIP_REG_24__SCAN_IN), .B2(n15946), .C1(n20023), 
        .C2(n15946), .A(n15929), .ZN(n15926) );
  OAI22_X1 U19062 ( .A1(n15924), .A2(n20014), .B1(n20935), .B2(n19997), .ZN(
        n15925) );
  AOI211_X1 U19063 ( .C1(n20034), .C2(n15927), .A(n15926), .B(n15925), .ZN(
        n15933) );
  OR2_X1 U19064 ( .A1(n15928), .A2(n16023), .ZN(n15931) );
  NAND3_X1 U19065 ( .A1(n15935), .A2(P1_REIP_REG_24__SCAN_IN), .A3(n15929), 
        .ZN(n15930) );
  AND2_X1 U19066 ( .A1(n15931), .A2(n15930), .ZN(n15932) );
  OAI211_X1 U19067 ( .C1(n15934), .C2(n20038), .A(n15933), .B(n15932), .ZN(
        P1_U2815) );
  INV_X1 U19068 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n20743) );
  NAND2_X1 U19069 ( .A1(n15935), .A2(n20743), .ZN(n15940) );
  OAI22_X1 U19070 ( .A1(n15937), .A2(n20006), .B1(n15936), .B2(n19997), .ZN(
        n15938) );
  AOI21_X1 U19071 ( .B1(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n20026), .A(
        n15938), .ZN(n15939) );
  OAI211_X1 U19072 ( .C1(n20743), .C2(n15946), .A(n15940), .B(n15939), .ZN(
        n15941) );
  AOI21_X1 U19073 ( .B1(n15942), .B2(n19992), .A(n15941), .ZN(n15943) );
  OAI21_X1 U19074 ( .B1(n15944), .B2(n20038), .A(n15943), .ZN(P1_U2816) );
  AOI22_X1 U19075 ( .A1(n15945), .A2(n20034), .B1(P1_EBX_REG_23__SCAN_IN), 
        .B2(n20025), .ZN(n15953) );
  INV_X1 U19076 ( .A(n15946), .ZN(n15951) );
  OAI22_X1 U19077 ( .A1(n15948), .A2(n16023), .B1(n15947), .B2(n20038), .ZN(
        n15949) );
  OAI211_X1 U19078 ( .C1(n15954), .C2(n20014), .A(n15953), .B(n15952), .ZN(
        P1_U2817) );
  INV_X1 U19079 ( .A(n15955), .ZN(n16040) );
  INV_X1 U19080 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n20739) );
  NOR3_X1 U19081 ( .A1(P1_REIP_REG_22__SCAN_IN), .A2(n15959), .A3(n20739), 
        .ZN(n15958) );
  AOI22_X1 U19082 ( .A1(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n20026), .B1(
        P1_EBX_REG_22__SCAN_IN), .B2(n20025), .ZN(n15956) );
  OAI21_X1 U19083 ( .B1(n16043), .B2(n20006), .A(n15956), .ZN(n15957) );
  AOI211_X1 U19084 ( .C1(n16040), .C2(n19992), .A(n15958), .B(n15957), .ZN(
        n15963) );
  NOR2_X1 U19085 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(n15959), .ZN(n15969) );
  OAI21_X1 U19086 ( .B1(n16020), .B2(n15961), .A(n15960), .ZN(n15976) );
  OAI21_X1 U19087 ( .B1(n15969), .B2(n15976), .A(P1_REIP_REG_22__SCAN_IN), 
        .ZN(n15962) );
  OAI211_X1 U19088 ( .C1(n15964), .C2(n20038), .A(n15963), .B(n15962), .ZN(
        P1_U2818) );
  AOI22_X1 U19089 ( .A1(n15965), .A2(n20034), .B1(P1_EBX_REG_21__SCAN_IN), 
        .B2(n20025), .ZN(n15971) );
  OAI22_X1 U19090 ( .A1(n15967), .A2(n16023), .B1(n15966), .B2(n20038), .ZN(
        n15968) );
  AOI211_X1 U19091 ( .C1(P1_REIP_REG_21__SCAN_IN), .C2(n15976), .A(n15969), 
        .B(n15968), .ZN(n15970) );
  OAI211_X1 U19092 ( .C1(n15972), .C2(n20014), .A(n15971), .B(n15970), .ZN(
        P1_U2819) );
  INV_X1 U19093 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n15973) );
  OAI22_X1 U19094 ( .A1(n15973), .A2(n20014), .B1(n16048), .B2(n20006), .ZN(
        n15974) );
  AOI21_X1 U19095 ( .B1(P1_EBX_REG_20__SCAN_IN), .B2(n20025), .A(n15974), .ZN(
        n15979) );
  INV_X1 U19096 ( .A(P1_REIP_REG_20__SCAN_IN), .ZN(n20736) );
  OAI21_X1 U19097 ( .B1(n15975), .B2(n15984), .A(n20736), .ZN(n15977) );
  AOI22_X1 U19098 ( .A1(n16044), .A2(n19992), .B1(n15977), .B2(n15976), .ZN(
        n15978) );
  OAI211_X1 U19099 ( .C1(n20038), .C2(n15980), .A(n15979), .B(n15978), .ZN(
        P1_U2820) );
  INV_X1 U19100 ( .A(n20011), .ZN(n19990) );
  OAI22_X1 U19101 ( .A1(n16056), .A2(n20006), .B1(n15981), .B2(n19997), .ZN(
        n15982) );
  AOI211_X1 U19102 ( .C1(n20026), .C2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n19990), .B(n15982), .ZN(n15988) );
  INV_X1 U19103 ( .A(n15983), .ZN(n16053) );
  INV_X1 U19104 ( .A(P1_REIP_REG_18__SCAN_IN), .ZN(n20733) );
  NAND2_X1 U19105 ( .A1(n20733), .A2(n15984), .ZN(n15986) );
  AOI22_X1 U19106 ( .A1(n16053), .A2(n19992), .B1(n15986), .B2(n15985), .ZN(
        n15987) );
  OAI211_X1 U19107 ( .C1(n20038), .C2(n16116), .A(n15988), .B(n15987), .ZN(
        P1_U2822) );
  AOI22_X1 U19108 ( .A1(P1_EBX_REG_16__SCAN_IN), .A2(n20025), .B1(
        P1_REIP_REG_16__SCAN_IN), .B2(n16007), .ZN(n15989) );
  OAI21_X1 U19109 ( .B1(n16061), .B2(n20006), .A(n15989), .ZN(n15990) );
  AOI211_X1 U19110 ( .C1(n20026), .C2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n19990), .B(n15990), .ZN(n15994) );
  INV_X1 U19111 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n20730) );
  AOI21_X1 U19112 ( .B1(n15055), .B2(n20730), .A(n16004), .ZN(n15992) );
  AOI22_X1 U19113 ( .A1(n16058), .A2(n19992), .B1(n15992), .B2(n15991), .ZN(
        n15993) );
  OAI211_X1 U19114 ( .C1(n20038), .C2(n15995), .A(n15994), .B(n15993), .ZN(
        P1_U2824) );
  INV_X1 U19115 ( .A(n15996), .ZN(n16132) );
  AOI22_X1 U19116 ( .A1(n15997), .A2(n20034), .B1(n20010), .B2(n16132), .ZN(
        n16003) );
  AOI22_X1 U19117 ( .A1(P1_EBX_REG_15__SCAN_IN), .A2(n20025), .B1(
        P1_REIP_REG_15__SCAN_IN), .B2(n16007), .ZN(n15998) );
  OAI211_X1 U19118 ( .C1(n15999), .C2(n20014), .A(n15998), .B(n20011), .ZN(
        n16000) );
  AOI21_X1 U19119 ( .B1(n16001), .B2(n19992), .A(n16000), .ZN(n16002) );
  OAI211_X1 U19120 ( .C1(P1_REIP_REG_15__SCAN_IN), .C2(n16004), .A(n16003), 
        .B(n16002), .ZN(P1_U2825) );
  OAI22_X1 U19121 ( .A1(n16005), .A2(n19997), .B1(n20038), .B2(n16137), .ZN(
        n16006) );
  AOI211_X1 U19122 ( .C1(n20026), .C2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n19990), .B(n16006), .ZN(n16011) );
  AOI22_X1 U19123 ( .A1(n16069), .A2(n19992), .B1(n20034), .B2(n16068), .ZN(
        n16010) );
  OAI21_X1 U19124 ( .B1(P1_REIP_REG_14__SCAN_IN), .B2(n16008), .A(n16007), 
        .ZN(n16009) );
  NAND3_X1 U19125 ( .A1(n16011), .A2(n16010), .A3(n16009), .ZN(P1_U2826) );
  OAI22_X1 U19126 ( .A1(n16012), .A2(n19997), .B1(n20038), .B2(n16160), .ZN(
        n16013) );
  AOI211_X1 U19127 ( .C1(n20026), .C2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n19990), .B(n16013), .ZN(n16017) );
  INV_X1 U19128 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n20725) );
  INV_X1 U19129 ( .A(P1_REIP_REG_12__SCAN_IN), .ZN(n20997) );
  OAI21_X1 U19130 ( .B1(n20725), .B2(n16027), .A(n20997), .ZN(n16014) );
  AOI22_X1 U19131 ( .A1(n16076), .A2(n20034), .B1(n16015), .B2(n16014), .ZN(
        n16016) );
  OAI211_X1 U19132 ( .C1(n16023), .C2(n16018), .A(n16017), .B(n16016), .ZN(
        P1_U2828) );
  INV_X1 U19133 ( .A(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n21151) );
  NOR2_X1 U19134 ( .A1(n16020), .A2(n16019), .ZN(n16032) );
  AOI22_X1 U19135 ( .A1(n20010), .A2(n16167), .B1(P1_REIP_REG_11__SCAN_IN), 
        .B2(n16032), .ZN(n16021) );
  OAI211_X1 U19136 ( .C1(n20014), .C2(n21151), .A(n16021), .B(n20011), .ZN(
        n16025) );
  OAI22_X1 U19137 ( .A1(n16088), .A2(n20006), .B1(n16023), .B2(n16022), .ZN(
        n16024) );
  AOI211_X1 U19138 ( .C1(P1_EBX_REG_11__SCAN_IN), .C2(n20025), .A(n16025), .B(
        n16024), .ZN(n16026) );
  OAI21_X1 U19139 ( .B1(P1_REIP_REG_11__SCAN_IN), .B2(n16027), .A(n16026), 
        .ZN(P1_U2829) );
  NAND2_X1 U19140 ( .A1(n19970), .A2(P1_REIP_REG_9__SCAN_IN), .ZN(n16038) );
  OAI21_X1 U19141 ( .B1(n20014), .B2(n21019), .A(n20011), .ZN(n16031) );
  OAI22_X1 U19142 ( .A1(n16029), .A2(n19997), .B1(n20038), .B2(n16028), .ZN(
        n16030) );
  AOI211_X1 U19143 ( .C1(P1_REIP_REG_10__SCAN_IN), .C2(n16032), .A(n16031), 
        .B(n16030), .ZN(n16037) );
  INV_X1 U19144 ( .A(n16033), .ZN(n16034) );
  AOI22_X1 U19145 ( .A1(n16035), .A2(n19992), .B1(n16034), .B2(n20034), .ZN(
        n16036) );
  OAI211_X1 U19146 ( .C1(P1_REIP_REG_10__SCAN_IN), .C2(n16038), .A(n16037), 
        .B(n16036), .ZN(P1_U2830) );
  AOI22_X1 U19147 ( .A1(n20091), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B1(
        n20103), .B2(P1_REIP_REG_22__SCAN_IN), .ZN(n16042) );
  AOI22_X1 U19148 ( .A1(n16040), .A2(n20097), .B1(n20098), .B2(n16039), .ZN(
        n16041) );
  OAI211_X1 U19149 ( .C1(n20102), .C2(n16043), .A(n16042), .B(n16041), .ZN(
        P1_U2977) );
  AOI22_X1 U19150 ( .A1(n20091), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B1(
        n20103), .B2(P1_REIP_REG_20__SCAN_IN), .ZN(n16047) );
  AOI22_X1 U19151 ( .A1(n16045), .A2(n20098), .B1(n20097), .B2(n16044), .ZN(
        n16046) );
  OAI211_X1 U19152 ( .C1(n20102), .C2(n16048), .A(n16047), .B(n16046), .ZN(
        P1_U2979) );
  AOI22_X1 U19153 ( .A1(n20091), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B1(
        n20103), .B2(P1_REIP_REG_18__SCAN_IN), .ZN(n16055) );
  INV_X1 U19154 ( .A(n16049), .ZN(n16052) );
  AOI21_X1 U19155 ( .B1(n16052), .B2(n10148), .A(n16051), .ZN(n16120) );
  AOI22_X1 U19156 ( .A1(n16120), .A2(n20098), .B1(n20097), .B2(n16053), .ZN(
        n16054) );
  OAI211_X1 U19157 ( .C1(n20102), .C2(n16056), .A(n16055), .B(n16054), .ZN(
        P1_U2981) );
  AOI22_X1 U19158 ( .A1(n20091), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B1(
        n20103), .B2(P1_REIP_REG_16__SCAN_IN), .ZN(n16060) );
  AOI22_X1 U19159 ( .A1(n16058), .A2(n20097), .B1(n20098), .B2(n16057), .ZN(
        n16059) );
  OAI211_X1 U19160 ( .C1(n20102), .C2(n16061), .A(n16060), .B(n16059), .ZN(
        P1_U2983) );
  INV_X1 U19161 ( .A(n16062), .ZN(n16063) );
  AOI21_X1 U19162 ( .B1(n16065), .B2(n16064), .A(n16063), .ZN(n16067) );
  AOI22_X1 U19163 ( .A1(n16081), .A2(n16143), .B1(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n9913), .ZN(n16066) );
  XNOR2_X1 U19164 ( .A(n16067), .B(n16066), .ZN(n16138) );
  AOI22_X1 U19165 ( .A1(n20091), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(
        n20103), .B2(P1_REIP_REG_14__SCAN_IN), .ZN(n16071) );
  AOI22_X1 U19166 ( .A1(n16069), .A2(n20097), .B1(n16077), .B2(n16068), .ZN(
        n16070) );
  OAI211_X1 U19167 ( .C1(n16138), .C2(n19949), .A(n16071), .B(n16070), .ZN(
        P1_U2985) );
  AOI21_X1 U19168 ( .B1(n16074), .B2(n16073), .A(n16072), .ZN(n16166) );
  AOI22_X1 U19169 ( .A1(n20091), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        n20103), .B2(P1_REIP_REG_12__SCAN_IN), .ZN(n16079) );
  AOI22_X1 U19170 ( .A1(n16077), .A2(n16076), .B1(n20097), .B2(n16075), .ZN(
        n16078) );
  OAI211_X1 U19171 ( .C1(n16166), .C2(n19949), .A(n16079), .B(n16078), .ZN(
        P1_U2987) );
  AOI22_X1 U19172 ( .A1(n20091), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B1(
        n20103), .B2(P1_REIP_REG_11__SCAN_IN), .ZN(n16087) );
  NOR3_X1 U19173 ( .A1(n14891), .A2(n16081), .A3(n16080), .ZN(n16083) );
  NOR2_X1 U19174 ( .A1(n16083), .A2(n16082), .ZN(n16084) );
  XNOR2_X1 U19175 ( .A(n16084), .B(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n16169) );
  AOI22_X1 U19176 ( .A1(n20098), .A2(n16169), .B1(n20097), .B2(n16085), .ZN(
        n16086) );
  OAI211_X1 U19177 ( .C1(n20102), .C2(n16088), .A(n16087), .B(n16086), .ZN(
        P1_U2988) );
  AOI22_X1 U19178 ( .A1(n20091), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B1(
        n20103), .B2(P1_REIP_REG_7__SCAN_IN), .ZN(n16094) );
  NAND2_X1 U19179 ( .A1(n16091), .A2(n16090), .ZN(n16092) );
  XNOR2_X1 U19180 ( .A(n16089), .B(n16092), .ZN(n16187) );
  AOI22_X1 U19181 ( .A1(n16187), .A2(n20098), .B1(n20097), .B2(n19982), .ZN(
        n16093) );
  OAI211_X1 U19182 ( .C1(n20102), .C2(n19985), .A(n16094), .B(n16093), .ZN(
        P1_U2992) );
  AOI22_X1 U19183 ( .A1(n20091), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B1(
        n20103), .B2(P1_REIP_REG_6__SCAN_IN), .ZN(n16097) );
  AOI22_X1 U19184 ( .A1(n16095), .A2(n20098), .B1(n20097), .B2(n19993), .ZN(
        n16096) );
  OAI211_X1 U19185 ( .C1(n20102), .C2(n19996), .A(n16097), .B(n16096), .ZN(
        P1_U2993) );
  AOI22_X1 U19186 ( .A1(n20091), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .B1(
        n20103), .B2(P1_REIP_REG_5__SCAN_IN), .ZN(n16103) );
  OAI21_X1 U19187 ( .B1(n16100), .B2(n16099), .A(n16098), .ZN(n16101) );
  INV_X1 U19188 ( .A(n16101), .ZN(n16196) );
  AOI22_X1 U19189 ( .A1(n16196), .A2(n20098), .B1(n20097), .B2(n20004), .ZN(
        n16102) );
  OAI211_X1 U19190 ( .C1(n20102), .C2(n20007), .A(n16103), .B(n16102), .ZN(
        P1_U2994) );
  INV_X1 U19191 ( .A(P1_REIP_REG_19__SCAN_IN), .ZN(n16114) );
  INV_X1 U19192 ( .A(n16104), .ZN(n16107) );
  INV_X1 U19193 ( .A(n16105), .ZN(n16106) );
  AOI22_X1 U19194 ( .A1(n16107), .A2(n20137), .B1(n20114), .B2(n16106), .ZN(
        n16113) );
  INV_X1 U19195 ( .A(n16108), .ZN(n16110) );
  AOI22_X1 U19196 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n16111), .B1(
        n16110), .B2(n16109), .ZN(n16112) );
  OAI211_X1 U19197 ( .C1(n16114), .C2(n20128), .A(n16113), .B(n16112), .ZN(
        P1_U3012) );
  INV_X1 U19198 ( .A(n16115), .ZN(n20140) );
  AOI21_X1 U19199 ( .B1(n20140), .B2(n16117), .A(n16148), .ZN(n16130) );
  NAND2_X1 U19200 ( .A1(n16140), .A2(n16123), .ZN(n16118) );
  OAI22_X1 U19201 ( .A1(n16118), .A2(n16117), .B1(n20145), .B2(n16116), .ZN(
        n16119) );
  AOI21_X1 U19202 ( .B1(n16120), .B2(n20137), .A(n16119), .ZN(n16122) );
  NAND2_X1 U19203 ( .A1(n20103), .A2(P1_REIP_REG_18__SCAN_IN), .ZN(n16121) );
  OAI211_X1 U19204 ( .C1(n16130), .C2(n16123), .A(n16122), .B(n16121), .ZN(
        P1_U3013) );
  AOI21_X1 U19205 ( .B1(n16124), .B2(n16140), .A(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n16129) );
  AOI22_X1 U19206 ( .A1(n16126), .A2(n20137), .B1(n20114), .B2(n16125), .ZN(
        n16128) );
  NAND2_X1 U19207 ( .A1(n20103), .A2(P1_REIP_REG_17__SCAN_IN), .ZN(n16127) );
  OAI211_X1 U19208 ( .C1(n16130), .C2(n16129), .A(n16128), .B(n16127), .ZN(
        P1_U3014) );
  AOI22_X1 U19209 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n16131), .B1(
        n20103), .B2(P1_REIP_REG_15__SCAN_IN), .ZN(n16135) );
  AOI22_X1 U19210 ( .A1(n16133), .A2(n20137), .B1(n20114), .B2(n16132), .ZN(
        n16134) );
  OAI211_X1 U19211 ( .C1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n16136), .A(
        n16135), .B(n16134), .ZN(P1_U3016) );
  OAI22_X1 U19212 ( .A1(n16138), .A2(n16177), .B1(n20145), .B2(n16137), .ZN(
        n16139) );
  AOI21_X1 U19213 ( .B1(n16140), .B2(n16143), .A(n16139), .ZN(n16142) );
  NAND2_X1 U19214 ( .A1(n20103), .A2(P1_REIP_REG_14__SCAN_IN), .ZN(n16141) );
  OAI211_X1 U19215 ( .C1(n16144), .C2(n16143), .A(n16142), .B(n16141), .ZN(
        P1_U3017) );
  INV_X1 U19216 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n21141) );
  NAND3_X1 U19217 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A3(n21141), .ZN(n16151) );
  AOI21_X1 U19218 ( .B1(n16146), .B2(n20114), .A(n16145), .ZN(n16150) );
  AOI22_X1 U19219 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n16148), .B1(
        n20137), .B2(n16147), .ZN(n16149) );
  OAI211_X1 U19220 ( .C1(n16152), .C2(n16151), .A(n16150), .B(n16149), .ZN(
        P1_U3018) );
  NOR3_X1 U19221 ( .A1(n12643), .A2(n16154), .A3(n16180), .ZN(n16164) );
  INV_X1 U19222 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n16163) );
  INV_X1 U19223 ( .A(n16153), .ZN(n16159) );
  INV_X1 U19224 ( .A(n16154), .ZN(n16155) );
  AOI21_X1 U19225 ( .B1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n16155), .A(
        n20121), .ZN(n16157) );
  AOI211_X1 U19226 ( .C1(n20125), .C2(n16158), .A(n16157), .B(n16156), .ZN(
        n16174) );
  OAI21_X1 U19227 ( .B1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n16159), .A(
        n16174), .ZN(n16162) );
  OAI22_X1 U19228 ( .A1(n16160), .A2(n20145), .B1(n20997), .B2(n20128), .ZN(
        n16161) );
  AOI221_X1 U19229 ( .B1(n16164), .B2(n16163), .C1(n16162), .C2(
        P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A(n16161), .ZN(n16165) );
  OAI21_X1 U19230 ( .B1(n16166), .B2(n16177), .A(n16165), .ZN(P1_U3019) );
  AOI22_X1 U19231 ( .A1(n16167), .A2(n20114), .B1(n20103), .B2(
        P1_REIP_REG_11__SCAN_IN), .ZN(n16173) );
  NOR2_X1 U19232 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n16168), .ZN(
        n16170) );
  AOI22_X1 U19233 ( .A1(n16171), .A2(n16170), .B1(n20137), .B2(n16169), .ZN(
        n16172) );
  OAI211_X1 U19234 ( .C1(n16174), .C2(n12643), .A(n16173), .B(n16172), .ZN(
        P1_U3020) );
  AOI21_X1 U19235 ( .B1(n16181), .B2(n20140), .A(n16175), .ZN(n16190) );
  OAI222_X1 U19236 ( .A1(n16178), .A2(n20145), .B1(n20128), .B2(n20721), .C1(
        n16177), .C2(n16176), .ZN(n16179) );
  INV_X1 U19237 ( .A(n16179), .ZN(n16183) );
  NOR2_X1 U19238 ( .A1(n16181), .A2(n16180), .ZN(n16186) );
  OAI221_X1 U19239 ( .B1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .C1(n16184), .C2(n16191), .A(
        n16186), .ZN(n16182) );
  OAI211_X1 U19240 ( .C1(n16190), .C2(n16184), .A(n16183), .B(n16182), .ZN(
        P1_U3023) );
  INV_X1 U19241 ( .A(n16185), .ZN(n19974) );
  AOI22_X1 U19242 ( .A1(n20114), .A2(n19974), .B1(n20103), .B2(
        P1_REIP_REG_7__SCAN_IN), .ZN(n16189) );
  AOI22_X1 U19243 ( .A1(n16187), .A2(n20137), .B1(n16186), .B2(n16191), .ZN(
        n16188) );
  OAI211_X1 U19244 ( .C1(n16191), .C2(n16190), .A(n16189), .B(n16188), .ZN(
        P1_U3024) );
  INV_X1 U19245 ( .A(P1_REIP_REG_5__SCAN_IN), .ZN(n16192) );
  OAI22_X1 U19246 ( .A1(n20145), .A2(n16193), .B1(n20128), .B2(n16192), .ZN(
        n16194) );
  INV_X1 U19247 ( .A(n16194), .ZN(n16198) );
  AOI22_X1 U19248 ( .A1(n16196), .A2(n20137), .B1(n16195), .B2(n20107), .ZN(
        n16197) );
  OAI211_X1 U19249 ( .C1(n16200), .C2(n16199), .A(n16198), .B(n16197), .ZN(
        P1_U3026) );
  NAND4_X1 U19250 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(
        P1_STATE2_REG_1__SCAN_IN), .A3(n20802), .A4(n20810), .ZN(n16201) );
  OAI21_X1 U19251 ( .B1(n16202), .B2(n20208), .A(n16201), .ZN(n20694) );
  OAI21_X1 U19252 ( .B1(n16204), .B2(n20694), .A(n16203), .ZN(n16205) );
  OAI221_X1 U19253 ( .B1(n20807), .B2(n20413), .C1(n20807), .C2(n20810), .A(
        n16205), .ZN(n16206) );
  AOI221_X1 U19254 ( .B1(n16207), .B2(n13782), .C1(n20806), .C2(n13782), .A(
        n16206), .ZN(P1_U3162) );
  NOR2_X1 U19255 ( .A1(n16207), .A2(n20806), .ZN(n16209) );
  OAI22_X1 U19256 ( .A1(n20413), .A2(n16209), .B1(n16208), .B2(n20806), .ZN(
        P1_U3466) );
  AOI22_X1 U19257 ( .A1(P2_EBX_REG_26__SCAN_IN), .A2(n19090), .B1(
        P2_REIP_REG_26__SCAN_IN), .B2(n19091), .ZN(n16223) );
  OAI22_X1 U19258 ( .A1(n16211), .A2(n19095), .B1(n16210), .B2(n19057), .ZN(
        n16212) );
  INV_X1 U19259 ( .A(n16212), .ZN(n16222) );
  INV_X1 U19260 ( .A(n16213), .ZN(n16214) );
  AOI22_X1 U19261 ( .A1(n16215), .A2(n19097), .B1(n16214), .B2(n19088), .ZN(
        n16221) );
  AOI21_X1 U19262 ( .B1(n16218), .B2(n16217), .A(n16216), .ZN(n16219) );
  NAND2_X1 U19263 ( .A1(n9868), .A2(n16219), .ZN(n16220) );
  NAND4_X1 U19264 ( .A1(n16223), .A2(n16222), .A3(n16221), .A4(n16220), .ZN(
        P2_U2829) );
  AOI22_X1 U19265 ( .A1(n19108), .A2(n16224), .B1(n19155), .B2(
        P2_EAX_REG_22__SCAN_IN), .ZN(n16229) );
  AOI22_X1 U19266 ( .A1(n19110), .A2(BUF1_REG_22__SCAN_IN), .B1(n19109), .B2(
        BUF2_REG_22__SCAN_IN), .ZN(n16228) );
  AOI22_X1 U19267 ( .A1(n16226), .A2(n19116), .B1(n19156), .B2(n16225), .ZN(
        n16227) );
  NAND3_X1 U19268 ( .A1(n16229), .A2(n16228), .A3(n16227), .ZN(P2_U2897) );
  AOI22_X1 U19269 ( .A1(n19108), .A2(n19282), .B1(n19155), .B2(
        P2_EAX_REG_20__SCAN_IN), .ZN(n16233) );
  AOI22_X1 U19270 ( .A1(n19110), .A2(BUF1_REG_20__SCAN_IN), .B1(n19109), .B2(
        BUF2_REG_20__SCAN_IN), .ZN(n16232) );
  AOI22_X1 U19271 ( .A1(n16230), .A2(n19116), .B1(n19156), .B2(n18951), .ZN(
        n16231) );
  NAND3_X1 U19272 ( .A1(n16233), .A2(n16232), .A3(n16231), .ZN(P2_U2899) );
  AOI22_X1 U19273 ( .A1(n19108), .A2(n16234), .B1(n19155), .B2(
        P2_EAX_REG_18__SCAN_IN), .ZN(n16238) );
  AOI22_X1 U19274 ( .A1(n19110), .A2(BUF1_REG_18__SCAN_IN), .B1(n19109), .B2(
        BUF2_REG_18__SCAN_IN), .ZN(n16237) );
  AOI22_X1 U19275 ( .A1(n16235), .A2(n19116), .B1(n19156), .B2(n18972), .ZN(
        n16236) );
  NAND3_X1 U19276 ( .A1(n16238), .A2(n16237), .A3(n16236), .ZN(P2_U2901) );
  AOI22_X1 U19277 ( .A1(n19246), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B1(
        n16302), .B2(n18991), .ZN(n16246) );
  AOI22_X1 U19278 ( .A1(n16239), .A2(n19248), .B1(n19250), .B2(n18995), .ZN(
        n16245) );
  INV_X1 U19279 ( .A(n16240), .ZN(n16242) );
  OAI211_X1 U19280 ( .C1(n16242), .C2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n19251), .B(n16241), .ZN(n16243) );
  NAND4_X1 U19281 ( .A1(n16246), .A2(n16245), .A3(n16244), .A4(n16243), .ZN(
        P2_U2998) );
  AOI22_X1 U19282 ( .A1(n19246), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(
        P2_REIP_REG_14__SCAN_IN), .B2(n19245), .ZN(n16250) );
  AOI222_X1 U19283 ( .A1(n16248), .A2(n19248), .B1(n19250), .B2(n19020), .C1(
        n19251), .C2(n16247), .ZN(n16249) );
  AOI22_X1 U19284 ( .A1(n19246), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        P2_REIP_REG_12__SCAN_IN), .B2(n19038), .ZN(n16257) );
  INV_X1 U19285 ( .A(n16251), .ZN(n16255) );
  INV_X1 U19286 ( .A(n16252), .ZN(n16253) );
  AOI222_X1 U19287 ( .A1(n16255), .A2(n19251), .B1(n19248), .B2(n16254), .C1(
        n19250), .C2(n16253), .ZN(n16256) );
  OAI211_X1 U19288 ( .C1(n19256), .C2(n16258), .A(n16257), .B(n16256), .ZN(
        P2_U3002) );
  AOI22_X1 U19289 ( .A1(P2_REIP_REG_11__SCAN_IN), .A2(n19245), .B1(n16302), 
        .B2(n16259), .ZN(n16265) );
  OAI22_X1 U19290 ( .A1(n16261), .A2(n16295), .B1(n16260), .B2(n16293), .ZN(
        n16262) );
  AOI21_X1 U19291 ( .B1(n19250), .B2(n16263), .A(n16262), .ZN(n16264) );
  OAI211_X1 U19292 ( .C1(n16310), .C2(n16266), .A(n16265), .B(n16264), .ZN(
        P2_U3003) );
  AOI22_X1 U19293 ( .A1(n19246), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B1(
        P2_REIP_REG_10__SCAN_IN), .B2(n19245), .ZN(n16270) );
  AOI222_X1 U19294 ( .A1(n16268), .A2(n19248), .B1(n19250), .B2(n19042), .C1(
        n19251), .C2(n16267), .ZN(n16269) );
  OAI211_X1 U19295 ( .C1(n19256), .C2(n19040), .A(n16270), .B(n16269), .ZN(
        P2_U3004) );
  AOI22_X1 U19296 ( .A1(P2_REIP_REG_9__SCAN_IN), .A2(n19038), .B1(n16302), 
        .B2(n16271), .ZN(n16277) );
  OAI22_X1 U19297 ( .A1(n16273), .A2(n16295), .B1(n16293), .B2(n16272), .ZN(
        n16274) );
  AOI21_X1 U19298 ( .B1(n19250), .B2(n16275), .A(n16274), .ZN(n16276) );
  OAI211_X1 U19299 ( .C1(n16310), .C2(n16278), .A(n16277), .B(n16276), .ZN(
        P2_U3005) );
  AOI22_X1 U19300 ( .A1(n19246), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B1(
        P2_REIP_REG_8__SCAN_IN), .B2(n19038), .ZN(n16291) );
  NAND2_X1 U19301 ( .A1(n16280), .A2(n16279), .ZN(n16286) );
  INV_X1 U19302 ( .A(n16281), .ZN(n16282) );
  AOI21_X1 U19303 ( .B1(n16284), .B2(n16283), .A(n16282), .ZN(n16285) );
  XOR2_X1 U19304 ( .A(n16286), .B(n16285), .Z(n16330) );
  XOR2_X1 U19305 ( .A(n16287), .B(n16288), .Z(n16324) );
  AOI222_X1 U19306 ( .A1(n16330), .A2(n19248), .B1(n19250), .B2(n16289), .C1(
        n19251), .C2(n16324), .ZN(n16290) );
  OAI211_X1 U19307 ( .C1(n19256), .C2(n16292), .A(n16291), .B(n16290), .ZN(
        P2_U3006) );
  AOI22_X1 U19308 ( .A1(P2_REIP_REG_5__SCAN_IN), .A2(n19245), .B1(n16302), 
        .B2(n19081), .ZN(n16299) );
  OAI22_X1 U19309 ( .A1(n16296), .A2(n16295), .B1(n16294), .B2(n16293), .ZN(
        n16297) );
  AOI21_X1 U19310 ( .B1(n19250), .B2(n19082), .A(n16297), .ZN(n16298) );
  OAI211_X1 U19311 ( .C1(n16310), .C2(n16300), .A(n16299), .B(n16298), .ZN(
        P2_U3009) );
  AOI22_X1 U19312 ( .A1(P2_REIP_REG_3__SCAN_IN), .A2(n19245), .B1(n16302), 
        .B2(n16301), .ZN(n16309) );
  NAND3_X1 U19313 ( .A1(n16303), .A2(n14102), .A3(n19251), .ZN(n16304) );
  OAI21_X1 U19314 ( .B1(n16305), .B2(n13842), .A(n16304), .ZN(n16306) );
  AOI21_X1 U19315 ( .B1(n16307), .B2(n19248), .A(n16306), .ZN(n16308) );
  OAI211_X1 U19316 ( .C1(n11328), .C2(n16310), .A(n16309), .B(n16308), .ZN(
        P2_U3011) );
  INV_X1 U19317 ( .A(n16311), .ZN(n16315) );
  OAI21_X1 U19318 ( .B1(n16312), .B2(n15632), .A(n15846), .ZN(n19118) );
  OAI22_X1 U19319 ( .A1(n16313), .A2(n19118), .B1(n15437), .B2(n12458), .ZN(
        n16314) );
  AOI221_X1 U19320 ( .B1(n16316), .B2(n12221), .C1(n16315), .C2(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(n16314), .ZN(n16320) );
  OAI22_X1 U19321 ( .A1(n16317), .A2(n16327), .B1(n16326), .B2(n19005), .ZN(
        n16318) );
  INV_X1 U19322 ( .A(n16318), .ZN(n16319) );
  OAI211_X1 U19323 ( .C1(n16322), .C2(n16321), .A(n16320), .B(n16319), .ZN(
        P2_U3031) );
  AOI22_X1 U19324 ( .A1(n16323), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .B1(
        n16344), .B2(n19135), .ZN(n16336) );
  INV_X1 U19325 ( .A(n16324), .ZN(n16328) );
  OAI22_X1 U19326 ( .A1(n16328), .A2(n16327), .B1(n16326), .B2(n16325), .ZN(
        n16329) );
  AOI21_X1 U19327 ( .B1(n16338), .B2(n16330), .A(n16329), .ZN(n16335) );
  NAND2_X1 U19328 ( .A1(P2_REIP_REG_8__SCAN_IN), .A2(n19038), .ZN(n16334) );
  OAI211_X1 U19329 ( .C1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A(n16332), .B(n16331), .ZN(n16333) );
  NAND4_X1 U19330 ( .A1(n16336), .A2(n16335), .A3(n16334), .A4(n16333), .ZN(
        P2_U3038) );
  AOI22_X1 U19331 ( .A1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n16339), .B1(
        n16338), .B2(n16337), .ZN(n16350) );
  NAND2_X1 U19332 ( .A1(n16340), .A2(n19098), .ZN(n16348) );
  NAND2_X1 U19333 ( .A1(n16342), .A2(n16341), .ZN(n16346) );
  INV_X1 U19334 ( .A(n16343), .ZN(n19089) );
  NAND2_X1 U19335 ( .A1(n16344), .A2(n19089), .ZN(n16345) );
  AND4_X1 U19336 ( .A1(n16348), .A2(n16347), .A3(n16346), .A4(n16345), .ZN(
        n16349) );
  OAI211_X1 U19337 ( .C1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(n16351), .A(
        n16350), .B(n16349), .ZN(P2_U3046) );
  MUX2_X1 U19338 ( .A(n15752), .B(n16358), .S(n16354), .Z(n16382) );
  MUX2_X1 U19339 ( .A(n11651), .B(n16357), .S(n16354), .Z(n16381) );
  INV_X1 U19340 ( .A(n16353), .ZN(n16356) );
  OAI211_X1 U19341 ( .C1(n16353), .C2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B(n16352), .ZN(n16355) );
  OAI211_X1 U19342 ( .C1(n16356), .C2(n19914), .A(n16355), .B(n16354), .ZN(
        n16361) );
  INV_X1 U19343 ( .A(n16357), .ZN(n16359) );
  OAI22_X1 U19344 ( .A1(n16359), .A2(n19898), .B1(n19905), .B2(n16358), .ZN(
        n16360) );
  OAI22_X1 U19345 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n16381), .B1(
        n16361), .B2(n16360), .ZN(n16362) );
  AOI21_X1 U19346 ( .B1(n19354), .B2(n16382), .A(n16362), .ZN(n16386) );
  AOI22_X1 U19347 ( .A1(n16365), .A2(n16364), .B1(n11616), .B2(n16363), .ZN(
        n16369) );
  NAND2_X1 U19348 ( .A1(n16367), .A2(n16366), .ZN(n16368) );
  AND2_X1 U19349 ( .A1(n16369), .A2(n16368), .ZN(n19932) );
  NAND2_X1 U19350 ( .A1(n16371), .A2(n16370), .ZN(n16378) );
  AND3_X1 U19351 ( .A1(n16374), .A2(n16373), .A3(n16372), .ZN(n16375) );
  AND2_X1 U19352 ( .A1(n11616), .A2(n16375), .ZN(n18915) );
  OAI21_X1 U19353 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(P2_MORE_REG_SCAN_IN), .A(
        n18915), .ZN(n16377) );
  NAND4_X1 U19354 ( .A1(n19932), .A2(n16378), .A3(n16377), .A4(n16376), .ZN(
        n16379) );
  AOI21_X1 U19355 ( .B1(n16380), .B2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(
        n16379), .ZN(n16385) );
  INV_X1 U19356 ( .A(n16381), .ZN(n16383) );
  NAND2_X1 U19357 ( .A1(n16383), .A2(n16382), .ZN(n16384) );
  OAI211_X1 U19358 ( .C1(n16386), .C2(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A(
        n16385), .B(n16384), .ZN(n16387) );
  INV_X1 U19359 ( .A(n16387), .ZN(n16402) );
  OAI21_X1 U19360 ( .B1(n16387), .B2(P2_STATE2_REG_1__SCAN_IN), .A(
        P2_STATE2_REG_0__SCAN_IN), .ZN(n16393) );
  NAND3_X1 U19361 ( .A1(n16390), .A2(n16389), .A3(n16388), .ZN(n16391) );
  NAND3_X1 U19362 ( .A1(n16393), .A2(n16392), .A3(n16391), .ZN(n19807) );
  OAI21_X1 U19363 ( .B1(n19916), .B2(n19915), .A(n19807), .ZN(n16396) );
  AOI211_X1 U19364 ( .C1(P2_STATE2_REG_0__SCAN_IN), .C2(n16396), .A(n16395), 
        .B(n16394), .ZN(n16401) );
  NOR2_X1 U19365 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n16397), .ZN(n16398) );
  OAI22_X1 U19366 ( .A1(n16399), .A2(n16398), .B1(n19803), .B2(n19807), .ZN(
        n16400) );
  OAI211_X1 U19367 ( .C1(n16402), .C2(n18914), .A(n16401), .B(n16400), .ZN(
        P2_U3176) );
  INV_X1 U19368 ( .A(n16403), .ZN(n16404) );
  OAI221_X1 U19369 ( .B1(n19917), .B2(P2_STATE2_REG_0__SCAN_IN), .C1(n19917), 
        .C2(n19807), .A(n16404), .ZN(P2_U3593) );
  XNOR2_X1 U19370 ( .A(n16417), .B(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16583) );
  INV_X1 U19371 ( .A(n16583), .ZN(n16601) );
  INV_X1 U19372 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n16602) );
  NAND2_X1 U19373 ( .A1(n18231), .A2(P3_REIP_REG_30__SCAN_IN), .ZN(n16405) );
  OAI221_X1 U19374 ( .B1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n16407), .C1(
        n16602), .C2(n16406), .A(n16405), .ZN(n16408) );
  AOI21_X1 U19375 ( .B1(n17767), .B2(n16601), .A(n16408), .ZN(n16413) );
  OAI22_X1 U19376 ( .A1(n16427), .A2(n17914), .B1(n16425), .B2(n17822), .ZN(
        n16411) );
  INV_X1 U19377 ( .A(n18022), .ZN(n18101) );
  NOR2_X1 U19378 ( .A1(n16409), .A2(n17721), .ZN(n17566) );
  AOI22_X1 U19379 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16411), .B1(
        n16410), .B2(n17566), .ZN(n16412) );
  OAI211_X1 U19380 ( .C1(n17808), .C2(n16414), .A(n16413), .B(n16412), .ZN(
        P3_U2800) );
  OAI21_X1 U19381 ( .B1(n18343), .B2(n16415), .A(n16610), .ZN(n16423) );
  INV_X1 U19382 ( .A(n16416), .ZN(n16420) );
  INV_X1 U19383 ( .A(n16417), .ZN(n16418) );
  OAI21_X1 U19384 ( .B1(n16419), .B2(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n16418), .ZN(n16616) );
  AOI21_X1 U19385 ( .B1(n17750), .B2(n16420), .A(n16616), .ZN(n16422) );
  AOI211_X1 U19386 ( .C1(n16424), .C2(n16423), .A(n16422), .B(n16421), .ZN(
        n16433) );
  NOR2_X1 U19387 ( .A1(n16425), .A2(n17822), .ZN(n16431) );
  INV_X1 U19388 ( .A(n16426), .ZN(n16448) );
  NOR2_X1 U19389 ( .A1(n16448), .A2(n17916), .ZN(n16451) );
  OR2_X1 U19390 ( .A1(n17917), .A2(n16448), .ZN(n16428) );
  AOI211_X1 U19391 ( .C1(n16429), .C2(n16428), .A(n16427), .B(n17914), .ZN(
        n16430) );
  AOI221_X1 U19392 ( .B1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n16431), 
        .C1(n16451), .C2(n16431), .A(n16430), .ZN(n16432) );
  OAI211_X1 U19393 ( .C1(n17808), .C2(n16434), .A(n16433), .B(n16432), .ZN(
        P3_U2801) );
  OAI21_X1 U19394 ( .B1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n18140), .A(
        n16435), .ZN(n16441) );
  NAND2_X1 U19395 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n18848), .ZN(
        n16437) );
  NOR4_X1 U19396 ( .A1(n16438), .A2(n16437), .A3(n16436), .A4(n18214), .ZN(
        n16439) );
  AOI211_X1 U19397 ( .C1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .C2(n16441), .A(
        n16440), .B(n16439), .ZN(n16445) );
  AOI22_X1 U19398 ( .A1(n16443), .A2(n18021), .B1(n16442), .B2(n18147), .ZN(
        n16444) );
  OAI211_X1 U19399 ( .C1(n16446), .C2(n18224), .A(n16445), .B(n16444), .ZN(
        P3_U2831) );
  NAND2_X1 U19400 ( .A1(n18231), .A2(P3_REIP_REG_28__SCAN_IN), .ZN(n17548) );
  AOI22_X1 U19401 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17757), .B1(
        n17818), .B2(n17553), .ZN(n17545) );
  AOI21_X1 U19402 ( .B1(n17818), .B2(n17561), .A(n17559), .ZN(n17544) );
  NOR2_X1 U19403 ( .A1(n17545), .A2(n17544), .ZN(n17543) );
  NOR4_X1 U19404 ( .A1(n16447), .A2(n17393), .A3(n17543), .A4(n18687), .ZN(
        n16453) );
  OAI21_X1 U19405 ( .B1(n17917), .B2(n16448), .A(n18681), .ZN(n16449) );
  OAI211_X1 U19406 ( .C1(n16451), .C2(n18083), .A(n16450), .B(n16449), .ZN(
        n16452) );
  OAI211_X1 U19407 ( .C1(n16453), .C2(n16452), .A(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B(n18218), .ZN(n16462) );
  NAND2_X1 U19408 ( .A1(n16454), .A2(n18227), .ZN(n18235) );
  NOR3_X1 U19409 ( .A1(n17543), .A2(n17757), .A3(n18235), .ZN(n16459) );
  INV_X1 U19410 ( .A(n17919), .ZN(n18016) );
  INV_X1 U19411 ( .A(n18692), .ZN(n18712) );
  AOI21_X1 U19412 ( .B1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n18712), .A(
        n18699), .ZN(n18200) );
  INV_X1 U19413 ( .A(n16455), .ZN(n16456) );
  OAI211_X1 U19414 ( .C1(n18016), .C2(n18200), .A(n16457), .B(n16456), .ZN(
        n17930) );
  NAND2_X1 U19415 ( .A1(n18227), .A2(n17930), .ZN(n17997) );
  NOR2_X1 U19416 ( .A1(n17639), .A2(n17997), .ZN(n17982) );
  OAI211_X1 U19417 ( .C1(n16459), .C2(n17982), .A(n16458), .B(n17553), .ZN(
        n16461) );
  NAND3_X1 U19418 ( .A1(n17559), .A2(n18147), .A3(n17545), .ZN(n16460) );
  NAND4_X1 U19419 ( .A1(n17548), .A2(n16462), .A3(n16461), .A4(n16460), .ZN(
        P3_U2834) );
  NOR3_X1 U19420 ( .A1(P3_BE_N_REG_3__SCAN_IN), .A2(P3_W_R_N_REG_SCAN_IN), 
        .A3(P3_BE_N_REG_0__SCAN_IN), .ZN(n16464) );
  NOR4_X1 U19421 ( .A1(P3_BE_N_REG_1__SCAN_IN), .A2(P3_BE_N_REG_2__SCAN_IN), 
        .A3(P3_D_C_N_REG_SCAN_IN), .A4(P3_ADS_N_REG_SCAN_IN), .ZN(n16463) );
  NAND4_X1 U19422 ( .A1(P3_M_IO_N_REG_SCAN_IN), .A2(n16464), .A3(n16463), .A4(
        U215), .ZN(U213) );
  INV_X2 U19423 ( .A(U212), .ZN(n16512) );
  INV_X2 U19424 ( .A(U214), .ZN(n16513) );
  NOR2_X1 U19425 ( .A1(n16513), .A2(n16465), .ZN(n16509) );
  AOI222_X1 U19426 ( .A1(n16512), .A2(P2_DATAO_REG_31__SCAN_IN), .B1(n16509), 
        .B2(BUF1_REG_31__SCAN_IN), .C1(n16513), .C2(P1_DATAO_REG_31__SCAN_IN), 
        .ZN(n16466) );
  INV_X1 U19427 ( .A(n16466), .ZN(U216) );
  INV_X1 U19428 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n19173) );
  INV_X1 U19429 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n16550) );
  OAI222_X1 U19430 ( .A1(U212), .A2(n19173), .B1(n16515), .B2(n16467), .C1(
        U214), .C2(n16550), .ZN(U217) );
  AOI222_X1 U19431 ( .A1(n16512), .A2(P2_DATAO_REG_29__SCAN_IN), .B1(n16509), 
        .B2(BUF1_REG_29__SCAN_IN), .C1(n16513), .C2(P1_DATAO_REG_29__SCAN_IN), 
        .ZN(n16468) );
  INV_X1 U19432 ( .A(n16468), .ZN(U218) );
  INV_X1 U19433 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n16470) );
  AOI22_X1 U19434 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(n16513), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(n16512), .ZN(n16469) );
  OAI21_X1 U19435 ( .B1(n16470), .B2(n16515), .A(n16469), .ZN(U219) );
  AOI222_X1 U19436 ( .A1(n16512), .A2(P2_DATAO_REG_27__SCAN_IN), .B1(n16509), 
        .B2(BUF1_REG_27__SCAN_IN), .C1(n16513), .C2(P1_DATAO_REG_27__SCAN_IN), 
        .ZN(n16471) );
  INV_X1 U19437 ( .A(n16471), .ZN(U220) );
  INV_X1 U19438 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n16473) );
  AOI22_X1 U19439 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(n16513), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(n16512), .ZN(n16472) );
  OAI21_X1 U19440 ( .B1(n16473), .B2(n16515), .A(n16472), .ZN(U221) );
  INV_X1 U19441 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n16475) );
  AOI22_X1 U19442 ( .A1(P1_DATAO_REG_25__SCAN_IN), .A2(n16513), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(n16512), .ZN(n16474) );
  OAI21_X1 U19443 ( .B1(n16475), .B2(n16515), .A(n16474), .ZN(U222) );
  INV_X1 U19444 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n16477) );
  AOI22_X1 U19445 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n16513), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(n16512), .ZN(n16476) );
  OAI21_X1 U19446 ( .B1(n16477), .B2(n16515), .A(n16476), .ZN(U223) );
  INV_X1 U19447 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n16479) );
  AOI22_X1 U19448 ( .A1(P1_DATAO_REG_23__SCAN_IN), .A2(n16513), .B1(
        P2_DATAO_REG_23__SCAN_IN), .B2(n16512), .ZN(n16478) );
  OAI21_X1 U19449 ( .B1(n16479), .B2(n16515), .A(n16478), .ZN(U224) );
  AOI22_X1 U19450 ( .A1(P1_DATAO_REG_22__SCAN_IN), .A2(n16513), .B1(
        P2_DATAO_REG_22__SCAN_IN), .B2(n16512), .ZN(n16480) );
  OAI21_X1 U19451 ( .B1(n14776), .B2(n16515), .A(n16480), .ZN(U225) );
  INV_X1 U19452 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n16482) );
  AOI22_X1 U19453 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(n16513), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(n16512), .ZN(n16481) );
  OAI21_X1 U19454 ( .B1(n16482), .B2(n16515), .A(n16481), .ZN(U226) );
  AOI22_X1 U19455 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n16513), .B1(
        P2_DATAO_REG_20__SCAN_IN), .B2(n16512), .ZN(n16483) );
  OAI21_X1 U19456 ( .B1(n16484), .B2(n16515), .A(n16483), .ZN(U227) );
  INV_X1 U19457 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n16486) );
  AOI22_X1 U19458 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(n16513), .B1(
        P2_DATAO_REG_19__SCAN_IN), .B2(n16512), .ZN(n16485) );
  OAI21_X1 U19459 ( .B1(n16486), .B2(n16515), .A(n16485), .ZN(U228) );
  AOI22_X1 U19460 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(n16513), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n16512), .ZN(n16487) );
  OAI21_X1 U19461 ( .B1(n14790), .B2(n16515), .A(n16487), .ZN(U229) );
  INV_X1 U19462 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n16489) );
  AOI22_X1 U19463 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(n16513), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n16512), .ZN(n16488) );
  OAI21_X1 U19464 ( .B1(n16489), .B2(n16515), .A(n16488), .ZN(U230) );
  AOI22_X1 U19465 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n16513), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n16512), .ZN(n16490) );
  OAI21_X1 U19466 ( .B1(n14801), .B2(n16515), .A(n16490), .ZN(U231) );
  AOI22_X1 U19467 ( .A1(P1_DATAO_REG_15__SCAN_IN), .A2(n16513), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n16512), .ZN(n16491) );
  OAI21_X1 U19468 ( .B1(n13588), .B2(n16515), .A(n16491), .ZN(U232) );
  AOI22_X1 U19469 ( .A1(P1_DATAO_REG_14__SCAN_IN), .A2(n16513), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n16512), .ZN(n16492) );
  OAI21_X1 U19470 ( .B1(n14371), .B2(n16515), .A(n16492), .ZN(U233) );
  AOI22_X1 U19471 ( .A1(P1_DATAO_REG_13__SCAN_IN), .A2(n16513), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n16512), .ZN(n16493) );
  OAI21_X1 U19472 ( .B1(n13503), .B2(n16515), .A(n16493), .ZN(U234) );
  AOI22_X1 U19473 ( .A1(P1_DATAO_REG_12__SCAN_IN), .A2(n16513), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n16512), .ZN(n16494) );
  OAI21_X1 U19474 ( .B1(n16495), .B2(n16515), .A(n16494), .ZN(U235) );
  AOI22_X1 U19475 ( .A1(P1_DATAO_REG_11__SCAN_IN), .A2(n16513), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n16512), .ZN(n16496) );
  OAI21_X1 U19476 ( .B1(n13457), .B2(n16515), .A(n16496), .ZN(U236) );
  AOI22_X1 U19477 ( .A1(P1_DATAO_REG_10__SCAN_IN), .A2(n16513), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n16512), .ZN(n16497) );
  OAI21_X1 U19478 ( .B1(n21071), .B2(n16515), .A(n16497), .ZN(U237) );
  AOI22_X1 U19479 ( .A1(P1_DATAO_REG_9__SCAN_IN), .A2(n16513), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n16512), .ZN(n16498) );
  OAI21_X1 U19480 ( .B1(n13440), .B2(n16515), .A(n16498), .ZN(U238) );
  AOI22_X1 U19481 ( .A1(P1_DATAO_REG_8__SCAN_IN), .A2(n16513), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n16512), .ZN(n16499) );
  OAI21_X1 U19482 ( .B1(n13450), .B2(n16515), .A(n16499), .ZN(U239) );
  INV_X1 U19483 ( .A(BUF1_REG_7__SCAN_IN), .ZN(n21152) );
  AOI22_X1 U19484 ( .A1(P1_DATAO_REG_7__SCAN_IN), .A2(n16513), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n16512), .ZN(n16500) );
  OAI21_X1 U19485 ( .B1(n21152), .B2(n16515), .A(n16500), .ZN(U240) );
  INV_X1 U19486 ( .A(BUF1_REG_6__SCAN_IN), .ZN(n16502) );
  AOI22_X1 U19487 ( .A1(P1_DATAO_REG_6__SCAN_IN), .A2(n16513), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n16512), .ZN(n16501) );
  OAI21_X1 U19488 ( .B1(n16502), .B2(n16515), .A(n16501), .ZN(U241) );
  INV_X1 U19489 ( .A(BUF1_REG_5__SCAN_IN), .ZN(n16504) );
  AOI22_X1 U19490 ( .A1(P1_DATAO_REG_5__SCAN_IN), .A2(n16513), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n16512), .ZN(n16503) );
  OAI21_X1 U19491 ( .B1(n16504), .B2(n16515), .A(n16503), .ZN(U242) );
  AOI22_X1 U19492 ( .A1(P1_DATAO_REG_4__SCAN_IN), .A2(n16513), .B1(
        P2_DATAO_REG_4__SCAN_IN), .B2(n16512), .ZN(n16505) );
  OAI21_X1 U19493 ( .B1(n16506), .B2(n16515), .A(n16505), .ZN(U243) );
  INV_X1 U19494 ( .A(BUF1_REG_3__SCAN_IN), .ZN(n16508) );
  AOI22_X1 U19495 ( .A1(P1_DATAO_REG_3__SCAN_IN), .A2(n16513), .B1(
        P2_DATAO_REG_3__SCAN_IN), .B2(n16512), .ZN(n16507) );
  OAI21_X1 U19496 ( .B1(n16508), .B2(n16515), .A(n16507), .ZN(U244) );
  AOI222_X1 U19497 ( .A1(n16512), .A2(P2_DATAO_REG_2__SCAN_IN), .B1(n16509), 
        .B2(BUF1_REG_2__SCAN_IN), .C1(n16513), .C2(P1_DATAO_REG_2__SCAN_IN), 
        .ZN(n16510) );
  INV_X1 U19498 ( .A(n16510), .ZN(U245) );
  INV_X1 U19499 ( .A(BUF1_REG_1__SCAN_IN), .ZN(n21010) );
  AOI22_X1 U19500 ( .A1(P1_DATAO_REG_1__SCAN_IN), .A2(n16513), .B1(
        P2_DATAO_REG_1__SCAN_IN), .B2(n16512), .ZN(n16511) );
  OAI21_X1 U19501 ( .B1(n21010), .B2(n16515), .A(n16511), .ZN(U246) );
  AOI22_X1 U19502 ( .A1(P1_DATAO_REG_0__SCAN_IN), .A2(n16513), .B1(
        P2_DATAO_REG_0__SCAN_IN), .B2(n16512), .ZN(n16514) );
  OAI21_X1 U19503 ( .B1(n16516), .B2(n16515), .A(n16514), .ZN(U247) );
  INV_X1 U19504 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n16517) );
  AOI22_X1 U19505 ( .A1(n16547), .A2(n16517), .B1(n21157), .B2(U215), .ZN(U251) );
  OAI22_X1 U19506 ( .A1(U215), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n16547), .ZN(n16518) );
  INV_X1 U19507 ( .A(n16518), .ZN(U252) );
  OAI22_X1 U19508 ( .A1(U215), .A2(P2_DATAO_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n16547), .ZN(n16519) );
  INV_X1 U19509 ( .A(n16519), .ZN(U253) );
  INV_X1 U19510 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n16520) );
  INV_X1 U19511 ( .A(BUF2_REG_3__SCAN_IN), .ZN(n18257) );
  AOI22_X1 U19512 ( .A1(n16547), .A2(n16520), .B1(n18257), .B2(U215), .ZN(U254) );
  INV_X1 U19513 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n16521) );
  AOI22_X1 U19514 ( .A1(n16547), .A2(n16521), .B1(n18261), .B2(U215), .ZN(U255) );
  INV_X1 U19515 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n16522) );
  INV_X1 U19516 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n18265) );
  AOI22_X1 U19517 ( .A1(n16536), .A2(n16522), .B1(n18265), .B2(U215), .ZN(U256) );
  INV_X1 U19518 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n16523) );
  INV_X1 U19519 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n18270) );
  AOI22_X1 U19520 ( .A1(n16547), .A2(n16523), .B1(n18270), .B2(U215), .ZN(U257) );
  INV_X1 U19521 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n16524) );
  INV_X1 U19522 ( .A(BUF2_REG_7__SCAN_IN), .ZN(n18274) );
  AOI22_X1 U19523 ( .A1(n16547), .A2(n16524), .B1(n18274), .B2(U215), .ZN(U258) );
  INV_X1 U19524 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n16525) );
  INV_X1 U19525 ( .A(BUF2_REG_8__SCAN_IN), .ZN(n21054) );
  AOI22_X1 U19526 ( .A1(n16536), .A2(n16525), .B1(n21054), .B2(U215), .ZN(U259) );
  INV_X1 U19527 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n16526) );
  INV_X1 U19528 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n17522) );
  AOI22_X1 U19529 ( .A1(n16547), .A2(n16526), .B1(n17522), .B2(U215), .ZN(U260) );
  INV_X1 U19530 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n16527) );
  INV_X1 U19531 ( .A(BUF2_REG_10__SCAN_IN), .ZN(n17524) );
  AOI22_X1 U19532 ( .A1(n16536), .A2(n16527), .B1(n17524), .B2(U215), .ZN(U261) );
  INV_X1 U19533 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n16528) );
  INV_X1 U19534 ( .A(BUF2_REG_11__SCAN_IN), .ZN(n17526) );
  AOI22_X1 U19535 ( .A1(n16536), .A2(n16528), .B1(n17526), .B2(U215), .ZN(U262) );
  INV_X1 U19536 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n16529) );
  INV_X1 U19537 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n17528) );
  AOI22_X1 U19538 ( .A1(n16547), .A2(n16529), .B1(n17528), .B2(U215), .ZN(U263) );
  INV_X1 U19539 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n16530) );
  INV_X1 U19540 ( .A(BUF2_REG_13__SCAN_IN), .ZN(n17533) );
  AOI22_X1 U19541 ( .A1(n16547), .A2(n16530), .B1(n17533), .B2(U215), .ZN(U264) );
  OAI22_X1 U19542 ( .A1(U215), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n16536), .ZN(n16531) );
  INV_X1 U19543 ( .A(n16531), .ZN(U265) );
  OAI22_X1 U19544 ( .A1(U215), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n16536), .ZN(n16532) );
  INV_X1 U19545 ( .A(n16532), .ZN(U266) );
  OAI22_X1 U19546 ( .A1(U215), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n16536), .ZN(n16533) );
  INV_X1 U19547 ( .A(n16533), .ZN(U267) );
  OAI22_X1 U19548 ( .A1(U215), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n16536), .ZN(n16534) );
  INV_X1 U19549 ( .A(n16534), .ZN(U268) );
  OAI22_X1 U19550 ( .A1(U215), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n16536), .ZN(n16535) );
  INV_X1 U19551 ( .A(n16535), .ZN(U269) );
  OAI22_X1 U19552 ( .A1(U215), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n16536), .ZN(n16537) );
  INV_X1 U19553 ( .A(n16537), .ZN(U270) );
  INV_X1 U19554 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n16538) );
  INV_X1 U19555 ( .A(BUF2_REG_20__SCAN_IN), .ZN(n17329) );
  AOI22_X1 U19556 ( .A1(n16547), .A2(n16538), .B1(n17329), .B2(U215), .ZN(U271) );
  OAI22_X1 U19557 ( .A1(U215), .A2(P2_DATAO_REG_21__SCAN_IN), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n16547), .ZN(n16539) );
  INV_X1 U19558 ( .A(n16539), .ZN(U272) );
  INV_X1 U19559 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n16540) );
  INV_X1 U19560 ( .A(BUF2_REG_22__SCAN_IN), .ZN(n17316) );
  AOI22_X1 U19561 ( .A1(n16547), .A2(n16540), .B1(n17316), .B2(U215), .ZN(U273) );
  OAI22_X1 U19562 ( .A1(U215), .A2(P2_DATAO_REG_23__SCAN_IN), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n16547), .ZN(n16541) );
  INV_X1 U19563 ( .A(n16541), .ZN(U274) );
  OAI22_X1 U19564 ( .A1(U215), .A2(P2_DATAO_REG_24__SCAN_IN), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n16547), .ZN(n16542) );
  INV_X1 U19565 ( .A(n16542), .ZN(U275) );
  OAI22_X1 U19566 ( .A1(U215), .A2(P2_DATAO_REG_25__SCAN_IN), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n16547), .ZN(n16543) );
  INV_X1 U19567 ( .A(n16543), .ZN(U276) );
  OAI22_X1 U19568 ( .A1(U215), .A2(P2_DATAO_REG_26__SCAN_IN), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n16547), .ZN(n16544) );
  INV_X1 U19569 ( .A(n16544), .ZN(U277) );
  INV_X1 U19570 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n20918) );
  INV_X1 U19571 ( .A(BUF2_REG_27__SCAN_IN), .ZN(n17294) );
  AOI22_X1 U19572 ( .A1(n16547), .A2(n20918), .B1(n17294), .B2(U215), .ZN(U278) );
  OAI22_X1 U19573 ( .A1(U215), .A2(P2_DATAO_REG_28__SCAN_IN), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n16547), .ZN(n16545) );
  INV_X1 U19574 ( .A(n16545), .ZN(U279) );
  INV_X1 U19575 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n21041) );
  INV_X1 U19576 ( .A(BUF2_REG_29__SCAN_IN), .ZN(n18266) );
  AOI22_X1 U19577 ( .A1(n16547), .A2(n21041), .B1(n18266), .B2(U215), .ZN(U280) );
  INV_X1 U19578 ( .A(BUF2_REG_30__SCAN_IN), .ZN(n16546) );
  AOI22_X1 U19579 ( .A1(n16547), .A2(n19173), .B1(n16546), .B2(U215), .ZN(U281) );
  OAI22_X1 U19580 ( .A1(U215), .A2(P2_DATAO_REG_31__SCAN_IN), .B1(
        BUF2_REG_31__SCAN_IN), .B2(n16547), .ZN(n16548) );
  INV_X1 U19581 ( .A(n16548), .ZN(U282) );
  INV_X1 U19582 ( .A(P3_DATAO_REG_30__SCAN_IN), .ZN(n16549) );
  OAI222_X1 U19583 ( .A1(P1_DATAO_REG_31__SCAN_IN), .A2(n16550), .B1(
        P2_DATAO_REG_31__SCAN_IN), .B2(n19173), .C1(P3_DATAO_REG_31__SCAN_IN), 
        .C2(n16549), .ZN(n16551) );
  INV_X1 U19584 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n18785) );
  INV_X1 U19585 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n19844) );
  AOI22_X1 U19586 ( .A1(n9840), .A2(n18785), .B1(n19844), .B2(n16552), .ZN(
        U347) );
  INV_X1 U19587 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n18783) );
  INV_X1 U19588 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n19843) );
  AOI22_X1 U19589 ( .A1(n9840), .A2(n18783), .B1(n19843), .B2(n16552), .ZN(
        U348) );
  INV_X1 U19590 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n18780) );
  INV_X1 U19591 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n19841) );
  AOI22_X1 U19592 ( .A1(n9840), .A2(n18780), .B1(n19841), .B2(n16552), .ZN(
        U349) );
  INV_X1 U19593 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n18779) );
  INV_X1 U19594 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n19840) );
  AOI22_X1 U19595 ( .A1(n9840), .A2(n18779), .B1(n19840), .B2(n16552), .ZN(
        U350) );
  INV_X1 U19596 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n21077) );
  INV_X1 U19597 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n19839) );
  AOI22_X1 U19598 ( .A1(n9840), .A2(n21077), .B1(n19839), .B2(n16552), .ZN(
        U351) );
  INV_X1 U19599 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n18776) );
  INV_X1 U19600 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n19837) );
  AOI22_X1 U19601 ( .A1(n9840), .A2(n18776), .B1(n19837), .B2(n16552), .ZN(
        U352) );
  INV_X1 U19602 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n18775) );
  INV_X1 U19603 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n19835) );
  AOI22_X1 U19604 ( .A1(n9840), .A2(n18775), .B1(n19835), .B2(n16552), .ZN(
        U353) );
  INV_X1 U19605 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n21127) );
  AOI22_X1 U19606 ( .A1(n9840), .A2(n21127), .B1(n19834), .B2(n16552), .ZN(
        U354) );
  INV_X1 U19607 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n18824) );
  INV_X1 U19608 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n21093) );
  AOI22_X1 U19609 ( .A1(n9840), .A2(n18824), .B1(n21093), .B2(n16551), .ZN(
        U355) );
  INV_X1 U19610 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n18820) );
  INV_X1 U19611 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n19872) );
  AOI22_X1 U19612 ( .A1(n9840), .A2(n18820), .B1(n19872), .B2(n16552), .ZN(
        U356) );
  INV_X1 U19613 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n18817) );
  INV_X1 U19614 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n19870) );
  AOI22_X1 U19615 ( .A1(n9840), .A2(n18817), .B1(n19870), .B2(n16552), .ZN(
        U357) );
  INV_X1 U19616 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n18816) );
  INV_X1 U19617 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n19868) );
  AOI22_X1 U19618 ( .A1(n9840), .A2(n18816), .B1(n19868), .B2(n16551), .ZN(
        U358) );
  INV_X1 U19619 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n18814) );
  INV_X1 U19620 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n19867) );
  AOI22_X1 U19621 ( .A1(n9840), .A2(n18814), .B1(n19867), .B2(n16551), .ZN(
        U359) );
  INV_X1 U19622 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n18812) );
  INV_X1 U19623 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n19865) );
  AOI22_X1 U19624 ( .A1(n9840), .A2(n18812), .B1(n19865), .B2(n16551), .ZN(
        U360) );
  INV_X1 U19625 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n18810) );
  INV_X1 U19626 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n19863) );
  AOI22_X1 U19627 ( .A1(n9840), .A2(n18810), .B1(n19863), .B2(n16551), .ZN(
        U361) );
  INV_X1 U19628 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n21080) );
  INV_X1 U19629 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n19861) );
  AOI22_X1 U19630 ( .A1(n9840), .A2(n21080), .B1(n19861), .B2(n16552), .ZN(
        U362) );
  INV_X1 U19631 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n18807) );
  INV_X1 U19632 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n19859) );
  AOI22_X1 U19633 ( .A1(n9840), .A2(n18807), .B1(n19859), .B2(n16552), .ZN(
        U363) );
  INV_X1 U19634 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n18805) );
  INV_X1 U19635 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n19858) );
  AOI22_X1 U19636 ( .A1(n9840), .A2(n18805), .B1(n19858), .B2(n16552), .ZN(
        U364) );
  INV_X1 U19637 ( .A(P3_ADDRESS_REG_1__SCAN_IN), .ZN(n18772) );
  INV_X1 U19638 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n19833) );
  AOI22_X1 U19639 ( .A1(n9840), .A2(n18772), .B1(n19833), .B2(n16552), .ZN(
        U365) );
  INV_X1 U19640 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n18802) );
  INV_X1 U19641 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n19857) );
  AOI22_X1 U19642 ( .A1(n9840), .A2(n18802), .B1(n19857), .B2(n16552), .ZN(
        U366) );
  INV_X1 U19643 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n18801) );
  INV_X1 U19644 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n19855) );
  AOI22_X1 U19645 ( .A1(n9840), .A2(n18801), .B1(n19855), .B2(n16552), .ZN(
        U367) );
  INV_X1 U19646 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n18799) );
  INV_X1 U19647 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n19853) );
  AOI22_X1 U19648 ( .A1(n9840), .A2(n18799), .B1(n19853), .B2(n16552), .ZN(
        U368) );
  INV_X1 U19649 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n18796) );
  INV_X1 U19650 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n19852) );
  AOI22_X1 U19651 ( .A1(n9840), .A2(n18796), .B1(n19852), .B2(n16552), .ZN(
        U369) );
  INV_X1 U19652 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n18795) );
  INV_X1 U19653 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n19851) );
  AOI22_X1 U19654 ( .A1(n9840), .A2(n18795), .B1(n19851), .B2(n16552), .ZN(
        U370) );
  INV_X1 U19655 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n18794) );
  INV_X1 U19656 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n19849) );
  AOI22_X1 U19657 ( .A1(n9840), .A2(n18794), .B1(n19849), .B2(n16552), .ZN(
        U371) );
  INV_X1 U19658 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n18792) );
  INV_X1 U19659 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n19848) );
  AOI22_X1 U19660 ( .A1(n9840), .A2(n18792), .B1(n19848), .B2(n16551), .ZN(
        U372) );
  INV_X1 U19661 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n18791) );
  INV_X1 U19662 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n19847) );
  AOI22_X1 U19663 ( .A1(n9840), .A2(n18791), .B1(n19847), .B2(n16552), .ZN(
        U373) );
  INV_X1 U19664 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n18788) );
  INV_X1 U19665 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n19846) );
  AOI22_X1 U19666 ( .A1(n9840), .A2(n18788), .B1(n19846), .B2(n16551), .ZN(
        U374) );
  INV_X1 U19667 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n18787) );
  INV_X1 U19668 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n19845) );
  AOI22_X1 U19669 ( .A1(n9840), .A2(n18787), .B1(n19845), .B2(n16551), .ZN(
        U375) );
  INV_X1 U19670 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n18770) );
  INV_X1 U19671 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n19832) );
  AOI22_X1 U19672 ( .A1(n9840), .A2(n18770), .B1(n19832), .B2(n16552), .ZN(
        U376) );
  INV_X1 U19673 ( .A(P3_ADS_N_REG_SCAN_IN), .ZN(n16553) );
  INV_X1 U19674 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n18769) );
  NAND2_X1 U19675 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(n18769), .ZN(n18757) );
  AOI22_X1 U19676 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n18757), .B1(
        P3_STATE_REG_1__SCAN_IN), .B2(n18767), .ZN(n18835) );
  OAI21_X1 U19677 ( .B1(n18767), .B2(n16553), .A(n18832), .ZN(P3_U2633) );
  INV_X1 U19678 ( .A(n16559), .ZN(n16554) );
  OAI21_X1 U19679 ( .B1(n16554), .B2(n17491), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n16555) );
  OAI21_X1 U19680 ( .B1(n16556), .B2(n18747), .A(n16555), .ZN(P3_U2634) );
  AOI21_X1 U19681 ( .B1(n18767), .B2(n18769), .A(P3_D_C_N_REG_SCAN_IN), .ZN(
        n16557) );
  AOI22_X1 U19682 ( .A1(n18898), .A2(P3_CODEFETCH_REG_SCAN_IN), .B1(n16557), 
        .B2(n18899), .ZN(P3_U2635) );
  NOR2_X1 U19683 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(P3_STATE_REG_2__SCAN_IN), 
        .ZN(n18754) );
  OAI21_X1 U19684 ( .B1(n18754), .B2(BS16), .A(n18835), .ZN(n18833) );
  OAI21_X1 U19685 ( .B1(n18835), .B2(n18887), .A(n18833), .ZN(P3_U2636) );
  AND3_X1 U19686 ( .A1(n18685), .A2(n16559), .A3(n16558), .ZN(n18688) );
  NOR2_X1 U19687 ( .A1(n18688), .A2(n18743), .ZN(n18878) );
  OAI21_X1 U19688 ( .B1(n18878), .B2(n21087), .A(n16560), .ZN(P3_U2637) );
  NOR4_X1 U19689 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_21__SCAN_IN), .A3(P3_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_23__SCAN_IN), .ZN(n16564) );
  NOR4_X1 U19690 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_17__SCAN_IN), .A3(P3_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_19__SCAN_IN), .ZN(n16563) );
  NOR4_X1 U19691 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_29__SCAN_IN), .A3(P3_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_31__SCAN_IN), .ZN(n16562) );
  NOR4_X1 U19692 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_25__SCAN_IN), .A3(P3_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_27__SCAN_IN), .ZN(n16561) );
  NAND4_X1 U19693 ( .A1(n16564), .A2(n16563), .A3(n16562), .A4(n16561), .ZN(
        n16570) );
  NOR4_X1 U19694 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_4__SCAN_IN), .A3(P3_DATAWIDTH_REG_5__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_6__SCAN_IN), .ZN(n16568) );
  AOI211_X1 U19695 ( .C1(P3_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_11__SCAN_IN), .B(
        P3_DATAWIDTH_REG_2__SCAN_IN), .ZN(n16567) );
  NOR4_X1 U19696 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_13__SCAN_IN), .A3(P3_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_15__SCAN_IN), .ZN(n16566) );
  NOR4_X1 U19697 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_8__SCAN_IN), .A3(P3_DATAWIDTH_REG_9__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_10__SCAN_IN), .ZN(n16565) );
  NAND4_X1 U19698 ( .A1(n16568), .A2(n16567), .A3(n16566), .A4(n16565), .ZN(
        n16569) );
  NOR2_X1 U19699 ( .A1(n16570), .A2(n16569), .ZN(n20816) );
  INV_X1 U19700 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n20815) );
  INV_X1 U19701 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n18834) );
  NOR3_X1 U19702 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A3(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n20818) );
  AOI21_X1 U19703 ( .B1(n20815), .B2(n18834), .A(n20818), .ZN(n16571) );
  INV_X1 U19704 ( .A(P3_BYTEENABLE_REG_3__SCAN_IN), .ZN(n18827) );
  INV_X1 U19705 ( .A(n20816), .ZN(n18872) );
  AOI22_X1 U19706 ( .A1(n20816), .A2(n16571), .B1(n18827), .B2(n18872), .ZN(
        P3_U2639) );
  INV_X1 U19707 ( .A(n16572), .ZN(n16575) );
  INV_X1 U19708 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n17563) );
  NOR2_X1 U19709 ( .A1(n16575), .A2(n17563), .ZN(n16574) );
  OAI21_X1 U19710 ( .B1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n16574), .A(
        n16573), .ZN(n17550) );
  AOI21_X1 U19711 ( .B1(n16575), .B2(n17563), .A(n16574), .ZN(n17558) );
  INV_X1 U19712 ( .A(n17558), .ZN(n16635) );
  INV_X1 U19713 ( .A(n17542), .ZN(n16576) );
  OAI21_X1 U19714 ( .B1(n16576), .B2(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n16575), .ZN(n17576) );
  INV_X1 U19715 ( .A(n16579), .ZN(n16578) );
  INV_X1 U19716 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n17603) );
  NOR2_X1 U19717 ( .A1(n16578), .A2(n17603), .ZN(n16577) );
  OAI21_X1 U19718 ( .B1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n16577), .A(
        n17542), .ZN(n17587) );
  AOI22_X1 U19719 ( .A1(n16579), .A2(n17603), .B1(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n16578), .ZN(n17600) );
  AOI21_X1 U19720 ( .B1(n17586), .B2(n17618), .A(n16579), .ZN(n17616) );
  INV_X1 U19721 ( .A(n17616), .ZN(n16678) );
  OAI21_X1 U19722 ( .B1(n16580), .B2(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n17586), .ZN(n17645) );
  OAI21_X1 U19723 ( .B1(n16582), .B2(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A(
        n16581), .ZN(n17646) );
  AOI21_X1 U19724 ( .B1(n17629), .B2(n17663), .A(n16582), .ZN(n17665) );
  INV_X1 U19725 ( .A(n17665), .ZN(n16713) );
  INV_X1 U19726 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n16888) );
  NAND2_X1 U19727 ( .A1(n16751), .A2(n16888), .ZN(n16753) );
  OAI21_X1 U19728 ( .B1(n17629), .B2(n16753), .A(n16789), .ZN(n16712) );
  NAND2_X1 U19729 ( .A1(n16713), .A2(n16712), .ZN(n16711) );
  NAND2_X1 U19730 ( .A1(n16789), .A2(n16711), .ZN(n16701) );
  NAND2_X1 U19731 ( .A1(n17646), .A2(n16701), .ZN(n16700) );
  NAND2_X1 U19732 ( .A1(n16789), .A2(n16700), .ZN(n16694) );
  NAND2_X1 U19733 ( .A1(n17645), .A2(n16694), .ZN(n16693) );
  NAND2_X1 U19734 ( .A1(n16789), .A2(n16693), .ZN(n16677) );
  NAND2_X1 U19735 ( .A1(n16678), .A2(n16677), .ZN(n16676) );
  NAND2_X1 U19736 ( .A1(n16789), .A2(n16676), .ZN(n16666) );
  NAND2_X1 U19737 ( .A1(n17600), .A2(n16666), .ZN(n16665) );
  NAND2_X1 U19738 ( .A1(n16789), .A2(n16665), .ZN(n16653) );
  NAND2_X1 U19739 ( .A1(n17587), .A2(n16653), .ZN(n16652) );
  NAND2_X1 U19740 ( .A1(n16789), .A2(n16652), .ZN(n16646) );
  NAND2_X1 U19741 ( .A1(n17576), .A2(n16646), .ZN(n16645) );
  NAND2_X1 U19742 ( .A1(n16789), .A2(n16645), .ZN(n16634) );
  NAND2_X1 U19743 ( .A1(n16635), .A2(n16634), .ZN(n16633) );
  NAND2_X1 U19744 ( .A1(n16789), .A2(n16633), .ZN(n16624) );
  NAND2_X1 U19745 ( .A1(n17550), .A2(n16624), .ZN(n16623) );
  NAND2_X1 U19746 ( .A1(n16789), .A2(n16623), .ZN(n16615) );
  NAND2_X1 U19747 ( .A1(n16616), .A2(n16615), .ZN(n16614) );
  NAND2_X1 U19748 ( .A1(n16789), .A2(n16614), .ZN(n16600) );
  NAND2_X1 U19749 ( .A1(n16583), .A2(n16600), .ZN(n16598) );
  NAND3_X1 U19750 ( .A1(n18891), .A2(n18901), .A3(n18887), .ZN(n18752) );
  NOR2_X1 U19751 ( .A1(n18236), .A2(n18752), .ZN(n16914) );
  INV_X1 U19752 ( .A(n16914), .ZN(n18750) );
  NAND2_X1 U19753 ( .A1(n16789), .A2(n16882), .ZN(n16826) );
  NAND2_X1 U19754 ( .A1(P3_EBX_REG_31__SCAN_IN), .A2(n16589), .ZN(n16586) );
  AOI211_X4 U19755 ( .C1(n18887), .C2(n18880), .A(n16587), .B(n16586), .ZN(
        n16936) );
  NOR3_X1 U19756 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .ZN(n16934) );
  NAND2_X1 U19757 ( .A1(n16934), .A2(n17252), .ZN(n16921) );
  NOR2_X1 U19758 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n16921), .ZN(n16904) );
  NAND2_X1 U19759 ( .A1(n16904), .A2(n17230), .ZN(n16894) );
  INV_X1 U19760 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n17237) );
  NAND2_X1 U19761 ( .A1(n16875), .A2(n17237), .ZN(n16867) );
  INV_X1 U19762 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n16842) );
  NAND2_X1 U19763 ( .A1(n16840), .A2(n16842), .ZN(n16824) );
  INV_X1 U19764 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n16821) );
  NAND2_X1 U19765 ( .A1(n16823), .A2(n16821), .ZN(n16813) );
  NAND2_X1 U19766 ( .A1(n16799), .A2(n16792), .ZN(n16790) );
  INV_X1 U19767 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n16768) );
  NAND2_X1 U19768 ( .A1(n16775), .A2(n16768), .ZN(n16766) );
  INV_X1 U19769 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n16746) );
  NAND2_X1 U19770 ( .A1(n16754), .A2(n16746), .ZN(n16745) );
  INV_X1 U19771 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n16721) );
  NAND2_X1 U19772 ( .A1(n16728), .A2(n16721), .ZN(n16719) );
  INV_X1 U19773 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n17026) );
  NAND2_X1 U19774 ( .A1(n16707), .A2(n17026), .ZN(n16702) );
  INV_X1 U19775 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n16680) );
  NAND2_X1 U19776 ( .A1(n16688), .A2(n16680), .ZN(n16679) );
  NAND2_X1 U19777 ( .A1(n16660), .A2(n16651), .ZN(n16650) );
  INV_X1 U19778 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n17005) );
  NAND2_X1 U19779 ( .A1(n16640), .A2(n17005), .ZN(n16632) );
  NOR2_X1 U19780 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n16632), .ZN(n16621) );
  INV_X1 U19781 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n16992) );
  NAND2_X1 U19782 ( .A1(n16621), .A2(n16992), .ZN(n16599) );
  NOR2_X1 U19783 ( .A1(n16954), .A2(n16599), .ZN(n16607) );
  INV_X1 U19784 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n16592) );
  INV_X1 U19785 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n18825) );
  AOI211_X1 U19786 ( .C1(n18885), .C2(n18886), .A(n18889), .B(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n16588) );
  INV_X1 U19787 ( .A(n16588), .ZN(n18736) );
  INV_X1 U19788 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n18813) );
  INV_X1 U19789 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n18809) );
  INV_X1 U19790 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n18786) );
  INV_X1 U19791 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n18774) );
  NAND3_X1 U19792 ( .A1(P3_REIP_REG_3__SCAN_IN), .A2(P3_REIP_REG_1__SCAN_IN), 
        .A3(P3_REIP_REG_2__SCAN_IN), .ZN(n16903) );
  NOR2_X1 U19793 ( .A1(n18774), .A2(n16903), .ZN(n16886) );
  NAND2_X1 U19794 ( .A1(P3_REIP_REG_5__SCAN_IN), .A2(n16886), .ZN(n16868) );
  NAND2_X1 U19795 ( .A1(P3_REIP_REG_6__SCAN_IN), .A2(P3_REIP_REG_7__SCAN_IN), 
        .ZN(n16869) );
  NOR2_X1 U19796 ( .A1(n16868), .A2(n16869), .ZN(n16853) );
  NAND2_X1 U19797 ( .A1(P3_REIP_REG_8__SCAN_IN), .A2(n16853), .ZN(n16809) );
  NAND2_X1 U19798 ( .A1(P3_REIP_REG_10__SCAN_IN), .A2(P3_REIP_REG_9__SCAN_IN), 
        .ZN(n16822) );
  NOR3_X1 U19799 ( .A1(n18786), .A2(n16809), .A3(n16822), .ZN(n16802) );
  NAND2_X1 U19800 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n16802), .ZN(n16671) );
  NAND2_X1 U19801 ( .A1(P3_REIP_REG_14__SCAN_IN), .A2(P3_REIP_REG_13__SCAN_IN), 
        .ZN(n16670) );
  NOR2_X1 U19802 ( .A1(n16671), .A2(n16670), .ZN(n16685) );
  NAND3_X1 U19803 ( .A1(P3_REIP_REG_17__SCAN_IN), .A2(P3_REIP_REG_16__SCAN_IN), 
        .A3(P3_REIP_REG_15__SCAN_IN), .ZN(n16687) );
  NAND3_X1 U19804 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(P3_REIP_REG_19__SCAN_IN), 
        .A3(P3_REIP_REG_18__SCAN_IN), .ZN(n16697) );
  NAND2_X1 U19805 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(P3_REIP_REG_21__SCAN_IN), 
        .ZN(n16691) );
  NOR3_X1 U19806 ( .A1(n16687), .A2(n16697), .A3(n16691), .ZN(n16674) );
  NAND3_X1 U19807 ( .A1(P3_REIP_REG_23__SCAN_IN), .A2(n16685), .A3(n16674), 
        .ZN(n16662) );
  NOR2_X1 U19808 ( .A1(n18809), .A2(n16662), .ZN(n16654) );
  NAND2_X1 U19809 ( .A1(P3_REIP_REG_25__SCAN_IN), .A2(n16654), .ZN(n16642) );
  NOR2_X1 U19810 ( .A1(n18813), .A2(n16642), .ZN(n16594) );
  NAND2_X1 U19811 ( .A1(n16939), .A2(n16594), .ZN(n16625) );
  NAND2_X1 U19812 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .ZN(n16595) );
  NOR2_X1 U19813 ( .A1(n16625), .A2(n16595), .ZN(n16613) );
  NAND2_X1 U19814 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(n16613), .ZN(n16593) );
  NOR3_X1 U19815 ( .A1(P3_REIP_REG_31__SCAN_IN), .A2(n18825), .A3(n16593), 
        .ZN(n16591) );
  INV_X1 U19816 ( .A(n18745), .ZN(n18620) );
  NOR2_X1 U19817 ( .A1(n18747), .A2(n18620), .ZN(n18740) );
  NOR4_X2 U19818 ( .A1(n18231), .A2(n18904), .A3(n16882), .A4(n18740), .ZN(
        n16930) );
  INV_X1 U19819 ( .A(P3_EBX_REG_31__SCAN_IN), .ZN(n21123) );
  AOI211_X4 U19820 ( .C1(P3_EBX_REG_31__SCAN_IN), .C2(n16589), .A(n16588), .B(
        n16587), .ZN(n16950) );
  OAI22_X1 U19821 ( .A1(n20969), .A2(n16925), .B1(n21123), .B2(n16955), .ZN(
        n16590) );
  AOI211_X1 U19822 ( .C1(n16607), .C2(n16592), .A(n16591), .B(n16590), .ZN(
        n16597) );
  NOR2_X1 U19823 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n16593), .ZN(n16605) );
  OR2_X1 U19824 ( .A1(n16946), .A2(n16594), .ZN(n16641) );
  NAND2_X1 U19825 ( .A1(n16958), .A2(n16641), .ZN(n16639) );
  AOI221_X1 U19826 ( .B1(n18819), .B2(n16939), .C1(n16595), .C2(n16939), .A(
        n16639), .ZN(n16603) );
  INV_X1 U19827 ( .A(n16603), .ZN(n16612) );
  OAI21_X1 U19828 ( .B1(n16605), .B2(n16612), .A(P3_REIP_REG_31__SCAN_IN), 
        .ZN(n16596) );
  OAI211_X1 U19829 ( .C1(n16598), .C2(n16826), .A(n16597), .B(n16596), .ZN(
        P3_U2640) );
  NAND2_X1 U19830 ( .A1(n16936), .A2(n16599), .ZN(n16619) );
  XNOR2_X1 U19831 ( .A(n16601), .B(n16600), .ZN(n16606) );
  OAI22_X1 U19832 ( .A1(n16603), .A2(n18825), .B1(n16602), .B2(n16925), .ZN(
        n16604) );
  AOI211_X1 U19833 ( .C1(n16606), .C2(n16882), .A(n16605), .B(n16604), .ZN(
        n16609) );
  OAI21_X1 U19834 ( .B1(n16950), .B2(n16607), .A(P3_EBX_REG_30__SCAN_IN), .ZN(
        n16608) );
  OAI211_X1 U19835 ( .C1(P3_EBX_REG_30__SCAN_IN), .C2(n16619), .A(n16609), .B(
        n16608), .ZN(P3_U2641) );
  NOR2_X1 U19836 ( .A1(n16621), .A2(n16992), .ZN(n16620) );
  OAI22_X1 U19837 ( .A1(n16610), .A2(n16925), .B1(n16955), .B2(n16992), .ZN(
        n16611) );
  AOI221_X1 U19838 ( .B1(n16613), .B2(n18819), .C1(n16612), .C2(
        P3_REIP_REG_29__SCAN_IN), .A(n16611), .ZN(n16618) );
  OAI211_X1 U19839 ( .C1(n16616), .C2(n16615), .A(n16882), .B(n16614), .ZN(
        n16617) );
  OAI211_X1 U19840 ( .C1(n16620), .C2(n16619), .A(n16618), .B(n16617), .ZN(
        P3_U2642) );
  AOI22_X1 U19841 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n16944), .B1(
        n16950), .B2(P3_EBX_REG_28__SCAN_IN), .ZN(n16629) );
  NOR2_X1 U19842 ( .A1(P3_REIP_REG_27__SCAN_IN), .A2(n16625), .ZN(n16631) );
  AOI211_X1 U19843 ( .C1(P3_EBX_REG_28__SCAN_IN), .C2(n16632), .A(n16621), .B(
        n16954), .ZN(n16622) );
  AOI221_X1 U19844 ( .B1(n16631), .B2(P3_REIP_REG_28__SCAN_IN), .C1(n16639), 
        .C2(P3_REIP_REG_28__SCAN_IN), .A(n16622), .ZN(n16628) );
  OAI211_X1 U19845 ( .C1(n17550), .C2(n16624), .A(n16882), .B(n16623), .ZN(
        n16627) );
  INV_X1 U19846 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n18815) );
  OR3_X1 U19847 ( .A1(n18815), .A2(n16625), .A3(P3_REIP_REG_28__SCAN_IN), .ZN(
        n16626) );
  NAND4_X1 U19848 ( .A1(n16629), .A2(n16628), .A3(n16627), .A4(n16626), .ZN(
        P3_U2643) );
  OAI22_X1 U19849 ( .A1(n17563), .A2(n16925), .B1(n16955), .B2(n17005), .ZN(
        n16630) );
  AOI211_X1 U19850 ( .C1(P3_REIP_REG_27__SCAN_IN), .C2(n16639), .A(n16631), 
        .B(n16630), .ZN(n16638) );
  OAI211_X1 U19851 ( .C1(n16640), .C2(n17005), .A(n16936), .B(n16632), .ZN(
        n16637) );
  OAI211_X1 U19852 ( .C1(n16635), .C2(n16634), .A(n16882), .B(n16633), .ZN(
        n16636) );
  NAND3_X1 U19853 ( .A1(n16638), .A2(n16637), .A3(n16636), .ZN(P3_U2644) );
  INV_X1 U19854 ( .A(n16639), .ZN(n16649) );
  AOI211_X1 U19855 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n16650), .A(n16640), .B(
        n16954), .ZN(n16644) );
  OAI22_X1 U19856 ( .A1(n17574), .A2(n16925), .B1(n16642), .B2(n16641), .ZN(
        n16643) );
  AOI211_X1 U19857 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n16950), .A(n16644), .B(
        n16643), .ZN(n16648) );
  OAI211_X1 U19858 ( .C1(n17576), .C2(n16646), .A(n16914), .B(n16645), .ZN(
        n16647) );
  OAI211_X1 U19859 ( .C1(n16649), .C2(n18813), .A(n16648), .B(n16647), .ZN(
        P3_U2645) );
  INV_X1 U19860 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n18811) );
  AOI21_X1 U19861 ( .B1(n16939), .B2(n16662), .A(n16930), .ZN(n16669) );
  NAND2_X1 U19862 ( .A1(n16939), .A2(n18809), .ZN(n16661) );
  AOI22_X1 U19863 ( .A1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n16944), .B1(
        n16950), .B2(P3_EBX_REG_25__SCAN_IN), .ZN(n16658) );
  OAI211_X1 U19864 ( .C1(n16660), .C2(n16651), .A(n16936), .B(n16650), .ZN(
        n16657) );
  OAI211_X1 U19865 ( .C1(n17587), .C2(n16653), .A(n16882), .B(n16652), .ZN(
        n16656) );
  NAND3_X1 U19866 ( .A1(n16939), .A2(n16654), .A3(n18811), .ZN(n16655) );
  AND4_X1 U19867 ( .A1(n16658), .A2(n16657), .A3(n16656), .A4(n16655), .ZN(
        n16659) );
  OAI221_X1 U19868 ( .B1(n18811), .B2(n16669), .C1(n18811), .C2(n16661), .A(
        n16659), .ZN(P3_U2646) );
  AOI211_X1 U19869 ( .C1(P3_EBX_REG_24__SCAN_IN), .C2(n16679), .A(n16660), .B(
        n16954), .ZN(n16664) );
  OAI22_X1 U19870 ( .A1(n17603), .A2(n16925), .B1(n16662), .B2(n16661), .ZN(
        n16663) );
  AOI211_X1 U19871 ( .C1(P3_EBX_REG_24__SCAN_IN), .C2(n16950), .A(n16664), .B(
        n16663), .ZN(n16668) );
  OAI211_X1 U19872 ( .C1(n17600), .C2(n16666), .A(n16882), .B(n16665), .ZN(
        n16667) );
  OAI211_X1 U19873 ( .C1(n16669), .C2(n18809), .A(n16668), .B(n16667), .ZN(
        P3_U2647) );
  AOI22_X1 U19874 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n16944), .B1(
        n16950), .B2(P3_EBX_REG_23__SCAN_IN), .ZN(n16684) );
  INV_X1 U19875 ( .A(n16669), .ZN(n16675) );
  INV_X1 U19876 ( .A(n16670), .ZN(n16672) );
  NOR2_X1 U19877 ( .A1(n16946), .A2(n16671), .ZN(n16786) );
  NAND2_X1 U19878 ( .A1(n16672), .A2(n16786), .ZN(n16765) );
  NOR2_X1 U19879 ( .A1(P3_REIP_REG_23__SCAN_IN), .A2(n16765), .ZN(n16673) );
  AOI22_X1 U19880 ( .A1(P3_REIP_REG_23__SCAN_IN), .A2(n16675), .B1(n16674), 
        .B2(n16673), .ZN(n16683) );
  OAI211_X1 U19881 ( .C1(n16678), .C2(n16677), .A(n16882), .B(n16676), .ZN(
        n16682) );
  OAI211_X1 U19882 ( .C1(n16688), .C2(n16680), .A(n16936), .B(n16679), .ZN(
        n16681) );
  NAND4_X1 U19883 ( .A1(n16684), .A2(n16683), .A3(n16682), .A4(n16681), .ZN(
        P3_U2648) );
  NAND2_X1 U19884 ( .A1(n16946), .A2(n16958), .ZN(n16956) );
  NAND2_X1 U19885 ( .A1(n16685), .A2(n16958), .ZN(n16776) );
  OAI21_X1 U19886 ( .B1(n16687), .B2(n16776), .A(n16956), .ZN(n16686) );
  INV_X1 U19887 ( .A(n16686), .ZN(n16744) );
  AOI21_X1 U19888 ( .B1(n16697), .B2(n16956), .A(n16744), .ZN(n16716) );
  INV_X1 U19889 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n18806) );
  INV_X1 U19890 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n18804) );
  AOI211_X1 U19891 ( .C1(n18806), .C2(n18804), .A(n16697), .B(n16724), .ZN(
        n16692) );
  AOI211_X1 U19892 ( .C1(P3_EBX_REG_22__SCAN_IN), .C2(n16702), .A(n16688), .B(
        n16954), .ZN(n16690) );
  INV_X1 U19893 ( .A(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n17632) );
  INV_X1 U19894 ( .A(P3_EBX_REG_22__SCAN_IN), .ZN(n17021) );
  OAI22_X1 U19895 ( .A1(n17632), .A2(n16925), .B1(n16955), .B2(n17021), .ZN(
        n16689) );
  AOI211_X1 U19896 ( .C1(n16692), .C2(n16691), .A(n16690), .B(n16689), .ZN(
        n16696) );
  OAI211_X1 U19897 ( .C1(n17645), .C2(n16694), .A(n16882), .B(n16693), .ZN(
        n16695) );
  OAI211_X1 U19898 ( .C1(n16716), .C2(n18806), .A(n16696), .B(n16695), .ZN(
        P3_U2649) );
  AOI22_X1 U19899 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n16944), .B1(
        n16950), .B2(P3_EBX_REG_21__SCAN_IN), .ZN(n16706) );
  INV_X1 U19900 ( .A(n16716), .ZN(n16699) );
  NOR2_X1 U19901 ( .A1(n16697), .A2(n16724), .ZN(n16698) );
  AOI22_X1 U19902 ( .A1(P3_REIP_REG_21__SCAN_IN), .A2(n16699), .B1(n16698), 
        .B2(n18804), .ZN(n16705) );
  OAI211_X1 U19903 ( .C1(n17646), .C2(n16701), .A(n16882), .B(n16700), .ZN(
        n16704) );
  OAI211_X1 U19904 ( .C1(n16707), .C2(n17026), .A(n16936), .B(n16702), .ZN(
        n16703) );
  NAND4_X1 U19905 ( .A1(n16706), .A2(n16705), .A3(n16704), .A4(n16703), .ZN(
        P3_U2650) );
  INV_X1 U19906 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n18803) );
  INV_X1 U19907 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n18800) );
  INV_X1 U19908 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n18798) );
  NOR4_X1 U19909 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(n18800), .A3(n18798), 
        .A4(n16724), .ZN(n16710) );
  AOI211_X1 U19910 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n16719), .A(n16707), .B(
        n16954), .ZN(n16709) );
  INV_X1 U19911 ( .A(P3_EBX_REG_20__SCAN_IN), .ZN(n16961) );
  OAI22_X1 U19912 ( .A1(n17663), .A2(n16925), .B1(n16955), .B2(n16961), .ZN(
        n16708) );
  NOR3_X1 U19913 ( .A1(n16710), .A2(n16709), .A3(n16708), .ZN(n16715) );
  OAI211_X1 U19914 ( .C1(n16713), .C2(n16712), .A(n16914), .B(n16711), .ZN(
        n16714) );
  OAI211_X1 U19915 ( .C1(n16716), .C2(n18803), .A(n16715), .B(n16714), .ZN(
        P3_U2651) );
  INV_X1 U19916 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n16738) );
  NOR2_X1 U19917 ( .A1(n16730), .A2(n16738), .ZN(n16717) );
  OAI21_X1 U19918 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n16717), .A(
        n17629), .ZN(n17674) );
  NAND2_X1 U19919 ( .A1(n17670), .A2(n16888), .ZN(n16731) );
  OAI21_X1 U19920 ( .B1(n16738), .B2(n16731), .A(n16789), .ZN(n16718) );
  XNOR2_X1 U19921 ( .A(n17674), .B(n16718), .ZN(n16727) );
  NOR3_X1 U19922 ( .A1(P3_REIP_REG_19__SCAN_IN), .A2(n18798), .A3(n16724), 
        .ZN(n16723) );
  OAI211_X1 U19923 ( .C1(n16728), .C2(n16721), .A(n16936), .B(n16719), .ZN(
        n16720) );
  OAI211_X1 U19924 ( .C1(n16955), .C2(n16721), .A(n18218), .B(n16720), .ZN(
        n16722) );
  AOI211_X1 U19925 ( .C1(n16944), .C2(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n16723), .B(n16722), .ZN(n16726) );
  NOR2_X1 U19926 ( .A1(P3_REIP_REG_18__SCAN_IN), .A2(n16724), .ZN(n16735) );
  OAI21_X1 U19927 ( .B1(n16744), .B2(n16735), .A(P3_REIP_REG_19__SCAN_IN), 
        .ZN(n16725) );
  OAI211_X1 U19928 ( .C1(n18750), .C2(n16727), .A(n16726), .B(n16725), .ZN(
        P3_U2652) );
  AOI211_X1 U19929 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n16745), .A(n16728), .B(
        n16954), .ZN(n16729) );
  AOI211_X1 U19930 ( .C1(n16950), .C2(P3_EBX_REG_18__SCAN_IN), .A(n18231), .B(
        n16729), .ZN(n16737) );
  AOI22_X1 U19931 ( .A1(n17670), .A2(n16738), .B1(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n16730), .ZN(n17681) );
  NAND2_X1 U19932 ( .A1(n16789), .A2(n16731), .ZN(n16733) );
  OAI21_X1 U19933 ( .B1(n17681), .B2(n16733), .A(n16914), .ZN(n16732) );
  AOI21_X1 U19934 ( .B1(n17681), .B2(n16733), .A(n16732), .ZN(n16734) );
  AOI211_X1 U19935 ( .C1(n16744), .C2(P3_REIP_REG_18__SCAN_IN), .A(n16735), 
        .B(n16734), .ZN(n16736) );
  OAI211_X1 U19936 ( .C1(n16738), .C2(n16925), .A(n16737), .B(n16736), .ZN(
        P3_U2653) );
  AOI22_X1 U19937 ( .A1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n16944), .B1(
        n16950), .B2(P3_EBX_REG_17__SCAN_IN), .ZN(n16749) );
  INV_X1 U19938 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n20933) );
  INV_X1 U19939 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n18793) );
  NOR4_X1 U19940 ( .A1(P3_REIP_REG_17__SCAN_IN), .A2(n20933), .A3(n18793), 
        .A4(n16765), .ZN(n16743) );
  AOI21_X1 U19941 ( .B1(n16750), .B2(n17693), .A(n17670), .ZN(n17698) );
  INV_X1 U19942 ( .A(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n17715) );
  OAI21_X1 U19943 ( .B1(n17715), .B2(n16753), .A(n16789), .ZN(n16739) );
  INV_X1 U19944 ( .A(n16739), .ZN(n16741) );
  OAI21_X1 U19945 ( .B1(n17698), .B2(n16741), .A(n16914), .ZN(n16740) );
  AOI21_X1 U19946 ( .B1(n17698), .B2(n16741), .A(n16740), .ZN(n16742) );
  AOI211_X1 U19947 ( .C1(n16744), .C2(P3_REIP_REG_17__SCAN_IN), .A(n16743), 
        .B(n16742), .ZN(n16748) );
  OAI211_X1 U19948 ( .C1(n16754), .C2(n16746), .A(n16936), .B(n16745), .ZN(
        n16747) );
  NAND4_X1 U19949 ( .A1(n16749), .A2(n16748), .A3(n18218), .A4(n16747), .ZN(
        P3_U2654) );
  OAI21_X1 U19950 ( .B1(n16751), .B2(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n16750), .ZN(n16752) );
  INV_X1 U19951 ( .A(n16752), .ZN(n17711) );
  INV_X1 U19952 ( .A(n16826), .ZN(n16945) );
  NAND2_X1 U19953 ( .A1(n16945), .A2(n16753), .ZN(n16773) );
  AOI22_X1 U19954 ( .A1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n16944), .B1(
        n16950), .B2(P3_EBX_REG_16__SCAN_IN), .ZN(n16761) );
  AOI211_X1 U19955 ( .C1(n16789), .C2(n16753), .A(n18750), .B(n16752), .ZN(
        n16759) );
  AOI211_X1 U19956 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n16766), .A(n16754), .B(
        n16954), .ZN(n16758) );
  NOR2_X1 U19957 ( .A1(n18793), .A2(n16765), .ZN(n16756) );
  OAI21_X1 U19958 ( .B1(n18793), .B2(n16776), .A(n16956), .ZN(n16764) );
  INV_X1 U19959 ( .A(n16764), .ZN(n16755) );
  MUX2_X1 U19960 ( .A(n16756), .B(n16755), .S(P3_REIP_REG_16__SCAN_IN), .Z(
        n16757) );
  NOR4_X1 U19961 ( .A1(n18231), .A2(n16759), .A3(n16758), .A4(n16757), .ZN(
        n16760) );
  OAI211_X1 U19962 ( .C1(n17711), .C2(n16773), .A(n16761), .B(n16760), .ZN(
        P3_U2655) );
  OAI21_X1 U19963 ( .B1(n17710), .B2(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A(
        n16762), .ZN(n17722) );
  INV_X1 U19964 ( .A(n17722), .ZN(n16774) );
  NOR2_X1 U19965 ( .A1(n18750), .A2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n16835) );
  NAND2_X1 U19966 ( .A1(n16882), .A2(n9843), .ZN(n16927) );
  INV_X1 U19967 ( .A(n16927), .ZN(n16763) );
  AOI21_X1 U19968 ( .B1(n17710), .B2(n16835), .A(n16763), .ZN(n16772) );
  AOI21_X1 U19969 ( .B1(n18793), .B2(n16765), .A(n16764), .ZN(n16770) );
  OAI211_X1 U19970 ( .C1(n16775), .C2(n16768), .A(n16936), .B(n16766), .ZN(
        n16767) );
  OAI211_X1 U19971 ( .C1(n16955), .C2(n16768), .A(n18218), .B(n16767), .ZN(
        n16769) );
  AOI211_X1 U19972 ( .C1(n16944), .C2(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A(
        n16770), .B(n16769), .ZN(n16771) );
  OAI221_X1 U19973 ( .B1(n16774), .B2(n16773), .C1(n17722), .C2(n16772), .A(
        n16771), .ZN(P3_U2656) );
  AOI211_X1 U19974 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n16790), .A(n16775), .B(
        n16954), .ZN(n16784) );
  INV_X1 U19975 ( .A(n16776), .ZN(n16782) );
  AOI22_X1 U19976 ( .A1(P3_REIP_REG_14__SCAN_IN), .A2(n16956), .B1(
        P3_REIP_REG_13__SCAN_IN), .B2(n16786), .ZN(n16781) );
  INV_X1 U19977 ( .A(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n16778) );
  INV_X1 U19978 ( .A(n17744), .ZN(n16788) );
  OR2_X1 U19979 ( .A1(n17748), .A2(n16788), .ZN(n16777) );
  AOI21_X1 U19980 ( .B1(n16778), .B2(n16777), .A(n17710), .ZN(n17734) );
  INV_X1 U19981 ( .A(n16779), .ZN(n16874) );
  NOR2_X1 U19982 ( .A1(n16874), .A2(n17810), .ZN(n16855) );
  NAND2_X1 U19983 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n16855), .ZN(
        n16839) );
  NOR2_X1 U19984 ( .A1(n16839), .A2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n16831) );
  AOI21_X1 U19985 ( .B1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n16831), .A(
        n9843), .ZN(n16811) );
  INV_X1 U19986 ( .A(n16811), .ZN(n16810) );
  OAI21_X1 U19987 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n9843), .A(
        n16810), .ZN(n16804) );
  AOI21_X1 U19988 ( .B1(n16789), .B2(n16788), .A(n16804), .ZN(n16787) );
  XOR2_X1 U19989 ( .A(n17734), .B(n16787), .Z(n16780) );
  OAI22_X1 U19990 ( .A1(n16782), .A2(n16781), .B1(n18750), .B2(n16780), .ZN(
        n16783) );
  AOI211_X1 U19991 ( .C1(n16944), .C2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n16784), .B(n16783), .ZN(n16785) );
  OAI211_X1 U19992 ( .C1(n16955), .C2(n20937), .A(n16785), .B(n18218), .ZN(
        P3_U2657) );
  INV_X1 U19993 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n18790) );
  AOI22_X1 U19994 ( .A1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n16944), .B1(
        n16786), .B2(n18790), .ZN(n16798) );
  NOR2_X1 U19995 ( .A1(n16787), .A2(n18750), .ZN(n16795) );
  NOR2_X1 U19996 ( .A1(n17748), .A2(n17763), .ZN(n16803) );
  OAI22_X1 U19997 ( .A1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n16803), .B1(
        n17748), .B2(n16788), .ZN(n17749) );
  OAI21_X1 U19998 ( .B1(n9843), .B2(n16888), .A(n16914), .ZN(n16953) );
  AOI211_X1 U19999 ( .C1(n16789), .C2(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A(
        n16953), .B(n17749), .ZN(n16794) );
  OAI211_X1 U20000 ( .C1(n16799), .C2(n16792), .A(n16936), .B(n16790), .ZN(
        n16791) );
  OAI21_X1 U20001 ( .B1(n16792), .B2(n16955), .A(n16791), .ZN(n16793) );
  AOI211_X1 U20002 ( .C1(n16795), .C2(n17749), .A(n16794), .B(n16793), .ZN(
        n16797) );
  OAI21_X1 U20003 ( .B1(n16802), .B2(n16946), .A(n16958), .ZN(n16819) );
  NOR2_X1 U20004 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n16946), .ZN(n16801) );
  OAI21_X1 U20005 ( .B1(n16819), .B2(n16801), .A(P3_REIP_REG_13__SCAN_IN), 
        .ZN(n16796) );
  NAND4_X1 U20006 ( .A1(n16798), .A2(n16797), .A3(n18218), .A4(n16796), .ZN(
        P3_U2658) );
  AOI211_X1 U20007 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n16813), .A(n16799), .B(
        n16954), .ZN(n16800) );
  AOI21_X1 U20008 ( .B1(n16944), .B2(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n16800), .ZN(n16808) );
  AOI22_X1 U20009 ( .A1(n16950), .A2(P3_EBX_REG_12__SCAN_IN), .B1(n16802), 
        .B2(n16801), .ZN(n16807) );
  AOI21_X1 U20010 ( .B1(n17748), .B2(n17763), .A(n16803), .ZN(n17766) );
  XOR2_X1 U20011 ( .A(n17766), .B(n16804), .Z(n16805) );
  AOI22_X1 U20012 ( .A1(n16914), .A2(n16805), .B1(P3_REIP_REG_12__SCAN_IN), 
        .B2(n16819), .ZN(n16806) );
  NAND4_X1 U20013 ( .A1(n16808), .A2(n16807), .A3(n16806), .A4(n18218), .ZN(
        P3_U2659) );
  INV_X1 U20014 ( .A(n16809), .ZN(n16827) );
  NAND2_X1 U20015 ( .A1(n16939), .A2(n16827), .ZN(n16849) );
  OAI21_X1 U20016 ( .B1(n16822), .B2(n16849), .A(n18786), .ZN(n16818) );
  NOR2_X1 U20017 ( .A1(n17789), .A2(n16839), .ZN(n16825) );
  OAI21_X1 U20018 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n16825), .A(
        n17748), .ZN(n17779) );
  INV_X1 U20019 ( .A(n17779), .ZN(n16812) );
  OAI221_X1 U20020 ( .B1(n16812), .B2(n16811), .C1(n17779), .C2(n16810), .A(
        n16914), .ZN(n16815) );
  OAI211_X1 U20021 ( .C1(n16823), .C2(n16821), .A(n16936), .B(n16813), .ZN(
        n16814) );
  OAI211_X1 U20022 ( .C1(n16925), .C2(n16816), .A(n16815), .B(n16814), .ZN(
        n16817) );
  AOI21_X1 U20023 ( .B1(n16819), .B2(n16818), .A(n16817), .ZN(n16820) );
  OAI211_X1 U20024 ( .C1(n16955), .C2(n16821), .A(n16820), .B(n18218), .ZN(
        P3_U2660) );
  OAI21_X1 U20025 ( .B1(P3_REIP_REG_10__SCAN_IN), .B2(P3_REIP_REG_9__SCAN_IN), 
        .A(n16822), .ZN(n16834) );
  AOI211_X1 U20026 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n16824), .A(n16823), .B(
        n16954), .ZN(n16830) );
  OAI22_X1 U20027 ( .A1(n17789), .A2(n16925), .B1(n16955), .B2(n17189), .ZN(
        n16829) );
  AOI21_X1 U20028 ( .B1(n17789), .B2(n16839), .A(n16825), .ZN(n17792) );
  OR2_X1 U20029 ( .A1(n16826), .A2(n16831), .ZN(n16843) );
  NOR2_X1 U20030 ( .A1(n16946), .A2(n16827), .ZN(n16852) );
  NOR2_X1 U20031 ( .A1(n16930), .A2(n16852), .ZN(n16838) );
  INV_X1 U20032 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n18784) );
  OAI22_X1 U20033 ( .A1(n17792), .A2(n16843), .B1(n16838), .B2(n18784), .ZN(
        n16828) );
  NOR4_X1 U20034 ( .A1(n18231), .A2(n16830), .A3(n16829), .A4(n16828), .ZN(
        n16833) );
  OAI211_X1 U20035 ( .C1(n16831), .C2(n9843), .A(n16914), .B(n17792), .ZN(
        n16832) );
  OAI211_X1 U20036 ( .C1(n16849), .C2(n16834), .A(n16833), .B(n16832), .ZN(
        P3_U2661) );
  AND2_X1 U20037 ( .A1(n16855), .A2(n16835), .ZN(n16837) );
  AOI221_X1 U20038 ( .B1(n16944), .B2(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .C1(
        n16837), .C2(n16836), .A(n18231), .ZN(n16848) );
  INV_X1 U20039 ( .A(n16838), .ZN(n16858) );
  OR2_X1 U20040 ( .A1(n16954), .A2(n16840), .ZN(n16850) );
  OAI21_X1 U20041 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n16855), .A(
        n16839), .ZN(n17803) );
  OAI22_X1 U20042 ( .A1(P3_EBX_REG_9__SCAN_IN), .A2(n16850), .B1(n16927), .B2(
        n17803), .ZN(n16846) );
  INV_X1 U20043 ( .A(n17803), .ZN(n16844) );
  AOI21_X1 U20044 ( .B1(n16936), .B2(n16840), .A(n16950), .ZN(n16841) );
  OAI22_X1 U20045 ( .A1(n16844), .A2(n16843), .B1(n16842), .B2(n16841), .ZN(
        n16845) );
  AOI211_X1 U20046 ( .C1(P3_REIP_REG_9__SCAN_IN), .C2(n16858), .A(n16846), .B(
        n16845), .ZN(n16847) );
  OAI211_X1 U20047 ( .C1(P3_REIP_REG_9__SCAN_IN), .C2(n16849), .A(n16848), .B(
        n16847), .ZN(P3_U2662) );
  AOI21_X1 U20048 ( .B1(n16867), .B2(P3_EBX_REG_8__SCAN_IN), .A(n16850), .ZN(
        n16851) );
  AOI21_X1 U20049 ( .B1(P3_EBX_REG_8__SCAN_IN), .B2(n16950), .A(n16851), .ZN(
        n16862) );
  AOI22_X1 U20050 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n16944), .B1(
        n16853), .B2(n16852), .ZN(n16861) );
  INV_X1 U20051 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n17827) );
  NOR2_X1 U20052 ( .A1(n16854), .A2(n17827), .ZN(n17811) );
  NOR2_X1 U20053 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n17904), .ZN(
        n16933) );
  AOI21_X1 U20054 ( .B1(n17811), .B2(n16933), .A(n9843), .ZN(n16857) );
  NOR2_X1 U20055 ( .A1(n16874), .A2(n17827), .ZN(n16863) );
  INV_X1 U20056 ( .A(n16855), .ZN(n16856) );
  OAI21_X1 U20057 ( .B1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n16863), .A(
        n16856), .ZN(n17813) );
  XNOR2_X1 U20058 ( .A(n16857), .B(n17813), .ZN(n16859) );
  AOI22_X1 U20059 ( .A1(n16914), .A2(n16859), .B1(P3_REIP_REG_8__SCAN_IN), 
        .B2(n16858), .ZN(n16860) );
  NAND4_X1 U20060 ( .A1(n16862), .A2(n16861), .A3(n16860), .A4(n18218), .ZN(
        P3_U2663) );
  AOI21_X1 U20061 ( .B1(n16868), .B2(n16939), .A(n16930), .ZN(n16891) );
  INV_X1 U20062 ( .A(n16891), .ZN(n16880) );
  AOI21_X1 U20063 ( .B1(n16874), .B2(n17827), .A(n16863), .ZN(n17831) );
  AOI21_X1 U20064 ( .B1(n17746), .B2(n16933), .A(n9843), .ZN(n16881) );
  OAI21_X1 U20065 ( .B1(n17831), .B2(n16881), .A(n16914), .ZN(n16864) );
  AOI21_X1 U20066 ( .B1(n17831), .B2(n16881), .A(n16864), .ZN(n16866) );
  OAI22_X1 U20067 ( .A1(n17827), .A2(n16925), .B1(n16955), .B2(n17237), .ZN(
        n16865) );
  AOI211_X1 U20068 ( .C1(n16880), .C2(P3_REIP_REG_7__SCAN_IN), .A(n16866), .B(
        n16865), .ZN(n16872) );
  OAI211_X1 U20069 ( .C1(n16875), .C2(n17237), .A(n16936), .B(n16867), .ZN(
        n16871) );
  NOR2_X1 U20070 ( .A1(n16946), .A2(n16868), .ZN(n16873) );
  OAI211_X1 U20071 ( .C1(P3_REIP_REG_6__SCAN_IN), .C2(P3_REIP_REG_7__SCAN_IN), 
        .A(n16873), .B(n16869), .ZN(n16870) );
  NAND4_X1 U20072 ( .A1(n16872), .A2(n18218), .A3(n16871), .A4(n16870), .ZN(
        P3_U2664) );
  INV_X1 U20073 ( .A(n16873), .ZN(n16885) );
  NOR2_X1 U20074 ( .A1(n17904), .A2(n17851), .ZN(n16889) );
  INV_X1 U20075 ( .A(n16889), .ZN(n16898) );
  NOR2_X1 U20076 ( .A1(n17852), .A2(n16898), .ZN(n16887) );
  OAI21_X1 U20077 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n16887), .A(
        n16874), .ZN(n17840) );
  AOI211_X1 U20078 ( .C1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .C2(n16927), .A(
        n16953), .B(n17840), .ZN(n16879) );
  INV_X1 U20079 ( .A(P3_EBX_REG_6__SCAN_IN), .ZN(n17239) );
  AOI211_X1 U20080 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n16894), .A(n16875), .B(
        n16954), .ZN(n16876) );
  AOI211_X1 U20081 ( .C1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .C2(n16944), .A(
        n18231), .B(n16876), .ZN(n16877) );
  OAI21_X1 U20082 ( .B1(n16955), .B2(n17239), .A(n16877), .ZN(n16878) );
  AOI211_X1 U20083 ( .C1(n16880), .C2(P3_REIP_REG_6__SCAN_IN), .A(n16879), .B(
        n16878), .ZN(n16884) );
  NAND3_X1 U20084 ( .A1(n16882), .A2(n16881), .A3(n17840), .ZN(n16883) );
  OAI211_X1 U20085 ( .C1(P3_REIP_REG_6__SCAN_IN), .C2(n16885), .A(n16884), .B(
        n16883), .ZN(P3_U2665) );
  AOI21_X1 U20086 ( .B1(n16939), .B2(n16886), .A(P3_REIP_REG_5__SCAN_IN), .ZN(
        n16892) );
  AOI21_X1 U20087 ( .B1(n17852), .B2(n16898), .A(n16887), .ZN(n17854) );
  AOI21_X1 U20088 ( .B1(n16889), .B2(n16888), .A(n9843), .ZN(n16899) );
  XNOR2_X1 U20089 ( .A(n17854), .B(n16899), .ZN(n16890) );
  OAI22_X1 U20090 ( .A1(n16892), .A2(n16891), .B1(n18750), .B2(n16890), .ZN(
        n16893) );
  AOI211_X1 U20091 ( .C1(n16950), .C2(P3_EBX_REG_5__SCAN_IN), .A(n18231), .B(
        n16893), .ZN(n16896) );
  OAI211_X1 U20092 ( .C1(n16904), .C2(n17230), .A(n16936), .B(n16894), .ZN(
        n16895) );
  OAI211_X1 U20093 ( .C1(n16925), .C2(n17852), .A(n16896), .B(n16895), .ZN(
        P3_U2666) );
  INV_X1 U20094 ( .A(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n16902) );
  NAND2_X1 U20095 ( .A1(n17868), .A2(n16902), .ZN(n17862) );
  INV_X1 U20096 ( .A(n17862), .ZN(n16900) );
  INV_X1 U20097 ( .A(n17868), .ZN(n16897) );
  NOR2_X1 U20098 ( .A1(n17904), .A2(n16897), .ZN(n16912) );
  OAI21_X1 U20099 ( .B1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n16912), .A(
        n16898), .ZN(n17871) );
  AOI22_X1 U20100 ( .A1(n16933), .A2(n16900), .B1(n16899), .B2(n17871), .ZN(
        n16911) );
  AOI21_X1 U20101 ( .B1(n16903), .B2(n16939), .A(n16930), .ZN(n16901) );
  INV_X1 U20102 ( .A(n16901), .ZN(n16920) );
  OAI22_X1 U20103 ( .A1(n16902), .A2(n16925), .B1(n17871), .B2(n16927), .ZN(
        n16909) );
  NAND2_X1 U20104 ( .A1(n18248), .A2(n18904), .ZN(n18907) );
  NOR3_X1 U20105 ( .A1(P3_REIP_REG_4__SCAN_IN), .A2(n16946), .A3(n16903), .ZN(
        n16906) );
  AOI211_X1 U20106 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n16921), .A(n16904), .B(
        n16954), .ZN(n16905) );
  AOI211_X1 U20107 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n16950), .A(n16906), .B(
        n16905), .ZN(n16907) );
  OAI221_X1 U20108 ( .B1(n18907), .B2(n9887), .C1(n18907), .C2(n18691), .A(
        n16907), .ZN(n16908) );
  AOI211_X1 U20109 ( .C1(P3_REIP_REG_4__SCAN_IN), .C2(n16920), .A(n16909), .B(
        n16908), .ZN(n16910) );
  OAI211_X1 U20110 ( .C1(n16911), .C2(n18750), .A(n16910), .B(n18218), .ZN(
        P3_U2667) );
  NAND2_X1 U20111 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_2__SCAN_IN), 
        .ZN(n16938) );
  INV_X1 U20112 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n18773) );
  OAI21_X1 U20113 ( .B1(n16946), .B2(n16938), .A(n18773), .ZN(n16919) );
  NAND2_X1 U20114 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n16926) );
  AOI21_X1 U20115 ( .B1(n16924), .B2(n16926), .A(n16912), .ZN(n17875) );
  NOR2_X1 U20116 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n16926), .ZN(
        n16931) );
  NOR2_X1 U20117 ( .A1(n16931), .A2(n9843), .ZN(n16916) );
  OAI21_X1 U20118 ( .B1(n17875), .B2(n16916), .A(n16914), .ZN(n16915) );
  AOI21_X1 U20119 ( .B1(n17875), .B2(n16916), .A(n16915), .ZN(n16918) );
  NOR2_X1 U20120 ( .A1(n18870), .A2(n18700), .ZN(n18697) );
  OAI21_X1 U20121 ( .B1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n18697), .A(
        n9887), .ZN(n18838) );
  OAI22_X1 U20122 ( .A1(n16955), .A2(n17252), .B1(n18907), .B2(n18838), .ZN(
        n16917) );
  AOI211_X1 U20123 ( .C1(n16920), .C2(n16919), .A(n16918), .B(n16917), .ZN(
        n16923) );
  OAI211_X1 U20124 ( .C1(n16934), .C2(n17252), .A(n16936), .B(n16921), .ZN(
        n16922) );
  OAI211_X1 U20125 ( .C1(n16925), .C2(n16924), .A(n16923), .B(n16922), .ZN(
        P3_U2668) );
  OAI22_X1 U20126 ( .A1(n17888), .A2(n16925), .B1(n16955), .B2(n17256), .ZN(
        n16929) );
  NAND2_X1 U20127 ( .A1(n18854), .A2(n18705), .ZN(n18696) );
  OAI21_X1 U20128 ( .B1(n18700), .B2(n18870), .A(n18696), .ZN(n18847) );
  OAI21_X1 U20129 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n16926), .ZN(n17896) );
  OAI22_X1 U20130 ( .A1(n18847), .A2(n18907), .B1(n17896), .B2(n16927), .ZN(
        n16928) );
  AOI211_X1 U20131 ( .C1(P3_REIP_REG_2__SCAN_IN), .C2(n16930), .A(n16929), .B(
        n16928), .ZN(n16943) );
  INV_X1 U20132 ( .A(n16931), .ZN(n16932) );
  OAI211_X1 U20133 ( .C1(n16933), .C2(n17896), .A(n16945), .B(n16932), .ZN(
        n16942) );
  NOR2_X1 U20134 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n16937) );
  INV_X1 U20135 ( .A(n16934), .ZN(n16935) );
  OAI211_X1 U20136 ( .C1(n16937), .C2(n17256), .A(n16936), .B(n16935), .ZN(
        n16941) );
  OAI211_X1 U20137 ( .C1(P3_REIP_REG_1__SCAN_IN), .C2(P3_REIP_REG_2__SCAN_IN), 
        .A(n16939), .B(n16938), .ZN(n16940) );
  NAND4_X1 U20138 ( .A1(n16943), .A2(n16942), .A3(n16941), .A4(n16940), .ZN(
        P3_U2669) );
  AOI21_X1 U20139 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16945), .A(
        n16944), .ZN(n16952) );
  OAI21_X1 U20140 ( .B1(P3_EBX_REG_0__SCAN_IN), .B2(P3_EBX_REG_1__SCAN_IN), 
        .A(n17257), .ZN(n17262) );
  OAI22_X1 U20141 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n16946), .B1(n16954), 
        .B2(n17262), .ZN(n16949) );
  NAND2_X1 U20142 ( .A1(n18705), .A2(n16947), .ZN(n18855) );
  OAI22_X1 U20143 ( .A1(n20815), .A2(n16958), .B1(n18855), .B2(n18907), .ZN(
        n16948) );
  AOI211_X1 U20144 ( .C1(n16950), .C2(P3_EBX_REG_1__SCAN_IN), .A(n16949), .B(
        n16948), .ZN(n16951) );
  OAI221_X1 U20145 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n16953), .C1(
        n17904), .C2(n16952), .A(n16951), .ZN(P3_U2670) );
  NAND2_X1 U20146 ( .A1(n16955), .A2(n16954), .ZN(n16957) );
  AOI22_X1 U20147 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(n16957), .B1(
        P3_REIP_REG_0__SCAN_IN), .B2(n16956), .ZN(n16960) );
  NAND3_X1 U20148 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n18849), .A3(
        n16958), .ZN(n16959) );
  OAI211_X1 U20149 ( .C1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .C2(n18907), .A(
        n16960), .B(n16959), .ZN(P3_U2671) );
  INV_X1 U20150 ( .A(P3_EBX_REG_26__SCAN_IN), .ZN(n16964) );
  NOR2_X1 U20151 ( .A1(n16961), .A2(n17076), .ZN(n17040) );
  NAND4_X1 U20152 ( .A1(P3_EBX_REG_25__SCAN_IN), .A2(P3_EBX_REG_24__SCAN_IN), 
        .A3(n16993), .A4(n17040), .ZN(n16962) );
  NOR4_X1 U20153 ( .A1(n16992), .A2(n16964), .A3(n16963), .A4(n16962), .ZN(
        n16990) );
  NAND2_X1 U20154 ( .A1(P3_EBX_REG_30__SCAN_IN), .A2(n16990), .ZN(n16989) );
  NAND2_X1 U20155 ( .A1(n16989), .A2(P3_EBX_REG_31__SCAN_IN), .ZN(n16966) );
  NAND2_X1 U20156 ( .A1(n18277), .A2(n21123), .ZN(n16965) );
  OAI22_X1 U20157 ( .A1(n17267), .A2(n16966), .B1(n16989), .B2(n16965), .ZN(
        P3_U2672) );
  AOI22_X1 U20158 ( .A1(n17220), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n9838), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n16976) );
  AOI22_X1 U20159 ( .A1(n9851), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(n9849), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n16975) );
  AOI22_X1 U20160 ( .A1(n17192), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n17148), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n16967) );
  OAI21_X1 U20161 ( .B1(n17136), .B2(n21192), .A(n16967), .ZN(n16973) );
  AOI22_X1 U20162 ( .A1(n17200), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17216), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n16971) );
  AOI22_X1 U20163 ( .A1(n17176), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n17211), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n16970) );
  AOI22_X1 U20164 ( .A1(n17199), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n17153), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n16969) );
  AOI22_X1 U20165 ( .A1(n9837), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n9839), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n16968) );
  NAND4_X1 U20166 ( .A1(n16971), .A2(n16970), .A3(n16969), .A4(n16968), .ZN(
        n16972) );
  AOI211_X1 U20167 ( .C1(n17193), .C2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A(
        n16973), .B(n16972), .ZN(n16974) );
  NAND3_X1 U20168 ( .A1(n16976), .A2(n16975), .A3(n16974), .ZN(n16988) );
  AOI22_X1 U20169 ( .A1(n9838), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17213), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n16980) );
  AOI22_X1 U20170 ( .A1(n17219), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17147), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n16979) );
  AOI22_X1 U20171 ( .A1(n17212), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n17148), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n16978) );
  AOI22_X1 U20172 ( .A1(n17193), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17194), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n16977) );
  NAND4_X1 U20173 ( .A1(n16980), .A2(n16979), .A3(n16978), .A4(n16977), .ZN(
        n16986) );
  AOI22_X1 U20174 ( .A1(n17176), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17211), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n16984) );
  AOI22_X1 U20175 ( .A1(n9849), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(n9839), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n16983) );
  AOI22_X1 U20176 ( .A1(n17200), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17098), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n16982) );
  AOI22_X1 U20177 ( .A1(n17220), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n9837), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n16981) );
  NAND4_X1 U20178 ( .A1(n16984), .A2(n16983), .A3(n16982), .A4(n16981), .ZN(
        n16985) );
  NOR2_X1 U20179 ( .A1(n16986), .A2(n16985), .ZN(n16996) );
  INV_X1 U20180 ( .A(n17001), .ZN(n16995) );
  NOR3_X1 U20181 ( .A1(n16996), .A2(n16994), .A3(n16995), .ZN(n16987) );
  XNOR2_X1 U20182 ( .A(n16988), .B(n16987), .ZN(n17280) );
  OAI211_X1 U20183 ( .C1(P3_EBX_REG_30__SCAN_IN), .C2(n16990), .A(n16989), .B(
        n14394), .ZN(n16991) );
  OAI21_X1 U20184 ( .B1(n17280), .B2(n17260), .A(n16991), .ZN(P3_U2673) );
  NAND2_X1 U20185 ( .A1(n16993), .A2(n16992), .ZN(n17000) );
  NOR2_X1 U20186 ( .A1(n16995), .A2(n16994), .ZN(n16997) );
  XNOR2_X1 U20187 ( .A(n16997), .B(n16996), .ZN(n17281) );
  AOI22_X1 U20188 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n16998), .B1(n17267), 
        .B2(n17281), .ZN(n16999) );
  OAI21_X1 U20189 ( .B1(n17006), .B2(n17000), .A(n16999), .ZN(P3_U2674) );
  AOI21_X1 U20190 ( .B1(n17002), .B2(n17007), .A(n17001), .ZN(n17290) );
  NAND2_X1 U20191 ( .A1(n17267), .A2(n17290), .ZN(n17003) );
  OAI221_X1 U20192 ( .B1(P3_EBX_REG_27__SCAN_IN), .B2(n17006), .C1(n17005), 
        .C2(n17004), .A(n17003), .ZN(P3_U2676) );
  AOI21_X1 U20193 ( .B1(P3_EBX_REG_26__SCAN_IN), .B2(n17260), .A(n17015), .ZN(
        n17010) );
  OAI21_X1 U20194 ( .B1(n17009), .B2(n17008), .A(n17007), .ZN(n17298) );
  OAI22_X1 U20195 ( .A1(n17011), .A2(n17010), .B1(n17260), .B2(n17298), .ZN(
        P3_U2677) );
  INV_X1 U20196 ( .A(n17012), .ZN(n17020) );
  AOI21_X1 U20197 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n17260), .A(n17020), .ZN(
        n17014) );
  XNOR2_X1 U20198 ( .A(n17013), .B(n17016), .ZN(n17303) );
  OAI22_X1 U20199 ( .A1(n17015), .A2(n17014), .B1(n17260), .B2(n17303), .ZN(
        P3_U2678) );
  AOI21_X1 U20200 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n17260), .A(n17025), .ZN(
        n17019) );
  OAI21_X1 U20201 ( .B1(n17018), .B2(n17017), .A(n17016), .ZN(n17308) );
  OAI22_X1 U20202 ( .A1(n17020), .A2(n17019), .B1(n17260), .B2(n17308), .ZN(
        P3_U2679) );
  NOR3_X1 U20203 ( .A1(n17021), .A2(n17026), .A3(n17052), .ZN(n17039) );
  AOI21_X1 U20204 ( .B1(P3_EBX_REG_23__SCAN_IN), .B2(n17260), .A(n17039), .ZN(
        n17024) );
  XNOR2_X1 U20205 ( .A(n17023), .B(n17022), .ZN(n17313) );
  OAI22_X1 U20206 ( .A1(n17025), .A2(n17024), .B1(n17260), .B2(n17313), .ZN(
        P3_U2680) );
  NOR2_X1 U20207 ( .A1(n17026), .A2(n17052), .ZN(n17027) );
  AOI21_X1 U20208 ( .B1(P3_EBX_REG_22__SCAN_IN), .B2(n17260), .A(n17027), .ZN(
        n17038) );
  AOI22_X1 U20209 ( .A1(n17199), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n17153), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17031) );
  AOI22_X1 U20210 ( .A1(n9849), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17213), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n17030) );
  AOI22_X1 U20211 ( .A1(n9851), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17200), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n17029) );
  AOI22_X1 U20212 ( .A1(n17220), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17148), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n17028) );
  NAND4_X1 U20213 ( .A1(n17031), .A2(n17030), .A3(n17029), .A4(n17028), .ZN(
        n17037) );
  AOI22_X1 U20214 ( .A1(n17193), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17211), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n17035) );
  AOI22_X1 U20215 ( .A1(n17176), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17147), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n17034) );
  AOI22_X1 U20216 ( .A1(n17194), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n9837), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n17033) );
  AOI22_X1 U20217 ( .A1(n9838), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(n9839), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n17032) );
  NAND4_X1 U20218 ( .A1(n17035), .A2(n17034), .A3(n17033), .A4(n17032), .ZN(
        n17036) );
  NOR2_X1 U20219 ( .A1(n17037), .A2(n17036), .ZN(n17317) );
  OAI22_X1 U20220 ( .A1(n17039), .A2(n17038), .B1(n17317), .B2(n14394), .ZN(
        P3_U2681) );
  NOR2_X1 U20221 ( .A1(n17267), .A2(n17040), .ZN(n17063) );
  AOI22_X1 U20222 ( .A1(n9849), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(n9838), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n17050) );
  AOI22_X1 U20223 ( .A1(n17147), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n9839), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n17049) );
  AOI22_X1 U20224 ( .A1(n17194), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n9837), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n17041) );
  OAI21_X1 U20225 ( .B1(n10259), .B2(n17246), .A(n17041), .ZN(n17047) );
  AOI22_X1 U20226 ( .A1(n17193), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17112), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n17045) );
  AOI22_X1 U20227 ( .A1(n17200), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17177), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n17044) );
  AOI22_X1 U20228 ( .A1(n17199), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17211), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n17043) );
  AOI22_X1 U20229 ( .A1(n17192), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17148), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n17042) );
  NAND4_X1 U20230 ( .A1(n17045), .A2(n17044), .A3(n17043), .A4(n17042), .ZN(
        n17046) );
  AOI211_X1 U20231 ( .C1(n17219), .C2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A(
        n17047), .B(n17046), .ZN(n17048) );
  NAND3_X1 U20232 ( .A1(n17050), .A2(n17049), .A3(n17048), .ZN(n17322) );
  AOI22_X1 U20233 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n17063), .B1(n17267), 
        .B2(n17322), .ZN(n17051) );
  OAI21_X1 U20234 ( .B1(P3_EBX_REG_21__SCAN_IN), .B2(n17052), .A(n17051), .ZN(
        P3_U2682) );
  AOI22_X1 U20235 ( .A1(n17199), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n17193), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n17056) );
  AOI22_X1 U20236 ( .A1(n9851), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17212), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17055) );
  AOI22_X1 U20237 ( .A1(n9838), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n15785), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n17054) );
  AOI22_X1 U20238 ( .A1(n9849), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(n9837), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n17053) );
  NAND4_X1 U20239 ( .A1(n17056), .A2(n17055), .A3(n17054), .A4(n17053), .ZN(
        n17062) );
  AOI22_X1 U20240 ( .A1(n17176), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n9839), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n17060) );
  AOI22_X1 U20241 ( .A1(n17200), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17213), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n17059) );
  AOI22_X1 U20242 ( .A1(n17220), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17194), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n17058) );
  AOI22_X1 U20243 ( .A1(n17147), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17211), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n17057) );
  NAND4_X1 U20244 ( .A1(n17060), .A2(n17059), .A3(n17058), .A4(n17057), .ZN(
        n17061) );
  NOR2_X1 U20245 ( .A1(n17062), .A2(n17061), .ZN(n17330) );
  OAI21_X1 U20246 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(n17064), .A(n17063), .ZN(
        n17065) );
  OAI21_X1 U20247 ( .B1(n17330), .B2(n17260), .A(n17065), .ZN(P3_U2683) );
  AOI22_X1 U20248 ( .A1(n17212), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n17112), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n17069) );
  AOI22_X1 U20249 ( .A1(n17220), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17194), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n17068) );
  AOI22_X1 U20250 ( .A1(n17193), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n9837), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n17067) );
  AOI22_X1 U20251 ( .A1(n17199), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n15785), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n17066) );
  NAND4_X1 U20252 ( .A1(n17069), .A2(n17068), .A3(n17067), .A4(n17066), .ZN(
        n17075) );
  AOI22_X1 U20253 ( .A1(n9851), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17147), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n17073) );
  AOI22_X1 U20254 ( .A1(n17211), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17213), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n17072) );
  AOI22_X1 U20255 ( .A1(n17200), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n9838), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n17071) );
  AOI22_X1 U20256 ( .A1(n9849), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(n9839), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n17070) );
  NAND4_X1 U20257 ( .A1(n17073), .A2(n17072), .A3(n17071), .A4(n17070), .ZN(
        n17074) );
  NOR2_X1 U20258 ( .A1(n17075), .A2(n17074), .ZN(n17337) );
  OAI21_X1 U20259 ( .B1(P3_EBX_REG_19__SCAN_IN), .B2(n17077), .A(n17076), .ZN(
        n17078) );
  AOI22_X1 U20260 ( .A1(n17267), .A2(n17337), .B1(n17078), .B2(n14394), .ZN(
        P3_U2684) );
  NAND2_X1 U20261 ( .A1(n17260), .A2(n17090), .ZN(n17105) );
  AOI22_X1 U20262 ( .A1(n17211), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17213), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n17089) );
  AOI22_X1 U20263 ( .A1(n17199), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n9839), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n17088) );
  AOI22_X1 U20264 ( .A1(n17217), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n9838), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n17079) );
  OAI21_X1 U20265 ( .B1(n17080), .B2(n21013), .A(n17079), .ZN(n17086) );
  AOI22_X1 U20266 ( .A1(n17219), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n17177), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n17084) );
  AOI22_X1 U20267 ( .A1(n9849), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(n9837), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n17083) );
  AOI22_X1 U20268 ( .A1(n17193), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17112), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n17082) );
  AOI22_X1 U20269 ( .A1(n17147), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17148), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n17081) );
  NAND4_X1 U20270 ( .A1(n17084), .A2(n17083), .A3(n17082), .A4(n17081), .ZN(
        n17085) );
  AOI211_X1 U20271 ( .C1(n17153), .C2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A(
        n17086), .B(n17085), .ZN(n17087) );
  NAND3_X1 U20272 ( .A1(n17089), .A2(n17088), .A3(n17087), .ZN(n17338) );
  NOR3_X1 U20273 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n17356), .A3(n17090), .ZN(
        n17091) );
  AOI21_X1 U20274 ( .B1(n17267), .B2(n17338), .A(n17091), .ZN(n17092) );
  OAI21_X1 U20275 ( .B1(n17093), .B2(n17105), .A(n17092), .ZN(P3_U2685) );
  AOI22_X1 U20276 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n17220), .B1(
        n17147), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n17097) );
  AOI22_X1 U20277 ( .A1(n17200), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n17193), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n17096) );
  AOI22_X1 U20278 ( .A1(n17219), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_6__1__SCAN_IN), .B2(n17112), .ZN(n17095) );
  AOI22_X1 U20279 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n15785), .B1(
        n9837), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n17094) );
  NAND4_X1 U20280 ( .A1(n17097), .A2(n17096), .A3(n17095), .A4(n17094), .ZN(
        n17104) );
  AOI22_X1 U20281 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n17194), .B1(
        n9838), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n17102) );
  AOI22_X1 U20282 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n9839), .B1(
        P3_INSTQUEUE_REG_13__1__SCAN_IN), .B2(n17211), .ZN(n17101) );
  AOI22_X1 U20283 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n17098), .B1(
        n9849), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n17100) );
  AOI22_X1 U20284 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n17153), .B1(
        n17213), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n17099) );
  NAND4_X1 U20285 ( .A1(n17102), .A2(n17101), .A3(n17100), .A4(n17099), .ZN(
        n17103) );
  NOR2_X1 U20286 ( .A1(n17104), .A2(n17103), .ZN(n17348) );
  NOR2_X1 U20287 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n17120), .ZN(n17106) );
  OAI22_X1 U20288 ( .A1(n17348), .A2(n14394), .B1(n17106), .B2(n17105), .ZN(
        P3_U2686) );
  AOI22_X1 U20289 ( .A1(n18277), .A2(n17107), .B1(P3_EBX_REG_16__SCAN_IN), 
        .B2(n14394), .ZN(n17119) );
  AOI22_X1 U20290 ( .A1(n17199), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n9849), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n17111) );
  AOI22_X1 U20291 ( .A1(n17200), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17193), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n17110) );
  AOI22_X1 U20292 ( .A1(n9851), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n17213), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n17109) );
  AOI22_X1 U20293 ( .A1(n17212), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n15785), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n17108) );
  NAND4_X1 U20294 ( .A1(n17111), .A2(n17110), .A3(n17109), .A4(n17108), .ZN(
        n17118) );
  AOI22_X1 U20295 ( .A1(n9837), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n9838), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n17116) );
  AOI22_X1 U20296 ( .A1(n17220), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17112), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n17115) );
  AOI22_X1 U20297 ( .A1(n17217), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n9839), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n17114) );
  AOI22_X1 U20298 ( .A1(n17147), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17211), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n17113) );
  NAND4_X1 U20299 ( .A1(n17116), .A2(n17115), .A3(n17114), .A4(n17113), .ZN(
        n17117) );
  NOR2_X1 U20300 ( .A1(n17118), .A2(n17117), .ZN(n17355) );
  OAI22_X1 U20301 ( .A1(n17120), .A2(n17119), .B1(n17355), .B2(n14394), .ZN(
        P3_U2687) );
  AOI22_X1 U20302 ( .A1(n9849), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n17177), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n17124) );
  AOI22_X1 U20303 ( .A1(n17176), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17213), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n17123) );
  AOI22_X1 U20304 ( .A1(n9851), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n17212), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n17122) );
  AOI22_X1 U20305 ( .A1(n17200), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n15785), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n17121) );
  NAND4_X1 U20306 ( .A1(n17124), .A2(n17123), .A3(n17122), .A4(n17121), .ZN(
        n17130) );
  AOI22_X1 U20307 ( .A1(n17147), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n9838), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n17128) );
  AOI22_X1 U20308 ( .A1(n17193), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n9837), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n17127) );
  AOI22_X1 U20309 ( .A1(n17217), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n17211), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n17126) );
  AOI22_X1 U20310 ( .A1(n17199), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n9839), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n17125) );
  NAND4_X1 U20311 ( .A1(n17128), .A2(n17127), .A3(n17126), .A4(n17125), .ZN(
        n17129) );
  NOR2_X1 U20312 ( .A1(n17130), .A2(n17129), .ZN(n17362) );
  OAI21_X1 U20313 ( .B1(P3_EBX_REG_15__SCAN_IN), .B2(n17133), .A(n17131), .ZN(
        n17132) );
  AOI22_X1 U20314 ( .A1(n17267), .A2(n17362), .B1(n17132), .B2(n14394), .ZN(
        P3_U2688) );
  AOI21_X1 U20315 ( .B1(n20937), .B2(n17134), .A(n17133), .ZN(n17146) );
  AOI22_X1 U20316 ( .A1(n17199), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17147), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n17145) );
  AOI22_X1 U20317 ( .A1(n17211), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17192), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n17144) );
  AOI22_X1 U20318 ( .A1(n17176), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n9839), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n17135) );
  OAI21_X1 U20319 ( .B1(n17136), .B2(n21007), .A(n17135), .ZN(n17142) );
  AOI22_X1 U20320 ( .A1(n9849), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(n9838), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n17140) );
  AOI22_X1 U20321 ( .A1(n17212), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n17177), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n17139) );
  AOI22_X1 U20322 ( .A1(n9837), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n15785), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17138) );
  AOI22_X1 U20323 ( .A1(n9851), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n17200), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n17137) );
  NAND4_X1 U20324 ( .A1(n17140), .A2(n17139), .A3(n17138), .A4(n17137), .ZN(
        n17141) );
  AOI211_X1 U20325 ( .C1(n17193), .C2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A(
        n17142), .B(n17141), .ZN(n17143) );
  NAND3_X1 U20326 ( .A1(n17145), .A2(n17144), .A3(n17143), .ZN(n17364) );
  MUX2_X1 U20327 ( .A(n17146), .B(n17364), .S(n17267), .Z(P3_U2689) );
  AOI22_X1 U20328 ( .A1(n17199), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n17194), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n17152) );
  AOI22_X1 U20329 ( .A1(n17176), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n9839), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n17151) );
  AOI22_X1 U20330 ( .A1(n17147), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n9837), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n17150) );
  AOI22_X1 U20331 ( .A1(n17211), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17148), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17149) );
  NAND4_X1 U20332 ( .A1(n17152), .A2(n17151), .A3(n17150), .A4(n17149), .ZN(
        n17159) );
  AOI22_X1 U20333 ( .A1(n9851), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(n9849), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n17157) );
  AOI22_X1 U20334 ( .A1(n17200), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17193), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n17156) );
  AOI22_X1 U20335 ( .A1(n9838), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17192), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n17155) );
  AOI22_X1 U20336 ( .A1(n17153), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n17177), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n17154) );
  NAND4_X1 U20337 ( .A1(n17157), .A2(n17156), .A3(n17155), .A4(n17154), .ZN(
        n17158) );
  NOR2_X1 U20338 ( .A1(n17159), .A2(n17158), .ZN(n17372) );
  OAI21_X1 U20339 ( .B1(P3_EBX_REG_12__SCAN_IN), .B2(n17161), .A(n17160), .ZN(
        n17162) );
  OAI21_X1 U20340 ( .B1(n17372), .B2(n14394), .A(n17162), .ZN(P3_U2691) );
  AOI22_X1 U20341 ( .A1(n9851), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(n9839), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n17166) );
  AOI22_X1 U20342 ( .A1(n17220), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17211), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n17165) );
  AOI22_X1 U20343 ( .A1(n17199), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n9849), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n17164) );
  AOI22_X1 U20344 ( .A1(n17193), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n15785), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17163) );
  NAND4_X1 U20345 ( .A1(n17166), .A2(n17165), .A3(n17164), .A4(n17163), .ZN(
        n17172) );
  AOI22_X1 U20346 ( .A1(n17176), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n9838), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n17170) );
  AOI22_X1 U20347 ( .A1(n17212), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17147), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n17169) );
  AOI22_X1 U20348 ( .A1(n17200), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n9837), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n17168) );
  AOI22_X1 U20349 ( .A1(n17217), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17192), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n17167) );
  NAND4_X1 U20350 ( .A1(n17170), .A2(n17169), .A3(n17168), .A4(n17167), .ZN(
        n17171) );
  NOR2_X1 U20351 ( .A1(n17172), .A2(n17171), .ZN(n17377) );
  OAI21_X1 U20352 ( .B1(P3_EBX_REG_11__SCAN_IN), .B2(n17174), .A(n17173), .ZN(
        n17175) );
  AOI22_X1 U20353 ( .A1(n17267), .A2(n17377), .B1(n17175), .B2(n14394), .ZN(
        P3_U2692) );
  AOI22_X1 U20354 ( .A1(n17200), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n9837), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n17181) );
  AOI22_X1 U20355 ( .A1(n17176), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n17213), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n17180) );
  AOI22_X1 U20356 ( .A1(n9849), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n17177), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n17179) );
  AOI22_X1 U20357 ( .A1(n9851), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n15785), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17178) );
  NAND4_X1 U20358 ( .A1(n17181), .A2(n17180), .A3(n17179), .A4(n17178), .ZN(
        n17187) );
  AOI22_X1 U20359 ( .A1(n17212), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n17194), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n17185) );
  AOI22_X1 U20360 ( .A1(n17193), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n9838), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n17184) );
  AOI22_X1 U20361 ( .A1(n17199), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n17147), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n17183) );
  AOI22_X1 U20362 ( .A1(n17211), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n9839), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n17182) );
  NAND4_X1 U20363 ( .A1(n17185), .A2(n17184), .A3(n17183), .A4(n17182), .ZN(
        n17186) );
  NOR2_X1 U20364 ( .A1(n17187), .A2(n17186), .ZN(n17383) );
  INV_X1 U20365 ( .A(n17207), .ZN(n17188) );
  OAI33_X1 U20366 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n17356), .A3(n17207), 
        .B1(n17189), .B2(n17267), .B3(n17188), .ZN(n17190) );
  INV_X1 U20367 ( .A(n17190), .ZN(n17191) );
  OAI21_X1 U20368 ( .B1(n17383), .B2(n17260), .A(n17191), .ZN(P3_U2693) );
  AOI22_X1 U20369 ( .A1(n17219), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_13__1__SCAN_IN), .B2(n17192), .ZN(n17198) );
  AOI22_X1 U20370 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n17211), .B1(
        n17220), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n17197) );
  AOI22_X1 U20371 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n15785), .B1(
        n17193), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n17196) );
  AOI22_X1 U20372 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n17194), .B1(
        P3_INSTQUEUE_REG_4__1__SCAN_IN), .B2(n9838), .ZN(n17195) );
  NAND4_X1 U20373 ( .A1(n17198), .A2(n17197), .A3(n17196), .A4(n17195), .ZN(
        n17206) );
  AOI22_X1 U20374 ( .A1(n9849), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_7__1__SCAN_IN), .B2(n9839), .ZN(n17204) );
  AOI22_X1 U20375 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n17147), .B1(
        n17112), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n17203) );
  AOI22_X1 U20376 ( .A1(n17199), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_9__1__SCAN_IN), .B2(n9837), .ZN(n17202) );
  AOI22_X1 U20377 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n17153), .B1(
        n17200), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n17201) );
  NAND4_X1 U20378 ( .A1(n17204), .A2(n17203), .A3(n17202), .A4(n17201), .ZN(
        n17205) );
  NOR2_X1 U20379 ( .A1(n17206), .A2(n17205), .ZN(n17385) );
  OAI211_X1 U20380 ( .C1(P3_EBX_REG_9__SCAN_IN), .C2(n17208), .A(n17207), .B(
        n14394), .ZN(n17209) );
  OAI21_X1 U20381 ( .B1(n17385), .B2(n17260), .A(n17209), .ZN(P3_U2694) );
  NAND2_X1 U20382 ( .A1(n17260), .A2(n17210), .ZN(n17236) );
  AOI22_X1 U20383 ( .A1(n17212), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17211), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n17229) );
  AOI22_X1 U20384 ( .A1(n17193), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n9838), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n17228) );
  AOI22_X1 U20385 ( .A1(n9849), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n17213), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n17214) );
  OAI21_X1 U20386 ( .B1(n17215), .B2(n21111), .A(n17214), .ZN(n17226) );
  AOI22_X1 U20387 ( .A1(n17217), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17216), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n17224) );
  AOI22_X1 U20388 ( .A1(n9832), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(n9837), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n17223) );
  AOI22_X1 U20389 ( .A1(n9851), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n17112), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n17222) );
  AOI22_X1 U20390 ( .A1(n17220), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n9839), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n17221) );
  NAND4_X1 U20391 ( .A1(n17224), .A2(n17223), .A3(n17222), .A4(n17221), .ZN(
        n17225) );
  AOI211_X1 U20392 ( .C1(n17098), .C2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A(
        n17226), .B(n17225), .ZN(n17227) );
  NAND3_X1 U20393 ( .A1(n17229), .A2(n17228), .A3(n17227), .ZN(n17389) );
  NOR3_X1 U20394 ( .A1(n17356), .A2(n17230), .A3(n17247), .ZN(n17240) );
  NOR3_X1 U20395 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n17237), .A3(n17239), .ZN(
        n17231) );
  AOI22_X1 U20396 ( .A1(n17267), .A2(n17389), .B1(n17240), .B2(n17231), .ZN(
        n17232) );
  OAI21_X1 U20397 ( .B1(n17233), .B2(n17236), .A(n17232), .ZN(P3_U2695) );
  NOR2_X1 U20398 ( .A1(P3_EBX_REG_7__SCAN_IN), .A2(n17239), .ZN(n17234) );
  AOI22_X1 U20399 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n17267), .B1(
        n17240), .B2(n17234), .ZN(n17235) );
  OAI21_X1 U20400 ( .B1(n17237), .B2(n17236), .A(n17235), .ZN(P3_U2696) );
  INV_X1 U20401 ( .A(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17242) );
  NOR2_X1 U20402 ( .A1(n17267), .A2(n17238), .ZN(n17243) );
  AOI22_X1 U20403 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n17243), .B1(n17240), .B2(
        n17239), .ZN(n17241) );
  OAI21_X1 U20404 ( .B1(n17242), .B2(n14394), .A(n17241), .ZN(P3_U2697) );
  INV_X1 U20405 ( .A(n17247), .ZN(n17244) );
  OAI21_X1 U20406 ( .B1(P3_EBX_REG_5__SCAN_IN), .B2(n17244), .A(n17243), .ZN(
        n17245) );
  OAI21_X1 U20407 ( .B1(n17260), .B2(n17246), .A(n17245), .ZN(P3_U2698) );
  NAND2_X1 U20408 ( .A1(n17248), .A2(n17263), .ZN(n17258) );
  NOR2_X1 U20409 ( .A1(n17252), .A2(n17258), .ZN(n17251) );
  AOI21_X1 U20410 ( .B1(P3_EBX_REG_4__SCAN_IN), .B2(n17260), .A(n17251), .ZN(
        n17250) );
  INV_X1 U20411 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17249) );
  OAI22_X1 U20412 ( .A1(n17244), .A2(n17250), .B1(n17249), .B2(n14394), .ZN(
        P3_U2699) );
  INV_X1 U20413 ( .A(n17251), .ZN(n17254) );
  OAI21_X1 U20414 ( .B1(n17252), .B2(n17267), .A(n17258), .ZN(n17253) );
  AOI22_X1 U20415 ( .A1(n17254), .A2(n17253), .B1(
        P3_INSTQUEUE_REG_0__3__SCAN_IN), .B2(n17267), .ZN(n17255) );
  INV_X1 U20416 ( .A(n17255), .ZN(P3_U2700) );
  OAI221_X1 U20417 ( .B1(n17257), .B2(n17266), .C1(n18277), .C2(n17266), .A(
        n17256), .ZN(n17259) );
  OAI211_X1 U20418 ( .C1(n17260), .C2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A(
        n17259), .B(n17258), .ZN(n17261) );
  INV_X1 U20419 ( .A(n17261), .ZN(P3_U2701) );
  INV_X1 U20420 ( .A(n17262), .ZN(n17264) );
  AOI222_X1 U20421 ( .A1(n17264), .A2(n17263), .B1(P3_EBX_REG_1__SCAN_IN), 
        .B2(n17266), .C1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .C2(n17267), .ZN(
        n17265) );
  INV_X1 U20422 ( .A(n17265), .ZN(P3_U2702) );
  AOI22_X1 U20423 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n17267), .B1(
        P3_EBX_REG_0__SCAN_IN), .B2(n17266), .ZN(n17268) );
  OAI21_X1 U20424 ( .B1(P3_EBX_REG_0__SCAN_IN), .B2(n17269), .A(n17268), .ZN(
        P3_U2703) );
  INV_X1 U20425 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n17434) );
  INV_X1 U20426 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n17438) );
  INV_X1 U20427 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n17444) );
  INV_X1 U20428 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n17448) );
  INV_X1 U20429 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n17450) );
  INV_X1 U20430 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n17540) );
  INV_X1 U20431 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n17474) );
  INV_X1 U20432 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n17512) );
  NAND4_X1 U20433 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(P3_EAX_REG_0__SCAN_IN), 
        .A3(P3_EAX_REG_4__SCAN_IN), .A4(P3_EAX_REG_3__SCAN_IN), .ZN(n17270) );
  NOR2_X1 U20434 ( .A1(n17512), .A2(n17270), .ZN(n17400) );
  NAND2_X1 U20435 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n17400), .ZN(n17396) );
  NAND3_X1 U20436 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(P3_EAX_REG_11__SCAN_IN), 
        .A3(P3_EAX_REG_10__SCAN_IN), .ZN(n17363) );
  INV_X1 U20437 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n17468) );
  INV_X1 U20438 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n17520) );
  NAND3_X1 U20439 ( .A1(P3_EAX_REG_14__SCAN_IN), .A2(P3_EAX_REG_13__SCAN_IN), 
        .A3(n17271), .ZN(n17357) );
  NAND2_X1 U20440 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(P3_EAX_REG_17__SCAN_IN), 
        .ZN(n17327) );
  NAND2_X1 U20441 ( .A1(P3_EAX_REG_24__SCAN_IN), .A2(n17305), .ZN(n17304) );
  NAND2_X1 U20442 ( .A1(P3_EAX_REG_29__SCAN_IN), .A2(n17286), .ZN(n17282) );
  NAND2_X1 U20443 ( .A1(n17277), .A2(P3_EAX_REG_30__SCAN_IN), .ZN(n17276) );
  NOR2_X2 U20444 ( .A1(n18271), .A2(n17413), .ZN(n17349) );
  OAI22_X1 U20445 ( .A1(P3_EAX_REG_30__SCAN_IN), .A2(n17404), .B1(n17375), 
        .B2(n17277), .ZN(n17273) );
  AOI22_X1 U20446 ( .A1(BUF2_REG_31__SCAN_IN), .A2(n17349), .B1(
        P3_EAX_REG_31__SCAN_IN), .B2(n17273), .ZN(n17274) );
  OAI21_X1 U20447 ( .B1(P3_EAX_REG_31__SCAN_IN), .B2(n17276), .A(n17274), .ZN(
        P3_U2704) );
  NOR2_X2 U20448 ( .A1(n17275), .A2(n17413), .ZN(n17350) );
  AOI22_X1 U20449 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17350), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n17349), .ZN(n17279) );
  OAI211_X1 U20450 ( .C1(n17277), .C2(P3_EAX_REG_30__SCAN_IN), .A(n17413), .B(
        n17276), .ZN(n17278) );
  OAI211_X1 U20451 ( .C1(n17280), .C2(n17415), .A(n17279), .B(n17278), .ZN(
        P3_U2705) );
  INV_X1 U20452 ( .A(n17349), .ZN(n17328) );
  AOI22_X1 U20453 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17350), .B1(n17281), .B2(
        n17422), .ZN(n17284) );
  OAI211_X1 U20454 ( .C1(n17286), .C2(P3_EAX_REG_29__SCAN_IN), .A(n17413), .B(
        n17282), .ZN(n17283) );
  OAI211_X1 U20455 ( .C1(n17328), .C2(n18266), .A(n17284), .B(n17283), .ZN(
        P3_U2706) );
  INV_X1 U20456 ( .A(n17350), .ZN(n17343) );
  AOI22_X1 U20457 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n17349), .B1(n17285), .B2(
        n17422), .ZN(n17289) );
  AOI211_X1 U20458 ( .C1(n17434), .C2(n17291), .A(n17286), .B(n17375), .ZN(
        n17287) );
  INV_X1 U20459 ( .A(n17287), .ZN(n17288) );
  OAI211_X1 U20460 ( .C1(n17343), .C2(n17528), .A(n17289), .B(n17288), .ZN(
        P3_U2707) );
  AOI22_X1 U20461 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17350), .B1(n17290), .B2(
        n17422), .ZN(n17293) );
  OAI211_X1 U20462 ( .C1(n9915), .C2(P3_EAX_REG_27__SCAN_IN), .A(n17413), .B(
        n17291), .ZN(n17292) );
  OAI211_X1 U20463 ( .C1(n17328), .C2(n17294), .A(n17293), .B(n17292), .ZN(
        P3_U2708) );
  AOI22_X1 U20464 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17350), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n17349), .ZN(n17297) );
  AOI211_X1 U20465 ( .C1(n17438), .C2(n17299), .A(n9915), .B(n17375), .ZN(
        n17295) );
  INV_X1 U20466 ( .A(n17295), .ZN(n17296) );
  OAI211_X1 U20467 ( .C1(n17298), .C2(n17415), .A(n17297), .B(n17296), .ZN(
        P3_U2709) );
  AOI22_X1 U20468 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17350), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n17349), .ZN(n17302) );
  OAI211_X1 U20469 ( .C1(n17300), .C2(P3_EAX_REG_25__SCAN_IN), .A(n17413), .B(
        n17299), .ZN(n17301) );
  OAI211_X1 U20470 ( .C1(n17303), .C2(n17415), .A(n17302), .B(n17301), .ZN(
        P3_U2710) );
  AOI22_X1 U20471 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17350), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n17349), .ZN(n17307) );
  OAI211_X1 U20472 ( .C1(n17305), .C2(P3_EAX_REG_24__SCAN_IN), .A(n17413), .B(
        n17304), .ZN(n17306) );
  OAI211_X1 U20473 ( .C1(n17308), .C2(n17415), .A(n17307), .B(n17306), .ZN(
        P3_U2711) );
  AOI22_X1 U20474 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17350), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n17349), .ZN(n17312) );
  OAI211_X1 U20475 ( .C1(P3_EAX_REG_23__SCAN_IN), .C2(n17310), .A(n17413), .B(
        n17309), .ZN(n17311) );
  OAI211_X1 U20476 ( .C1(n17313), .C2(n17415), .A(n17312), .B(n17311), .ZN(
        P3_U2712) );
  NOR2_X1 U20477 ( .A1(n17356), .A2(n17314), .ZN(n17320) );
  NAND2_X1 U20478 ( .A1(n18277), .A2(n17315), .ZN(n17326) );
  NAND2_X1 U20479 ( .A1(n17413), .A2(n17326), .ZN(n17333) );
  OAI21_X1 U20480 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n17404), .A(n17333), .ZN(
        n17319) );
  OAI22_X1 U20481 ( .A1(n17317), .A2(n17415), .B1(n17316), .B2(n17328), .ZN(
        n17318) );
  AOI221_X1 U20482 ( .B1(n17320), .B2(n17444), .C1(n17319), .C2(
        P3_EAX_REG_22__SCAN_IN), .A(n17318), .ZN(n17321) );
  OAI21_X1 U20483 ( .B1(n18270), .B2(n17343), .A(n17321), .ZN(P3_U2713) );
  AOI22_X1 U20484 ( .A1(BUF2_REG_21__SCAN_IN), .A2(n17349), .B1(n17422), .B2(
        n17322), .ZN(n17325) );
  INV_X1 U20485 ( .A(n17333), .ZN(n17323) );
  AOI22_X1 U20486 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17350), .B1(
        P3_EAX_REG_21__SCAN_IN), .B2(n17323), .ZN(n17324) );
  OAI211_X1 U20487 ( .C1(P3_EAX_REG_21__SCAN_IN), .C2(n17326), .A(n17325), .B(
        n17324), .ZN(P3_U2714) );
  NOR3_X1 U20488 ( .A1(n17356), .A2(n17351), .A3(n17327), .ZN(n17339) );
  NAND2_X1 U20489 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(n17339), .ZN(n17334) );
  OAI22_X1 U20490 ( .A1(n17330), .A2(n17415), .B1(n17329), .B2(n17328), .ZN(
        n17331) );
  AOI21_X1 U20491 ( .B1(BUF2_REG_4__SCAN_IN), .B2(n17350), .A(n17331), .ZN(
        n17332) );
  OAI221_X1 U20492 ( .B1(P3_EAX_REG_20__SCAN_IN), .B2(n17334), .C1(n17448), 
        .C2(n17333), .A(n17332), .ZN(P3_U2715) );
  AOI22_X1 U20493 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17350), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n17349), .ZN(n17336) );
  OAI211_X1 U20494 ( .C1(n17339), .C2(P3_EAX_REG_19__SCAN_IN), .A(n17413), .B(
        n17334), .ZN(n17335) );
  OAI211_X1 U20495 ( .C1(n17337), .C2(n17415), .A(n17336), .B(n17335), .ZN(
        P3_U2716) );
  INV_X1 U20496 ( .A(BUF2_REG_2__SCAN_IN), .ZN(n18253) );
  AOI22_X1 U20497 ( .A1(BUF2_REG_18__SCAN_IN), .A2(n17349), .B1(n17422), .B2(
        n17338), .ZN(n17342) );
  INV_X1 U20498 ( .A(P3_EAX_REG_18__SCAN_IN), .ZN(n17452) );
  INV_X1 U20499 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n17494) );
  OR2_X1 U20500 ( .A1(n17494), .A2(n17351), .ZN(n17344) );
  AOI211_X1 U20501 ( .C1(n17452), .C2(n17344), .A(n17339), .B(n17375), .ZN(
        n17340) );
  INV_X1 U20502 ( .A(n17340), .ZN(n17341) );
  OAI211_X1 U20503 ( .C1(n17343), .C2(n18253), .A(n17342), .B(n17341), .ZN(
        P3_U2717) );
  AOI22_X1 U20504 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17350), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n17349), .ZN(n17347) );
  INV_X1 U20505 ( .A(n17351), .ZN(n17345) );
  OAI211_X1 U20506 ( .C1(n17345), .C2(P3_EAX_REG_17__SCAN_IN), .A(n17413), .B(
        n17344), .ZN(n17346) );
  OAI211_X1 U20507 ( .C1(n17348), .C2(n17415), .A(n17347), .B(n17346), .ZN(
        P3_U2718) );
  AOI22_X1 U20508 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17350), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n17349), .ZN(n17354) );
  OAI211_X1 U20509 ( .C1(P3_EAX_REG_16__SCAN_IN), .C2(n17352), .A(n17413), .B(
        n17351), .ZN(n17353) );
  OAI211_X1 U20510 ( .C1(n17355), .C2(n17415), .A(n17354), .B(n17353), .ZN(
        P3_U2719) );
  NOR2_X1 U20511 ( .A1(n17356), .A2(n17357), .ZN(n17359) );
  NAND2_X1 U20512 ( .A1(n17413), .A2(n17357), .ZN(n17366) );
  INV_X1 U20513 ( .A(n17366), .ZN(n17358) );
  MUX2_X1 U20514 ( .A(n17359), .B(n17358), .S(P3_EAX_REG_15__SCAN_IN), .Z(
        n17360) );
  AOI21_X1 U20515 ( .B1(BUF2_REG_15__SCAN_IN), .B2(n17423), .A(n17360), .ZN(
        n17361) );
  OAI21_X1 U20516 ( .B1(n17362), .B2(n17415), .A(n17361), .ZN(P3_U2720) );
  NAND3_X1 U20517 ( .A1(n18277), .A2(P3_EAX_REG_7__SCAN_IN), .A3(n17399), .ZN(
        n17392) );
  NOR2_X1 U20518 ( .A1(n17520), .A2(n17392), .ZN(n17384) );
  NAND2_X1 U20519 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(n17384), .ZN(n17371) );
  NOR2_X1 U20520 ( .A1(n17363), .A2(n17371), .ZN(n17374) );
  NAND2_X1 U20521 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(n17374), .ZN(n17367) );
  INV_X1 U20522 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n17535) );
  AOI22_X1 U20523 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17423), .B1(n17422), .B2(
        n17364), .ZN(n17365) );
  OAI221_X1 U20524 ( .B1(P3_EAX_REG_14__SCAN_IN), .B2(n17367), .C1(n17535), 
        .C2(n17366), .A(n17365), .ZN(P3_U2721) );
  INV_X1 U20525 ( .A(n17367), .ZN(n17370) );
  AOI21_X1 U20526 ( .B1(P3_EAX_REG_13__SCAN_IN), .B2(n17413), .A(n17374), .ZN(
        n17369) );
  OAI222_X1 U20527 ( .A1(n17418), .A2(n17533), .B1(n17370), .B2(n17369), .C1(
        n17415), .C2(n17368), .ZN(P3_U2722) );
  INV_X1 U20528 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n17464) );
  INV_X1 U20529 ( .A(n17371), .ZN(n17387) );
  NAND2_X1 U20530 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n17387), .ZN(n17380) );
  NOR2_X1 U20531 ( .A1(n17464), .A2(n17380), .ZN(n17379) );
  AOI21_X1 U20532 ( .B1(P3_EAX_REG_12__SCAN_IN), .B2(n17413), .A(n17379), .ZN(
        n17373) );
  OAI222_X1 U20533 ( .A1(n17418), .A2(n17528), .B1(n17374), .B2(n17373), .C1(
        n17415), .C2(n17372), .ZN(P3_U2723) );
  OAI21_X1 U20534 ( .B1(n17464), .B2(n17375), .A(n17380), .ZN(n17376) );
  INV_X1 U20535 ( .A(n17376), .ZN(n17378) );
  OAI222_X1 U20536 ( .A1(n17418), .A2(n17526), .B1(n17379), .B2(n17378), .C1(
        n17415), .C2(n17377), .ZN(P3_U2724) );
  NAND2_X1 U20537 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17423), .ZN(n17382) );
  OAI211_X1 U20538 ( .C1(P3_EAX_REG_10__SCAN_IN), .C2(n17387), .A(n17413), .B(
        n17380), .ZN(n17381) );
  OAI211_X1 U20539 ( .C1(n17383), .C2(n17415), .A(n17382), .B(n17381), .ZN(
        P3_U2725) );
  AOI21_X1 U20540 ( .B1(P3_EAX_REG_9__SCAN_IN), .B2(n17413), .A(n17384), .ZN(
        n17386) );
  OAI222_X1 U20541 ( .A1(n17418), .A2(n17522), .B1(n17387), .B2(n17386), .C1(
        n17415), .C2(n17385), .ZN(P3_U2726) );
  NAND2_X1 U20542 ( .A1(n17413), .A2(n17388), .ZN(n17391) );
  AOI22_X1 U20543 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17423), .B1(n17422), .B2(
        n17389), .ZN(n17390) );
  OAI221_X1 U20544 ( .B1(P3_EAX_REG_8__SCAN_IN), .B2(n17392), .C1(n17520), 
        .C2(n17391), .A(n17390), .ZN(P3_U2727) );
  INV_X1 U20545 ( .A(n17392), .ZN(n17395) );
  AOI22_X1 U20546 ( .A1(n18277), .A2(n17399), .B1(P3_EAX_REG_7__SCAN_IN), .B2(
        n17413), .ZN(n17394) );
  OAI222_X1 U20547 ( .A1(n17418), .A2(n18274), .B1(n17395), .B2(n17394), .C1(
        n17415), .C2(n17393), .ZN(P3_U2728) );
  NOR2_X1 U20548 ( .A1(n17396), .A2(n17404), .ZN(n17402) );
  AOI21_X1 U20549 ( .B1(P3_EAX_REG_6__SCAN_IN), .B2(n17413), .A(n17402), .ZN(
        n17398) );
  OAI222_X1 U20550 ( .A1(n17418), .A2(n18270), .B1(n17399), .B2(n17398), .C1(
        n17415), .C2(n17397), .ZN(P3_U2729) );
  INV_X1 U20551 ( .A(n17404), .ZN(n17419) );
  AND2_X1 U20552 ( .A1(n17400), .A2(n17419), .ZN(n17407) );
  AOI21_X1 U20553 ( .B1(P3_EAX_REG_5__SCAN_IN), .B2(n17413), .A(n17407), .ZN(
        n17403) );
  OAI222_X1 U20554 ( .A1(n17418), .A2(n18265), .B1(n17403), .B2(n17402), .C1(
        n17415), .C2(n17401), .ZN(P3_U2730) );
  INV_X1 U20555 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n17480) );
  NOR3_X1 U20556 ( .A1(n17512), .A2(n17488), .A3(n17404), .ZN(n17412) );
  NAND2_X1 U20557 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(n17412), .ZN(n17408) );
  NOR2_X1 U20558 ( .A1(n17480), .A2(n17408), .ZN(n17411) );
  AOI21_X1 U20559 ( .B1(P3_EAX_REG_4__SCAN_IN), .B2(n17413), .A(n17411), .ZN(
        n17406) );
  OAI222_X1 U20560 ( .A1(n18261), .A2(n17418), .B1(n17407), .B2(n17406), .C1(
        n17415), .C2(n17405), .ZN(P3_U2731) );
  INV_X1 U20561 ( .A(n17408), .ZN(n17417) );
  AOI21_X1 U20562 ( .B1(P3_EAX_REG_3__SCAN_IN), .B2(n17413), .A(n17417), .ZN(
        n17410) );
  OAI222_X1 U20563 ( .A1(n18257), .A2(n17418), .B1(n17411), .B2(n17410), .C1(
        n17415), .C2(n17409), .ZN(P3_U2732) );
  AOI21_X1 U20564 ( .B1(P3_EAX_REG_2__SCAN_IN), .B2(n17413), .A(n17412), .ZN(
        n17416) );
  OAI222_X1 U20565 ( .A1(n18253), .A2(n17418), .B1(n17417), .B2(n17416), .C1(
        n17415), .C2(n17414), .ZN(P3_U2733) );
  NAND2_X1 U20566 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(n17419), .ZN(n17426) );
  AOI21_X1 U20567 ( .B1(n18277), .B2(n17488), .A(n17420), .ZN(n17425) );
  AOI22_X1 U20568 ( .A1(n17423), .A2(BUF2_REG_1__SCAN_IN), .B1(n17422), .B2(
        n17421), .ZN(n17424) );
  OAI221_X1 U20569 ( .B1(P3_EAX_REG_1__SCAN_IN), .B2(n17426), .C1(n17512), 
        .C2(n17425), .A(n17424), .ZN(P3_U2734) );
  AND2_X1 U20570 ( .A1(n17470), .A2(P3_DATAO_REG_31__SCAN_IN), .ZN(P3_U2736)
         );
  INV_X1 U20571 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n17509) );
  NAND2_X1 U20572 ( .A1(n17429), .A2(n17428), .ZN(n17455) );
  AOI22_X1 U20573 ( .A1(n18881), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(n17484), 
        .B2(P3_DATAO_REG_30__SCAN_IN), .ZN(n17430) );
  OAI21_X1 U20574 ( .B1(n17509), .B2(n17455), .A(n17430), .ZN(P3_U2737) );
  INV_X1 U20575 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n17432) );
  AOI22_X1 U20576 ( .A1(n18881), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n17470), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n17431) );
  OAI21_X1 U20577 ( .B1(n17432), .B2(n17455), .A(n17431), .ZN(P3_U2738) );
  AOI22_X1 U20578 ( .A1(n18881), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n17470), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n17433) );
  OAI21_X1 U20579 ( .B1(n17434), .B2(n17455), .A(n17433), .ZN(P3_U2739) );
  INV_X1 U20580 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n17436) );
  AOI22_X1 U20581 ( .A1(n18881), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n17470), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n17435) );
  OAI21_X1 U20582 ( .B1(n17436), .B2(n17455), .A(n17435), .ZN(P3_U2740) );
  AOI22_X1 U20583 ( .A1(n18881), .A2(P3_UWORD_REG_10__SCAN_IN), .B1(n17470), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n17437) );
  OAI21_X1 U20584 ( .B1(n17438), .B2(n17455), .A(n17437), .ZN(P3_U2741) );
  AOI22_X1 U20585 ( .A1(n18881), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n17470), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n17439) );
  OAI21_X1 U20586 ( .B1(n10012), .B2(n17455), .A(n17439), .ZN(P3_U2742) );
  INV_X1 U20587 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n17502) );
  AOI22_X1 U20588 ( .A1(n18881), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n17470), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n17440) );
  OAI21_X1 U20589 ( .B1(n17502), .B2(n17455), .A(n17440), .ZN(P3_U2743) );
  INV_X1 U20590 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n17442) );
  AOI22_X1 U20591 ( .A1(n17485), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n17484), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n17441) );
  OAI21_X1 U20592 ( .B1(n17442), .B2(n17455), .A(n17441), .ZN(P3_U2744) );
  AOI22_X1 U20593 ( .A1(n17485), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n17484), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n17443) );
  OAI21_X1 U20594 ( .B1(n17444), .B2(n17455), .A(n17443), .ZN(P3_U2745) );
  INV_X1 U20595 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n17446) );
  AOI22_X1 U20596 ( .A1(n17485), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n17484), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n17445) );
  OAI21_X1 U20597 ( .B1(n17446), .B2(n17455), .A(n17445), .ZN(P3_U2746) );
  AOI22_X1 U20598 ( .A1(n17485), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n17484), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n17447) );
  OAI21_X1 U20599 ( .B1(n17448), .B2(n17455), .A(n17447), .ZN(P3_U2747) );
  AOI22_X1 U20600 ( .A1(n17485), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n17484), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n17449) );
  OAI21_X1 U20601 ( .B1(n17450), .B2(n17455), .A(n17449), .ZN(P3_U2748) );
  AOI22_X1 U20602 ( .A1(n17485), .A2(P3_UWORD_REG_2__SCAN_IN), .B1(n17484), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n17451) );
  OAI21_X1 U20603 ( .B1(n17452), .B2(n17455), .A(n17451), .ZN(P3_U2749) );
  AOI22_X1 U20604 ( .A1(n17485), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n17484), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n17453) );
  OAI21_X1 U20605 ( .B1(n17494), .B2(n17455), .A(n17453), .ZN(P3_U2750) );
  INV_X1 U20606 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n17456) );
  AOI22_X1 U20607 ( .A1(n17485), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n17484), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n17454) );
  OAI21_X1 U20608 ( .B1(n17456), .B2(n17455), .A(n17454), .ZN(P3_U2751) );
  AOI22_X1 U20609 ( .A1(n17485), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n17484), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n17457) );
  OAI21_X1 U20610 ( .B1(n17540), .B2(n17487), .A(n17457), .ZN(P3_U2752) );
  AOI22_X1 U20611 ( .A1(n17485), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n17484), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n17458) );
  OAI21_X1 U20612 ( .B1(n17535), .B2(n17487), .A(n17458), .ZN(P3_U2753) );
  INV_X1 U20613 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n17460) );
  AOI22_X1 U20614 ( .A1(n17485), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n17484), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n17459) );
  OAI21_X1 U20615 ( .B1(n17460), .B2(n17487), .A(n17459), .ZN(P3_U2754) );
  INV_X1 U20616 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n17462) );
  AOI22_X1 U20617 ( .A1(n17485), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n17484), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n17461) );
  OAI21_X1 U20618 ( .B1(n17462), .B2(n17487), .A(n17461), .ZN(P3_U2755) );
  AOI22_X1 U20619 ( .A1(n17485), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n17470), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n17463) );
  OAI21_X1 U20620 ( .B1(n17464), .B2(n17487), .A(n17463), .ZN(P3_U2756) );
  INV_X1 U20621 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n17466) );
  AOI22_X1 U20622 ( .A1(n17485), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n17470), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n17465) );
  OAI21_X1 U20623 ( .B1(n17466), .B2(n17487), .A(n17465), .ZN(P3_U2757) );
  AOI22_X1 U20624 ( .A1(n17485), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n17470), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n17467) );
  OAI21_X1 U20625 ( .B1(n17468), .B2(n17487), .A(n17467), .ZN(P3_U2758) );
  AOI22_X1 U20626 ( .A1(n17485), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n17484), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n17469) );
  OAI21_X1 U20627 ( .B1(n17520), .B2(n17487), .A(n17469), .ZN(P3_U2759) );
  INV_X1 U20628 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n17472) );
  AOI22_X1 U20629 ( .A1(n17485), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n17470), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n17471) );
  OAI21_X1 U20630 ( .B1(n17472), .B2(n17487), .A(n17471), .ZN(P3_U2760) );
  AOI22_X1 U20631 ( .A1(n17485), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n17484), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n17473) );
  OAI21_X1 U20632 ( .B1(n17474), .B2(n17487), .A(n17473), .ZN(P3_U2761) );
  INV_X1 U20633 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n17476) );
  AOI22_X1 U20634 ( .A1(n17485), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n17484), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n17475) );
  OAI21_X1 U20635 ( .B1(n17476), .B2(n17487), .A(n17475), .ZN(P3_U2762) );
  INV_X1 U20636 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n17478) );
  AOI22_X1 U20637 ( .A1(n17485), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n17484), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n17477) );
  OAI21_X1 U20638 ( .B1(n17478), .B2(n17487), .A(n17477), .ZN(P3_U2763) );
  AOI22_X1 U20639 ( .A1(n17485), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n17484), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n17479) );
  OAI21_X1 U20640 ( .B1(n17480), .B2(n17487), .A(n17479), .ZN(P3_U2764) );
  INV_X1 U20641 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n17482) );
  AOI22_X1 U20642 ( .A1(n17485), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n17484), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n17481) );
  OAI21_X1 U20643 ( .B1(n17482), .B2(n17487), .A(n17481), .ZN(P3_U2765) );
  AOI22_X1 U20644 ( .A1(n17485), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n17484), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n17483) );
  OAI21_X1 U20645 ( .B1(n17512), .B2(n17487), .A(n17483), .ZN(P3_U2766) );
  AOI22_X1 U20646 ( .A1(n17485), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n17484), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n17486) );
  OAI21_X1 U20647 ( .B1(n17488), .B2(n17487), .A(n17486), .ZN(P3_U2767) );
  OAI211_X1 U20648 ( .C1(n18880), .C2(n18886), .A(n17490), .B(n17489), .ZN(
        n17536) );
  NAND2_X1 U20649 ( .A1(n18886), .A2(n17490), .ZN(n18735) );
  AOI22_X1 U20650 ( .A1(P3_EAX_REG_16__SCAN_IN), .A2(n17530), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n17529), .ZN(n17492) );
  OAI21_X1 U20651 ( .B1(n21157), .B2(n17532), .A(n17492), .ZN(P3_U2768) );
  AOI22_X1 U20652 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17537), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n17529), .ZN(n17493) );
  OAI21_X1 U20653 ( .B1(n17494), .B2(n17539), .A(n17493), .ZN(P3_U2769) );
  AOI22_X1 U20654 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n17530), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n17529), .ZN(n17495) );
  OAI21_X1 U20655 ( .B1(n18253), .B2(n17532), .A(n17495), .ZN(P3_U2770) );
  AOI22_X1 U20656 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(n17530), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n17529), .ZN(n17496) );
  OAI21_X1 U20657 ( .B1(n18257), .B2(n17532), .A(n17496), .ZN(P3_U2771) );
  AOI22_X1 U20658 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n17530), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n17529), .ZN(n17497) );
  OAI21_X1 U20659 ( .B1(n18261), .B2(n17532), .A(n17497), .ZN(P3_U2772) );
  AOI22_X1 U20660 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(n17530), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n17529), .ZN(n17498) );
  OAI21_X1 U20661 ( .B1(n18265), .B2(n17532), .A(n17498), .ZN(P3_U2773) );
  AOI22_X1 U20662 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(n17530), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n17529), .ZN(n17499) );
  OAI21_X1 U20663 ( .B1(n18270), .B2(n17532), .A(n17499), .ZN(P3_U2774) );
  AOI22_X1 U20664 ( .A1(P3_EAX_REG_23__SCAN_IN), .A2(n17530), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n17529), .ZN(n17500) );
  OAI21_X1 U20665 ( .B1(n18274), .B2(n17532), .A(n17500), .ZN(P3_U2775) );
  AOI22_X1 U20666 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17537), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n17529), .ZN(n17501) );
  OAI21_X1 U20667 ( .B1(n17502), .B2(n17539), .A(n17501), .ZN(P3_U2776) );
  AOI22_X1 U20668 ( .A1(P3_EAX_REG_25__SCAN_IN), .A2(n17530), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n17529), .ZN(n17503) );
  OAI21_X1 U20669 ( .B1(n17522), .B2(n17532), .A(n17503), .ZN(P3_U2777) );
  AOI22_X1 U20670 ( .A1(P3_EAX_REG_26__SCAN_IN), .A2(n17530), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n17529), .ZN(n17504) );
  OAI21_X1 U20671 ( .B1(n17524), .B2(n17532), .A(n17504), .ZN(P3_U2778) );
  AOI22_X1 U20672 ( .A1(P3_EAX_REG_27__SCAN_IN), .A2(n17530), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n17529), .ZN(n17505) );
  OAI21_X1 U20673 ( .B1(n17526), .B2(n17532), .A(n17505), .ZN(P3_U2779) );
  AOI22_X1 U20674 ( .A1(P3_EAX_REG_28__SCAN_IN), .A2(n17530), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n17529), .ZN(n17506) );
  OAI21_X1 U20675 ( .B1(n17528), .B2(n17532), .A(n17506), .ZN(P3_U2780) );
  AOI22_X1 U20676 ( .A1(P3_EAX_REG_29__SCAN_IN), .A2(n17530), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n17529), .ZN(n17507) );
  OAI21_X1 U20677 ( .B1(n17533), .B2(n17532), .A(n17507), .ZN(P3_U2781) );
  AOI22_X1 U20678 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17537), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n17529), .ZN(n17508) );
  OAI21_X1 U20679 ( .B1(n17509), .B2(n17539), .A(n17508), .ZN(P3_U2782) );
  AOI22_X1 U20680 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(n17530), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n17529), .ZN(n17510) );
  OAI21_X1 U20681 ( .B1(n21157), .B2(n17532), .A(n17510), .ZN(P3_U2783) );
  AOI22_X1 U20682 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17537), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n17529), .ZN(n17511) );
  OAI21_X1 U20683 ( .B1(n17512), .B2(n17539), .A(n17511), .ZN(P3_U2784) );
  AOI22_X1 U20684 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(n17530), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n17529), .ZN(n17513) );
  OAI21_X1 U20685 ( .B1(n18253), .B2(n17532), .A(n17513), .ZN(P3_U2785) );
  AOI22_X1 U20686 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n17530), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n17529), .ZN(n17514) );
  OAI21_X1 U20687 ( .B1(n18257), .B2(n17532), .A(n17514), .ZN(P3_U2786) );
  AOI22_X1 U20688 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(n17530), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n17536), .ZN(n17515) );
  OAI21_X1 U20689 ( .B1(n18261), .B2(n17532), .A(n17515), .ZN(P3_U2787) );
  AOI22_X1 U20690 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n17530), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n17536), .ZN(n17516) );
  OAI21_X1 U20691 ( .B1(n18265), .B2(n17532), .A(n17516), .ZN(P3_U2788) );
  AOI22_X1 U20692 ( .A1(P3_EAX_REG_6__SCAN_IN), .A2(n17530), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n17536), .ZN(n17517) );
  OAI21_X1 U20693 ( .B1(n18270), .B2(n17532), .A(n17517), .ZN(P3_U2789) );
  AOI22_X1 U20694 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(n17530), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n17536), .ZN(n17518) );
  OAI21_X1 U20695 ( .B1(n18274), .B2(n17532), .A(n17518), .ZN(P3_U2790) );
  AOI22_X1 U20696 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17537), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n17536), .ZN(n17519) );
  OAI21_X1 U20697 ( .B1(n17520), .B2(n17539), .A(n17519), .ZN(P3_U2791) );
  AOI22_X1 U20698 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(n17530), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n17536), .ZN(n17521) );
  OAI21_X1 U20699 ( .B1(n17522), .B2(n17532), .A(n17521), .ZN(P3_U2792) );
  AOI22_X1 U20700 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n17530), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n17536), .ZN(n17523) );
  OAI21_X1 U20701 ( .B1(n17524), .B2(n17532), .A(n17523), .ZN(P3_U2793) );
  AOI22_X1 U20702 ( .A1(P3_EAX_REG_11__SCAN_IN), .A2(n17530), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n17536), .ZN(n17525) );
  OAI21_X1 U20703 ( .B1(n17526), .B2(n17532), .A(n17525), .ZN(P3_U2794) );
  AOI22_X1 U20704 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n17530), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n17529), .ZN(n17527) );
  OAI21_X1 U20705 ( .B1(n17528), .B2(n17532), .A(n17527), .ZN(P3_U2795) );
  AOI22_X1 U20706 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(n17530), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n17529), .ZN(n17531) );
  OAI21_X1 U20707 ( .B1(n17533), .B2(n17532), .A(n17531), .ZN(P3_U2796) );
  AOI22_X1 U20708 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17537), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n17536), .ZN(n17534) );
  OAI21_X1 U20709 ( .B1(n17535), .B2(n17539), .A(n17534), .ZN(P3_U2797) );
  AOI22_X1 U20710 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n17537), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n17536), .ZN(n17538) );
  OAI21_X1 U20711 ( .B1(n17540), .B2(n17539), .A(n17538), .ZN(P3_U2798) );
  OAI21_X1 U20712 ( .B1(n17546), .B2(n17867), .A(n17910), .ZN(n17541) );
  AOI21_X1 U20713 ( .B1(n17630), .B2(n17542), .A(n17541), .ZN(n17572) );
  OAI21_X1 U20714 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n17697), .A(
        n17572), .ZN(n17557) );
  AOI211_X1 U20715 ( .C1(n17545), .C2(n17544), .A(n17543), .B(n17808), .ZN(
        n17552) );
  AND2_X1 U20716 ( .A1(n17546), .A2(n17712), .ZN(n17564) );
  NAND2_X1 U20717 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n17547) );
  OAI211_X1 U20718 ( .C1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A(n17564), .B(n17547), .ZN(n17549) );
  OAI211_X1 U20719 ( .C1(n17750), .C2(n17550), .A(n17549), .B(n17548), .ZN(
        n17551) );
  AOI211_X1 U20720 ( .C1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .C2(n17557), .A(
        n17552), .B(n17551), .ZN(n17556) );
  NAND2_X1 U20721 ( .A1(n17914), .A2(n17822), .ZN(n17658) );
  AOI22_X1 U20722 ( .A1(n17894), .A2(n17917), .B1(n17598), .B2(n17916), .ZN(
        n17577) );
  NAND2_X1 U20723 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n17577), .ZN(
        n17565) );
  NAND3_X1 U20724 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17658), .A3(
        n17565), .ZN(n17555) );
  NAND3_X1 U20725 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n17566), .A3(
        n17553), .ZN(n17554) );
  NAND3_X1 U20726 ( .A1(n17556), .A2(n17555), .A3(n17554), .ZN(P3_U2802) );
  AOI22_X1 U20727 ( .A1(n17767), .A2(n17558), .B1(
        P3_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n17557), .ZN(n17569) );
  INV_X1 U20728 ( .A(n17559), .ZN(n17560) );
  NAND2_X1 U20729 ( .A1(n17561), .A2(n17560), .ZN(n17562) );
  XNOR2_X1 U20730 ( .A(n17562), .B(n17757), .ZN(n17926) );
  AOI22_X1 U20731 ( .A1(n17819), .A2(n17926), .B1(n17564), .B2(n17563), .ZN(
        n17568) );
  OAI21_X1 U20732 ( .B1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n17566), .A(
        n17565), .ZN(n17567) );
  NAND2_X1 U20733 ( .A1(n18231), .A2(P3_REIP_REG_27__SCAN_IN), .ZN(n17927) );
  NAND4_X1 U20734 ( .A1(n17569), .A2(n17568), .A3(n17567), .A4(n17927), .ZN(
        P3_U2803) );
  AOI21_X1 U20735 ( .B1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n17571), .A(
        n17570), .ZN(n17939) );
  NOR2_X1 U20736 ( .A1(n18218), .A2(n18813), .ZN(n17936) );
  AOI221_X1 U20737 ( .B1(n18343), .B2(n17574), .C1(n17573), .C2(n17574), .A(
        n17572), .ZN(n17582) );
  INV_X1 U20738 ( .A(n17697), .ZN(n17575) );
  AOI21_X1 U20739 ( .B1(n17750), .B2(n17697), .A(n17576), .ZN(n17581) );
  NAND2_X1 U20740 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n17918), .ZN(
        n17931) );
  NOR2_X1 U20741 ( .A1(n17721), .A2(n17931), .ZN(n17579) );
  INV_X1 U20742 ( .A(n17577), .ZN(n17578) );
  MUX2_X1 U20743 ( .A(n17579), .B(n17578), .S(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .Z(n17580) );
  NOR4_X1 U20744 ( .A1(n17936), .A2(n17582), .A3(n17581), .A4(n17580), .ZN(
        n17583) );
  OAI21_X1 U20745 ( .B1(n17939), .B2(n17808), .A(n17583), .ZN(P3_U2804) );
  INV_X1 U20746 ( .A(n18048), .ZN(n17585) );
  NAND2_X1 U20747 ( .A1(n18048), .A2(n17608), .ZN(n17956) );
  OAI21_X1 U20748 ( .B1(n17611), .B2(n17956), .A(n17594), .ZN(n17584) );
  OAI21_X1 U20749 ( .B1(n17931), .B2(n17585), .A(n17584), .ZN(n17953) );
  INV_X1 U20750 ( .A(n17910), .ZN(n17876) );
  NOR2_X1 U20751 ( .A1(n17599), .A2(n18343), .ZN(n17625) );
  AOI211_X1 U20752 ( .C1(n17630), .C2(n17586), .A(n17876), .B(n17625), .ZN(
        n17619) );
  OAI21_X1 U20753 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n17697), .A(
        n17619), .ZN(n17602) );
  NOR2_X1 U20754 ( .A1(n18218), .A2(n18811), .ZN(n17948) );
  AND2_X1 U20755 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n17589) );
  OAI211_X1 U20756 ( .C1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A(n17599), .B(n17712), .ZN(n17588) );
  OAI22_X1 U20757 ( .A1(n17589), .A2(n17588), .B1(n17750), .B2(n17587), .ZN(
        n17590) );
  AOI211_X1 U20758 ( .C1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .C2(n17602), .A(
        n17948), .B(n17590), .ZN(n17597) );
  NAND2_X1 U20759 ( .A1(n17918), .A2(n18058), .ZN(n17591) );
  XNOR2_X1 U20760 ( .A(n17591), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n17950) );
  AOI21_X1 U20761 ( .B1(n17593), .B2(n17757), .A(n17592), .ZN(n17595) );
  XNOR2_X1 U20762 ( .A(n17595), .B(n17594), .ZN(n17949) );
  AOI22_X1 U20763 ( .A1(n17894), .A2(n17950), .B1(n17819), .B2(n17949), .ZN(
        n17596) );
  OAI211_X1 U20764 ( .C1(n17822), .C2(n17953), .A(n17597), .B(n17596), .ZN(
        P3_U2805) );
  NAND2_X1 U20765 ( .A1(n18058), .A2(n17608), .ZN(n17957) );
  AOI22_X1 U20766 ( .A1(n17894), .A2(n17957), .B1(n17598), .B2(n17956), .ZN(
        n17620) );
  AND2_X1 U20767 ( .A1(n17599), .A2(n17712), .ZN(n17604) );
  OAI22_X1 U20768 ( .A1(n18218), .A2(n18809), .B1(n17750), .B2(n17600), .ZN(
        n17601) );
  AOI221_X1 U20769 ( .B1(n17604), .B2(n17603), .C1(n17602), .C2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A(n17601), .ZN(n17610) );
  AOI21_X1 U20770 ( .B1(n17606), .B2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n17605), .ZN(n17607) );
  INV_X1 U20771 ( .A(n17607), .ZN(n17955) );
  AND2_X1 U20772 ( .A1(n17611), .A2(n17608), .ZN(n17954) );
  AOI22_X1 U20773 ( .A1(n17819), .A2(n17955), .B1(n17690), .B2(n17954), .ZN(
        n17609) );
  OAI211_X1 U20774 ( .C1(n17620), .C2(n17611), .A(n17610), .B(n17609), .ZN(
        P3_U2806) );
  AOI22_X1 U20775 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n17757), .B1(
        n17612), .B2(n17635), .ZN(n17613) );
  NAND2_X1 U20776 ( .A1(n17659), .A2(n17613), .ZN(n17614) );
  XNOR2_X1 U20777 ( .A(n17614), .B(n20983), .ZN(n17970) );
  INV_X1 U20778 ( .A(n17615), .ZN(n17626) );
  NAND2_X1 U20779 ( .A1(n18231), .A2(P3_REIP_REG_23__SCAN_IN), .ZN(n17969) );
  OAI21_X1 U20780 ( .B1(n17767), .B2(n17575), .A(n17616), .ZN(n17617) );
  OAI211_X1 U20781 ( .C1(n17619), .C2(n17618), .A(n17969), .B(n17617), .ZN(
        n17624) );
  NOR2_X1 U20782 ( .A1(n17964), .A2(n17721), .ZN(n17622) );
  INV_X1 U20783 ( .A(n17620), .ZN(n17621) );
  MUX2_X1 U20784 ( .A(n17622), .B(n17621), .S(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .Z(n17623) );
  AOI211_X1 U20785 ( .C1(n17626), .C2(n17625), .A(n17624), .B(n17623), .ZN(
        n17627) );
  OAI21_X1 U20786 ( .B1(n17808), .B2(n17970), .A(n17627), .ZN(P3_U2807) );
  OAI21_X1 U20787 ( .B1(n17631), .B2(n17867), .A(n17910), .ZN(n17628) );
  AOI21_X1 U20788 ( .B1(n17630), .B2(n17629), .A(n17628), .ZN(n17661) );
  OAI21_X1 U20789 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n17697), .A(
        n17661), .ZN(n17649) );
  INV_X1 U20790 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n17633) );
  NAND2_X1 U20791 ( .A1(n17631), .A2(n17712), .ZN(n17647) );
  AOI221_X1 U20792 ( .B1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .C1(n17633), .C2(n17632), .A(
        n17647), .ZN(n17634) );
  NOR2_X1 U20793 ( .A1(n18218), .A2(n18806), .ZN(n17971) );
  AOI211_X1 U20794 ( .C1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .C2(n17649), .A(
        n17634), .B(n17971), .ZN(n17644) );
  INV_X1 U20795 ( .A(n17635), .ZN(n17636) );
  OAI21_X1 U20796 ( .B1(n17637), .B2(n17636), .A(n17659), .ZN(n17638) );
  XNOR2_X1 U20797 ( .A(n17638), .B(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n17972) );
  NOR2_X1 U20798 ( .A1(n17639), .A2(n17721), .ZN(n17641) );
  OAI22_X1 U20799 ( .A1(n18058), .A2(n17914), .B1(n18048), .B2(n17822), .ZN(
        n17703) );
  AOI21_X1 U20800 ( .B1(n17639), .B2(n17658), .A(n17703), .ZN(n17657) );
  INV_X1 U20801 ( .A(n17657), .ZN(n17640) );
  MUX2_X1 U20802 ( .A(n17641), .B(n17640), .S(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .Z(n17642) );
  AOI21_X1 U20803 ( .B1(n17819), .B2(n17972), .A(n17642), .ZN(n17643) );
  OAI211_X1 U20804 ( .C1(n17750), .C2(n17645), .A(n17644), .B(n17643), .ZN(
        P3_U2808) );
  NOR2_X1 U20805 ( .A1(n18218), .A2(n18804), .ZN(n17993) );
  OAI22_X1 U20806 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n17647), .B1(
        n17750), .B2(n17646), .ZN(n17648) );
  AOI211_X1 U20807 ( .C1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .C2(n17649), .A(
        n17993), .B(n17648), .ZN(n17656) );
  AND3_X1 U20808 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17818), .A3(
        n17650), .ZN(n17676) );
  AOI22_X1 U20809 ( .A1(n17653), .A2(n17676), .B1(n17687), .B2(n17651), .ZN(
        n17652) );
  XNOR2_X1 U20810 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .B(n17652), .ZN(
        n17994) );
  INV_X1 U20811 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n18031) );
  NOR2_X1 U20812 ( .A1(n18018), .A2(n18031), .ZN(n17986) );
  NAND3_X1 U20813 ( .A1(n17989), .A2(n17653), .A3(n17986), .ZN(n17996) );
  INV_X1 U20814 ( .A(n17996), .ZN(n17654) );
  AOI22_X1 U20815 ( .A1(n17819), .A2(n17994), .B1(n17690), .B2(n17654), .ZN(
        n17655) );
  OAI211_X1 U20816 ( .C1(n17657), .C2(n17989), .A(n17656), .B(n17655), .ZN(
        P3_U2809) );
  NAND2_X1 U20817 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17986), .ZN(
        n18000) );
  AOI21_X1 U20818 ( .B1(n17658), .B2(n18000), .A(n17703), .ZN(n17680) );
  INV_X1 U20819 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n21160) );
  NOR2_X1 U20820 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n18000), .ZN(
        n18003) );
  OAI221_X1 U20821 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n17685), 
        .C1(n18015), .C2(n17676), .A(n17659), .ZN(n17660) );
  XOR2_X1 U20822 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .B(n17660), .Z(
        n18007) );
  AOI221_X1 U20823 ( .B1(n18343), .B2(n17663), .C1(n17662), .C2(n17663), .A(
        n17661), .ZN(n17664) );
  AOI221_X1 U20824 ( .B1(n17767), .B2(n17665), .C1(n17575), .C2(n17665), .A(
        n17664), .ZN(n17666) );
  NAND2_X1 U20825 ( .A1(n18231), .A2(P3_REIP_REG_20__SCAN_IN), .ZN(n18005) );
  OAI211_X1 U20826 ( .C1(n17808), .C2(n18007), .A(n17666), .B(n18005), .ZN(
        n17667) );
  AOI21_X1 U20827 ( .B1(n17690), .B2(n18003), .A(n17667), .ZN(n17668) );
  OAI21_X1 U20828 ( .B1(n17680), .B2(n21160), .A(n17668), .ZN(P3_U2810) );
  INV_X1 U20829 ( .A(n17671), .ZN(n17669) );
  OAI21_X1 U20830 ( .B1(n17876), .B2(n17669), .A(n17905), .ZN(n17691) );
  OAI21_X1 U20831 ( .B1(n17670), .B2(n17909), .A(n17691), .ZN(n17684) );
  NOR2_X1 U20832 ( .A1(n18218), .A2(n18800), .ZN(n18011) );
  NAND2_X1 U20833 ( .A1(n17671), .A2(n17712), .ZN(n17682) );
  OAI21_X1 U20834 ( .B1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(n17672), .ZN(n17673) );
  OAI22_X1 U20835 ( .A1(n17750), .A2(n17674), .B1(n17682), .B2(n17673), .ZN(
        n17675) );
  AOI211_X1 U20836 ( .C1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .C2(n17684), .A(
        n18011), .B(n17675), .ZN(n17679) );
  AOI21_X1 U20837 ( .B1(n17685), .B2(n17687), .A(n17676), .ZN(n17677) );
  XNOR2_X1 U20838 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B(n17677), .ZN(
        n18010) );
  AND2_X1 U20839 ( .A1(n18015), .A2(n17986), .ZN(n18008) );
  AOI22_X1 U20840 ( .A1(n17819), .A2(n18010), .B1(n17690), .B2(n18008), .ZN(
        n17678) );
  OAI211_X1 U20841 ( .C1(n17680), .C2(n18015), .A(n17679), .B(n17678), .ZN(
        P3_U2811) );
  AOI21_X1 U20842 ( .B1(n17690), .B2(n18018), .A(n17703), .ZN(n17702) );
  NOR2_X1 U20843 ( .A1(n18218), .A2(n18798), .ZN(n18027) );
  OAI22_X1 U20844 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n17682), .B1(
        n17750), .B2(n17681), .ZN(n17683) );
  AOI211_X1 U20845 ( .C1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(n17684), .A(
        n18027), .B(n17683), .ZN(n17689) );
  AOI21_X1 U20846 ( .B1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n17818), .A(
        n17685), .ZN(n17686) );
  XOR2_X1 U20847 ( .A(n17687), .B(n17686), .Z(n18026) );
  NOR2_X1 U20848 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n18018), .ZN(
        n18025) );
  AOI22_X1 U20849 ( .A1(n17819), .A2(n18026), .B1(n17690), .B2(n18025), .ZN(
        n17688) );
  OAI211_X1 U20850 ( .C1(n17702), .C2(n18031), .A(n17689), .B(n17688), .ZN(
        P3_U2812) );
  AOI21_X1 U20851 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n17690), .A(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n17701) );
  AOI221_X1 U20852 ( .B1(n18343), .B2(n17693), .C1(n17692), .C2(n17693), .A(
        n17691), .ZN(n17694) );
  AOI21_X1 U20853 ( .B1(P3_REIP_REG_17__SCAN_IN), .B2(n18231), .A(n17694), 
        .ZN(n17700) );
  OAI21_X1 U20854 ( .B1(n17696), .B2(n21008), .A(n17695), .ZN(n18032) );
  AOI22_X1 U20855 ( .A1(n17819), .A2(n18032), .B1(n17698), .B2(n17903), .ZN(
        n17699) );
  OAI211_X1 U20856 ( .C1(n17702), .C2(n17701), .A(n17700), .B(n17699), .ZN(
        P3_U2813) );
  INV_X1 U20857 ( .A(n17703), .ZN(n17720) );
  AOI21_X1 U20858 ( .B1(n17818), .B2(n17705), .A(n17704), .ZN(n17706) );
  XNOR2_X1 U20859 ( .A(n17706), .B(n18043), .ZN(n18045) );
  INV_X1 U20860 ( .A(n17707), .ZN(n17708) );
  AOI21_X1 U20861 ( .B1(n17709), .B2(n17708), .A(n17876), .ZN(n17743) );
  OAI21_X1 U20862 ( .B1(n17710), .B2(n17909), .A(n17743), .ZN(n17724) );
  AOI22_X1 U20863 ( .A1(n17767), .A2(n17711), .B1(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n17724), .ZN(n17717) );
  INV_X1 U20864 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n17725) );
  INV_X1 U20865 ( .A(n17733), .ZN(n17713) );
  NAND2_X1 U20866 ( .A1(n17713), .A2(n17712), .ZN(n17764) );
  NOR2_X1 U20867 ( .A1(n17714), .A2(n17764), .ZN(n17726) );
  OAI221_X1 U20868 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .C1(n17725), .C2(n17715), .A(
        n17726), .ZN(n17716) );
  OAI211_X1 U20869 ( .C1(n20933), .C2(n18218), .A(n17717), .B(n17716), .ZN(
        n17718) );
  AOI21_X1 U20870 ( .B1(n17819), .B2(n18045), .A(n17718), .ZN(n17719) );
  OAI221_X1 U20871 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n17721), 
        .C1(n18043), .C2(n17720), .A(n17719), .ZN(P3_U2814) );
  INV_X1 U20872 ( .A(n18103), .ZN(n18023) );
  AOI21_X1 U20873 ( .B1(n18041), .B2(n18023), .A(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n18057) );
  OR2_X1 U20874 ( .A1(n17914), .A2(n18058), .ZN(n17732) );
  OAI22_X1 U20875 ( .A1(n18218), .A2(n18793), .B1(n17750), .B2(n17722), .ZN(
        n17723) );
  AOI221_X1 U20876 ( .B1(n17726), .B2(n17725), .C1(n17724), .C2(
        P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A(n17723), .ZN(n17731) );
  NAND4_X1 U20877 ( .A1(n17775), .A2(n17774), .A3(n18144), .A4(n13132), .ZN(
        n17768) );
  NOR2_X1 U20878 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n17768), .ZN(
        n17736) );
  INV_X1 U20879 ( .A(n18070), .ZN(n17755) );
  NOR3_X1 U20880 ( .A1(n17755), .A2(n17757), .A3(n17754), .ZN(n17727) );
  INV_X1 U20881 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n18067) );
  NAND2_X1 U20882 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n18067), .ZN(
        n18092) );
  OAI221_X1 U20883 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n17736), 
        .C1(n18074), .C2(n17727), .A(n18092), .ZN(n17728) );
  XNOR2_X1 U20884 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B(n17728), .ZN(
        n18062) );
  NOR2_X1 U20885 ( .A1(n18048), .A2(n17822), .ZN(n17729) );
  NAND2_X1 U20886 ( .A1(n18059), .A2(n17738), .ZN(n18055) );
  AOI22_X1 U20887 ( .A1(n17819), .A2(n18062), .B1(n17729), .B2(n18055), .ZN(
        n17730) );
  OAI211_X1 U20888 ( .C1(n18057), .C2(n17732), .A(n17731), .B(n17730), .ZN(
        P3_U2815) );
  NOR2_X1 U20889 ( .A1(n18343), .A2(n17733), .ZN(n17781) );
  AOI21_X1 U20890 ( .B1(n17744), .B2(n17781), .A(
        P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n17742) );
  AOI22_X1 U20891 ( .A1(n18231), .A2(P3_REIP_REG_14__SCAN_IN), .B1(n17734), 
        .B2(n17903), .ZN(n17741) );
  AND2_X1 U20892 ( .A1(n18023), .A2(n18041), .ZN(n17735) );
  AOI221_X1 U20893 ( .B1(n18103), .B2(n18074), .C1(n18068), .C2(n18074), .A(
        n17735), .ZN(n18065) );
  NAND2_X1 U20894 ( .A1(n17818), .A2(n9870), .ZN(n17798) );
  INV_X1 U20895 ( .A(n17798), .ZN(n17777) );
  INV_X1 U20896 ( .A(n18068), .ZN(n18051) );
  AOI22_X1 U20897 ( .A1(n17777), .A2(n18051), .B1(n17736), .B2(n18100), .ZN(
        n17737) );
  XNOR2_X1 U20898 ( .A(n17737), .B(n18074), .ZN(n18076) );
  OAI221_X1 U20899 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n18051), 
        .C1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n18022), .A(n17738), .ZN(
        n18075) );
  OAI22_X1 U20900 ( .A1(n18076), .A2(n17808), .B1(n17822), .B2(n18075), .ZN(
        n17739) );
  AOI21_X1 U20901 ( .B1(n17894), .B2(n18065), .A(n17739), .ZN(n17740) );
  OAI211_X1 U20902 ( .C1(n17743), .C2(n17742), .A(n17741), .B(n17740), .ZN(
        P3_U2816) );
  INV_X1 U20903 ( .A(n18108), .ZN(n18081) );
  NAND2_X1 U20904 ( .A1(n18081), .A2(n17805), .ZN(n17773) );
  AOI211_X1 U20905 ( .C1(n17763), .C2(n17751), .A(n17744), .B(n17764), .ZN(
        n17753) );
  OAI21_X1 U20906 ( .B1(n17745), .B2(n17867), .A(n17909), .ZN(n17747) );
  OAI21_X1 U20907 ( .B1(n17746), .B2(n17867), .A(n17910), .ZN(n17826) );
  AOI21_X1 U20908 ( .B1(n17748), .B2(n17747), .A(n17826), .ZN(n17762) );
  OAI22_X1 U20909 ( .A1(n17762), .A2(n17751), .B1(n17750), .B2(n17749), .ZN(
        n17752) );
  AOI211_X1 U20910 ( .C1(P3_REIP_REG_13__SCAN_IN), .C2(n18231), .A(n17753), 
        .B(n17752), .ZN(n17761) );
  NOR2_X1 U20911 ( .A1(n18103), .A2(n17755), .ZN(n18086) );
  NOR2_X1 U20912 ( .A1(n17755), .A2(n18101), .ZN(n18084) );
  OAI22_X1 U20913 ( .A1(n18086), .A2(n17914), .B1(n18084), .B2(n17822), .ZN(
        n17770) );
  NOR2_X1 U20914 ( .A1(n17755), .A2(n17754), .ZN(n17758) );
  OAI221_X1 U20915 ( .B1(n17758), .B2(n18100), .C1(n17758), .C2(n17757), .A(
        n17756), .ZN(n17759) );
  XNOR2_X1 U20916 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B(n17759), .ZN(
        n18082) );
  AOI22_X1 U20917 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n17770), .B1(
        n17819), .B2(n18082), .ZN(n17760) );
  OAI211_X1 U20918 ( .C1(n18092), .C2(n17773), .A(n17761), .B(n17760), .ZN(
        P3_U2817) );
  NAND2_X1 U20919 ( .A1(n18231), .A2(P3_REIP_REG_12__SCAN_IN), .ZN(n18098) );
  OAI221_X1 U20920 ( .B1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n17764), .C1(
        n17763), .C2(n17762), .A(n18098), .ZN(n17765) );
  AOI21_X1 U20921 ( .B1(n17767), .B2(n17766), .A(n17765), .ZN(n17772) );
  OAI21_X1 U20922 ( .B1(n18108), .B2(n17798), .A(n17768), .ZN(n17769) );
  XNOR2_X1 U20923 ( .A(n17769), .B(n18100), .ZN(n18097) );
  AOI22_X1 U20924 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n17770), .B1(
        n17819), .B2(n18097), .ZN(n17771) );
  OAI211_X1 U20925 ( .C1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .C2(n17773), .A(
        n17772), .B(n17771), .ZN(P3_U2818) );
  INV_X1 U20926 ( .A(n17774), .ZN(n17793) );
  NAND2_X1 U20927 ( .A1(n17775), .A2(n18144), .ZN(n17797) );
  NOR2_X1 U20928 ( .A1(n17793), .A2(n17797), .ZN(n17776) );
  AOI21_X1 U20929 ( .B1(n17777), .B2(n17784), .A(n17776), .ZN(n17778) );
  XNOR2_X1 U20930 ( .A(n17778), .B(n13132), .ZN(n18115) );
  INV_X1 U20931 ( .A(n17784), .ZN(n18107) );
  NOR2_X1 U20932 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n18107), .ZN(
        n18113) );
  NOR2_X1 U20933 ( .A1(n18218), .A2(n18786), .ZN(n18111) );
  INV_X2 U20934 ( .A(n18343), .ZN(n18626) );
  NAND3_X1 U20935 ( .A1(n17853), .A2(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A3(
        n18626), .ZN(n17825) );
  NOR2_X1 U20936 ( .A1(n17810), .A2(n17825), .ZN(n17801) );
  NAND2_X1 U20937 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n17801), .ZN(
        n17800) );
  NOR2_X1 U20938 ( .A1(n17789), .A2(n17800), .ZN(n17788) );
  AOI21_X1 U20939 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n17905), .A(
        n17788), .ZN(n17780) );
  OAI22_X1 U20940 ( .A1(n17781), .A2(n17780), .B1(n17897), .B2(n17779), .ZN(
        n17782) );
  AOI211_X1 U20941 ( .C1(n18113), .C2(n17805), .A(n18111), .B(n17782), .ZN(
        n17786) );
  NOR2_X1 U20942 ( .A1(n17784), .A2(n17783), .ZN(n17794) );
  OAI22_X1 U20943 ( .A1(n18022), .A2(n17822), .B1(n17914), .B2(n18023), .ZN(
        n17806) );
  OAI21_X1 U20944 ( .B1(n17794), .B2(n17806), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n17785) );
  OAI211_X1 U20945 ( .C1(n18115), .C2(n17808), .A(n17786), .B(n17785), .ZN(
        P3_U2819) );
  AOI22_X1 U20946 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n17798), .B1(
        n17797), .B2(n18127), .ZN(n17787) );
  XNOR2_X1 U20947 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B(n17787), .ZN(
        n18124) );
  INV_X1 U20948 ( .A(n17905), .ZN(n17850) );
  AOI211_X1 U20949 ( .C1(n17800), .C2(n17789), .A(n17850), .B(n17788), .ZN(
        n17791) );
  NOR2_X1 U20950 ( .A1(n18218), .A2(n18784), .ZN(n17790) );
  AOI211_X1 U20951 ( .C1(n17792), .C2(n17903), .A(n17791), .B(n17790), .ZN(
        n17796) );
  AOI22_X1 U20952 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n17806), .B1(
        n17794), .B2(n17793), .ZN(n17795) );
  OAI211_X1 U20953 ( .C1(n18124), .C2(n17808), .A(n17796), .B(n17795), .ZN(
        P3_U2820) );
  NAND2_X1 U20954 ( .A1(n17798), .A2(n17797), .ZN(n17799) );
  XNOR2_X1 U20955 ( .A(n17799), .B(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n18125) );
  OAI211_X1 U20956 ( .C1(n17801), .C2(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A(
        n17905), .B(n17800), .ZN(n17802) );
  NAND2_X1 U20957 ( .A1(n18231), .A2(P3_REIP_REG_9__SCAN_IN), .ZN(n18134) );
  OAI211_X1 U20958 ( .C1(n17897), .C2(n17803), .A(n17802), .B(n18134), .ZN(
        n17804) );
  AOI221_X1 U20959 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n17806), .C1(
        n18127), .C2(n17805), .A(n17804), .ZN(n17807) );
  OAI21_X1 U20960 ( .B1(n18125), .B2(n17808), .A(n17807), .ZN(P3_U2821) );
  INV_X1 U20961 ( .A(n17809), .ZN(n18152) );
  OAI211_X1 U20962 ( .C1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .C2(n17811), .A(
        n18626), .B(n17810), .ZN(n17812) );
  NAND2_X1 U20963 ( .A1(n18231), .A2(P3_REIP_REG_8__SCAN_IN), .ZN(n18141) );
  OAI211_X1 U20964 ( .C1(n17897), .C2(n17813), .A(n17812), .B(n18141), .ZN(
        n17814) );
  AOI21_X1 U20965 ( .B1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n17826), .A(
        n17814), .ZN(n17821) );
  AOI21_X1 U20966 ( .B1(n17816), .B2(n18144), .A(n17815), .ZN(n18148) );
  OAI21_X1 U20967 ( .B1(n17818), .B2(n17809), .A(n17817), .ZN(n18146) );
  AOI22_X1 U20968 ( .A1(n17894), .A2(n18148), .B1(n17819), .B2(n18146), .ZN(
        n17820) );
  OAI211_X1 U20969 ( .C1(n17822), .C2(n18152), .A(n17821), .B(n17820), .ZN(
        P3_U2822) );
  OAI21_X1 U20970 ( .B1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n17824), .A(
        n17823), .ZN(n18160) );
  INV_X1 U20971 ( .A(n17825), .ZN(n17842) );
  INV_X1 U20972 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n18778) );
  NOR2_X1 U20973 ( .A1(n18218), .A2(n18778), .ZN(n18158) );
  AOI221_X1 U20974 ( .B1(n17842), .B2(n17827), .C1(n17826), .C2(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A(n18158), .ZN(n17834) );
  NAND2_X1 U20975 ( .A1(n17829), .A2(n17828), .ZN(n17830) );
  XOR2_X1 U20976 ( .A(n17830), .B(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .Z(
        n18154) );
  INV_X1 U20977 ( .A(n18154), .ZN(n17832) );
  AOI22_X1 U20978 ( .A1(n17894), .A2(n17832), .B1(n17831), .B2(n17903), .ZN(
        n17833) );
  OAI211_X1 U20979 ( .C1(n17913), .C2(n18160), .A(n17834), .B(n17833), .ZN(
        P3_U2823) );
  OAI21_X1 U20980 ( .B1(n17837), .B2(n17836), .A(n17835), .ZN(n18168) );
  AOI21_X1 U20981 ( .B1(n18163), .B2(n17839), .A(n17838), .ZN(n18166) );
  AOI22_X1 U20982 ( .A1(n18626), .A2(n17853), .B1(
        P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n17905), .ZN(n17841) );
  OAI22_X1 U20983 ( .A1(n17842), .A2(n17841), .B1(n17897), .B2(n17840), .ZN(
        n17843) );
  AOI21_X1 U20984 ( .B1(n17894), .B2(n18166), .A(n17843), .ZN(n17844) );
  NAND2_X1 U20985 ( .A1(n18231), .A2(P3_REIP_REG_6__SCAN_IN), .ZN(n18162) );
  OAI211_X1 U20986 ( .C1(n17913), .C2(n18168), .A(n17844), .B(n18162), .ZN(
        P3_U2824) );
  OAI21_X1 U20987 ( .B1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n17846), .A(
        n17845), .ZN(n18176) );
  AOI21_X1 U20988 ( .B1(n17849), .B2(n17848), .A(n17847), .ZN(n18174) );
  AOI22_X1 U20989 ( .A1(n17894), .A2(n18174), .B1(n18231), .B2(
        P3_REIP_REG_5__SCAN_IN), .ZN(n17858) );
  AOI221_X1 U20990 ( .B1(n17876), .B2(n17852), .C1(n17851), .C2(n17852), .A(
        n17850), .ZN(n17856) );
  NAND2_X1 U20991 ( .A1(n17853), .A2(n18626), .ZN(n17855) );
  AOI22_X1 U20992 ( .A1(n17856), .A2(n17855), .B1(n17854), .B2(n17903), .ZN(
        n17857) );
  OAI211_X1 U20993 ( .C1(n17913), .C2(n18176), .A(n17858), .B(n17857), .ZN(
        P3_U2825) );
  OAI21_X1 U20994 ( .B1(n17861), .B2(n17860), .A(n17859), .ZN(n18182) );
  OAI22_X1 U20995 ( .A1(n17913), .A2(n18182), .B1(n18343), .B2(n17862), .ZN(
        n17863) );
  AOI21_X1 U20996 ( .B1(n18231), .B2(P3_REIP_REG_4__SCAN_IN), .A(n17863), .ZN(
        n17870) );
  AOI21_X1 U20997 ( .B1(n17866), .B2(n17865), .A(n17864), .ZN(n18184) );
  OAI21_X1 U20998 ( .B1(n17868), .B2(n17867), .A(n17910), .ZN(n17877) );
  AOI22_X1 U20999 ( .A1(n17894), .A2(n18184), .B1(
        P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n17877), .ZN(n17869) );
  OAI211_X1 U21000 ( .C1(n17897), .C2(n17871), .A(n17870), .B(n17869), .ZN(
        P3_U2826) );
  AOI21_X1 U21001 ( .B1(n17874), .B2(n17873), .A(n17872), .ZN(n18197) );
  AOI22_X1 U21002 ( .A1(n17894), .A2(n18197), .B1(n17875), .B2(n17903), .ZN(
        n17883) );
  NOR2_X1 U21003 ( .A1(n17876), .A2(n17888), .ZN(n17887) );
  OAI21_X1 U21004 ( .B1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n17887), .A(
        n17877), .ZN(n17882) );
  NAND2_X1 U21005 ( .A1(n18231), .A2(P3_REIP_REG_3__SCAN_IN), .ZN(n18194) );
  INV_X1 U21006 ( .A(n17913), .ZN(n17880) );
  OAI211_X1 U21007 ( .C1(n17878), .C2(n18190), .A(n17880), .B(n18189), .ZN(
        n17881) );
  NAND4_X1 U21008 ( .A1(n17883), .A2(n17882), .A3(n18194), .A4(n17881), .ZN(
        P3_U2827) );
  AOI21_X1 U21009 ( .B1(n17886), .B2(n17885), .A(n17884), .ZN(n18212) );
  AOI21_X1 U21010 ( .B1(n17888), .B2(n18343), .A(n17887), .ZN(n17893) );
  OAI21_X1 U21011 ( .B1(n17891), .B2(n17890), .A(n17889), .ZN(n18209) );
  INV_X1 U21012 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n18771) );
  OAI22_X1 U21013 ( .A1(n17913), .A2(n18209), .B1(n18218), .B2(n18771), .ZN(
        n17892) );
  AOI211_X1 U21014 ( .C1(n18212), .C2(n17894), .A(n17893), .B(n17892), .ZN(
        n17895) );
  OAI21_X1 U21015 ( .B1(n17897), .B2(n17896), .A(n17895), .ZN(P3_U2828) );
  NOR2_X1 U21016 ( .A1(n17898), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n17899) );
  XNOR2_X1 U21017 ( .A(n17899), .B(n17901), .ZN(n18225) );
  OAI21_X1 U21018 ( .B1(n17901), .B2(n17907), .A(n17900), .ZN(n18217) );
  OAI22_X1 U21019 ( .A1(n17913), .A2(n18217), .B1(n18218), .B2(n20815), .ZN(
        n17902) );
  AOI221_X1 U21020 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n17905), .C1(
        n17904), .C2(n17903), .A(n17902), .ZN(n17906) );
  OAI21_X1 U21021 ( .B1(n18225), .B2(n17914), .A(n17906), .ZN(P3_U2829) );
  AOI21_X1 U21022 ( .B1(n17908), .B2(n18226), .A(n17907), .ZN(n17915) );
  INV_X1 U21023 ( .A(n17915), .ZN(n18234) );
  NAND3_X1 U21024 ( .A1(n18236), .A2(n17910), .A3(n17909), .ZN(n17911) );
  AOI22_X1 U21025 ( .A1(n18231), .A2(P3_REIP_REG_0__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17911), .ZN(n17912) );
  OAI221_X1 U21026 ( .B1(n17915), .B2(n17914), .C1(n18234), .C2(n17913), .A(
        n17912), .ZN(P3_U2830) );
  NAND2_X1 U21027 ( .A1(n18692), .A2(n18203), .ZN(n18216) );
  OAI21_X1 U21028 ( .B1(n18714), .B2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n17940), .ZN(n17922) );
  AOI22_X1 U21029 ( .A1(n18681), .A2(n17917), .B1(n18102), .B2(n17916), .ZN(
        n17920) );
  NOR2_X1 U21030 ( .A1(n18692), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n18206) );
  NAND2_X1 U21031 ( .A1(n17919), .A2(n17918), .ZN(n17941) );
  NAND2_X1 U21032 ( .A1(n18714), .A2(n18692), .ZN(n18178) );
  OAI21_X1 U21033 ( .B1(n18206), .B2(n17941), .A(n18178), .ZN(n17945) );
  NAND2_X1 U21034 ( .A1(n17920), .A2(n17945), .ZN(n17921) );
  AOI211_X1 U21035 ( .C1(n17923), .C2(n18216), .A(n17922), .B(n17921), .ZN(
        n17932) );
  OAI211_X1 U21036 ( .C1(n18714), .C2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B(n17932), .ZN(n17924) );
  OAI221_X1 U21037 ( .B1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n17925), 
        .C1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n17930), .A(n17924), .ZN(
        n17929) );
  AOI22_X1 U21038 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n18220), .B1(
        n18147), .B2(n17926), .ZN(n17928) );
  OAI211_X1 U21039 ( .C1(n18214), .C2(n17929), .A(n17928), .B(n17927), .ZN(
        P3_U2835) );
  INV_X1 U21040 ( .A(n17930), .ZN(n17965) );
  NOR2_X1 U21041 ( .A1(n17965), .A2(n17931), .ZN(n17934) );
  INV_X1 U21042 ( .A(n17932), .ZN(n17933) );
  MUX2_X1 U21043 ( .A(n17934), .B(n17933), .S(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .Z(n17935) );
  AOI22_X1 U21044 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n18220), .B1(
        n18227), .B2(n17935), .ZN(n17938) );
  INV_X1 U21045 ( .A(n17936), .ZN(n17937) );
  OAI211_X1 U21046 ( .C1(n17939), .C2(n18123), .A(n17938), .B(n17937), .ZN(
        P3_U2836) );
  AND2_X1 U21047 ( .A1(n17940), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n17946) );
  OAI22_X1 U21048 ( .A1(n18203), .A2(n17942), .B1(n18200), .B2(n17941), .ZN(
        n17943) );
  OAI21_X1 U21049 ( .B1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n17943), .A(
        n18227), .ZN(n17944) );
  AOI21_X1 U21050 ( .B1(n17946), .B2(n17945), .A(n17944), .ZN(n17947) );
  AOI211_X1 U21051 ( .C1(n18220), .C2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n17948), .B(n17947), .ZN(n17952) );
  AOI22_X1 U21052 ( .A1(n18230), .A2(n17950), .B1(n18147), .B2(n17949), .ZN(
        n17951) );
  OAI211_X1 U21053 ( .C1(n18151), .C2(n17953), .A(n17952), .B(n17951), .ZN(
        P3_U2837) );
  INV_X1 U21054 ( .A(n17997), .ZN(n18009) );
  AOI22_X1 U21055 ( .A1(n18147), .A2(n17955), .B1(n18009), .B2(n17954), .ZN(
        n17963) );
  AOI22_X1 U21056 ( .A1(n18681), .A2(n17957), .B1(n18102), .B2(n17956), .ZN(
        n17959) );
  INV_X1 U21057 ( .A(n18206), .ZN(n18180) );
  OAI21_X1 U21058 ( .B1(n18016), .B2(n17964), .A(n18178), .ZN(n17958) );
  NAND4_X1 U21059 ( .A1(n17959), .A2(n18195), .A3(n18180), .A4(n17958), .ZN(
        n17961) );
  AOI221_X1 U21060 ( .B1(n17964), .B2(n18710), .C1(n18017), .C2(n18710), .A(
        n17961), .ZN(n17960) );
  AOI21_X1 U21061 ( .B1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n17960), .A(
        n18231), .ZN(n17966) );
  OAI211_X1 U21062 ( .C1(n18139), .C2(n17961), .A(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B(n17966), .ZN(n17962) );
  OAI211_X1 U21063 ( .C1(n18809), .C2(n18218), .A(n17963), .B(n17962), .ZN(
        P3_U2838) );
  NOR3_X1 U21064 ( .A1(n18220), .A2(n17965), .A3(n17964), .ZN(n17967) );
  OAI21_X1 U21065 ( .B1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n17967), .A(
        n17966), .ZN(n17968) );
  OAI211_X1 U21066 ( .C1(n17970), .C2(n18123), .A(n17969), .B(n17968), .ZN(
        P3_U2839) );
  INV_X1 U21067 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n21139) );
  AOI21_X1 U21068 ( .B1(n17972), .B2(n18147), .A(n17971), .ZN(n17984) );
  OAI21_X1 U21069 ( .B1(n18016), .B2(n18000), .A(n18699), .ZN(n17973) );
  OAI221_X1 U21070 ( .B1(n18203), .B2(n17974), .C1(n18203), .C2(n17986), .A(
        n17973), .ZN(n17999) );
  INV_X1 U21071 ( .A(n18681), .ZN(n18085) );
  NAND2_X1 U21072 ( .A1(n18085), .A2(n18083), .ZN(n18106) );
  INV_X1 U21073 ( .A(n18106), .ZN(n17975) );
  OAI22_X1 U21074 ( .A1(n18714), .A2(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .B1(
        n17976), .B2(n17975), .ZN(n17977) );
  NOR2_X1 U21075 ( .A1(n17999), .A2(n17977), .ZN(n17991) );
  OAI22_X1 U21076 ( .A1(n18058), .A2(n18085), .B1(n18048), .B2(n18083), .ZN(
        n17985) );
  OAI21_X1 U21077 ( .B1(n18118), .B2(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n17978) );
  AOI211_X1 U21078 ( .C1(n18710), .C2(n17988), .A(n17985), .B(n17978), .ZN(
        n17979) );
  OAI211_X1 U21079 ( .C1(n18692), .C2(n17980), .A(n17991), .B(n17979), .ZN(
        n17981) );
  OAI211_X1 U21080 ( .C1(n17982), .C2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n18227), .B(n17981), .ZN(n17983) );
  OAI211_X1 U21081 ( .C1(n18195), .C2(n21139), .A(n17984), .B(n17983), .ZN(
        P3_U2840) );
  INV_X1 U21082 ( .A(n18039), .ZN(n17987) );
  NOR2_X1 U21083 ( .A1(n18214), .A2(n17985), .ZN(n18037) );
  OAI221_X1 U21084 ( .B1(n18692), .B2(n17987), .C1(n18692), .C2(n17986), .A(
        n18037), .ZN(n17998) );
  AOI21_X1 U21085 ( .B1(n17988), .B2(n18216), .A(n17998), .ZN(n17990) );
  AOI211_X1 U21086 ( .C1(n17991), .C2(n17990), .A(n18231), .B(n17989), .ZN(
        n17992) );
  AOI211_X1 U21087 ( .C1(n18147), .C2(n17994), .A(n17993), .B(n17992), .ZN(
        n17995) );
  OAI21_X1 U21088 ( .B1(n17997), .B2(n17996), .A(n17995), .ZN(P3_U2841) );
  NAND3_X1 U21089 ( .A1(n18015), .A2(P3_STATE2_REG_2__SCAN_IN), .A3(n18216), 
        .ZN(n18002) );
  AOI211_X1 U21090 ( .C1(n18000), .C2(n18106), .A(n17999), .B(n17998), .ZN(
        n18001) );
  OR2_X1 U21091 ( .A1(n18231), .A2(n18001), .ZN(n18014) );
  NAND2_X1 U21092 ( .A1(n18002), .A2(n18014), .ZN(n18004) );
  AOI22_X1 U21093 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n18004), .B1(
        n18009), .B2(n18003), .ZN(n18006) );
  OAI211_X1 U21094 ( .C1(n18123), .C2(n18007), .A(n18006), .B(n18005), .ZN(
        P3_U2842) );
  AOI22_X1 U21095 ( .A1(n18147), .A2(n18010), .B1(n18009), .B2(n18008), .ZN(
        n18013) );
  INV_X1 U21096 ( .A(n18011), .ZN(n18012) );
  OAI211_X1 U21097 ( .C1(n18015), .C2(n18014), .A(n18013), .B(n18012), .ZN(
        P3_U2843) );
  INV_X1 U21098 ( .A(n18178), .ZN(n18204) );
  NOR3_X1 U21099 ( .A1(n18206), .A2(n18016), .A3(n18043), .ZN(n18020) );
  AOI222_X1 U21100 ( .A1(n18710), .A2(n18018), .B1(n18710), .B2(n18017), .C1(
        n18018), .C2(n18106), .ZN(n18019) );
  OAI211_X1 U21101 ( .C1(n18204), .C2(n18020), .A(n18037), .B(n18019), .ZN(
        n18033) );
  OAI221_X1 U21102 ( .B1(n18033), .B2(n21008), .C1(n18033), .C2(n18178), .A(
        n18218), .ZN(n18030) );
  INV_X1 U21103 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n18171) );
  OAI22_X1 U21104 ( .A1(n18203), .A2(n18201), .B1(n18179), .B2(n18200), .ZN(
        n18192) );
  AND2_X1 U21105 ( .A1(n18192), .A2(n18227), .ZN(n18177) );
  NAND3_X1 U21106 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(n18177), .ZN(n18172) );
  NOR2_X1 U21107 ( .A1(n18171), .A2(n18172), .ZN(n18153) );
  AOI222_X1 U21108 ( .A1(n18023), .A2(n18230), .B1(n18022), .B2(n18021), .C1(
        n18050), .C2(n18153), .ZN(n18119) );
  NOR2_X1 U21109 ( .A1(n18119), .A2(n18024), .ZN(n18044) );
  AOI22_X1 U21110 ( .A1(n18147), .A2(n18026), .B1(n18025), .B2(n18044), .ZN(
        n18029) );
  INV_X1 U21111 ( .A(n18027), .ZN(n18028) );
  OAI211_X1 U21112 ( .C1(n18031), .C2(n18030), .A(n18029), .B(n18028), .ZN(
        P3_U2844) );
  AOI22_X1 U21113 ( .A1(n18231), .A2(P3_REIP_REG_17__SCAN_IN), .B1(n18147), 
        .B2(n18032), .ZN(n18036) );
  NAND3_X1 U21114 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n18218), .A3(
        n18033), .ZN(n18035) );
  NAND3_X1 U21115 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n18044), .A3(
        n21008), .ZN(n18034) );
  NAND3_X1 U21116 ( .A1(n18036), .A2(n18035), .A3(n18034), .ZN(P3_U2845) );
  INV_X1 U21117 ( .A(n18037), .ZN(n18042) );
  AOI22_X1 U21118 ( .A1(n18710), .A2(n18038), .B1(n18699), .B2(n18066), .ZN(
        n18130) );
  OAI21_X1 U21119 ( .B1(n18059), .B2(n18712), .A(n18039), .ZN(n18040) );
  OAI211_X1 U21120 ( .C1(n18118), .C2(n18041), .A(n18130), .B(n18040), .ZN(
        n18053) );
  OAI221_X1 U21121 ( .B1(n18042), .B2(n18139), .C1(n18042), .C2(n18053), .A(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n18047) );
  AOI22_X1 U21122 ( .A1(n18045), .A2(n18147), .B1(n18044), .B2(n18043), .ZN(
        n18046) );
  OAI221_X1 U21123 ( .B1(n18231), .B2(n18047), .C1(n18218), .C2(n20933), .A(
        n18046), .ZN(P3_U2846) );
  NOR2_X1 U21124 ( .A1(n18048), .A2(n18083), .ZN(n18056) );
  INV_X1 U21125 ( .A(n18049), .ZN(n18052) );
  NAND4_X1 U21126 ( .A1(n18192), .A2(n18052), .A3(n18051), .A4(n18050), .ZN(
        n18072) );
  OAI21_X1 U21127 ( .B1(n18074), .B2(n18072), .A(n18059), .ZN(n18054) );
  AOI22_X1 U21128 ( .A1(n18056), .A2(n18055), .B1(n18054), .B2(n18053), .ZN(
        n18064) );
  NOR3_X1 U21129 ( .A1(n18058), .A2(n18057), .A3(n18224), .ZN(n18061) );
  OAI22_X1 U21130 ( .A1(n18059), .A2(n18195), .B1(n18218), .B2(n18793), .ZN(
        n18060) );
  AOI211_X1 U21131 ( .C1(n18062), .C2(n18147), .A(n18061), .B(n18060), .ZN(
        n18063) );
  OAI21_X1 U21132 ( .B1(n18064), .B2(n18214), .A(n18063), .ZN(P3_U2847) );
  INV_X1 U21133 ( .A(n18065), .ZN(n18080) );
  NOR2_X1 U21134 ( .A1(n18226), .A2(n18066), .ZN(n18129) );
  OAI221_X1 U21135 ( .B1(n18692), .B2(n18070), .C1(n18692), .C2(n18129), .A(
        n18130), .ZN(n18088) );
  AOI22_X1 U21136 ( .A1(n18699), .A2(n18068), .B1(n18067), .B2(n18216), .ZN(
        n18069) );
  OAI211_X1 U21137 ( .C1(n18070), .C2(n18203), .A(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B(n18069), .ZN(n18071) );
  OAI21_X1 U21138 ( .B1(n18088), .B2(n18071), .A(n18227), .ZN(n18073) );
  AOI222_X1 U21139 ( .A1(n18074), .A2(n18073), .B1(n18074), .B2(n18072), .C1(
        n18073), .C2(n18195), .ZN(n18078) );
  OAI22_X1 U21140 ( .A1(n18076), .A2(n18123), .B1(n18151), .B2(n18075), .ZN(
        n18077) );
  AOI211_X1 U21141 ( .C1(n18231), .C2(P3_REIP_REG_14__SCAN_IN), .A(n18078), 
        .B(n18077), .ZN(n18079) );
  OAI21_X1 U21142 ( .B1(n18224), .B2(n18080), .A(n18079), .ZN(P3_U2848) );
  INV_X1 U21143 ( .A(n18119), .ZN(n18126) );
  NAND2_X1 U21144 ( .A1(n18081), .A2(n18126), .ZN(n18094) );
  AOI22_X1 U21145 ( .A1(n18231), .A2(P3_REIP_REG_13__SCAN_IN), .B1(n18147), 
        .B2(n18082), .ZN(n18091) );
  OAI22_X1 U21146 ( .A1(n18086), .A2(n18085), .B1(n18084), .B2(n18083), .ZN(
        n18087) );
  AOI211_X1 U21147 ( .C1(n18109), .C2(n18108), .A(n18088), .B(n18087), .ZN(
        n18095) );
  OAI211_X1 U21148 ( .C1(n18118), .C2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n18227), .B(n18095), .ZN(n18089) );
  NAND3_X1 U21149 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n18218), .A3(
        n18089), .ZN(n18090) );
  OAI211_X1 U21150 ( .C1(n18094), .C2(n18092), .A(n18091), .B(n18090), .ZN(
        P3_U2849) );
  NAND2_X1 U21151 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n18227), .ZN(
        n18093) );
  AOI22_X1 U21152 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n18095), .B1(
        n18094), .B2(n18093), .ZN(n18096) );
  AOI21_X1 U21153 ( .B1(n18147), .B2(n18097), .A(n18096), .ZN(n18099) );
  OAI211_X1 U21154 ( .C1(n18195), .C2(n18100), .A(n18099), .B(n18098), .ZN(
        P3_U2850) );
  AOI22_X1 U21155 ( .A1(n18681), .A2(n18103), .B1(n18102), .B2(n18101), .ZN(
        n18104) );
  NAND2_X1 U21156 ( .A1(n18227), .A2(n18104), .ZN(n18131) );
  OAI221_X1 U21157 ( .B1(n18692), .B2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .C1(
        n18692), .C2(n18129), .A(n18130), .ZN(n18105) );
  AOI211_X1 U21158 ( .C1(n18107), .C2(n18106), .A(n18131), .B(n18105), .ZN(
        n18117) );
  AOI22_X1 U21159 ( .A1(n18109), .A2(n18108), .B1(n18712), .B2(n18116), .ZN(
        n18110) );
  AOI211_X1 U21160 ( .C1(n18117), .C2(n18110), .A(n18231), .B(n13132), .ZN(
        n18112) );
  AOI211_X1 U21161 ( .C1(n18113), .C2(n18126), .A(n18112), .B(n18111), .ZN(
        n18114) );
  OAI21_X1 U21162 ( .B1(n18115), .B2(n18123), .A(n18114), .ZN(P3_U2851) );
  AOI221_X1 U21163 ( .B1(n18118), .B2(n18117), .C1(
        P3_INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n18117), .A(n18116), .ZN(
        n18121) );
  NOR3_X1 U21164 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n18119), .A3(
        n18127), .ZN(n18120) );
  AOI221_X1 U21165 ( .B1(P3_REIP_REG_10__SCAN_IN), .B2(n18231), .C1(n18121), 
        .C2(n18218), .A(n18120), .ZN(n18122) );
  OAI21_X1 U21166 ( .B1(n18124), .B2(n18123), .A(n18122), .ZN(P3_U2852) );
  INV_X1 U21167 ( .A(n18125), .ZN(n18128) );
  AOI22_X1 U21168 ( .A1(n18147), .A2(n18128), .B1(n18127), .B2(n18126), .ZN(
        n18135) );
  AOI21_X1 U21169 ( .B1(n18130), .B2(n18692), .A(n18129), .ZN(n18132) );
  OAI211_X1 U21170 ( .C1(n18132), .C2(n18131), .A(
        P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B(n18218), .ZN(n18133) );
  NAND3_X1 U21171 ( .A1(n18135), .A2(n18134), .A3(n18133), .ZN(P3_U2853) );
  INV_X1 U21172 ( .A(n18153), .ZN(n18164) );
  NOR3_X1 U21173 ( .A1(n20916), .A2(n18163), .A3(n18164), .ZN(n18145) );
  OAI22_X1 U21174 ( .A1(n18137), .A2(n18204), .B1(n18136), .B2(n18203), .ZN(
        n18138) );
  OR2_X1 U21175 ( .A1(n18206), .A2(n18138), .ZN(n18161) );
  AOI211_X1 U21176 ( .C1(n18139), .C2(n18163), .A(n20916), .B(n18161), .ZN(
        n18156) );
  OAI21_X1 U21177 ( .B1(n18156), .B2(n18140), .A(n18195), .ZN(n18143) );
  INV_X1 U21178 ( .A(n18141), .ZN(n18142) );
  AOI221_X1 U21179 ( .B1(n18145), .B2(n18144), .C1(n18143), .C2(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A(n18142), .ZN(n18150) );
  AOI22_X1 U21180 ( .A1(n18230), .A2(n18148), .B1(n18147), .B2(n18146), .ZN(
        n18149) );
  OAI211_X1 U21181 ( .C1(n18152), .C2(n18151), .A(n18150), .B(n18149), .ZN(
        P3_U2854) );
  AOI22_X1 U21182 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n18227), .B1(
        P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n18153), .ZN(n18155) );
  OAI22_X1 U21183 ( .A1(n18156), .A2(n18155), .B1(n18224), .B2(n18154), .ZN(
        n18157) );
  AOI211_X1 U21184 ( .C1(n18220), .C2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n18158), .B(n18157), .ZN(n18159) );
  OAI21_X1 U21185 ( .B1(n18235), .B2(n18160), .A(n18159), .ZN(P3_U2855) );
  AOI21_X1 U21186 ( .B1(n18227), .B2(n18161), .A(n18220), .ZN(n18170) );
  OAI221_X1 U21187 ( .B1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n18164), .C1(
        n18163), .C2(n18170), .A(n18162), .ZN(n18165) );
  AOI21_X1 U21188 ( .B1(n18230), .B2(n18166), .A(n18165), .ZN(n18167) );
  OAI21_X1 U21189 ( .B1(n18235), .B2(n18168), .A(n18167), .ZN(P3_U2856) );
  NAND2_X1 U21190 ( .A1(n18231), .A2(P3_REIP_REG_5__SCAN_IN), .ZN(n18169) );
  OAI221_X1 U21191 ( .B1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n18172), .C1(
        n18171), .C2(n18170), .A(n18169), .ZN(n18173) );
  AOI21_X1 U21192 ( .B1(n18230), .B2(n18174), .A(n18173), .ZN(n18175) );
  OAI21_X1 U21193 ( .B1(n18235), .B2(n18176), .A(n18175), .ZN(P3_U2857) );
  NAND2_X1 U21194 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n18177), .ZN(
        n18188) );
  AOI22_X1 U21195 ( .A1(n18710), .A2(n18201), .B1(n18179), .B2(n18178), .ZN(
        n18181) );
  NAND3_X1 U21196 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n18181), .A3(
        n18180), .ZN(n18191) );
  AOI21_X1 U21197 ( .B1(n18221), .B2(n18191), .A(n18220), .ZN(n18186) );
  OAI22_X1 U21198 ( .A1(n18218), .A2(n18774), .B1(n18235), .B2(n18182), .ZN(
        n18183) );
  AOI21_X1 U21199 ( .B1(n18230), .B2(n18184), .A(n18183), .ZN(n18185) );
  OAI221_X1 U21200 ( .B1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n18188), .C1(
        n18187), .C2(n18186), .A(n18185), .ZN(P3_U2858) );
  OAI21_X1 U21201 ( .B1(n17878), .B2(n18190), .A(n18189), .ZN(n18199) );
  OAI211_X1 U21202 ( .C1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .C2(n18192), .A(
        n18227), .B(n18191), .ZN(n18193) );
  OAI211_X1 U21203 ( .C1(n18195), .C2(n13112), .A(n18194), .B(n18193), .ZN(
        n18196) );
  AOI21_X1 U21204 ( .B1(n18230), .B2(n18197), .A(n18196), .ZN(n18198) );
  OAI21_X1 U21205 ( .B1(n18235), .B2(n18199), .A(n18198), .ZN(P3_U2859) );
  NOR3_X1 U21206 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n13107), .A3(
        n18200), .ZN(n18211) );
  NAND2_X1 U21207 ( .A1(n18710), .A2(n18201), .ZN(n18208) );
  NAND2_X1 U21208 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18202) );
  OAI22_X1 U21209 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n18204), .B1(
        n18203), .B2(n18202), .ZN(n18205) );
  OAI21_X1 U21210 ( .B1(n18206), .B2(n18205), .A(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18207) );
  OAI211_X1 U21211 ( .C1(n18209), .C2(n18687), .A(n18208), .B(n18207), .ZN(
        n18210) );
  AOI211_X1 U21212 ( .C1(n18212), .C2(n18681), .A(n18211), .B(n18210), .ZN(
        n18215) );
  AOI22_X1 U21213 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n18220), .B1(
        n18231), .B2(P3_REIP_REG_2__SCAN_IN), .ZN(n18213) );
  OAI21_X1 U21214 ( .B1(n18215), .B2(n18214), .A(n18213), .ZN(P3_U2860) );
  AND3_X1 U21215 ( .A1(n18226), .A2(n18216), .A3(n18227), .ZN(n18229) );
  OAI22_X1 U21216 ( .A1(n18218), .A2(n20815), .B1(n18235), .B2(n18217), .ZN(
        n18219) );
  AOI221_X1 U21217 ( .B1(n18220), .B2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .C1(
        n18229), .C2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A(n18219), .ZN(
        n18223) );
  OAI211_X1 U21218 ( .C1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(n18699), .A(
        n18221), .B(n13107), .ZN(n18222) );
  OAI211_X1 U21219 ( .C1(n18225), .C2(n18224), .A(n18223), .B(n18222), .ZN(
        P3_U2861) );
  AOI211_X1 U21220 ( .C1(n18714), .C2(n18227), .A(n18231), .B(n18226), .ZN(
        n18228) );
  AOI211_X1 U21221 ( .C1(n18230), .C2(n18234), .A(n18229), .B(n18228), .ZN(
        n18233) );
  NAND2_X1 U21222 ( .A1(n18231), .A2(P3_REIP_REG_0__SCAN_IN), .ZN(n18232) );
  OAI211_X1 U21223 ( .C1(n18235), .C2(n18234), .A(n18233), .B(n18232), .ZN(
        P3_U2862) );
  INV_X1 U21224 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18527) );
  AOI211_X1 U21225 ( .C1(n21087), .C2(n18237), .A(n18901), .B(n18236), .ZN(
        n18737) );
  OAI21_X1 U21226 ( .B1(n18737), .B2(n18281), .A(n18242), .ZN(n18238) );
  OAI221_X1 U21227 ( .B1(n18527), .B2(n18883), .C1(n18527), .C2(n18242), .A(
        n18238), .ZN(P3_U2863) );
  INV_X1 U21228 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18726) );
  NOR2_X1 U21229 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18726), .ZN(
        n18528) );
  NOR2_X1 U21230 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18723), .ZN(
        n18412) );
  NOR2_X1 U21231 ( .A1(n18528), .A2(n18412), .ZN(n18240) );
  OAI22_X1 U21232 ( .A1(n18241), .A2(n18726), .B1(n18240), .B2(n18239), .ZN(
        P3_U2866) );
  NOR2_X1 U21233 ( .A1(n18727), .A2(n18242), .ZN(P3_U2867) );
  NAND2_X1 U21234 ( .A1(n18626), .A2(BUF2_REG_16__SCAN_IN), .ZN(n18630) );
  NOR2_X1 U21235 ( .A1(n18723), .A2(n18726), .ZN(n18563) );
  NOR2_X1 U21236 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18718), .ZN(
        n18481) );
  NAND2_X1 U21237 ( .A1(n18563), .A2(n18481), .ZN(n18604) );
  NOR2_X2 U21238 ( .A1(n18342), .A2(n21157), .ZN(n18622) );
  NAND2_X1 U21239 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18717) );
  INV_X1 U21240 ( .A(n18563), .ZN(n18243) );
  NOR2_X2 U21241 ( .A1(n18717), .A2(n18243), .ZN(n18675) );
  NAND2_X1 U21242 ( .A1(n18718), .A2(n18527), .ZN(n18719) );
  NAND2_X1 U21243 ( .A1(n18723), .A2(n18726), .ZN(n18366) );
  NOR2_X2 U21244 ( .A1(n18719), .A2(n18366), .ZN(n18338) );
  NOR2_X1 U21245 ( .A1(n18675), .A2(n18338), .ZN(n18300) );
  NOR2_X1 U21246 ( .A1(n18745), .A2(n18300), .ZN(n18275) );
  NAND2_X1 U21247 ( .A1(n18563), .A2(n18718), .ZN(n18561) );
  NOR2_X2 U21248 ( .A1(n18527), .A2(n18561), .ZN(n18652) );
  AND2_X1 U21249 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n18626), .ZN(n18621) );
  AOI22_X1 U21250 ( .A1(n18622), .A2(n18275), .B1(n18652), .B2(n18621), .ZN(
        n18250) );
  NOR2_X1 U21251 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18527), .ZN(
        n18457) );
  NOR2_X1 U21252 ( .A1(n18481), .A2(n18457), .ZN(n18530) );
  NOR2_X1 U21253 ( .A1(n18530), .A2(n18243), .ZN(n18594) );
  AOI21_X1 U21254 ( .B1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(
        P3_STATE2_REG_3__SCAN_IN), .A(n18342), .ZN(n18591) );
  INV_X1 U21255 ( .A(n18300), .ZN(n18244) );
  AOI22_X1 U21256 ( .A1(n18626), .A2(n18594), .B1(n18591), .B2(n18244), .ZN(
        n18278) );
  INV_X1 U21257 ( .A(n18245), .ZN(n18246) );
  NAND2_X1 U21258 ( .A1(n18247), .A2(n18246), .ZN(n18276) );
  NOR2_X1 U21259 ( .A1(n18248), .A2(n18276), .ZN(n18627) );
  AOI22_X1 U21260 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n18278), .B1(
        n18338), .B2(n18627), .ZN(n18249) );
  OAI211_X1 U21261 ( .C1(n18630), .C2(n18604), .A(n18250), .B(n18249), .ZN(
        P3_U2868) );
  INV_X1 U21262 ( .A(n18652), .ZN(n18680) );
  NAND2_X1 U21263 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n18626), .ZN(n18601) );
  INV_X1 U21264 ( .A(n18604), .ZN(n18616) );
  NAND2_X1 U21265 ( .A1(n18626), .A2(BUF2_REG_17__SCAN_IN), .ZN(n18636) );
  INV_X1 U21266 ( .A(n18636), .ZN(n18598) );
  AND2_X1 U21267 ( .A1(n18532), .A2(BUF2_REG_1__SCAN_IN), .ZN(n18631) );
  AOI22_X1 U21268 ( .A1(n18616), .A2(n18598), .B1(n18275), .B2(n18631), .ZN(
        n18252) );
  NOR2_X2 U21269 ( .A1(n18886), .A2(n18276), .ZN(n18633) );
  AOI22_X1 U21270 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n18278), .B1(
        n18338), .B2(n18633), .ZN(n18251) );
  OAI211_X1 U21271 ( .C1(n18680), .C2(n18601), .A(n18252), .B(n18251), .ZN(
        P3_U2869) );
  NAND2_X1 U21272 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n18626), .ZN(n18572) );
  AND2_X1 U21273 ( .A1(n18626), .A2(BUF2_REG_18__SCAN_IN), .ZN(n18639) );
  NOR2_X2 U21274 ( .A1(n18342), .A2(n18253), .ZN(n18637) );
  AOI22_X1 U21275 ( .A1(n18616), .A2(n18639), .B1(n18275), .B2(n18637), .ZN(
        n18256) );
  AOI22_X1 U21276 ( .A1(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n18278), .B1(
        n18338), .B2(n18569), .ZN(n18255) );
  OAI211_X1 U21277 ( .C1(n18680), .C2(n18572), .A(n18256), .B(n18255), .ZN(
        P3_U2870) );
  NAND2_X1 U21278 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n18626), .ZN(n18649) );
  NAND2_X1 U21279 ( .A1(n18626), .A2(BUF2_REG_19__SCAN_IN), .ZN(n18576) );
  INV_X1 U21280 ( .A(n18576), .ZN(n18645) );
  NOR2_X2 U21281 ( .A1(n18342), .A2(n18257), .ZN(n18644) );
  AOI22_X1 U21282 ( .A1(n18616), .A2(n18645), .B1(n18275), .B2(n18644), .ZN(
        n18260) );
  NOR2_X2 U21283 ( .A1(n18258), .A2(n18276), .ZN(n18646) );
  AOI22_X1 U21284 ( .A1(P3_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n18278), .B1(
        n18338), .B2(n18646), .ZN(n18259) );
  OAI211_X1 U21285 ( .C1(n18680), .C2(n18649), .A(n18260), .B(n18259), .ZN(
        P3_U2871) );
  NAND2_X1 U21286 ( .A1(n18626), .A2(BUF2_REG_20__SCAN_IN), .ZN(n18545) );
  NOR2_X2 U21287 ( .A1(n18342), .A2(n18261), .ZN(n18650) );
  NAND2_X1 U21288 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n18626), .ZN(n18657) );
  INV_X1 U21289 ( .A(n18657), .ZN(n18542) );
  AOI22_X1 U21290 ( .A1(n18275), .A2(n18650), .B1(n18652), .B2(n18542), .ZN(
        n18264) );
  NOR2_X2 U21291 ( .A1(n18262), .A2(n18276), .ZN(n18653) );
  AOI22_X1 U21292 ( .A1(P3_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n18278), .B1(
        n18338), .B2(n18653), .ZN(n18263) );
  OAI211_X1 U21293 ( .C1(n18604), .C2(n18545), .A(n18264), .B(n18263), .ZN(
        P3_U2872) );
  NAND2_X1 U21294 ( .A1(BUF2_REG_21__SCAN_IN), .A2(n18626), .ZN(n18663) );
  NOR2_X2 U21295 ( .A1(n18265), .A2(n18342), .ZN(n18658) );
  NOR2_X1 U21296 ( .A1(n18266), .A2(n18343), .ZN(n18659) );
  AOI22_X1 U21297 ( .A1(n18275), .A2(n18658), .B1(n18652), .B2(n18659), .ZN(
        n18269) );
  NOR2_X2 U21298 ( .A1(n18267), .A2(n18276), .ZN(n18660) );
  AOI22_X1 U21299 ( .A1(P3_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n18278), .B1(
        n18338), .B2(n18660), .ZN(n18268) );
  OAI211_X1 U21300 ( .C1(n18604), .C2(n18663), .A(n18269), .B(n18268), .ZN(
        P3_U2873) );
  NAND2_X1 U21301 ( .A1(BUF2_REG_22__SCAN_IN), .A2(n18626), .ZN(n18669) );
  NOR2_X2 U21302 ( .A1(n18270), .A2(n18342), .ZN(n18664) );
  NAND2_X1 U21303 ( .A1(BUF2_REG_30__SCAN_IN), .A2(n18626), .ZN(n18553) );
  INV_X1 U21304 ( .A(n18553), .ZN(n18665) );
  AOI22_X1 U21305 ( .A1(n18275), .A2(n18664), .B1(n18652), .B2(n18665), .ZN(
        n18273) );
  NOR2_X2 U21306 ( .A1(n18271), .A2(n18276), .ZN(n18666) );
  AOI22_X1 U21307 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n18278), .B1(
        n18338), .B2(n18666), .ZN(n18272) );
  OAI211_X1 U21308 ( .C1(n18604), .C2(n18669), .A(n18273), .B(n18272), .ZN(
        P3_U2874) );
  NAND2_X1 U21309 ( .A1(BUF2_REG_23__SCAN_IN), .A2(n18626), .ZN(n18679) );
  NOR2_X2 U21310 ( .A1(n18274), .A2(n18342), .ZN(n18671) );
  NAND2_X1 U21311 ( .A1(n18626), .A2(BUF2_REG_31__SCAN_IN), .ZN(n18560) );
  INV_X1 U21312 ( .A(n18560), .ZN(n18673) );
  AOI22_X1 U21313 ( .A1(n18275), .A2(n18671), .B1(n18652), .B2(n18673), .ZN(
        n18280) );
  NOR2_X2 U21314 ( .A1(n18277), .A2(n18276), .ZN(n18674) );
  AOI22_X1 U21315 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n18278), .B1(
        n18338), .B2(n18674), .ZN(n18279) );
  OAI211_X1 U21316 ( .C1(n18604), .C2(n18679), .A(n18280), .B(n18279), .ZN(
        P3_U2875) );
  INV_X1 U21317 ( .A(n18675), .ZN(n18643) );
  NAND2_X1 U21318 ( .A1(n18718), .A2(n18620), .ZN(n18458) );
  NOR2_X1 U21319 ( .A1(n18366), .A2(n18458), .ZN(n18296) );
  AOI22_X1 U21320 ( .A1(n18616), .A2(n18621), .B1(n18622), .B2(n18296), .ZN(
        n18283) );
  NOR2_X1 U21321 ( .A1(n18726), .A2(n18459), .ZN(n18623) );
  INV_X1 U21322 ( .A(n18366), .ZN(n18321) );
  NOR2_X1 U21323 ( .A1(n18342), .A2(n18281), .ZN(n18624) );
  AND2_X1 U21324 ( .A1(n18718), .A2(n18624), .ZN(n18562) );
  AOI22_X1 U21325 ( .A1(n18626), .A2(n18623), .B1(n18321), .B2(n18562), .ZN(
        n18297) );
  NAND2_X1 U21326 ( .A1(n18321), .A2(n18457), .ZN(n18365) );
  INV_X1 U21327 ( .A(n18365), .ZN(n18356) );
  AOI22_X1 U21328 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n18297), .B1(
        n18627), .B2(n18356), .ZN(n18282) );
  OAI211_X1 U21329 ( .C1(n18630), .C2(n18643), .A(n18283), .B(n18282), .ZN(
        P3_U2876) );
  INV_X1 U21330 ( .A(n18601), .ZN(n18632) );
  AOI22_X1 U21331 ( .A1(n18616), .A2(n18632), .B1(n18631), .B2(n18296), .ZN(
        n18285) );
  AOI22_X1 U21332 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n18297), .B1(
        n18633), .B2(n18356), .ZN(n18284) );
  OAI211_X1 U21333 ( .C1(n18643), .C2(n18636), .A(n18285), .B(n18284), .ZN(
        P3_U2877) );
  AOI22_X1 U21334 ( .A1(n18675), .A2(n18639), .B1(n18637), .B2(n18296), .ZN(
        n18287) );
  AOI22_X1 U21335 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n18297), .B1(
        n18569), .B2(n18356), .ZN(n18286) );
  OAI211_X1 U21336 ( .C1(n18604), .C2(n18572), .A(n18287), .B(n18286), .ZN(
        P3_U2878) );
  AOI22_X1 U21337 ( .A1(n18675), .A2(n18645), .B1(n18644), .B2(n18296), .ZN(
        n18289) );
  AOI22_X1 U21338 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n18297), .B1(
        n18646), .B2(n18356), .ZN(n18288) );
  OAI211_X1 U21339 ( .C1(n18604), .C2(n18649), .A(n18289), .B(n18288), .ZN(
        P3_U2879) );
  INV_X1 U21340 ( .A(n18545), .ZN(n18651) );
  AOI22_X1 U21341 ( .A1(n18675), .A2(n18651), .B1(n18650), .B2(n18296), .ZN(
        n18291) );
  AOI22_X1 U21342 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n18297), .B1(
        n18653), .B2(n18356), .ZN(n18290) );
  OAI211_X1 U21343 ( .C1(n18604), .C2(n18657), .A(n18291), .B(n18290), .ZN(
        P3_U2880) );
  INV_X1 U21344 ( .A(n18659), .ZN(n18549) );
  INV_X1 U21345 ( .A(n18663), .ZN(n18546) );
  AOI22_X1 U21346 ( .A1(n18675), .A2(n18546), .B1(n18658), .B2(n18296), .ZN(
        n18293) );
  AOI22_X1 U21347 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n18297), .B1(
        n18660), .B2(n18356), .ZN(n18292) );
  OAI211_X1 U21348 ( .C1(n18604), .C2(n18549), .A(n18293), .B(n18292), .ZN(
        P3_U2881) );
  INV_X1 U21349 ( .A(n18669), .ZN(n18550) );
  AOI22_X1 U21350 ( .A1(n18675), .A2(n18550), .B1(n18664), .B2(n18296), .ZN(
        n18295) );
  AOI22_X1 U21351 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n18297), .B1(
        n18666), .B2(n18356), .ZN(n18294) );
  OAI211_X1 U21352 ( .C1(n18604), .C2(n18553), .A(n18295), .B(n18294), .ZN(
        P3_U2882) );
  INV_X1 U21353 ( .A(n18679), .ZN(n18555) );
  AOI22_X1 U21354 ( .A1(n18675), .A2(n18555), .B1(n18671), .B2(n18296), .ZN(
        n18299) );
  AOI22_X1 U21355 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n18297), .B1(
        n18674), .B2(n18356), .ZN(n18298) );
  OAI211_X1 U21356 ( .C1(n18604), .C2(n18560), .A(n18299), .B(n18298), .ZN(
        P3_U2883) );
  INV_X1 U21357 ( .A(n18627), .ZN(n18597) );
  NAND2_X1 U21358 ( .A1(n18481), .A2(n18321), .ZN(n18382) );
  INV_X1 U21359 ( .A(n18630), .ZN(n18589) );
  INV_X1 U21360 ( .A(n18382), .ZN(n18384) );
  NOR2_X1 U21361 ( .A1(n18356), .A2(n18384), .ZN(n18344) );
  NOR2_X1 U21362 ( .A1(n18745), .A2(n18344), .ZN(n18316) );
  AOI22_X1 U21363 ( .A1(n18589), .A2(n18338), .B1(n18622), .B2(n18316), .ZN(
        n18303) );
  OAI22_X1 U21364 ( .A1(n18300), .A2(n18343), .B1(n18344), .B2(n18342), .ZN(
        n18301) );
  OAI21_X1 U21365 ( .B1(n18384), .B2(n18864), .A(n18301), .ZN(n18317) );
  AOI22_X1 U21366 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n18317), .B1(
        n18675), .B2(n18621), .ZN(n18302) );
  OAI211_X1 U21367 ( .C1(n18597), .C2(n18382), .A(n18303), .B(n18302), .ZN(
        P3_U2884) );
  INV_X1 U21368 ( .A(n18338), .ZN(n18334) );
  AOI22_X1 U21369 ( .A1(n18675), .A2(n18632), .B1(n18631), .B2(n18316), .ZN(
        n18305) );
  AOI22_X1 U21370 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n18317), .B1(
        n18633), .B2(n18384), .ZN(n18304) );
  OAI211_X1 U21371 ( .C1(n18334), .C2(n18636), .A(n18305), .B(n18304), .ZN(
        P3_U2885) );
  AOI22_X1 U21372 ( .A1(n18338), .A2(n18639), .B1(n18637), .B2(n18316), .ZN(
        n18307) );
  AOI22_X1 U21373 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n18317), .B1(
        n18569), .B2(n18384), .ZN(n18306) );
  OAI211_X1 U21374 ( .C1(n18643), .C2(n18572), .A(n18307), .B(n18306), .ZN(
        P3_U2886) );
  INV_X1 U21375 ( .A(n18649), .ZN(n18573) );
  AOI22_X1 U21376 ( .A1(n18675), .A2(n18573), .B1(n18644), .B2(n18316), .ZN(
        n18309) );
  AOI22_X1 U21377 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n18317), .B1(
        n18646), .B2(n18384), .ZN(n18308) );
  OAI211_X1 U21378 ( .C1(n18334), .C2(n18576), .A(n18309), .B(n18308), .ZN(
        P3_U2887) );
  AOI22_X1 U21379 ( .A1(n18338), .A2(n18651), .B1(n18650), .B2(n18316), .ZN(
        n18311) );
  AOI22_X1 U21380 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n18317), .B1(
        n18653), .B2(n18384), .ZN(n18310) );
  OAI211_X1 U21381 ( .C1(n18643), .C2(n18657), .A(n18311), .B(n18310), .ZN(
        P3_U2888) );
  AOI22_X1 U21382 ( .A1(n18675), .A2(n18659), .B1(n18658), .B2(n18316), .ZN(
        n18313) );
  AOI22_X1 U21383 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n18317), .B1(
        n18660), .B2(n18384), .ZN(n18312) );
  OAI211_X1 U21384 ( .C1(n18334), .C2(n18663), .A(n18313), .B(n18312), .ZN(
        P3_U2889) );
  AOI22_X1 U21385 ( .A1(n18675), .A2(n18665), .B1(n18664), .B2(n18316), .ZN(
        n18315) );
  AOI22_X1 U21386 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n18317), .B1(
        n18666), .B2(n18384), .ZN(n18314) );
  OAI211_X1 U21387 ( .C1(n18334), .C2(n18669), .A(n18315), .B(n18314), .ZN(
        P3_U2890) );
  AOI22_X1 U21388 ( .A1(n18338), .A2(n18555), .B1(n18671), .B2(n18316), .ZN(
        n18319) );
  AOI22_X1 U21389 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n18317), .B1(
        n18674), .B2(n18384), .ZN(n18318) );
  OAI211_X1 U21390 ( .C1(n18643), .C2(n18560), .A(n18319), .B(n18318), .ZN(
        P3_U2891) );
  INV_X1 U21391 ( .A(n18717), .ZN(n18505) );
  NAND2_X1 U21392 ( .A1(n18505), .A2(n18321), .ZN(n18405) );
  AOI22_X1 U21393 ( .A1(n18589), .A2(n18356), .B1(n18622), .B2(n18337), .ZN(
        n18323) );
  OAI21_X1 U21394 ( .B1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n18593), .A(
        n18532), .ZN(n18320) );
  AOI21_X1 U21395 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n18717), .A(n18320), 
        .ZN(n18411) );
  NAND2_X1 U21396 ( .A1(n18321), .A2(n18411), .ZN(n18339) );
  AOI22_X1 U21397 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n18339), .B1(
        n18338), .B2(n18621), .ZN(n18322) );
  OAI211_X1 U21398 ( .C1(n18597), .C2(n18405), .A(n18323), .B(n18322), .ZN(
        P3_U2892) );
  AOI22_X1 U21399 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n18339), .B1(
        n18631), .B2(n18337), .ZN(n18325) );
  INV_X1 U21400 ( .A(n18405), .ZN(n18407) );
  AOI22_X1 U21401 ( .A1(n18633), .A2(n18407), .B1(n18598), .B2(n18356), .ZN(
        n18324) );
  OAI211_X1 U21402 ( .C1(n18334), .C2(n18601), .A(n18325), .B(n18324), .ZN(
        P3_U2893) );
  INV_X1 U21403 ( .A(n18569), .ZN(n18642) );
  INV_X1 U21404 ( .A(n18572), .ZN(n18638) );
  AOI22_X1 U21405 ( .A1(n18338), .A2(n18638), .B1(n18637), .B2(n18337), .ZN(
        n18327) );
  AOI22_X1 U21406 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n18339), .B1(
        n18639), .B2(n18356), .ZN(n18326) );
  OAI211_X1 U21407 ( .C1(n18642), .C2(n18405), .A(n18327), .B(n18326), .ZN(
        P3_U2894) );
  AOI22_X1 U21408 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n18339), .B1(
        n18644), .B2(n18337), .ZN(n18329) );
  AOI22_X1 U21409 ( .A1(n18646), .A2(n18407), .B1(n18645), .B2(n18356), .ZN(
        n18328) );
  OAI211_X1 U21410 ( .C1(n18334), .C2(n18649), .A(n18329), .B(n18328), .ZN(
        P3_U2895) );
  AOI22_X1 U21411 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n18339), .B1(
        n18650), .B2(n18337), .ZN(n18331) );
  AOI22_X1 U21412 ( .A1(n18651), .A2(n18356), .B1(n18653), .B2(n18407), .ZN(
        n18330) );
  OAI211_X1 U21413 ( .C1(n18334), .C2(n18657), .A(n18331), .B(n18330), .ZN(
        P3_U2896) );
  AOI22_X1 U21414 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n18339), .B1(
        n18658), .B2(n18337), .ZN(n18333) );
  AOI22_X1 U21415 ( .A1(n18546), .A2(n18356), .B1(n18660), .B2(n18407), .ZN(
        n18332) );
  OAI211_X1 U21416 ( .C1(n18334), .C2(n18549), .A(n18333), .B(n18332), .ZN(
        P3_U2897) );
  AOI22_X1 U21417 ( .A1(n18338), .A2(n18665), .B1(n18664), .B2(n18337), .ZN(
        n18336) );
  AOI22_X1 U21418 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n18339), .B1(
        n18666), .B2(n18407), .ZN(n18335) );
  OAI211_X1 U21419 ( .C1(n18669), .C2(n18365), .A(n18336), .B(n18335), .ZN(
        P3_U2898) );
  AOI22_X1 U21420 ( .A1(n18338), .A2(n18673), .B1(n18671), .B2(n18337), .ZN(
        n18341) );
  AOI22_X1 U21421 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n18339), .B1(
        n18674), .B2(n18407), .ZN(n18340) );
  OAI211_X1 U21422 ( .C1(n18679), .C2(n18365), .A(n18341), .B(n18340), .ZN(
        P3_U2899) );
  INV_X1 U21423 ( .A(n18719), .ZN(n18434) );
  NAND2_X1 U21424 ( .A1(n18434), .A2(n18412), .ZN(n18426) );
  INV_X1 U21425 ( .A(n18426), .ZN(n18430) );
  NOR2_X1 U21426 ( .A1(n18407), .A2(n18430), .ZN(n18388) );
  NOR2_X1 U21427 ( .A1(n18745), .A2(n18388), .ZN(n18361) );
  AOI22_X1 U21428 ( .A1(n18589), .A2(n18384), .B1(n18622), .B2(n18361), .ZN(
        n18347) );
  OAI22_X1 U21429 ( .A1(n18344), .A2(n18343), .B1(n18388), .B2(n18342), .ZN(
        n18345) );
  OAI21_X1 U21430 ( .B1(n18430), .B2(n18864), .A(n18345), .ZN(n18362) );
  AOI22_X1 U21431 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n18362), .B1(
        n18621), .B2(n18356), .ZN(n18346) );
  OAI211_X1 U21432 ( .C1(n18597), .C2(n18426), .A(n18347), .B(n18346), .ZN(
        P3_U2900) );
  AOI22_X1 U21433 ( .A1(n18632), .A2(n18356), .B1(n18631), .B2(n18361), .ZN(
        n18349) );
  AOI22_X1 U21434 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n18362), .B1(
        n18633), .B2(n18430), .ZN(n18348) );
  OAI211_X1 U21435 ( .C1(n18636), .C2(n18382), .A(n18349), .B(n18348), .ZN(
        P3_U2901) );
  AOI22_X1 U21436 ( .A1(n18639), .A2(n18384), .B1(n18637), .B2(n18361), .ZN(
        n18351) );
  AOI22_X1 U21437 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n18362), .B1(
        n18569), .B2(n18430), .ZN(n18350) );
  OAI211_X1 U21438 ( .C1(n18572), .C2(n18365), .A(n18351), .B(n18350), .ZN(
        P3_U2902) );
  AOI22_X1 U21439 ( .A1(n18644), .A2(n18361), .B1(n18645), .B2(n18384), .ZN(
        n18353) );
  AOI22_X1 U21440 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n18362), .B1(
        n18646), .B2(n18430), .ZN(n18352) );
  OAI211_X1 U21441 ( .C1(n18649), .C2(n18365), .A(n18353), .B(n18352), .ZN(
        P3_U2903) );
  AOI22_X1 U21442 ( .A1(n18650), .A2(n18361), .B1(n18542), .B2(n18356), .ZN(
        n18355) );
  AOI22_X1 U21443 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n18362), .B1(
        n18653), .B2(n18430), .ZN(n18354) );
  OAI211_X1 U21444 ( .C1(n18545), .C2(n18382), .A(n18355), .B(n18354), .ZN(
        P3_U2904) );
  AOI22_X1 U21445 ( .A1(n18659), .A2(n18356), .B1(n18658), .B2(n18361), .ZN(
        n18358) );
  AOI22_X1 U21446 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n18362), .B1(
        n18660), .B2(n18430), .ZN(n18357) );
  OAI211_X1 U21447 ( .C1(n18663), .C2(n18382), .A(n18358), .B(n18357), .ZN(
        P3_U2905) );
  AOI22_X1 U21448 ( .A1(n18550), .A2(n18384), .B1(n18664), .B2(n18361), .ZN(
        n18360) );
  AOI22_X1 U21449 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n18362), .B1(
        n18666), .B2(n18430), .ZN(n18359) );
  OAI211_X1 U21450 ( .C1(n18553), .C2(n18365), .A(n18360), .B(n18359), .ZN(
        P3_U2906) );
  AOI22_X1 U21451 ( .A1(n18555), .A2(n18384), .B1(n18671), .B2(n18361), .ZN(
        n18364) );
  AOI22_X1 U21452 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n18362), .B1(
        n18674), .B2(n18430), .ZN(n18363) );
  OAI211_X1 U21453 ( .C1(n18560), .C2(n18365), .A(n18364), .B(n18363), .ZN(
        P3_U2907) );
  NAND2_X1 U21454 ( .A1(n18412), .A2(n18457), .ZN(n18456) );
  INV_X1 U21455 ( .A(n18412), .ZN(n18413) );
  NOR2_X1 U21456 ( .A1(n18413), .A2(n18458), .ZN(n18383) );
  AOI22_X1 U21457 ( .A1(n18589), .A2(n18407), .B1(n18622), .B2(n18383), .ZN(
        n18369) );
  NOR2_X1 U21458 ( .A1(n18718), .A2(n18366), .ZN(n18367) );
  AOI22_X1 U21459 ( .A1(n18626), .A2(n18367), .B1(n18412), .B2(n18562), .ZN(
        n18385) );
  AOI22_X1 U21460 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n18385), .B1(
        n18621), .B2(n18384), .ZN(n18368) );
  OAI211_X1 U21461 ( .C1(n18597), .C2(n18456), .A(n18369), .B(n18368), .ZN(
        P3_U2908) );
  AOI22_X1 U21462 ( .A1(n18632), .A2(n18384), .B1(n18631), .B2(n18383), .ZN(
        n18371) );
  INV_X1 U21463 ( .A(n18456), .ZN(n18445) );
  AOI22_X1 U21464 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n18385), .B1(
        n18633), .B2(n18445), .ZN(n18370) );
  OAI211_X1 U21465 ( .C1(n18636), .C2(n18405), .A(n18371), .B(n18370), .ZN(
        P3_U2909) );
  AOI22_X1 U21466 ( .A1(n18639), .A2(n18407), .B1(n18637), .B2(n18383), .ZN(
        n18373) );
  AOI22_X1 U21467 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n18385), .B1(
        n18569), .B2(n18445), .ZN(n18372) );
  OAI211_X1 U21468 ( .C1(n18572), .C2(n18382), .A(n18373), .B(n18372), .ZN(
        P3_U2910) );
  AOI22_X1 U21469 ( .A1(n18573), .A2(n18384), .B1(n18644), .B2(n18383), .ZN(
        n18375) );
  AOI22_X1 U21470 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n18385), .B1(
        n18646), .B2(n18445), .ZN(n18374) );
  OAI211_X1 U21471 ( .C1(n18576), .C2(n18405), .A(n18375), .B(n18374), .ZN(
        P3_U2911) );
  AOI22_X1 U21472 ( .A1(n18650), .A2(n18383), .B1(n18542), .B2(n18384), .ZN(
        n18377) );
  AOI22_X1 U21473 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n18385), .B1(
        n18653), .B2(n18445), .ZN(n18376) );
  OAI211_X1 U21474 ( .C1(n18545), .C2(n18405), .A(n18377), .B(n18376), .ZN(
        P3_U2912) );
  AOI22_X1 U21475 ( .A1(n18546), .A2(n18407), .B1(n18658), .B2(n18383), .ZN(
        n18379) );
  AOI22_X1 U21476 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n18385), .B1(
        n18660), .B2(n18445), .ZN(n18378) );
  OAI211_X1 U21477 ( .C1(n18549), .C2(n18382), .A(n18379), .B(n18378), .ZN(
        P3_U2913) );
  AOI22_X1 U21478 ( .A1(n18550), .A2(n18407), .B1(n18664), .B2(n18383), .ZN(
        n18381) );
  AOI22_X1 U21479 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n18385), .B1(
        n18666), .B2(n18445), .ZN(n18380) );
  OAI211_X1 U21480 ( .C1(n18553), .C2(n18382), .A(n18381), .B(n18380), .ZN(
        P3_U2914) );
  AOI22_X1 U21481 ( .A1(n18673), .A2(n18384), .B1(n18671), .B2(n18383), .ZN(
        n18387) );
  AOI22_X1 U21482 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n18385), .B1(
        n18674), .B2(n18445), .ZN(n18386) );
  OAI211_X1 U21483 ( .C1(n18679), .C2(n18405), .A(n18387), .B(n18386), .ZN(
        P3_U2915) );
  NAND2_X1 U21484 ( .A1(n18412), .A2(n18481), .ZN(n18475) );
  INV_X1 U21485 ( .A(n18475), .ZN(n18477) );
  NOR2_X1 U21486 ( .A1(n18445), .A2(n18477), .ZN(n18435) );
  NOR2_X1 U21487 ( .A1(n18745), .A2(n18435), .ZN(n18406) );
  AOI22_X1 U21488 ( .A1(n18589), .A2(n18430), .B1(n18622), .B2(n18406), .ZN(
        n18392) );
  INV_X1 U21489 ( .A(n18435), .ZN(n18390) );
  INV_X1 U21490 ( .A(n18388), .ZN(n18389) );
  OAI221_X1 U21491 ( .B1(n18390), .B2(n18593), .C1(n18390), .C2(n18389), .A(
        n18591), .ZN(n18408) );
  AOI22_X1 U21492 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n18408), .B1(
        n18621), .B2(n18407), .ZN(n18391) );
  OAI211_X1 U21493 ( .C1(n18597), .C2(n18475), .A(n18392), .B(n18391), .ZN(
        P3_U2916) );
  AOI22_X1 U21494 ( .A1(n18598), .A2(n18430), .B1(n18631), .B2(n18406), .ZN(
        n18394) );
  AOI22_X1 U21495 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n18408), .B1(
        n18633), .B2(n18477), .ZN(n18393) );
  OAI211_X1 U21496 ( .C1(n18601), .C2(n18405), .A(n18394), .B(n18393), .ZN(
        P3_U2917) );
  AOI22_X1 U21497 ( .A1(n18639), .A2(n18430), .B1(n18637), .B2(n18406), .ZN(
        n18396) );
  AOI22_X1 U21498 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n18408), .B1(
        n18569), .B2(n18477), .ZN(n18395) );
  OAI211_X1 U21499 ( .C1(n18572), .C2(n18405), .A(n18396), .B(n18395), .ZN(
        P3_U2918) );
  AOI22_X1 U21500 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n18408), .B1(
        n18644), .B2(n18406), .ZN(n18398) );
  AOI22_X1 U21501 ( .A1(n18573), .A2(n18407), .B1(n18646), .B2(n18477), .ZN(
        n18397) );
  OAI211_X1 U21502 ( .C1(n18576), .C2(n18426), .A(n18398), .B(n18397), .ZN(
        P3_U2919) );
  AOI22_X1 U21503 ( .A1(n18650), .A2(n18406), .B1(n18542), .B2(n18407), .ZN(
        n18400) );
  AOI22_X1 U21504 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n18408), .B1(
        n18653), .B2(n18477), .ZN(n18399) );
  OAI211_X1 U21505 ( .C1(n18545), .C2(n18426), .A(n18400), .B(n18399), .ZN(
        P3_U2920) );
  AOI22_X1 U21506 ( .A1(n18659), .A2(n18407), .B1(n18658), .B2(n18406), .ZN(
        n18402) );
  AOI22_X1 U21507 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n18408), .B1(
        n18660), .B2(n18477), .ZN(n18401) );
  OAI211_X1 U21508 ( .C1(n18663), .C2(n18426), .A(n18402), .B(n18401), .ZN(
        P3_U2921) );
  AOI22_X1 U21509 ( .A1(n18550), .A2(n18430), .B1(n18664), .B2(n18406), .ZN(
        n18404) );
  AOI22_X1 U21510 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n18408), .B1(
        n18666), .B2(n18477), .ZN(n18403) );
  OAI211_X1 U21511 ( .C1(n18553), .C2(n18405), .A(n18404), .B(n18403), .ZN(
        P3_U2922) );
  AOI22_X1 U21512 ( .A1(n18673), .A2(n18407), .B1(n18671), .B2(n18406), .ZN(
        n18410) );
  AOI22_X1 U21513 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n18408), .B1(
        n18674), .B2(n18477), .ZN(n18409) );
  OAI211_X1 U21514 ( .C1(n18679), .C2(n18426), .A(n18410), .B(n18409), .ZN(
        P3_U2923) );
  AOI22_X1 U21515 ( .A1(n18622), .A2(n18429), .B1(n18621), .B2(n18430), .ZN(
        n18415) );
  NAND2_X1 U21516 ( .A1(n18412), .A2(n18411), .ZN(n18431) );
  NOR2_X2 U21517 ( .A1(n18717), .A2(n18413), .ZN(n18493) );
  AOI22_X1 U21518 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n18431), .B1(
        n18627), .B2(n18493), .ZN(n18414) );
  OAI211_X1 U21519 ( .C1(n18630), .C2(n18456), .A(n18415), .B(n18414), .ZN(
        P3_U2924) );
  AOI22_X1 U21520 ( .A1(n18632), .A2(n18430), .B1(n18631), .B2(n18429), .ZN(
        n18417) );
  AOI22_X1 U21521 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n18431), .B1(
        n18633), .B2(n18493), .ZN(n18416) );
  OAI211_X1 U21522 ( .C1(n18636), .C2(n18456), .A(n18417), .B(n18416), .ZN(
        P3_U2925) );
  INV_X1 U21523 ( .A(n18493), .ZN(n18504) );
  AOI22_X1 U21524 ( .A1(n18638), .A2(n18430), .B1(n18637), .B2(n18429), .ZN(
        n18419) );
  AOI22_X1 U21525 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n18431), .B1(
        n18639), .B2(n18445), .ZN(n18418) );
  OAI211_X1 U21526 ( .C1(n18642), .C2(n18504), .A(n18419), .B(n18418), .ZN(
        P3_U2926) );
  AOI22_X1 U21527 ( .A1(n18573), .A2(n18430), .B1(n18644), .B2(n18429), .ZN(
        n18421) );
  AOI22_X1 U21528 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n18431), .B1(
        n18646), .B2(n18493), .ZN(n18420) );
  OAI211_X1 U21529 ( .C1(n18576), .C2(n18456), .A(n18421), .B(n18420), .ZN(
        P3_U2927) );
  AOI22_X1 U21530 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n18431), .B1(
        n18650), .B2(n18429), .ZN(n18423) );
  AOI22_X1 U21531 ( .A1(n18653), .A2(n18493), .B1(n18542), .B2(n18430), .ZN(
        n18422) );
  OAI211_X1 U21532 ( .C1(n18545), .C2(n18456), .A(n18423), .B(n18422), .ZN(
        P3_U2928) );
  AOI22_X1 U21533 ( .A1(n18546), .A2(n18445), .B1(n18658), .B2(n18429), .ZN(
        n18425) );
  AOI22_X1 U21534 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n18431), .B1(
        n18660), .B2(n18493), .ZN(n18424) );
  OAI211_X1 U21535 ( .C1(n18549), .C2(n18426), .A(n18425), .B(n18424), .ZN(
        P3_U2929) );
  AOI22_X1 U21536 ( .A1(n18665), .A2(n18430), .B1(n18664), .B2(n18429), .ZN(
        n18428) );
  AOI22_X1 U21537 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n18431), .B1(
        n18666), .B2(n18493), .ZN(n18427) );
  OAI211_X1 U21538 ( .C1(n18669), .C2(n18456), .A(n18428), .B(n18427), .ZN(
        P3_U2930) );
  AOI22_X1 U21539 ( .A1(n18673), .A2(n18430), .B1(n18671), .B2(n18429), .ZN(
        n18433) );
  AOI22_X1 U21540 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n18431), .B1(
        n18674), .B2(n18493), .ZN(n18432) );
  OAI211_X1 U21541 ( .C1(n18679), .C2(n18456), .A(n18433), .B(n18432), .ZN(
        P3_U2931) );
  NAND2_X1 U21542 ( .A1(n18434), .A2(n18528), .ZN(n18517) );
  INV_X1 U21543 ( .A(n18593), .ZN(n18482) );
  NOR2_X1 U21544 ( .A1(n18493), .A2(n18523), .ZN(n18483) );
  OAI21_X1 U21545 ( .B1(n18435), .B2(n18482), .A(n18483), .ZN(n18436) );
  OAI211_X1 U21546 ( .C1(n18523), .C2(n18864), .A(n18532), .B(n18436), .ZN(
        n18453) );
  NOR2_X1 U21547 ( .A1(n18745), .A2(n18483), .ZN(n18452) );
  AOI22_X1 U21548 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n18453), .B1(
        n18622), .B2(n18452), .ZN(n18438) );
  AOI22_X1 U21549 ( .A1(n18589), .A2(n18477), .B1(n18621), .B2(n18445), .ZN(
        n18437) );
  OAI211_X1 U21550 ( .C1(n18597), .C2(n18517), .A(n18438), .B(n18437), .ZN(
        P3_U2932) );
  AOI22_X1 U21551 ( .A1(n18632), .A2(n18445), .B1(n18631), .B2(n18452), .ZN(
        n18440) );
  AOI22_X1 U21552 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n18453), .B1(
        n18633), .B2(n18523), .ZN(n18439) );
  OAI211_X1 U21553 ( .C1(n18636), .C2(n18475), .A(n18440), .B(n18439), .ZN(
        P3_U2933) );
  AOI22_X1 U21554 ( .A1(n18639), .A2(n18477), .B1(n18637), .B2(n18452), .ZN(
        n18442) );
  AOI22_X1 U21555 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n18453), .B1(
        n18569), .B2(n18523), .ZN(n18441) );
  OAI211_X1 U21556 ( .C1(n18572), .C2(n18456), .A(n18442), .B(n18441), .ZN(
        P3_U2934) );
  AOI22_X1 U21557 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n18453), .B1(
        n18644), .B2(n18452), .ZN(n18444) );
  AOI22_X1 U21558 ( .A1(n18573), .A2(n18445), .B1(n18646), .B2(n18523), .ZN(
        n18443) );
  OAI211_X1 U21559 ( .C1(n18576), .C2(n18475), .A(n18444), .B(n18443), .ZN(
        P3_U2935) );
  AOI22_X1 U21560 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n18453), .B1(
        n18650), .B2(n18452), .ZN(n18447) );
  AOI22_X1 U21561 ( .A1(n18653), .A2(n18523), .B1(n18542), .B2(n18445), .ZN(
        n18446) );
  OAI211_X1 U21562 ( .C1(n18545), .C2(n18475), .A(n18447), .B(n18446), .ZN(
        P3_U2936) );
  AOI22_X1 U21563 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n18453), .B1(
        n18658), .B2(n18452), .ZN(n18449) );
  AOI22_X1 U21564 ( .A1(n18546), .A2(n18477), .B1(n18660), .B2(n18523), .ZN(
        n18448) );
  OAI211_X1 U21565 ( .C1(n18549), .C2(n18456), .A(n18449), .B(n18448), .ZN(
        P3_U2937) );
  AOI22_X1 U21566 ( .A1(n18550), .A2(n18477), .B1(n18664), .B2(n18452), .ZN(
        n18451) );
  AOI22_X1 U21567 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n18453), .B1(
        n18666), .B2(n18523), .ZN(n18450) );
  OAI211_X1 U21568 ( .C1(n18553), .C2(n18456), .A(n18451), .B(n18450), .ZN(
        P3_U2938) );
  AOI22_X1 U21569 ( .A1(n18555), .A2(n18477), .B1(n18671), .B2(n18452), .ZN(
        n18455) );
  AOI22_X1 U21570 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n18453), .B1(
        n18674), .B2(n18523), .ZN(n18454) );
  OAI211_X1 U21571 ( .C1(n18560), .C2(n18456), .A(n18455), .B(n18454), .ZN(
        P3_U2939) );
  NAND2_X1 U21572 ( .A1(n18528), .A2(n18457), .ZN(n18559) );
  INV_X1 U21573 ( .A(n18528), .ZN(n18506) );
  NOR2_X1 U21574 ( .A1(n18506), .A2(n18458), .ZN(n18476) );
  AOI22_X1 U21575 ( .A1(n18589), .A2(n18493), .B1(n18622), .B2(n18476), .ZN(
        n18462) );
  NOR2_X1 U21576 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18459), .ZN(
        n18460) );
  AOI22_X1 U21577 ( .A1(n18626), .A2(n18460), .B1(n18528), .B2(n18562), .ZN(
        n18478) );
  AOI22_X1 U21578 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n18478), .B1(
        n18621), .B2(n18477), .ZN(n18461) );
  OAI211_X1 U21579 ( .C1(n18597), .C2(n18559), .A(n18462), .B(n18461), .ZN(
        P3_U2940) );
  AOI22_X1 U21580 ( .A1(n18598), .A2(n18493), .B1(n18631), .B2(n18476), .ZN(
        n18464) );
  INV_X1 U21581 ( .A(n18559), .ZN(n18541) );
  AOI22_X1 U21582 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n18478), .B1(
        n18633), .B2(n18541), .ZN(n18463) );
  OAI211_X1 U21583 ( .C1(n18601), .C2(n18475), .A(n18464), .B(n18463), .ZN(
        P3_U2941) );
  AOI22_X1 U21584 ( .A1(n18639), .A2(n18493), .B1(n18637), .B2(n18476), .ZN(
        n18466) );
  AOI22_X1 U21585 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n18478), .B1(
        n18569), .B2(n18541), .ZN(n18465) );
  OAI211_X1 U21586 ( .C1(n18572), .C2(n18475), .A(n18466), .B(n18465), .ZN(
        P3_U2942) );
  AOI22_X1 U21587 ( .A1(n18644), .A2(n18476), .B1(n18645), .B2(n18493), .ZN(
        n18468) );
  AOI22_X1 U21588 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n18478), .B1(
        n18646), .B2(n18541), .ZN(n18467) );
  OAI211_X1 U21589 ( .C1(n18649), .C2(n18475), .A(n18468), .B(n18467), .ZN(
        P3_U2943) );
  AOI22_X1 U21590 ( .A1(n18651), .A2(n18493), .B1(n18650), .B2(n18476), .ZN(
        n18470) );
  AOI22_X1 U21591 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n18478), .B1(
        n18653), .B2(n18541), .ZN(n18469) );
  OAI211_X1 U21592 ( .C1(n18657), .C2(n18475), .A(n18470), .B(n18469), .ZN(
        P3_U2944) );
  AOI22_X1 U21593 ( .A1(n18546), .A2(n18493), .B1(n18658), .B2(n18476), .ZN(
        n18472) );
  AOI22_X1 U21594 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n18478), .B1(
        n18660), .B2(n18541), .ZN(n18471) );
  OAI211_X1 U21595 ( .C1(n18549), .C2(n18475), .A(n18472), .B(n18471), .ZN(
        P3_U2945) );
  AOI22_X1 U21596 ( .A1(n18550), .A2(n18493), .B1(n18664), .B2(n18476), .ZN(
        n18474) );
  AOI22_X1 U21597 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n18478), .B1(
        n18666), .B2(n18541), .ZN(n18473) );
  OAI211_X1 U21598 ( .C1(n18553), .C2(n18475), .A(n18474), .B(n18473), .ZN(
        P3_U2946) );
  AOI22_X1 U21599 ( .A1(n18673), .A2(n18477), .B1(n18671), .B2(n18476), .ZN(
        n18480) );
  AOI22_X1 U21600 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n18478), .B1(
        n18674), .B2(n18541), .ZN(n18479) );
  OAI211_X1 U21601 ( .C1(n18679), .C2(n18504), .A(n18480), .B(n18479), .ZN(
        P3_U2947) );
  NAND2_X1 U21602 ( .A1(n18528), .A2(n18481), .ZN(n18579) );
  AOI21_X1 U21603 ( .B1(n18559), .B2(n18579), .A(n18745), .ZN(n18500) );
  AOI22_X1 U21604 ( .A1(n18622), .A2(n18500), .B1(n18621), .B2(n18493), .ZN(
        n18486) );
  OAI211_X1 U21605 ( .C1(n18483), .C2(n18482), .A(n18559), .B(n18579), .ZN(
        n18484) );
  NAND2_X1 U21606 ( .A1(n18591), .A2(n18484), .ZN(n18501) );
  AOI22_X1 U21607 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n18501), .B1(
        n18589), .B2(n18523), .ZN(n18485) );
  OAI211_X1 U21608 ( .C1(n18597), .C2(n18579), .A(n18486), .B(n18485), .ZN(
        P3_U2948) );
  AOI22_X1 U21609 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n18501), .B1(
        n18631), .B2(n18500), .ZN(n18488) );
  INV_X1 U21610 ( .A(n18579), .ZN(n18585) );
  AOI22_X1 U21611 ( .A1(n18632), .A2(n18493), .B1(n18633), .B2(n18585), .ZN(
        n18487) );
  OAI211_X1 U21612 ( .C1(n18636), .C2(n18517), .A(n18488), .B(n18487), .ZN(
        P3_U2949) );
  AOI22_X1 U21613 ( .A1(n18639), .A2(n18523), .B1(n18637), .B2(n18500), .ZN(
        n18490) );
  AOI22_X1 U21614 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n18501), .B1(
        n18569), .B2(n18585), .ZN(n18489) );
  OAI211_X1 U21615 ( .C1(n18572), .C2(n18504), .A(n18490), .B(n18489), .ZN(
        P3_U2950) );
  AOI22_X1 U21616 ( .A1(n18644), .A2(n18500), .B1(n18645), .B2(n18523), .ZN(
        n18492) );
  AOI22_X1 U21617 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n18501), .B1(
        n18646), .B2(n18585), .ZN(n18491) );
  OAI211_X1 U21618 ( .C1(n18649), .C2(n18504), .A(n18492), .B(n18491), .ZN(
        P3_U2951) );
  AOI22_X1 U21619 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n18501), .B1(
        n18650), .B2(n18500), .ZN(n18495) );
  AOI22_X1 U21620 ( .A1(n18653), .A2(n18585), .B1(n18542), .B2(n18493), .ZN(
        n18494) );
  OAI211_X1 U21621 ( .C1(n18545), .C2(n18517), .A(n18495), .B(n18494), .ZN(
        P3_U2952) );
  AOI22_X1 U21622 ( .A1(n18546), .A2(n18523), .B1(n18658), .B2(n18500), .ZN(
        n18497) );
  AOI22_X1 U21623 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n18501), .B1(
        n18660), .B2(n18585), .ZN(n18496) );
  OAI211_X1 U21624 ( .C1(n18549), .C2(n18504), .A(n18497), .B(n18496), .ZN(
        P3_U2953) );
  AOI22_X1 U21625 ( .A1(n18550), .A2(n18523), .B1(n18664), .B2(n18500), .ZN(
        n18499) );
  AOI22_X1 U21626 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n18501), .B1(
        n18666), .B2(n18585), .ZN(n18498) );
  OAI211_X1 U21627 ( .C1(n18553), .C2(n18504), .A(n18499), .B(n18498), .ZN(
        P3_U2954) );
  AOI22_X1 U21628 ( .A1(n18555), .A2(n18523), .B1(n18671), .B2(n18500), .ZN(
        n18503) );
  AOI22_X1 U21629 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n18501), .B1(
        n18674), .B2(n18585), .ZN(n18502) );
  OAI211_X1 U21630 ( .C1(n18560), .C2(n18504), .A(n18503), .B(n18502), .ZN(
        P3_U2955) );
  NAND2_X1 U21631 ( .A1(n18505), .A2(n18528), .ZN(n18609) );
  NOR2_X1 U21632 ( .A1(n18718), .A2(n18506), .ZN(n18564) );
  AND2_X1 U21633 ( .A1(n18620), .A2(n18564), .ZN(n18522) );
  AOI22_X1 U21634 ( .A1(n18589), .A2(n18541), .B1(n18622), .B2(n18522), .ZN(
        n18508) );
  OAI211_X1 U21635 ( .C1(n18626), .C2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(
        n18624), .B(n18528), .ZN(n18524) );
  AOI22_X1 U21636 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n18524), .B1(
        n18621), .B2(n18523), .ZN(n18507) );
  OAI211_X1 U21637 ( .C1(n18597), .C2(n18609), .A(n18508), .B(n18507), .ZN(
        P3_U2956) );
  AOI22_X1 U21638 ( .A1(n18598), .A2(n18541), .B1(n18631), .B2(n18522), .ZN(
        n18510) );
  INV_X1 U21639 ( .A(n18609), .ZN(n18615) );
  AOI22_X1 U21640 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n18524), .B1(
        n18633), .B2(n18615), .ZN(n18509) );
  OAI211_X1 U21641 ( .C1(n18601), .C2(n18517), .A(n18510), .B(n18509), .ZN(
        P3_U2957) );
  AOI22_X1 U21642 ( .A1(n18639), .A2(n18541), .B1(n18637), .B2(n18522), .ZN(
        n18512) );
  AOI22_X1 U21643 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n18524), .B1(
        n18569), .B2(n18615), .ZN(n18511) );
  OAI211_X1 U21644 ( .C1(n18572), .C2(n18517), .A(n18512), .B(n18511), .ZN(
        P3_U2958) );
  AOI22_X1 U21645 ( .A1(n18573), .A2(n18523), .B1(n18644), .B2(n18522), .ZN(
        n18514) );
  AOI22_X1 U21646 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n18524), .B1(
        n18646), .B2(n18615), .ZN(n18513) );
  OAI211_X1 U21647 ( .C1(n18576), .C2(n18559), .A(n18514), .B(n18513), .ZN(
        P3_U2959) );
  AOI22_X1 U21648 ( .A1(n18651), .A2(n18541), .B1(n18650), .B2(n18522), .ZN(
        n18516) );
  AOI22_X1 U21649 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n18524), .B1(
        n18653), .B2(n18615), .ZN(n18515) );
  OAI211_X1 U21650 ( .C1(n18657), .C2(n18517), .A(n18516), .B(n18515), .ZN(
        P3_U2960) );
  AOI22_X1 U21651 ( .A1(n18659), .A2(n18523), .B1(n18658), .B2(n18522), .ZN(
        n18519) );
  AOI22_X1 U21652 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n18524), .B1(
        n18660), .B2(n18615), .ZN(n18518) );
  OAI211_X1 U21653 ( .C1(n18663), .C2(n18559), .A(n18519), .B(n18518), .ZN(
        P3_U2961) );
  AOI22_X1 U21654 ( .A1(n18665), .A2(n18523), .B1(n18664), .B2(n18522), .ZN(
        n18521) );
  AOI22_X1 U21655 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n18524), .B1(
        n18666), .B2(n18615), .ZN(n18520) );
  OAI211_X1 U21656 ( .C1(n18669), .C2(n18559), .A(n18521), .B(n18520), .ZN(
        P3_U2962) );
  AOI22_X1 U21657 ( .A1(n18673), .A2(n18523), .B1(n18671), .B2(n18522), .ZN(
        n18526) );
  AOI22_X1 U21658 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n18524), .B1(
        n18674), .B2(n18615), .ZN(n18525) );
  OAI211_X1 U21659 ( .C1(n18679), .C2(n18559), .A(n18526), .B(n18525), .ZN(
        P3_U2963) );
  INV_X1 U21660 ( .A(n18561), .ZN(n18625) );
  NAND2_X1 U21661 ( .A1(n18625), .A2(n18527), .ZN(n18656) );
  INV_X1 U21662 ( .A(n18656), .ZN(n18672) );
  NOR2_X1 U21663 ( .A1(n18615), .A2(n18672), .ZN(n18590) );
  NOR2_X1 U21664 ( .A1(n18745), .A2(n18590), .ZN(n18554) );
  AOI22_X1 U21665 ( .A1(n18589), .A2(n18585), .B1(n18622), .B2(n18554), .ZN(
        n18534) );
  NAND2_X1 U21666 ( .A1(n18593), .A2(n18528), .ZN(n18529) );
  OAI21_X1 U21667 ( .B1(n18530), .B2(n18529), .A(n18590), .ZN(n18531) );
  OAI211_X1 U21668 ( .C1(n18672), .C2(n18864), .A(n18532), .B(n18531), .ZN(
        n18556) );
  AOI22_X1 U21669 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n18556), .B1(
        n18621), .B2(n18541), .ZN(n18533) );
  OAI211_X1 U21670 ( .C1(n18597), .C2(n18656), .A(n18534), .B(n18533), .ZN(
        P3_U2964) );
  AOI22_X1 U21671 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n18556), .B1(
        n18631), .B2(n18554), .ZN(n18536) );
  AOI22_X1 U21672 ( .A1(n18633), .A2(n18672), .B1(n18598), .B2(n18585), .ZN(
        n18535) );
  OAI211_X1 U21673 ( .C1(n18601), .C2(n18559), .A(n18536), .B(n18535), .ZN(
        P3_U2965) );
  AOI22_X1 U21674 ( .A1(n18639), .A2(n18585), .B1(n18637), .B2(n18554), .ZN(
        n18538) );
  AOI22_X1 U21675 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n18556), .B1(
        n18569), .B2(n18672), .ZN(n18537) );
  OAI211_X1 U21676 ( .C1(n18572), .C2(n18559), .A(n18538), .B(n18537), .ZN(
        P3_U2966) );
  AOI22_X1 U21677 ( .A1(n18644), .A2(n18554), .B1(n18645), .B2(n18585), .ZN(
        n18540) );
  AOI22_X1 U21678 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n18556), .B1(
        n18646), .B2(n18672), .ZN(n18539) );
  OAI211_X1 U21679 ( .C1(n18649), .C2(n18559), .A(n18540), .B(n18539), .ZN(
        P3_U2967) );
  AOI22_X1 U21680 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n18556), .B1(
        n18650), .B2(n18554), .ZN(n18544) );
  AOI22_X1 U21681 ( .A1(n18653), .A2(n18672), .B1(n18542), .B2(n18541), .ZN(
        n18543) );
  OAI211_X1 U21682 ( .C1(n18545), .C2(n18579), .A(n18544), .B(n18543), .ZN(
        P3_U2968) );
  AOI22_X1 U21683 ( .A1(n18546), .A2(n18585), .B1(n18658), .B2(n18554), .ZN(
        n18548) );
  AOI22_X1 U21684 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n18556), .B1(
        n18660), .B2(n18672), .ZN(n18547) );
  OAI211_X1 U21685 ( .C1(n18549), .C2(n18559), .A(n18548), .B(n18547), .ZN(
        P3_U2969) );
  AOI22_X1 U21686 ( .A1(n18550), .A2(n18585), .B1(n18664), .B2(n18554), .ZN(
        n18552) );
  AOI22_X1 U21687 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n18556), .B1(
        n18666), .B2(n18672), .ZN(n18551) );
  OAI211_X1 U21688 ( .C1(n18553), .C2(n18559), .A(n18552), .B(n18551), .ZN(
        P3_U2970) );
  AOI22_X1 U21689 ( .A1(n18555), .A2(n18585), .B1(n18671), .B2(n18554), .ZN(
        n18558) );
  AOI22_X1 U21690 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n18556), .B1(
        n18674), .B2(n18672), .ZN(n18557) );
  OAI211_X1 U21691 ( .C1(n18560), .C2(n18559), .A(n18558), .B(n18557), .ZN(
        P3_U2971) );
  NOR2_X1 U21692 ( .A1(n18745), .A2(n18561), .ZN(n18584) );
  AOI22_X1 U21693 ( .A1(n18589), .A2(n18615), .B1(n18622), .B2(n18584), .ZN(
        n18566) );
  AOI22_X1 U21694 ( .A1(n18626), .A2(n18564), .B1(n18563), .B2(n18562), .ZN(
        n18586) );
  AOI22_X1 U21695 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n18586), .B1(
        n18621), .B2(n18585), .ZN(n18565) );
  OAI211_X1 U21696 ( .C1(n18597), .C2(n18680), .A(n18566), .B(n18565), .ZN(
        P3_U2972) );
  AOI22_X1 U21697 ( .A1(n18632), .A2(n18585), .B1(n18631), .B2(n18584), .ZN(
        n18568) );
  AOI22_X1 U21698 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n18586), .B1(
        n18652), .B2(n18633), .ZN(n18567) );
  OAI211_X1 U21699 ( .C1(n18636), .C2(n18609), .A(n18568), .B(n18567), .ZN(
        P3_U2973) );
  AOI22_X1 U21700 ( .A1(n18639), .A2(n18615), .B1(n18637), .B2(n18584), .ZN(
        n18571) );
  AOI22_X1 U21701 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n18586), .B1(
        n18652), .B2(n18569), .ZN(n18570) );
  OAI211_X1 U21702 ( .C1(n18572), .C2(n18579), .A(n18571), .B(n18570), .ZN(
        P3_U2974) );
  AOI22_X1 U21703 ( .A1(n18573), .A2(n18585), .B1(n18644), .B2(n18584), .ZN(
        n18575) );
  AOI22_X1 U21704 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n18586), .B1(
        n18652), .B2(n18646), .ZN(n18574) );
  OAI211_X1 U21705 ( .C1(n18576), .C2(n18609), .A(n18575), .B(n18574), .ZN(
        P3_U2975) );
  AOI22_X1 U21706 ( .A1(n18651), .A2(n18615), .B1(n18650), .B2(n18584), .ZN(
        n18578) );
  AOI22_X1 U21707 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n18586), .B1(
        n18652), .B2(n18653), .ZN(n18577) );
  OAI211_X1 U21708 ( .C1(n18657), .C2(n18579), .A(n18578), .B(n18577), .ZN(
        P3_U2976) );
  AOI22_X1 U21709 ( .A1(n18659), .A2(n18585), .B1(n18658), .B2(n18584), .ZN(
        n18581) );
  AOI22_X1 U21710 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n18586), .B1(
        n18652), .B2(n18660), .ZN(n18580) );
  OAI211_X1 U21711 ( .C1(n18663), .C2(n18609), .A(n18581), .B(n18580), .ZN(
        P3_U2977) );
  AOI22_X1 U21712 ( .A1(n18665), .A2(n18585), .B1(n18664), .B2(n18584), .ZN(
        n18583) );
  AOI22_X1 U21713 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n18586), .B1(
        n18652), .B2(n18666), .ZN(n18582) );
  OAI211_X1 U21714 ( .C1(n18669), .C2(n18609), .A(n18583), .B(n18582), .ZN(
        P3_U2978) );
  AOI22_X1 U21715 ( .A1(n18673), .A2(n18585), .B1(n18671), .B2(n18584), .ZN(
        n18588) );
  AOI22_X1 U21716 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n18586), .B1(
        n18652), .B2(n18674), .ZN(n18587) );
  OAI211_X1 U21717 ( .C1(n18679), .C2(n18609), .A(n18588), .B(n18587), .ZN(
        P3_U2979) );
  AND2_X1 U21718 ( .A1(n18620), .A2(n18594), .ZN(n18614) );
  AOI22_X1 U21719 ( .A1(n18589), .A2(n18672), .B1(n18622), .B2(n18614), .ZN(
        n18596) );
  INV_X1 U21720 ( .A(n18590), .ZN(n18592) );
  OAI221_X1 U21721 ( .B1(n18594), .B2(n18593), .C1(n18594), .C2(n18592), .A(
        n18591), .ZN(n18617) );
  AOI22_X1 U21722 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n18617), .B1(
        n18621), .B2(n18615), .ZN(n18595) );
  OAI211_X1 U21723 ( .C1(n18604), .C2(n18597), .A(n18596), .B(n18595), .ZN(
        P3_U2980) );
  AOI22_X1 U21724 ( .A1(n18598), .A2(n18672), .B1(n18631), .B2(n18614), .ZN(
        n18600) );
  AOI22_X1 U21725 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n18617), .B1(
        n18616), .B2(n18633), .ZN(n18599) );
  OAI211_X1 U21726 ( .C1(n18601), .C2(n18609), .A(n18600), .B(n18599), .ZN(
        P3_U2981) );
  AOI22_X1 U21727 ( .A1(n18638), .A2(n18615), .B1(n18637), .B2(n18614), .ZN(
        n18603) );
  AOI22_X1 U21728 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n18617), .B1(
        n18639), .B2(n18672), .ZN(n18602) );
  OAI211_X1 U21729 ( .C1(n18604), .C2(n18642), .A(n18603), .B(n18602), .ZN(
        P3_U2982) );
  AOI22_X1 U21730 ( .A1(n18644), .A2(n18614), .B1(n18645), .B2(n18672), .ZN(
        n18606) );
  AOI22_X1 U21731 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n18617), .B1(
        n18616), .B2(n18646), .ZN(n18605) );
  OAI211_X1 U21732 ( .C1(n18649), .C2(n18609), .A(n18606), .B(n18605), .ZN(
        P3_U2983) );
  AOI22_X1 U21733 ( .A1(n18651), .A2(n18672), .B1(n18650), .B2(n18614), .ZN(
        n18608) );
  AOI22_X1 U21734 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n18617), .B1(
        n18616), .B2(n18653), .ZN(n18607) );
  OAI211_X1 U21735 ( .C1(n18657), .C2(n18609), .A(n18608), .B(n18607), .ZN(
        P3_U2984) );
  AOI22_X1 U21736 ( .A1(n18659), .A2(n18615), .B1(n18658), .B2(n18614), .ZN(
        n18611) );
  AOI22_X1 U21737 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n18617), .B1(
        n18616), .B2(n18660), .ZN(n18610) );
  OAI211_X1 U21738 ( .C1(n18663), .C2(n18656), .A(n18611), .B(n18610), .ZN(
        P3_U2985) );
  AOI22_X1 U21739 ( .A1(n18665), .A2(n18615), .B1(n18664), .B2(n18614), .ZN(
        n18613) );
  AOI22_X1 U21740 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n18617), .B1(
        n18616), .B2(n18666), .ZN(n18612) );
  OAI211_X1 U21741 ( .C1(n18669), .C2(n18656), .A(n18613), .B(n18612), .ZN(
        P3_U2986) );
  AOI22_X1 U21742 ( .A1(n18673), .A2(n18615), .B1(n18671), .B2(n18614), .ZN(
        n18619) );
  AOI22_X1 U21743 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n18617), .B1(
        n18616), .B2(n18674), .ZN(n18618) );
  OAI211_X1 U21744 ( .C1(n18679), .C2(n18656), .A(n18619), .B(n18618), .ZN(
        P3_U2987) );
  AND2_X1 U21745 ( .A1(n18620), .A2(n18623), .ZN(n18670) );
  AOI22_X1 U21746 ( .A1(n18622), .A2(n18670), .B1(n18621), .B2(n18672), .ZN(
        n18629) );
  AOI22_X1 U21747 ( .A1(n18626), .A2(n18625), .B1(n18624), .B2(n18623), .ZN(
        n18676) );
  AOI22_X1 U21748 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n18676), .B1(
        n18675), .B2(n18627), .ZN(n18628) );
  OAI211_X1 U21749 ( .C1(n18630), .C2(n18680), .A(n18629), .B(n18628), .ZN(
        P3_U2988) );
  AOI22_X1 U21750 ( .A1(n18632), .A2(n18672), .B1(n18631), .B2(n18670), .ZN(
        n18635) );
  AOI22_X1 U21751 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n18676), .B1(
        n18675), .B2(n18633), .ZN(n18634) );
  OAI211_X1 U21752 ( .C1(n18680), .C2(n18636), .A(n18635), .B(n18634), .ZN(
        P3_U2989) );
  AOI22_X1 U21753 ( .A1(n18638), .A2(n18672), .B1(n18637), .B2(n18670), .ZN(
        n18641) );
  AOI22_X1 U21754 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n18676), .B1(
        n18652), .B2(n18639), .ZN(n18640) );
  OAI211_X1 U21755 ( .C1(n18643), .C2(n18642), .A(n18641), .B(n18640), .ZN(
        P3_U2990) );
  AOI22_X1 U21756 ( .A1(n18652), .A2(n18645), .B1(n18644), .B2(n18670), .ZN(
        n18648) );
  AOI22_X1 U21757 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n18676), .B1(
        n18675), .B2(n18646), .ZN(n18647) );
  OAI211_X1 U21758 ( .C1(n18649), .C2(n18656), .A(n18648), .B(n18647), .ZN(
        P3_U2991) );
  AOI22_X1 U21759 ( .A1(n18652), .A2(n18651), .B1(n18650), .B2(n18670), .ZN(
        n18655) );
  AOI22_X1 U21760 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n18676), .B1(
        n18675), .B2(n18653), .ZN(n18654) );
  OAI211_X1 U21761 ( .C1(n18657), .C2(n18656), .A(n18655), .B(n18654), .ZN(
        P3_U2992) );
  AOI22_X1 U21762 ( .A1(n18659), .A2(n18672), .B1(n18658), .B2(n18670), .ZN(
        n18662) );
  AOI22_X1 U21763 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n18676), .B1(
        n18675), .B2(n18660), .ZN(n18661) );
  OAI211_X1 U21764 ( .C1(n18680), .C2(n18663), .A(n18662), .B(n18661), .ZN(
        P3_U2993) );
  AOI22_X1 U21765 ( .A1(n18665), .A2(n18672), .B1(n18664), .B2(n18670), .ZN(
        n18668) );
  AOI22_X1 U21766 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n18676), .B1(
        n18675), .B2(n18666), .ZN(n18667) );
  OAI211_X1 U21767 ( .C1(n18680), .C2(n18669), .A(n18668), .B(n18667), .ZN(
        P3_U2994) );
  AOI22_X1 U21768 ( .A1(n18673), .A2(n18672), .B1(n18671), .B2(n18670), .ZN(
        n18678) );
  AOI22_X1 U21769 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n18676), .B1(
        n18675), .B2(n18674), .ZN(n18677) );
  OAI211_X1 U21770 ( .C1(n18680), .C2(n18679), .A(n18678), .B(n18677), .ZN(
        P3_U2995) );
  NOR2_X1 U21771 ( .A1(n18710), .A2(n18681), .ZN(n18683) );
  OAI222_X1 U21772 ( .A1(n18687), .A2(n18686), .B1(n18685), .B2(n18684), .C1(
        n18683), .C2(n18682), .ZN(n18879) );
  OAI21_X1 U21773 ( .B1(P3_FLUSH_REG_SCAN_IN), .B2(P3_MORE_REG_SCAN_IN), .A(
        n18688), .ZN(n18689) );
  OAI211_X1 U21774 ( .C1(n18691), .C2(n18711), .A(n18690), .B(n18689), .ZN(
        n18732) );
  OAI21_X1 U21775 ( .B1(n18692), .B2(n18870), .A(n18714), .ZN(n18703) );
  AOI22_X1 U21776 ( .A1(n18704), .A2(n18703), .B1(n18710), .B2(n18696), .ZN(
        n18839) );
  NOR2_X1 U21777 ( .A1(n18721), .A2(n18839), .ZN(n18702) );
  AOI21_X1 U21778 ( .B1(n18695), .B2(n18694), .A(n18693), .ZN(n18706) );
  OAI21_X1 U21779 ( .B1(n18697), .B2(n18706), .A(n18696), .ZN(n18698) );
  AOI21_X1 U21780 ( .B1(n18700), .B2(n18699), .A(n18698), .ZN(n18842) );
  NAND2_X1 U21781 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n18842), .ZN(
        n18701) );
  OAI22_X1 U21782 ( .A1(n18702), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n18721), .B2(n18701), .ZN(n18730) );
  INV_X1 U21783 ( .A(n18703), .ZN(n18715) );
  AOI211_X1 U21784 ( .C1(n18854), .C2(n18862), .A(n18704), .B(n18715), .ZN(
        n18709) );
  INV_X1 U21785 ( .A(n18705), .ZN(n18707) );
  NOR3_X1 U21786 ( .A1(n18707), .A2(n18706), .A3(n18854), .ZN(n18708) );
  AOI211_X1 U21787 ( .C1(n18710), .C2(n18847), .A(n18709), .B(n18708), .ZN(
        n18850) );
  AOI22_X1 U21788 ( .A1(n18721), .A2(n18854), .B1(n18850), .B2(n18711), .ZN(
        n18725) );
  NOR2_X1 U21789 ( .A1(n18713), .A2(n18712), .ZN(n18716) );
  AOI22_X1 U21790 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18714), .B1(
        n18716), .B2(n18870), .ZN(n18865) );
  OAI22_X1 U21791 ( .A1(n18716), .A2(n18855), .B1(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n18715), .ZN(n18859) );
  AOI222_X1 U21792 ( .A1(n18865), .A2(n18859), .B1(n18865), .B2(n18718), .C1(
        n18859), .C2(n18717), .ZN(n18720) );
  OAI21_X1 U21793 ( .B1(n18721), .B2(n18720), .A(n18719), .ZN(n18724) );
  AND2_X1 U21794 ( .A1(n18725), .A2(n18724), .ZN(n18722) );
  OAI221_X1 U21795 ( .B1(n18725), .B2(n18724), .C1(n18723), .C2(n18722), .A(
        n18727), .ZN(n18729) );
  AOI21_X1 U21796 ( .B1(n18727), .B2(n18726), .A(n18725), .ZN(n18728) );
  AOI222_X1 U21797 ( .A1(n18730), .A2(n18729), .B1(n18730), .B2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C1(n18729), .C2(n18728), .ZN(
        n18731) );
  NOR4_X1 U21798 ( .A1(n18733), .A2(n18879), .A3(n18732), .A4(n18731), .ZN(
        n18744) );
  NOR2_X1 U21799 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n18894) );
  AOI22_X1 U21800 ( .A1(n18866), .A2(n18894), .B1(n18889), .B2(n18881), .ZN(
        n18734) );
  INV_X1 U21801 ( .A(n18734), .ZN(n18739) );
  OAI211_X1 U21802 ( .C1(n18736), .C2(n18735), .A(n18884), .B(n18744), .ZN(
        n18837) );
  OAI21_X1 U21803 ( .B1(P3_STATE2_REG_2__SCAN_IN), .B2(n18880), .A(n18837), 
        .ZN(n18746) );
  NOR2_X1 U21804 ( .A1(n18737), .A2(n18746), .ZN(n18738) );
  MUX2_X1 U21805 ( .A(n18739), .B(n18738), .S(P3_STATE2_REG_0__SCAN_IN), .Z(
        n18742) );
  INV_X1 U21806 ( .A(n18740), .ZN(n18741) );
  OAI211_X1 U21807 ( .C1(n18744), .C2(n18743), .A(n18742), .B(n18741), .ZN(
        P3_U2996) );
  NAND2_X1 U21808 ( .A1(n18889), .A2(n18881), .ZN(n18749) );
  NAND4_X1 U21809 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(
        P3_STATE2_REG_1__SCAN_IN), .A3(n18889), .A4(n18901), .ZN(n18751) );
  OR3_X1 U21810 ( .A1(n18747), .A2(n18746), .A3(n18745), .ZN(n18748) );
  NAND4_X1 U21811 ( .A1(n18750), .A2(n18749), .A3(n18751), .A4(n18748), .ZN(
        P3_U2997) );
  INV_X1 U21812 ( .A(n18894), .ZN(n18753) );
  AND4_X1 U21813 ( .A1(n18753), .A2(n18752), .A3(n18751), .A4(n18836), .ZN(
        P3_U2998) );
  AND2_X1 U21814 ( .A1(P3_DATAWIDTH_REG_31__SCAN_IN), .A2(n18832), .ZN(
        P3_U2999) );
  AND2_X1 U21815 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n18832), .ZN(
        P3_U3000) );
  AND2_X1 U21816 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n18832), .ZN(
        P3_U3001) );
  AND2_X1 U21817 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n18832), .ZN(
        P3_U3002) );
  AND2_X1 U21818 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n18832), .ZN(
        P3_U3003) );
  AND2_X1 U21819 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n18832), .ZN(
        P3_U3004) );
  AND2_X1 U21820 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n18832), .ZN(
        P3_U3005) );
  AND2_X1 U21821 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n18832), .ZN(
        P3_U3006) );
  AND2_X1 U21822 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n18832), .ZN(
        P3_U3007) );
  AND2_X1 U21823 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n18832), .ZN(
        P3_U3008) );
  AND2_X1 U21824 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n18832), .ZN(
        P3_U3009) );
  AND2_X1 U21825 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n18832), .ZN(
        P3_U3010) );
  AND2_X1 U21826 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n18832), .ZN(
        P3_U3011) );
  AND2_X1 U21827 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n18832), .ZN(
        P3_U3012) );
  AND2_X1 U21828 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n18832), .ZN(
        P3_U3013) );
  AND2_X1 U21829 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n18832), .ZN(
        P3_U3014) );
  AND2_X1 U21830 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n18832), .ZN(
        P3_U3015) );
  AND2_X1 U21831 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n18832), .ZN(
        P3_U3016) );
  AND2_X1 U21832 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n18832), .ZN(
        P3_U3017) );
  AND2_X1 U21833 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n18832), .ZN(
        P3_U3018) );
  INV_X1 U21834 ( .A(P3_DATAWIDTH_REG_11__SCAN_IN), .ZN(n21107) );
  NOR2_X1 U21835 ( .A1(n21107), .A2(n18835), .ZN(P3_U3019) );
  AND2_X1 U21836 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n18832), .ZN(
        P3_U3020) );
  AND2_X1 U21837 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n18832), .ZN(P3_U3021) );
  AND2_X1 U21838 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n18832), .ZN(P3_U3022) );
  AND2_X1 U21839 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n18832), .ZN(P3_U3023) );
  AND2_X1 U21840 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n18832), .ZN(P3_U3024) );
  AND2_X1 U21841 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n18832), .ZN(P3_U3025) );
  AND2_X1 U21842 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n18832), .ZN(P3_U3026) );
  AND2_X1 U21843 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n18832), .ZN(P3_U3027) );
  AND2_X1 U21844 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n18832), .ZN(P3_U3028) );
  OAI21_X1 U21845 ( .B1(n18754), .B2(n19822), .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n18755) );
  AOI22_X1 U21846 ( .A1(n18767), .A2(n18769), .B1(n18899), .B2(n18755), .ZN(
        n18756) );
  NAND3_X1 U21847 ( .A1(NA), .A2(n18767), .A3(n18759), .ZN(n18762) );
  OAI211_X1 U21848 ( .C1(n18880), .C2(n18757), .A(n18756), .B(n18762), .ZN(
        P3_U3029) );
  INV_X1 U21849 ( .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n18896) );
  NOR2_X1 U21850 ( .A1(n18769), .A2(n19822), .ZN(n18765) );
  OAI22_X1 U21851 ( .A1(n18896), .A2(n18765), .B1(n19822), .B2(n18757), .ZN(
        n18758) );
  INV_X1 U21852 ( .A(n18758), .ZN(n18760) );
  NOR2_X1 U21853 ( .A1(n18880), .A2(n18759), .ZN(n18761) );
  INV_X1 U21854 ( .A(n18761), .ZN(n18763) );
  OAI211_X1 U21855 ( .C1(n18760), .C2(n18767), .A(n18763), .B(n18885), .ZN(
        P3_U3030) );
  AOI21_X1 U21856 ( .B1(n18767), .B2(n18762), .A(n18761), .ZN(n18768) );
  OAI22_X1 U21857 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(
        P3_REQUESTPENDING_REG_SCAN_IN), .B1(NA), .B2(n18763), .ZN(n18764) );
  OAI22_X1 U21858 ( .A1(n18765), .A2(n18764), .B1(
        P3_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .ZN(n18766) );
  OAI22_X1 U21859 ( .A1(n18768), .A2(n18769), .B1(n18767), .B2(n18766), .ZN(
        P3_U3031) );
  NAND2_X1 U21860 ( .A1(n18898), .A2(n18769), .ZN(n18821) );
  CLKBUF_X1 U21861 ( .A(n18821), .Z(n18822) );
  OAI222_X1 U21862 ( .A1(n20815), .A2(n18826), .B1(n18770), .B2(n18898), .C1(
        n18771), .C2(n18822), .ZN(P3_U3032) );
  OAI222_X1 U21863 ( .A1(n18822), .A2(n18773), .B1(n18772), .B2(n18898), .C1(
        n18771), .C2(n18826), .ZN(P3_U3033) );
  OAI222_X1 U21864 ( .A1(n18821), .A2(n18774), .B1(n21127), .B2(n18898), .C1(
        n18773), .C2(n18826), .ZN(P3_U3034) );
  INV_X1 U21865 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n18777) );
  OAI222_X1 U21866 ( .A1(n18821), .A2(n18777), .B1(n18775), .B2(n18898), .C1(
        n18774), .C2(n18826), .ZN(P3_U3035) );
  INV_X1 U21867 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n21023) );
  OAI222_X1 U21868 ( .A1(n18777), .A2(n18826), .B1(n18776), .B2(n18898), .C1(
        n21023), .C2(n18822), .ZN(P3_U3036) );
  OAI222_X1 U21869 ( .A1(n21023), .A2(n18826), .B1(n21077), .B2(n18898), .C1(
        n18778), .C2(n18822), .ZN(P3_U3037) );
  INV_X1 U21870 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n18781) );
  OAI222_X1 U21871 ( .A1(n18821), .A2(n18781), .B1(n18779), .B2(n18898), .C1(
        n18778), .C2(n18826), .ZN(P3_U3038) );
  INV_X1 U21872 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n18782) );
  OAI222_X1 U21873 ( .A1(n18781), .A2(n18826), .B1(n18780), .B2(n18898), .C1(
        n18782), .C2(n18822), .ZN(P3_U3039) );
  OAI222_X1 U21874 ( .A1(n18821), .A2(n18784), .B1(n18783), .B2(n18898), .C1(
        n18782), .C2(n18826), .ZN(P3_U3040) );
  OAI222_X1 U21875 ( .A1(n18821), .A2(n18786), .B1(n18785), .B2(n18898), .C1(
        n18784), .C2(n18826), .ZN(P3_U3041) );
  INV_X1 U21876 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n18789) );
  OAI222_X1 U21877 ( .A1(n18822), .A2(n18789), .B1(n18787), .B2(n18898), .C1(
        n18786), .C2(n18826), .ZN(P3_U3042) );
  OAI222_X1 U21878 ( .A1(n18789), .A2(n18826), .B1(n18788), .B2(n18898), .C1(
        n18790), .C2(n18822), .ZN(P3_U3043) );
  INV_X1 U21879 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n21144) );
  OAI222_X1 U21880 ( .A1(n18822), .A2(n21144), .B1(n18791), .B2(n18898), .C1(
        n18790), .C2(n18826), .ZN(P3_U3044) );
  OAI222_X1 U21881 ( .A1(n21144), .A2(n18826), .B1(n18792), .B2(n18898), .C1(
        n18793), .C2(n18822), .ZN(P3_U3045) );
  OAI222_X1 U21882 ( .A1(n18822), .A2(n20933), .B1(n18794), .B2(n18898), .C1(
        n18793), .C2(n18826), .ZN(P3_U3046) );
  INV_X1 U21883 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n18797) );
  OAI222_X1 U21884 ( .A1(n18822), .A2(n18797), .B1(n18795), .B2(n18898), .C1(
        n20933), .C2(n18826), .ZN(P3_U3047) );
  OAI222_X1 U21885 ( .A1(n18797), .A2(n18826), .B1(n18796), .B2(n18898), .C1(
        n18798), .C2(n18822), .ZN(P3_U3048) );
  OAI222_X1 U21886 ( .A1(n18822), .A2(n18800), .B1(n18799), .B2(n18898), .C1(
        n18798), .C2(n18826), .ZN(P3_U3049) );
  OAI222_X1 U21887 ( .A1(n18822), .A2(n18803), .B1(n18801), .B2(n18898), .C1(
        n18800), .C2(n18826), .ZN(P3_U3050) );
  OAI222_X1 U21888 ( .A1(n18803), .A2(n18826), .B1(n18802), .B2(n18898), .C1(
        n18804), .C2(n18822), .ZN(P3_U3051) );
  OAI222_X1 U21889 ( .A1(n18821), .A2(n18806), .B1(n18805), .B2(n18898), .C1(
        n18804), .C2(n18826), .ZN(P3_U3052) );
  INV_X1 U21890 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n18808) );
  OAI222_X1 U21891 ( .A1(n18821), .A2(n18808), .B1(n18807), .B2(n18898), .C1(
        n18806), .C2(n18826), .ZN(P3_U3053) );
  OAI222_X1 U21892 ( .A1(n18808), .A2(n18826), .B1(n21080), .B2(n18898), .C1(
        n18809), .C2(n18822), .ZN(P3_U3054) );
  OAI222_X1 U21893 ( .A1(n18821), .A2(n18811), .B1(n18810), .B2(n18898), .C1(
        n18809), .C2(n18826), .ZN(P3_U3055) );
  OAI222_X1 U21894 ( .A1(n18821), .A2(n18813), .B1(n18812), .B2(n18898), .C1(
        n18811), .C2(n18826), .ZN(P3_U3056) );
  OAI222_X1 U21895 ( .A1(n18821), .A2(n18815), .B1(n18814), .B2(n18898), .C1(
        n18813), .C2(n18826), .ZN(P3_U3057) );
  INV_X1 U21896 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n18818) );
  OAI222_X1 U21897 ( .A1(n18821), .A2(n18818), .B1(n18816), .B2(n18898), .C1(
        n18815), .C2(n18826), .ZN(P3_U3058) );
  OAI222_X1 U21898 ( .A1(n18818), .A2(n18826), .B1(n18817), .B2(n18898), .C1(
        n18819), .C2(n18822), .ZN(P3_U3059) );
  OAI222_X1 U21899 ( .A1(n18821), .A2(n18825), .B1(n18820), .B2(n18898), .C1(
        n18819), .C2(n18826), .ZN(P3_U3060) );
  OAI222_X1 U21900 ( .A1(n18826), .A2(n18825), .B1(n18824), .B2(n18898), .C1(
        n18823), .C2(n18822), .ZN(P3_U3061) );
  INV_X1 U21901 ( .A(P3_BE_N_REG_3__SCAN_IN), .ZN(n20967) );
  AOI22_X1 U21902 ( .A1(n18898), .A2(n18827), .B1(n20967), .B2(n18899), .ZN(
        P3_U3274) );
  INV_X1 U21903 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n18873) );
  INV_X1 U21904 ( .A(P3_BE_N_REG_2__SCAN_IN), .ZN(n18828) );
  AOI22_X1 U21905 ( .A1(n18898), .A2(n18873), .B1(n18828), .B2(n18899), .ZN(
        P3_U3275) );
  MUX2_X1 U21906 ( .A(P3_BE_N_REG_1__SCAN_IN), .B(P3_BYTEENABLE_REG_1__SCAN_IN), .S(n18898), .Z(P3_U3276) );
  INV_X1 U21907 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n18876) );
  INV_X1 U21908 ( .A(P3_BE_N_REG_0__SCAN_IN), .ZN(n18829) );
  AOI22_X1 U21909 ( .A1(n18898), .A2(n18876), .B1(n18829), .B2(n18899), .ZN(
        P3_U3277) );
  INV_X1 U21910 ( .A(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(n18831) );
  INV_X1 U21911 ( .A(n18833), .ZN(n18830) );
  AOI21_X1 U21912 ( .B1(n18832), .B2(n18831), .A(n18830), .ZN(P3_U3280) );
  OAI21_X1 U21913 ( .B1(n18835), .B2(n18834), .A(n18833), .ZN(P3_U3281) );
  OAI221_X1 U21914 ( .B1(n18864), .B2(P3_STATE2_REG_0__SCAN_IN), .C1(n18864), 
        .C2(n18837), .A(n18836), .ZN(P3_U3282) );
  INV_X1 U21915 ( .A(n18838), .ZN(n18841) );
  NOR3_X1 U21916 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n18839), .A3(
        n18849), .ZN(n18840) );
  AOI21_X1 U21917 ( .B1(n18841), .B2(n18866), .A(n18840), .ZN(n18846) );
  INV_X1 U21918 ( .A(n18842), .ZN(n18843) );
  AOI21_X1 U21919 ( .B1(n18902), .B2(n18843), .A(n18869), .ZN(n18845) );
  OAI22_X1 U21920 ( .A1(n18869), .A2(n18846), .B1(n18845), .B2(n18844), .ZN(
        P3_U3285) );
  INV_X1 U21921 ( .A(n18847), .ZN(n18852) );
  NAND2_X1 U21922 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n18863) );
  AOI22_X1 U21923 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n13107), .B1(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n18848), .ZN(n18857) );
  OAI22_X1 U21924 ( .A1(n18850), .A2(n18849), .B1(n18863), .B2(n18857), .ZN(
        n18851) );
  AOI21_X1 U21925 ( .B1(n18866), .B2(n18852), .A(n18851), .ZN(n18853) );
  AOI22_X1 U21926 ( .A1(n18869), .A2(n18854), .B1(n18853), .B2(n18860), .ZN(
        P3_U3288) );
  INV_X1 U21927 ( .A(n18855), .ZN(n18858) );
  INV_X1 U21928 ( .A(n18863), .ZN(n18856) );
  AOI222_X1 U21929 ( .A1(n18859), .A2(n18902), .B1(n18866), .B2(n18858), .C1(
        n18857), .C2(n18856), .ZN(n18861) );
  AOI22_X1 U21930 ( .A1(n18869), .A2(n18862), .B1(n18861), .B2(n18860), .ZN(
        P3_U3289) );
  OAI221_X1 U21931 ( .B1(P3_STATE2_REG_1__SCAN_IN), .B2(n18865), .C1(
        P3_STATE2_REG_1__SCAN_IN), .C2(n18864), .A(n18863), .ZN(n18868) );
  AOI21_X1 U21932 ( .B1(n18870), .B2(n18866), .A(n18869), .ZN(n18867) );
  AOI22_X1 U21933 ( .A1(n18870), .A2(n18869), .B1(n18868), .B2(n18867), .ZN(
        P3_U3290) );
  AOI21_X1 U21934 ( .B1(P3_REIP_REG_0__SCAN_IN), .B2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n18871) );
  AOI22_X1 U21935 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_0__SCAN_IN), 
        .B1(n18871), .B2(n20815), .ZN(n18874) );
  AOI22_X1 U21936 ( .A1(n20816), .A2(n18874), .B1(n18873), .B2(n18872), .ZN(
        P3_U3292) );
  OAI21_X1 U21937 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(P3_REIP_REG_0__SCAN_IN), 
        .A(n20816), .ZN(n18875) );
  OAI21_X1 U21938 ( .B1(n20816), .B2(n18876), .A(n18875), .ZN(P3_U3293) );
  INV_X1 U21939 ( .A(P3_W_R_N_REG_SCAN_IN), .ZN(n18877) );
  AOI22_X1 U21940 ( .A1(n18898), .A2(P3_READREQUEST_REG_SCAN_IN), .B1(n18877), 
        .B2(n18899), .ZN(P3_U3294) );
  MUX2_X1 U21941 ( .A(P3_MORE_REG_SCAN_IN), .B(n18879), .S(n18878), .Z(
        P3_U3295) );
  AOI21_X1 U21942 ( .B1(n18881), .B2(n18880), .A(n18904), .ZN(n18882) );
  OAI21_X1 U21943 ( .B1(n18884), .B2(n18883), .A(n18882), .ZN(n18897) );
  AOI21_X1 U21944 ( .B1(n18887), .B2(n18886), .A(n18885), .ZN(n18888) );
  INV_X1 U21945 ( .A(n18888), .ZN(n18890) );
  AOI211_X1 U21946 ( .C1(n18903), .C2(n18890), .A(n18889), .B(n18901), .ZN(
        n18892) );
  NOR2_X1 U21947 ( .A1(n18892), .A2(n18891), .ZN(n18893) );
  OAI21_X1 U21948 ( .B1(n18894), .B2(n18893), .A(n18897), .ZN(n18895) );
  OAI21_X1 U21949 ( .B1(n18897), .B2(n18896), .A(n18895), .ZN(P3_U3296) );
  OAI22_X1 U21950 ( .A1(n18899), .A2(P3_MEMORYFETCH_REG_SCAN_IN), .B1(
        P3_M_IO_N_REG_SCAN_IN), .B2(n18898), .ZN(n18900) );
  INV_X1 U21951 ( .A(n18900), .ZN(P3_U3297) );
  AOI21_X1 U21952 ( .B1(n18902), .B2(n18901), .A(n18904), .ZN(n18906) );
  INV_X1 U21953 ( .A(P3_READREQUEST_REG_SCAN_IN), .ZN(n18905) );
  AOI22_X1 U21954 ( .A1(n18906), .A2(n18905), .B1(n18904), .B2(n18903), .ZN(
        P3_U3298) );
  INV_X1 U21955 ( .A(n18906), .ZN(n18908) );
  OAI21_X1 U21956 ( .B1(n18908), .B2(P3_MEMORYFETCH_REG_SCAN_IN), .A(n18907), 
        .ZN(n18909) );
  INV_X1 U21957 ( .A(n18909), .ZN(P3_U3299) );
  INV_X1 U21958 ( .A(P2_ADS_N_REG_SCAN_IN), .ZN(n18911) );
  INV_X1 U21959 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n19830) );
  NAND2_X1 U21960 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n19830), .ZN(n19823) );
  INV_X1 U21961 ( .A(P2_STATE_REG_1__SCAN_IN), .ZN(n18910) );
  NAND2_X1 U21962 ( .A1(n21058), .A2(n18910), .ZN(n19819) );
  OAI21_X1 U21963 ( .B1(n21058), .B2(n19823), .A(n19819), .ZN(n19885) );
  OAI21_X1 U21964 ( .B1(n21058), .B2(n18911), .A(n19811), .ZN(P2_U2815) );
  AOI22_X1 U21965 ( .A1(P2_D_C_N_REG_SCAN_IN), .A2(n19937), .B1(n18913), .B2(
        n21058), .ZN(n18912) );
  OAI21_X1 U21966 ( .B1(P2_CODEFETCH_REG_SCAN_IN), .B2(n19937), .A(n18912), 
        .ZN(P2_U2817) );
  OAI21_X1 U21967 ( .B1(n18913), .B2(BS16), .A(n19885), .ZN(n19883) );
  OAI21_X1 U21968 ( .B1(n19885), .B2(n19573), .A(n19883), .ZN(P2_U2818) );
  NOR2_X1 U21969 ( .A1(n18915), .A2(n18914), .ZN(n19933) );
  INV_X1 U21970 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n18917) );
  OAI21_X1 U21971 ( .B1(n19933), .B2(n18917), .A(n18916), .ZN(P2_U2819) );
  INV_X1 U21972 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n19881) );
  NOR4_X1 U21973 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_10__SCAN_IN), .A3(P2_DATAWIDTH_REG_11__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_12__SCAN_IN), .ZN(n18927) );
  NOR4_X1 U21974 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_5__SCAN_IN), .A3(P2_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_7__SCAN_IN), .ZN(n18926) );
  AOI211_X1 U21975 ( .C1(P2_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_0__SCAN_IN), .A(P2_DATAWIDTH_REG_9__SCAN_IN), .B(
        P2_DATAWIDTH_REG_3__SCAN_IN), .ZN(n18918) );
  INV_X1 U21976 ( .A(P2_DATAWIDTH_REG_17__SCAN_IN), .ZN(n21063) );
  INV_X1 U21977 ( .A(P2_DATAWIDTH_REG_14__SCAN_IN), .ZN(n20947) );
  NAND3_X1 U21978 ( .A1(n18918), .A2(n21063), .A3(n20947), .ZN(n18924) );
  NOR4_X1 U21979 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_20__SCAN_IN), .A3(P2_DATAWIDTH_REG_21__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_22__SCAN_IN), .ZN(n18922) );
  NOR4_X1 U21980 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_15__SCAN_IN), .A3(P2_DATAWIDTH_REG_16__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_18__SCAN_IN), .ZN(n18921) );
  NOR4_X1 U21981 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_29__SCAN_IN), .A3(P2_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_31__SCAN_IN), .ZN(n18920) );
  NOR4_X1 U21982 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_24__SCAN_IN), .A3(P2_DATAWIDTH_REG_25__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_26__SCAN_IN), .ZN(n18919) );
  NAND4_X1 U21983 ( .A1(n18922), .A2(n18921), .A3(n18920), .A4(n18919), .ZN(
        n18923) );
  NOR4_X1 U21984 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_2__SCAN_IN), .A3(n18924), .A4(n18923), .ZN(n18925) );
  NAND3_X1 U21985 ( .A1(n18927), .A2(n18926), .A3(n18925), .ZN(n18934) );
  NOR2_X1 U21986 ( .A1(n18934), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n18928) );
  AOI22_X1 U21987 ( .A1(n19881), .A2(n18934), .B1(n19831), .B2(n18928), .ZN(
        P2_U2820) );
  INV_X1 U21988 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n19879) );
  NOR2_X1 U21989 ( .A1(P2_DATAWIDTH_REG_1__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n18931) );
  NAND2_X1 U21990 ( .A1(n18931), .A2(n18929), .ZN(n18936) );
  NOR2_X1 U21991 ( .A1(n18934), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n18930) );
  AOI22_X1 U21992 ( .A1(n19879), .A2(n18934), .B1(n18936), .B2(n18930), .ZN(
        P2_U2821) );
  INV_X1 U21993 ( .A(n18934), .ZN(n18940) );
  NOR2_X1 U21994 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n18937) );
  INV_X1 U21995 ( .A(n18937), .ZN(n18933) );
  NOR2_X1 U21996 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n18931), .ZN(n18932) );
  MUX2_X1 U21997 ( .A(n18933), .B(n18932), .S(P2_REIP_REG_0__SCAN_IN), .Z(
        n18935) );
  INV_X1 U21998 ( .A(P2_BYTEENABLE_REG_2__SCAN_IN), .ZN(n19877) );
  AOI22_X1 U21999 ( .A1(n18940), .A2(n18935), .B1(n19877), .B2(n18934), .ZN(
        P2_U2822) );
  INV_X1 U22000 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n21195) );
  INV_X1 U22001 ( .A(n18936), .ZN(n18938) );
  OAI21_X1 U22002 ( .B1(n18938), .B2(n18937), .A(n18940), .ZN(n18939) );
  OAI21_X1 U22003 ( .B1(n18940), .B2(n21195), .A(n18939), .ZN(P2_U2823) );
  AOI211_X1 U22004 ( .C1(n18943), .C2(n18942), .A(n18941), .B(n19809), .ZN(
        n18950) );
  OAI22_X1 U22005 ( .A1(n19072), .A2(n10079), .B1(n19856), .B2(n19074), .ZN(
        n18944) );
  AOI21_X1 U22006 ( .B1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n19101), .A(
        n18944), .ZN(n18947) );
  NAND2_X1 U22007 ( .A1(n18945), .A2(n19049), .ZN(n18946) );
  OAI211_X1 U22008 ( .C1(n18948), .C2(n19067), .A(n18947), .B(n18946), .ZN(
        n18949) );
  AOI211_X1 U22009 ( .C1(n19088), .C2(n18951), .A(n18950), .B(n18949), .ZN(
        n18952) );
  INV_X1 U22010 ( .A(n18952), .ZN(P2_U2835) );
  INV_X1 U22011 ( .A(n18953), .ZN(n18963) );
  AOI21_X1 U22012 ( .B1(n19090), .B2(P2_EBX_REG_19__SCAN_IN), .A(n19245), .ZN(
        n18954) );
  OAI21_X1 U22013 ( .B1(n19854), .B2(n19074), .A(n18954), .ZN(n18955) );
  AOI21_X1 U22014 ( .B1(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n19101), .A(
        n18955), .ZN(n18956) );
  OAI21_X1 U22015 ( .B1(n18957), .B2(n19067), .A(n18956), .ZN(n18962) );
  AOI211_X1 U22016 ( .C1(n18960), .C2(n18959), .A(n19809), .B(n18958), .ZN(
        n18961) );
  AOI211_X1 U22017 ( .C1(n19049), .C2(n18963), .A(n18962), .B(n18961), .ZN(
        n18964) );
  OAI21_X1 U22018 ( .B1(n18965), .B2(n19087), .A(n18964), .ZN(P2_U2836) );
  NOR2_X1 U22019 ( .A1(n10053), .A2(n18966), .ZN(n18983) );
  XOR2_X1 U22020 ( .A(n18983), .B(n18967), .Z(n18976) );
  INV_X1 U22021 ( .A(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n18969) );
  OAI222_X1 U22022 ( .A1(n19095), .A2(n18970), .B1(n19057), .B2(n18969), .C1(
        n18968), .C2(n19072), .ZN(n18971) );
  AOI211_X1 U22023 ( .C1(P2_REIP_REG_18__SCAN_IN), .C2(n19091), .A(n19038), 
        .B(n18971), .ZN(n18975) );
  AOI22_X1 U22024 ( .A1(n18973), .A2(n19097), .B1(n19088), .B2(n18972), .ZN(
        n18974) );
  OAI211_X1 U22025 ( .C1(n19809), .C2(n18976), .A(n18975), .B(n18974), .ZN(
        P2_U2837) );
  AOI22_X1 U22026 ( .A1(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n19101), .B1(
        P2_REIP_REG_17__SCAN_IN), .B2(n19091), .ZN(n18989) );
  OAI22_X1 U22027 ( .A1(n18978), .A2(n19095), .B1(n18977), .B2(n18984), .ZN(
        n18979) );
  AOI211_X1 U22028 ( .C1(P2_EBX_REG_17__SCAN_IN), .C2(n19090), .A(n19245), .B(
        n18979), .ZN(n18988) );
  INV_X1 U22029 ( .A(n18980), .ZN(n18981) );
  AOI22_X1 U22030 ( .A1(n18982), .A2(n19097), .B1(n19088), .B2(n18981), .ZN(
        n18987) );
  OAI211_X1 U22031 ( .C1(n18985), .C2(n18984), .A(n9868), .B(n18983), .ZN(
        n18986) );
  NAND4_X1 U22032 ( .A1(n18989), .A2(n18988), .A3(n18987), .A4(n18986), .ZN(
        P2_U2838) );
  AND2_X1 U22033 ( .A1(n19079), .A2(n18990), .ZN(n19008) );
  XNOR2_X1 U22034 ( .A(n18991), .B(n19008), .ZN(n18998) );
  OAI222_X1 U22035 ( .A1(n19095), .A2(n18993), .B1(n19057), .B2(n11332), .C1(
        n18992), .C2(n19072), .ZN(n18994) );
  AOI211_X1 U22036 ( .C1(P2_REIP_REG_16__SCAN_IN), .C2(n19091), .A(n19038), 
        .B(n18994), .ZN(n18997) );
  AOI22_X1 U22037 ( .A1(n18995), .A2(n19097), .B1(n19088), .B2(n19111), .ZN(
        n18996) );
  OAI211_X1 U22038 ( .C1(n19809), .C2(n18998), .A(n18997), .B(n18996), .ZN(
        P2_U2839) );
  INV_X1 U22039 ( .A(n18999), .ZN(n19007) );
  INV_X1 U22040 ( .A(n19009), .ZN(n19003) );
  AOI22_X1 U22041 ( .A1(P2_EBX_REG_15__SCAN_IN), .A2(n19090), .B1(
        P2_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n19101), .ZN(n19000) );
  OAI211_X1 U22042 ( .C1(n19074), .C2(n15437), .A(n19000), .B(n15684), .ZN(
        n19001) );
  AOI21_X1 U22043 ( .B1(n19003), .B2(n19002), .A(n19001), .ZN(n19004) );
  OAI21_X1 U22044 ( .B1(n19005), .B2(n19067), .A(n19004), .ZN(n19006) );
  AOI21_X1 U22045 ( .B1(n19007), .B2(n19049), .A(n19006), .ZN(n19012) );
  OAI211_X1 U22046 ( .C1(n19010), .C2(n19009), .A(n9868), .B(n19008), .ZN(
        n19011) );
  OAI211_X1 U22047 ( .C1(n19087), .C2(n19118), .A(n19012), .B(n19011), .ZN(
        P2_U2840) );
  NOR2_X1 U22048 ( .A1(n10053), .A2(n19013), .ZN(n19016) );
  XOR2_X1 U22049 ( .A(n19016), .B(n19015), .Z(n19023) );
  AOI222_X1 U22050 ( .A1(n19017), .A2(n19049), .B1(
        P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n19101), .C1(
        P2_EBX_REG_14__SCAN_IN), .C2(n19090), .ZN(n19018) );
  INV_X1 U22051 ( .A(n19018), .ZN(n19019) );
  AOI211_X1 U22052 ( .C1(P2_REIP_REG_14__SCAN_IN), .C2(n19091), .A(n19038), 
        .B(n19019), .ZN(n19022) );
  AOI22_X1 U22053 ( .A1(n19020), .A2(n19097), .B1(n19088), .B2(n19119), .ZN(
        n19021) );
  OAI211_X1 U22054 ( .C1(n19809), .C2(n19023), .A(n19022), .B(n19021), .ZN(
        P2_U2841) );
  NAND2_X1 U22055 ( .A1(n19079), .A2(n19024), .ZN(n19026) );
  XOR2_X1 U22056 ( .A(n19026), .B(n19025), .Z(n19033) );
  AOI22_X1 U22057 ( .A1(n19027), .A2(n19049), .B1(
        P2_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n19101), .ZN(n19028) );
  OAI211_X1 U22058 ( .C1(n15449), .C2(n19074), .A(n19028), .B(n15684), .ZN(
        n19031) );
  OAI22_X1 U22059 ( .A1(n19029), .A2(n19067), .B1(n19087), .B2(n19123), .ZN(
        n19030) );
  AOI211_X1 U22060 ( .C1(P2_EBX_REG_13__SCAN_IN), .C2(n19090), .A(n19031), .B(
        n19030), .ZN(n19032) );
  OAI21_X1 U22061 ( .B1(n19033), .B2(n19809), .A(n19032), .ZN(P2_U2842) );
  INV_X1 U22062 ( .A(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n19035) );
  OAI222_X1 U22063 ( .A1(n19095), .A2(n19036), .B1(n19057), .B2(n19035), .C1(
        n19034), .C2(n19072), .ZN(n19037) );
  AOI211_X1 U22064 ( .C1(P2_REIP_REG_10__SCAN_IN), .C2(n19091), .A(n19038), 
        .B(n19037), .ZN(n19045) );
  NOR2_X1 U22065 ( .A1(n10053), .A2(n19039), .ZN(n19041) );
  XNOR2_X1 U22066 ( .A(n19041), .B(n19040), .ZN(n19043) );
  AOI22_X1 U22067 ( .A1(n19043), .A2(n9868), .B1(n19097), .B2(n19042), .ZN(
        n19044) );
  OAI211_X1 U22068 ( .C1(n19132), .C2(n19087), .A(n19045), .B(n19044), .ZN(
        P2_U2845) );
  NAND2_X1 U22069 ( .A1(n19079), .A2(n19046), .ZN(n19048) );
  XOR2_X1 U22070 ( .A(n19048), .B(n19047), .Z(n19056) );
  AOI22_X1 U22071 ( .A1(n19050), .A2(n19049), .B1(n19101), .B2(
        P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n19051) );
  OAI211_X1 U22072 ( .C1(n11530), .C2(n19074), .A(n19051), .B(n15684), .ZN(
        n19054) );
  OAI22_X1 U22073 ( .A1(n19138), .A2(n19087), .B1(n19067), .B2(n19052), .ZN(
        n19053) );
  AOI211_X1 U22074 ( .C1(P2_EBX_REG_7__SCAN_IN), .C2(n19090), .A(n19054), .B(
        n19053), .ZN(n19055) );
  OAI21_X1 U22075 ( .B1(n19056), .B2(n19809), .A(n19055), .ZN(P2_U2848) );
  INV_X1 U22076 ( .A(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n19058) );
  OAI22_X1 U22077 ( .A1(n19059), .A2(n19095), .B1(n19058), .B2(n19057), .ZN(
        n19060) );
  INV_X1 U22078 ( .A(n19060), .ZN(n19061) );
  OAI211_X1 U22079 ( .C1(n19838), .C2(n19074), .A(n12458), .B(n19061), .ZN(
        n19062) );
  INV_X1 U22080 ( .A(n19062), .ZN(n19071) );
  NOR2_X1 U22081 ( .A1(n10053), .A2(n19063), .ZN(n19064) );
  XNOR2_X1 U22082 ( .A(n19065), .B(n19064), .ZN(n19069) );
  OAI22_X1 U22083 ( .A1(n19139), .A2(n19087), .B1(n19067), .B2(n19066), .ZN(
        n19068) );
  AOI21_X1 U22084 ( .B1(n19069), .B2(n9868), .A(n19068), .ZN(n19070) );
  OAI211_X1 U22085 ( .C1(n11524), .C2(n19072), .A(n19071), .B(n19070), .ZN(
        P2_U2849) );
  OAI21_X1 U22086 ( .B1(n19073), .B2(n19072), .A(n12458), .ZN(n19077) );
  OAI22_X1 U22087 ( .A1(n19075), .A2(n19095), .B1(n19836), .B2(n19074), .ZN(
        n19076) );
  AOI211_X1 U22088 ( .C1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .C2(n19101), .A(
        n19077), .B(n19076), .ZN(n19086) );
  NAND2_X1 U22089 ( .A1(n19079), .A2(n19078), .ZN(n19080) );
  XNOR2_X1 U22090 ( .A(n19081), .B(n19080), .ZN(n19084) );
  AOI22_X1 U22091 ( .A1(n19084), .A2(n9868), .B1(n19097), .B2(n19082), .ZN(
        n19085) );
  OAI211_X1 U22092 ( .C1(n19087), .C2(n19146), .A(n19086), .B(n19085), .ZN(
        P2_U2850) );
  NAND2_X1 U22093 ( .A1(n19089), .A2(n19088), .ZN(n19093) );
  AOI22_X1 U22094 ( .A1(n19091), .A2(P2_REIP_REG_0__SCAN_IN), .B1(n19090), 
        .B2(P2_EBX_REG_0__SCAN_IN), .ZN(n19092) );
  OAI211_X1 U22095 ( .C1(n19095), .C2(n19094), .A(n19093), .B(n19092), .ZN(
        n19096) );
  AOI21_X1 U22096 ( .B1(n19098), .B2(n19097), .A(n19096), .ZN(n19104) );
  AOI22_X1 U22097 ( .A1(n19921), .A2(n19100), .B1(n19099), .B2(n9868), .ZN(
        n19103) );
  NAND2_X1 U22098 ( .A1(P2_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n19101), .ZN(
        n19102) );
  NAND3_X1 U22099 ( .A1(n19104), .A2(n19103), .A3(n19102), .ZN(P2_U2855) );
  AOI22_X1 U22100 ( .A1(n12453), .A2(n19156), .B1(n19109), .B2(
        BUF2_REG_31__SCAN_IN), .ZN(n19106) );
  AOI22_X1 U22101 ( .A1(P2_EAX_REG_31__SCAN_IN), .A2(n19155), .B1(n19110), 
        .B2(BUF1_REG_31__SCAN_IN), .ZN(n19105) );
  NAND2_X1 U22102 ( .A1(n19106), .A2(n19105), .ZN(P2_U2888) );
  AOI22_X1 U22103 ( .A1(n19108), .A2(n19107), .B1(n19155), .B2(
        P2_EAX_REG_16__SCAN_IN), .ZN(n19115) );
  AOI22_X1 U22104 ( .A1(n19110), .A2(BUF1_REG_16__SCAN_IN), .B1(n19109), .B2(
        BUF2_REG_16__SCAN_IN), .ZN(n19114) );
  AOI22_X1 U22105 ( .A1(n19112), .A2(n19116), .B1(n19156), .B2(n19111), .ZN(
        n19113) );
  NAND3_X1 U22106 ( .A1(n19115), .A2(n19114), .A3(n19113), .ZN(P2_U2903) );
  INV_X1 U22107 ( .A(n19129), .ZN(n19164) );
  OAI222_X1 U22108 ( .A1(n19118), .A2(n19147), .B1(n13474), .B2(n19140), .C1(
        n19117), .C2(n19164), .ZN(P2_U2904) );
  INV_X1 U22109 ( .A(n19119), .ZN(n19121) );
  AOI22_X1 U22110 ( .A1(P2_EAX_REG_14__SCAN_IN), .A2(n19155), .B1(n19238), 
        .B2(n19129), .ZN(n19120) );
  OAI21_X1 U22111 ( .B1(n19147), .B2(n19121), .A(n19120), .ZN(P2_U2905) );
  INV_X1 U22112 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n19208) );
  OAI222_X1 U22113 ( .A1(n19123), .A2(n19147), .B1(n19208), .B2(n19140), .C1(
        n19164), .C2(n19122), .ZN(P2_U2906) );
  AOI22_X1 U22114 ( .A1(P2_EAX_REG_12__SCAN_IN), .A2(n19155), .B1(n19124), 
        .B2(n19129), .ZN(n19125) );
  OAI21_X1 U22115 ( .B1(n19147), .B2(n19126), .A(n19125), .ZN(P2_U2907) );
  INV_X1 U22116 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n19212) );
  OAI222_X1 U22117 ( .A1(n19128), .A2(n19147), .B1(n19212), .B2(n19140), .C1(
        n19164), .C2(n19127), .ZN(P2_U2908) );
  AOI22_X1 U22118 ( .A1(P2_EAX_REG_10__SCAN_IN), .A2(n19155), .B1(n19130), 
        .B2(n19129), .ZN(n19131) );
  OAI21_X1 U22119 ( .B1(n19147), .B2(n19132), .A(n19131), .ZN(P2_U2909) );
  INV_X1 U22120 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n19216) );
  OAI222_X1 U22121 ( .A1(n19134), .A2(n19147), .B1(n19216), .B2(n19140), .C1(
        n19164), .C2(n19133), .ZN(P2_U2910) );
  INV_X1 U22122 ( .A(n19135), .ZN(n19137) );
  INV_X1 U22123 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n19218) );
  OAI222_X1 U22124 ( .A1(n19137), .A2(n19147), .B1(n19218), .B2(n19140), .C1(
        n19164), .C2(n19136), .ZN(P2_U2911) );
  INV_X1 U22125 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n19220) );
  OAI222_X1 U22126 ( .A1(n19138), .A2(n19147), .B1(n19220), .B2(n19140), .C1(
        n19164), .C2(n19299), .ZN(P2_U2912) );
  INV_X1 U22127 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n19222) );
  OAI222_X1 U22128 ( .A1(n19139), .A2(n19147), .B1(n19222), .B2(n19140), .C1(
        n19164), .C2(n19291), .ZN(P2_U2913) );
  INV_X1 U22129 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n19224) );
  OAI22_X1 U22130 ( .A1(n19224), .A2(n19140), .B1(n19287), .B2(n19164), .ZN(
        n19141) );
  INV_X1 U22131 ( .A(n19141), .ZN(n19145) );
  OR3_X1 U22132 ( .A1(n19143), .A2(n19142), .A3(n19160), .ZN(n19144) );
  OAI211_X1 U22133 ( .C1(n19147), .C2(n19146), .A(n19145), .B(n19144), .ZN(
        P2_U2914) );
  AOI22_X1 U22134 ( .A1(n19892), .A2(n19156), .B1(P2_EAX_REG_3__SCAN_IN), .B2(
        n19155), .ZN(n19153) );
  AOI21_X1 U22135 ( .B1(n19150), .B2(n19149), .A(n19148), .ZN(n19151) );
  OR2_X1 U22136 ( .A1(n19151), .A2(n19160), .ZN(n19152) );
  OAI211_X1 U22137 ( .C1(n19154), .C2(n19164), .A(n19153), .B(n19152), .ZN(
        P2_U2916) );
  AOI22_X1 U22138 ( .A1(n19156), .A2(n19906), .B1(P2_EAX_REG_1__SCAN_IN), .B2(
        n19155), .ZN(n19163) );
  AOI21_X1 U22139 ( .B1(n19159), .B2(n19158), .A(n19157), .ZN(n19161) );
  OR2_X1 U22140 ( .A1(n19161), .A2(n19160), .ZN(n19162) );
  OAI211_X1 U22141 ( .C1(n19272), .C2(n19164), .A(n19163), .B(n19162), .ZN(
        P2_U2918) );
  NAND2_X1 U22142 ( .A1(n19165), .A2(n19808), .ZN(n19167) );
  NAND2_X1 U22143 ( .A1(n19167), .A2(n19166), .ZN(n19168) );
  NAND2_X1 U22144 ( .A1(n19236), .A2(n19169), .ZN(n19174) );
  INV_X2 U22145 ( .A(n19174), .ZN(n19233) );
  AND2_X1 U22146 ( .A1(n19233), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(P2_U2920)
         );
  INV_X1 U22147 ( .A(n19202), .ZN(n19171) );
  AOI22_X1 U22148 ( .A1(P2_EAX_REG_30__SCAN_IN), .A2(n19171), .B1(n19234), 
        .B2(P2_UWORD_REG_14__SCAN_IN), .ZN(n19172) );
  OAI21_X1 U22149 ( .B1(n19174), .B2(n19173), .A(n19172), .ZN(P2_U2921) );
  AOI22_X1 U22150 ( .A1(n19234), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(n19233), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n19175) );
  OAI21_X1 U22151 ( .B1(n19176), .B2(n19202), .A(n19175), .ZN(P2_U2922) );
  AOI22_X1 U22152 ( .A1(n19234), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(n19233), 
        .B2(P2_DATAO_REG_28__SCAN_IN), .ZN(n19177) );
  OAI21_X1 U22153 ( .B1(n19178), .B2(n19202), .A(n19177), .ZN(P2_U2923) );
  AOI22_X1 U22154 ( .A1(n19196), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(n19233), 
        .B2(P2_DATAO_REG_27__SCAN_IN), .ZN(n19179) );
  OAI21_X1 U22155 ( .B1(n19180), .B2(n19202), .A(n19179), .ZN(P2_U2924) );
  AOI22_X1 U22156 ( .A1(n19196), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(n19233), 
        .B2(P2_DATAO_REG_26__SCAN_IN), .ZN(n19181) );
  OAI21_X1 U22157 ( .B1(n19182), .B2(n19202), .A(n19181), .ZN(P2_U2925) );
  AOI22_X1 U22158 ( .A1(n19196), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(n19233), 
        .B2(P2_DATAO_REG_25__SCAN_IN), .ZN(n19183) );
  OAI21_X1 U22159 ( .B1(n19184), .B2(n19202), .A(n19183), .ZN(P2_U2926) );
  AOI22_X1 U22160 ( .A1(n19196), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(n19233), 
        .B2(P2_DATAO_REG_24__SCAN_IN), .ZN(n19185) );
  OAI21_X1 U22161 ( .B1(n19186), .B2(n19202), .A(n19185), .ZN(P2_U2927) );
  INV_X1 U22162 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n19188) );
  AOI22_X1 U22163 ( .A1(n19196), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n19233), 
        .B2(P2_DATAO_REG_23__SCAN_IN), .ZN(n19187) );
  OAI21_X1 U22164 ( .B1(n19188), .B2(n19202), .A(n19187), .ZN(P2_U2928) );
  INV_X1 U22165 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n19190) );
  AOI22_X1 U22166 ( .A1(n19196), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(n19233), 
        .B2(P2_DATAO_REG_22__SCAN_IN), .ZN(n19189) );
  OAI21_X1 U22167 ( .B1(n19190), .B2(n19202), .A(n19189), .ZN(P2_U2929) );
  INV_X1 U22168 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n19192) );
  AOI22_X1 U22169 ( .A1(n19196), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n19233), 
        .B2(P2_DATAO_REG_21__SCAN_IN), .ZN(n19191) );
  OAI21_X1 U22170 ( .B1(n19192), .B2(n19202), .A(n19191), .ZN(P2_U2930) );
  INV_X1 U22171 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n19194) );
  AOI22_X1 U22172 ( .A1(n19196), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n19233), 
        .B2(P2_DATAO_REG_20__SCAN_IN), .ZN(n19193) );
  OAI21_X1 U22173 ( .B1(n19194), .B2(n19202), .A(n19193), .ZN(P2_U2931) );
  INV_X1 U22174 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n21012) );
  AOI22_X1 U22175 ( .A1(n19196), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n19233), 
        .B2(P2_DATAO_REG_19__SCAN_IN), .ZN(n19195) );
  OAI21_X1 U22176 ( .B1(n21012), .B2(n19202), .A(n19195), .ZN(P2_U2932) );
  INV_X1 U22177 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n19198) );
  AOI22_X1 U22178 ( .A1(n19196), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n19233), 
        .B2(P2_DATAO_REG_18__SCAN_IN), .ZN(n19197) );
  OAI21_X1 U22179 ( .B1(n19198), .B2(n19202), .A(n19197), .ZN(P2_U2933) );
  INV_X1 U22180 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n19200) );
  AOI22_X1 U22181 ( .A1(n19234), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n19233), 
        .B2(P2_DATAO_REG_17__SCAN_IN), .ZN(n19199) );
  OAI21_X1 U22182 ( .B1(n19200), .B2(n19202), .A(n19199), .ZN(P2_U2934) );
  INV_X1 U22183 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n19203) );
  AOI22_X1 U22184 ( .A1(n19234), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(n19233), 
        .B2(P2_DATAO_REG_16__SCAN_IN), .ZN(n19201) );
  OAI21_X1 U22185 ( .B1(n19203), .B2(n19202), .A(n19201), .ZN(P2_U2935) );
  AOI22_X1 U22186 ( .A1(n19234), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n19233), 
        .B2(P2_DATAO_REG_15__SCAN_IN), .ZN(n19204) );
  OAI21_X1 U22187 ( .B1(n13474), .B2(n19236), .A(n19204), .ZN(P2_U2936) );
  INV_X1 U22188 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n19206) );
  AOI22_X1 U22189 ( .A1(n19234), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n19233), 
        .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n19205) );
  OAI21_X1 U22190 ( .B1(n19206), .B2(n19236), .A(n19205), .ZN(P2_U2937) );
  AOI22_X1 U22191 ( .A1(n19234), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n19233), 
        .B2(P2_DATAO_REG_13__SCAN_IN), .ZN(n19207) );
  OAI21_X1 U22192 ( .B1(n19208), .B2(n19236), .A(n19207), .ZN(P2_U2938) );
  AOI22_X1 U22193 ( .A1(n19234), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(n19233), 
        .B2(P2_DATAO_REG_12__SCAN_IN), .ZN(n19209) );
  OAI21_X1 U22194 ( .B1(n19210), .B2(n19236), .A(n19209), .ZN(P2_U2939) );
  AOI22_X1 U22195 ( .A1(n19234), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n19233), 
        .B2(P2_DATAO_REG_11__SCAN_IN), .ZN(n19211) );
  OAI21_X1 U22196 ( .B1(n19212), .B2(n19236), .A(n19211), .ZN(P2_U2940) );
  AOI22_X1 U22197 ( .A1(n19234), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(n19233), 
        .B2(P2_DATAO_REG_10__SCAN_IN), .ZN(n19213) );
  OAI21_X1 U22198 ( .B1(n19214), .B2(n19236), .A(n19213), .ZN(P2_U2941) );
  AOI22_X1 U22199 ( .A1(n19234), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n19233), 
        .B2(P2_DATAO_REG_9__SCAN_IN), .ZN(n19215) );
  OAI21_X1 U22200 ( .B1(n19216), .B2(n19236), .A(n19215), .ZN(P2_U2942) );
  AOI22_X1 U22201 ( .A1(n19234), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n19233), 
        .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n19217) );
  OAI21_X1 U22202 ( .B1(n19218), .B2(n19236), .A(n19217), .ZN(P2_U2943) );
  AOI22_X1 U22203 ( .A1(n19234), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n19233), 
        .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n19219) );
  OAI21_X1 U22204 ( .B1(n19220), .B2(n19236), .A(n19219), .ZN(P2_U2944) );
  AOI22_X1 U22205 ( .A1(n19234), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n19233), 
        .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n19221) );
  OAI21_X1 U22206 ( .B1(n19222), .B2(n19236), .A(n19221), .ZN(P2_U2945) );
  AOI22_X1 U22207 ( .A1(n19234), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n19233), 
        .B2(P2_DATAO_REG_5__SCAN_IN), .ZN(n19223) );
  OAI21_X1 U22208 ( .B1(n19224), .B2(n19236), .A(n19223), .ZN(P2_U2946) );
  INV_X1 U22209 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n19226) );
  AOI22_X1 U22210 ( .A1(n19234), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n19233), 
        .B2(P2_DATAO_REG_4__SCAN_IN), .ZN(n19225) );
  OAI21_X1 U22211 ( .B1(n19226), .B2(n19236), .A(n19225), .ZN(P2_U2947) );
  INV_X1 U22212 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n19228) );
  AOI22_X1 U22213 ( .A1(n19234), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n19233), 
        .B2(P2_DATAO_REG_3__SCAN_IN), .ZN(n19227) );
  OAI21_X1 U22214 ( .B1(n19228), .B2(n19236), .A(n19227), .ZN(P2_U2948) );
  INV_X1 U22215 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n19230) );
  AOI22_X1 U22216 ( .A1(n19234), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n19233), 
        .B2(P2_DATAO_REG_2__SCAN_IN), .ZN(n19229) );
  OAI21_X1 U22217 ( .B1(n19230), .B2(n19236), .A(n19229), .ZN(P2_U2949) );
  INV_X1 U22218 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n19232) );
  AOI22_X1 U22219 ( .A1(n19234), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n19233), 
        .B2(P2_DATAO_REG_1__SCAN_IN), .ZN(n19231) );
  OAI21_X1 U22220 ( .B1(n19232), .B2(n19236), .A(n19231), .ZN(P2_U2950) );
  AOI22_X1 U22221 ( .A1(n19234), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n19233), 
        .B2(P2_DATAO_REG_0__SCAN_IN), .ZN(n19235) );
  OAI21_X1 U22222 ( .B1(n13576), .B2(n19236), .A(n19235), .ZN(P2_U2951) );
  AOI22_X1 U22223 ( .A1(n19237), .A2(P2_UWORD_REG_14__SCAN_IN), .B1(
        P2_EAX_REG_30__SCAN_IN), .B2(n19241), .ZN(n19240) );
  NAND2_X1 U22224 ( .A1(n19239), .A2(n19238), .ZN(n19243) );
  NAND2_X1 U22225 ( .A1(n19240), .A2(n19243), .ZN(P2_U2966) );
  AOI22_X1 U22226 ( .A1(n19242), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n19241), 
        .B2(P2_EAX_REG_14__SCAN_IN), .ZN(n19244) );
  NAND2_X1 U22227 ( .A1(n19244), .A2(n19243), .ZN(P2_U2981) );
  AOI22_X1 U22228 ( .A1(n19246), .A2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B1(
        P2_REIP_REG_4__SCAN_IN), .B2(n19245), .ZN(n19254) );
  AOI222_X1 U22229 ( .A1(n19252), .A2(n19251), .B1(n19250), .B2(n19249), .C1(
        n19248), .C2(n19247), .ZN(n19253) );
  OAI211_X1 U22230 ( .C1(n19256), .C2(n19255), .A(n19254), .B(n19253), .ZN(
        P2_U3010) );
  NAND2_X1 U22231 ( .A1(n19354), .A2(n19914), .ZN(n19310) );
  NOR2_X1 U22232 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19310), .ZN(
        n19298) );
  AOI22_X1 U22233 ( .A1(n19780), .A2(n19749), .B1(n19740), .B2(n19298), .ZN(
        n19269) );
  INV_X1 U22234 ( .A(n19332), .ZN(n19258) );
  NOR2_X1 U22235 ( .A1(n19780), .A2(n19258), .ZN(n19259) );
  OAI21_X1 U22236 ( .B1(n19259), .B2(n19573), .A(n19691), .ZN(n19267) );
  NOR2_X1 U22237 ( .A1(n19898), .A2(n19260), .ZN(n19791) );
  NOR2_X1 U22238 ( .A1(n19791), .A2(n19298), .ZN(n19266) );
  INV_X1 U22239 ( .A(n19266), .ZN(n19263) );
  INV_X1 U22240 ( .A(n19298), .ZN(n19261) );
  OAI211_X1 U22241 ( .C1(n12072), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19886), 
        .B(n19261), .ZN(n19262) );
  OAI211_X1 U22242 ( .C1(n19267), .C2(n19263), .A(n19747), .B(n19262), .ZN(
        n19301) );
  INV_X1 U22243 ( .A(n12072), .ZN(n19264) );
  OAI21_X1 U22244 ( .B1(n19264), .B2(n19298), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19265) );
  AOI22_X1 U22245 ( .A1(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n19301), .B1(
        n19741), .B2(n19300), .ZN(n19268) );
  OAI211_X1 U22246 ( .C1(n19752), .C2(n19332), .A(n19269), .B(n19268), .ZN(
        P2_U3048) );
  AOI22_X1 U22247 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n19295), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n19294), .ZN(n19758) );
  AOI22_X1 U22248 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n19294), .B1(
        BUF1_REG_25__SCAN_IN), .B2(n19295), .ZN(n19707) );
  NOR2_X2 U22249 ( .A1(n19271), .A2(n19270), .ZN(n19753) );
  AOI22_X1 U22250 ( .A1(n19780), .A2(n19755), .B1(n19753), .B2(n19298), .ZN(
        n19274) );
  NOR2_X2 U22251 ( .A1(n19272), .A2(n19389), .ZN(n19754) );
  AOI22_X1 U22252 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n19301), .B1(
        n19754), .B2(n19300), .ZN(n19273) );
  OAI211_X1 U22253 ( .C1(n19758), .C2(n19332), .A(n19274), .B(n19273), .ZN(
        P2_U3049) );
  AOI22_X1 U22254 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n19295), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n19294), .ZN(n19764) );
  AOI22_X1 U22255 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n19295), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n19294), .ZN(n19711) );
  AOI22_X1 U22256 ( .A1(n19780), .A2(n19761), .B1(n19759), .B2(n19298), .ZN(
        n19278) );
  NOR2_X2 U22257 ( .A1(n19276), .A2(n19389), .ZN(n19760) );
  AOI22_X1 U22258 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n19301), .B1(
        n19760), .B2(n19300), .ZN(n19277) );
  OAI211_X1 U22259 ( .C1(n19764), .C2(n19332), .A(n19278), .B(n19277), .ZN(
        P2_U3050) );
  AOI22_X1 U22260 ( .A1(n19780), .A2(n19767), .B1(n19765), .B2(n19298), .ZN(
        n19280) );
  AOI22_X1 U22261 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n19301), .B1(
        n19766), .B2(n19300), .ZN(n19279) );
  OAI211_X1 U22262 ( .C1(n19770), .C2(n19332), .A(n19280), .B(n19279), .ZN(
        P2_U3051) );
  AOI22_X1 U22263 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n19295), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n19294), .ZN(n19717) );
  AOI22_X1 U22264 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n19295), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n19294), .ZN(n19776) );
  INV_X1 U22265 ( .A(n19776), .ZN(n19714) );
  AOI22_X1 U22266 ( .A1(n19714), .A2(n19780), .B1(n19771), .B2(n19298), .ZN(
        n19285) );
  INV_X1 U22267 ( .A(n19282), .ZN(n19283) );
  NOR2_X2 U22268 ( .A1(n19283), .A2(n19389), .ZN(n19772) );
  AOI22_X1 U22269 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n19301), .B1(
        n19772), .B2(n19300), .ZN(n19284) );
  OAI211_X1 U22270 ( .C1(n19717), .C2(n19332), .A(n19285), .B(n19284), .ZN(
        P2_U3052) );
  AOI22_X1 U22271 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n19294), .B1(
        BUF1_REG_29__SCAN_IN), .B2(n19295), .ZN(n19784) );
  AOI22_X1 U22272 ( .A1(n19780), .A2(n19719), .B1(n19777), .B2(n19298), .ZN(
        n19289) );
  NOR2_X2 U22273 ( .A1(n19287), .A2(n19389), .ZN(n19778) );
  AOI22_X1 U22274 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n19301), .B1(
        n19778), .B2(n19300), .ZN(n19288) );
  OAI211_X1 U22275 ( .C1(n19722), .C2(n19332), .A(n19289), .B(n19288), .ZN(
        P2_U3053) );
  AOI22_X1 U22276 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n19295), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n19294), .ZN(n19726) );
  AND2_X1 U22277 ( .A1(n19290), .A2(n19296), .ZN(n19785) );
  AOI22_X1 U22278 ( .A1(n19780), .A2(n19787), .B1(n19785), .B2(n19298), .ZN(
        n19293) );
  NOR2_X2 U22279 ( .A1(n19291), .A2(n19389), .ZN(n19786) );
  AOI22_X1 U22280 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n19301), .B1(
        n19786), .B2(n19300), .ZN(n19292) );
  OAI211_X1 U22281 ( .C1(n19790), .C2(n19332), .A(n19293), .B(n19292), .ZN(
        P2_U3054) );
  AOI22_X1 U22282 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n19295), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n19294), .ZN(n19801) );
  AOI22_X1 U22283 ( .A1(BUF1_REG_31__SCAN_IN), .A2(n19295), .B1(
        BUF2_REG_31__SCAN_IN), .B2(n19294), .ZN(n19734) );
  AND2_X1 U22284 ( .A1(n19297), .A2(n19296), .ZN(n19792) );
  AOI22_X1 U22285 ( .A1(n19780), .A2(n19795), .B1(n19792), .B2(n19298), .ZN(
        n19303) );
  NOR2_X2 U22286 ( .A1(n19299), .A2(n19389), .ZN(n19793) );
  AOI22_X1 U22287 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n19301), .B1(
        n19793), .B2(n19300), .ZN(n19302) );
  OAI211_X1 U22288 ( .C1(n19801), .C2(n19332), .A(n19303), .B(n19302), .ZN(
        P2_U3055) );
  INV_X1 U22289 ( .A(n19304), .ZN(n19306) );
  NOR2_X1 U22290 ( .A1(n19538), .A2(n19305), .ZN(n19327) );
  NOR3_X1 U22291 ( .A1(n19306), .A2(n19327), .A3(n19735), .ZN(n19309) );
  INV_X1 U22292 ( .A(n19310), .ZN(n19307) );
  AOI21_X1 U22293 ( .B1(n19917), .B2(n19307), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19308) );
  NOR2_X1 U22294 ( .A1(n19309), .A2(n19308), .ZN(n19328) );
  AOI22_X1 U22295 ( .A1(n19328), .A2(n19741), .B1(n19740), .B2(n19327), .ZN(
        n19314) );
  AND2_X1 U22296 ( .A1(n19539), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19480) );
  INV_X1 U22297 ( .A(n19540), .ZN(n19536) );
  NAND2_X1 U22298 ( .A1(n19480), .A2(n19536), .ZN(n19311) );
  AOI21_X1 U22299 ( .B1(n19311), .B2(n19310), .A(n19309), .ZN(n19312) );
  OAI211_X1 U22300 ( .C1(n19327), .C2(n19917), .A(n19312), .B(n19747), .ZN(
        n19329) );
  AOI22_X1 U22301 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19329), .B1(
        n19349), .B2(n19690), .ZN(n19313) );
  OAI211_X1 U22302 ( .C1(n19703), .C2(n19332), .A(n19314), .B(n19313), .ZN(
        P2_U3056) );
  AOI22_X1 U22303 ( .A1(n19328), .A2(n19754), .B1(n19753), .B2(n19327), .ZN(
        n19316) );
  AOI22_X1 U22304 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19329), .B1(
        n19349), .B2(n19704), .ZN(n19315) );
  OAI211_X1 U22305 ( .C1(n19707), .C2(n19332), .A(n19316), .B(n19315), .ZN(
        P2_U3057) );
  AOI22_X1 U22306 ( .A1(n19328), .A2(n19760), .B1(n19759), .B2(n19327), .ZN(
        n19318) );
  INV_X1 U22307 ( .A(n19764), .ZN(n19708) );
  AOI22_X1 U22308 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19329), .B1(
        n19349), .B2(n19708), .ZN(n19317) );
  OAI211_X1 U22309 ( .C1(n19711), .C2(n19332), .A(n19318), .B(n19317), .ZN(
        P2_U3058) );
  AOI22_X1 U22310 ( .A1(n19328), .A2(n19766), .B1(n19765), .B2(n19327), .ZN(
        n19320) );
  AOI22_X1 U22311 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19329), .B1(
        n19349), .B2(n19620), .ZN(n19319) );
  OAI211_X1 U22312 ( .C1(n19623), .C2(n19332), .A(n19320), .B(n19319), .ZN(
        P2_U3059) );
  AOI22_X1 U22313 ( .A1(n19328), .A2(n19772), .B1(n19771), .B2(n19327), .ZN(
        n19322) );
  AOI22_X1 U22314 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19329), .B1(
        n19349), .B2(n19773), .ZN(n19321) );
  OAI211_X1 U22315 ( .C1(n19776), .C2(n19332), .A(n19322), .B(n19321), .ZN(
        P2_U3060) );
  AOI22_X1 U22316 ( .A1(n19328), .A2(n19778), .B1(n19777), .B2(n19327), .ZN(
        n19324) );
  INV_X1 U22317 ( .A(n19722), .ZN(n19779) );
  AOI22_X1 U22318 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19329), .B1(
        n19349), .B2(n19779), .ZN(n19323) );
  OAI211_X1 U22319 ( .C1(n19784), .C2(n19332), .A(n19324), .B(n19323), .ZN(
        P2_U3061) );
  AOI22_X1 U22320 ( .A1(n19328), .A2(n19786), .B1(n19785), .B2(n19327), .ZN(
        n19326) );
  INV_X1 U22321 ( .A(n19790), .ZN(n19723) );
  AOI22_X1 U22322 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19329), .B1(
        n19349), .B2(n19723), .ZN(n19325) );
  OAI211_X1 U22323 ( .C1(n19726), .C2(n19332), .A(n19326), .B(n19325), .ZN(
        P2_U3062) );
  AOI22_X1 U22324 ( .A1(n19328), .A2(n19793), .B1(n19792), .B2(n19327), .ZN(
        n19331) );
  INV_X1 U22325 ( .A(n19801), .ZN(n19728) );
  AOI22_X1 U22326 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19329), .B1(
        n19349), .B2(n19728), .ZN(n19330) );
  OAI211_X1 U22327 ( .C1(n19734), .C2(n19332), .A(n19331), .B(n19330), .ZN(
        P2_U3063) );
  AOI22_X1 U22328 ( .A1(n19348), .A2(n19754), .B1(n19753), .B2(n19347), .ZN(
        n19334) );
  AOI22_X1 U22329 ( .A1(n19379), .A2(n19704), .B1(n19349), .B2(n19755), .ZN(
        n19333) );
  OAI211_X1 U22330 ( .C1(n19338), .C2(n19335), .A(n19334), .B(n19333), .ZN(
        P2_U3065) );
  AOI22_X1 U22331 ( .A1(n19348), .A2(n19760), .B1(n19759), .B2(n19347), .ZN(
        n19337) );
  AOI22_X1 U22332 ( .A1(n19349), .A2(n19761), .B1(n19379), .B2(n19708), .ZN(
        n19336) );
  OAI211_X1 U22333 ( .C1(n19338), .C2(n21044), .A(n19337), .B(n19336), .ZN(
        P2_U3066) );
  AOI22_X1 U22334 ( .A1(n19348), .A2(n19766), .B1(n19765), .B2(n19347), .ZN(
        n19340) );
  AOI22_X1 U22335 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19350), .B1(
        n19349), .B2(n19767), .ZN(n19339) );
  OAI211_X1 U22336 ( .C1(n19770), .C2(n19373), .A(n19340), .B(n19339), .ZN(
        P2_U3067) );
  AOI22_X1 U22337 ( .A1(n19348), .A2(n19772), .B1(n19771), .B2(n19347), .ZN(
        n19342) );
  AOI22_X1 U22338 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19350), .B1(
        n19349), .B2(n19714), .ZN(n19341) );
  OAI211_X1 U22339 ( .C1(n19717), .C2(n19373), .A(n19342), .B(n19341), .ZN(
        P2_U3068) );
  AOI22_X1 U22340 ( .A1(n19348), .A2(n19778), .B1(n19777), .B2(n19347), .ZN(
        n19344) );
  AOI22_X1 U22341 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19350), .B1(
        n19349), .B2(n19719), .ZN(n19343) );
  OAI211_X1 U22342 ( .C1(n19722), .C2(n19373), .A(n19344), .B(n19343), .ZN(
        P2_U3069) );
  AOI22_X1 U22343 ( .A1(n19348), .A2(n19786), .B1(n19785), .B2(n19347), .ZN(
        n19346) );
  AOI22_X1 U22344 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19350), .B1(
        n19349), .B2(n19787), .ZN(n19345) );
  OAI211_X1 U22345 ( .C1(n19790), .C2(n19373), .A(n19346), .B(n19345), .ZN(
        P2_U3070) );
  AOI22_X1 U22346 ( .A1(n19348), .A2(n19793), .B1(n19792), .B2(n19347), .ZN(
        n19352) );
  AOI22_X1 U22347 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19350), .B1(
        n19349), .B2(n19795), .ZN(n19351) );
  OAI211_X1 U22348 ( .C1(n19801), .C2(n19373), .A(n19352), .B(n19351), .ZN(
        P2_U3071) );
  AND2_X1 U22349 ( .A1(n19606), .A2(n19354), .ZN(n19378) );
  AOI22_X1 U22350 ( .A1(n19749), .A2(n19379), .B1(n19740), .B2(n19378), .ZN(
        n19364) );
  INV_X1 U22351 ( .A(n19480), .ZN(n19353) );
  OAI21_X1 U22352 ( .B1(n19353), .B2(n19889), .A(n19691), .ZN(n19362) );
  NAND2_X1 U22353 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19354), .ZN(
        n19361) );
  INV_X1 U22354 ( .A(n19361), .ZN(n19357) );
  INV_X1 U22355 ( .A(n19378), .ZN(n19355) );
  OAI211_X1 U22356 ( .C1(n19358), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19886), 
        .B(n19355), .ZN(n19356) );
  OAI211_X1 U22357 ( .C1(n19362), .C2(n19357), .A(n19747), .B(n19356), .ZN(
        n19381) );
  INV_X1 U22358 ( .A(n19358), .ZN(n19359) );
  OAI21_X1 U22359 ( .B1(n19359), .B2(n19378), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19360) );
  OAI21_X1 U22360 ( .B1(n19362), .B2(n19361), .A(n19360), .ZN(n19380) );
  AOI22_X1 U22361 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19381), .B1(
        n19741), .B2(n19380), .ZN(n19363) );
  OAI211_X1 U22362 ( .C1(n19752), .C2(n19387), .A(n19364), .B(n19363), .ZN(
        P2_U3072) );
  AOI22_X1 U22363 ( .A1(n19755), .A2(n19379), .B1(n19378), .B2(n19753), .ZN(
        n19366) );
  AOI22_X1 U22364 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19381), .B1(
        n19754), .B2(n19380), .ZN(n19365) );
  OAI211_X1 U22365 ( .C1(n19758), .C2(n19387), .A(n19366), .B(n19365), .ZN(
        P2_U3073) );
  AOI22_X1 U22366 ( .A1(n19708), .A2(n19410), .B1(n19378), .B2(n19759), .ZN(
        n19368) );
  AOI22_X1 U22367 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19381), .B1(
        n19760), .B2(n19380), .ZN(n19367) );
  OAI211_X1 U22368 ( .C1(n19711), .C2(n19373), .A(n19368), .B(n19367), .ZN(
        P2_U3074) );
  AOI22_X1 U22369 ( .A1(n19767), .A2(n19379), .B1(n19765), .B2(n19378), .ZN(
        n19370) );
  AOI22_X1 U22370 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19381), .B1(
        n19766), .B2(n19380), .ZN(n19369) );
  OAI211_X1 U22371 ( .C1(n19770), .C2(n19387), .A(n19370), .B(n19369), .ZN(
        P2_U3075) );
  AOI22_X1 U22372 ( .A1(n19773), .A2(n19410), .B1(n19378), .B2(n19771), .ZN(
        n19372) );
  AOI22_X1 U22373 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19381), .B1(
        n19772), .B2(n19380), .ZN(n19371) );
  OAI211_X1 U22374 ( .C1(n19776), .C2(n19373), .A(n19372), .B(n19371), .ZN(
        P2_U3076) );
  AOI22_X1 U22375 ( .A1(n19719), .A2(n19379), .B1(n19378), .B2(n19777), .ZN(
        n19375) );
  AOI22_X1 U22376 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19381), .B1(
        n19778), .B2(n19380), .ZN(n19374) );
  OAI211_X1 U22377 ( .C1(n19722), .C2(n19387), .A(n19375), .B(n19374), .ZN(
        P2_U3077) );
  AOI22_X1 U22378 ( .A1(n19787), .A2(n19379), .B1(n19378), .B2(n19785), .ZN(
        n19377) );
  AOI22_X1 U22379 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19381), .B1(
        n19786), .B2(n19380), .ZN(n19376) );
  OAI211_X1 U22380 ( .C1(n19790), .C2(n19387), .A(n19377), .B(n19376), .ZN(
        P2_U3078) );
  AOI22_X1 U22381 ( .A1(n19795), .A2(n19379), .B1(n19378), .B2(n19792), .ZN(
        n19383) );
  AOI22_X1 U22382 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19381), .B1(
        n19793), .B2(n19380), .ZN(n19382) );
  OAI211_X1 U22383 ( .C1(n19801), .C2(n19387), .A(n19383), .B(n19382), .ZN(
        P2_U3079) );
  OR2_X1 U22384 ( .A1(n19449), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19421) );
  NOR2_X1 U22385 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19421), .ZN(
        n19408) );
  NOR3_X1 U22386 ( .A1(n19384), .A2(n19408), .A3(n19735), .ZN(n19388) );
  AND3_X1 U22387 ( .A1(n19385), .A2(n19450), .A3(n19898), .ZN(n19393) );
  AOI21_X1 U22388 ( .B1(n19393), .B2(n19917), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19386) );
  AOI22_X1 U22389 ( .A1(n19409), .A2(n19741), .B1(n19740), .B2(n19408), .ZN(
        n19395) );
  AOI21_X1 U22390 ( .B1(n19387), .B2(n19433), .A(n19573), .ZN(n19392) );
  INV_X1 U22391 ( .A(n19408), .ZN(n19390) );
  AOI211_X1 U22392 ( .C1(P2_STATE2_REG_3__SCAN_IN), .C2(n19390), .A(n19389), 
        .B(n19388), .ZN(n19391) );
  AOI22_X1 U22393 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n19411), .B1(
        n19410), .B2(n19749), .ZN(n19394) );
  OAI211_X1 U22394 ( .C1(n19752), .C2(n19433), .A(n19395), .B(n19394), .ZN(
        P2_U3080) );
  AOI22_X1 U22395 ( .A1(n19409), .A2(n19754), .B1(n19753), .B2(n19408), .ZN(
        n19397) );
  AOI22_X1 U22396 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19411), .B1(
        n19410), .B2(n19755), .ZN(n19396) );
  OAI211_X1 U22397 ( .C1(n19758), .C2(n19433), .A(n19397), .B(n19396), .ZN(
        P2_U3081) );
  AOI22_X1 U22398 ( .A1(n19409), .A2(n19760), .B1(n19759), .B2(n19408), .ZN(
        n19399) );
  AOI22_X1 U22399 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19411), .B1(
        n19410), .B2(n19761), .ZN(n19398) );
  OAI211_X1 U22400 ( .C1(n19764), .C2(n19433), .A(n19399), .B(n19398), .ZN(
        P2_U3082) );
  AOI22_X1 U22401 ( .A1(n19409), .A2(n19766), .B1(n19765), .B2(n19408), .ZN(
        n19401) );
  AOI22_X1 U22402 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19411), .B1(
        n19410), .B2(n19767), .ZN(n19400) );
  OAI211_X1 U22403 ( .C1(n19770), .C2(n19433), .A(n19401), .B(n19400), .ZN(
        P2_U3083) );
  AOI22_X1 U22404 ( .A1(n19409), .A2(n19772), .B1(n19771), .B2(n19408), .ZN(
        n19403) );
  AOI22_X1 U22405 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19411), .B1(
        n19410), .B2(n19714), .ZN(n19402) );
  OAI211_X1 U22406 ( .C1(n19717), .C2(n19433), .A(n19403), .B(n19402), .ZN(
        P2_U3084) );
  AOI22_X1 U22407 ( .A1(n19409), .A2(n19778), .B1(n19777), .B2(n19408), .ZN(
        n19405) );
  AOI22_X1 U22408 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19411), .B1(
        n19410), .B2(n19719), .ZN(n19404) );
  OAI211_X1 U22409 ( .C1(n19722), .C2(n19433), .A(n19405), .B(n19404), .ZN(
        P2_U3085) );
  AOI22_X1 U22410 ( .A1(n19409), .A2(n19786), .B1(n19785), .B2(n19408), .ZN(
        n19407) );
  AOI22_X1 U22411 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19411), .B1(
        n19410), .B2(n19787), .ZN(n19406) );
  OAI211_X1 U22412 ( .C1(n19790), .C2(n19433), .A(n19407), .B(n19406), .ZN(
        P2_U3086) );
  AOI22_X1 U22413 ( .A1(n19409), .A2(n19793), .B1(n19792), .B2(n19408), .ZN(
        n19413) );
  AOI22_X1 U22414 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19411), .B1(
        n19410), .B2(n19795), .ZN(n19412) );
  OAI211_X1 U22415 ( .C1(n19801), .C2(n19433), .A(n19413), .B(n19412), .ZN(
        P2_U3087) );
  NOR2_X1 U22416 ( .A1(n19449), .A2(n19538), .ZN(n19438) );
  AOI22_X1 U22417 ( .A1(n19749), .A2(n19439), .B1(n19740), .B2(n19438), .ZN(
        n19424) );
  INV_X1 U22418 ( .A(n19658), .ZN(n19664) );
  AOI21_X1 U22419 ( .B1(n19480), .B2(n19664), .A(n19886), .ZN(n19418) );
  INV_X1 U22420 ( .A(n19438), .ZN(n19414) );
  NAND2_X1 U22421 ( .A1(n19415), .A2(n19414), .ZN(n19419) );
  NOR2_X1 U22422 ( .A1(n19419), .A2(n19735), .ZN(n19416) );
  AOI21_X1 U22423 ( .B1(n19418), .B2(n19421), .A(n19416), .ZN(n19417) );
  OAI211_X1 U22424 ( .C1(n19438), .C2(n19917), .A(n19417), .B(n19747), .ZN(
        n19441) );
  INV_X1 U22425 ( .A(n19418), .ZN(n19422) );
  INV_X1 U22426 ( .A(n19419), .ZN(n19420) );
  OAI22_X1 U22427 ( .A1(n19422), .A2(n19421), .B1(n19420), .B2(n19735), .ZN(
        n19440) );
  AOI22_X1 U22428 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n19441), .B1(
        n19741), .B2(n19440), .ZN(n19423) );
  OAI211_X1 U22429 ( .C1(n19752), .C2(n19461), .A(n19424), .B(n19423), .ZN(
        P2_U3088) );
  AOI22_X1 U22430 ( .A1(n19704), .A2(n19472), .B1(n19438), .B2(n19753), .ZN(
        n19426) );
  AOI22_X1 U22431 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19441), .B1(
        n19754), .B2(n19440), .ZN(n19425) );
  OAI211_X1 U22432 ( .C1(n19707), .C2(n19433), .A(n19426), .B(n19425), .ZN(
        P2_U3089) );
  AOI22_X1 U22433 ( .A1(n19761), .A2(n19439), .B1(n19438), .B2(n19759), .ZN(
        n19428) );
  AOI22_X1 U22434 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19441), .B1(
        n19760), .B2(n19440), .ZN(n19427) );
  OAI211_X1 U22435 ( .C1(n19764), .C2(n19461), .A(n19428), .B(n19427), .ZN(
        P2_U3090) );
  AOI22_X1 U22436 ( .A1(n19767), .A2(n19439), .B1(n19765), .B2(n19438), .ZN(
        n19430) );
  AOI22_X1 U22437 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19441), .B1(
        n19766), .B2(n19440), .ZN(n19429) );
  OAI211_X1 U22438 ( .C1(n19770), .C2(n19461), .A(n19430), .B(n19429), .ZN(
        P2_U3091) );
  AOI22_X1 U22439 ( .A1(n19773), .A2(n19472), .B1(n19438), .B2(n19771), .ZN(
        n19432) );
  AOI22_X1 U22440 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19441), .B1(
        n19772), .B2(n19440), .ZN(n19431) );
  OAI211_X1 U22441 ( .C1(n19776), .C2(n19433), .A(n19432), .B(n19431), .ZN(
        P2_U3092) );
  AOI22_X1 U22442 ( .A1(n19719), .A2(n19439), .B1(n19438), .B2(n19777), .ZN(
        n19435) );
  AOI22_X1 U22443 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19441), .B1(
        n19778), .B2(n19440), .ZN(n19434) );
  OAI211_X1 U22444 ( .C1(n19722), .C2(n19461), .A(n19435), .B(n19434), .ZN(
        P2_U3093) );
  AOI22_X1 U22445 ( .A1(n19787), .A2(n19439), .B1(n19438), .B2(n19785), .ZN(
        n19437) );
  AOI22_X1 U22446 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19441), .B1(
        n19786), .B2(n19440), .ZN(n19436) );
  OAI211_X1 U22447 ( .C1(n19790), .C2(n19461), .A(n19437), .B(n19436), .ZN(
        P2_U3094) );
  AOI22_X1 U22448 ( .A1(n19795), .A2(n19439), .B1(n19438), .B2(n19792), .ZN(
        n19443) );
  AOI22_X1 U22449 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19441), .B1(
        n19793), .B2(n19440), .ZN(n19442) );
  OAI211_X1 U22450 ( .C1(n19801), .C2(n19461), .A(n19443), .B(n19442), .ZN(
        P2_U3095) );
  NOR2_X1 U22451 ( .A1(n19449), .A2(n19572), .ZN(n19470) );
  OAI21_X1 U22452 ( .B1(n19444), .B2(n19470), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19445) );
  OAI21_X1 U22453 ( .B1(n19449), .B2(n19446), .A(n19445), .ZN(n19471) );
  AOI22_X1 U22454 ( .A1(n19471), .A2(n19741), .B1(n19740), .B2(n19470), .ZN(
        n19456) );
  OAI21_X1 U22455 ( .B1(n19472), .B2(n19498), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19448) );
  OAI21_X1 U22456 ( .B1(n19450), .B2(n19449), .A(n19448), .ZN(n19454) );
  INV_X1 U22457 ( .A(n19470), .ZN(n19451) );
  OAI211_X1 U22458 ( .C1(n19452), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19886), 
        .B(n19451), .ZN(n19453) );
  NAND3_X1 U22459 ( .A1(n19454), .A2(n19747), .A3(n19453), .ZN(n19473) );
  AOI22_X1 U22460 ( .A1(P2_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n19473), .B1(
        n19498), .B2(n19690), .ZN(n19455) );
  OAI211_X1 U22461 ( .C1(n19703), .C2(n19461), .A(n19456), .B(n19455), .ZN(
        P2_U3096) );
  AOI22_X1 U22462 ( .A1(n19471), .A2(n19754), .B1(n19753), .B2(n19470), .ZN(
        n19458) );
  AOI22_X1 U22463 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19473), .B1(
        n19498), .B2(n19704), .ZN(n19457) );
  OAI211_X1 U22464 ( .C1(n19707), .C2(n19461), .A(n19458), .B(n19457), .ZN(
        P2_U3097) );
  AOI22_X1 U22465 ( .A1(n19471), .A2(n19760), .B1(n19759), .B2(n19470), .ZN(
        n19460) );
  AOI22_X1 U22466 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19473), .B1(
        n19498), .B2(n19708), .ZN(n19459) );
  OAI211_X1 U22467 ( .C1(n19711), .C2(n19461), .A(n19460), .B(n19459), .ZN(
        P2_U3098) );
  AOI22_X1 U22468 ( .A1(n19471), .A2(n19766), .B1(n19765), .B2(n19470), .ZN(
        n19463) );
  AOI22_X1 U22469 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19473), .B1(
        n19472), .B2(n19767), .ZN(n19462) );
  OAI211_X1 U22470 ( .C1(n19770), .C2(n19505), .A(n19463), .B(n19462), .ZN(
        P2_U3099) );
  AOI22_X1 U22471 ( .A1(n19471), .A2(n19772), .B1(n19771), .B2(n19470), .ZN(
        n19465) );
  AOI22_X1 U22472 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19473), .B1(
        n19472), .B2(n19714), .ZN(n19464) );
  OAI211_X1 U22473 ( .C1(n19717), .C2(n19505), .A(n19465), .B(n19464), .ZN(
        P2_U3100) );
  AOI22_X1 U22474 ( .A1(n19471), .A2(n19778), .B1(n19777), .B2(n19470), .ZN(
        n19467) );
  AOI22_X1 U22475 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19473), .B1(
        n19472), .B2(n19719), .ZN(n19466) );
  OAI211_X1 U22476 ( .C1(n19722), .C2(n19505), .A(n19467), .B(n19466), .ZN(
        P2_U3101) );
  AOI22_X1 U22477 ( .A1(n19471), .A2(n19786), .B1(n19785), .B2(n19470), .ZN(
        n19469) );
  AOI22_X1 U22478 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19473), .B1(
        n19472), .B2(n19787), .ZN(n19468) );
  OAI211_X1 U22479 ( .C1(n19790), .C2(n19505), .A(n19469), .B(n19468), .ZN(
        P2_U3102) );
  AOI22_X1 U22480 ( .A1(n19471), .A2(n19793), .B1(n19792), .B2(n19470), .ZN(
        n19475) );
  AOI22_X1 U22481 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19473), .B1(
        n19472), .B2(n19795), .ZN(n19474) );
  OAI211_X1 U22482 ( .C1(n19801), .C2(n19505), .A(n19475), .B(n19474), .ZN(
        P2_U3103) );
  NOR2_X1 U22483 ( .A1(n19737), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19484) );
  INV_X1 U22484 ( .A(n19484), .ZN(n19479) );
  INV_X1 U22485 ( .A(n19482), .ZN(n19477) );
  INV_X1 U22486 ( .A(n19481), .ZN(n19510) );
  OAI21_X1 U22487 ( .B1(n19477), .B2(n19510), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19478) );
  OAI21_X1 U22488 ( .B1(n19479), .B2(n19886), .A(n19478), .ZN(n19501) );
  AOI22_X1 U22489 ( .A1(n19501), .A2(n19741), .B1(n19510), .B2(n19740), .ZN(
        n19487) );
  NAND2_X1 U22490 ( .A1(n19480), .A2(n19742), .ZN(n19887) );
  INV_X1 U22491 ( .A(n19887), .ZN(n19485) );
  OAI211_X1 U22492 ( .C1(n19482), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19481), 
        .B(n19886), .ZN(n19483) );
  OAI211_X1 U22493 ( .C1(n19485), .C2(n19484), .A(n19747), .B(n19483), .ZN(
        n19502) );
  AOI22_X1 U22494 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n19502), .B1(
        n19498), .B2(n19749), .ZN(n19486) );
  OAI211_X1 U22495 ( .C1(n19752), .C2(n19525), .A(n19487), .B(n19486), .ZN(
        P2_U3104) );
  AOI22_X1 U22496 ( .A1(n19501), .A2(n19754), .B1(n19510), .B2(n19753), .ZN(
        n19489) );
  AOI22_X1 U22497 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19502), .B1(
        n19498), .B2(n19755), .ZN(n19488) );
  OAI211_X1 U22498 ( .C1(n19758), .C2(n19525), .A(n19489), .B(n19488), .ZN(
        P2_U3105) );
  AOI22_X1 U22499 ( .A1(n19501), .A2(n19760), .B1(n19510), .B2(n19759), .ZN(
        n19491) );
  AOI22_X1 U22500 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19502), .B1(
        n19531), .B2(n19708), .ZN(n19490) );
  OAI211_X1 U22501 ( .C1(n19711), .C2(n19505), .A(n19491), .B(n19490), .ZN(
        P2_U3106) );
  AOI22_X1 U22502 ( .A1(n19501), .A2(n19766), .B1(n19510), .B2(n19765), .ZN(
        n19493) );
  AOI22_X1 U22503 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19502), .B1(
        n19498), .B2(n19767), .ZN(n19492) );
  OAI211_X1 U22504 ( .C1(n19770), .C2(n19525), .A(n19493), .B(n19492), .ZN(
        P2_U3107) );
  AOI22_X1 U22505 ( .A1(n19501), .A2(n19772), .B1(n19510), .B2(n19771), .ZN(
        n19495) );
  AOI22_X1 U22506 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19502), .B1(
        n19498), .B2(n19714), .ZN(n19494) );
  OAI211_X1 U22507 ( .C1(n19717), .C2(n19525), .A(n19495), .B(n19494), .ZN(
        P2_U3108) );
  AOI22_X1 U22508 ( .A1(n19501), .A2(n19778), .B1(n19510), .B2(n19777), .ZN(
        n19497) );
  AOI22_X1 U22509 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19502), .B1(
        n19498), .B2(n19719), .ZN(n19496) );
  OAI211_X1 U22510 ( .C1(n19722), .C2(n19525), .A(n19497), .B(n19496), .ZN(
        P2_U3109) );
  AOI22_X1 U22511 ( .A1(n19501), .A2(n19786), .B1(n19510), .B2(n19785), .ZN(
        n19500) );
  AOI22_X1 U22512 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19502), .B1(
        n19498), .B2(n19787), .ZN(n19499) );
  OAI211_X1 U22513 ( .C1(n19790), .C2(n19525), .A(n19500), .B(n19499), .ZN(
        P2_U3110) );
  AOI22_X1 U22514 ( .A1(n19501), .A2(n19793), .B1(n19510), .B2(n19792), .ZN(
        n19504) );
  AOI22_X1 U22515 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19502), .B1(
        n19531), .B2(n19728), .ZN(n19503) );
  OAI211_X1 U22516 ( .C1(n19734), .C2(n19505), .A(n19504), .B(n19503), .ZN(
        P2_U3111) );
  NAND2_X1 U22517 ( .A1(n19905), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19608) );
  NOR2_X1 U22518 ( .A1(n19608), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19544) );
  INV_X1 U22519 ( .A(n19544), .ZN(n19547) );
  NOR2_X1 U22520 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19547), .ZN(
        n19530) );
  AOI22_X1 U22521 ( .A1(n19749), .A2(n19531), .B1(n19740), .B2(n19530), .ZN(
        n19516) );
  OAI21_X1 U22522 ( .B1(n19553), .B2(n19531), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19506) );
  NAND2_X1 U22523 ( .A1(n19506), .A2(n19691), .ZN(n19514) );
  NOR2_X1 U22524 ( .A1(n19514), .A2(n19510), .ZN(n19507) );
  AOI211_X1 U22525 ( .C1(P2_STATE2_REG_2__SCAN_IN), .C2(n19508), .A(
        P2_STATE2_REG_3__SCAN_IN), .B(n19507), .ZN(n19509) );
  NOR2_X1 U22526 ( .A1(n19510), .A2(n19530), .ZN(n19513) );
  OAI21_X1 U22527 ( .B1(n19511), .B2(n19530), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19512) );
  AOI22_X1 U22528 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19533), .B1(
        n19741), .B2(n19532), .ZN(n19515) );
  OAI211_X1 U22529 ( .C1(n19752), .C2(n19569), .A(n19516), .B(n19515), .ZN(
        P2_U3112) );
  AOI22_X1 U22530 ( .A1(n19704), .A2(n19553), .B1(n19753), .B2(n19530), .ZN(
        n19518) );
  AOI22_X1 U22531 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19533), .B1(
        n19754), .B2(n19532), .ZN(n19517) );
  OAI211_X1 U22532 ( .C1(n19707), .C2(n19525), .A(n19518), .B(n19517), .ZN(
        P2_U3113) );
  AOI22_X1 U22533 ( .A1(n19761), .A2(n19531), .B1(n19759), .B2(n19530), .ZN(
        n19520) );
  AOI22_X1 U22534 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19533), .B1(
        n19760), .B2(n19532), .ZN(n19519) );
  OAI211_X1 U22535 ( .C1(n19764), .C2(n19569), .A(n19520), .B(n19519), .ZN(
        P2_U3114) );
  AOI22_X1 U22536 ( .A1(n19767), .A2(n19531), .B1(n19765), .B2(n19530), .ZN(
        n19522) );
  AOI22_X1 U22537 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19533), .B1(
        n19766), .B2(n19532), .ZN(n19521) );
  OAI211_X1 U22538 ( .C1(n19770), .C2(n19569), .A(n19522), .B(n19521), .ZN(
        P2_U3115) );
  AOI22_X1 U22539 ( .A1(n19773), .A2(n19553), .B1(n19771), .B2(n19530), .ZN(
        n19524) );
  AOI22_X1 U22540 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19533), .B1(
        n19772), .B2(n19532), .ZN(n19523) );
  OAI211_X1 U22541 ( .C1(n19776), .C2(n19525), .A(n19524), .B(n19523), .ZN(
        P2_U3116) );
  AOI22_X1 U22542 ( .A1(n19719), .A2(n19531), .B1(n19777), .B2(n19530), .ZN(
        n19527) );
  AOI22_X1 U22543 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19533), .B1(
        n19778), .B2(n19532), .ZN(n19526) );
  OAI211_X1 U22544 ( .C1(n19722), .C2(n19569), .A(n19527), .B(n19526), .ZN(
        P2_U3117) );
  AOI22_X1 U22545 ( .A1(n19787), .A2(n19531), .B1(n19785), .B2(n19530), .ZN(
        n19529) );
  AOI22_X1 U22546 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19533), .B1(
        n19786), .B2(n19532), .ZN(n19528) );
  OAI211_X1 U22547 ( .C1(n19790), .C2(n19569), .A(n19529), .B(n19528), .ZN(
        P2_U3118) );
  AOI22_X1 U22548 ( .A1(n19795), .A2(n19531), .B1(n19792), .B2(n19530), .ZN(
        n19535) );
  AOI22_X1 U22549 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19533), .B1(
        n19793), .B2(n19532), .ZN(n19534) );
  OAI211_X1 U22550 ( .C1(n19801), .C2(n19569), .A(n19535), .B(n19534), .ZN(
        P2_U3119) );
  NOR2_X1 U22551 ( .A1(n19538), .A2(n19608), .ZN(n19564) );
  AOI22_X1 U22552 ( .A1(n19749), .A2(n19553), .B1(n19740), .B2(n19564), .ZN(
        n19550) );
  INV_X1 U22553 ( .A(n19539), .ZN(n19894) );
  NAND2_X1 U22554 ( .A1(n19894), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19663) );
  OAI21_X1 U22555 ( .B1(n19663), .B2(n19540), .A(n19691), .ZN(n19548) );
  INV_X1 U22556 ( .A(n19564), .ZN(n19541) );
  OAI211_X1 U22557 ( .C1(n19542), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19886), 
        .B(n19541), .ZN(n19543) );
  OAI211_X1 U22558 ( .C1(n19548), .C2(n19544), .A(n19747), .B(n19543), .ZN(
        n19566) );
  OAI21_X1 U22559 ( .B1(n19545), .B2(n19564), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19546) );
  OAI21_X1 U22560 ( .B1(n19548), .B2(n19547), .A(n19546), .ZN(n19565) );
  AOI22_X1 U22561 ( .A1(P2_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n19566), .B1(
        n19741), .B2(n19565), .ZN(n19549) );
  OAI211_X1 U22562 ( .C1(n19752), .C2(n19604), .A(n19550), .B(n19549), .ZN(
        P2_U3120) );
  AOI22_X1 U22563 ( .A1(n19755), .A2(n19553), .B1(n19753), .B2(n19564), .ZN(
        n19552) );
  AOI22_X1 U22564 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19566), .B1(
        n19754), .B2(n19565), .ZN(n19551) );
  OAI211_X1 U22565 ( .C1(n19758), .C2(n19604), .A(n19552), .B(n19551), .ZN(
        P2_U3121) );
  AOI22_X1 U22566 ( .A1(n19761), .A2(n19553), .B1(n19759), .B2(n19564), .ZN(
        n19555) );
  AOI22_X1 U22567 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19566), .B1(
        n19760), .B2(n19565), .ZN(n19554) );
  OAI211_X1 U22568 ( .C1(n19764), .C2(n19604), .A(n19555), .B(n19554), .ZN(
        P2_U3122) );
  AOI22_X1 U22569 ( .A1(n19620), .A2(n19595), .B1(n19765), .B2(n19564), .ZN(
        n19557) );
  AOI22_X1 U22570 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19566), .B1(
        n19766), .B2(n19565), .ZN(n19556) );
  OAI211_X1 U22571 ( .C1(n19623), .C2(n19569), .A(n19557), .B(n19556), .ZN(
        P2_U3123) );
  AOI22_X1 U22572 ( .A1(n19595), .A2(n19773), .B1(n19771), .B2(n19564), .ZN(
        n19559) );
  AOI22_X1 U22573 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19566), .B1(
        n19772), .B2(n19565), .ZN(n19558) );
  OAI211_X1 U22574 ( .C1(n19776), .C2(n19569), .A(n19559), .B(n19558), .ZN(
        P2_U3124) );
  AOI22_X1 U22575 ( .A1(n19779), .A2(n19595), .B1(n19777), .B2(n19564), .ZN(
        n19561) );
  AOI22_X1 U22576 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19566), .B1(
        n19778), .B2(n19565), .ZN(n19560) );
  OAI211_X1 U22577 ( .C1(n19784), .C2(n19569), .A(n19561), .B(n19560), .ZN(
        P2_U3125) );
  AOI22_X1 U22578 ( .A1(n19723), .A2(n19595), .B1(n19785), .B2(n19564), .ZN(
        n19563) );
  AOI22_X1 U22579 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19566), .B1(
        n19786), .B2(n19565), .ZN(n19562) );
  OAI211_X1 U22580 ( .C1(n19726), .C2(n19569), .A(n19563), .B(n19562), .ZN(
        P2_U3126) );
  AOI22_X1 U22581 ( .A1(n19728), .A2(n19595), .B1(n19792), .B2(n19564), .ZN(
        n19568) );
  AOI22_X1 U22582 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19566), .B1(
        n19793), .B2(n19565), .ZN(n19567) );
  OAI211_X1 U22583 ( .C1(n19734), .C2(n19569), .A(n19568), .B(n19567), .ZN(
        P2_U3127) );
  INV_X1 U22584 ( .A(n19689), .ZN(n19571) );
  INV_X1 U22585 ( .A(n19889), .ZN(n19570) );
  NOR2_X1 U22586 ( .A1(n19572), .A2(n19608), .ZN(n19598) );
  AOI22_X1 U22587 ( .A1(n19690), .A2(n19599), .B1(n19740), .B2(n19598), .ZN(
        n19584) );
  NOR2_X1 U22588 ( .A1(n19599), .A2(n19595), .ZN(n19574) );
  OAI21_X1 U22589 ( .B1(n19574), .B2(n19573), .A(n19691), .ZN(n19582) );
  INV_X1 U22590 ( .A(n19608), .ZN(n19605) );
  AND2_X1 U22591 ( .A1(n19575), .A2(n19605), .ZN(n19578) );
  INV_X1 U22592 ( .A(n19598), .ZN(n19576) );
  OAI211_X1 U22593 ( .C1(n12064), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19886), 
        .B(n19576), .ZN(n19577) );
  OAI211_X1 U22594 ( .C1(n19582), .C2(n19578), .A(n19747), .B(n19577), .ZN(
        n19601) );
  INV_X1 U22595 ( .A(n19578), .ZN(n19581) );
  OAI21_X1 U22596 ( .B1(n19579), .B2(n19598), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19580) );
  AOI22_X1 U22597 ( .A1(P2_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19601), .B1(
        n19741), .B2(n19600), .ZN(n19583) );
  OAI211_X1 U22598 ( .C1(n19703), .C2(n19604), .A(n19584), .B(n19583), .ZN(
        P2_U3128) );
  AOI22_X1 U22599 ( .A1(n19599), .A2(n19704), .B1(n19753), .B2(n19598), .ZN(
        n19586) );
  AOI22_X1 U22600 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19601), .B1(
        n19754), .B2(n19600), .ZN(n19585) );
  OAI211_X1 U22601 ( .C1(n19707), .C2(n19604), .A(n19586), .B(n19585), .ZN(
        P2_U3129) );
  AOI22_X1 U22602 ( .A1(n19595), .A2(n19761), .B1(n19759), .B2(n19598), .ZN(
        n19588) );
  AOI22_X1 U22603 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19601), .B1(
        n19760), .B2(n19600), .ZN(n19587) );
  OAI211_X1 U22604 ( .C1(n19764), .C2(n19635), .A(n19588), .B(n19587), .ZN(
        P2_U3130) );
  AOI22_X1 U22605 ( .A1(n19595), .A2(n19767), .B1(n19765), .B2(n19598), .ZN(
        n19590) );
  AOI22_X1 U22606 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19601), .B1(
        n19766), .B2(n19600), .ZN(n19589) );
  OAI211_X1 U22607 ( .C1(n19770), .C2(n19635), .A(n19590), .B(n19589), .ZN(
        P2_U3131) );
  AOI22_X1 U22608 ( .A1(n19599), .A2(n19773), .B1(n19771), .B2(n19598), .ZN(
        n19592) );
  AOI22_X1 U22609 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19601), .B1(
        n19772), .B2(n19600), .ZN(n19591) );
  OAI211_X1 U22610 ( .C1(n19776), .C2(n19604), .A(n19592), .B(n19591), .ZN(
        P2_U3132) );
  AOI22_X1 U22611 ( .A1(n19595), .A2(n19719), .B1(n19777), .B2(n19598), .ZN(
        n19594) );
  AOI22_X1 U22612 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19601), .B1(
        n19778), .B2(n19600), .ZN(n19593) );
  OAI211_X1 U22613 ( .C1(n19722), .C2(n19635), .A(n19594), .B(n19593), .ZN(
        P2_U3133) );
  AOI22_X1 U22614 ( .A1(n19595), .A2(n19787), .B1(n19785), .B2(n19598), .ZN(
        n19597) );
  AOI22_X1 U22615 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19601), .B1(
        n19786), .B2(n19600), .ZN(n19596) );
  OAI211_X1 U22616 ( .C1(n19790), .C2(n19635), .A(n19597), .B(n19596), .ZN(
        P2_U3134) );
  AOI22_X1 U22617 ( .A1(n19728), .A2(n19599), .B1(n19792), .B2(n19598), .ZN(
        n19603) );
  AOI22_X1 U22618 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19601), .B1(
        n19793), .B2(n19600), .ZN(n19602) );
  OAI211_X1 U22619 ( .C1(n19734), .C2(n19604), .A(n19603), .B(n19602), .ZN(
        P2_U3135) );
  AND2_X1 U22620 ( .A1(n19606), .A2(n19605), .ZN(n19630) );
  NOR2_X1 U22621 ( .A1(n19630), .A2(n19735), .ZN(n19607) );
  NAND2_X1 U22622 ( .A1(n12085), .A2(n19607), .ZN(n19611) );
  OR2_X1 U22623 ( .A1(n19914), .A2(n19608), .ZN(n19610) );
  OAI21_X1 U22624 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19610), .A(n19735), 
        .ZN(n19609) );
  AOI22_X1 U22625 ( .A1(n19631), .A2(n19741), .B1(n19740), .B2(n19630), .ZN(
        n19615) );
  OAI21_X1 U22626 ( .B1(n19663), .B2(n19889), .A(n19610), .ZN(n19612) );
  AND2_X1 U22627 ( .A1(n19612), .A2(n19611), .ZN(n19613) );
  OAI211_X1 U22628 ( .C1(n19630), .C2(n19917), .A(n19613), .B(n19747), .ZN(
        n19632) );
  AOI22_X1 U22629 ( .A1(P2_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19632), .B1(
        n19654), .B2(n19690), .ZN(n19614) );
  OAI211_X1 U22630 ( .C1(n19703), .C2(n19635), .A(n19615), .B(n19614), .ZN(
        P2_U3136) );
  AOI22_X1 U22631 ( .A1(n19631), .A2(n19754), .B1(n19753), .B2(n19630), .ZN(
        n19617) );
  AOI22_X1 U22632 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19632), .B1(
        n19654), .B2(n19704), .ZN(n19616) );
  OAI211_X1 U22633 ( .C1(n19707), .C2(n19635), .A(n19617), .B(n19616), .ZN(
        P2_U3137) );
  AOI22_X1 U22634 ( .A1(n19631), .A2(n19760), .B1(n19759), .B2(n19630), .ZN(
        n19619) );
  AOI22_X1 U22635 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19632), .B1(
        n19654), .B2(n19708), .ZN(n19618) );
  OAI211_X1 U22636 ( .C1(n19711), .C2(n19635), .A(n19619), .B(n19618), .ZN(
        P2_U3138) );
  AOI22_X1 U22637 ( .A1(n19631), .A2(n19766), .B1(n19765), .B2(n19630), .ZN(
        n19622) );
  AOI22_X1 U22638 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19632), .B1(
        n19654), .B2(n19620), .ZN(n19621) );
  OAI211_X1 U22639 ( .C1(n19623), .C2(n19635), .A(n19622), .B(n19621), .ZN(
        P2_U3139) );
  AOI22_X1 U22640 ( .A1(n19631), .A2(n19772), .B1(n19771), .B2(n19630), .ZN(
        n19625) );
  AOI22_X1 U22641 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19632), .B1(
        n19654), .B2(n19773), .ZN(n19624) );
  OAI211_X1 U22642 ( .C1(n19776), .C2(n19635), .A(n19625), .B(n19624), .ZN(
        P2_U3140) );
  AOI22_X1 U22643 ( .A1(n19631), .A2(n19778), .B1(n19777), .B2(n19630), .ZN(
        n19627) );
  AOI22_X1 U22644 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19632), .B1(
        n19654), .B2(n19779), .ZN(n19626) );
  OAI211_X1 U22645 ( .C1(n19784), .C2(n19635), .A(n19627), .B(n19626), .ZN(
        P2_U3141) );
  AOI22_X1 U22646 ( .A1(n19631), .A2(n19786), .B1(n19785), .B2(n19630), .ZN(
        n19629) );
  AOI22_X1 U22647 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19632), .B1(
        n19654), .B2(n19723), .ZN(n19628) );
  OAI211_X1 U22648 ( .C1(n19726), .C2(n19635), .A(n19629), .B(n19628), .ZN(
        P2_U3142) );
  AOI22_X1 U22649 ( .A1(n19631), .A2(n19793), .B1(n19792), .B2(n19630), .ZN(
        n19634) );
  AOI22_X1 U22650 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19632), .B1(
        n19654), .B2(n19728), .ZN(n19633) );
  OAI211_X1 U22651 ( .C1(n19734), .C2(n19635), .A(n19634), .B(n19633), .ZN(
        P2_U3143) );
  INV_X1 U22652 ( .A(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n19638) );
  AOI22_X1 U22653 ( .A1(n19653), .A2(n19741), .B1(n19652), .B2(n19740), .ZN(
        n19637) );
  AOI22_X1 U22654 ( .A1(n19654), .A2(n19749), .B1(n19684), .B2(n19690), .ZN(
        n19636) );
  OAI211_X1 U22655 ( .C1(n19657), .C2(n19638), .A(n19637), .B(n19636), .ZN(
        P2_U3144) );
  INV_X1 U22656 ( .A(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n19641) );
  AOI22_X1 U22657 ( .A1(n19653), .A2(n19754), .B1(n19652), .B2(n19753), .ZN(
        n19640) );
  AOI22_X1 U22658 ( .A1(n19684), .A2(n19704), .B1(n19654), .B2(n19755), .ZN(
        n19639) );
  OAI211_X1 U22659 ( .C1(n19657), .C2(n19641), .A(n19640), .B(n19639), .ZN(
        P2_U3145) );
  INV_X1 U22660 ( .A(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n19644) );
  AOI22_X1 U22661 ( .A1(n19653), .A2(n19760), .B1(n19652), .B2(n19759), .ZN(
        n19643) );
  AOI22_X1 U22662 ( .A1(n19654), .A2(n19761), .B1(n19684), .B2(n19708), .ZN(
        n19642) );
  OAI211_X1 U22663 ( .C1(n19657), .C2(n19644), .A(n19643), .B(n19642), .ZN(
        P2_U3146) );
  INV_X1 U22664 ( .A(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n19647) );
  AOI22_X1 U22665 ( .A1(n19653), .A2(n19772), .B1(n19652), .B2(n19771), .ZN(
        n19646) );
  AOI22_X1 U22666 ( .A1(n19684), .A2(n19773), .B1(n19654), .B2(n19714), .ZN(
        n19645) );
  OAI211_X1 U22667 ( .C1(n19657), .C2(n19647), .A(n19646), .B(n19645), .ZN(
        P2_U3148) );
  AOI22_X1 U22668 ( .A1(n19653), .A2(n19778), .B1(n19652), .B2(n19777), .ZN(
        n19649) );
  AOI22_X1 U22669 ( .A1(n19654), .A2(n19719), .B1(n19684), .B2(n19779), .ZN(
        n19648) );
  OAI211_X1 U22670 ( .C1(n19657), .C2(n12073), .A(n19649), .B(n19648), .ZN(
        P2_U3149) );
  AOI22_X1 U22671 ( .A1(n19653), .A2(n19786), .B1(n19652), .B2(n19785), .ZN(
        n19651) );
  AOI22_X1 U22672 ( .A1(n19654), .A2(n19787), .B1(n19684), .B2(n19723), .ZN(
        n19650) );
  OAI211_X1 U22673 ( .C1(n19657), .C2(n12139), .A(n19651), .B(n19650), .ZN(
        P2_U3150) );
  AOI22_X1 U22674 ( .A1(n19653), .A2(n19793), .B1(n19652), .B2(n19792), .ZN(
        n19656) );
  AOI22_X1 U22675 ( .A1(n19654), .A2(n19795), .B1(n19684), .B2(n19728), .ZN(
        n19655) );
  OAI211_X1 U22676 ( .C1(n19657), .C2(n11728), .A(n19656), .B(n19655), .ZN(
        P2_U3151) );
  NOR2_X1 U22677 ( .A1(n19924), .A2(n19666), .ZN(n19693) );
  NOR3_X1 U22678 ( .A1(n19660), .A2(n19693), .A3(n19735), .ZN(n19665) );
  INV_X1 U22679 ( .A(n19666), .ZN(n19661) );
  AOI21_X1 U22680 ( .B1(n19917), .B2(n19661), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19662) );
  AOI22_X1 U22681 ( .A1(n19683), .A2(n19741), .B1(n19740), .B2(n19693), .ZN(
        n19670) );
  INV_X1 U22682 ( .A(n19663), .ZN(n19743) );
  NAND2_X1 U22683 ( .A1(n19743), .A2(n19664), .ZN(n19667) );
  AOI21_X1 U22684 ( .B1(n19667), .B2(n19666), .A(n19665), .ZN(n19668) );
  OAI211_X1 U22685 ( .C1(n19693), .C2(n19917), .A(n19668), .B(n19747), .ZN(
        n19685) );
  AOI22_X1 U22686 ( .A1(P2_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n19685), .B1(
        n19684), .B2(n19749), .ZN(n19669) );
  OAI211_X1 U22687 ( .C1(n19752), .C2(n19733), .A(n19670), .B(n19669), .ZN(
        P2_U3152) );
  AOI22_X1 U22688 ( .A1(n19683), .A2(n19754), .B1(n19753), .B2(n19693), .ZN(
        n19672) );
  AOI22_X1 U22689 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19685), .B1(
        n19684), .B2(n19755), .ZN(n19671) );
  OAI211_X1 U22690 ( .C1(n19758), .C2(n19733), .A(n19672), .B(n19671), .ZN(
        P2_U3153) );
  AOI22_X1 U22691 ( .A1(n19683), .A2(n19760), .B1(n19759), .B2(n19693), .ZN(
        n19674) );
  AOI22_X1 U22692 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19685), .B1(
        n19684), .B2(n19761), .ZN(n19673) );
  OAI211_X1 U22693 ( .C1(n19764), .C2(n19733), .A(n19674), .B(n19673), .ZN(
        P2_U3154) );
  AOI22_X1 U22694 ( .A1(n19683), .A2(n19766), .B1(n19765), .B2(n19693), .ZN(
        n19676) );
  AOI22_X1 U22695 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19685), .B1(
        n19684), .B2(n19767), .ZN(n19675) );
  OAI211_X1 U22696 ( .C1(n19770), .C2(n19733), .A(n19676), .B(n19675), .ZN(
        P2_U3155) );
  AOI22_X1 U22697 ( .A1(n19683), .A2(n19772), .B1(n19771), .B2(n19693), .ZN(
        n19678) );
  AOI22_X1 U22698 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19685), .B1(
        n19684), .B2(n19714), .ZN(n19677) );
  OAI211_X1 U22699 ( .C1(n19717), .C2(n19733), .A(n19678), .B(n19677), .ZN(
        P2_U3156) );
  AOI22_X1 U22700 ( .A1(n19683), .A2(n19778), .B1(n19777), .B2(n19693), .ZN(
        n19680) );
  AOI22_X1 U22701 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19685), .B1(
        n19684), .B2(n19719), .ZN(n19679) );
  OAI211_X1 U22702 ( .C1(n19722), .C2(n19733), .A(n19680), .B(n19679), .ZN(
        P2_U3157) );
  AOI22_X1 U22703 ( .A1(n19683), .A2(n19786), .B1(n19785), .B2(n19693), .ZN(
        n19682) );
  AOI22_X1 U22704 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19685), .B1(
        n19684), .B2(n19787), .ZN(n19681) );
  OAI211_X1 U22705 ( .C1(n19790), .C2(n19733), .A(n19682), .B(n19681), .ZN(
        P2_U3158) );
  AOI22_X1 U22706 ( .A1(n19683), .A2(n19793), .B1(n19792), .B2(n19693), .ZN(
        n19687) );
  AOI22_X1 U22707 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n19685), .B1(
        n19684), .B2(n19795), .ZN(n19686) );
  OAI211_X1 U22708 ( .C1(n19801), .C2(n19733), .A(n19687), .B(n19686), .ZN(
        P2_U3159) );
  NOR3_X2 U22709 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19898), .A3(
        n19737), .ZN(n19727) );
  AOI22_X1 U22710 ( .A1(n19690), .A2(n19796), .B1(n19740), .B2(n19727), .ZN(
        n19702) );
  OAI21_X1 U22711 ( .B1(n19796), .B2(n19718), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19692) );
  NAND2_X1 U22712 ( .A1(n19692), .A2(n19691), .ZN(n19700) );
  NOR2_X1 U22713 ( .A1(n19727), .A2(n19693), .ZN(n19699) );
  INV_X1 U22714 ( .A(n19699), .ZN(n19696) );
  INV_X1 U22715 ( .A(n19727), .ZN(n19694) );
  OAI211_X1 U22716 ( .C1(n12063), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19886), 
        .B(n19694), .ZN(n19695) );
  OAI211_X1 U22717 ( .C1(n19700), .C2(n19696), .A(n19747), .B(n19695), .ZN(
        n19730) );
  OAI21_X1 U22718 ( .B1(n19697), .B2(n19727), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19698) );
  AOI22_X1 U22719 ( .A1(P2_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n19730), .B1(
        n19741), .B2(n19729), .ZN(n19701) );
  OAI211_X1 U22720 ( .C1(n19703), .C2(n19733), .A(n19702), .B(n19701), .ZN(
        P2_U3160) );
  AOI22_X1 U22721 ( .A1(n19704), .A2(n19796), .B1(n19753), .B2(n19727), .ZN(
        n19706) );
  AOI22_X1 U22722 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n19730), .B1(
        n19754), .B2(n19729), .ZN(n19705) );
  OAI211_X1 U22723 ( .C1(n19707), .C2(n19733), .A(n19706), .B(n19705), .ZN(
        P2_U3161) );
  AOI22_X1 U22724 ( .A1(n19708), .A2(n19796), .B1(n19759), .B2(n19727), .ZN(
        n19710) );
  AOI22_X1 U22725 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n19730), .B1(
        n19760), .B2(n19729), .ZN(n19709) );
  OAI211_X1 U22726 ( .C1(n19711), .C2(n19733), .A(n19710), .B(n19709), .ZN(
        P2_U3162) );
  INV_X1 U22727 ( .A(n19796), .ZN(n19783) );
  AOI22_X1 U22728 ( .A1(n19718), .A2(n19767), .B1(n19765), .B2(n19727), .ZN(
        n19713) );
  AOI22_X1 U22729 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n19730), .B1(
        n19766), .B2(n19729), .ZN(n19712) );
  OAI211_X1 U22730 ( .C1(n19770), .C2(n19783), .A(n19713), .B(n19712), .ZN(
        P2_U3163) );
  AOI22_X1 U22731 ( .A1(n19714), .A2(n19718), .B1(n19771), .B2(n19727), .ZN(
        n19716) );
  AOI22_X1 U22732 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n19730), .B1(
        n19772), .B2(n19729), .ZN(n19715) );
  OAI211_X1 U22733 ( .C1(n19717), .C2(n19783), .A(n19716), .B(n19715), .ZN(
        P2_U3164) );
  AOI22_X1 U22734 ( .A1(n19719), .A2(n19718), .B1(n19777), .B2(n19727), .ZN(
        n19721) );
  AOI22_X1 U22735 ( .A1(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n19730), .B1(
        n19778), .B2(n19729), .ZN(n19720) );
  OAI211_X1 U22736 ( .C1(n19722), .C2(n19783), .A(n19721), .B(n19720), .ZN(
        P2_U3165) );
  AOI22_X1 U22737 ( .A1(n19723), .A2(n19796), .B1(n19785), .B2(n19727), .ZN(
        n19725) );
  AOI22_X1 U22738 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n19730), .B1(
        n19786), .B2(n19729), .ZN(n19724) );
  OAI211_X1 U22739 ( .C1(n19726), .C2(n19733), .A(n19725), .B(n19724), .ZN(
        P2_U3166) );
  AOI22_X1 U22740 ( .A1(n19728), .A2(n19796), .B1(n19792), .B2(n19727), .ZN(
        n19732) );
  AOI22_X1 U22741 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n19730), .B1(
        n19793), .B2(n19729), .ZN(n19731) );
  OAI211_X1 U22742 ( .C1(n19734), .C2(n19733), .A(n19732), .B(n19731), .ZN(
        P2_U3167) );
  INV_X1 U22743 ( .A(n12080), .ZN(n19736) );
  NOR3_X1 U22744 ( .A1(n19736), .A2(n19791), .A3(n19735), .ZN(n19744) );
  OR2_X1 U22745 ( .A1(n19898), .A2(n19737), .ZN(n19745) );
  INV_X1 U22746 ( .A(n19745), .ZN(n19738) );
  AOI21_X1 U22747 ( .B1(n19917), .B2(n19738), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19739) );
  AOI22_X1 U22748 ( .A1(n19794), .A2(n19741), .B1(n19740), .B2(n19791), .ZN(
        n19751) );
  NAND2_X1 U22749 ( .A1(n19743), .A2(n19742), .ZN(n19746) );
  AOI21_X1 U22750 ( .B1(n19746), .B2(n19745), .A(n19744), .ZN(n19748) );
  OAI211_X1 U22751 ( .C1(n19791), .C2(n19917), .A(n19748), .B(n19747), .ZN(
        n19797) );
  AOI22_X1 U22752 ( .A1(P2_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n19797), .B1(
        n19796), .B2(n19749), .ZN(n19750) );
  OAI211_X1 U22753 ( .C1(n19752), .C2(n19800), .A(n19751), .B(n19750), .ZN(
        P2_U3168) );
  AOI22_X1 U22754 ( .A1(n19794), .A2(n19754), .B1(n19753), .B2(n19791), .ZN(
        n19757) );
  AOI22_X1 U22755 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n19797), .B1(
        n19796), .B2(n19755), .ZN(n19756) );
  OAI211_X1 U22756 ( .C1(n19758), .C2(n19800), .A(n19757), .B(n19756), .ZN(
        P2_U3169) );
  AOI22_X1 U22757 ( .A1(n19794), .A2(n19760), .B1(n19759), .B2(n19791), .ZN(
        n19763) );
  AOI22_X1 U22758 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n19797), .B1(
        n19796), .B2(n19761), .ZN(n19762) );
  OAI211_X1 U22759 ( .C1(n19764), .C2(n19800), .A(n19763), .B(n19762), .ZN(
        P2_U3170) );
  AOI22_X1 U22760 ( .A1(n19794), .A2(n19766), .B1(n19765), .B2(n19791), .ZN(
        n19769) );
  AOI22_X1 U22761 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n19797), .B1(
        n19796), .B2(n19767), .ZN(n19768) );
  OAI211_X1 U22762 ( .C1(n19770), .C2(n19800), .A(n19769), .B(n19768), .ZN(
        P2_U3171) );
  AOI22_X1 U22763 ( .A1(n19794), .A2(n19772), .B1(n19771), .B2(n19791), .ZN(
        n19775) );
  AOI22_X1 U22764 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n19797), .B1(
        n19780), .B2(n19773), .ZN(n19774) );
  OAI211_X1 U22765 ( .C1(n19776), .C2(n19783), .A(n19775), .B(n19774), .ZN(
        P2_U3172) );
  AOI22_X1 U22766 ( .A1(n19794), .A2(n19778), .B1(n19777), .B2(n19791), .ZN(
        n19782) );
  AOI22_X1 U22767 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n19797), .B1(
        n19780), .B2(n19779), .ZN(n19781) );
  OAI211_X1 U22768 ( .C1(n19784), .C2(n19783), .A(n19782), .B(n19781), .ZN(
        P2_U3173) );
  AOI22_X1 U22769 ( .A1(n19794), .A2(n19786), .B1(n19785), .B2(n19791), .ZN(
        n19789) );
  AOI22_X1 U22770 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n19797), .B1(
        n19796), .B2(n19787), .ZN(n19788) );
  OAI211_X1 U22771 ( .C1(n19790), .C2(n19800), .A(n19789), .B(n19788), .ZN(
        P2_U3174) );
  AOI22_X1 U22772 ( .A1(n19794), .A2(n19793), .B1(n19792), .B2(n19791), .ZN(
        n19799) );
  AOI22_X1 U22773 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n19797), .B1(
        n19796), .B2(n19795), .ZN(n19798) );
  OAI211_X1 U22774 ( .C1(n19801), .C2(n19800), .A(n19799), .B(n19798), .ZN(
        P2_U3175) );
  NOR3_X1 U22775 ( .A1(n19812), .A2(n19890), .A3(n13537), .ZN(n19806) );
  AOI211_X1 U22776 ( .C1(n19807), .C2(n19804), .A(n19803), .B(n19802), .ZN(
        n19805) );
  AOI221_X1 U22777 ( .B1(n19808), .B2(n19807), .C1(n19806), .C2(n19807), .A(
        n19805), .ZN(n19810) );
  NAND2_X1 U22778 ( .A1(n19810), .A2(n19809), .ZN(P2_U3177) );
  AND2_X1 U22779 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n19811), .ZN(
        P2_U3179) );
  AND2_X1 U22780 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n19811), .ZN(
        P2_U3180) );
  AND2_X1 U22781 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n19811), .ZN(
        P2_U3181) );
  AND2_X1 U22782 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n19811), .ZN(
        P2_U3182) );
  AND2_X1 U22783 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n19811), .ZN(
        P2_U3183) );
  AND2_X1 U22784 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n19811), .ZN(
        P2_U3184) );
  AND2_X1 U22785 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n19811), .ZN(
        P2_U3185) );
  AND2_X1 U22786 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n19811), .ZN(
        P2_U3186) );
  AND2_X1 U22787 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n19811), .ZN(
        P2_U3187) );
  AND2_X1 U22788 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n19811), .ZN(
        P2_U3188) );
  AND2_X1 U22789 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n19811), .ZN(
        P2_U3189) );
  AND2_X1 U22790 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n19811), .ZN(
        P2_U3190) );
  AND2_X1 U22791 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n19811), .ZN(
        P2_U3191) );
  AND2_X1 U22792 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n19811), .ZN(
        P2_U3192) );
  NOR2_X1 U22793 ( .A1(n21063), .A2(n19885), .ZN(P2_U3193) );
  AND2_X1 U22794 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n19811), .ZN(
        P2_U3194) );
  AND2_X1 U22795 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n19811), .ZN(
        P2_U3195) );
  NOR2_X1 U22796 ( .A1(n20947), .A2(n19885), .ZN(P2_U3196) );
  AND2_X1 U22797 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n19811), .ZN(
        P2_U3197) );
  AND2_X1 U22798 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n19811), .ZN(
        P2_U3198) );
  AND2_X1 U22799 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n19811), .ZN(
        P2_U3199) );
  AND2_X1 U22800 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n19811), .ZN(
        P2_U3200) );
  INV_X1 U22801 ( .A(P2_DATAWIDTH_REG_9__SCAN_IN), .ZN(n21154) );
  NOR2_X1 U22802 ( .A1(n21154), .A2(n19885), .ZN(P2_U3201) );
  AND2_X1 U22803 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n19811), .ZN(P2_U3202) );
  AND2_X1 U22804 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n19811), .ZN(P2_U3203) );
  AND2_X1 U22805 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n19811), .ZN(P2_U3204) );
  AND2_X1 U22806 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n19811), .ZN(P2_U3205) );
  AND2_X1 U22807 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n19811), .ZN(P2_U3206) );
  AND2_X1 U22808 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n19811), .ZN(P2_U3207) );
  INV_X1 U22809 ( .A(P2_DATAWIDTH_REG_2__SCAN_IN), .ZN(n20931) );
  NOR2_X1 U22810 ( .A1(n20931), .A2(n19885), .ZN(P2_U3208) );
  INV_X1 U22811 ( .A(NA), .ZN(n20706) );
  OAI21_X1 U22812 ( .B1(n20706), .B2(n19819), .A(P2_STATE_REG_2__SCAN_IN), 
        .ZN(n19829) );
  INV_X1 U22813 ( .A(n19829), .ZN(n19816) );
  NAND2_X1 U22814 ( .A1(n19812), .A2(P2_STATE_REG_1__SCAN_IN), .ZN(n19827) );
  INV_X1 U22815 ( .A(n19827), .ZN(n19817) );
  NOR3_X1 U22816 ( .A1(n19817), .A2(n19813), .A3(n21058), .ZN(n19815) );
  OAI211_X1 U22817 ( .C1(HOLD), .C2(n19813), .A(n19937), .B(n19824), .ZN(
        n19814) );
  OAI21_X1 U22818 ( .B1(n19816), .B2(n19815), .A(n19814), .ZN(P2_U3209) );
  NOR2_X1 U22819 ( .A1(n19818), .A2(n19817), .ZN(n19821) );
  NOR2_X1 U22820 ( .A1(HOLD), .A2(n21058), .ZN(n19828) );
  OAI211_X1 U22821 ( .C1(n19828), .C2(n19830), .A(
        P2_REQUESTPENDING_REG_SCAN_IN), .B(n19819), .ZN(n19820) );
  OAI211_X1 U22822 ( .C1(n19823), .C2(n19822), .A(n19821), .B(n19820), .ZN(
        P2_U3210) );
  OAI22_X1 U22823 ( .A1(P2_REQUESTPENDING_REG_SCAN_IN), .A2(n19824), .B1(NA), 
        .B2(n19827), .ZN(n19825) );
  OAI211_X1 U22824 ( .C1(P2_REQUESTPENDING_REG_SCAN_IN), .C2(HOLD), .A(
        P2_STATE_REG_0__SCAN_IN), .B(n19825), .ZN(n19826) );
  OAI221_X1 U22825 ( .B1(n19829), .B2(n19828), .C1(n19829), .C2(n19827), .A(
        n19826), .ZN(P2_U3211) );
  OAI222_X1 U22826 ( .A1(n19875), .A2(n21092), .B1(n19832), .B2(n19940), .C1(
        n19831), .C2(n19873), .ZN(P2_U3212) );
  OAI222_X1 U22827 ( .A1(n19875), .A2(n11812), .B1(n19833), .B2(n19940), .C1(
        n21092), .C2(n19873), .ZN(P2_U3213) );
  OAI222_X1 U22828 ( .A1(n19875), .A2(n11816), .B1(n19834), .B2(n19940), .C1(
        n11812), .C2(n19873), .ZN(P2_U3214) );
  OAI222_X1 U22829 ( .A1(n19875), .A2(n19836), .B1(n19835), .B2(n19940), .C1(
        n11816), .C2(n19873), .ZN(P2_U3215) );
  OAI222_X1 U22830 ( .A1(n19875), .A2(n19838), .B1(n19837), .B2(n19940), .C1(
        n19836), .C2(n19873), .ZN(P2_U3216) );
  OAI222_X1 U22831 ( .A1(n19875), .A2(n11530), .B1(n19839), .B2(n19940), .C1(
        n19838), .C2(n19873), .ZN(P2_U3217) );
  OAI222_X1 U22832 ( .A1(n19875), .A2(n14190), .B1(n19840), .B2(n19940), .C1(
        n11530), .C2(n19873), .ZN(P2_U3218) );
  INV_X1 U22833 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n19842) );
  OAI222_X1 U22834 ( .A1(n19875), .A2(n19842), .B1(n19841), .B2(n19940), .C1(
        n14190), .C2(n19873), .ZN(P2_U3219) );
  OAI222_X1 U22835 ( .A1(n19875), .A2(n11864), .B1(n19843), .B2(n19940), .C1(
        n19842), .C2(n19873), .ZN(P2_U3220) );
  OAI222_X1 U22836 ( .A1(n19875), .A2(n11878), .B1(n19844), .B2(n19940), .C1(
        n11864), .C2(n19873), .ZN(P2_U3221) );
  OAI222_X1 U22837 ( .A1(n19875), .A2(n11892), .B1(n19845), .B2(n19940), .C1(
        n11878), .C2(n19873), .ZN(P2_U3222) );
  OAI222_X1 U22838 ( .A1(n19875), .A2(n15449), .B1(n19846), .B2(n19940), .C1(
        n11892), .C2(n19873), .ZN(P2_U3223) );
  OAI222_X1 U22839 ( .A1(n19875), .A2(n11919), .B1(n19847), .B2(n19940), .C1(
        n15449), .C2(n19873), .ZN(P2_U3224) );
  OAI222_X1 U22840 ( .A1(n19875), .A2(n15437), .B1(n19848), .B2(n19940), .C1(
        n11919), .C2(n19873), .ZN(P2_U3225) );
  INV_X1 U22841 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n19850) );
  OAI222_X1 U22842 ( .A1(n19875), .A2(n19850), .B1(n19849), .B2(n19940), .C1(
        n15437), .C2(n19873), .ZN(P2_U3226) );
  OAI222_X1 U22843 ( .A1(n19875), .A2(n21095), .B1(n19851), .B2(n19940), .C1(
        n19850), .C2(n19873), .ZN(P2_U3227) );
  OAI222_X1 U22844 ( .A1(n19875), .A2(n15411), .B1(n19852), .B2(n19940), .C1(
        n21095), .C2(n19873), .ZN(P2_U3228) );
  OAI222_X1 U22845 ( .A1(n19875), .A2(n19854), .B1(n19853), .B2(n19940), .C1(
        n15411), .C2(n19873), .ZN(P2_U3229) );
  OAI222_X1 U22846 ( .A1(n19875), .A2(n19856), .B1(n19855), .B2(n19940), .C1(
        n19854), .C2(n19873), .ZN(P2_U3230) );
  OAI222_X1 U22847 ( .A1(n19875), .A2(n21126), .B1(n19857), .B2(n19940), .C1(
        n19856), .C2(n19873), .ZN(P2_U3231) );
  OAI222_X1 U22848 ( .A1(n19875), .A2(n15861), .B1(n19858), .B2(n19940), .C1(
        n21126), .C2(n19873), .ZN(P2_U3232) );
  OAI222_X1 U22849 ( .A1(n19875), .A2(n19860), .B1(n19859), .B2(n19940), .C1(
        n15861), .C2(n19873), .ZN(P2_U3233) );
  OAI222_X1 U22850 ( .A1(n19875), .A2(n19862), .B1(n19861), .B2(n19940), .C1(
        n19860), .C2(n19873), .ZN(P2_U3234) );
  OAI222_X1 U22851 ( .A1(n19875), .A2(n19864), .B1(n19863), .B2(n19940), .C1(
        n19862), .C2(n19873), .ZN(P2_U3235) );
  OAI222_X1 U22852 ( .A1(n19875), .A2(n19866), .B1(n19865), .B2(n19940), .C1(
        n19864), .C2(n19873), .ZN(P2_U3236) );
  OAI222_X1 U22853 ( .A1(n19875), .A2(n21193), .B1(n19867), .B2(n19940), .C1(
        n19866), .C2(n19873), .ZN(P2_U3237) );
  OAI222_X1 U22854 ( .A1(n19873), .A2(n21193), .B1(n19868), .B2(n19940), .C1(
        n19869), .C2(n19875), .ZN(P2_U3238) );
  OAI222_X1 U22855 ( .A1(n19875), .A2(n19871), .B1(n19870), .B2(n19940), .C1(
        n19869), .C2(n19873), .ZN(P2_U3239) );
  OAI222_X1 U22856 ( .A1(n19875), .A2(n12509), .B1(n19872), .B2(n19940), .C1(
        n19871), .C2(n19873), .ZN(P2_U3240) );
  OAI222_X1 U22857 ( .A1(n19875), .A2(n19874), .B1(n21093), .B2(n19940), .C1(
        n12509), .C2(n19873), .ZN(P2_U3241) );
  AOI22_X1 U22858 ( .A1(n19940), .A2(n21195), .B1(n20943), .B2(n19937), .ZN(
        P2_U3585) );
  INV_X1 U22859 ( .A(P2_BE_N_REG_2__SCAN_IN), .ZN(n19876) );
  AOI22_X1 U22860 ( .A1(n19940), .A2(n19877), .B1(n19876), .B2(n19937), .ZN(
        P2_U3586) );
  INV_X1 U22861 ( .A(P2_BE_N_REG_1__SCAN_IN), .ZN(n19878) );
  AOI22_X1 U22862 ( .A1(n19940), .A2(n19879), .B1(n19878), .B2(n19937), .ZN(
        P2_U3587) );
  INV_X1 U22863 ( .A(P2_BE_N_REG_0__SCAN_IN), .ZN(n19880) );
  AOI22_X1 U22864 ( .A1(n19940), .A2(n19881), .B1(n19880), .B2(n19937), .ZN(
        P2_U3588) );
  OAI21_X1 U22865 ( .B1(n19885), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .A(n19883), 
        .ZN(n19882) );
  INV_X1 U22866 ( .A(n19882), .ZN(P2_U3591) );
  INV_X1 U22867 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n19884) );
  OAI21_X1 U22868 ( .B1(n19885), .B2(n19884), .A(n19883), .ZN(P2_U3592) );
  OR2_X1 U22869 ( .A1(n19887), .A2(n19886), .ZN(n19896) );
  INV_X1 U22870 ( .A(n19907), .ZN(n19888) );
  OR2_X1 U22871 ( .A1(n19889), .A2(n19888), .ZN(n19899) );
  NAND2_X1 U22872 ( .A1(n19890), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19891) );
  OAI21_X1 U22873 ( .B1(n19910), .B2(n19891), .A(n19920), .ZN(n19900) );
  NAND2_X1 U22874 ( .A1(n19899), .A2(n19900), .ZN(n19893) );
  AOI22_X1 U22875 ( .A1(n19894), .A2(n19893), .B1(P2_STATE2_REG_3__SCAN_IN), 
        .B2(n19892), .ZN(n19895) );
  AND2_X1 U22876 ( .A1(n19896), .A2(n19895), .ZN(n19897) );
  AOI22_X1 U22877 ( .A1(n19925), .A2(n19898), .B1(n19897), .B2(n19922), .ZN(
        P2_U3602) );
  OAI21_X1 U22878 ( .B1(n19901), .B2(n19900), .A(n19899), .ZN(n19902) );
  AOI21_X1 U22879 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19903), .A(n19902), 
        .ZN(n19904) );
  AOI22_X1 U22880 ( .A1(n19925), .A2(n19905), .B1(n19904), .B2(n19922), .ZN(
        P2_U3603) );
  AOI22_X1 U22881 ( .A1(n19910), .A2(n19907), .B1(P2_STATE2_REG_3__SCAN_IN), 
        .B2(n19906), .ZN(n19913) );
  INV_X1 U22882 ( .A(n19920), .ZN(n19909) );
  AND2_X1 U22883 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19908) );
  NOR3_X1 U22884 ( .A1(n19910), .A2(n19909), .A3(n19908), .ZN(n19911) );
  NOR2_X1 U22885 ( .A1(n19925), .A2(n19911), .ZN(n19912) );
  AOI22_X1 U22886 ( .A1(n19914), .A2(n19925), .B1(n19913), .B2(n19912), .ZN(
        P2_U3604) );
  NOR2_X1 U22887 ( .A1(n19916), .A2(n19915), .ZN(n19919) );
  NOR2_X1 U22888 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19917), .ZN(
        n19918) );
  AOI211_X1 U22889 ( .C1(n19921), .C2(n19920), .A(n19919), .B(n19918), .ZN(
        n19923) );
  AOI22_X1 U22890 ( .A1(n19925), .A2(n19924), .B1(n19923), .B2(n19922), .ZN(
        P2_U3605) );
  AOI22_X1 U22891 ( .A1(n19940), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n19926), 
        .B2(n19937), .ZN(P2_U3608) );
  INV_X1 U22892 ( .A(P2_MORE_REG_SCAN_IN), .ZN(n21138) );
  INV_X1 U22893 ( .A(n19933), .ZN(n19936) );
  INV_X1 U22894 ( .A(n19927), .ZN(n19931) );
  AOI22_X1 U22895 ( .A1(n19931), .A2(n19930), .B1(n19929), .B2(n19928), .ZN(
        n19935) );
  AND2_X1 U22896 ( .A1(n19933), .A2(n19932), .ZN(n19934) );
  AOI22_X1 U22897 ( .A1(n21138), .A2(n19936), .B1(n19935), .B2(n19934), .ZN(
        P2_U3609) );
  INV_X1 U22898 ( .A(P2_M_IO_N_REG_SCAN_IN), .ZN(n19938) );
  AOI22_X1 U22899 ( .A1(n19940), .A2(n19939), .B1(n19938), .B2(n19937), .ZN(
        P2_U3611) );
  AND2_X1 U22900 ( .A1(n20700), .A2(P1_STATE_REG_0__SCAN_IN), .ZN(n19942) );
  INV_X1 U22901 ( .A(P1_ADS_N_REG_SCAN_IN), .ZN(n19941) );
  INV_X1 U22902 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n20704) );
  AOI21_X1 U22903 ( .B1(n19942), .B2(n19941), .A(n20814), .ZN(P1_U2802) );
  OAI21_X1 U22904 ( .B1(n19944), .B2(n19943), .A(P1_CODEFETCH_REG_SCAN_IN), 
        .ZN(n19945) );
  OAI21_X1 U22905 ( .B1(n19946), .B2(n20806), .A(n19945), .ZN(P1_U2803) );
  NOR2_X1 U22906 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(P1_STATE_REG_0__SCAN_IN), 
        .ZN(n19948) );
  OAI21_X1 U22907 ( .B1(n19948), .B2(P1_D_C_N_REG_SCAN_IN), .A(n9834), .ZN(
        n19947) );
  OAI21_X1 U22908 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(n9834), .A(n19947), 
        .ZN(P1_U2804) );
  AOI21_X1 U22909 ( .B1(P1_STATE_REG_0__SCAN_IN), .B2(n20700), .A(n20814), 
        .ZN(n20770) );
  OAI21_X1 U22910 ( .B1(BS16), .B2(n19948), .A(n20770), .ZN(n20768) );
  OAI21_X1 U22911 ( .B1(n20770), .B2(n20208), .A(n20768), .ZN(P1_U2805) );
  OAI21_X1 U22912 ( .B1(n19951), .B2(n19950), .A(n19949), .ZN(P1_U2806) );
  NOR4_X1 U22913 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_20__SCAN_IN), .A3(P1_DATAWIDTH_REG_21__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_22__SCAN_IN), .ZN(n19955) );
  NOR4_X1 U22914 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_16__SCAN_IN), .A3(P1_DATAWIDTH_REG_17__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_18__SCAN_IN), .ZN(n19954) );
  NOR4_X1 U22915 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_29__SCAN_IN), .A3(P1_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_31__SCAN_IN), .ZN(n19953) );
  NOR4_X1 U22916 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_24__SCAN_IN), .A3(P1_DATAWIDTH_REG_25__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_26__SCAN_IN), .ZN(n19952) );
  NAND4_X1 U22917 ( .A1(n19955), .A2(n19954), .A3(n19953), .A4(n19952), .ZN(
        n19961) );
  NOR4_X1 U22918 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_27__SCAN_IN), .A3(P1_DATAWIDTH_REG_2__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_3__SCAN_IN), .ZN(n19959) );
  AOI211_X1 U22919 ( .C1(P1_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_7__SCAN_IN), .B(
        P1_DATAWIDTH_REG_5__SCAN_IN), .ZN(n19958) );
  NOR4_X1 U22920 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_12__SCAN_IN), .A3(P1_DATAWIDTH_REG_13__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_14__SCAN_IN), .ZN(n19957) );
  NOR4_X1 U22921 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_6__SCAN_IN), .A3(P1_DATAWIDTH_REG_8__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_9__SCAN_IN), .ZN(n19956) );
  NAND4_X1 U22922 ( .A1(n19959), .A2(n19958), .A3(n19957), .A4(n19956), .ZN(
        n19960) );
  NOR2_X1 U22923 ( .A1(n19961), .A2(n19960), .ZN(n20798) );
  INV_X1 U22924 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n20763) );
  NOR3_X1 U22925 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A3(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n19963) );
  OAI21_X1 U22926 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n19963), .A(n20798), .ZN(
        n19962) );
  OAI21_X1 U22927 ( .B1(n20798), .B2(n20763), .A(n19962), .ZN(P1_U2807) );
  INV_X1 U22928 ( .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20769) );
  AOI21_X1 U22929 ( .B1(n13701), .B2(n20769), .A(n19963), .ZN(n19964) );
  INV_X1 U22930 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n20760) );
  INV_X1 U22931 ( .A(n20798), .ZN(n20795) );
  AOI22_X1 U22932 ( .A1(n20798), .A2(n19964), .B1(n20760), .B2(n20795), .ZN(
        P1_U2808) );
  AOI22_X1 U22933 ( .A1(P1_EBX_REG_9__SCAN_IN), .A2(n20025), .B1(n20010), .B2(
        n19965), .ZN(n19966) );
  OAI211_X1 U22934 ( .C1(n20014), .C2(n19967), .A(n19966), .B(n20011), .ZN(
        n19968) );
  AOI221_X1 U22935 ( .B1(n19970), .B2(n21039), .C1(n19969), .C2(
        P1_REIP_REG_9__SCAN_IN), .A(n19968), .ZN(n19973) );
  AOI22_X1 U22936 ( .A1(n20041), .A2(n19992), .B1(n20034), .B2(n19971), .ZN(
        n19972) );
  NAND2_X1 U22937 ( .A1(n19973), .A2(n19972), .ZN(P1_U2831) );
  NAND2_X1 U22938 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(P1_REIP_REG_5__SCAN_IN), 
        .ZN(n19978) );
  NOR3_X1 U22939 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(n19978), .A3(n19999), .ZN(
        n19977) );
  AOI22_X1 U22940 ( .A1(P1_EBX_REG_7__SCAN_IN), .A2(n20025), .B1(n20010), .B2(
        n19974), .ZN(n19975) );
  OAI211_X1 U22941 ( .C1(n20014), .C2(n10662), .A(n19975), .B(n20011), .ZN(
        n19976) );
  NOR2_X1 U22942 ( .A1(n19977), .A2(n19976), .ZN(n19984) );
  INV_X1 U22943 ( .A(n19978), .ZN(n19981) );
  INV_X1 U22944 ( .A(n20023), .ZN(n20028) );
  AOI21_X1 U22945 ( .B1(n20028), .B2(n19980), .A(n19979), .ZN(n20021) );
  OAI21_X1 U22946 ( .B1(n19981), .B2(n20023), .A(n20021), .ZN(n19991) );
  AOI22_X1 U22947 ( .A1(n19982), .A2(n19992), .B1(n19991), .B2(
        P1_REIP_REG_7__SCAN_IN), .ZN(n19983) );
  OAI211_X1 U22948 ( .C1(n19985), .C2(n20006), .A(n19984), .B(n19983), .ZN(
        P1_U2833) );
  NOR2_X1 U22949 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(n19999), .ZN(n19986) );
  AOI22_X1 U22950 ( .A1(P1_EBX_REG_6__SCAN_IN), .A2(n20025), .B1(
        P1_REIP_REG_5__SCAN_IN), .B2(n19986), .ZN(n19987) );
  OAI21_X1 U22951 ( .B1(n20038), .B2(n19988), .A(n19987), .ZN(n19989) );
  AOI211_X1 U22952 ( .C1(n20026), .C2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n19990), .B(n19989), .ZN(n19995) );
  AOI22_X1 U22953 ( .A1(n19993), .A2(n19992), .B1(n19991), .B2(
        P1_REIP_REG_6__SCAN_IN), .ZN(n19994) );
  OAI211_X1 U22954 ( .C1(n19996), .C2(n20006), .A(n19995), .B(n19994), .ZN(
        P1_U2834) );
  OAI22_X1 U22955 ( .A1(n19999), .A2(P1_REIP_REG_5__SCAN_IN), .B1(n19998), 
        .B2(n19997), .ZN(n20003) );
  AOI22_X1 U22956 ( .A1(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n20026), .B1(
        n20010), .B2(n20000), .ZN(n20001) );
  OAI211_X1 U22957 ( .C1(n20021), .C2(n16192), .A(n20001), .B(n20011), .ZN(
        n20002) );
  AOI211_X1 U22958 ( .C1(n20004), .C2(n20017), .A(n20003), .B(n20002), .ZN(
        n20005) );
  OAI21_X1 U22959 ( .B1(n20007), .B2(n20006), .A(n20005), .ZN(P1_U2835) );
  NOR3_X1 U22960 ( .A1(n13701), .A2(n13935), .A3(n13774), .ZN(n20008) );
  AOI21_X1 U22961 ( .B1(n20028), .B2(n20008), .A(P1_REIP_REG_4__SCAN_IN), .ZN(
        n20020) );
  AOI22_X1 U22962 ( .A1(n20010), .A2(n20104), .B1(n20009), .B2(n20027), .ZN(
        n20012) );
  OAI211_X1 U22963 ( .C1(n20014), .C2(n20013), .A(n20012), .B(n20011), .ZN(
        n20015) );
  AOI21_X1 U22964 ( .B1(P1_EBX_REG_4__SCAN_IN), .B2(n20025), .A(n20015), .ZN(
        n20019) );
  INV_X1 U22965 ( .A(n20101), .ZN(n20016) );
  AOI22_X1 U22966 ( .A1(n20096), .A2(n20017), .B1(n20034), .B2(n20016), .ZN(
        n20018) );
  OAI211_X1 U22967 ( .C1(n20021), .C2(n20020), .A(n20019), .B(n20018), .ZN(
        P1_U2836) );
  OAI21_X1 U22968 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n20023), .A(n20022), .ZN(
        n20024) );
  AOI22_X1 U22969 ( .A1(P1_EBX_REG_2__SCAN_IN), .A2(n20025), .B1(
        P1_REIP_REG_2__SCAN_IN), .B2(n20024), .ZN(n20037) );
  INV_X1 U22970 ( .A(n13707), .ZN(n20154) );
  AOI22_X1 U22971 ( .A1(n20154), .A2(n20027), .B1(n20026), .B2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n20030) );
  NAND3_X1 U22972 ( .A1(n20028), .A2(n13774), .A3(P1_REIP_REG_1__SCAN_IN), 
        .ZN(n20029) );
  OAI211_X1 U22973 ( .C1(n20032), .C2(n20031), .A(n20030), .B(n20029), .ZN(
        n20033) );
  AOI21_X1 U22974 ( .B1(n20035), .B2(n20034), .A(n20033), .ZN(n20036) );
  OAI211_X1 U22975 ( .C1(n20038), .C2(n20129), .A(n20037), .B(n20036), .ZN(
        P1_U2838) );
  INV_X1 U22976 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n21047) );
  AOI22_X1 U22977 ( .A1(n20041), .A2(n20040), .B1(n20039), .B2(n20076), .ZN(
        n20042) );
  OAI21_X1 U22978 ( .B1(n20043), .B2(n21047), .A(n20042), .ZN(P1_U2895) );
  AOI22_X1 U22979 ( .A1(P1_EAX_REG_15__SCAN_IN), .A2(n20047), .B1(n20064), 
        .B2(P1_DATAO_REG_15__SCAN_IN), .ZN(n20044) );
  OAI21_X1 U22980 ( .B1(n20046), .B2(n20045), .A(n20044), .ZN(P1_U2921) );
  AOI22_X1 U22981 ( .A1(P1_LWORD_REG_14__SCAN_IN), .A2(n20811), .B1(n20064), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n20048) );
  OAI21_X1 U22982 ( .B1(n14373), .B2(n20073), .A(n20048), .ZN(P1_U2922) );
  AOI22_X1 U22983 ( .A1(P1_LWORD_REG_13__SCAN_IN), .A2(n20811), .B1(n20064), 
        .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n20049) );
  OAI21_X1 U22984 ( .B1(n20971), .B2(n20073), .A(n20049), .ZN(P1_U2923) );
  INV_X1 U22985 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n20051) );
  AOI22_X1 U22986 ( .A1(P1_LWORD_REG_12__SCAN_IN), .A2(n20811), .B1(n20064), 
        .B2(P1_DATAO_REG_12__SCAN_IN), .ZN(n20050) );
  OAI21_X1 U22987 ( .B1(n20051), .B2(n20073), .A(n20050), .ZN(P1_U2924) );
  AOI22_X1 U22988 ( .A1(P1_LWORD_REG_11__SCAN_IN), .A2(n20811), .B1(n20071), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n20052) );
  OAI21_X1 U22989 ( .B1(n20053), .B2(n20073), .A(n20052), .ZN(P1_U2925) );
  AOI22_X1 U22990 ( .A1(P1_LWORD_REG_10__SCAN_IN), .A2(n20811), .B1(n20064), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n20054) );
  OAI21_X1 U22991 ( .B1(n21136), .B2(n20073), .A(n20054), .ZN(P1_U2926) );
  AOI22_X1 U22992 ( .A1(P1_LWORD_REG_9__SCAN_IN), .A2(n20811), .B1(n20064), 
        .B2(P1_DATAO_REG_9__SCAN_IN), .ZN(n20055) );
  OAI21_X1 U22993 ( .B1(n21047), .B2(n20073), .A(n20055), .ZN(P1_U2927) );
  AOI22_X1 U22994 ( .A1(P1_LWORD_REG_8__SCAN_IN), .A2(n20811), .B1(n20064), 
        .B2(P1_DATAO_REG_8__SCAN_IN), .ZN(n20056) );
  OAI21_X1 U22995 ( .B1(n20057), .B2(n20073), .A(n20056), .ZN(P1_U2928) );
  AOI22_X1 U22996 ( .A1(P1_LWORD_REG_7__SCAN_IN), .A2(n20811), .B1(n20064), 
        .B2(P1_DATAO_REG_7__SCAN_IN), .ZN(n20058) );
  OAI21_X1 U22997 ( .B1(n20059), .B2(n20073), .A(n20058), .ZN(P1_U2929) );
  AOI22_X1 U22998 ( .A1(P1_LWORD_REG_6__SCAN_IN), .A2(n20811), .B1(n20064), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n20060) );
  OAI21_X1 U22999 ( .B1(n14014), .B2(n20073), .A(n20060), .ZN(P1_U2930) );
  AOI22_X1 U23000 ( .A1(P1_LWORD_REG_5__SCAN_IN), .A2(n20811), .B1(n20064), 
        .B2(P1_DATAO_REG_5__SCAN_IN), .ZN(n20061) );
  OAI21_X1 U23001 ( .B1(n10638), .B2(n20073), .A(n20061), .ZN(P1_U2931) );
  AOI22_X1 U23002 ( .A1(P1_LWORD_REG_4__SCAN_IN), .A2(n20811), .B1(n20064), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .ZN(n20062) );
  OAI21_X1 U23003 ( .B1(n20063), .B2(n20073), .A(n20062), .ZN(P1_U2932) );
  AOI22_X1 U23004 ( .A1(P1_LWORD_REG_3__SCAN_IN), .A2(n20811), .B1(n20064), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n20065) );
  OAI21_X1 U23005 ( .B1(n20066), .B2(n20073), .A(n20065), .ZN(P1_U2933) );
  AOI22_X1 U23006 ( .A1(P1_LWORD_REG_2__SCAN_IN), .A2(n20811), .B1(n20071), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n20067) );
  OAI21_X1 U23007 ( .B1(n20068), .B2(n20073), .A(n20067), .ZN(P1_U2934) );
  AOI22_X1 U23008 ( .A1(P1_LWORD_REG_1__SCAN_IN), .A2(n20811), .B1(n20071), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n20069) );
  OAI21_X1 U23009 ( .B1(n20070), .B2(n20073), .A(n20069), .ZN(P1_U2935) );
  AOI22_X1 U23010 ( .A1(P1_LWORD_REG_0__SCAN_IN), .A2(n20811), .B1(n20071), 
        .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n20072) );
  OAI21_X1 U23011 ( .B1(n20074), .B2(n20073), .A(n20072), .ZN(P1_U2936) );
  AOI22_X1 U23012 ( .A1(n20088), .A2(P1_EAX_REG_25__SCAN_IN), .B1(
        P1_UWORD_REG_9__SCAN_IN), .B2(n20075), .ZN(n20077) );
  NAND2_X1 U23013 ( .A1(n20082), .A2(n20076), .ZN(n20084) );
  NAND2_X1 U23014 ( .A1(n20077), .A2(n20084), .ZN(P1_U2946) );
  AOI22_X1 U23015 ( .A1(n20088), .A2(P1_EAX_REG_28__SCAN_IN), .B1(
        P1_UWORD_REG_12__SCAN_IN), .B2(n13688), .ZN(n20079) );
  NAND2_X1 U23016 ( .A1(n20082), .A2(n20078), .ZN(n20086) );
  NAND2_X1 U23017 ( .A1(n20079), .A2(n20086), .ZN(P1_U2949) );
  AOI22_X1 U23018 ( .A1(n20088), .A2(P1_EAX_REG_30__SCAN_IN), .B1(
        P1_UWORD_REG_14__SCAN_IN), .B2(n13688), .ZN(n20083) );
  INV_X1 U23019 ( .A(n20080), .ZN(n20081) );
  NAND2_X1 U23020 ( .A1(n20082), .A2(n20081), .ZN(n20089) );
  NAND2_X1 U23021 ( .A1(n20083), .A2(n20089), .ZN(P1_U2951) );
  AOI22_X1 U23022 ( .A1(n20088), .A2(P1_EAX_REG_9__SCAN_IN), .B1(
        P1_LWORD_REG_9__SCAN_IN), .B2(n20075), .ZN(n20085) );
  NAND2_X1 U23023 ( .A1(n20085), .A2(n20084), .ZN(P1_U2961) );
  AOI22_X1 U23024 ( .A1(n20088), .A2(P1_EAX_REG_12__SCAN_IN), .B1(
        P1_LWORD_REG_12__SCAN_IN), .B2(n20075), .ZN(n20087) );
  NAND2_X1 U23025 ( .A1(n20087), .A2(n20086), .ZN(P1_U2964) );
  AOI22_X1 U23026 ( .A1(n20088), .A2(P1_EAX_REG_14__SCAN_IN), .B1(
        P1_LWORD_REG_14__SCAN_IN), .B2(n20075), .ZN(n20090) );
  NAND2_X1 U23027 ( .A1(n20090), .A2(n20089), .ZN(P1_U2966) );
  AOI22_X1 U23028 ( .A1(n20091), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .B1(
        n20103), .B2(P1_REIP_REG_4__SCAN_IN), .ZN(n20100) );
  OAI21_X1 U23029 ( .B1(n20094), .B2(n20093), .A(n20092), .ZN(n20095) );
  INV_X1 U23030 ( .A(n20095), .ZN(n20105) );
  AOI22_X1 U23031 ( .A1(n20105), .A2(n20098), .B1(n20097), .B2(n20096), .ZN(
        n20099) );
  OAI211_X1 U23032 ( .C1(n20102), .C2(n20101), .A(n20100), .B(n20099), .ZN(
        P1_U2995) );
  AOI22_X1 U23033 ( .A1(n20114), .A2(n20104), .B1(n20103), .B2(
        P1_REIP_REG_4__SCAN_IN), .ZN(n20110) );
  AOI22_X1 U23034 ( .A1(n20105), .A2(n20137), .B1(
        P1_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n20116), .ZN(n20109) );
  OAI211_X1 U23035 ( .C1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A(n20107), .B(n20106), .ZN(n20108) );
  NAND3_X1 U23036 ( .A1(n20110), .A2(n20109), .A3(n20108), .ZN(P1_U3027) );
  INV_X1 U23037 ( .A(n20111), .ZN(n20113) );
  AOI21_X1 U23038 ( .B1(n20114), .B2(n20113), .A(n20112), .ZN(n20118) );
  AOI22_X1 U23039 ( .A1(n20116), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .B1(
        n20115), .B2(n20137), .ZN(n20117) );
  OAI211_X1 U23040 ( .C1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .C2(n20119), .A(
        n20118), .B(n20117), .ZN(P1_U3028) );
  OR2_X1 U23041 ( .A1(n20151), .A2(n20120), .ZN(n20136) );
  NOR3_X1 U23042 ( .A1(n20122), .A2(n20151), .A3(n20121), .ZN(n20124) );
  AOI211_X1 U23043 ( .C1(n20151), .C2(n20125), .A(n20124), .B(n20123), .ZN(
        n20134) );
  AND3_X1 U23044 ( .A1(n20127), .A2(n20126), .A3(n20137), .ZN(n20132) );
  OAI22_X1 U23045 ( .A1(n20145), .A2(n20129), .B1(n13774), .B2(n20128), .ZN(
        n20130) );
  NOR3_X1 U23046 ( .A1(n20132), .A2(n20131), .A3(n20130), .ZN(n20133) );
  OAI221_X1 U23047 ( .B1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n20136), .C1(
        n20135), .C2(n20134), .A(n20133), .ZN(P1_U3029) );
  AND3_X1 U23048 ( .A1(n13704), .A2(n20138), .A3(n20137), .ZN(n20147) );
  NAND3_X1 U23049 ( .A1(n20151), .A2(n20140), .A3(n20139), .ZN(n20143) );
  INV_X1 U23050 ( .A(n20141), .ZN(n20142) );
  OAI211_X1 U23051 ( .C1(n20145), .C2(n20144), .A(n20143), .B(n20142), .ZN(
        n20146) );
  NOR2_X1 U23052 ( .A1(n20147), .A2(n20146), .ZN(n20148) );
  OAI221_X1 U23053 ( .B1(n20151), .B2(n20150), .C1(n20151), .C2(n20149), .A(
        n20148), .ZN(P1_U3030) );
  NOR2_X1 U23054 ( .A1(n20152), .A2(n20791), .ZN(P1_U3032) );
  NAND2_X1 U23055 ( .A1(n20465), .A2(n20406), .ZN(n20293) );
  NAND2_X1 U23056 ( .A1(n20163), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20593) );
  NAND2_X1 U23057 ( .A1(n20297), .A2(n20593), .ZN(n20232) );
  OR2_X1 U23058 ( .A1(n13917), .A2(n20294), .ZN(n20569) );
  NAND2_X1 U23059 ( .A1(n20637), .A2(n20562), .ZN(n20681) );
  OAI21_X1 U23060 ( .B1(n20221), .B2(n20688), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20153) );
  INV_X1 U23061 ( .A(n20786), .ZN(n20500) );
  NAND2_X1 U23062 ( .A1(n20153), .A2(n20500), .ZN(n20165) );
  OR2_X1 U23063 ( .A1(n20234), .A2(n20591), .ZN(n20164) );
  INV_X1 U23064 ( .A(n20164), .ZN(n20155) );
  NAND3_X1 U23065 ( .A1(n20783), .A2(n20461), .A3(n20523), .ZN(n20207) );
  NOR2_X1 U23066 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20207), .ZN(
        n20197) );
  OAI22_X1 U23067 ( .A1(n20165), .A2(n20155), .B1(n20197), .B2(n20413), .ZN(
        n20156) );
  INV_X1 U23068 ( .A(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n21074) );
  NOR2_X2 U23069 ( .A1(n20195), .A2(n20157), .ZN(n20636) );
  NOR2_X2 U23070 ( .A1(n20159), .A2(n20158), .ZN(n20196) );
  AOI22_X1 U23071 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n20196), .B1(DATAI_24_), 
        .B2(n20161), .ZN(n20539) );
  INV_X1 U23072 ( .A(n20539), .ZN(n20641) );
  AOI22_X1 U23073 ( .A1(n20636), .A2(n20197), .B1(n20688), .B2(n20641), .ZN(
        n20167) );
  NOR2_X2 U23074 ( .A1(n20162), .A2(n20198), .ZN(n20635) );
  OR2_X1 U23075 ( .A1(n20163), .A2(n20802), .ZN(n20469) );
  AOI22_X1 U23076 ( .A1(DATAI_16_), .A2(n20161), .B1(BUF1_REG_16__SCAN_IN), 
        .B2(n20196), .ZN(n20644) );
  INV_X1 U23077 ( .A(n20644), .ZN(n20524) );
  AOI22_X1 U23078 ( .A1(n20635), .A2(n20200), .B1(n20221), .B2(n20524), .ZN(
        n20166) );
  OAI211_X1 U23079 ( .C1(n20183), .C2(n21074), .A(n20167), .B(n20166), .ZN(
        P1_U3033) );
  NOR2_X2 U23080 ( .A1(n20195), .A2(n20168), .ZN(n20646) );
  AOI22_X1 U23081 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n20196), .B1(DATAI_25_), 
        .B2(n20161), .ZN(n20650) );
  INV_X1 U23082 ( .A(n20650), .ZN(n20602) );
  AOI22_X1 U23083 ( .A1(n20646), .A2(n20197), .B1(n20688), .B2(n20602), .ZN(
        n20171) );
  NOR2_X2 U23084 ( .A1(n20169), .A2(n20198), .ZN(n20645) );
  AOI22_X1 U23085 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n20196), .B1(DATAI_17_), 
        .B2(n20161), .ZN(n20605) );
  INV_X1 U23086 ( .A(n20605), .ZN(n20647) );
  AOI22_X1 U23087 ( .A1(n20645), .A2(n20200), .B1(n20221), .B2(n20647), .ZN(
        n20170) );
  OAI211_X1 U23088 ( .C1(n20183), .C2(n20172), .A(n20171), .B(n20170), .ZN(
        P1_U3034) );
  INV_X1 U23089 ( .A(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n20176) );
  NOR2_X2 U23090 ( .A1(n20195), .A2(n13376), .ZN(n20652) );
  AOI22_X1 U23091 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n20196), .B1(DATAI_26_), 
        .B2(n20161), .ZN(n20545) );
  INV_X1 U23092 ( .A(n20545), .ZN(n20653) );
  AOI22_X1 U23093 ( .A1(n20652), .A2(n20197), .B1(n20688), .B2(n20653), .ZN(
        n20175) );
  NOR2_X2 U23094 ( .A1(n20173), .A2(n20198), .ZN(n20651) );
  AOI22_X1 U23095 ( .A1(DATAI_18_), .A2(n20161), .B1(BUF1_REG_18__SCAN_IN), 
        .B2(n20196), .ZN(n20656) );
  INV_X1 U23096 ( .A(n20656), .ZN(n20542) );
  AOI22_X1 U23097 ( .A1(n20651), .A2(n20200), .B1(n20221), .B2(n20542), .ZN(
        n20174) );
  OAI211_X1 U23098 ( .C1(n20183), .C2(n20176), .A(n20175), .B(n20174), .ZN(
        P1_U3035) );
  INV_X1 U23099 ( .A(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n20181) );
  NOR2_X2 U23100 ( .A1(n20195), .A2(n20177), .ZN(n20658) );
  AOI22_X1 U23101 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n20196), .B1(DATAI_27_), 
        .B2(n20161), .ZN(n20662) );
  INV_X1 U23102 ( .A(n20662), .ZN(n20608) );
  AOI22_X1 U23103 ( .A1(n20658), .A2(n20197), .B1(n20688), .B2(n20608), .ZN(
        n20180) );
  NOR2_X2 U23104 ( .A1(n20178), .A2(n20198), .ZN(n20657) );
  AOI22_X1 U23105 ( .A1(DATAI_19_), .A2(n20161), .B1(BUF1_REG_19__SCAN_IN), 
        .B2(n20196), .ZN(n20611) );
  INV_X1 U23106 ( .A(n20611), .ZN(n20659) );
  AOI22_X1 U23107 ( .A1(n20657), .A2(n20200), .B1(n20221), .B2(n20659), .ZN(
        n20179) );
  OAI211_X1 U23108 ( .C1(n20183), .C2(n20181), .A(n20180), .B(n20179), .ZN(
        P1_U3036) );
  AOI22_X1 U23109 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n20196), .B1(DATAI_20_), 
        .B2(n20161), .ZN(n20615) );
  NOR2_X2 U23110 ( .A1(n20195), .A2(n20182), .ZN(n20664) );
  AOI22_X1 U23111 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n20196), .B1(DATAI_28_), 
        .B2(n20161), .ZN(n20668) );
  INV_X1 U23112 ( .A(n20668), .ZN(n20612) );
  AOI22_X1 U23113 ( .A1(n20664), .A2(n20197), .B1(n20688), .B2(n20612), .ZN(
        n20186) );
  INV_X1 U23114 ( .A(n20183), .ZN(n20201) );
  NOR2_X2 U23115 ( .A1(n20184), .A2(n20198), .ZN(n20663) );
  AOI22_X1 U23116 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n20201), .B1(
        n20663), .B2(n20200), .ZN(n20185) );
  OAI211_X1 U23117 ( .C1(n20615), .C2(n20231), .A(n20186), .B(n20185), .ZN(
        P1_U3037) );
  AOI22_X1 U23118 ( .A1(DATAI_21_), .A2(n20161), .B1(BUF1_REG_21__SCAN_IN), 
        .B2(n20196), .ZN(n20619) );
  AOI22_X1 U23119 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n20196), .B1(DATAI_29_), 
        .B2(n20161), .ZN(n20674) );
  INV_X1 U23120 ( .A(n20674), .ZN(n20616) );
  AOI22_X1 U23121 ( .A1(n9828), .A2(n20197), .B1(n20688), .B2(n20616), .ZN(
        n20189) );
  NOR2_X2 U23122 ( .A1(n20187), .A2(n20198), .ZN(n20669) );
  AOI22_X1 U23123 ( .A1(P1_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n20201), .B1(
        n20669), .B2(n20200), .ZN(n20188) );
  OAI211_X1 U23124 ( .C1(n20619), .C2(n20231), .A(n20189), .B(n20188), .ZN(
        P1_U3038) );
  NOR2_X2 U23125 ( .A1(n20195), .A2(n20190), .ZN(n20676) );
  AOI22_X1 U23126 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n20196), .B1(DATAI_30_), 
        .B2(n20161), .ZN(n20555) );
  INV_X1 U23127 ( .A(n20555), .ZN(n20677) );
  AOI22_X1 U23128 ( .A1(n20676), .A2(n20197), .B1(n20688), .B2(n20677), .ZN(
        n20193) );
  NOR2_X2 U23129 ( .A1(n20191), .A2(n20198), .ZN(n20675) );
  AOI22_X1 U23130 ( .A1(P1_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n20201), .B1(
        n20675), .B2(n20200), .ZN(n20192) );
  OAI211_X1 U23131 ( .C1(n20682), .C2(n20231), .A(n20193), .B(n20192), .ZN(
        P1_U3039) );
  AOI22_X1 U23132 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n20196), .B1(DATAI_23_), 
        .B2(n20161), .ZN(n20629) );
  NOR2_X2 U23133 ( .A1(n20195), .A2(n20194), .ZN(n20686) );
  AOI22_X1 U23134 ( .A1(BUF1_REG_31__SCAN_IN), .A2(n20196), .B1(DATAI_31_), 
        .B2(n20161), .ZN(n20693) );
  INV_X1 U23135 ( .A(n20693), .ZN(n20624) );
  AOI22_X1 U23136 ( .A1(n20686), .A2(n20197), .B1(n20688), .B2(n20624), .ZN(
        n20203) );
  NOR2_X2 U23137 ( .A1(n20199), .A2(n20198), .ZN(n20684) );
  AOI22_X1 U23138 ( .A1(P1_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n20201), .B1(
        n20684), .B2(n20200), .ZN(n20202) );
  OAI211_X1 U23139 ( .C1(n20629), .C2(n20231), .A(n20203), .B(n20202), .ZN(
        P1_U3040) );
  NOR2_X1 U23140 ( .A1(n20790), .A2(n20207), .ZN(n20227) );
  INV_X1 U23141 ( .A(n20205), .ZN(n20434) );
  NAND2_X1 U23142 ( .A1(n20434), .A2(n20500), .ZN(n20565) );
  INV_X1 U23143 ( .A(n20227), .ZN(n20206) );
  OAI222_X1 U23144 ( .A1(n20234), .A2(n20565), .B1(n20206), .B2(n20786), .C1(
        n20802), .C2(n20207), .ZN(n20226) );
  AOI22_X1 U23145 ( .A1(n20636), .A2(n20227), .B1(n20635), .B2(n20226), .ZN(
        n20212) );
  INV_X1 U23146 ( .A(n20207), .ZN(n20210) );
  OR3_X1 U23147 ( .A1(n9866), .A2(n20786), .A3(n20208), .ZN(n20568) );
  NOR2_X1 U23148 ( .A1(n20263), .A2(n20568), .ZN(n20209) );
  OAI21_X1 U23149 ( .B1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n20413), .A(
        n20297), .ZN(n20266) );
  OAI21_X1 U23150 ( .B1(n20210), .B2(n20209), .A(n20638), .ZN(n20228) );
  AOI22_X1 U23151 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n20228), .B1(
        n20221), .B2(n20641), .ZN(n20211) );
  OAI211_X1 U23152 ( .C1(n20644), .C2(n20260), .A(n20212), .B(n20211), .ZN(
        P1_U3041) );
  AOI22_X1 U23153 ( .A1(n20646), .A2(n20227), .B1(n20645), .B2(n20226), .ZN(
        n20214) );
  AOI22_X1 U23154 ( .A1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n20228), .B1(
        n20252), .B2(n20647), .ZN(n20213) );
  OAI211_X1 U23155 ( .C1(n20650), .C2(n20231), .A(n20214), .B(n20213), .ZN(
        P1_U3042) );
  AOI22_X1 U23156 ( .A1(n20652), .A2(n20227), .B1(n20651), .B2(n20226), .ZN(
        n20216) );
  AOI22_X1 U23157 ( .A1(P1_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n20228), .B1(
        n20252), .B2(n20542), .ZN(n20215) );
  OAI211_X1 U23158 ( .C1(n20545), .C2(n20231), .A(n20216), .B(n20215), .ZN(
        P1_U3043) );
  AOI22_X1 U23159 ( .A1(n20658), .A2(n20227), .B1(n20657), .B2(n20226), .ZN(
        n20218) );
  AOI22_X1 U23160 ( .A1(P1_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n20228), .B1(
        n20252), .B2(n20659), .ZN(n20217) );
  OAI211_X1 U23161 ( .C1(n20662), .C2(n20231), .A(n20218), .B(n20217), .ZN(
        P1_U3044) );
  AOI22_X1 U23162 ( .A1(n20664), .A2(n20227), .B1(n20663), .B2(n20226), .ZN(
        n20220) );
  AOI22_X1 U23163 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n20228), .B1(
        n20221), .B2(n20612), .ZN(n20219) );
  OAI211_X1 U23164 ( .C1(n20615), .C2(n20260), .A(n20220), .B(n20219), .ZN(
        P1_U3045) );
  AOI22_X1 U23165 ( .A1(n9828), .A2(n20227), .B1(n20669), .B2(n20226), .ZN(
        n20223) );
  AOI22_X1 U23166 ( .A1(P1_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n20228), .B1(
        n20221), .B2(n20616), .ZN(n20222) );
  OAI211_X1 U23167 ( .C1(n20619), .C2(n20260), .A(n20223), .B(n20222), .ZN(
        P1_U3046) );
  AOI22_X1 U23168 ( .A1(n20676), .A2(n20227), .B1(n20675), .B2(n20226), .ZN(
        n20225) );
  INV_X1 U23169 ( .A(n20682), .ZN(n20552) );
  AOI22_X1 U23170 ( .A1(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n20228), .B1(
        n20252), .B2(n20552), .ZN(n20224) );
  OAI211_X1 U23171 ( .C1(n20555), .C2(n20231), .A(n20225), .B(n20224), .ZN(
        P1_U3047) );
  AOI22_X1 U23172 ( .A1(n20686), .A2(n20227), .B1(n20684), .B2(n20226), .ZN(
        n20230) );
  INV_X1 U23173 ( .A(n20629), .ZN(n20687) );
  AOI22_X1 U23174 ( .A1(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n20228), .B1(
        n20252), .B2(n20687), .ZN(n20229) );
  OAI211_X1 U23175 ( .C1(n20693), .C2(n20231), .A(n20230), .B(n20229), .ZN(
        P1_U3048) );
  NAND3_X1 U23176 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20783), .A3(
        n20461), .ZN(n20269) );
  NOR2_X1 U23177 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20269), .ZN(
        n20255) );
  NAND2_X1 U23178 ( .A1(n9866), .A2(n12574), .ZN(n20348) );
  AOI22_X1 U23179 ( .A1(n20636), .A2(n20255), .B1(n20287), .B2(n20524), .ZN(
        n20241) );
  NAND2_X1 U23180 ( .A1(n20260), .A2(n20286), .ZN(n20233) );
  AOI21_X1 U23181 ( .B1(n20233), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n20786), 
        .ZN(n20237) );
  INV_X1 U23182 ( .A(n20234), .ZN(n20265) );
  NAND2_X1 U23183 ( .A1(n20265), .A2(n20591), .ZN(n20238) );
  INV_X1 U23184 ( .A(n20255), .ZN(n20235) );
  AOI22_X1 U23185 ( .A1(n20237), .A2(n20238), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20235), .ZN(n20236) );
  OAI21_X1 U23186 ( .B1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n20465), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n20351) );
  NAND3_X1 U23187 ( .A1(n20467), .A2(n20236), .A3(n20351), .ZN(n20257) );
  INV_X1 U23188 ( .A(n20237), .ZN(n20239) );
  INV_X1 U23189 ( .A(n20465), .ZN(n20407) );
  NAND2_X1 U23190 ( .A1(n20407), .A2(n20783), .ZN(n20354) );
  OAI22_X1 U23191 ( .A1(n20239), .A2(n20238), .B1(n20469), .B2(n20354), .ZN(
        n20256) );
  AOI22_X1 U23192 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n20257), .B1(
        n20635), .B2(n20256), .ZN(n20240) );
  OAI211_X1 U23193 ( .C1(n20539), .C2(n20260), .A(n20241), .B(n20240), .ZN(
        P1_U3049) );
  AOI22_X1 U23194 ( .A1(n20646), .A2(n20255), .B1(n20287), .B2(n20647), .ZN(
        n20243) );
  AOI22_X1 U23195 ( .A1(P1_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n20257), .B1(
        n20645), .B2(n20256), .ZN(n20242) );
  OAI211_X1 U23196 ( .C1(n20650), .C2(n20260), .A(n20243), .B(n20242), .ZN(
        P1_U3050) );
  AOI22_X1 U23197 ( .A1(n20652), .A2(n20255), .B1(n20287), .B2(n20542), .ZN(
        n20245) );
  AOI22_X1 U23198 ( .A1(P1_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n20257), .B1(
        n20651), .B2(n20256), .ZN(n20244) );
  OAI211_X1 U23199 ( .C1(n20545), .C2(n20260), .A(n20245), .B(n20244), .ZN(
        P1_U3051) );
  AOI22_X1 U23200 ( .A1(n20658), .A2(n20255), .B1(n20287), .B2(n20659), .ZN(
        n20247) );
  AOI22_X1 U23201 ( .A1(P1_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n20257), .B1(
        n20657), .B2(n20256), .ZN(n20246) );
  OAI211_X1 U23202 ( .C1(n20662), .C2(n20260), .A(n20247), .B(n20246), .ZN(
        P1_U3052) );
  INV_X1 U23203 ( .A(n20615), .ZN(n20665) );
  AOI22_X1 U23204 ( .A1(n20664), .A2(n20255), .B1(n20287), .B2(n20665), .ZN(
        n20249) );
  AOI22_X1 U23205 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n20257), .B1(
        n20663), .B2(n20256), .ZN(n20248) );
  OAI211_X1 U23206 ( .C1(n20668), .C2(n20260), .A(n20249), .B(n20248), .ZN(
        P1_U3053) );
  AOI22_X1 U23207 ( .A1(n9828), .A2(n20255), .B1(n20252), .B2(n20616), .ZN(
        n20251) );
  AOI22_X1 U23208 ( .A1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n20257), .B1(
        n20669), .B2(n20256), .ZN(n20250) );
  OAI211_X1 U23209 ( .C1(n20619), .C2(n20286), .A(n20251), .B(n20250), .ZN(
        P1_U3054) );
  AOI22_X1 U23210 ( .A1(n20676), .A2(n20255), .B1(n20252), .B2(n20677), .ZN(
        n20254) );
  AOI22_X1 U23211 ( .A1(P1_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n20257), .B1(
        n20675), .B2(n20256), .ZN(n20253) );
  OAI211_X1 U23212 ( .C1(n20682), .C2(n20286), .A(n20254), .B(n20253), .ZN(
        P1_U3055) );
  AOI22_X1 U23213 ( .A1(n20686), .A2(n20255), .B1(n20287), .B2(n20687), .ZN(
        n20259) );
  AOI22_X1 U23214 ( .A1(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n20257), .B1(
        n20684), .B2(n20256), .ZN(n20258) );
  OAI211_X1 U23215 ( .C1(n20693), .C2(n20260), .A(n20259), .B(n20258), .ZN(
        P1_U3056) );
  INV_X1 U23216 ( .A(n20501), .ZN(n20261) );
  AOI22_X1 U23217 ( .A1(n20636), .A2(n10275), .B1(n20311), .B2(n20524), .ZN(
        n20273) );
  AOI21_X1 U23218 ( .B1(n20263), .B2(n20500), .A(n20262), .ZN(n20270) );
  AND2_X1 U23219 ( .A1(n20264), .A2(n10551), .ZN(n20631) );
  AOI21_X1 U23220 ( .B1(n20265), .B2(n20631), .A(n10275), .ZN(n20271) );
  INV_X1 U23221 ( .A(n20271), .ZN(n20268) );
  AOI21_X1 U23222 ( .B1(n20786), .B2(n20269), .A(n20266), .ZN(n20267) );
  OAI21_X1 U23223 ( .B1(n20270), .B2(n20268), .A(n20267), .ZN(n20289) );
  OAI22_X1 U23224 ( .A1(n20271), .A2(n20270), .B1(n20802), .B2(n20269), .ZN(
        n20288) );
  AOI22_X1 U23225 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n20289), .B1(
        n20635), .B2(n20288), .ZN(n20272) );
  OAI211_X1 U23226 ( .C1(n20539), .C2(n20286), .A(n20273), .B(n20272), .ZN(
        P1_U3057) );
  AOI22_X1 U23227 ( .A1(n20646), .A2(n10275), .B1(n20311), .B2(n20647), .ZN(
        n20275) );
  AOI22_X1 U23228 ( .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n20289), .B1(
        n20645), .B2(n20288), .ZN(n20274) );
  OAI211_X1 U23229 ( .C1(n20650), .C2(n20286), .A(n20275), .B(n20274), .ZN(
        P1_U3058) );
  AOI22_X1 U23230 ( .A1(n20652), .A2(n10275), .B1(n20287), .B2(n20653), .ZN(
        n20277) );
  AOI22_X1 U23231 ( .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n20289), .B1(
        n20651), .B2(n20288), .ZN(n20276) );
  OAI211_X1 U23232 ( .C1(n20656), .C2(n20319), .A(n20277), .B(n20276), .ZN(
        P1_U3059) );
  AOI22_X1 U23233 ( .A1(n20658), .A2(n10275), .B1(n20311), .B2(n20659), .ZN(
        n20279) );
  AOI22_X1 U23234 ( .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20289), .B1(
        n20657), .B2(n20288), .ZN(n20278) );
  OAI211_X1 U23235 ( .C1(n20662), .C2(n20286), .A(n20279), .B(n20278), .ZN(
        P1_U3060) );
  AOI22_X1 U23236 ( .A1(n20664), .A2(n10275), .B1(n20311), .B2(n20665), .ZN(
        n20281) );
  AOI22_X1 U23237 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n20289), .B1(
        n20663), .B2(n20288), .ZN(n20280) );
  OAI211_X1 U23238 ( .C1(n20668), .C2(n20286), .A(n20281), .B(n20280), .ZN(
        P1_U3061) );
  INV_X1 U23239 ( .A(n20619), .ZN(n20671) );
  AOI22_X1 U23240 ( .A1(n9828), .A2(n10275), .B1(n20311), .B2(n20671), .ZN(
        n20283) );
  AOI22_X1 U23241 ( .A1(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n20289), .B1(
        n20669), .B2(n20288), .ZN(n20282) );
  OAI211_X1 U23242 ( .C1(n20674), .C2(n20286), .A(n20283), .B(n20282), .ZN(
        P1_U3062) );
  AOI22_X1 U23243 ( .A1(n20676), .A2(n10275), .B1(n20311), .B2(n20552), .ZN(
        n20285) );
  AOI22_X1 U23244 ( .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20289), .B1(
        n20675), .B2(n20288), .ZN(n20284) );
  OAI211_X1 U23245 ( .C1(n20555), .C2(n20286), .A(n20285), .B(n20284), .ZN(
        P1_U3063) );
  AOI22_X1 U23246 ( .A1(n20686), .A2(n10275), .B1(n20287), .B2(n20624), .ZN(
        n20291) );
  AOI22_X1 U23247 ( .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n20289), .B1(
        n20684), .B2(n20288), .ZN(n20290) );
  OAI211_X1 U23248 ( .C1(n20629), .C2(n20319), .A(n20291), .B(n20290), .ZN(
        P1_U3064) );
  NAND3_X1 U23249 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n20783), .A3(
        n20523), .ZN(n20323) );
  NOR2_X1 U23250 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20323), .ZN(
        n20315) );
  NOR2_X1 U23251 ( .A1(n13707), .A2(n20292), .ZN(n20379) );
  NAND2_X1 U23252 ( .A1(n20379), .A2(n20529), .ZN(n20295) );
  OAI22_X1 U23253 ( .A1(n20295), .A2(n20786), .B1(n20593), .B2(n20293), .ZN(
        n20314) );
  AOI22_X1 U23254 ( .A1(n20636), .A2(n20315), .B1(n20635), .B2(n20314), .ZN(
        n20300) );
  NAND2_X1 U23255 ( .A1(n20320), .A2(n12574), .ZN(n20335) );
  OAI21_X1 U23256 ( .B1(n20344), .B2(n20311), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20296) );
  AOI21_X1 U23257 ( .B1(n20296), .B2(n20295), .A(P1_STATE2_REG_3__SCAN_IN), 
        .ZN(n20298) );
  AOI22_X1 U23258 ( .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n20316), .B1(
        n20344), .B2(n20524), .ZN(n20299) );
  OAI211_X1 U23259 ( .C1(n20539), .C2(n20319), .A(n20300), .B(n20299), .ZN(
        P1_U3065) );
  AOI22_X1 U23260 ( .A1(n20646), .A2(n20315), .B1(n20645), .B2(n20314), .ZN(
        n20302) );
  AOI22_X1 U23261 ( .A1(P1_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n20316), .B1(
        n20344), .B2(n20647), .ZN(n20301) );
  OAI211_X1 U23262 ( .C1(n20650), .C2(n20319), .A(n20302), .B(n20301), .ZN(
        P1_U3066) );
  AOI22_X1 U23263 ( .A1(n20652), .A2(n20315), .B1(n20651), .B2(n20314), .ZN(
        n20304) );
  AOI22_X1 U23264 ( .A1(P1_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n20316), .B1(
        n20344), .B2(n20542), .ZN(n20303) );
  OAI211_X1 U23265 ( .C1(n20545), .C2(n20319), .A(n20304), .B(n20303), .ZN(
        P1_U3067) );
  AOI22_X1 U23266 ( .A1(n20658), .A2(n20315), .B1(n20657), .B2(n20314), .ZN(
        n20306) );
  AOI22_X1 U23267 ( .A1(P1_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n20316), .B1(
        n20344), .B2(n20659), .ZN(n20305) );
  OAI211_X1 U23268 ( .C1(n20662), .C2(n20319), .A(n20306), .B(n20305), .ZN(
        P1_U3068) );
  AOI22_X1 U23269 ( .A1(n20664), .A2(n20315), .B1(n20663), .B2(n20314), .ZN(
        n20308) );
  AOI22_X1 U23270 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n20316), .B1(
        n20344), .B2(n20665), .ZN(n20307) );
  OAI211_X1 U23271 ( .C1(n20668), .C2(n20319), .A(n20308), .B(n20307), .ZN(
        P1_U3069) );
  AOI22_X1 U23272 ( .A1(n9828), .A2(n20315), .B1(n20669), .B2(n20314), .ZN(
        n20310) );
  AOI22_X1 U23273 ( .A1(P1_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n20316), .B1(
        n20311), .B2(n20616), .ZN(n20309) );
  OAI211_X1 U23274 ( .C1(n20619), .C2(n20335), .A(n20310), .B(n20309), .ZN(
        P1_U3070) );
  AOI22_X1 U23275 ( .A1(n20676), .A2(n20315), .B1(n20675), .B2(n20314), .ZN(
        n20313) );
  AOI22_X1 U23276 ( .A1(P1_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n20316), .B1(
        n20311), .B2(n20677), .ZN(n20312) );
  OAI211_X1 U23277 ( .C1(n20682), .C2(n20335), .A(n20313), .B(n20312), .ZN(
        P1_U3071) );
  AOI22_X1 U23278 ( .A1(n20686), .A2(n20315), .B1(n20684), .B2(n20314), .ZN(
        n20318) );
  AOI22_X1 U23279 ( .A1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n20316), .B1(
        n20344), .B2(n20687), .ZN(n20317) );
  OAI211_X1 U23280 ( .C1(n20693), .C2(n20319), .A(n20318), .B(n20317), .ZN(
        P1_U3072) );
  NOR2_X1 U23281 ( .A1(n20790), .A2(n20323), .ZN(n20343) );
  INV_X1 U23282 ( .A(n20379), .ZN(n20322) );
  INV_X1 U23283 ( .A(n20343), .ZN(n20321) );
  OAI222_X1 U23284 ( .A1(n20322), .A2(n20565), .B1(n20321), .B2(n20786), .C1(
        n20802), .C2(n20323), .ZN(n20342) );
  AOI22_X1 U23285 ( .A1(n20636), .A2(n20343), .B1(n20635), .B2(n20342), .ZN(
        n20328) );
  INV_X1 U23286 ( .A(n20323), .ZN(n20326) );
  INV_X1 U23287 ( .A(n20383), .ZN(n20324) );
  NOR2_X1 U23288 ( .A1(n20324), .A2(n20568), .ZN(n20325) );
  OAI21_X1 U23289 ( .B1(n20326), .B2(n20325), .A(n20638), .ZN(n20345) );
  AOI22_X1 U23290 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n20345), .B1(
        n20344), .B2(n20641), .ZN(n20327) );
  OAI211_X1 U23291 ( .C1(n20644), .C2(n20378), .A(n20328), .B(n20327), .ZN(
        P1_U3073) );
  AOI22_X1 U23292 ( .A1(n20646), .A2(n20343), .B1(n20645), .B2(n20342), .ZN(
        n20330) );
  AOI22_X1 U23293 ( .A1(P1_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n20345), .B1(
        n20344), .B2(n20602), .ZN(n20329) );
  OAI211_X1 U23294 ( .C1(n20605), .C2(n20378), .A(n20330), .B(n20329), .ZN(
        P1_U3074) );
  AOI22_X1 U23295 ( .A1(n20652), .A2(n20343), .B1(n20651), .B2(n20342), .ZN(
        n20332) );
  AOI22_X1 U23296 ( .A1(P1_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n20345), .B1(
        n20369), .B2(n20542), .ZN(n20331) );
  OAI211_X1 U23297 ( .C1(n20545), .C2(n20335), .A(n20332), .B(n20331), .ZN(
        P1_U3075) );
  AOI22_X1 U23298 ( .A1(n20658), .A2(n20343), .B1(n20657), .B2(n20342), .ZN(
        n20334) );
  AOI22_X1 U23299 ( .A1(P1_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n20345), .B1(
        n20369), .B2(n20659), .ZN(n20333) );
  OAI211_X1 U23300 ( .C1(n20662), .C2(n20335), .A(n20334), .B(n20333), .ZN(
        P1_U3076) );
  AOI22_X1 U23301 ( .A1(n20664), .A2(n20343), .B1(n20663), .B2(n20342), .ZN(
        n20337) );
  AOI22_X1 U23302 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n20345), .B1(
        n20344), .B2(n20612), .ZN(n20336) );
  OAI211_X1 U23303 ( .C1(n20615), .C2(n20378), .A(n20337), .B(n20336), .ZN(
        P1_U3077) );
  AOI22_X1 U23304 ( .A1(n9828), .A2(n20343), .B1(n20669), .B2(n20342), .ZN(
        n20339) );
  AOI22_X1 U23305 ( .A1(P1_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n20345), .B1(
        n20344), .B2(n20616), .ZN(n20338) );
  OAI211_X1 U23306 ( .C1(n20619), .C2(n20378), .A(n20339), .B(n20338), .ZN(
        P1_U3078) );
  AOI22_X1 U23307 ( .A1(n20676), .A2(n20343), .B1(n20675), .B2(n20342), .ZN(
        n20341) );
  AOI22_X1 U23308 ( .A1(P1_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n20345), .B1(
        n20344), .B2(n20677), .ZN(n20340) );
  OAI211_X1 U23309 ( .C1(n20682), .C2(n20378), .A(n20341), .B(n20340), .ZN(
        P1_U3079) );
  AOI22_X1 U23310 ( .A1(n20686), .A2(n20343), .B1(n20684), .B2(n20342), .ZN(
        n20347) );
  AOI22_X1 U23311 ( .A1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n20345), .B1(
        n20344), .B2(n20624), .ZN(n20346) );
  OAI211_X1 U23312 ( .C1(n20629), .C2(n20378), .A(n20347), .B(n20346), .ZN(
        P1_U3080) );
  INV_X1 U23313 ( .A(n20348), .ZN(n20462) );
  NOR2_X1 U23314 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20380), .ZN(
        n20373) );
  AOI22_X1 U23315 ( .A1(n20636), .A2(n20373), .B1(n20369), .B2(n20641), .ZN(
        n20358) );
  NAND3_X1 U23316 ( .A1(n20378), .A2(n20500), .A3(n20372), .ZN(n20349) );
  NAND2_X1 U23317 ( .A1(n20349), .A2(n20526), .ZN(n20353) );
  NAND2_X1 U23318 ( .A1(n20379), .A2(n20591), .ZN(n20355) );
  INV_X1 U23319 ( .A(n20373), .ZN(n20350) );
  AOI22_X1 U23320 ( .A1(n20353), .A2(n20355), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20350), .ZN(n20352) );
  NAND3_X1 U23321 ( .A1(n20598), .A2(n20352), .A3(n20351), .ZN(n20375) );
  INV_X1 U23322 ( .A(n20353), .ZN(n20356) );
  OAI22_X1 U23323 ( .A1(n20356), .A2(n20355), .B1(n20354), .B2(n20593), .ZN(
        n20374) );
  AOI22_X1 U23324 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n20375), .B1(
        n20635), .B2(n20374), .ZN(n20357) );
  OAI211_X1 U23325 ( .C1(n20644), .C2(n20372), .A(n20358), .B(n20357), .ZN(
        P1_U3081) );
  AOI22_X1 U23326 ( .A1(n20646), .A2(n20373), .B1(n20369), .B2(n20602), .ZN(
        n20360) );
  AOI22_X1 U23327 ( .A1(P1_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n20375), .B1(
        n20645), .B2(n20374), .ZN(n20359) );
  OAI211_X1 U23328 ( .C1(n20605), .C2(n20372), .A(n20360), .B(n20359), .ZN(
        P1_U3082) );
  AOI22_X1 U23329 ( .A1(n20652), .A2(n20373), .B1(n20369), .B2(n20653), .ZN(
        n20362) );
  AOI22_X1 U23330 ( .A1(P1_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n20375), .B1(
        n20651), .B2(n20374), .ZN(n20361) );
  OAI211_X1 U23331 ( .C1(n20656), .C2(n20372), .A(n20362), .B(n20361), .ZN(
        P1_U3083) );
  AOI22_X1 U23332 ( .A1(n20658), .A2(n20373), .B1(n20369), .B2(n20608), .ZN(
        n20364) );
  AOI22_X1 U23333 ( .A1(P1_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n20375), .B1(
        n20657), .B2(n20374), .ZN(n20363) );
  OAI211_X1 U23334 ( .C1(n20611), .C2(n20372), .A(n20364), .B(n20363), .ZN(
        P1_U3084) );
  AOI22_X1 U23335 ( .A1(n20664), .A2(n20373), .B1(n20402), .B2(n20665), .ZN(
        n20366) );
  AOI22_X1 U23336 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n20375), .B1(
        n20663), .B2(n20374), .ZN(n20365) );
  OAI211_X1 U23337 ( .C1(n20668), .C2(n20378), .A(n20366), .B(n20365), .ZN(
        P1_U3085) );
  AOI22_X1 U23338 ( .A1(n9828), .A2(n20373), .B1(n20369), .B2(n20616), .ZN(
        n20368) );
  AOI22_X1 U23339 ( .A1(P1_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n20375), .B1(
        n20669), .B2(n20374), .ZN(n20367) );
  OAI211_X1 U23340 ( .C1(n20619), .C2(n20372), .A(n20368), .B(n20367), .ZN(
        P1_U3086) );
  AOI22_X1 U23341 ( .A1(n20676), .A2(n20373), .B1(n20369), .B2(n20677), .ZN(
        n20371) );
  AOI22_X1 U23342 ( .A1(P1_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n20375), .B1(
        n20675), .B2(n20374), .ZN(n20370) );
  OAI211_X1 U23343 ( .C1(n20682), .C2(n20372), .A(n20371), .B(n20370), .ZN(
        P1_U3087) );
  AOI22_X1 U23344 ( .A1(n20686), .A2(n20373), .B1(n20402), .B2(n20687), .ZN(
        n20377) );
  AOI22_X1 U23345 ( .A1(P1_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n20375), .B1(
        n20684), .B2(n20374), .ZN(n20376) );
  OAI211_X1 U23346 ( .C1(n20693), .C2(n20378), .A(n20377), .B(n20376), .ZN(
        P1_U3088) );
  AOI21_X1 U23347 ( .B1(n20379), .B2(n20631), .A(n20401), .ZN(n20381) );
  OAI22_X1 U23348 ( .A1(n20381), .A2(n20786), .B1(n20380), .B2(n20802), .ZN(
        n20400) );
  AOI22_X1 U23349 ( .A1(n20636), .A2(n20401), .B1(n20635), .B2(n20400), .ZN(
        n20387) );
  NAND2_X1 U23350 ( .A1(n20383), .A2(n20382), .ZN(n20778) );
  INV_X1 U23351 ( .A(n20778), .ZN(n20385) );
  OAI21_X1 U23352 ( .B1(n20385), .B2(n20384), .A(n20638), .ZN(n20403) );
  AOI22_X1 U23353 ( .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n20403), .B1(
        n20402), .B2(n20641), .ZN(n20386) );
  OAI211_X1 U23354 ( .C1(n20644), .C2(n20433), .A(n20387), .B(n20386), .ZN(
        P1_U3089) );
  AOI22_X1 U23355 ( .A1(n20646), .A2(n20401), .B1(n20645), .B2(n20400), .ZN(
        n20389) );
  AOI22_X1 U23356 ( .A1(P1_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n20403), .B1(
        n20402), .B2(n20602), .ZN(n20388) );
  OAI211_X1 U23357 ( .C1(n20605), .C2(n20433), .A(n20389), .B(n20388), .ZN(
        P1_U3090) );
  AOI22_X1 U23358 ( .A1(n20652), .A2(n20401), .B1(n20651), .B2(n20400), .ZN(
        n20391) );
  AOI22_X1 U23359 ( .A1(P1_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n20403), .B1(
        n20402), .B2(n20653), .ZN(n20390) );
  OAI211_X1 U23360 ( .C1(n20656), .C2(n20433), .A(n20391), .B(n20390), .ZN(
        P1_U3091) );
  AOI22_X1 U23361 ( .A1(n20658), .A2(n20401), .B1(n20657), .B2(n20400), .ZN(
        n20393) );
  AOI22_X1 U23362 ( .A1(P1_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n20403), .B1(
        n20402), .B2(n20608), .ZN(n20392) );
  OAI211_X1 U23363 ( .C1(n20611), .C2(n20433), .A(n20393), .B(n20392), .ZN(
        P1_U3092) );
  AOI22_X1 U23364 ( .A1(n20664), .A2(n20401), .B1(n20663), .B2(n20400), .ZN(
        n20395) );
  AOI22_X1 U23365 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n20403), .B1(
        n20402), .B2(n20612), .ZN(n20394) );
  OAI211_X1 U23366 ( .C1(n20615), .C2(n20433), .A(n20395), .B(n20394), .ZN(
        P1_U3093) );
  AOI22_X1 U23367 ( .A1(n9828), .A2(n20401), .B1(n20669), .B2(n20400), .ZN(
        n20397) );
  AOI22_X1 U23368 ( .A1(P1_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n20403), .B1(
        n20402), .B2(n20616), .ZN(n20396) );
  OAI211_X1 U23369 ( .C1(n20619), .C2(n20433), .A(n20397), .B(n20396), .ZN(
        P1_U3094) );
  AOI22_X1 U23370 ( .A1(n20676), .A2(n20401), .B1(n20675), .B2(n20400), .ZN(
        n20399) );
  AOI22_X1 U23371 ( .A1(P1_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n20403), .B1(
        n20402), .B2(n20677), .ZN(n20398) );
  OAI211_X1 U23372 ( .C1(n20682), .C2(n20433), .A(n20399), .B(n20398), .ZN(
        P1_U3095) );
  AOI22_X1 U23373 ( .A1(n20686), .A2(n20401), .B1(n20684), .B2(n20400), .ZN(
        n20405) );
  AOI22_X1 U23374 ( .A1(P1_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n20403), .B1(
        n20402), .B2(n20624), .ZN(n20404) );
  OAI211_X1 U23375 ( .C1(n20629), .C2(n20433), .A(n20405), .B(n20404), .ZN(
        P1_U3096) );
  NAND3_X1 U23376 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n20461), .A3(
        n20523), .ZN(n20435) );
  NOR2_X1 U23377 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20435), .ZN(
        n20429) );
  AOI21_X1 U23378 ( .B1(n9934), .B2(n20529), .A(n20429), .ZN(n20410) );
  NOR2_X1 U23379 ( .A1(n20407), .A2(n20406), .ZN(n20532) );
  INV_X1 U23380 ( .A(n20532), .ZN(n20534) );
  OAI22_X1 U23381 ( .A1(n20410), .A2(n20786), .B1(n20534), .B2(n20469), .ZN(
        n20428) );
  AOI22_X1 U23382 ( .A1(n20636), .A2(n20429), .B1(n20635), .B2(n20428), .ZN(
        n20415) );
  INV_X1 U23383 ( .A(n13917), .ZN(n20408) );
  NAND2_X1 U23384 ( .A1(n20439), .A2(n12574), .ZN(n20460) );
  INV_X1 U23385 ( .A(n20433), .ZN(n20409) );
  OAI21_X1 U23386 ( .B1(n20446), .B2(n20409), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20411) );
  NAND2_X1 U23387 ( .A1(n20411), .A2(n20410), .ZN(n20412) );
  AOI22_X1 U23388 ( .A1(P1_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n20430), .B1(
        n20446), .B2(n20524), .ZN(n20414) );
  OAI211_X1 U23389 ( .C1(n20539), .C2(n20433), .A(n20415), .B(n20414), .ZN(
        P1_U3097) );
  AOI22_X1 U23390 ( .A1(n20646), .A2(n20429), .B1(n20645), .B2(n20428), .ZN(
        n20417) );
  AOI22_X1 U23391 ( .A1(P1_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n20430), .B1(
        n20446), .B2(n20647), .ZN(n20416) );
  OAI211_X1 U23392 ( .C1(n20650), .C2(n20433), .A(n20417), .B(n20416), .ZN(
        P1_U3098) );
  AOI22_X1 U23393 ( .A1(n20652), .A2(n20429), .B1(n20651), .B2(n20428), .ZN(
        n20419) );
  AOI22_X1 U23394 ( .A1(P1_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n20430), .B1(
        n20446), .B2(n20542), .ZN(n20418) );
  OAI211_X1 U23395 ( .C1(n20545), .C2(n20433), .A(n20419), .B(n20418), .ZN(
        P1_U3099) );
  AOI22_X1 U23396 ( .A1(n20658), .A2(n20429), .B1(n20657), .B2(n20428), .ZN(
        n20421) );
  AOI22_X1 U23397 ( .A1(P1_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n20430), .B1(
        n20446), .B2(n20659), .ZN(n20420) );
  OAI211_X1 U23398 ( .C1(n20662), .C2(n20433), .A(n20421), .B(n20420), .ZN(
        P1_U3100) );
  AOI22_X1 U23399 ( .A1(n20664), .A2(n20429), .B1(n20663), .B2(n20428), .ZN(
        n20423) );
  AOI22_X1 U23400 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n20430), .B1(
        n20446), .B2(n20665), .ZN(n20422) );
  OAI211_X1 U23401 ( .C1(n20668), .C2(n20433), .A(n20423), .B(n20422), .ZN(
        P1_U3101) );
  AOI22_X1 U23402 ( .A1(n9828), .A2(n20429), .B1(n20669), .B2(n20428), .ZN(
        n20425) );
  AOI22_X1 U23403 ( .A1(P1_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n20430), .B1(
        n20446), .B2(n20671), .ZN(n20424) );
  OAI211_X1 U23404 ( .C1(n20674), .C2(n20433), .A(n20425), .B(n20424), .ZN(
        P1_U3102) );
  AOI22_X1 U23405 ( .A1(n20676), .A2(n20429), .B1(n20675), .B2(n20428), .ZN(
        n20427) );
  AOI22_X1 U23406 ( .A1(P1_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n20430), .B1(
        n20446), .B2(n20552), .ZN(n20426) );
  OAI211_X1 U23407 ( .C1(n20555), .C2(n20433), .A(n20427), .B(n20426), .ZN(
        P1_U3103) );
  AOI22_X1 U23408 ( .A1(n20686), .A2(n20429), .B1(n20684), .B2(n20428), .ZN(
        n20432) );
  AOI22_X1 U23409 ( .A1(P1_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n20430), .B1(
        n20446), .B2(n20687), .ZN(n20431) );
  OAI211_X1 U23410 ( .C1(n20693), .C2(n20433), .A(n20432), .B(n20431), .ZN(
        P1_U3104) );
  NOR2_X1 U23411 ( .A1(n20790), .A2(n20435), .ZN(n20456) );
  AOI21_X1 U23412 ( .B1(n9934), .B2(n20434), .A(n20456), .ZN(n20436) );
  OAI22_X1 U23413 ( .A1(n20436), .A2(n20786), .B1(n20435), .B2(n20802), .ZN(
        n20455) );
  AOI22_X1 U23414 ( .A1(n20636), .A2(n20456), .B1(n20635), .B2(n20455), .ZN(
        n20441) );
  INV_X1 U23415 ( .A(n20435), .ZN(n20438) );
  NAND2_X1 U23416 ( .A1(n20776), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n20497) );
  NAND2_X1 U23417 ( .A1(n20436), .A2(n20497), .ZN(n20437) );
  OAI221_X1 U23418 ( .B1(n20500), .B2(n20438), .C1(n20786), .C2(n20437), .A(
        n20638), .ZN(n20457) );
  AOI22_X1 U23419 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n20457), .B1(
        n20484), .B2(n20524), .ZN(n20440) );
  OAI211_X1 U23420 ( .C1(n20539), .C2(n20460), .A(n20441), .B(n20440), .ZN(
        P1_U3105) );
  AOI22_X1 U23421 ( .A1(n20646), .A2(n20456), .B1(n20645), .B2(n20455), .ZN(
        n20443) );
  AOI22_X1 U23422 ( .A1(P1_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n20457), .B1(
        n20484), .B2(n20647), .ZN(n20442) );
  OAI211_X1 U23423 ( .C1(n20650), .C2(n20460), .A(n20443), .B(n20442), .ZN(
        P1_U3106) );
  AOI22_X1 U23424 ( .A1(n20652), .A2(n20456), .B1(n20651), .B2(n20455), .ZN(
        n20445) );
  AOI22_X1 U23425 ( .A1(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n20457), .B1(
        n20446), .B2(n20653), .ZN(n20444) );
  OAI211_X1 U23426 ( .C1(n20656), .C2(n20492), .A(n20445), .B(n20444), .ZN(
        P1_U3107) );
  AOI22_X1 U23427 ( .A1(n20658), .A2(n20456), .B1(n20657), .B2(n20455), .ZN(
        n20448) );
  AOI22_X1 U23428 ( .A1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n20457), .B1(
        n20446), .B2(n20608), .ZN(n20447) );
  OAI211_X1 U23429 ( .C1(n20611), .C2(n20492), .A(n20448), .B(n20447), .ZN(
        P1_U3108) );
  AOI22_X1 U23430 ( .A1(n20664), .A2(n20456), .B1(n20663), .B2(n20455), .ZN(
        n20450) );
  AOI22_X1 U23431 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n20457), .B1(
        n20484), .B2(n20665), .ZN(n20449) );
  OAI211_X1 U23432 ( .C1(n20668), .C2(n20460), .A(n20450), .B(n20449), .ZN(
        P1_U3109) );
  AOI22_X1 U23433 ( .A1(n9828), .A2(n20456), .B1(n20669), .B2(n20455), .ZN(
        n20452) );
  AOI22_X1 U23434 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n20457), .B1(
        n20484), .B2(n20671), .ZN(n20451) );
  OAI211_X1 U23435 ( .C1(n20674), .C2(n20460), .A(n20452), .B(n20451), .ZN(
        P1_U3110) );
  AOI22_X1 U23436 ( .A1(n20676), .A2(n20456), .B1(n20675), .B2(n20455), .ZN(
        n20454) );
  AOI22_X1 U23437 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n20457), .B1(
        n20484), .B2(n20552), .ZN(n20453) );
  OAI211_X1 U23438 ( .C1(n20555), .C2(n20460), .A(n20454), .B(n20453), .ZN(
        P1_U3111) );
  AOI22_X1 U23439 ( .A1(n20686), .A2(n20456), .B1(n20684), .B2(n20455), .ZN(
        n20459) );
  AOI22_X1 U23440 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n20457), .B1(
        n20484), .B2(n20687), .ZN(n20458) );
  OAI211_X1 U23441 ( .C1(n20693), .C2(n20460), .A(n20459), .B(n20458), .ZN(
        P1_U3112) );
  NAND3_X1 U23442 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n20461), .ZN(n20494) );
  NOR2_X1 U23443 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20494), .ZN(
        n20487) );
  AOI22_X1 U23444 ( .A1(n20636), .A2(n20487), .B1(n20519), .B2(n20524), .ZN(
        n20473) );
  NAND3_X1 U23445 ( .A1(n20492), .A2(n20500), .A3(n20513), .ZN(n20463) );
  NAND2_X1 U23446 ( .A1(n20463), .A2(n20526), .ZN(n20468) );
  NAND2_X1 U23447 ( .A1(n9934), .A2(n20591), .ZN(n20470) );
  INV_X1 U23448 ( .A(n20487), .ZN(n20464) );
  AOI22_X1 U23449 ( .A1(n20468), .A2(n20470), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20464), .ZN(n20466) );
  OR2_X1 U23450 ( .A1(n20465), .A2(n20783), .ZN(n20592) );
  NAND2_X1 U23451 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20592), .ZN(n20597) );
  NAND3_X1 U23452 ( .A1(n20467), .A2(n20466), .A3(n20597), .ZN(n20489) );
  INV_X1 U23453 ( .A(n20468), .ZN(n20471) );
  AOI22_X1 U23454 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n20489), .B1(
        n20635), .B2(n20488), .ZN(n20472) );
  OAI211_X1 U23455 ( .C1(n20539), .C2(n20492), .A(n20473), .B(n20472), .ZN(
        P1_U3113) );
  AOI22_X1 U23456 ( .A1(n20646), .A2(n20487), .B1(n20484), .B2(n20602), .ZN(
        n20475) );
  AOI22_X1 U23457 ( .A1(P1_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n20489), .B1(
        n20645), .B2(n20488), .ZN(n20474) );
  OAI211_X1 U23458 ( .C1(n20605), .C2(n20513), .A(n20475), .B(n20474), .ZN(
        P1_U3114) );
  AOI22_X1 U23459 ( .A1(n20652), .A2(n20487), .B1(n20484), .B2(n20653), .ZN(
        n20477) );
  AOI22_X1 U23460 ( .A1(P1_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n20489), .B1(
        n20651), .B2(n20488), .ZN(n20476) );
  OAI211_X1 U23461 ( .C1(n20656), .C2(n20513), .A(n20477), .B(n20476), .ZN(
        P1_U3115) );
  AOI22_X1 U23462 ( .A1(n20658), .A2(n20487), .B1(n20519), .B2(n20659), .ZN(
        n20479) );
  AOI22_X1 U23463 ( .A1(P1_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n20489), .B1(
        n20657), .B2(n20488), .ZN(n20478) );
  OAI211_X1 U23464 ( .C1(n20662), .C2(n20492), .A(n20479), .B(n20478), .ZN(
        P1_U3116) );
  AOI22_X1 U23465 ( .A1(n20664), .A2(n20487), .B1(n20484), .B2(n20612), .ZN(
        n20481) );
  AOI22_X1 U23466 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n20489), .B1(
        n20663), .B2(n20488), .ZN(n20480) );
  OAI211_X1 U23467 ( .C1(n20615), .C2(n20513), .A(n20481), .B(n20480), .ZN(
        P1_U3117) );
  AOI22_X1 U23468 ( .A1(n9828), .A2(n20487), .B1(n20519), .B2(n20671), .ZN(
        n20483) );
  AOI22_X1 U23469 ( .A1(P1_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n20489), .B1(
        n20669), .B2(n20488), .ZN(n20482) );
  OAI211_X1 U23470 ( .C1(n20674), .C2(n20492), .A(n20483), .B(n20482), .ZN(
        P1_U3118) );
  AOI22_X1 U23471 ( .A1(n20676), .A2(n20487), .B1(n20484), .B2(n20677), .ZN(
        n20486) );
  AOI22_X1 U23472 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n20489), .B1(
        n20675), .B2(n20488), .ZN(n20485) );
  OAI211_X1 U23473 ( .C1(n20682), .C2(n20513), .A(n20486), .B(n20485), .ZN(
        P1_U3119) );
  AOI22_X1 U23474 ( .A1(n20686), .A2(n20487), .B1(n20519), .B2(n20687), .ZN(
        n20491) );
  AOI22_X1 U23475 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n20489), .B1(
        n20684), .B2(n20488), .ZN(n20490) );
  OAI211_X1 U23476 ( .C1(n20693), .C2(n20492), .A(n20491), .B(n20490), .ZN(
        P1_U3120) );
  AOI21_X1 U23477 ( .B1(n9934), .B2(n20631), .A(n10263), .ZN(n20495) );
  OAI22_X1 U23478 ( .A1(n20495), .A2(n20786), .B1(n20494), .B2(n20802), .ZN(
        n20518) );
  AOI22_X1 U23479 ( .A1(n20636), .A2(n10263), .B1(n20635), .B2(n20518), .ZN(
        n20503) );
  INV_X1 U23480 ( .A(n20494), .ZN(n20499) );
  OAI21_X1 U23481 ( .B1(n20497), .B2(n20496), .A(n20495), .ZN(n20498) );
  OAI221_X1 U23482 ( .B1(n20500), .B2(n20499), .C1(n20786), .C2(n20498), .A(
        n20638), .ZN(n20520) );
  INV_X1 U23483 ( .A(n20561), .ZN(n20510) );
  AOI22_X1 U23484 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n20520), .B1(
        n20510), .B2(n20524), .ZN(n20502) );
  OAI211_X1 U23485 ( .C1(n20539), .C2(n20513), .A(n20503), .B(n20502), .ZN(
        P1_U3121) );
  AOI22_X1 U23486 ( .A1(n20646), .A2(n10263), .B1(n20645), .B2(n20518), .ZN(
        n20505) );
  AOI22_X1 U23487 ( .A1(P1_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n20520), .B1(
        n20519), .B2(n20602), .ZN(n20504) );
  OAI211_X1 U23488 ( .C1(n20605), .C2(n20561), .A(n20505), .B(n20504), .ZN(
        P1_U3122) );
  AOI22_X1 U23489 ( .A1(n20652), .A2(n10263), .B1(n20651), .B2(n20518), .ZN(
        n20507) );
  AOI22_X1 U23490 ( .A1(P1_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n20520), .B1(
        n20519), .B2(n20653), .ZN(n20506) );
  OAI211_X1 U23491 ( .C1(n20656), .C2(n20561), .A(n20507), .B(n20506), .ZN(
        P1_U3123) );
  AOI22_X1 U23492 ( .A1(n20658), .A2(n10263), .B1(n20657), .B2(n20518), .ZN(
        n20509) );
  AOI22_X1 U23493 ( .A1(P1_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n20520), .B1(
        n20510), .B2(n20659), .ZN(n20508) );
  OAI211_X1 U23494 ( .C1(n20662), .C2(n20513), .A(n20509), .B(n20508), .ZN(
        P1_U3124) );
  AOI22_X1 U23495 ( .A1(n20664), .A2(n10263), .B1(n20663), .B2(n20518), .ZN(
        n20512) );
  AOI22_X1 U23496 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n20520), .B1(
        n20510), .B2(n20665), .ZN(n20511) );
  OAI211_X1 U23497 ( .C1(n20668), .C2(n20513), .A(n20512), .B(n20511), .ZN(
        P1_U3125) );
  AOI22_X1 U23498 ( .A1(n9828), .A2(n10263), .B1(n20669), .B2(n20518), .ZN(
        n20515) );
  AOI22_X1 U23499 ( .A1(P1_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n20520), .B1(
        n20519), .B2(n20616), .ZN(n20514) );
  OAI211_X1 U23500 ( .C1(n20619), .C2(n20561), .A(n20515), .B(n20514), .ZN(
        P1_U3126) );
  AOI22_X1 U23501 ( .A1(n20676), .A2(n10263), .B1(n20675), .B2(n20518), .ZN(
        n20517) );
  AOI22_X1 U23502 ( .A1(P1_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n20520), .B1(
        n20519), .B2(n20677), .ZN(n20516) );
  OAI211_X1 U23503 ( .C1(n20682), .C2(n20561), .A(n20517), .B(n20516), .ZN(
        P1_U3127) );
  AOI22_X1 U23504 ( .A1(n20686), .A2(n10263), .B1(n20684), .B2(n20518), .ZN(
        n20522) );
  AOI22_X1 U23505 ( .A1(P1_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n20520), .B1(
        n20519), .B2(n20624), .ZN(n20521) );
  OAI211_X1 U23506 ( .C1(n20629), .C2(n20561), .A(n20522), .B(n20521), .ZN(
        P1_U3128) );
  NAND3_X1 U23507 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n20523), .ZN(n20567) );
  NOR2_X1 U23508 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20567), .ZN(
        n20556) );
  NOR2_X1 U23509 ( .A1(n20569), .A2(n9866), .ZN(n20563) );
  AOI22_X1 U23510 ( .A1(n20636), .A2(n20556), .B1(n20587), .B2(n20524), .ZN(
        n20538) );
  INV_X1 U23511 ( .A(n20587), .ZN(n20525) );
  NAND3_X1 U23512 ( .A1(n20525), .A2(n20500), .A3(n20561), .ZN(n20527) );
  NAND2_X1 U23513 ( .A1(n20527), .A2(n20526), .ZN(n20533) );
  NOR2_X1 U23514 ( .A1(n13707), .A2(n20528), .ZN(n20632) );
  NAND2_X1 U23515 ( .A1(n20632), .A2(n20529), .ZN(n20535) );
  INV_X1 U23516 ( .A(n20556), .ZN(n20530) );
  AOI22_X1 U23517 ( .A1(n20533), .A2(n20535), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20530), .ZN(n20531) );
  OAI211_X1 U23518 ( .C1(n20532), .C2(n20802), .A(n20598), .B(n20531), .ZN(
        n20558) );
  INV_X1 U23519 ( .A(n20533), .ZN(n20536) );
  OAI22_X1 U23520 ( .A1(n20536), .A2(n20535), .B1(n20593), .B2(n20534), .ZN(
        n20557) );
  AOI22_X1 U23521 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n20558), .B1(
        n20635), .B2(n20557), .ZN(n20537) );
  OAI211_X1 U23522 ( .C1(n20539), .C2(n20561), .A(n20538), .B(n20537), .ZN(
        P1_U3129) );
  AOI22_X1 U23523 ( .A1(n20646), .A2(n20556), .B1(n20587), .B2(n20647), .ZN(
        n20541) );
  AOI22_X1 U23524 ( .A1(P1_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n20558), .B1(
        n20645), .B2(n20557), .ZN(n20540) );
  OAI211_X1 U23525 ( .C1(n20650), .C2(n20561), .A(n20541), .B(n20540), .ZN(
        P1_U3130) );
  AOI22_X1 U23526 ( .A1(n20652), .A2(n20556), .B1(n20587), .B2(n20542), .ZN(
        n20544) );
  AOI22_X1 U23527 ( .A1(P1_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n20558), .B1(
        n20651), .B2(n20557), .ZN(n20543) );
  OAI211_X1 U23528 ( .C1(n20545), .C2(n20561), .A(n20544), .B(n20543), .ZN(
        P1_U3131) );
  AOI22_X1 U23529 ( .A1(n20658), .A2(n20556), .B1(n20587), .B2(n20659), .ZN(
        n20547) );
  AOI22_X1 U23530 ( .A1(P1_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n20558), .B1(
        n20657), .B2(n20557), .ZN(n20546) );
  OAI211_X1 U23531 ( .C1(n20662), .C2(n20561), .A(n20547), .B(n20546), .ZN(
        P1_U3132) );
  AOI22_X1 U23532 ( .A1(n20664), .A2(n20556), .B1(n20587), .B2(n20665), .ZN(
        n20549) );
  AOI22_X1 U23533 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n20558), .B1(
        n20663), .B2(n20557), .ZN(n20548) );
  OAI211_X1 U23534 ( .C1(n20668), .C2(n20561), .A(n20549), .B(n20548), .ZN(
        P1_U3133) );
  AOI22_X1 U23535 ( .A1(n9828), .A2(n20556), .B1(n20587), .B2(n20671), .ZN(
        n20551) );
  AOI22_X1 U23536 ( .A1(P1_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n20558), .B1(
        n20669), .B2(n20557), .ZN(n20550) );
  OAI211_X1 U23537 ( .C1(n20674), .C2(n20561), .A(n20551), .B(n20550), .ZN(
        P1_U3134) );
  AOI22_X1 U23538 ( .A1(n20676), .A2(n20556), .B1(n20587), .B2(n20552), .ZN(
        n20554) );
  AOI22_X1 U23539 ( .A1(P1_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n20558), .B1(
        n20675), .B2(n20557), .ZN(n20553) );
  OAI211_X1 U23540 ( .C1(n20555), .C2(n20561), .A(n20554), .B(n20553), .ZN(
        P1_U3135) );
  AOI22_X1 U23541 ( .A1(n20686), .A2(n20556), .B1(n20587), .B2(n20687), .ZN(
        n20560) );
  AOI22_X1 U23542 ( .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n20558), .B1(
        n20684), .B2(n20557), .ZN(n20559) );
  OAI211_X1 U23543 ( .C1(n20693), .C2(n20561), .A(n20560), .B(n20559), .ZN(
        P1_U3136) );
  NAND2_X1 U23544 ( .A1(n20563), .A2(n20562), .ZN(n20594) );
  NOR2_X1 U23545 ( .A1(n20790), .A2(n20567), .ZN(n20586) );
  INV_X1 U23546 ( .A(n20632), .ZN(n20566) );
  INV_X1 U23547 ( .A(n20586), .ZN(n20564) );
  OAI222_X1 U23548 ( .A1(n20566), .A2(n20565), .B1(n20564), .B2(n20786), .C1(
        n20802), .C2(n20567), .ZN(n20585) );
  AOI22_X1 U23549 ( .A1(n20636), .A2(n20586), .B1(n20635), .B2(n20585), .ZN(
        n20572) );
  INV_X1 U23550 ( .A(n20567), .ZN(n20570) );
  NOR2_X1 U23551 ( .A1(n20569), .A2(n20568), .ZN(n20771) );
  OAI21_X1 U23552 ( .B1(n20570), .B2(n20771), .A(n20638), .ZN(n20588) );
  AOI22_X1 U23553 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n20588), .B1(
        n20587), .B2(n20641), .ZN(n20571) );
  OAI211_X1 U23554 ( .C1(n20644), .C2(n20594), .A(n20572), .B(n20571), .ZN(
        P1_U3137) );
  AOI22_X1 U23555 ( .A1(n20646), .A2(n20586), .B1(n20645), .B2(n20585), .ZN(
        n20574) );
  AOI22_X1 U23556 ( .A1(P1_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n20588), .B1(
        n20587), .B2(n20602), .ZN(n20573) );
  OAI211_X1 U23557 ( .C1(n20605), .C2(n20594), .A(n20574), .B(n20573), .ZN(
        P1_U3138) );
  AOI22_X1 U23558 ( .A1(n20652), .A2(n20586), .B1(n20651), .B2(n20585), .ZN(
        n20576) );
  AOI22_X1 U23559 ( .A1(P1_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n20588), .B1(
        n20587), .B2(n20653), .ZN(n20575) );
  OAI211_X1 U23560 ( .C1(n20656), .C2(n20594), .A(n20576), .B(n20575), .ZN(
        P1_U3139) );
  AOI22_X1 U23561 ( .A1(n20658), .A2(n20586), .B1(n20657), .B2(n20585), .ZN(
        n20578) );
  AOI22_X1 U23562 ( .A1(P1_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n20588), .B1(
        n20587), .B2(n20608), .ZN(n20577) );
  OAI211_X1 U23563 ( .C1(n20611), .C2(n20594), .A(n20578), .B(n20577), .ZN(
        P1_U3140) );
  AOI22_X1 U23564 ( .A1(n20664), .A2(n20586), .B1(n20663), .B2(n20585), .ZN(
        n20580) );
  AOI22_X1 U23565 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n20588), .B1(
        n20587), .B2(n20612), .ZN(n20579) );
  OAI211_X1 U23566 ( .C1(n20615), .C2(n20594), .A(n20580), .B(n20579), .ZN(
        P1_U3141) );
  AOI22_X1 U23567 ( .A1(n9828), .A2(n20586), .B1(n20669), .B2(n20585), .ZN(
        n20582) );
  AOI22_X1 U23568 ( .A1(P1_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n20588), .B1(
        n20587), .B2(n20616), .ZN(n20581) );
  OAI211_X1 U23569 ( .C1(n20619), .C2(n20594), .A(n20582), .B(n20581), .ZN(
        P1_U3142) );
  AOI22_X1 U23570 ( .A1(n20676), .A2(n20586), .B1(n20675), .B2(n20585), .ZN(
        n20584) );
  AOI22_X1 U23571 ( .A1(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n20588), .B1(
        n20587), .B2(n20677), .ZN(n20583) );
  OAI211_X1 U23572 ( .C1(n20682), .C2(n20594), .A(n20584), .B(n20583), .ZN(
        P1_U3143) );
  AOI22_X1 U23573 ( .A1(n20686), .A2(n20586), .B1(n20684), .B2(n20585), .ZN(
        n20590) );
  AOI22_X1 U23574 ( .A1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n20588), .B1(
        n20587), .B2(n20624), .ZN(n20589) );
  OAI211_X1 U23575 ( .C1(n20629), .C2(n20594), .A(n20590), .B(n20589), .ZN(
        P1_U3144) );
  NOR2_X1 U23576 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20633), .ZN(
        n20623) );
  NAND2_X1 U23577 ( .A1(n20632), .A2(n20591), .ZN(n20595) );
  OAI22_X1 U23578 ( .A1(n20595), .A2(n20786), .B1(n20593), .B2(n20592), .ZN(
        n20622) );
  AOI22_X1 U23579 ( .A1(n20636), .A2(n20623), .B1(n20635), .B2(n20622), .ZN(
        n20601) );
  INV_X1 U23580 ( .A(n20692), .ZN(n20678) );
  OAI21_X1 U23581 ( .B1(n20678), .B2(n20625), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20596) );
  AOI21_X1 U23582 ( .B1(n20596), .B2(n20595), .A(P1_STATE2_REG_3__SCAN_IN), 
        .ZN(n20599) );
  AOI22_X1 U23583 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n20626), .B1(
        n20625), .B2(n20641), .ZN(n20600) );
  OAI211_X1 U23584 ( .C1(n20644), .C2(n20692), .A(n20601), .B(n20600), .ZN(
        P1_U3145) );
  AOI22_X1 U23585 ( .A1(n20646), .A2(n20623), .B1(n20645), .B2(n20622), .ZN(
        n20604) );
  AOI22_X1 U23586 ( .A1(P1_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n20626), .B1(
        n20625), .B2(n20602), .ZN(n20603) );
  OAI211_X1 U23587 ( .C1(n20605), .C2(n20692), .A(n20604), .B(n20603), .ZN(
        P1_U3146) );
  AOI22_X1 U23588 ( .A1(n20652), .A2(n20623), .B1(n20651), .B2(n20622), .ZN(
        n20607) );
  AOI22_X1 U23589 ( .A1(P1_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n20626), .B1(
        n20625), .B2(n20653), .ZN(n20606) );
  OAI211_X1 U23590 ( .C1(n20656), .C2(n20692), .A(n20607), .B(n20606), .ZN(
        P1_U3147) );
  AOI22_X1 U23591 ( .A1(n20658), .A2(n20623), .B1(n20657), .B2(n20622), .ZN(
        n20610) );
  AOI22_X1 U23592 ( .A1(P1_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n20626), .B1(
        n20625), .B2(n20608), .ZN(n20609) );
  OAI211_X1 U23593 ( .C1(n20611), .C2(n20692), .A(n20610), .B(n20609), .ZN(
        P1_U3148) );
  AOI22_X1 U23594 ( .A1(n20664), .A2(n20623), .B1(n20663), .B2(n20622), .ZN(
        n20614) );
  AOI22_X1 U23595 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n20626), .B1(
        n20625), .B2(n20612), .ZN(n20613) );
  OAI211_X1 U23596 ( .C1(n20615), .C2(n20692), .A(n20614), .B(n20613), .ZN(
        P1_U3149) );
  AOI22_X1 U23597 ( .A1(n9828), .A2(n20623), .B1(n20669), .B2(n20622), .ZN(
        n20618) );
  AOI22_X1 U23598 ( .A1(P1_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n20626), .B1(
        n20625), .B2(n20616), .ZN(n20617) );
  OAI211_X1 U23599 ( .C1(n20619), .C2(n20692), .A(n20618), .B(n20617), .ZN(
        P1_U3150) );
  AOI22_X1 U23600 ( .A1(n20676), .A2(n20623), .B1(n20675), .B2(n20622), .ZN(
        n20621) );
  AOI22_X1 U23601 ( .A1(P1_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n20626), .B1(
        n20625), .B2(n20677), .ZN(n20620) );
  OAI211_X1 U23602 ( .C1(n20682), .C2(n20692), .A(n20621), .B(n20620), .ZN(
        P1_U3151) );
  AOI22_X1 U23603 ( .A1(n20686), .A2(n20623), .B1(n20684), .B2(n20622), .ZN(
        n20628) );
  AOI22_X1 U23604 ( .A1(P1_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n20626), .B1(
        n20625), .B2(n20624), .ZN(n20627) );
  OAI211_X1 U23605 ( .C1(n20629), .C2(n20692), .A(n20628), .B(n20627), .ZN(
        P1_U3152) );
  INV_X1 U23606 ( .A(n20630), .ZN(n20685) );
  AOI21_X1 U23607 ( .B1(n20632), .B2(n20631), .A(n20685), .ZN(n20634) );
  OAI22_X1 U23608 ( .A1(n20634), .A2(n20786), .B1(n20633), .B2(n20802), .ZN(
        n20683) );
  AOI22_X1 U23609 ( .A1(n20636), .A2(n20685), .B1(n20635), .B2(n20683), .ZN(
        n20643) );
  AND2_X1 U23610 ( .A1(n20637), .A2(n20775), .ZN(n20639) );
  OAI21_X1 U23611 ( .B1(n20640), .B2(n20639), .A(n20638), .ZN(n20689) );
  AOI22_X1 U23612 ( .A1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n20689), .B1(
        n20678), .B2(n20641), .ZN(n20642) );
  OAI211_X1 U23613 ( .C1(n20644), .C2(n20681), .A(n20643), .B(n20642), .ZN(
        P1_U3153) );
  AOI22_X1 U23614 ( .A1(n20646), .A2(n20685), .B1(n20645), .B2(n20683), .ZN(
        n20649) );
  AOI22_X1 U23615 ( .A1(P1_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n20689), .B1(
        n20688), .B2(n20647), .ZN(n20648) );
  OAI211_X1 U23616 ( .C1(n20650), .C2(n20692), .A(n20649), .B(n20648), .ZN(
        P1_U3154) );
  AOI22_X1 U23617 ( .A1(n20652), .A2(n20685), .B1(n20651), .B2(n20683), .ZN(
        n20655) );
  AOI22_X1 U23618 ( .A1(P1_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n20689), .B1(
        n20678), .B2(n20653), .ZN(n20654) );
  OAI211_X1 U23619 ( .C1(n20656), .C2(n20681), .A(n20655), .B(n20654), .ZN(
        P1_U3155) );
  AOI22_X1 U23620 ( .A1(n20658), .A2(n20685), .B1(n20657), .B2(n20683), .ZN(
        n20661) );
  AOI22_X1 U23621 ( .A1(P1_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n20689), .B1(
        n20688), .B2(n20659), .ZN(n20660) );
  OAI211_X1 U23622 ( .C1(n20662), .C2(n20692), .A(n20661), .B(n20660), .ZN(
        P1_U3156) );
  AOI22_X1 U23623 ( .A1(n20664), .A2(n20685), .B1(n20663), .B2(n20683), .ZN(
        n20667) );
  AOI22_X1 U23624 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n20689), .B1(
        n20688), .B2(n20665), .ZN(n20666) );
  OAI211_X1 U23625 ( .C1(n20668), .C2(n20692), .A(n20667), .B(n20666), .ZN(
        P1_U3157) );
  AOI22_X1 U23626 ( .A1(n9828), .A2(n20685), .B1(n20669), .B2(n20683), .ZN(
        n20673) );
  AOI22_X1 U23627 ( .A1(P1_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n20689), .B1(
        n20688), .B2(n20671), .ZN(n20672) );
  OAI211_X1 U23628 ( .C1(n20674), .C2(n20692), .A(n20673), .B(n20672), .ZN(
        P1_U3158) );
  AOI22_X1 U23629 ( .A1(n20676), .A2(n20685), .B1(n20675), .B2(n20683), .ZN(
        n20680) );
  AOI22_X1 U23630 ( .A1(P1_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n20689), .B1(
        n20678), .B2(n20677), .ZN(n20679) );
  OAI211_X1 U23631 ( .C1(n20682), .C2(n20681), .A(n20680), .B(n20679), .ZN(
        P1_U3159) );
  AOI22_X1 U23632 ( .A1(n20686), .A2(n20685), .B1(n20684), .B2(n20683), .ZN(
        n20691) );
  AOI22_X1 U23633 ( .A1(P1_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n20689), .B1(
        n20688), .B2(n20687), .ZN(n20690) );
  OAI211_X1 U23634 ( .C1(n20693), .C2(n20692), .A(n20691), .B(n20690), .ZN(
        P1_U3160) );
  AOI21_X1 U23635 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n20806), .A(n20694), 
        .ZN(n20696) );
  NAND2_X1 U23636 ( .A1(n20696), .A2(n20695), .ZN(P1_U3163) );
  AND2_X1 U23637 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n20766), .ZN(
        P1_U3164) );
  AND2_X1 U23638 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n20766), .ZN(
        P1_U3165) );
  AND2_X1 U23639 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n20766), .ZN(
        P1_U3166) );
  AND2_X1 U23640 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n20766), .ZN(
        P1_U3167) );
  INV_X1 U23641 ( .A(P1_DATAWIDTH_REG_27__SCAN_IN), .ZN(n21121) );
  NOR2_X1 U23642 ( .A1(n20770), .A2(n21121), .ZN(P1_U3168) );
  AND2_X1 U23643 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n20766), .ZN(
        P1_U3169) );
  AND2_X1 U23644 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n20766), .ZN(
        P1_U3170) );
  AND2_X1 U23645 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n20766), .ZN(
        P1_U3171) );
  AND2_X1 U23646 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n20766), .ZN(
        P1_U3172) );
  AND2_X1 U23647 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n20766), .ZN(
        P1_U3173) );
  AND2_X1 U23648 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n20766), .ZN(
        P1_U3174) );
  AND2_X1 U23649 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n20766), .ZN(
        P1_U3175) );
  AND2_X1 U23650 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n20766), .ZN(
        P1_U3176) );
  AND2_X1 U23651 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n20766), .ZN(
        P1_U3177) );
  AND2_X1 U23652 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n20766), .ZN(
        P1_U3178) );
  AND2_X1 U23653 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n20766), .ZN(
        P1_U3179) );
  AND2_X1 U23654 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n20766), .ZN(
        P1_U3180) );
  AND2_X1 U23655 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n20766), .ZN(
        P1_U3181) );
  AND2_X1 U23656 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(n20766), .ZN(
        P1_U3182) );
  AND2_X1 U23657 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n20766), .ZN(
        P1_U3183) );
  INV_X1 U23658 ( .A(P1_DATAWIDTH_REG_11__SCAN_IN), .ZN(n21096) );
  NOR2_X1 U23659 ( .A1(n20770), .A2(n21096), .ZN(P1_U3184) );
  AND2_X1 U23660 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n20766), .ZN(
        P1_U3185) );
  AND2_X1 U23661 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n20766), .ZN(P1_U3186) );
  AND2_X1 U23662 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n20766), .ZN(P1_U3187) );
  INV_X1 U23663 ( .A(P1_DATAWIDTH_REG_7__SCAN_IN), .ZN(n21196) );
  NOR2_X1 U23664 ( .A1(n20770), .A2(n21196), .ZN(P1_U3188) );
  AND2_X1 U23665 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n20766), .ZN(P1_U3189) );
  INV_X1 U23666 ( .A(P1_DATAWIDTH_REG_5__SCAN_IN), .ZN(n21042) );
  NOR2_X1 U23667 ( .A1(n20770), .A2(n21042), .ZN(P1_U3190) );
  AND2_X1 U23668 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n20766), .ZN(P1_U3191) );
  AND2_X1 U23669 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n20766), .ZN(P1_U3192) );
  AND2_X1 U23670 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n20766), .ZN(P1_U3193) );
  AOI21_X1 U23671 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n20701), .A(n20704), 
        .ZN(n20709) );
  OR2_X1 U23672 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n20698) );
  OAI21_X1 U23673 ( .B1(P1_STATE_REG_0__SCAN_IN), .B2(n20706), .A(
        P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n20697) );
  AOI21_X1 U23674 ( .B1(HOLD), .B2(n20698), .A(n20697), .ZN(n20699) );
  OAI22_X1 U23675 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20709), .B1(n20814), 
        .B2(n20699), .ZN(P1_U3194) );
  AOI21_X1 U23676 ( .B1(n20701), .B2(n20706), .A(n20700), .ZN(n20711) );
  INV_X1 U23677 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n20703) );
  OAI211_X1 U23678 ( .C1(P1_STATE_REG_2__SCAN_IN), .C2(n20703), .A(
        P1_STATE_REG_0__SCAN_IN), .B(HOLD), .ZN(n20710) );
  INV_X1 U23679 ( .A(n20702), .ZN(n20707) );
  NOR2_X1 U23680 ( .A1(n20704), .A2(n20703), .ZN(n20705) );
  OAI22_X1 U23681 ( .A1(n20707), .A2(n20706), .B1(P1_STATE_REG_2__SCAN_IN), 
        .B2(n20705), .ZN(n20708) );
  OAI22_X1 U23682 ( .A1(n20711), .A2(n20710), .B1(n20709), .B2(n20708), .ZN(
        P1_U3196) );
  NAND2_X1 U23683 ( .A1(n20814), .A2(n20712), .ZN(n20750) );
  INV_X1 U23684 ( .A(P1_ADDRESS_REG_0__SCAN_IN), .ZN(n20713) );
  NAND2_X1 U23685 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20814), .ZN(n20754) );
  OAI222_X1 U23686 ( .A1(n20750), .A2(n13774), .B1(n20713), .B2(n20814), .C1(
        n13701), .C2(n20754), .ZN(P1_U3197) );
  INV_X1 U23687 ( .A(P1_ADDRESS_REG_1__SCAN_IN), .ZN(n20714) );
  OAI222_X1 U23688 ( .A1(n20754), .A2(n13774), .B1(n20714), .B2(n20814), .C1(
        n13935), .C2(n20750), .ZN(P1_U3198) );
  INV_X1 U23689 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n20716) );
  OAI222_X1 U23690 ( .A1(n20754), .A2(n13935), .B1(n20715), .B2(n20814), .C1(
        n20716), .C2(n20750), .ZN(P1_U3199) );
  INV_X1 U23691 ( .A(P1_ADDRESS_REG_3__SCAN_IN), .ZN(n21124) );
  OAI222_X1 U23692 ( .A1(n20750), .A2(n16192), .B1(n21124), .B2(n20814), .C1(
        n20716), .C2(n20754), .ZN(P1_U3200) );
  INV_X1 U23693 ( .A(n20750), .ZN(n20756) );
  AOI22_X1 U23694 ( .A1(P1_ADDRESS_REG_4__SCAN_IN), .A2(n9834), .B1(
        P1_REIP_REG_6__SCAN_IN), .B2(n20756), .ZN(n20717) );
  OAI21_X1 U23695 ( .B1(n16192), .B2(n20754), .A(n20717), .ZN(P1_U3201) );
  INV_X1 U23696 ( .A(P1_REIP_REG_6__SCAN_IN), .ZN(n20719) );
  AOI22_X1 U23697 ( .A1(P1_ADDRESS_REG_5__SCAN_IN), .A2(n9834), .B1(
        P1_REIP_REG_7__SCAN_IN), .B2(n20756), .ZN(n20718) );
  OAI21_X1 U23698 ( .B1(n20719), .B2(n20754), .A(n20718), .ZN(P1_U3202) );
  INV_X1 U23699 ( .A(n20754), .ZN(n20757) );
  AOI22_X1 U23700 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(n9834), .B1(
        P1_REIP_REG_7__SCAN_IN), .B2(n20757), .ZN(n20720) );
  OAI21_X1 U23701 ( .B1(n20721), .B2(n20750), .A(n20720), .ZN(P1_U3203) );
  INV_X1 U23702 ( .A(P1_ADDRESS_REG_7__SCAN_IN), .ZN(n20722) );
  OAI222_X1 U23703 ( .A1(n20750), .A2(n21039), .B1(n20722), .B2(n20814), .C1(
        n20721), .C2(n20754), .ZN(P1_U3204) );
  AOI22_X1 U23704 ( .A1(P1_ADDRESS_REG_8__SCAN_IN), .A2(n9834), .B1(
        P1_REIP_REG_10__SCAN_IN), .B2(n20756), .ZN(n20723) );
  OAI21_X1 U23705 ( .B1(n21039), .B2(n20754), .A(n20723), .ZN(P1_U3205) );
  AOI22_X1 U23706 ( .A1(P1_ADDRESS_REG_9__SCAN_IN), .A2(n9834), .B1(
        P1_REIP_REG_10__SCAN_IN), .B2(n20757), .ZN(n20724) );
  OAI21_X1 U23707 ( .B1(n20725), .B2(n20750), .A(n20724), .ZN(P1_U3206) );
  INV_X1 U23708 ( .A(P1_ADDRESS_REG_10__SCAN_IN), .ZN(n21048) );
  OAI222_X1 U23709 ( .A1(n20754), .A2(n20725), .B1(n21048), .B2(n20814), .C1(
        n20997), .C2(n20750), .ZN(P1_U3207) );
  AOI22_X1 U23710 ( .A1(P1_ADDRESS_REG_11__SCAN_IN), .A2(n9834), .B1(
        P1_REIP_REG_13__SCAN_IN), .B2(n20756), .ZN(n20726) );
  OAI21_X1 U23711 ( .B1(n20997), .B2(n20754), .A(n20726), .ZN(P1_U3208) );
  AOI22_X1 U23712 ( .A1(P1_ADDRESS_REG_12__SCAN_IN), .A2(n9834), .B1(
        P1_REIP_REG_14__SCAN_IN), .B2(n20756), .ZN(n20727) );
  OAI21_X1 U23713 ( .B1(n14928), .B2(n20754), .A(n20727), .ZN(P1_U3209) );
  AOI22_X1 U23714 ( .A1(P1_ADDRESS_REG_13__SCAN_IN), .A2(n9834), .B1(
        P1_REIP_REG_14__SCAN_IN), .B2(n20757), .ZN(n20728) );
  OAI21_X1 U23715 ( .B1(n20730), .B2(n20750), .A(n20728), .ZN(P1_U3210) );
  INV_X1 U23716 ( .A(P1_ADDRESS_REG_14__SCAN_IN), .ZN(n20729) );
  OAI222_X1 U23717 ( .A1(n20754), .A2(n20730), .B1(n20729), .B2(n20814), .C1(
        n15055), .C2(n20750), .ZN(P1_U3211) );
  AOI22_X1 U23718 ( .A1(P1_ADDRESS_REG_15__SCAN_IN), .A2(n9834), .B1(
        P1_REIP_REG_17__SCAN_IN), .B2(n20756), .ZN(n20731) );
  OAI21_X1 U23719 ( .B1(n15055), .B2(n20754), .A(n20731), .ZN(P1_U3212) );
  AOI22_X1 U23720 ( .A1(P1_ADDRESS_REG_16__SCAN_IN), .A2(n9834), .B1(
        P1_REIP_REG_17__SCAN_IN), .B2(n20757), .ZN(n20732) );
  OAI21_X1 U23721 ( .B1(n20733), .B2(n20750), .A(n20732), .ZN(P1_U3213) );
  AOI222_X1 U23722 ( .A1(n20757), .A2(P1_REIP_REG_18__SCAN_IN), .B1(
        P1_ADDRESS_REG_17__SCAN_IN), .B2(n9834), .C1(P1_REIP_REG_19__SCAN_IN), 
        .C2(n20756), .ZN(n20734) );
  INV_X1 U23723 ( .A(n20734), .ZN(P1_U3214) );
  AOI222_X1 U23724 ( .A1(n20756), .A2(P1_REIP_REG_20__SCAN_IN), .B1(
        P1_ADDRESS_REG_18__SCAN_IN), .B2(n9834), .C1(P1_REIP_REG_19__SCAN_IN), 
        .C2(n20757), .ZN(n20735) );
  INV_X1 U23725 ( .A(n20735), .ZN(P1_U3215) );
  INV_X1 U23726 ( .A(P1_ADDRESS_REG_19__SCAN_IN), .ZN(n20737) );
  OAI222_X1 U23727 ( .A1(n20750), .A2(n20739), .B1(n20737), .B2(n20814), .C1(
        n20736), .C2(n20754), .ZN(P1_U3216) );
  INV_X1 U23728 ( .A(P1_ADDRESS_REG_20__SCAN_IN), .ZN(n20738) );
  OAI222_X1 U23729 ( .A1(n20754), .A2(n20739), .B1(n20738), .B2(n20814), .C1(
        n20741), .C2(n20750), .ZN(P1_U3217) );
  AOI22_X1 U23730 ( .A1(P1_ADDRESS_REG_21__SCAN_IN), .A2(n9834), .B1(
        P1_REIP_REG_23__SCAN_IN), .B2(n20756), .ZN(n20740) );
  OAI21_X1 U23731 ( .B1(n20741), .B2(n20754), .A(n20740), .ZN(P1_U3218) );
  AOI22_X1 U23732 ( .A1(P1_ADDRESS_REG_22__SCAN_IN), .A2(n9834), .B1(
        P1_REIP_REG_23__SCAN_IN), .B2(n20757), .ZN(n20742) );
  OAI21_X1 U23733 ( .B1(n20743), .B2(n20750), .A(n20742), .ZN(P1_U3219) );
  AOI222_X1 U23734 ( .A1(n20757), .A2(P1_REIP_REG_24__SCAN_IN), .B1(
        P1_ADDRESS_REG_23__SCAN_IN), .B2(n9834), .C1(P1_REIP_REG_25__SCAN_IN), 
        .C2(n20756), .ZN(n20744) );
  INV_X1 U23735 ( .A(n20744), .ZN(P1_U3220) );
  AOI222_X1 U23736 ( .A1(n20757), .A2(P1_REIP_REG_25__SCAN_IN), .B1(
        P1_ADDRESS_REG_24__SCAN_IN), .B2(n9834), .C1(P1_REIP_REG_26__SCAN_IN), 
        .C2(n20756), .ZN(n20745) );
  INV_X1 U23737 ( .A(n20745), .ZN(P1_U3221) );
  INV_X1 U23738 ( .A(P1_ADDRESS_REG_25__SCAN_IN), .ZN(n20746) );
  OAI222_X1 U23739 ( .A1(n20754), .A2(n20747), .B1(n20746), .B2(n20814), .C1(
        n20749), .C2(n20750), .ZN(P1_U3222) );
  INV_X1 U23740 ( .A(P1_ADDRESS_REG_26__SCAN_IN), .ZN(n20748) );
  OAI222_X1 U23741 ( .A1(n20754), .A2(n20749), .B1(n20748), .B2(n20814), .C1(
        n20753), .C2(n20750), .ZN(P1_U3223) );
  INV_X1 U23742 ( .A(P1_ADDRESS_REG_27__SCAN_IN), .ZN(n20752) );
  OAI222_X1 U23743 ( .A1(n20754), .A2(n20753), .B1(n20752), .B2(n20814), .C1(
        n20751), .C2(n20750), .ZN(P1_U3224) );
  AOI222_X1 U23744 ( .A1(n20756), .A2(P1_REIP_REG_30__SCAN_IN), .B1(
        P1_ADDRESS_REG_28__SCAN_IN), .B2(n9834), .C1(P1_REIP_REG_29__SCAN_IN), 
        .C2(n20757), .ZN(n20755) );
  INV_X1 U23745 ( .A(n20755), .ZN(P1_U3225) );
  AOI222_X1 U23746 ( .A1(n20757), .A2(P1_REIP_REG_30__SCAN_IN), .B1(
        P1_ADDRESS_REG_29__SCAN_IN), .B2(n9834), .C1(P1_REIP_REG_31__SCAN_IN), 
        .C2(n20756), .ZN(n20758) );
  INV_X1 U23747 ( .A(n20758), .ZN(P1_U3226) );
  INV_X1 U23748 ( .A(P1_BE_N_REG_3__SCAN_IN), .ZN(n20759) );
  AOI22_X1 U23749 ( .A1(n20814), .A2(n20760), .B1(n20759), .B2(n9834), .ZN(
        P1_U3458) );
  INV_X1 U23750 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n20793) );
  INV_X1 U23751 ( .A(P1_BE_N_REG_2__SCAN_IN), .ZN(n20761) );
  AOI22_X1 U23752 ( .A1(n20814), .A2(n20793), .B1(n20761), .B2(n9834), .ZN(
        P1_U3459) );
  INV_X1 U23753 ( .A(P1_BE_N_REG_1__SCAN_IN), .ZN(n20762) );
  AOI22_X1 U23754 ( .A1(n20814), .A2(n20763), .B1(n20762), .B2(n9834), .ZN(
        P1_U3460) );
  INV_X1 U23755 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n20796) );
  INV_X1 U23756 ( .A(P1_BE_N_REG_0__SCAN_IN), .ZN(n20764) );
  AOI22_X1 U23757 ( .A1(n20814), .A2(n20796), .B1(n20764), .B2(n9834), .ZN(
        P1_U3461) );
  INV_X1 U23758 ( .A(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(n20767) );
  INV_X1 U23759 ( .A(n20768), .ZN(n20765) );
  AOI21_X1 U23760 ( .B1(n20767), .B2(n20766), .A(n20765), .ZN(P1_U3464) );
  OAI21_X1 U23761 ( .B1(n20770), .B2(n20769), .A(n20768), .ZN(P1_U3465) );
  INV_X1 U23762 ( .A(n20771), .ZN(n20780) );
  NAND2_X1 U23763 ( .A1(n20776), .A2(n20775), .ZN(n20777) );
  NAND4_X1 U23764 ( .A1(n20780), .A2(n20779), .A3(n20778), .A4(n20777), .ZN(
        n20781) );
  NAND2_X1 U23765 ( .A1(n20791), .A2(n20781), .ZN(n20782) );
  OAI21_X1 U23766 ( .B1(n20791), .B2(n20783), .A(n20782), .ZN(P1_U3475) );
  OAI22_X1 U23767 ( .A1(n12574), .A2(n20786), .B1(n20785), .B2(n20784), .ZN(
        n20787) );
  OAI21_X1 U23768 ( .B1(n20788), .B2(n20787), .A(n20791), .ZN(n20789) );
  OAI21_X1 U23769 ( .B1(n20791), .B2(n20790), .A(n20789), .ZN(P1_U3478) );
  AOI211_X1 U23770 ( .C1(P1_REIP_REG_0__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_REIP_REG_1__SCAN_IN), .B(
        P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20792) );
  AOI21_X1 U23771 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(P1_REIP_REG_0__SCAN_IN), 
        .A(n20792), .ZN(n20794) );
  AOI22_X1 U23772 ( .A1(n20798), .A2(n20794), .B1(n20793), .B2(n20795), .ZN(
        P1_U3481) );
  NOR2_X1 U23773 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_0__SCAN_IN), 
        .ZN(n20797) );
  AOI22_X1 U23774 ( .A1(n20798), .A2(n20797), .B1(n20796), .B2(n20795), .ZN(
        P1_U3482) );
  AOI22_X1 U23775 ( .A1(n20814), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n20799), 
        .B2(n9834), .ZN(P1_U3483) );
  AOI21_X1 U23776 ( .B1(n20801), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n20800), 
        .ZN(n20804) );
  NOR3_X1 U23777 ( .A1(n20804), .A2(n20803), .A3(n20802), .ZN(n20805) );
  AOI21_X1 U23778 ( .B1(n20807), .B2(n20806), .A(n20805), .ZN(n20813) );
  AOI211_X1 U23779 ( .C1(n20811), .C2(n20810), .A(n20809), .B(n20808), .ZN(
        n20812) );
  MUX2_X1 U23780 ( .A(n20813), .B(P1_REQUESTPENDING_REG_SCAN_IN), .S(n20812), 
        .Z(P1_U3485) );
  MUX2_X1 U23781 ( .A(P1_M_IO_N_REG_SCAN_IN), .B(P1_MEMORYFETCH_REG_SCAN_IN), 
        .S(n20814), .Z(P1_U3486) );
  NAND2_X1 U23782 ( .A1(n20815), .A2(n20816), .ZN(n20817) );
  OAI22_X1 U23783 ( .A1(n20818), .A2(n20817), .B1(P3_BYTEENABLE_REG_1__SCAN_IN), .B2(n20816), .ZN(n21217) );
  OAI22_X1 U23784 ( .A1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(keyinput75), 
        .B1(P1_EBX_REG_11__SCAN_IN), .B2(keyinput77), .ZN(n20819) );
  AOI221_X1 U23785 ( .B1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(keyinput75), 
        .C1(keyinput77), .C2(P1_EBX_REG_11__SCAN_IN), .A(n20819), .ZN(n20826)
         );
  OAI22_X1 U23786 ( .A1(P2_EBX_REG_29__SCAN_IN), .A2(keyinput33), .B1(
        P1_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(keyinput15), .ZN(n20820) );
  AOI221_X1 U23787 ( .B1(P2_EBX_REG_29__SCAN_IN), .B2(keyinput33), .C1(
        keyinput15), .C2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A(n20820), .ZN(
        n20825) );
  OAI22_X1 U23788 ( .A1(DATAI_8_), .A2(keyinput50), .B1(keyinput32), .B2(
        BUF1_REG_1__SCAN_IN), .ZN(n20821) );
  AOI221_X1 U23789 ( .B1(DATAI_8_), .B2(keyinput50), .C1(BUF1_REG_1__SCAN_IN), 
        .C2(keyinput32), .A(n20821), .ZN(n20824) );
  OAI22_X1 U23790 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(keyinput58), .B1(
        keyinput95), .B2(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n20822) );
  AOI221_X1 U23791 ( .B1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B2(keyinput58), 
        .C1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .C2(keyinput95), .A(n20822), 
        .ZN(n20823) );
  NAND4_X1 U23792 ( .A1(n20826), .A2(n20825), .A3(n20824), .A4(n20823), .ZN(
        n20854) );
  OAI22_X1 U23793 ( .A1(P1_INSTQUEUE_REG_15__6__SCAN_IN), .A2(keyinput83), 
        .B1(P2_BE_N_REG_3__SCAN_IN), .B2(keyinput105), .ZN(n20827) );
  AOI221_X1 U23794 ( .B1(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B2(keyinput83), 
        .C1(keyinput105), .C2(P2_BE_N_REG_3__SCAN_IN), .A(n20827), .ZN(n20834)
         );
  OAI22_X1 U23795 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(keyinput90), .B1(keyinput7), .B2(P2_DATAO_REG_27__SCAN_IN), .ZN(n20828) );
  AOI221_X1 U23796 ( .B1(P3_EAX_REG_5__SCAN_IN), .B2(keyinput90), .C1(
        P2_DATAO_REG_27__SCAN_IN), .C2(keyinput7), .A(n20828), .ZN(n20833) );
  OAI22_X1 U23797 ( .A1(P2_INSTQUEUE_REG_13__0__SCAN_IN), .A2(keyinput43), 
        .B1(P1_EBX_REG_25__SCAN_IN), .B2(keyinput37), .ZN(n20829) );
  AOI221_X1 U23798 ( .B1(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B2(keyinput43), 
        .C1(keyinput37), .C2(P1_EBX_REG_25__SCAN_IN), .A(n20829), .ZN(n20832)
         );
  OAI22_X1 U23799 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(keyinput48), .B1(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(keyinput5), .ZN(n20830) );
  AOI221_X1 U23800 ( .B1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B2(keyinput48), 
        .C1(keyinput5), .C2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A(n20830), 
        .ZN(n20831) );
  NAND4_X1 U23801 ( .A1(n20834), .A2(n20833), .A3(n20832), .A4(n20831), .ZN(
        n20853) );
  OAI22_X1 U23802 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(keyinput61), .B1(
        P2_EBX_REG_17__SCAN_IN), .B2(keyinput14), .ZN(n20835) );
  AOI221_X1 U23803 ( .B1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B2(keyinput61), 
        .C1(keyinput14), .C2(P2_EBX_REG_17__SCAN_IN), .A(n20835), .ZN(n20842)
         );
  OAI22_X1 U23804 ( .A1(P1_EBX_REG_12__SCAN_IN), .A2(keyinput34), .B1(
        DATAI_18_), .B2(keyinput20), .ZN(n20836) );
  AOI221_X1 U23805 ( .B1(P1_EBX_REG_12__SCAN_IN), .B2(keyinput34), .C1(
        keyinput20), .C2(DATAI_18_), .A(n20836), .ZN(n20841) );
  OAI22_X1 U23806 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(keyinput49), 
        .B1(keyinput22), .B2(P3_REIP_REG_6__SCAN_IN), .ZN(n20837) );
  AOI221_X1 U23807 ( .B1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(keyinput49), 
        .C1(P3_REIP_REG_6__SCAN_IN), .C2(keyinput22), .A(n20837), .ZN(n20840)
         );
  OAI22_X1 U23808 ( .A1(P1_EAX_REG_13__SCAN_IN), .A2(keyinput0), .B1(
        P2_DATAWIDTH_REG_28__SCAN_IN), .B2(keyinput26), .ZN(n20838) );
  AOI221_X1 U23809 ( .B1(P1_EAX_REG_13__SCAN_IN), .B2(keyinput0), .C1(
        keyinput26), .C2(P2_DATAWIDTH_REG_28__SCAN_IN), .A(n20838), .ZN(n20839) );
  NAND4_X1 U23810 ( .A1(n20842), .A2(n20841), .A3(n20840), .A4(n20839), .ZN(
        n20852) );
  OAI22_X1 U23811 ( .A1(P2_EBX_REG_16__SCAN_IN), .A2(keyinput121), .B1(
        keyinput112), .B2(P1_EAX_REG_29__SCAN_IN), .ZN(n20843) );
  AOI221_X1 U23812 ( .B1(P2_EBX_REG_16__SCAN_IN), .B2(keyinput121), .C1(
        P1_EAX_REG_29__SCAN_IN), .C2(keyinput112), .A(n20843), .ZN(n20850) );
  OAI22_X1 U23813 ( .A1(P1_DATAO_REG_0__SCAN_IN), .A2(keyinput60), .B1(
        keyinput57), .B2(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n20844) );
  AOI221_X1 U23814 ( .B1(P1_DATAO_REG_0__SCAN_IN), .B2(keyinput60), .C1(
        P3_BYTEENABLE_REG_2__SCAN_IN), .C2(keyinput57), .A(n20844), .ZN(n20849) );
  OAI22_X1 U23815 ( .A1(P2_EAX_REG_2__SCAN_IN), .A2(keyinput92), .B1(
        P1_INSTQUEUE_REG_8__5__SCAN_IN), .B2(keyinput97), .ZN(n20845) );
  AOI221_X1 U23816 ( .B1(P2_EAX_REG_2__SCAN_IN), .B2(keyinput92), .C1(
        keyinput97), .C2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .A(n20845), .ZN(
        n20848) );
  OAI22_X1 U23817 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(keyinput63), 
        .B1(keyinput109), .B2(P3_UWORD_REG_11__SCAN_IN), .ZN(n20846) );
  AOI221_X1 U23818 ( .B1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(keyinput63), 
        .C1(P3_UWORD_REG_11__SCAN_IN), .C2(keyinput109), .A(n20846), .ZN(
        n20847) );
  NAND4_X1 U23819 ( .A1(n20850), .A2(n20849), .A3(n20848), .A4(n20847), .ZN(
        n20851) );
  NOR4_X1 U23820 ( .A1(n20854), .A2(n20853), .A3(n20852), .A4(n20851), .ZN(
        n21215) );
  AOI22_X1 U23821 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(keyinput194), .B1(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(keyinput130), .ZN(n20855) );
  OAI221_X1 U23822 ( .B1(P1_DATAWIDTH_REG_7__SCAN_IN), .B2(keyinput194), .C1(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .C2(keyinput130), .A(n20855), .ZN(
        n20862) );
  AOI22_X1 U23823 ( .A1(DATAI_18_), .A2(keyinput148), .B1(
        P1_EAX_REG_29__SCAN_IN), .B2(keyinput240), .ZN(n20856) );
  OAI221_X1 U23824 ( .B1(DATAI_18_), .B2(keyinput148), .C1(
        P1_EAX_REG_29__SCAN_IN), .C2(keyinput240), .A(n20856), .ZN(n20861) );
  AOI22_X1 U23825 ( .A1(P3_DATAO_REG_7__SCAN_IN), .A2(keyinput168), .B1(
        P2_INSTQUEUE_REG_2__2__SCAN_IN), .B2(keyinput235), .ZN(n20857) );
  OAI221_X1 U23826 ( .B1(P3_DATAO_REG_7__SCAN_IN), .B2(keyinput168), .C1(
        P2_INSTQUEUE_REG_2__2__SCAN_IN), .C2(keyinput235), .A(n20857), .ZN(
        n20860) );
  AOI22_X1 U23827 ( .A1(P3_UWORD_REG_11__SCAN_IN), .A2(keyinput237), .B1(
        P3_EAX_REG_5__SCAN_IN), .B2(keyinput218), .ZN(n20858) );
  OAI221_X1 U23828 ( .B1(P3_UWORD_REG_11__SCAN_IN), .B2(keyinput237), .C1(
        P3_EAX_REG_5__SCAN_IN), .C2(keyinput218), .A(n20858), .ZN(n20859) );
  NOR4_X1 U23829 ( .A1(n20862), .A2(n20861), .A3(n20860), .A4(n20859), .ZN(
        n20890) );
  AOI22_X1 U23830 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(keyinput154), .B1(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(keyinput169), .ZN(n20863) );
  OAI221_X1 U23831 ( .B1(P2_DATAWIDTH_REG_28__SCAN_IN), .B2(keyinput154), .C1(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .C2(keyinput169), .A(n20863), 
        .ZN(n20870) );
  AOI22_X1 U23832 ( .A1(P1_DATAO_REG_0__SCAN_IN), .A2(keyinput188), .B1(
        READY11_REG_SCAN_IN), .B2(keyinput231), .ZN(n20864) );
  OAI221_X1 U23833 ( .B1(P1_DATAO_REG_0__SCAN_IN), .B2(keyinput188), .C1(
        READY11_REG_SCAN_IN), .C2(keyinput231), .A(n20864), .ZN(n20869) );
  AOI22_X1 U23834 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(keyinput177), 
        .B1(P1_ADDRESS_REG_10__SCAN_IN), .B2(keyinput196), .ZN(n20865) );
  OAI221_X1 U23835 ( .B1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(keyinput177), 
        .C1(P1_ADDRESS_REG_10__SCAN_IN), .C2(keyinput196), .A(n20865), .ZN(
        n20868) );
  AOI22_X1 U23836 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(keyinput189), 
        .B1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B2(keyinput176), .ZN(n20866) );
  OAI221_X1 U23837 ( .B1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B2(keyinput189), 
        .C1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .C2(keyinput176), .A(n20866), 
        .ZN(n20867) );
  NOR4_X1 U23838 ( .A1(n20870), .A2(n20869), .A3(n20868), .A4(n20867), .ZN(
        n20889) );
  AOI22_X1 U23839 ( .A1(P3_DATAO_REG_21__SCAN_IN), .A2(keyinput213), .B1(
        P1_ADDRESS_REG_3__SCAN_IN), .B2(keyinput138), .ZN(n20871) );
  OAI221_X1 U23840 ( .B1(P3_DATAO_REG_21__SCAN_IN), .B2(keyinput213), .C1(
        P1_ADDRESS_REG_3__SCAN_IN), .C2(keyinput138), .A(n20871), .ZN(n20878)
         );
  AOI22_X1 U23841 ( .A1(P3_ADDRESS_REG_24__SCAN_IN), .A2(keyinput182), .B1(
        P3_EAX_REG_24__SCAN_IN), .B2(keyinput255), .ZN(n20872) );
  OAI221_X1 U23842 ( .B1(P3_ADDRESS_REG_24__SCAN_IN), .B2(keyinput182), .C1(
        P3_EAX_REG_24__SCAN_IN), .C2(keyinput255), .A(n20872), .ZN(n20877) );
  AOI22_X1 U23843 ( .A1(P3_ADDRESS_REG_22__SCAN_IN), .A2(keyinput206), .B1(
        P2_EAX_REG_27__SCAN_IN), .B2(keyinput239), .ZN(n20873) );
  OAI221_X1 U23844 ( .B1(P3_ADDRESS_REG_22__SCAN_IN), .B2(keyinput206), .C1(
        P2_EAX_REG_27__SCAN_IN), .C2(keyinput239), .A(n20873), .ZN(n20876) );
  AOI22_X1 U23845 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(keyinput172), .B1(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(keyinput200), .ZN(n20874) );
  OAI221_X1 U23846 ( .B1(P2_DATAWIDTH_REG_17__SCAN_IN), .B2(keyinput172), .C1(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .C2(keyinput200), .A(n20874), 
        .ZN(n20875) );
  NOR4_X1 U23847 ( .A1(n20878), .A2(n20877), .A3(n20876), .A4(n20875), .ZN(
        n20888) );
  AOI22_X1 U23848 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(keyinput230), .B1(
        P2_INSTQUEUE_REG_7__3__SCAN_IN), .B2(keyinput145), .ZN(n20879) );
  OAI221_X1 U23849 ( .B1(P2_ADDRESS_REG_29__SCAN_IN), .B2(keyinput230), .C1(
        P2_INSTQUEUE_REG_7__3__SCAN_IN), .C2(keyinput145), .A(n20879), .ZN(
        n20886) );
  AOI22_X1 U23850 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(keyinput129), 
        .B1(P1_EBX_REG_12__SCAN_IN), .B2(keyinput162), .ZN(n20880) );
  OAI221_X1 U23851 ( .B1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B2(keyinput129), 
        .C1(P1_EBX_REG_12__SCAN_IN), .C2(keyinput162), .A(n20880), .ZN(n20885)
         );
  AOI22_X1 U23852 ( .A1(P3_BYTEENABLE_REG_2__SCAN_IN), .A2(keyinput185), .B1(
        P1_INSTQUEUE_REG_0__0__SCAN_IN), .B2(keyinput198), .ZN(n20881) );
  OAI221_X1 U23853 ( .B1(P3_BYTEENABLE_REG_2__SCAN_IN), .B2(keyinput185), .C1(
        P1_INSTQUEUE_REG_0__0__SCAN_IN), .C2(keyinput198), .A(n20881), .ZN(
        n20884) );
  AOI22_X1 U23854 ( .A1(P1_D_C_N_REG_SCAN_IN), .A2(keyinput164), .B1(
        P2_INSTQUEUE_REG_11__6__SCAN_IN), .B2(keyinput222), .ZN(n20882) );
  OAI221_X1 U23855 ( .B1(P1_D_C_N_REG_SCAN_IN), .B2(keyinput164), .C1(
        P2_INSTQUEUE_REG_11__6__SCAN_IN), .C2(keyinput222), .A(n20882), .ZN(
        n20883) );
  NOR4_X1 U23856 ( .A1(n20886), .A2(n20885), .A3(n20884), .A4(n20883), .ZN(
        n20887) );
  NAND4_X1 U23857 ( .A1(n20890), .A2(n20889), .A3(n20888), .A4(n20887), .ZN(
        n21037) );
  AOI22_X1 U23858 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(keyinput216), 
        .B1(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(keyinput226), .ZN(n20891)
         );
  OAI221_X1 U23859 ( .B1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .B2(keyinput216), 
        .C1(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .C2(keyinput226), .A(n20891), 
        .ZN(n20898) );
  AOI22_X1 U23860 ( .A1(P3_REQUESTPENDING_REG_SCAN_IN), .A2(keyinput209), .B1(
        P1_INSTQUEUE_REG_0__6__SCAN_IN), .B2(keyinput132), .ZN(n20892) );
  OAI221_X1 U23861 ( .B1(P3_REQUESTPENDING_REG_SCAN_IN), .B2(keyinput209), 
        .C1(P1_INSTQUEUE_REG_0__6__SCAN_IN), .C2(keyinput132), .A(n20892), 
        .ZN(n20897) );
  AOI22_X1 U23862 ( .A1(P2_BYTEENABLE_REG_3__SCAN_IN), .A2(keyinput151), .B1(
        BUF2_REG_8__SCAN_IN), .B2(keyinput219), .ZN(n20893) );
  OAI221_X1 U23863 ( .B1(P2_BYTEENABLE_REG_3__SCAN_IN), .B2(keyinput151), .C1(
        BUF2_REG_8__SCAN_IN), .C2(keyinput219), .A(n20893), .ZN(n20896) );
  AOI22_X1 U23864 ( .A1(P2_REIP_REG_27__SCAN_IN), .A2(keyinput136), .B1(
        P2_EBX_REG_29__SCAN_IN), .B2(keyinput161), .ZN(n20894) );
  OAI221_X1 U23865 ( .B1(P2_REIP_REG_27__SCAN_IN), .B2(keyinput136), .C1(
        P2_EBX_REG_29__SCAN_IN), .C2(keyinput161), .A(n20894), .ZN(n20895) );
  NOR4_X1 U23866 ( .A1(n20898), .A2(n20897), .A3(n20896), .A4(n20895), .ZN(
        n20929) );
  AOI22_X1 U23867 ( .A1(P2_DATAWIDTH_REG_1__SCAN_IN), .A2(keyinput192), .B1(
        P3_INSTQUEUE_REG_10__7__SCAN_IN), .B2(keyinput170), .ZN(n20899) );
  OAI221_X1 U23868 ( .B1(P2_DATAWIDTH_REG_1__SCAN_IN), .B2(keyinput192), .C1(
        P3_INSTQUEUE_REG_10__7__SCAN_IN), .C2(keyinput170), .A(n20899), .ZN(
        n20906) );
  AOI22_X1 U23869 ( .A1(P1_EBX_REG_30__SCAN_IN), .A2(keyinput157), .B1(
        P1_EBX_REG_11__SCAN_IN), .B2(keyinput205), .ZN(n20900) );
  OAI221_X1 U23870 ( .B1(P1_EBX_REG_30__SCAN_IN), .B2(keyinput157), .C1(
        P1_EBX_REG_11__SCAN_IN), .C2(keyinput205), .A(n20900), .ZN(n20905) );
  AOI22_X1 U23871 ( .A1(P1_EAX_REG_11__SCAN_IN), .A2(keyinput253), .B1(
        P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(keyinput131), .ZN(n20901) );
  OAI221_X1 U23872 ( .B1(P1_EAX_REG_11__SCAN_IN), .B2(keyinput253), .C1(
        P1_PHYADDRPOINTER_REG_11__SCAN_IN), .C2(keyinput131), .A(n20901), .ZN(
        n20904) );
  AOI22_X1 U23873 ( .A1(P1_LWORD_REG_5__SCAN_IN), .A2(keyinput141), .B1(
        P1_UWORD_REG_0__SCAN_IN), .B2(keyinput254), .ZN(n20902) );
  OAI221_X1 U23874 ( .B1(P1_LWORD_REG_5__SCAN_IN), .B2(keyinput141), .C1(
        P1_UWORD_REG_0__SCAN_IN), .C2(keyinput254), .A(n20902), .ZN(n20903) );
  NOR4_X1 U23875 ( .A1(n20906), .A2(n20905), .A3(n20904), .A4(n20903), .ZN(
        n20928) );
  AOI22_X1 U23876 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(keyinput208), .B1(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(keyinput144), .ZN(n20907) );
  OAI221_X1 U23877 ( .B1(P1_DATAWIDTH_REG_11__SCAN_IN), .B2(keyinput208), .C1(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .C2(keyinput144), .A(n20907), 
        .ZN(n20914) );
  AOI22_X1 U23878 ( .A1(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(keyinput248), 
        .B1(P2_EBX_REG_17__SCAN_IN), .B2(keyinput142), .ZN(n20908) );
  OAI221_X1 U23879 ( .B1(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(keyinput248), 
        .C1(P2_EBX_REG_17__SCAN_IN), .C2(keyinput142), .A(n20908), .ZN(n20913)
         );
  AOI22_X1 U23880 ( .A1(P1_EBX_REG_8__SCAN_IN), .A2(keyinput193), .B1(
        P2_REIP_REG_2__SCAN_IN), .B2(keyinput180), .ZN(n20909) );
  OAI221_X1 U23881 ( .B1(P1_EBX_REG_8__SCAN_IN), .B2(keyinput193), .C1(
        P2_REIP_REG_2__SCAN_IN), .C2(keyinput180), .A(n20909), .ZN(n20912) );
  AOI22_X1 U23882 ( .A1(P3_ADDRESS_REG_5__SCAN_IN), .A2(keyinput244), .B1(
        BUF1_REG_10__SCAN_IN), .B2(keyinput207), .ZN(n20910) );
  OAI221_X1 U23883 ( .B1(P3_ADDRESS_REG_5__SCAN_IN), .B2(keyinput244), .C1(
        BUF1_REG_10__SCAN_IN), .C2(keyinput207), .A(n20910), .ZN(n20911) );
  NOR4_X1 U23884 ( .A1(n20914), .A2(n20913), .A3(n20912), .A4(n20911), .ZN(
        n20927) );
  AOI22_X1 U23885 ( .A1(n20916), .A2(keyinput133), .B1(keyinput187), .B2(
        n21144), .ZN(n20915) );
  OAI221_X1 U23886 ( .B1(n20916), .B2(keyinput133), .C1(n21144), .C2(
        keyinput187), .A(n20915), .ZN(n20925) );
  AOI22_X1 U23887 ( .A1(P2_EAX_REG_2__SCAN_IN), .A2(keyinput220), .B1(n20918), 
        .B2(keyinput135), .ZN(n20917) );
  OAI221_X1 U23888 ( .B1(P2_EAX_REG_2__SCAN_IN), .B2(keyinput220), .C1(n20918), 
        .C2(keyinput135), .A(n20917), .ZN(n20924) );
  AOI22_X1 U23889 ( .A1(n21111), .A2(keyinput224), .B1(n21141), .B2(
        keyinput146), .ZN(n20919) );
  OAI221_X1 U23890 ( .B1(n21111), .B2(keyinput224), .C1(n21141), .C2(
        keyinput146), .A(n20919), .ZN(n20923) );
  XNOR2_X1 U23891 ( .A(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B(keyinput158), .ZN(
        n20921) );
  XNOR2_X1 U23892 ( .A(keyinput175), .B(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n20920) );
  NAND2_X1 U23893 ( .A1(n20921), .A2(n20920), .ZN(n20922) );
  NOR4_X1 U23894 ( .A1(n20925), .A2(n20924), .A3(n20923), .A4(n20922), .ZN(
        n20926) );
  NAND4_X1 U23895 ( .A1(n20929), .A2(n20928), .A3(n20927), .A4(n20926), .ZN(
        n21036) );
  AOI22_X1 U23896 ( .A1(n21095), .A2(keyinput246), .B1(keyinput201), .B2(
        n20931), .ZN(n20930) );
  OAI221_X1 U23897 ( .B1(n21095), .B2(keyinput246), .C1(n20931), .C2(
        keyinput201), .A(n20930), .ZN(n20941) );
  AOI22_X1 U23898 ( .A1(n20933), .A2(keyinput227), .B1(n21136), .B2(
        keyinput247), .ZN(n20932) );
  OAI221_X1 U23899 ( .B1(n20933), .B2(keyinput227), .C1(n21136), .C2(
        keyinput247), .A(n20932), .ZN(n20940) );
  INV_X1 U23900 ( .A(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n21073) );
  AOI22_X1 U23901 ( .A1(n20935), .A2(keyinput165), .B1(n21073), .B2(
        keyinput179), .ZN(n20934) );
  OAI221_X1 U23902 ( .B1(n20935), .B2(keyinput165), .C1(n21073), .C2(
        keyinput179), .A(n20934), .ZN(n20939) );
  AOI22_X1 U23903 ( .A1(n20937), .A2(keyinput156), .B1(n21142), .B2(
        keyinput243), .ZN(n20936) );
  OAI221_X1 U23904 ( .B1(n20937), .B2(keyinput156), .C1(n21142), .C2(
        keyinput243), .A(n20936), .ZN(n20938) );
  NOR4_X1 U23905 ( .A1(n20941), .A2(n20940), .A3(n20939), .A4(n20938), .ZN(
        n20979) );
  AOI22_X1 U23906 ( .A1(n20943), .A2(keyinput233), .B1(keyinput238), .B2(
        n21107), .ZN(n20942) );
  OAI221_X1 U23907 ( .B1(n20943), .B2(keyinput233), .C1(n21107), .C2(
        keyinput238), .A(n20942), .ZN(n20951) );
  AOI22_X1 U23908 ( .A1(n21045), .A2(keyinput199), .B1(keyinput163), .B2(
        n21042), .ZN(n20944) );
  OAI221_X1 U23909 ( .B1(n21045), .B2(keyinput199), .C1(n21042), .C2(
        keyinput163), .A(n20944), .ZN(n20950) );
  AOI22_X1 U23910 ( .A1(n21120), .A2(keyinput197), .B1(keyinput140), .B2(
        n21041), .ZN(n20945) );
  OAI221_X1 U23911 ( .B1(n21120), .B2(keyinput197), .C1(n21041), .C2(
        keyinput140), .A(n20945), .ZN(n20949) );
  AOI22_X1 U23912 ( .A1(n20947), .A2(keyinput139), .B1(n21145), .B2(
        keyinput241), .ZN(n20946) );
  OAI221_X1 U23913 ( .B1(n20947), .B2(keyinput139), .C1(n21145), .C2(
        keyinput241), .A(n20946), .ZN(n20948) );
  NOR4_X1 U23914 ( .A1(n20951), .A2(n20950), .A3(n20949), .A4(n20948), .ZN(
        n20978) );
  INV_X1 U23915 ( .A(P2_LWORD_REG_13__SCAN_IN), .ZN(n20953) );
  AOI22_X1 U23916 ( .A1(n13974), .A2(keyinput190), .B1(keyinput252), .B2(
        n20953), .ZN(n20952) );
  OAI221_X1 U23917 ( .B1(n13974), .B2(keyinput190), .C1(n20953), .C2(
        keyinput252), .A(n20952), .ZN(n20963) );
  INV_X1 U23918 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n21155) );
  AOI22_X1 U23919 ( .A1(n21155), .A2(keyinput228), .B1(keyinput155), .B2(
        n21127), .ZN(n20954) );
  OAI221_X1 U23920 ( .B1(n21155), .B2(keyinput228), .C1(n21127), .C2(
        keyinput155), .A(n20954), .ZN(n20962) );
  INV_X1 U23921 ( .A(P3_UWORD_REG_7__SCAN_IN), .ZN(n20956) );
  AOI22_X1 U23922 ( .A1(n21060), .A2(keyinput184), .B1(keyinput214), .B2(
        n20956), .ZN(n20955) );
  OAI221_X1 U23923 ( .B1(n21060), .B2(keyinput184), .C1(n20956), .C2(
        keyinput214), .A(n20955), .ZN(n20961) );
  INV_X1 U23924 ( .A(P2_LWORD_REG_0__SCAN_IN), .ZN(n20957) );
  XOR2_X1 U23925 ( .A(n20957), .B(keyinput166), .Z(n20959) );
  XNOR2_X1 U23926 ( .A(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B(keyinput171), .ZN(
        n20958) );
  NAND2_X1 U23927 ( .A1(n20959), .A2(n20958), .ZN(n20960) );
  NOR4_X1 U23928 ( .A1(n20963), .A2(n20962), .A3(n20961), .A4(n20960), .ZN(
        n20977) );
  INV_X1 U23929 ( .A(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n21158) );
  AOI22_X1 U23930 ( .A1(n21087), .A2(keyinput204), .B1(n21158), .B2(
        keyinput232), .ZN(n20964) );
  OAI221_X1 U23931 ( .B1(n21087), .B2(keyinput204), .C1(n21158), .C2(
        keyinput232), .A(n20964), .ZN(n20975) );
  INV_X1 U23932 ( .A(P1_UWORD_REG_4__SCAN_IN), .ZN(n20966) );
  AOI22_X1 U23933 ( .A1(n20967), .A2(keyinput242), .B1(n20966), .B2(
        keyinput173), .ZN(n20965) );
  OAI221_X1 U23934 ( .B1(n20967), .B2(keyinput242), .C1(n20966), .C2(
        keyinput173), .A(n20965), .ZN(n20974) );
  AOI22_X1 U23935 ( .A1(n20969), .A2(keyinput153), .B1(keyinput149), .B2(
        n21154), .ZN(n20968) );
  OAI221_X1 U23936 ( .B1(n20969), .B2(keyinput153), .C1(n21154), .C2(
        keyinput149), .A(n20968), .ZN(n20973) );
  AOI22_X1 U23937 ( .A1(n21138), .A2(keyinput152), .B1(n20971), .B2(
        keyinput128), .ZN(n20970) );
  OAI221_X1 U23938 ( .B1(n21138), .B2(keyinput152), .C1(n20971), .C2(
        keyinput128), .A(n20970), .ZN(n20972) );
  NOR4_X1 U23939 ( .A1(n20975), .A2(n20974), .A3(n20973), .A4(n20972), .ZN(
        n20976) );
  NAND4_X1 U23940 ( .A1(n20979), .A2(n20978), .A3(n20977), .A4(n20976), .ZN(
        n21035) );
  INV_X1 U23941 ( .A(DATAI_8_), .ZN(n20981) );
  AOI22_X1 U23942 ( .A1(n20981), .A2(keyinput178), .B1(keyinput195), .B2(
        n21121), .ZN(n20980) );
  OAI221_X1 U23943 ( .B1(n20981), .B2(keyinput178), .C1(n21121), .C2(
        keyinput195), .A(n20980), .ZN(n20991) );
  AOI22_X1 U23944 ( .A1(n20983), .A2(keyinput191), .B1(n18992), .B2(
        keyinput249), .ZN(n20982) );
  OAI221_X1 U23945 ( .B1(n20983), .B2(keyinput191), .C1(n18992), .C2(
        keyinput249), .A(n20982), .ZN(n20990) );
  INV_X1 U23946 ( .A(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n20984) );
  XOR2_X1 U23947 ( .A(n20984), .B(keyinput186), .Z(n20987) );
  XNOR2_X1 U23948 ( .A(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B(keyinput159), .ZN(
        n20986) );
  XNOR2_X1 U23949 ( .A(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B(keyinput174), .ZN(
        n20985) );
  NAND3_X1 U23950 ( .A1(n20987), .A2(n20986), .A3(n20985), .ZN(n20989) );
  XNOR2_X1 U23951 ( .A(n21058), .B(keyinput212), .ZN(n20988) );
  NOR4_X1 U23952 ( .A1(n20991), .A2(n20990), .A3(n20989), .A4(n20988), .ZN(
        n21033) );
  INV_X1 U23953 ( .A(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n20993) );
  AOI22_X1 U23954 ( .A1(n21123), .A2(keyinput202), .B1(n20993), .B2(
        keyinput225), .ZN(n20992) );
  OAI221_X1 U23955 ( .B1(n21123), .B2(keyinput202), .C1(n20993), .C2(
        keyinput225), .A(n20992), .ZN(n21002) );
  AOI22_X1 U23956 ( .A1(n21047), .A2(keyinput134), .B1(keyinput250), .B2(
        n21055), .ZN(n20994) );
  OAI221_X1 U23957 ( .B1(n21047), .B2(keyinput134), .C1(n21055), .C2(
        keyinput250), .A(n20994), .ZN(n21001) );
  AOI22_X1 U23958 ( .A1(n21039), .A2(keyinput210), .B1(n21089), .B2(
        keyinput245), .ZN(n20995) );
  OAI221_X1 U23959 ( .B1(n21039), .B2(keyinput210), .C1(n21089), .C2(
        keyinput245), .A(n20995), .ZN(n21000) );
  AOI22_X1 U23960 ( .A1(n20998), .A2(keyinput167), .B1(keyinput221), .B2(
        n20997), .ZN(n20996) );
  OAI221_X1 U23961 ( .B1(n20998), .B2(keyinput167), .C1(n20997), .C2(
        keyinput221), .A(n20996), .ZN(n20999) );
  NOR4_X1 U23962 ( .A1(n21002), .A2(n21001), .A3(n21000), .A4(n20999), .ZN(
        n21032) );
  INV_X1 U23963 ( .A(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n21005) );
  INV_X1 U23964 ( .A(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n21004) );
  AOI22_X1 U23965 ( .A1(n21005), .A2(keyinput211), .B1(n21004), .B2(
        keyinput217), .ZN(n21003) );
  OAI221_X1 U23966 ( .B1(n21005), .B2(keyinput211), .C1(n21004), .C2(
        keyinput217), .A(n21003), .ZN(n21017) );
  AOI22_X1 U23967 ( .A1(n21008), .A2(keyinput223), .B1(n21007), .B2(
        keyinput251), .ZN(n21006) );
  OAI221_X1 U23968 ( .B1(n21008), .B2(keyinput223), .C1(n21007), .C2(
        keyinput251), .A(n21006), .ZN(n21016) );
  AOI22_X1 U23969 ( .A1(n21010), .A2(keyinput160), .B1(n21152), .B2(
        keyinput215), .ZN(n21009) );
  OAI221_X1 U23970 ( .B1(n21010), .B2(keyinput160), .C1(n21152), .C2(
        keyinput215), .A(n21009), .ZN(n21015) );
  AOI22_X1 U23971 ( .A1(n21013), .A2(keyinput236), .B1(n21012), .B2(
        keyinput137), .ZN(n21011) );
  OAI221_X1 U23972 ( .B1(n21013), .B2(keyinput236), .C1(n21012), .C2(
        keyinput137), .A(n21011), .ZN(n21014) );
  NOR4_X1 U23973 ( .A1(n21017), .A2(n21016), .A3(n21015), .A4(n21014), .ZN(
        n21031) );
  AOI22_X1 U23974 ( .A1(n21019), .A2(keyinput143), .B1(n11753), .B2(
        keyinput147), .ZN(n21018) );
  OAI221_X1 U23975 ( .B1(n21019), .B2(keyinput143), .C1(n11753), .C2(
        keyinput147), .A(n21018), .ZN(n21029) );
  AOI22_X1 U23976 ( .A1(n21021), .A2(keyinput183), .B1(n21161), .B2(
        keyinput234), .ZN(n21020) );
  OAI221_X1 U23977 ( .B1(n21021), .B2(keyinput183), .C1(n21161), .C2(
        keyinput234), .A(n21020), .ZN(n21028) );
  AOI22_X1 U23978 ( .A1(n21024), .A2(keyinput203), .B1(keyinput150), .B2(
        n21023), .ZN(n21022) );
  OAI221_X1 U23979 ( .B1(n21024), .B2(keyinput203), .C1(n21023), .C2(
        keyinput150), .A(n21022), .ZN(n21027) );
  AOI22_X1 U23980 ( .A1(n21157), .A2(keyinput181), .B1(n21126), .B2(
        keyinput229), .ZN(n21025) );
  OAI221_X1 U23981 ( .B1(n21157), .B2(keyinput181), .C1(n21126), .C2(
        keyinput229), .A(n21025), .ZN(n21026) );
  NOR4_X1 U23982 ( .A1(n21029), .A2(n21028), .A3(n21027), .A4(n21026), .ZN(
        n21030) );
  NAND4_X1 U23983 ( .A1(n21033), .A2(n21032), .A3(n21031), .A4(n21030), .ZN(
        n21034) );
  NOR4_X1 U23984 ( .A1(n21037), .A2(n21036), .A3(n21035), .A4(n21034), .ZN(
        n21172) );
  AOI22_X1 U23985 ( .A1(n21039), .A2(keyinput82), .B1(n13974), .B2(keyinput62), 
        .ZN(n21038) );
  OAI221_X1 U23986 ( .B1(n21039), .B2(keyinput82), .C1(n13974), .C2(keyinput62), .A(n21038), .ZN(n21052) );
  AOI22_X1 U23987 ( .A1(n21042), .A2(keyinput35), .B1(n21041), .B2(keyinput12), 
        .ZN(n21040) );
  OAI221_X1 U23988 ( .B1(n21042), .B2(keyinput35), .C1(n21041), .C2(keyinput12), .A(n21040), .ZN(n21051) );
  AOI22_X1 U23989 ( .A1(n21045), .A2(keyinput71), .B1(n21044), .B2(keyinput107), .ZN(n21043) );
  OAI221_X1 U23990 ( .B1(n21045), .B2(keyinput71), .C1(n21044), .C2(
        keyinput107), .A(n21043), .ZN(n21050) );
  AOI22_X1 U23991 ( .A1(n21048), .A2(keyinput68), .B1(n21047), .B2(keyinput6), 
        .ZN(n21046) );
  OAI221_X1 U23992 ( .B1(n21048), .B2(keyinput68), .C1(n21047), .C2(keyinput6), 
        .A(n21046), .ZN(n21049) );
  NOR4_X1 U23993 ( .A1(n21052), .A2(n21051), .A3(n21050), .A4(n21049), .ZN(
        n21104) );
  AOI22_X1 U23994 ( .A1(n21055), .A2(keyinput122), .B1(n21054), .B2(keyinput91), .ZN(n21053) );
  OAI221_X1 U23995 ( .B1(n21055), .B2(keyinput122), .C1(n21054), .C2(
        keyinput91), .A(n21053), .ZN(n21068) );
  INV_X1 U23996 ( .A(P1_UWORD_REG_0__SCAN_IN), .ZN(n21057) );
  AOI22_X1 U23997 ( .A1(n21058), .A2(keyinput84), .B1(keyinput126), .B2(n21057), .ZN(n21056) );
  OAI221_X1 U23998 ( .B1(n21058), .B2(keyinput84), .C1(n21057), .C2(
        keyinput126), .A(n21056), .ZN(n21067) );
  AOI22_X1 U23999 ( .A1(n21061), .A2(keyinput65), .B1(n21060), .B2(keyinput56), 
        .ZN(n21059) );
  OAI221_X1 U24000 ( .B1(n21061), .B2(keyinput65), .C1(n21060), .C2(keyinput56), .A(n21059), .ZN(n21066) );
  INV_X1 U24001 ( .A(P3_DATAO_REG_21__SCAN_IN), .ZN(n21064) );
  AOI22_X1 U24002 ( .A1(n21064), .A2(keyinput85), .B1(keyinput44), .B2(n21063), 
        .ZN(n21062) );
  OAI221_X1 U24003 ( .B1(n21064), .B2(keyinput85), .C1(n21063), .C2(keyinput44), .A(n21062), .ZN(n21065) );
  NOR4_X1 U24004 ( .A1(n21068), .A2(n21067), .A3(n21066), .A4(n21065), .ZN(
        n21103) );
  AOI22_X1 U24005 ( .A1(n21071), .A2(keyinput79), .B1(n21070), .B2(keyinput16), 
        .ZN(n21069) );
  OAI221_X1 U24006 ( .B1(n21071), .B2(keyinput79), .C1(n21070), .C2(keyinput16), .A(n21069), .ZN(n21084) );
  AOI22_X1 U24007 ( .A1(n21074), .A2(keyinput70), .B1(keyinput51), .B2(n21073), 
        .ZN(n21072) );
  OAI221_X1 U24008 ( .B1(n21074), .B2(keyinput70), .C1(n21073), .C2(keyinput51), .A(n21072), .ZN(n21083) );
  INV_X1 U24009 ( .A(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n21076) );
  AOI22_X1 U24010 ( .A1(n21077), .A2(keyinput116), .B1(n21076), .B2(keyinput4), 
        .ZN(n21075) );
  OAI221_X1 U24011 ( .B1(n21077), .B2(keyinput116), .C1(n21076), .C2(keyinput4), .A(n21075), .ZN(n21082) );
  INV_X1 U24012 ( .A(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n21079) );
  AOI22_X1 U24013 ( .A1(n21080), .A2(keyinput78), .B1(n21079), .B2(keyinput1), 
        .ZN(n21078) );
  OAI221_X1 U24014 ( .B1(n21080), .B2(keyinput78), .C1(n21079), .C2(keyinput1), 
        .A(n21078), .ZN(n21081) );
  NOR4_X1 U24015 ( .A1(n21084), .A2(n21083), .A3(n21082), .A4(n21081), .ZN(
        n21102) );
  AOI22_X1 U24016 ( .A1(n21087), .A2(keyinput76), .B1(n21086), .B2(keyinput41), 
        .ZN(n21085) );
  OAI221_X1 U24017 ( .B1(n21087), .B2(keyinput76), .C1(n21086), .C2(keyinput41), .A(n21085), .ZN(n21100) );
  AOI22_X1 U24018 ( .A1(n21090), .A2(keyinput2), .B1(keyinput117), .B2(n21089), 
        .ZN(n21088) );
  OAI221_X1 U24019 ( .B1(n21090), .B2(keyinput2), .C1(n21089), .C2(keyinput117), .A(n21088), .ZN(n21099) );
  AOI22_X1 U24020 ( .A1(n21093), .A2(keyinput102), .B1(n21092), .B2(keyinput52), .ZN(n21091) );
  OAI221_X1 U24021 ( .B1(n21093), .B2(keyinput102), .C1(n21092), .C2(
        keyinput52), .A(n21091), .ZN(n21098) );
  AOI22_X1 U24022 ( .A1(n21096), .A2(keyinput80), .B1(n21095), .B2(keyinput118), .ZN(n21094) );
  OAI221_X1 U24023 ( .B1(n21096), .B2(keyinput80), .C1(n21095), .C2(
        keyinput118), .A(n21094), .ZN(n21097) );
  NOR4_X1 U24024 ( .A1(n21100), .A2(n21099), .A3(n21098), .A4(n21097), .ZN(
        n21101) );
  NAND4_X1 U24025 ( .A1(n21104), .A2(n21103), .A3(n21102), .A4(n21101), .ZN(
        n21171) );
  AOI22_X1 U24026 ( .A1(n12152), .A2(keyinput94), .B1(keyinput19), .B2(n11753), 
        .ZN(n21105) );
  OAI221_X1 U24027 ( .B1(n12152), .B2(keyinput94), .C1(n11753), .C2(keyinput19), .A(n21105), .ZN(n21118) );
  AOI22_X1 U24028 ( .A1(n21108), .A2(keyinput98), .B1(keyinput110), .B2(n21107), .ZN(n21106) );
  OAI221_X1 U24029 ( .B1(n21108), .B2(keyinput98), .C1(n21107), .C2(
        keyinput110), .A(n21106), .ZN(n21117) );
  AOI22_X1 U24030 ( .A1(n21111), .A2(keyinput96), .B1(n21110), .B2(keyinput29), 
        .ZN(n21109) );
  OAI221_X1 U24031 ( .B1(n21111), .B2(keyinput96), .C1(n21110), .C2(keyinput29), .A(n21109), .ZN(n21116) );
  INV_X1 U24032 ( .A(P3_DATAO_REG_7__SCAN_IN), .ZN(n21114) );
  INV_X1 U24033 ( .A(READY11_REG_SCAN_IN), .ZN(n21113) );
  AOI22_X1 U24034 ( .A1(n21114), .A2(keyinput40), .B1(n21113), .B2(keyinput103), .ZN(n21112) );
  OAI221_X1 U24035 ( .B1(n21114), .B2(keyinput40), .C1(n21113), .C2(
        keyinput103), .A(n21112), .ZN(n21115) );
  NOR4_X1 U24036 ( .A1(n21118), .A2(n21117), .A3(n21116), .A4(n21115), .ZN(
        n21169) );
  AOI22_X1 U24037 ( .A1(n21121), .A2(keyinput67), .B1(n21120), .B2(keyinput69), 
        .ZN(n21119) );
  OAI221_X1 U24038 ( .B1(n21121), .B2(keyinput67), .C1(n21120), .C2(keyinput69), .A(n21119), .ZN(n21133) );
  AOI22_X1 U24039 ( .A1(n21124), .A2(keyinput10), .B1(keyinput74), .B2(n21123), 
        .ZN(n21122) );
  OAI221_X1 U24040 ( .B1(n21124), .B2(keyinput10), .C1(n21123), .C2(keyinput74), .A(n21122), .ZN(n21132) );
  AOI22_X1 U24041 ( .A1(n21127), .A2(keyinput27), .B1(n21126), .B2(keyinput101), .ZN(n21125) );
  OAI221_X1 U24042 ( .B1(n21127), .B2(keyinput27), .C1(n21126), .C2(
        keyinput101), .A(n21125), .ZN(n21131) );
  XNOR2_X1 U24043 ( .A(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B(keyinput30), .ZN(
        n21129) );
  XNOR2_X1 U24044 ( .A(keyinput9), .B(P2_EAX_REG_19__SCAN_IN), .ZN(n21128) );
  NAND2_X1 U24045 ( .A1(n21129), .A2(n21128), .ZN(n21130) );
  NOR4_X1 U24046 ( .A1(n21133), .A2(n21132), .A3(n21131), .A4(n21130), .ZN(
        n21168) );
  AOI22_X1 U24047 ( .A1(n21136), .A2(keyinput119), .B1(n21135), .B2(keyinput47), .ZN(n21134) );
  OAI221_X1 U24048 ( .B1(n21136), .B2(keyinput119), .C1(n21135), .C2(
        keyinput47), .A(n21134), .ZN(n21149) );
  AOI22_X1 U24049 ( .A1(n21139), .A2(keyinput72), .B1(keyinput24), .B2(n21138), 
        .ZN(n21137) );
  OAI221_X1 U24050 ( .B1(n21139), .B2(keyinput72), .C1(n21138), .C2(keyinput24), .A(n21137), .ZN(n21148) );
  AOI22_X1 U24051 ( .A1(n21142), .A2(keyinput115), .B1(keyinput18), .B2(n21141), .ZN(n21140) );
  OAI221_X1 U24052 ( .B1(n21142), .B2(keyinput115), .C1(n21141), .C2(
        keyinput18), .A(n21140), .ZN(n21147) );
  AOI22_X1 U24053 ( .A1(n21145), .A2(keyinput113), .B1(keyinput59), .B2(n21144), .ZN(n21143) );
  OAI221_X1 U24054 ( .B1(n21145), .B2(keyinput113), .C1(n21144), .C2(
        keyinput59), .A(n21143), .ZN(n21146) );
  NOR4_X1 U24055 ( .A1(n21149), .A2(n21148), .A3(n21147), .A4(n21146), .ZN(
        n21167) );
  AOI22_X1 U24056 ( .A1(n21152), .A2(keyinput87), .B1(n21151), .B2(keyinput3), 
        .ZN(n21150) );
  OAI221_X1 U24057 ( .B1(n21152), .B2(keyinput87), .C1(n21151), .C2(keyinput3), 
        .A(n21150), .ZN(n21165) );
  AOI22_X1 U24058 ( .A1(n21155), .A2(keyinput100), .B1(keyinput21), .B2(n21154), .ZN(n21153) );
  OAI221_X1 U24059 ( .B1(n21155), .B2(keyinput100), .C1(n21154), .C2(
        keyinput21), .A(n21153), .ZN(n21164) );
  AOI22_X1 U24060 ( .A1(n21158), .A2(keyinput104), .B1(keyinput53), .B2(n21157), .ZN(n21156) );
  OAI221_X1 U24061 ( .B1(n21158), .B2(keyinput104), .C1(n21157), .C2(
        keyinput53), .A(n21156), .ZN(n21163) );
  AOI22_X1 U24062 ( .A1(n21161), .A2(keyinput106), .B1(keyinput88), .B2(n21160), .ZN(n21159) );
  OAI221_X1 U24063 ( .B1(n21161), .B2(keyinput106), .C1(n21160), .C2(
        keyinput88), .A(n21159), .ZN(n21162) );
  NOR4_X1 U24064 ( .A1(n21165), .A2(n21164), .A3(n21163), .A4(n21162), .ZN(
        n21166) );
  NAND4_X1 U24065 ( .A1(n21169), .A2(n21168), .A3(n21167), .A4(n21166), .ZN(
        n21170) );
  NOR3_X1 U24066 ( .A1(n21172), .A2(n21171), .A3(n21170), .ZN(n21214) );
  OAI22_X1 U24067 ( .A1(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(keyinput39), 
        .B1(keyinput111), .B2(P2_EAX_REG_27__SCAN_IN), .ZN(n21173) );
  AOI221_X1 U24068 ( .B1(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(keyinput39), 
        .C1(P2_EAX_REG_27__SCAN_IN), .C2(keyinput111), .A(n21173), .ZN(n21180)
         );
  OAI22_X1 U24069 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(keyinput31), 
        .B1(P1_REIP_REG_12__SCAN_IN), .B2(keyinput93), .ZN(n21174) );
  AOI221_X1 U24070 ( .B1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B2(keyinput31), 
        .C1(keyinput93), .C2(P1_REIP_REG_12__SCAN_IN), .A(n21174), .ZN(n21179)
         );
  OAI22_X1 U24071 ( .A1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(keyinput55), 
        .B1(P1_D_C_N_REG_SCAN_IN), .B2(keyinput36), .ZN(n21175) );
  AOI221_X1 U24072 ( .B1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(keyinput55), 
        .C1(keyinput36), .C2(P1_D_C_N_REG_SCAN_IN), .A(n21175), .ZN(n21178) );
  OAI22_X1 U24073 ( .A1(P1_INSTQUEUE_REG_8__7__SCAN_IN), .A2(keyinput89), .B1(
        P3_INSTQUEUE_REG_8__6__SCAN_IN), .B2(keyinput123), .ZN(n21176) );
  AOI221_X1 U24074 ( .B1(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B2(keyinput89), 
        .C1(keyinput123), .C2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A(n21176), 
        .ZN(n21177) );
  NAND4_X1 U24075 ( .A1(n21180), .A2(n21179), .A3(n21178), .A4(n21177), .ZN(
        n21212) );
  OAI22_X1 U24076 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(keyinput46), .B1(
        P2_INSTQUEUE_REG_7__3__SCAN_IN), .B2(keyinput17), .ZN(n21181) );
  AOI221_X1 U24077 ( .B1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B2(keyinput46), 
        .C1(keyinput17), .C2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A(n21181), .ZN(
        n21188) );
  OAI22_X1 U24078 ( .A1(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(keyinput120), 
        .B1(keyinput73), .B2(P2_DATAWIDTH_REG_2__SCAN_IN), .ZN(n21182) );
  AOI221_X1 U24079 ( .B1(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(keyinput120), 
        .C1(P2_DATAWIDTH_REG_2__SCAN_IN), .C2(keyinput73), .A(n21182), .ZN(
        n21187) );
  OAI22_X1 U24080 ( .A1(P1_EAX_REG_11__SCAN_IN), .A2(keyinput125), .B1(
        keyinput64), .B2(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n21183) );
  AOI221_X1 U24081 ( .B1(P1_EAX_REG_11__SCAN_IN), .B2(keyinput125), .C1(
        P2_DATAWIDTH_REG_1__SCAN_IN), .C2(keyinput64), .A(n21183), .ZN(n21186)
         );
  OAI22_X1 U24082 ( .A1(P2_LWORD_REG_0__SCAN_IN), .A2(keyinput38), .B1(
        keyinput54), .B2(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n21184) );
  AOI221_X1 U24083 ( .B1(P2_LWORD_REG_0__SCAN_IN), .B2(keyinput38), .C1(
        P3_ADDRESS_REG_24__SCAN_IN), .C2(keyinput54), .A(n21184), .ZN(n21185)
         );
  NAND4_X1 U24084 ( .A1(n21188), .A2(n21187), .A3(n21186), .A4(n21185), .ZN(
        n21211) );
  OAI22_X1 U24085 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(keyinput28), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(keyinput86), .ZN(n21189) );
  AOI221_X1 U24086 ( .B1(P3_EBX_REG_14__SCAN_IN), .B2(keyinput28), .C1(
        keyinput86), .C2(P3_UWORD_REG_7__SCAN_IN), .A(n21189), .ZN(n21200) );
  OAI22_X1 U24087 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(keyinput99), .B1(
        keyinput81), .B2(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n21190) );
  AOI221_X1 U24088 ( .B1(P3_REIP_REG_16__SCAN_IN), .B2(keyinput99), .C1(
        P3_REQUESTPENDING_REG_SCAN_IN), .C2(keyinput81), .A(n21190), .ZN(
        n21199) );
  OAI22_X1 U24089 ( .A1(n21193), .A2(keyinput8), .B1(n21192), .B2(keyinput42), 
        .ZN(n21191) );
  AOI221_X1 U24090 ( .B1(n21193), .B2(keyinput8), .C1(keyinput42), .C2(n21192), 
        .A(n21191), .ZN(n21198) );
  OAI22_X1 U24091 ( .A1(n21196), .A2(keyinput66), .B1(n21195), .B2(keyinput23), 
        .ZN(n21194) );
  AOI221_X1 U24092 ( .B1(n21196), .B2(keyinput66), .C1(keyinput23), .C2(n21195), .A(n21194), .ZN(n21197) );
  NAND4_X1 U24093 ( .A1(n21200), .A2(n21199), .A3(n21198), .A4(n21197), .ZN(
        n21210) );
  OAI22_X1 U24094 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(keyinput108), 
        .B1(keyinput45), .B2(P1_UWORD_REG_4__SCAN_IN), .ZN(n21201) );
  AOI221_X1 U24095 ( .B1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B2(keyinput108), 
        .C1(P1_UWORD_REG_4__SCAN_IN), .C2(keyinput45), .A(n21201), .ZN(n21208)
         );
  OAI22_X1 U24096 ( .A1(P1_LWORD_REG_5__SCAN_IN), .A2(keyinput13), .B1(
        P2_DATAWIDTH_REG_14__SCAN_IN), .B2(keyinput11), .ZN(n21202) );
  AOI221_X1 U24097 ( .B1(P1_LWORD_REG_5__SCAN_IN), .B2(keyinput13), .C1(
        keyinput11), .C2(P2_DATAWIDTH_REG_14__SCAN_IN), .A(n21202), .ZN(n21207) );
  OAI22_X1 U24098 ( .A1(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .A2(keyinput25), 
        .B1(P2_LWORD_REG_13__SCAN_IN), .B2(keyinput124), .ZN(n21203) );
  AOI221_X1 U24099 ( .B1(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(keyinput25), 
        .C1(keyinput124), .C2(P2_LWORD_REG_13__SCAN_IN), .A(n21203), .ZN(
        n21206) );
  OAI22_X1 U24100 ( .A1(P3_EAX_REG_24__SCAN_IN), .A2(keyinput127), .B1(
        keyinput114), .B2(P3_BE_N_REG_3__SCAN_IN), .ZN(n21204) );
  AOI221_X1 U24101 ( .B1(P3_EAX_REG_24__SCAN_IN), .B2(keyinput127), .C1(
        P3_BE_N_REG_3__SCAN_IN), .C2(keyinput114), .A(n21204), .ZN(n21205) );
  NAND4_X1 U24102 ( .A1(n21208), .A2(n21207), .A3(n21206), .A4(n21205), .ZN(
        n21209) );
  NOR4_X1 U24103 ( .A1(n21212), .A2(n21211), .A3(n21210), .A4(n21209), .ZN(
        n21213) );
  NAND3_X1 U24104 ( .A1(n21215), .A2(n21214), .A3(n21213), .ZN(n21216) );
  XOR2_X1 U24105 ( .A(n21217), .B(n21216), .Z(P3_U2638) );
  INV_X2 U11412 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10289) );
  BUF_X1 U11373 ( .A(n17218), .Z(n9832) );
  AND2_X1 U12878 ( .A1(n10575), .A2(n10574), .ZN(n20294) );
  AND2_X2 U14685 ( .A1(n11653), .A2(n12799), .ZN(n11776) );
  NAND3_X1 U11307 ( .A1(n10028), .A2(n13758), .A3(n20806), .ZN(n10027) );
  CLKBUF_X1 U11326 ( .A(n11508), .Z(n11613) );
  CLKBUF_X1 U11361 ( .A(n11184), .Z(n9860) );
  CLKBUF_X1 U11386 ( .A(n13371), .Z(n15892) );
  CLKBUF_X1 U11523 ( .A(n13911), .Z(n9866) );
  CLKBUF_X1 U11571 ( .A(n10422), .Z(n20190) );
  CLKBUF_X1 U11589 ( .A(n14567), .Z(n14581) );
  AND2_X1 U11693 ( .A1(n20704), .A2(P1_STATE_REG_1__SCAN_IN), .ZN(n20814) );
  CLKBUF_X1 U11835 ( .A(n16536), .Z(n16547) );
  OR2_X1 U12105 ( .A1(n20195), .A2(n10418), .ZN(n21218) );
  CLKBUF_X1 U12429 ( .A(n18881), .Z(n17485) );
endmodule

