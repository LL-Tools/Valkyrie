

module b22_C_2inp_gates_syn ( P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, 
        P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, 
        P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, 
        P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, 
        P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, 
        P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, 
        P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, 
        P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, 
        P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, 
        P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, SUB_1596_U4, 
        SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65, SUB_1596_U66, 
        SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70, SUB_1596_U54, 
        SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58, SUB_1596_U59, 
        SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53, U29, U28, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, P1_U3474, 
        P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, P1_U3495, 
        P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513, P1_U3515, 
        P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, 
        P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, 
        P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, 
        P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, 
        P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, 
        P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556, P1_U3557, 
        P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560, P1_U3561, 
        P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, 
        P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, 
        P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, 
        P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588, P1_U3589, 
        P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U4016, 
        P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321, 
        P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314, 
        P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307, 
        P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300, 
        P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417, P2_U3295, 
        P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, 
        P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, 
        P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, 
        P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, 
        P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442, P2_U3445, 
        P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, P2_U3466, 
        P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, P2_U3486, 
        P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492, P2_U3493, 
        P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, 
        P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, 
        P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, 
        P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, 
        P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, P2_U3528, 
        P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, 
        P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, 
        P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, 
        P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, 
        P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531, P2_U3532, 
        P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, 
        P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, 
        P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552, P2_U3553, 
        P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, P2_U3560, 
        P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211, P2_U3210, 
        P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, 
        P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, 
        P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, 
        P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087, P2_U3947, 
        P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290, P3_U3289, 
        P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283, P3_U3282, 
        P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276, P3_U3275, 
        P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269, P3_U3268, 
        P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377, P3_U3263, 
        P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257, P3_U3256, 
        P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250, P3_U3249, 
        P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243, P3_U3242, 
        P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236, P3_U3235, 
        P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402, P3_U3405, 
        P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423, P3_U3426, 
        P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444, P3_U3446, 
        P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452, P3_U3453, 
        P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459, P3_U3460, 
        P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466, P3_U3467, 
        P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473, P3_U3474, 
        P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480, P3_U3481, 
        P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487, P3_U3488, 
        P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230, P3_U3229, 
        P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223, P3_U3222, 
        P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216, P3_U3215, 
        P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209, P3_U3208, 
        P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202, P3_U3201, 
        P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195, P3_U3194, 
        P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188, P3_U3187, 
        P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491, P3_U3492, 
        P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498, P3_U3499, 
        P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505, P3_U3506, 
        P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512, P3_U3513, 
        P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519, P3_U3520, 
        P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179, P3_U3178, 
        P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172, P3_U3171, 
        P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165, P3_U3164, 
        P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158, P3_U3157, 
        P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150, P3_U3897, 
        keyinput127, keyinput126, keyinput125, keyinput124, keyinput123, 
        keyinput122, keyinput121, keyinput120, keyinput119, keyinput118, 
        keyinput117, keyinput116, keyinput115, keyinput114, keyinput113, 
        keyinput112, keyinput111, keyinput110, keyinput109, keyinput108, 
        keyinput107, keyinput106, keyinput105, keyinput104, keyinput103, 
        keyinput102, keyinput101, keyinput100, keyinput99, keyinput98, 
        keyinput97, keyinput96, keyinput95, keyinput94, keyinput93, keyinput92, 
        keyinput91, keyinput90, keyinput89, keyinput88, keyinput87, keyinput86, 
        keyinput85, keyinput84, keyinput83, keyinput82, keyinput81, keyinput80, 
        keyinput79, keyinput78, keyinput77, keyinput76, keyinput75, keyinput74, 
        keyinput73, keyinput72, keyinput71, keyinput70, keyinput69, keyinput68, 
        keyinput67, keyinput66, keyinput65, keyinput64, keyinput63, keyinput62, 
        keyinput61, keyinput60, keyinput59, keyinput58, keyinput57, keyinput56, 
        keyinput55, keyinput54, keyinput53, keyinput52, keyinput51, keyinput50, 
        keyinput49, keyinput48, keyinput47, keyinput46, keyinput45, keyinput44, 
        keyinput43, keyinput42, keyinput41, keyinput40, keyinput39, keyinput38, 
        keyinput37, keyinput36, keyinput35, keyinput34, keyinput33, keyinput32, 
        keyinput31, keyinput30, keyinput29, keyinput28, keyinput27, keyinput26, 
        keyinput25, keyinput24, keyinput23, keyinput22, keyinput21, keyinput20, 
        keyinput19, keyinput18, keyinput17, keyinput16, keyinput15, keyinput14, 
        keyinput13, keyinput12, keyinput11, keyinput10, keyinput9, keyinput8, 
        keyinput7, keyinput6, keyinput5, keyinput4, keyinput3, keyinput2, 
        keyinput1, keyinput0 );
  input P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
         P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
         P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
         P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
         P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
         P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
         P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
         P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
         P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
         P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN,
         P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN,
         P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN,
         P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN,
         P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN,
         P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN,
         P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
         P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN,
         P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN,
         P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN,
         P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN,
         P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN,
         P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
         P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN,
         P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN,
         P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN,
         P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN,
         P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN,
         P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN,
         P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN,
         P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN,
         P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN,
         P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN,
         P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
         P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN,
         P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN,
         P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN,
         P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
         P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
         P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
         P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
         P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
         P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
         P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
         P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
         P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
         P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
         P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
         P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
         P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
         P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
         P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
         P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
         P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
         P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
         P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
         P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
         P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
         P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN,
         P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN,
         P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN,
         P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN,
         P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN,
         P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN,
         P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN,
         P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN,
         P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN,
         P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN,
         P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN,
         P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN,
         P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN,
         P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN,
         P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN,
         P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN,
         P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN,
         P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN,
         P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN,
         P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN,
         P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN,
         P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN,
         P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN,
         P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
         P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN,
         P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN,
         P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
         P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
         P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
         P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
         P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
         P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
         P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
         P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
         P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
         P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
         P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
         P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
         P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN,
         P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN,
         P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
         P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN,
         P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN,
         P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN,
         P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN,
         P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN,
         P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN,
         P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN,
         P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN,
         P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN,
         P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN,
         P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN,
         P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN,
         P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN,
         P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN,
         P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
         P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN,
         P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN,
         P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
         P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
         P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
         P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
         P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
         P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
         P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
         P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
         P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
         P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
         P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
         P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
         P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
         P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
         P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
         P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
         P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput127,
         keyinput126, keyinput125, keyinput124, keyinput123, keyinput122,
         keyinput121, keyinput120, keyinput119, keyinput118, keyinput117,
         keyinput116, keyinput115, keyinput114, keyinput113, keyinput112,
         keyinput111, keyinput110, keyinput109, keyinput108, keyinput107,
         keyinput106, keyinput105, keyinput104, keyinput103, keyinput102,
         keyinput101, keyinput100, keyinput99, keyinput98, keyinput97,
         keyinput96, keyinput95, keyinput94, keyinput93, keyinput92,
         keyinput91, keyinput90, keyinput89, keyinput88, keyinput87,
         keyinput86, keyinput85, keyinput84, keyinput83, keyinput82,
         keyinput81, keyinput80, keyinput79, keyinput78, keyinput77,
         keyinput76, keyinput75, keyinput74, keyinput73, keyinput72,
         keyinput71, keyinput70, keyinput69, keyinput68, keyinput67,
         keyinput66, keyinput65, keyinput64, keyinput63, keyinput62,
         keyinput61, keyinput60, keyinput59, keyinput58, keyinput57,
         keyinput56, keyinput55, keyinput54, keyinput53, keyinput52,
         keyinput51, keyinput50, keyinput49, keyinput48, keyinput47,
         keyinput46, keyinput45, keyinput44, keyinput43, keyinput42,
         keyinput41, keyinput40, keyinput39, keyinput38, keyinput37,
         keyinput36, keyinput35, keyinput34, keyinput33, keyinput32,
         keyinput31, keyinput30, keyinput29, keyinput28, keyinput27,
         keyinput26, keyinput25, keyinput24, keyinput23, keyinput22,
         keyinput21, keyinput20, keyinput19, keyinput18, keyinput17,
         keyinput16, keyinput15, keyinput14, keyinput13, keyinput12,
         keyinput11, keyinput10, keyinput9, keyinput8, keyinput7, keyinput6,
         keyinput5, keyinput4, keyinput3, keyinput2, keyinput1, keyinput0;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n6516, n6517, n6518, n6519, n6520, n6522, n6523, n6525, n6526, n6527,
         n6529, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539,
         n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549,
         n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559,
         n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569,
         n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579,
         n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589,
         n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599,
         n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609,
         n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619,
         n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629,
         n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639,
         n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649,
         n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659,
         n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669,
         n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679,
         n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689,
         n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699,
         n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709,
         n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719,
         n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729,
         n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739,
         n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749,
         n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759,
         n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769,
         n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779,
         n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789,
         n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799,
         n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809,
         n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819,
         n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829,
         n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839,
         n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849,
         n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859,
         n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869,
         n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879,
         n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889,
         n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899,
         n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909,
         n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919,
         n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929,
         n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939,
         n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949,
         n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959,
         n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969,
         n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979,
         n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989,
         n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999,
         n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009,
         n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019,
         n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029,
         n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039,
         n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049,
         n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059,
         n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069,
         n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079,
         n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089,
         n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099,
         n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109,
         n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119,
         n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129,
         n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139,
         n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149,
         n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159,
         n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169,
         n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179,
         n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189,
         n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199,
         n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209,
         n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219,
         n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229,
         n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239,
         n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249,
         n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259,
         n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269,
         n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279,
         n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289,
         n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299,
         n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309,
         n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319,
         n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329,
         n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339,
         n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349,
         n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359,
         n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369,
         n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379,
         n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389,
         n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399,
         n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409,
         n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419,
         n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429,
         n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439,
         n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449,
         n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459,
         n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469,
         n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479,
         n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489,
         n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499,
         n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509,
         n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519,
         n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529,
         n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539,
         n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549,
         n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559,
         n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569,
         n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579,
         n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589,
         n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599,
         n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609,
         n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619,
         n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629,
         n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639,
         n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649,
         n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659,
         n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669,
         n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679,
         n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689,
         n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699,
         n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709,
         n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719,
         n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729,
         n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739,
         n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749,
         n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759,
         n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769,
         n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779,
         n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789,
         n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799,
         n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809,
         n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819,
         n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829,
         n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839,
         n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849,
         n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859,
         n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869,
         n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879,
         n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889,
         n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899,
         n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909,
         n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919,
         n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929,
         n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939,
         n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949,
         n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959,
         n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969,
         n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979,
         n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989,
         n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999,
         n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009,
         n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019,
         n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029,
         n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039,
         n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049,
         n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059,
         n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069,
         n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079,
         n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089,
         n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099,
         n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109,
         n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119,
         n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129,
         n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139,
         n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149,
         n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159,
         n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169,
         n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179,
         n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189,
         n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199,
         n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209,
         n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219,
         n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229,
         n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239,
         n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249,
         n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259,
         n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269,
         n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279,
         n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290,
         n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300,
         n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310,
         n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320,
         n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330,
         n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340,
         n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350,
         n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360,
         n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370,
         n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380,
         n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390,
         n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400,
         n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410,
         n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420,
         n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430,
         n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440,
         n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450,
         n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460,
         n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470,
         n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480,
         n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490,
         n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500,
         n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510,
         n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520,
         n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530,
         n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540,
         n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550,
         n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560,
         n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570,
         n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580,
         n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590,
         n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600,
         n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610,
         n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620,
         n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630,
         n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640,
         n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650,
         n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660,
         n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670,
         n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680,
         n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690,
         n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700,
         n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710,
         n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720,
         n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730,
         n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740,
         n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750,
         n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760,
         n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770,
         n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780,
         n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790,
         n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800,
         n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810,
         n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820,
         n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830,
         n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840,
         n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850,
         n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860,
         n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870,
         n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880,
         n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890,
         n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900,
         n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910,
         n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920,
         n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930,
         n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940,
         n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950,
         n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960,
         n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970,
         n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980,
         n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990,
         n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000,
         n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010,
         n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020,
         n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030,
         n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040,
         n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050,
         n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060,
         n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070,
         n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080,
         n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090,
         n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100,
         n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110,
         n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120,
         n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130,
         n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140,
         n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150,
         n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160,
         n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170,
         n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180,
         n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190,
         n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200,
         n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210,
         n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220,
         n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230,
         n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240,
         n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250,
         n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260,
         n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270,
         n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280,
         n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290,
         n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300,
         n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310,
         n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320,
         n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330,
         n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340,
         n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350,
         n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360,
         n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370,
         n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380,
         n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390,
         n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400,
         n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410,
         n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420,
         n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430,
         n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440,
         n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450,
         n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460,
         n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470,
         n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480,
         n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490,
         n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500,
         n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510,
         n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520,
         n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530,
         n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540,
         n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550,
         n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560,
         n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570,
         n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580,
         n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590,
         n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600,
         n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610,
         n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620,
         n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630,
         n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640,
         n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650,
         n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660,
         n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670,
         n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680,
         n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690,
         n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700,
         n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710,
         n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720,
         n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730,
         n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740,
         n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750,
         n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760,
         n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770,
         n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780,
         n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790,
         n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800,
         n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810,
         n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820,
         n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830,
         n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840,
         n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850,
         n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860,
         n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870,
         n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880,
         n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890,
         n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900,
         n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910,
         n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920,
         n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930,
         n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940,
         n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950,
         n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960,
         n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970,
         n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980,
         n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990,
         n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
         n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
         n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
         n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
         n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
         n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
         n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280,
         n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288,
         n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296,
         n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304,
         n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
         n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320,
         n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328,
         n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336,
         n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344,
         n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352,
         n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360,
         n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368,
         n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376,
         n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384,
         n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392,
         n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400,
         n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408,
         n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416,
         n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424,
         n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432,
         n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440,
         n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448,
         n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456,
         n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464,
         n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472,
         n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480,
         n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488,
         n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496,
         n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504,
         n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512,
         n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520,
         n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528,
         n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536,
         n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544,
         n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552,
         n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560,
         n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568,
         n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576,
         n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584,
         n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592,
         n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600,
         n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608,
         n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616,
         n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624,
         n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632,
         n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640,
         n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648,
         n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656,
         n10657, n10658, n10659, n10660, n10661, n10662, n10663, n10664,
         n10665, n10666, n10667, n10668, n10669, n10670, n10671, n10672,
         n10673, n10674, n10675, n10676, n10677, n10678, n10679, n10680,
         n10681, n10682, n10683, n10684, n10685, n10686, n10687, n10688,
         n10689, n10690, n10691, n10692, n10693, n10694, n10695, n10696,
         n10697, n10698, n10699, n10700, n10701, n10702, n10703, n10704,
         n10705, n10706, n10707, n10708, n10709, n10710, n10711, n10712,
         n10713, n10714, n10715, n10716, n10717, n10718, n10719, n10720,
         n10721, n10722, n10723, n10724, n10725, n10726, n10727, n10728,
         n10729, n10730, n10731, n10732, n10733, n10734, n10735, n10736,
         n10737, n10738, n10739, n10740, n10741, n10742, n10743, n10744,
         n10745, n10746, n10747, n10748, n10749, n10750, n10751, n10752,
         n10753, n10754, n10755, n10756, n10757, n10758, n10759, n10760,
         n10761, n10762, n10763, n10764, n10765, n10766, n10767, n10768,
         n10769, n10770, n10771, n10772, n10773, n10774, n10775, n10776,
         n10777, n10778, n10779, n10780, n10781, n10782, n10783, n10784,
         n10785, n10786, n10787, n10788, n10789, n10790, n10791, n10792,
         n10793, n10794, n10795, n10796, n10797, n10798, n10799, n10800,
         n10801, n10802, n10803, n10804, n10805, n10806, n10807, n10808,
         n10809, n10810, n10811, n10812, n10813, n10814, n10815, n10816,
         n10817, n10818, n10819, n10820, n10821, n10822, n10823, n10824,
         n10825, n10826, n10827, n10828, n10829, n10830, n10831, n10832,
         n10833, n10834, n10835, n10836, n10837, n10838, n10839, n10840,
         n10841, n10842, n10843, n10844, n10845, n10846, n10847, n10848,
         n10849, n10850, n10851, n10852, n10853, n10854, n10855, n10856,
         n10857, n10858, n10859, n10860, n10861, n10862, n10863, n10864,
         n10865, n10866, n10867, n10868, n10869, n10870, n10871, n10872,
         n10873, n10874, n10875, n10876, n10877, n10878, n10879, n10880,
         n10881, n10882, n10883, n10884, n10885, n10886, n10887, n10888,
         n10889, n10890, n10891, n10892, n10893, n10894, n10895, n10896,
         n10897, n10898, n10899, n10900, n10901, n10902, n10903, n10904,
         n10905, n10906, n10907, n10908, n10909, n10910, n10911, n10912,
         n10913, n10914, n10915, n10916, n10917, n10918, n10919, n10920,
         n10921, n10922, n10923, n10924, n10925, n10926, n10927, n10928,
         n10929, n10930, n10931, n10932, n10933, n10934, n10935, n10936,
         n10937, n10938, n10939, n10940, n10941, n10942, n10943, n10944,
         n10945, n10946, n10947, n10948, n10949, n10950, n10951, n10952,
         n10953, n10954, n10955, n10956, n10957, n10958, n10959, n10960,
         n10961, n10962, n10963, n10964, n10965, n10966, n10967, n10968,
         n10969, n10970, n10971, n10972, n10973, n10974, n10975, n10976,
         n10977, n10978, n10979, n10980, n10981, n10982, n10983, n10984,
         n10985, n10986, n10987, n10988, n10989, n10990, n10991, n10992,
         n10993, n10994, n10995, n10996, n10997, n10998, n10999, n11000,
         n11001, n11002, n11003, n11004, n11005, n11006, n11007, n11008,
         n11009, n11010, n11011, n11012, n11013, n11014, n11015, n11016,
         n11017, n11018, n11019, n11020, n11021, n11022, n11023, n11024,
         n11025, n11026, n11027, n11028, n11029, n11030, n11031, n11032,
         n11033, n11034, n11035, n11036, n11037, n11038, n11039, n11040,
         n11041, n11042, n11043, n11044, n11045, n11046, n11047, n11048,
         n11049, n11050, n11051, n11052, n11053, n11054, n11055, n11056,
         n11057, n11058, n11059, n11060, n11061, n11062, n11063, n11064,
         n11065, n11066, n11067, n11068, n11069, n11070, n11071, n11072,
         n11073, n11074, n11075, n11076, n11077, n11078, n11079, n11080,
         n11081, n11082, n11083, n11084, n11085, n11086, n11087, n11088,
         n11089, n11090, n11091, n11092, n11093, n11094, n11095, n11096,
         n11097, n11098, n11099, n11100, n11101, n11102, n11103, n11104,
         n11105, n11106, n11107, n11108, n11109, n11110, n11111, n11112,
         n11113, n11114, n11115, n11116, n11117, n11118, n11119, n11120,
         n11121, n11122, n11123, n11124, n11125, n11126, n11127, n11128,
         n11129, n11130, n11131, n11132, n11133, n11134, n11135, n11136,
         n11137, n11138, n11139, n11140, n11141, n11142, n11143, n11144,
         n11145, n11146, n11147, n11148, n11149, n11150, n11151, n11152,
         n11153, n11154, n11155, n11156, n11157, n11158, n11159, n11160,
         n11161, n11162, n11163, n11164, n11165, n11166, n11167, n11168,
         n11169, n11170, n11171, n11172, n11173, n11174, n11175, n11176,
         n11177, n11178, n11179, n11180, n11181, n11182, n11183, n11184,
         n11185, n11186, n11187, n11188, n11189, n11190, n11191, n11192,
         n11193, n11194, n11195, n11196, n11197, n11198, n11199, n11200,
         n11201, n11202, n11203, n11204, n11205, n11206, n11207, n11208,
         n11209, n11210, n11211, n11212, n11213, n11214, n11215, n11216,
         n11217, n11218, n11219, n11220, n11221, n11222, n11223, n11224,
         n11225, n11226, n11227, n11228, n11229, n11230, n11231, n11232,
         n11233, n11234, n11235, n11236, n11237, n11238, n11239, n11240,
         n11241, n11242, n11243, n11244, n11245, n11246, n11247, n11248,
         n11249, n11250, n11251, n11252, n11253, n11254, n11255, n11256,
         n11257, n11258, n11259, n11260, n11261, n11262, n11263, n11264,
         n11265, n11266, n11267, n11268, n11269, n11270, n11271, n11272,
         n11273, n11274, n11275, n11276, n11277, n11278, n11279, n11280,
         n11281, n11282, n11283, n11284, n11285, n11286, n11287, n11288,
         n11289, n11290, n11291, n11292, n11293, n11294, n11295, n11296,
         n11297, n11298, n11299, n11300, n11301, n11302, n11303, n11304,
         n11305, n11306, n11307, n11308, n11309, n11310, n11311, n11312,
         n11313, n11314, n11315, n11316, n11317, n11318, n11319, n11320,
         n11321, n11322, n11323, n11324, n11325, n11326, n11327, n11328,
         n11329, n11330, n11331, n11332, n11333, n11334, n11335, n11336,
         n11337, n11338, n11339, n11340, n11341, n11342, n11343, n11344,
         n11345, n11346, n11347, n11348, n11349, n11350, n11351, n11352,
         n11353, n11354, n11355, n11356, n11357, n11358, n11359, n11360,
         n11361, n11362, n11363, n11364, n11365, n11366, n11367, n11368,
         n11369, n11370, n11371, n11372, n11373, n11374, n11375, n11376,
         n11377, n11378, n11379, n11380, n11381, n11382, n11383, n11384,
         n11385, n11386, n11387, n11388, n11389, n11390, n11391, n11392,
         n11393, n11394, n11395, n11396, n11397, n11398, n11399, n11400,
         n11401, n11402, n11403, n11404, n11405, n11406, n11407, n11408,
         n11409, n11410, n11411, n11412, n11413, n11414, n11415, n11416,
         n11417, n11418, n11419, n11420, n11421, n11422, n11423, n11424,
         n11425, n11426, n11427, n11428, n11429, n11430, n11431, n11432,
         n11433, n11434, n11435, n11436, n11437, n11438, n11439, n11440,
         n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448,
         n11449, n11450, n11451, n11452, n11453, n11454, n11455, n11456,
         n11457, n11458, n11459, n11460, n11461, n11462, n11463, n11464,
         n11465, n11466, n11467, n11468, n11469, n11470, n11471, n11472,
         n11473, n11474, n11475, n11476, n11477, n11478, n11479, n11480,
         n11481, n11482, n11483, n11484, n11485, n11486, n11487, n11488,
         n11489, n11490, n11491, n11492, n11493, n11494, n11495, n11496,
         n11497, n11498, n11499, n11500, n11501, n11502, n11503, n11504,
         n11505, n11506, n11507, n11508, n11509, n11510, n11511, n11512,
         n11513, n11514, n11515, n11516, n11517, n11518, n11519, n11520,
         n11521, n11522, n11523, n11524, n11525, n11526, n11527, n11528,
         n11529, n11530, n11531, n11532, n11533, n11534, n11535, n11536,
         n11537, n11538, n11539, n11540, n11541, n11542, n11543, n11544,
         n11545, n11546, n11547, n11548, n11549, n11550, n11551, n11552,
         n11553, n11554, n11555, n11556, n11557, n11558, n11559, n11560,
         n11561, n11562, n11563, n11564, n11565, n11566, n11567, n11568,
         n11569, n11570, n11571, n11572, n11573, n11574, n11575, n11576,
         n11577, n11578, n11579, n11580, n11581, n11582, n11583, n11584,
         n11585, n11586, n11587, n11588, n11589, n11590, n11591, n11592,
         n11593, n11594, n11595, n11596, n11597, n11598, n11599, n11600,
         n11601, n11602, n11603, n11604, n11605, n11606, n11607, n11608,
         n11609, n11610, n11611, n11612, n11613, n11614, n11615, n11616,
         n11617, n11618, n11619, n11620, n11621, n11622, n11623, n11624,
         n11625, n11626, n11627, n11628, n11629, n11630, n11631, n11632,
         n11633, n11634, n11635, n11636, n11637, n11638, n11639, n11640,
         n11641, n11642, n11643, n11644, n11645, n11646, n11647, n11648,
         n11649, n11650, n11651, n11652, n11653, n11654, n11655, n11656,
         n11657, n11658, n11659, n11660, n11661, n11662, n11663, n11664,
         n11665, n11666, n11667, n11668, n11669, n11670, n11671, n11672,
         n11673, n11674, n11675, n11676, n11677, n11678, n11679, n11680,
         n11681, n11682, n11683, n11684, n11685, n11686, n11687, n11688,
         n11689, n11690, n11691, n11692, n11693, n11694, n11695, n11696,
         n11697, n11698, n11699, n11700, n11701, n11702, n11703, n11704,
         n11705, n11706, n11707, n11708, n11709, n11710, n11711, n11712,
         n11713, n11714, n11715, n11716, n11717, n11718, n11719, n11720,
         n11721, n11722, n11723, n11724, n11725, n11726, n11727, n11728,
         n11729, n11730, n11731, n11732, n11733, n11734, n11735, n11736,
         n11737, n11738, n11739, n11740, n11741, n11742, n11743, n11744,
         n11745, n11746, n11747, n11748, n11749, n11750, n11751, n11752,
         n11753, n11754, n11755, n11756, n11757, n11758, n11759, n11760,
         n11761, n11762, n11763, n11764, n11765, n11766, n11767, n11768,
         n11769, n11770, n11771, n11772, n11773, n11774, n11775, n11776,
         n11777, n11778, n11779, n11780, n11781, n11782, n11783, n11784,
         n11785, n11786, n11787, n11788, n11789, n11790, n11791, n11792,
         n11793, n11794, n11795, n11796, n11797, n11798, n11799, n11800,
         n11801, n11802, n11803, n11804, n11805, n11806, n11807, n11808,
         n11809, n11810, n11811, n11812, n11813, n11814, n11815, n11816,
         n11817, n11818, n11819, n11820, n11821, n11822, n11823, n11824,
         n11825, n11826, n11827, n11828, n11829, n11830, n11831, n11832,
         n11833, n11834, n11835, n11836, n11837, n11838, n11839, n11840,
         n11841, n11842, n11843, n11844, n11845, n11846, n11847, n11848,
         n11849, n11850, n11851, n11852, n11853, n11854, n11855, n11856,
         n11857, n11858, n11859, n11860, n11861, n11862, n11863, n11864,
         n11865, n11866, n11867, n11868, n11869, n11870, n11871, n11872,
         n11873, n11874, n11875, n11876, n11877, n11878, n11879, n11880,
         n11881, n11882, n11883, n11884, n11885, n11886, n11887, n11888,
         n11889, n11890, n11891, n11892, n11893, n11894, n11895, n11896,
         n11897, n11898, n11899, n11900, n11901, n11902, n11903, n11904,
         n11905, n11906, n11907, n11908, n11909, n11910, n11911, n11912,
         n11913, n11914, n11915, n11916, n11917, n11918, n11919, n11920,
         n11921, n11922, n11923, n11924, n11925, n11926, n11927, n11928,
         n11929, n11930, n11931, n11932, n11933, n11934, n11935, n11936,
         n11937, n11938, n11939, n11940, n11941, n11942, n11943, n11944,
         n11945, n11946, n11947, n11948, n11949, n11950, n11951, n11952,
         n11953, n11954, n11955, n11956, n11957, n11958, n11959, n11960,
         n11961, n11962, n11963, n11964, n11965, n11966, n11967, n11968,
         n11969, n11970, n11971, n11972, n11973, n11974, n11975, n11976,
         n11977, n11978, n11979, n11980, n11981, n11982, n11983, n11984,
         n11985, n11986, n11987, n11988, n11989, n11990, n11991, n11992,
         n11993, n11994, n11995, n11996, n11997, n11998, n11999, n12000,
         n12001, n12002, n12003, n12004, n12005, n12006, n12007, n12008,
         n12009, n12010, n12011, n12012, n12013, n12014, n12015, n12016,
         n12017, n12018, n12019, n12020, n12021, n12022, n12023, n12024,
         n12025, n12026, n12027, n12028, n12029, n12030, n12031, n12032,
         n12033, n12034, n12035, n12036, n12037, n12038, n12039, n12040,
         n12041, n12042, n12043, n12044, n12045, n12046, n12047, n12048,
         n12049, n12050, n12051, n12052, n12053, n12054, n12055, n12056,
         n12057, n12058, n12059, n12060, n12061, n12062, n12063, n12064,
         n12065, n12066, n12067, n12068, n12069, n12070, n12071, n12072,
         n12073, n12074, n12075, n12076, n12077, n12078, n12079, n12080,
         n12081, n12082, n12083, n12084, n12085, n12086, n12087, n12088,
         n12089, n12090, n12091, n12092, n12093, n12094, n12095, n12096,
         n12097, n12098, n12099, n12100, n12101, n12102, n12103, n12104,
         n12105, n12106, n12107, n12108, n12109, n12110, n12111, n12112,
         n12113, n12114, n12115, n12116, n12117, n12118, n12119, n12120,
         n12121, n12122, n12123, n12124, n12125, n12126, n12127, n12128,
         n12129, n12130, n12131, n12132, n12133, n12134, n12135, n12136,
         n12137, n12138, n12139, n12140, n12141, n12142, n12143, n12144,
         n12145, n12146, n12147, n12148, n12149, n12150, n12151, n12152,
         n12153, n12154, n12155, n12156, n12157, n12158, n12159, n12160,
         n12161, n12162, n12163, n12164, n12165, n12166, n12167, n12168,
         n12169, n12170, n12171, n12172, n12173, n12174, n12175, n12176,
         n12177, n12178, n12179, n12180, n12181, n12182, n12183, n12184,
         n12185, n12186, n12187, n12188, n12189, n12190, n12191, n12192,
         n12193, n12194, n12195, n12196, n12197, n12198, n12199, n12200,
         n12201, n12202, n12203, n12204, n12205, n12206, n12207, n12208,
         n12209, n12210, n12211, n12212, n12213, n12214, n12215, n12216,
         n12217, n12218, n12219, n12220, n12221, n12222, n12223, n12224,
         n12225, n12226, n12227, n12228, n12229, n12230, n12231, n12232,
         n12233, n12234, n12235, n12236, n12237, n12238, n12239, n12240,
         n12241, n12242, n12243, n12244, n12245, n12246, n12247, n12248,
         n12249, n12250, n12251, n12252, n12253, n12254, n12255, n12256,
         n12257, n12258, n12259, n12260, n12261, n12262, n12263, n12264,
         n12265, n12266, n12267, n12268, n12269, n12270, n12271, n12272,
         n12273, n12274, n12275, n12276, n12277, n12278, n12279, n12280,
         n12281, n12282, n12283, n12284, n12285, n12286, n12287, n12288,
         n12289, n12290, n12291, n12292, n12293, n12294, n12295, n12296,
         n12297, n12298, n12299, n12300, n12301, n12302, n12303, n12304,
         n12305, n12306, n12307, n12308, n12309, n12310, n12311, n12312,
         n12313, n12314, n12315, n12316, n12317, n12318, n12319, n12320,
         n12321, n12322, n12323, n12324, n12325, n12326, n12327, n12328,
         n12329, n12330, n12331, n12332, n12333, n12334, n12335, n12336,
         n12337, n12338, n12339, n12340, n12341, n12342, n12343, n12344,
         n12345, n12346, n12347, n12348, n12349, n12350, n12351, n12352,
         n12353, n12354, n12355, n12356, n12357, n12358, n12359, n12360,
         n12361, n12362, n12363, n12364, n12365, n12366, n12367, n12368,
         n12369, n12370, n12371, n12372, n12373, n12374, n12375, n12376,
         n12377, n12378, n12379, n12380, n12381, n12382, n12383, n12384,
         n12385, n12386, n12387, n12388, n12389, n12390, n12391, n12392,
         n12393, n12394, n12395, n12396, n12397, n12398, n12399, n12400,
         n12401, n12402, n12403, n12404, n12405, n12406, n12407, n12408,
         n12409, n12410, n12411, n12412, n12413, n12414, n12415, n12416,
         n12417, n12418, n12419, n12420, n12421, n12422, n12423, n12424,
         n12425, n12426, n12427, n12428, n12429, n12430, n12431, n12432,
         n12433, n12434, n12435, n12436, n12437, n12438, n12439, n12440,
         n12441, n12442, n12443, n12444, n12445, n12446, n12447, n12448,
         n12449, n12450, n12451, n12452, n12453, n12454, n12455, n12456,
         n12457, n12458, n12459, n12460, n12461, n12462, n12463, n12464,
         n12465, n12466, n12467, n12468, n12469, n12470, n12471, n12472,
         n12473, n12474, n12475, n12476, n12477, n12478, n12479, n12480,
         n12481, n12482, n12483, n12484, n12485, n12486, n12487, n12488,
         n12489, n12490, n12491, n12492, n12493, n12494, n12495, n12496,
         n12497, n12498, n12499, n12500, n12501, n12502, n12503, n12504,
         n12505, n12506, n12507, n12508, n12509, n12510, n12511, n12512,
         n12513, n12514, n12515, n12516, n12517, n12518, n12519, n12520,
         n12521, n12522, n12523, n12524, n12525, n12526, n12527, n12528,
         n12529, n12530, n12531, n12532, n12533, n12534, n12535, n12536,
         n12537, n12538, n12539, n12540, n12541, n12542, n12543, n12544,
         n12545, n12546, n12547, n12548, n12549, n12550, n12551, n12552,
         n12553, n12554, n12555, n12556, n12557, n12558, n12559, n12560,
         n12561, n12562, n12563, n12564, n12565, n12566, n12567, n12568,
         n12569, n12570, n12571, n12572, n12573, n12574, n12575, n12576,
         n12577, n12578, n12579, n12580, n12581, n12582, n12583, n12584,
         n12585, n12586, n12587, n12588, n12589, n12590, n12591, n12592,
         n12593, n12594, n12595, n12596, n12597, n12598, n12599, n12600,
         n12601, n12602, n12603, n12604, n12605, n12606, n12607, n12608,
         n12609, n12610, n12611, n12612, n12613, n12614, n12615, n12616,
         n12617, n12618, n12619, n12620, n12621, n12622, n12623, n12624,
         n12625, n12626, n12627, n12628, n12629, n12630, n12631, n12632,
         n12633, n12634, n12635, n12636, n12637, n12638, n12639, n12640,
         n12641, n12642, n12643, n12644, n12645, n12646, n12647, n12648,
         n12649, n12650, n12651, n12652, n12653, n12654, n12655, n12656,
         n12657, n12658, n12659, n12660, n12661, n12662, n12663, n12664,
         n12665, n12666, n12667, n12668, n12669, n12670, n12671, n12672,
         n12673, n12674, n12675, n12676, n12677, n12678, n12679, n12680,
         n12681, n12682, n12683, n12684, n12685, n12686, n12687, n12688,
         n12689, n12690, n12691, n12692, n12693, n12694, n12695, n12696,
         n12697, n12698, n12699, n12700, n12701, n12702, n12703, n12704,
         n12705, n12706, n12707, n12708, n12709, n12710, n12711, n12712,
         n12713, n12714, n12715, n12716, n12717, n12718, n12719, n12720,
         n12721, n12722, n12723, n12724, n12725, n12726, n12727, n12728,
         n12729, n12730, n12731, n12732, n12733, n12734, n12735, n12736,
         n12737, n12738, n12739, n12740, n12741, n12742, n12743, n12744,
         n12745, n12746, n12747, n12748, n12749, n12750, n12751, n12752,
         n12753, n12754, n12755, n12756, n12757, n12758, n12759, n12760,
         n12761, n12762, n12763, n12764, n12765, n12766, n12767, n12768,
         n12769, n12770, n12771, n12772, n12773, n12774, n12775, n12776,
         n12777, n12778, n12779, n12780, n12781, n12782, n12783, n12784,
         n12785, n12786, n12787, n12788, n12789, n12790, n12791, n12792,
         n12793, n12794, n12795, n12796, n12797, n12798, n12799, n12800,
         n12801, n12802, n12803, n12804, n12805, n12806, n12807, n12808,
         n12809, n12810, n12811, n12812, n12813, n12814, n12815, n12816,
         n12817, n12818, n12819, n12820, n12821, n12822, n12823, n12824,
         n12825, n12826, n12827, n12828, n12829, n12830, n12831, n12832,
         n12833, n12834, n12835, n12836, n12837, n12838, n12839, n12840,
         n12841, n12842, n12843, n12844, n12845, n12846, n12847, n12848,
         n12849, n12850, n12851, n12852, n12853, n12854, n12855, n12856,
         n12857, n12858, n12859, n12860, n12861, n12862, n12863, n12864,
         n12865, n12866, n12867, n12868, n12869, n12870, n12871, n12872,
         n12873, n12874, n12875, n12876, n12877, n12878, n12879, n12880,
         n12881, n12882, n12883, n12884, n12885, n12886, n12887, n12888,
         n12889, n12890, n12891, n12892, n12893, n12894, n12895, n12896,
         n12897, n12898, n12899, n12900, n12901, n12902, n12903, n12904,
         n12905, n12906, n12907, n12908, n12909, n12910, n12911, n12912,
         n12913, n12914, n12915, n12916, n12917, n12918, n12919, n12920,
         n12921, n12922, n12923, n12924, n12925, n12926, n12927, n12928,
         n12929, n12930, n12931, n12932, n12933, n12934, n12935, n12936,
         n12937, n12938, n12939, n12940, n12941, n12942, n12943, n12944,
         n12945, n12946, n12947, n12948, n12949, n12950, n12951, n12952,
         n12953, n12954, n12955, n12956, n12957, n12958, n12959, n12960,
         n12961, n12962, n12963, n12964, n12965, n12966, n12967, n12968,
         n12969, n12970, n12971, n12972, n12973, n12974, n12975, n12976,
         n12977, n12978, n12979, n12980, n12981, n12982, n12983, n12984,
         n12985, n12986, n12987, n12988, n12989, n12990, n12991, n12992,
         n12993, n12994, n12995, n12996, n12997, n12998, n12999, n13000,
         n13001, n13002, n13003, n13004, n13005, n13006, n13007, n13008,
         n13009, n13010, n13011, n13012, n13013, n13014, n13015, n13016,
         n13017, n13018, n13019, n13020, n13021, n13022, n13023, n13024,
         n13025, n13026, n13027, n13028, n13029, n13030, n13031, n13032,
         n13033, n13034, n13035, n13036, n13037, n13038, n13039, n13040,
         n13041, n13042, n13043, n13044, n13045, n13046, n13047, n13048,
         n13049, n13050, n13051, n13052, n13053, n13054, n13055, n13056,
         n13057, n13058, n13059, n13060, n13061, n13062, n13063, n13064,
         n13065, n13066, n13067, n13068, n13069, n13070, n13071, n13072,
         n13073, n13074, n13075, n13076, n13077, n13078, n13079, n13080,
         n13081, n13082, n13083, n13084, n13085, n13086, n13087, n13088,
         n13089, n13090, n13091, n13092, n13093, n13094, n13095, n13096,
         n13097, n13098, n13099, n13100, n13101, n13102, n13103, n13104,
         n13105, n13106, n13107, n13108, n13109, n13110, n13111, n13112,
         n13113, n13114, n13115, n13116, n13117, n13118, n13119, n13120,
         n13121, n13122, n13123, n13124, n13125, n13126, n13127, n13128,
         n13129, n13130, n13131, n13132, n13133, n13134, n13135, n13136,
         n13137, n13138, n13139, n13140, n13141, n13142, n13143, n13144,
         n13145, n13146, n13147, n13148, n13149, n13150, n13151, n13152,
         n13153, n13154, n13155, n13156, n13157, n13158, n13159, n13160,
         n13161, n13162, n13163, n13164, n13165, n13166, n13167, n13168,
         n13169, n13170, n13171, n13172, n13173, n13174, n13175, n13176,
         n13177, n13178, n13179, n13180, n13181, n13182, n13183, n13184,
         n13185, n13186, n13187, n13188, n13189, n13190, n13191, n13192,
         n13193, n13194, n13195, n13196, n13197, n13198, n13199, n13200,
         n13201, n13202, n13203, n13204, n13205, n13206, n13207, n13208,
         n13209, n13210, n13211, n13212, n13213, n13214, n13215, n13216,
         n13217, n13218, n13219, n13220, n13221, n13222, n13223, n13224,
         n13225, n13226, n13227, n13228, n13229, n13230, n13231, n13232,
         n13233, n13234, n13235, n13236, n13237, n13238, n13239, n13240,
         n13241, n13242, n13243, n13244, n13245, n13246, n13247, n13248,
         n13249, n13250, n13251, n13252, n13253, n13254, n13255, n13256,
         n13257, n13258, n13259, n13260, n13261, n13262, n13263, n13264,
         n13265, n13266, n13267, n13268, n13269, n13270, n13271, n13272,
         n13273, n13274, n13275, n13276, n13277, n13278, n13279, n13280,
         n13281, n13282, n13283, n13284, n13285, n13286, n13287, n13288,
         n13289, n13290, n13291, n13292, n13293, n13294, n13295, n13296,
         n13297, n13298, n13299, n13300, n13301, n13302, n13303, n13304,
         n13305, n13306, n13307, n13308, n13309, n13310, n13311, n13312,
         n13313, n13314, n13315, n13316, n13317, n13318, n13319, n13320,
         n13321, n13322, n13323, n13324, n13325, n13326, n13327, n13328,
         n13329, n13330, n13331, n13332, n13333, n13334, n13335, n13336,
         n13337, n13338, n13339, n13340, n13341, n13342, n13343, n13344,
         n13345, n13346, n13347, n13348, n13349, n13350, n13351, n13352,
         n13353, n13354, n13355, n13356, n13357, n13358, n13359, n13360,
         n13361, n13362, n13363, n13364, n13365, n13366, n13367, n13368,
         n13369, n13370, n13371, n13372, n13373, n13374, n13375, n13376,
         n13377, n13378, n13379, n13380, n13381, n13382, n13383, n13384,
         n13385, n13386, n13387, n13388, n13389, n13390, n13391, n13392,
         n13393, n13394, n13395, n13396, n13397, n13398, n13399, n13400,
         n13401, n13402, n13403, n13404, n13405, n13406, n13407, n13408,
         n13409, n13410, n13411, n13412, n13413, n13414, n13415, n13416,
         n13417, n13418, n13419, n13420, n13421, n13422, n13423, n13424,
         n13425, n13426, n13427, n13428, n13429, n13430, n13431, n13432,
         n13433, n13434, n13435, n13436, n13437, n13438, n13439, n13440,
         n13441, n13442, n13443, n13444, n13445, n13446, n13447, n13448,
         n13449, n13450, n13451, n13452, n13453, n13454, n13455, n13456,
         n13457, n13458, n13459, n13460, n13461, n13462, n13463, n13464,
         n13465, n13466, n13467, n13468, n13469, n13470, n13471, n13472,
         n13473, n13474, n13475, n13476, n13477, n13478, n13479, n13480,
         n13481, n13482, n13483, n13484, n13485, n13486, n13487, n13488,
         n13489, n13490, n13491, n13492, n13493, n13494, n13495, n13496,
         n13497, n13498, n13499, n13500, n13501, n13502, n13503, n13504,
         n13505, n13506, n13507, n13508, n13509, n13510, n13511, n13512,
         n13513, n13514, n13515, n13516, n13517, n13518, n13519, n13520,
         n13521, n13522, n13523, n13524, n13525, n13526, n13527, n13528,
         n13529, n13530, n13531, n13532, n13533, n13534, n13535, n13536,
         n13537, n13538, n13539, n13540, n13541, n13542, n13543, n13544,
         n13545, n13546, n13547, n13548, n13549, n13550, n13551, n13552,
         n13553, n13554, n13555, n13556, n13557, n13558, n13559, n13560,
         n13561, n13562, n13563, n13564, n13565, n13566, n13567, n13568,
         n13569, n13570, n13571, n13572, n13573, n13574, n13575, n13576,
         n13577, n13578, n13579, n13580, n13581, n13582, n13583, n13584,
         n13585, n13586, n13587, n13588, n13589, n13590, n13591, n13592,
         n13593, n13594, n13595, n13596, n13597, n13599, n13600, n13601,
         n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609,
         n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617,
         n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625,
         n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633,
         n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641,
         n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649,
         n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657,
         n13658, n13659, n13660, n13661, n13662, n13663, n13664, n13665,
         n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673,
         n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681,
         n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689,
         n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697,
         n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705,
         n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713,
         n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721,
         n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729,
         n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737,
         n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745,
         n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753,
         n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761,
         n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769,
         n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777,
         n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785,
         n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793,
         n13794, n13795, n13796, n13797, n13798, n13799, n13800, n13801,
         n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809,
         n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817,
         n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825,
         n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833,
         n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841,
         n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849,
         n13850, n13851, n13852, n13853, n13854, n13855, n13856, n13857,
         n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865,
         n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873,
         n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881,
         n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889,
         n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897,
         n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905,
         n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913,
         n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921,
         n13922, n13923, n13924, n13925, n13926, n13927, n13928, n13929,
         n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937,
         n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945,
         n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953,
         n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961,
         n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969,
         n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977,
         n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985,
         n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993,
         n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001,
         n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009,
         n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017,
         n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025,
         n14026, n14027, n14028, n14029, n14030, n14031, n14032, n14033,
         n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041,
         n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049,
         n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057,
         n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065,
         n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073,
         n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081,
         n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089,
         n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097,
         n14098, n14099, n14100, n14101, n14102, n14103, n14104, n14105,
         n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113,
         n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121,
         n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129,
         n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137,
         n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145,
         n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153,
         n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161,
         n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169,
         n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177,
         n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185,
         n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193,
         n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201,
         n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209,
         n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217,
         n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225,
         n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233,
         n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241,
         n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249,
         n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257,
         n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265,
         n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273,
         n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281,
         n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289,
         n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297,
         n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305,
         n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313,
         n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321,
         n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329,
         n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337,
         n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345,
         n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353,
         n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361,
         n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369,
         n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377,
         n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385,
         n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393,
         n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401,
         n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409,
         n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417,
         n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425,
         n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433,
         n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441,
         n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449,
         n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457,
         n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465,
         n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473,
         n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481,
         n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489,
         n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497,
         n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505,
         n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513,
         n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521,
         n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529,
         n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537,
         n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545,
         n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553,
         n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561,
         n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569,
         n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577,
         n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585,
         n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593,
         n14594, n14595, n14596, n14597, n14598, n14599, n14600, n14601,
         n14602, n14603, n14604, n14605, n14606, n14607, n14608, n14609,
         n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617,
         n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625,
         n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633,
         n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641,
         n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649,
         n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657,
         n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665,
         n14666, n14667, n14668, n14669, n14670, n14671, n14672, n14673,
         n14674, n14675, n14676, n14677, n14678, n14679, n14680, n14681,
         n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689,
         n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697,
         n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705,
         n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713,
         n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721,
         n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729,
         n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737,
         n14738, n14739, n14740, n14741, n14742, n14743, n14744, n14745,
         n14746, n14747, n14748, n14749, n14750, n14751, n14752, n14753,
         n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761,
         n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769,
         n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777,
         n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785,
         n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793,
         n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801,
         n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809,
         n14810, n14811, n14812, n14813, n14814, n14815, n14816, n14817,
         n14818, n14819, n14820, n14821, n14822, n14823, n14824, n14825,
         n14826, n14827, n14828, n14829, n14830, n14831, n14832, n14833,
         n14834, n14835, n14836, n14837, n14838, n14839, n14840, n14841,
         n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849,
         n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857,
         n14858, n14859, n14860, n14861, n14862, n14863, n14864, n14865,
         n14866, n14867, n14868, n14869, n14870, n14871, n14872, n14873,
         n14874, n14875, n14876, n14877, n14878, n14879, n14880, n14881,
         n14882, n14883, n14884, n14885, n14886, n14887, n14888, n14889,
         n14890, n14891, n14892, n14893, n14894, n14895, n14896, n14897,
         n14898, n14899, n14900, n14901, n14902, n14903, n14904, n14905,
         n14906, n14907, n14908, n14909, n14910, n14911, n14912, n14913,
         n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921,
         n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929,
         n14930, n14931, n14932, n14933, n14934, n14935, n14936, n14937,
         n14938, n14939, n14940, n14941, n14942, n14943, n14944, n14945,
         n14946, n14947, n14948, n14949, n14950, n14951, n14952, n14953,
         n14954, n14955, n14956, n14957, n14958, n14959, n14960, n14961,
         n14962, n14963, n14964, n14965, n14966, n14967, n14968, n14969,
         n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14977,
         n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985,
         n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993,
         n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001,
         n15002, n15003, n15004, n15005, n15006, n15007, n15008, n15009,
         n15010, n15011, n15012, n15013, n15014, n15015, n15016, n15017,
         n15018, n15019, n15020, n15021, n15022, n15023, n15024, n15025,
         n15026, n15027, n15028, n15029, n15030, n15031, n15032, n15033,
         n15034, n15035, n15036, n15037, n15038, n15039, n15040, n15041,
         n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049,
         n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057,
         n15058, n15059, n15060, n15061, n15062, n15063, n15064, n15065,
         n15066, n15067, n15068, n15069, n15070, n15071, n15072, n15073,
         n15074, n15075, n15076, n15077, n15078, n15079, n15080, n15081,
         n15082, n15083, n15084, n15085, n15086, n15087, n15088, n15089,
         n15090, n15091, n15092, n15093, n15094, n15095, n15096, n15097,
         n15098, n15099, n15100, n15101, n15102, n15103, n15104, n15105,
         n15106, n15107, n15108, n15109, n15110, n15111, n15112, n15113,
         n15114, n15115, n15116, n15117, n15118, n15119, n15120, n15121,
         n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129,
         n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137,
         n15138, n15139, n15140, n15141, n15142, n15143, n15144, n15145,
         n15146, n15147, n15148, n15149, n15150, n15151, n15152, n15153,
         n15154, n15155, n15156, n15157, n15158, n15159, n15160, n15161,
         n15162, n15163, n15164, n15165, n15166, n15167, n15168, n15169,
         n15170, n15171, n15172, n15173, n15174, n15175, n15176, n15177,
         n15178, n15179, n15180, n15181, n15182, n15183, n15184, n15185,
         n15186, n15187, n15188, n15189, n15190, n15191, n15192, n15193,
         n15194, n15195, n15196, n15197, n15198, n15199, n15200, n15201,
         n15202, n15203, n15204, n15205, n15206, n15207, n15208, n15209,
         n15210, n15211, n15212, n15213, n15214, n15215, n15216, n15217,
         n15218, n15219, n15220, n15221, n15222, n15223, n15224, n15225,
         n15226, n15227, n15228, n15229, n15230, n15231, n15232, n15233,
         n15234, n15235, n15236, n15237, n15238, n15239, n15240, n15241,
         n15242, n15243, n15244, n15245, n15246, n15247, n15248, n15249,
         n15250, n15251, n15252, n15253, n15254, n15255, n15256, n15257,
         n15258, n15259, n15260, n15261, n15262, n15263, n15264, n15265,
         n15266, n15267, n15268, n15269, n15270, n15271, n15272, n15273,
         n15274, n15275, n15276, n15277, n15278, n15279, n15280, n15281,
         n15282, n15283, n15284, n15285, n15286, n15287, n15288, n15289,
         n15290, n15291, n15292, n15293, n15294, n15295, n15296, n15297,
         n15298, n15299, n15300, n15301, n15302, n15303, n15304, n15305,
         n15306, n15307, n15308, n15309, n15310, n15311, n15312, n15313,
         n15314, n15315, n15316, n15317, n15318, n15319, n15320, n15321,
         n15322, n15323, n15324, n15325, n15326, n15327, n15328, n15329,
         n15330, n15331, n15332, n15333, n15334, n15335, n15336, n15337,
         n15338, n15339, n15340, n15341, n15342, n15343, n15344, n15345,
         n15346, n15347, n15348, n15349, n15350, n15351, n15352, n15353,
         n15354, n15355, n15356, n15357, n15358, n15359, n15360, n15361,
         n15362, n15363, n15364, n15365, n15366, n15367, n15368, n15369,
         n15370, n15371, n15372, n15373, n15374, n15375, n15376, n15377,
         n15378, n15379, n15380, n15381, n15382, n15383, n15384, n15385,
         n15386, n15387, n15388, n15389, n15390, n15391, n15392, n15393,
         n15394, n15395, n15396, n15397, n15398, n15399, n15400, n15401,
         n15402, n15403, n15404, n15405, n15406, n15407, n15408, n15409,
         n15410, n15411, n15412, n15413, n15414, n15415, n15416, n15417,
         n15418, n15419, n15420, n15421, n15422, n15423, n15424, n15425,
         n15426, n15427, n15428, n15429, n15430, n15431, n15432, n15433,
         n15434, n15435, n15436, n15437;

  AND2_X1 U7264 ( .A1(n6976), .A2(n6975), .ZN(n8556) );
  INV_X1 U7265 ( .A(n6516), .ZN(n13992) );
  OR2_X1 U7266 ( .A1(n11870), .A2(n6941), .ZN(n6940) );
  NAND2_X1 U7267 ( .A1(n8139), .A2(n8138), .ZN(n13277) );
  NAND2_X1 U7268 ( .A1(n8482), .A2(n8481), .ZN(n8505) );
  AOI21_X1 U7269 ( .B1(n12793), .B2(n11809), .A(n7605), .ZN(n12781) );
  OAI22_X1 U7270 ( .A1(n12861), .A2(n11802), .B1(n12851), .B2(n12918), .ZN(
        n12850) );
  NOR2_X2 U7271 ( .A1(n10550), .A2(n10779), .ZN(n7403) );
  NAND2_X1 U7272 ( .A1(n13700), .A2(n13699), .ZN(n11662) );
  XNOR2_X1 U7273 ( .A(n6832), .B(n8100), .ZN(n11573) );
  NAND2_X1 U7274 ( .A1(n8098), .A2(n8097), .ZN(n6832) );
  OR2_X1 U7275 ( .A1(n14665), .A2(n14664), .ZN(n14666) );
  NAND2_X1 U7276 ( .A1(n8914), .A2(n8913), .ZN(n8936) );
  CLKBUF_X2 U7277 ( .A(n12087), .Z(n6529) );
  INV_X1 U7278 ( .A(n12003), .ZN(n7134) );
  INV_X1 U7279 ( .A(n9197), .ZN(n9271) );
  NAND4_X2 U7280 ( .A1(n8739), .A2(n8738), .A3(n8737), .A4(n8736), .ZN(n15054)
         );
  NAND4_X2 U7282 ( .A1(n8727), .A2(n8726), .A3(n8725), .A4(n8724), .ZN(n12557)
         );
  BUF_X2 U7283 ( .A(n8973), .Z(n6542) );
  AND2_X1 U7285 ( .A1(n8603), .A2(n11466), .ZN(n8698) );
  NAND2_X2 U7286 ( .A1(n9116), .A2(n9721), .ZN(n9724) );
  INV_X1 U7287 ( .A(n8302), .ZN(n8348) );
  AND2_X2 U7288 ( .A1(n9181), .A2(n9185), .ZN(n11428) );
  NAND4_X2 U7289 ( .A1(n9329), .A2(n9328), .A3(n9327), .A4(n9326), .ZN(n13776)
         );
  NAND2_X1 U7290 ( .A1(n8653), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8655) );
  XNOR2_X1 U7291 ( .A(n8601), .B(P3_IR_REG_30__SCAN_IN), .ZN(n8603) );
  CLKBUF_X1 U7292 ( .A(n9734), .Z(n6532) );
  CLKBUF_X2 U7293 ( .A(n8549), .Z(n6527) );
  INV_X1 U7294 ( .A(n8162), .ZN(n7769) );
  NAND2_X1 U7295 ( .A1(n11572), .A2(n9473), .ZN(n9402) );
  NAND2_X1 U7296 ( .A1(n9366), .A2(n9365), .ZN(n9652) );
  AND2_X1 U7297 ( .A1(n8227), .A2(n8549), .ZN(n8553) );
  OR2_X1 U7298 ( .A1(n7730), .A2(n7728), .ZN(n7408) );
  OAI21_X1 U7299 ( .B1(n9187), .B2(n7540), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n9339) );
  INV_X2 U7300 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n7728) );
  NOR2_X2 U7301 ( .A1(n13848), .A2(n13849), .ZN(n13855) );
  NOR2_X1 U7302 ( .A1(n14140), .A2(n6572), .ZN(n13922) );
  AND2_X1 U7303 ( .A1(n11855), .A2(n12084), .ZN(n12747) );
  NOR2_X2 U7304 ( .A1(n12276), .A2(n14010), .ZN(n6516) );
  OAI22_X1 U7305 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(n15253), .B1(n11465), 
        .B2(n11819), .ZN(n6517) );
  OAI22_X1 U7306 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(n15253), .B1(n11465), 
        .B2(n11819), .ZN(n11824) );
  AOI21_X2 U7307 ( .B1(n11463), .B2(n11464), .A(n6804), .ZN(n11819) );
  AOI21_X1 U7308 ( .B1(n13693), .B2(n13692), .A(n11706), .ZN(n6518) );
  AOI21_X1 U7309 ( .B1(n13693), .B2(n13692), .A(n11706), .ZN(n13634) );
  XNOR2_X1 U7310 ( .A(n6813), .B(n6812), .ZN(n6519) );
  XNOR2_X1 U7311 ( .A(n6813), .B(n6812), .ZN(n14137) );
  AND2_X1 U7312 ( .A1(n7110), .A2(n12582), .ZN(n6520) );
  NAND2_X2 U7314 ( .A1(n13341), .A2(n13342), .ZN(n13340) );
  OAI21_X2 U7315 ( .B1(n10728), .B2(n10727), .A(n7880), .ZN(n10542) );
  CLKBUF_X1 U7316 ( .A(n14385), .Z(n6522) );
  XNOR2_X1 U7317 ( .A(n14316), .B(n14317), .ZN(n14385) );
  OR2_X2 U7318 ( .A1(n8360), .A2(n8359), .ZN(n8365) );
  INV_X2 U7319 ( .A(n8310), .ZN(n8439) );
  AND2_X2 U7320 ( .A1(n6850), .A2(n8678), .ZN(n8596) );
  OAI21_X2 U7321 ( .B1(n10937), .B2(n12019), .A(n12018), .ZN(n11173) );
  OAI21_X2 U7322 ( .B1(n14431), .B2(n7162), .A(n6628), .ZN(n11361) );
  INV_X1 U7324 ( .A(n12087), .ZN(n12095) );
  INV_X2 U7325 ( .A(n12328), .ZN(n12330) );
  AOI22_X1 U7326 ( .A1(n9814), .A2(P3_REG2_REG_2__SCAN_IN), .B1(n14362), .B2(
        n10051), .ZN(n9804) );
  INV_X1 U7327 ( .A(n8717), .ZN(n11896) );
  INV_X2 U7328 ( .A(n9271), .ZN(n9239) );
  BUF_X1 U7329 ( .A(n7746), .Z(n6537) );
  BUF_X1 U7330 ( .A(n7766), .Z(n9535) );
  INV_X1 U7331 ( .A(n6720), .ZN(n11700) );
  INV_X2 U7332 ( .A(n11745), .ZN(n11775) );
  CLKBUF_X3 U7333 ( .A(n9402), .Z(n12317) );
  INV_X1 U7334 ( .A(n8709), .ZN(n8989) );
  XNOR2_X1 U7335 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n8983), .ZN(n8984) );
  AOI22_X1 U7336 ( .A1(n8045), .A2(P1_DATAO_REG_3__SCAN_IN), .B1(n8044), .B2(
        n13184), .ZN(n7795) );
  INV_X1 U7337 ( .A(n12387), .ZN(n9322) );
  XNOR2_X1 U7340 ( .A(n14256), .B(n14956), .ZN(n14301) );
  INV_X1 U7341 ( .A(P3_IR_REG_4__SCAN_IN), .ZN(n8679) );
  NAND2_X1 U7342 ( .A1(n11774), .A2(n11773), .ZN(n14140) );
  NAND2_X1 U7343 ( .A1(n11051), .A2(n11050), .ZN(n12225) );
  XNOR2_X1 U7344 ( .A(n9342), .B(n9341), .ZN(n9599) );
  INV_X4 U7345 ( .A(n7626), .ZN(n9473) );
  CLKBUF_X3 U7346 ( .A(n9721), .Z(n12670) );
  BUF_X1 U7348 ( .A(n8227), .Z(n6531) );
  XOR2_X1 U7349 ( .A(n14295), .B(P2_ADDR_REG_1__SCAN_IN), .Z(n15436) );
  NAND2_X1 U7350 ( .A1(n9323), .A2(n12387), .ZN(n11601) );
  NAND2_X1 U7351 ( .A1(n7479), .A2(n11221), .ZN(n11313) );
  NOR3_X4 U7352 ( .A1(n11062), .A2(n14534), .A3(n7262), .ZN(n7264) );
  XNOR2_X1 U7353 ( .A(n8301), .B(n10839), .ZN(n10232) );
  NAND4_X2 U7354 ( .A1(n7773), .A2(n7772), .A3(n7771), .A4(n7770), .ZN(n8301)
         );
  NAND4_X2 U7355 ( .A1(n7765), .A2(n7764), .A3(n7763), .A4(n7762), .ZN(n8305)
         );
  NAND4_X4 U7356 ( .A1(n9401), .A2(n9400), .A3(n9399), .A4(n9398), .ZN(n13778)
         );
  OAI22_X2 U7357 ( .A1(n14790), .A2(n15358), .B1(n9544), .B2(n14791), .ZN(
        n13165) );
  NAND2_X2 U7358 ( .A1(n11915), .A2(n11914), .ZN(n14437) );
  NAND2_X2 U7360 ( .A1(n14104), .A2(n11498), .ZN(n14080) );
  AOI22_X2 U7361 ( .A1(n12185), .A2(n12184), .B1(n12183), .B2(n12182), .ZN(
        n12191) );
  XNOR2_X1 U7362 ( .A(n8635), .B(n6896), .ZN(n10724) );
  NAND2_X2 U7363 ( .A1(n6705), .A2(n10676), .ZN(n14629) );
  OR2_X2 U7364 ( .A1(n14037), .A2(n14048), .ZN(n14035) );
  OAI21_X2 U7365 ( .B1(n7644), .B2(n7881), .A(n7319), .ZN(n7895) );
  NAND2_X2 U7366 ( .A1(n7477), .A2(n10423), .ZN(n10675) );
  INV_X2 U7367 ( .A(n9323), .ZN(n11637) );
  BUF_X8 U7369 ( .A(n8946), .Z(n6525) );
  NAND2_X2 U7370 ( .A1(n11466), .A2(n13012), .ZN(n8946) );
  XNOR2_X2 U7371 ( .A(n14291), .B(P1_ADDR_REG_4__SCAN_IN), .ZN(n14292) );
  XNOR2_X2 U7372 ( .A(n14257), .B(n14258), .ZN(n14291) );
  NAND2_X2 U7373 ( .A1(n11428), .A2(n7260), .ZN(n9443) );
  BUF_X4 U7374 ( .A(n11601), .Z(n6526) );
  XNOR2_X2 U7375 ( .A(n14294), .B(n6737), .ZN(n14295) );
  NOR2_X2 U7376 ( .A1(n14259), .A2(n14260), .ZN(n14261) );
  NAND2_X2 U7377 ( .A1(n11315), .A2(n7483), .ZN(n14552) );
  AOI21_X2 U7378 ( .B1(n8822), .B2(n7364), .A(n7361), .ZN(n8863) );
  OAI21_X2 U7379 ( .B1(n12813), .B2(n12814), .A(n12067), .ZN(n12804) );
  NOR2_X4 U7380 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n9584) );
  XNOR2_X2 U7381 ( .A(n7105), .B(n7104), .ZN(n14958) );
  OR2_X2 U7382 ( .A1(n10067), .A2(n6590), .ZN(n7105) );
  OAI21_X2 U7383 ( .B1(n12823), .B2(n11849), .A(n12062), .ZN(n12813) );
  NAND2_X2 U7384 ( .A1(n12842), .A2(n11958), .ZN(n12823) );
  OR2_X2 U7385 ( .A1(n13776), .A2(n14714), .ZN(n12172) );
  AND2_X4 U7386 ( .A1(n8603), .A2(n8604), .ZN(n8697) );
  AND2_X2 U7387 ( .A1(n7756), .A2(n7721), .ZN(n7722) );
  NOR2_X4 U7388 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n7756) );
  OAI21_X2 U7389 ( .B1(n12850), .B2(n12849), .A(n11803), .ZN(n12836) );
  NAND2_X2 U7390 ( .A1(n14242), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9317) );
  NOR2_X1 U7391 ( .A1(n11288), .A2(n6523), .ZN(n12087) );
  AOI21_X2 U7392 ( .B1(n7347), .B2(n6678), .A(n6805), .ZN(n8983) );
  OR2_X2 U7393 ( .A1(n8936), .A2(n7349), .ZN(n7347) );
  NOR2_X2 U7394 ( .A1(n14957), .A2(n10069), .ZN(n14977) );
  NOR2_X2 U7395 ( .A1(n14958), .A2(n15156), .ZN(n14957) );
  XNOR2_X2 U7396 ( .A(n9045), .B(P1_DATAO_REG_24__SCAN_IN), .ZN(n9047) );
  INV_X2 U7397 ( .A(n9475), .ZN(n7626) );
  XNOR2_X1 U7398 ( .A(n8220), .B(n8221), .ZN(n8227) );
  AOI21_X2 U7399 ( .B1(n7035), .B2(n6739), .A(n7032), .ZN(n14256) );
  AND2_X2 U7401 ( .A1(n7027), .A2(n7026), .ZN(n14585) );
  OAI22_X2 U7402 ( .A1(n9134), .A2(n9133), .B1(P2_DATAO_REG_25__SCAN_IN), .B2(
        n11427), .ZN(n11463) );
  XNOR2_X2 U7403 ( .A(n12557), .B(n10096), .ZN(n11975) );
  NAND2_X2 U7404 ( .A1(n7033), .A2(n14324), .ZN(n14388) );
  XOR2_X2 U7405 ( .A(n14292), .B(P2_ADDR_REG_4__SCAN_IN), .Z(n15426) );
  INV_X1 U7406 ( .A(n7626), .ZN(n6533) );
  OAI21_X2 U7408 ( .B1(n14300), .B2(n14299), .A(n14348), .ZN(n15432) );
  OAI21_X1 U7409 ( .B1(n7556), .B2(n6579), .A(n7557), .ZN(n8498) );
  NAND2_X1 U7410 ( .A1(n13625), .A2(n13624), .ZN(n13623) );
  NAND2_X1 U7411 ( .A1(n13987), .A2(n13988), .ZN(n13986) );
  NAND2_X1 U7412 ( .A1(n8156), .A2(n8155), .ZN(n13469) );
  AND2_X1 U7413 ( .A1(n14001), .A2(n14006), .ZN(n14003) );
  NAND2_X1 U7414 ( .A1(n11149), .A2(n11150), .ZN(n11262) );
  AND2_X1 U7415 ( .A1(n11260), .A2(n11263), .ZN(n11261) );
  OAI21_X1 U7416 ( .B1(n8074), .B2(n7019), .A(n7016), .ZN(n7699) );
  OAI21_X1 U7417 ( .B1(n10897), .B2(n7949), .A(n7950), .ZN(n11073) );
  OR2_X1 U7418 ( .A1(n8821), .A2(n8820), .ZN(n11297) );
  NAND2_X1 U7419 ( .A1(n11496), .A2(n11495), .ZN(n14115) );
  AND2_X1 U7420 ( .A1(n11501), .A2(n11500), .ZN(n14215) );
  NAND2_X1 U7421 ( .A1(n9958), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14467) );
  NAND2_X1 U7422 ( .A1(n7307), .A2(n7306), .ZN(n7861) );
  CLKBUF_X1 U7423 ( .A(n10071), .Z(n10072) );
  AND2_X2 U7424 ( .A1(n10559), .A2(n11884), .ZN(n6902) );
  NOR2_X1 U7425 ( .A1(n12556), .A2(n10584), .ZN(n12005) );
  INV_X2 U7426 ( .A(n12179), .ZN(n12173) );
  NAND2_X2 U7427 ( .A1(n12166), .A2(n12167), .ZN(n12340) );
  XNOR2_X2 U7428 ( .A(n13159), .B(n13050), .ZN(n10254) );
  NAND2_X1 U7429 ( .A1(n13776), .A2(n14714), .ZN(n12171) );
  INV_X2 U7430 ( .A(n10439), .ZN(n11701) );
  INV_X2 U7431 ( .A(n10041), .ZN(n7482) );
  NAND2_X1 U7432 ( .A1(n13780), .A2(n10530), .ZN(n10528) );
  INV_X2 U7433 ( .A(n9535), .ZN(n8044) );
  INV_X4 U7434 ( .A(n8348), .ZN(n6534) );
  NAND2_X2 U7435 ( .A1(n9357), .A2(n12143), .ZN(n12159) );
  INV_X1 U7436 ( .A(n10724), .ZN(n11968) );
  CLKBUF_X1 U7437 ( .A(n8973), .Z(n6541) );
  INV_X1 U7438 ( .A(n11534), .ZN(n13868) );
  NAND2_X1 U7439 ( .A1(n11637), .A2(n9322), .ZN(n12325) );
  INV_X1 U7440 ( .A(n8023), .ZN(n6535) );
  BUF_X1 U7441 ( .A(P2_IR_REG_0__SCAN_IN), .Z(n15330) );
  AND2_X1 U7442 ( .A1(n12379), .A2(n12150), .ZN(n7289) );
  AOI211_X1 U7443 ( .C1(n13474), .C2(n14479), .A(n13135), .B(n13134), .ZN(
        n13136) );
  NAND2_X1 U7444 ( .A1(n8274), .A2(n7205), .ZN(n13249) );
  MUX2_X1 U7445 ( .A(n12931), .B(P3_REG1_REG_28__SCAN_IN), .S(n15129), .Z(
        n12876) );
  OR2_X1 U7446 ( .A1(n7573), .A2(n8462), .ZN(n6968) );
  NAND2_X1 U7447 ( .A1(n7526), .A2(n7524), .ZN(n13942) );
  MUX2_X1 U7448 ( .A(n12926), .B(n12710), .S(n15066), .Z(n12714) );
  NAND2_X1 U7449 ( .A1(n13243), .A2(n13246), .ZN(n13245) );
  NAND2_X1 U7450 ( .A1(n7156), .A2(n7158), .ZN(n12733) );
  NAND2_X1 U7451 ( .A1(n7440), .A2(n7441), .ZN(n13243) );
  NAND2_X1 U7452 ( .A1(n12747), .A2(n7160), .ZN(n7156) );
  NAND2_X1 U7453 ( .A1(n13277), .A2(n7442), .ZN(n7440) );
  NAND2_X1 U7454 ( .A1(n12139), .A2(n12138), .ZN(n13880) );
  NAND2_X1 U7455 ( .A1(n8267), .A2(n8266), .ZN(n13293) );
  XNOR2_X1 U7456 ( .A(n7370), .B(n6576), .ZN(n11870) );
  INV_X1 U7457 ( .A(n13914), .ZN(n6812) );
  XNOR2_X1 U7458 ( .A(n6743), .B(n12672), .ZN(n12650) );
  NAND2_X1 U7459 ( .A1(n12319), .A2(n12318), .ZN(n13887) );
  NAND2_X1 U7460 ( .A1(n7371), .A2(n6618), .ZN(n7370) );
  AOI21_X1 U7461 ( .B1(n12126), .B2(n12125), .A(n6632), .ZN(n12390) );
  NAND2_X1 U7462 ( .A1(n13107), .A2(n13106), .ZN(n7371) );
  NAND2_X1 U7463 ( .A1(n7128), .A2(n7127), .ZN(n6743) );
  OAI22_X1 U7464 ( .A1(n8505), .A2(n8504), .B1(n8503), .B2(n13010), .ZN(n8508)
         );
  XNOR2_X1 U7465 ( .A(n11869), .B(n11867), .ZN(n13107) );
  AND2_X1 U7466 ( .A1(n11916), .A2(n12099), .ZN(n11943) );
  AND2_X1 U7467 ( .A1(n6893), .A2(n6891), .ZN(n12126) );
  NAND2_X1 U7468 ( .A1(n11816), .A2(n6610), .ZN(n12734) );
  NAND2_X1 U7469 ( .A1(n8172), .A2(n8171), .ZN(n13464) );
  AOI21_X1 U7470 ( .B1(n7442), .B2(n8151), .A(n6555), .ZN(n7441) );
  NAND2_X1 U7471 ( .A1(n7208), .A2(n7209), .ZN(n13354) );
  XNOR2_X1 U7472 ( .A(n14405), .B(n14404), .ZN(n14403) );
  OAI21_X1 U7473 ( .B1(n12547), .B2(n14422), .A(n11907), .ZN(n12096) );
  NAND2_X1 U7474 ( .A1(n13986), .A2(n7075), .ZN(n13974) );
  OR2_X1 U7475 ( .A1(n14076), .A2(n7498), .ZN(n7497) );
  NAND2_X1 U7476 ( .A1(n7023), .A2(n14399), .ZN(n14405) );
  CLKBUF_X1 U7477 ( .A(n13745), .Z(n6745) );
  AND2_X1 U7478 ( .A1(n11898), .A2(n11897), .ZN(n14422) );
  NAND2_X1 U7479 ( .A1(n11330), .A2(n9268), .ZN(n14473) );
  NAND2_X1 U7480 ( .A1(n7464), .A2(n7462), .ZN(n13396) );
  OR2_X1 U7481 ( .A1(n12723), .A2(n12711), .ZN(n11907) );
  NAND2_X1 U7482 ( .A1(n12089), .A2(n11846), .ZN(n12717) );
  AND2_X1 U7483 ( .A1(n11835), .A2(n11834), .ZN(n12711) );
  NAND2_X1 U7484 ( .A1(n6831), .A2(n11575), .ZN(n13981) );
  NAND2_X1 U7485 ( .A1(n11946), .A2(n11949), .ZN(n12772) );
  NAND2_X1 U7486 ( .A1(n9138), .A2(n9137), .ZN(n12940) );
  NAND2_X1 U7487 ( .A1(n14552), .A2(n11493), .ZN(n14103) );
  NAND2_X1 U7488 ( .A1(n9051), .A2(n9050), .ZN(n12886) );
  NOR2_X1 U7489 ( .A1(n14589), .A2(n14588), .ZN(n14335) );
  NAND2_X1 U7490 ( .A1(n7110), .A2(n12582), .ZN(n7107) );
  NAND2_X1 U7491 ( .A1(n6870), .A2(n6867), .ZN(n12400) );
  CLKBUF_X1 U7492 ( .A(n11240), .Z(n6763) );
  NAND2_X1 U7493 ( .A1(n8060), .A2(n6847), .ZN(n8074) );
  NAND2_X1 U7494 ( .A1(n9030), .A2(n9029), .ZN(n9045) );
  NAND2_X1 U7495 ( .A1(n7030), .A2(n7031), .ZN(n7029) );
  OAI21_X1 U7496 ( .B1(n8997), .B2(n8998), .A(n7357), .ZN(n7356) );
  NAND2_X1 U7497 ( .A1(n11522), .A2(n11521), .ZN(n14204) );
  NAND2_X1 U7498 ( .A1(n8007), .A2(n8006), .ZN(n14480) );
  NAND2_X1 U7499 ( .A1(n6803), .A2(n8985), .ZN(n8997) );
  NAND2_X1 U7500 ( .A1(n10876), .A2(n6607), .ZN(n10997) );
  NAND2_X1 U7501 ( .A1(n8030), .A2(n8028), .ZN(n7002) );
  AOI21_X2 U7502 ( .B1(n10173), .B2(n14325), .A(n14387), .ZN(n14577) );
  NAND2_X1 U7503 ( .A1(n10615), .A2(n7486), .ZN(n10814) );
  NAND2_X2 U7504 ( .A1(n6712), .A2(n7898), .ZN(n10779) );
  NAND2_X1 U7505 ( .A1(n9986), .A2(n6574), .ZN(n10450) );
  NAND2_X1 U7506 ( .A1(n9987), .A2(n9988), .ZN(n9986) );
  NAND2_X1 U7507 ( .A1(n6704), .A2(n6670), .ZN(n10641) );
  OAI21_X1 U7508 ( .B1(n7861), .B2(n7011), .A(n6550), .ZN(n7932) );
  AND2_X2 U7509 ( .A1(n9872), .A2(n12868), .ZN(n15066) );
  AND2_X1 U7510 ( .A1(n7126), .A2(n10072), .ZN(n10075) );
  INV_X1 U7511 ( .A(n14647), .ZN(n6536) );
  INV_X2 U7512 ( .A(n13429), .ZN(n13419) );
  NAND2_X1 U7513 ( .A1(n10301), .A2(n10300), .ZN(n10421) );
  NAND2_X1 U7514 ( .A1(n7038), .A2(n14311), .ZN(n14312) );
  NAND2_X1 U7515 ( .A1(n7822), .A2(n7821), .ZN(n10479) );
  NAND2_X1 U7516 ( .A1(n10391), .A2(n10390), .ZN(n14649) );
  NAND2_X1 U7517 ( .A1(n6998), .A2(n7636), .ZN(n7833) );
  NAND2_X2 U7518 ( .A1(n12172), .A2(n12171), .ZN(n14654) );
  BUF_X2 U7519 ( .A(n10452), .Z(n6720) );
  NOR2_X1 U7520 ( .A1(n14267), .A2(n14266), .ZN(n14290) );
  XNOR2_X1 U7521 ( .A(n14307), .B(n7039), .ZN(n14376) );
  AND2_X1 U7522 ( .A1(n10364), .A2(n10363), .ZN(n15059) );
  AND2_X1 U7523 ( .A1(n12001), .A2(n12004), .ZN(n11924) );
  AND2_X1 U7524 ( .A1(n6800), .A2(n6596), .ZN(n14307) );
  NAND2_X1 U7525 ( .A1(n6999), .A2(n7633), .ZN(n7816) );
  OR2_X1 U7526 ( .A1(n13780), .A2(n14677), .ZN(n12339) );
  NAND4_X2 U7527 ( .A1(n8687), .A2(n8686), .A3(n8685), .A4(n8684), .ZN(n15037)
         );
  NAND4_X2 U7528 ( .A1(n9382), .A2(n9381), .A3(n9380), .A4(n9379), .ZN(n13780)
         );
  NAND4_X2 U7529 ( .A1(n9362), .A2(n9361), .A3(n9360), .A4(n9359), .ZN(n13779)
         );
  OR2_X1 U7530 ( .A1(n6539), .A2(n9596), .ZN(n9359) );
  CLKBUF_X1 U7531 ( .A(n7791), .Z(n8509) );
  AND3_X1 U7532 ( .A1(n8722), .A2(n8721), .A3(n8720), .ZN(n10096) );
  INV_X4 U7533 ( .A(n11896), .ZN(n11913) );
  XNOR2_X1 U7534 ( .A(P1_ADDR_REG_5__SCAN_IN), .B(n14304), .ZN(n14305) );
  NAND2_X1 U7535 ( .A1(n7766), .A2(n9473), .ZN(n7800) );
  XNOR2_X1 U7536 ( .A(n14261), .B(n14974), .ZN(n14304) );
  OR2_X1 U7537 ( .A1(n8669), .A2(n8644), .ZN(n8646) );
  NAND2_X2 U7538 ( .A1(n7741), .A2(n7740), .ZN(n8130) );
  NOR2_X1 U7539 ( .A1(n9783), .A2(n14941), .ZN(n9786) );
  INV_X2 U7540 ( .A(n12321), .ZN(n11784) );
  CLKBUF_X3 U7541 ( .A(n12325), .Z(n6540) );
  CLKBUF_X3 U7542 ( .A(n12325), .Z(n6539) );
  OR2_X1 U7543 ( .A1(n11601), .A2(n9358), .ZN(n9360) );
  OAI21_X1 U7544 ( .B1(n9350), .B2(P1_IR_REG_21__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n7074) );
  AND2_X2 U7545 ( .A1(n12387), .A2(n11637), .ZN(n12321) );
  AND2_X1 U7546 ( .A1(n13012), .A2(n8604), .ZN(n8973) );
  AND2_X1 U7547 ( .A1(n14876), .A2(n11796), .ZN(n8298) );
  XNOR2_X1 U7548 ( .A(n9337), .B(n9336), .ZN(n12143) );
  INV_X1 U7549 ( .A(n8603), .ZN(n13012) );
  NAND2_X1 U7550 ( .A1(n7732), .A2(n7731), .ZN(n9541) );
  XNOR2_X1 U7551 ( .A(n8602), .B(P3_IR_REG_29__SCAN_IN), .ZN(n8604) );
  MUX2_X1 U7552 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7729), .S(
        P2_IR_REG_27__SCAN_IN), .Z(n7732) );
  XNOR2_X1 U7553 ( .A(n8225), .B(n8224), .ZN(n11796) );
  XNOR2_X1 U7554 ( .A(n7736), .B(n13576), .ZN(n7746) );
  OR2_X1 U7555 ( .A1(n9805), .A2(n9804), .ZN(n7116) );
  OR2_X1 U7556 ( .A1(n9188), .A2(n9318), .ZN(n9342) );
  NAND2_X2 U7557 ( .A1(n9473), .A2(P1_U3086), .ZN(n14247) );
  INV_X1 U7558 ( .A(n6802), .ZN(n14257) );
  NAND2_X1 U7559 ( .A1(n6985), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8218) );
  NAND2_X1 U7560 ( .A1(n7468), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7736) );
  NOR2_X1 U7561 ( .A1(n8632), .A2(P3_IR_REG_19__SCAN_IN), .ZN(n8628) );
  NAND2_X1 U7562 ( .A1(n8219), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8220) );
  XNOR2_X1 U7563 ( .A(n8746), .B(P3_IR_REG_5__SCAN_IN), .ZN(n14966) );
  XNOR2_X1 U7564 ( .A(n6917), .B(P2_IR_REG_21__SCAN_IN), .ZN(n8549) );
  OAI21_X1 U7565 ( .B1(n9475), .B2(P2_DATAO_REG_1__SCAN_IN), .A(n6766), .ZN(
        n7621) );
  NOR2_X1 U7566 ( .A1(n10500), .A2(P1_IR_REG_18__SCAN_IN), .ZN(n9351) );
  OAI21_X1 U7567 ( .B1(n8023), .B2(n7396), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n6917) );
  NAND2_X1 U7568 ( .A1(n7779), .A2(n7793), .ZN(n13162) );
  AND2_X1 U7569 ( .A1(n6849), .A2(n8594), .ZN(n8678) );
  NAND2_X2 U7570 ( .A1(n7619), .A2(n7618), .ZN(n9475) );
  XNOR2_X1 U7571 ( .A(n8732), .B(P3_IR_REG_3__SCAN_IN), .ZN(n14952) );
  OAI21_X1 U7572 ( .B1(n14293), .B2(n14254), .A(n7036), .ZN(n7035) );
  NOR2_X1 U7573 ( .A1(n6568), .A2(n7543), .ZN(n7542) );
  AND4_X1 U7574 ( .A1(n15356), .A2(n8194), .A3(n8043), .A4(n8200), .ZN(n7724)
         );
  XNOR2_X1 U7575 ( .A(n6754), .B(P3_ADDR_REG_1__SCAN_IN), .ZN(n14293) );
  NOR3_X1 U7576 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), .A3(
        n9873), .ZN(n9781) );
  NAND2_X1 U7577 ( .A1(P3_ADDR_REG_0__SCAN_IN), .A2(n6752), .ZN(n14254) );
  AND2_X1 U7578 ( .A1(n14255), .A2(P3_ADDR_REG_2__SCAN_IN), .ZN(n7032) );
  AND2_X1 U7579 ( .A1(n9496), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n8644) );
  AND2_X1 U7580 ( .A1(n15262), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n8704) );
  XNOR2_X1 U7581 ( .A(n7102), .B(n6826), .ZN(n9734) );
  AND4_X1 U7582 ( .A1(n15380), .A2(n7720), .A3(n7719), .A4(n7718), .ZN(n7723)
         );
  INV_X1 U7583 ( .A(P3_IR_REG_1__SCAN_IN), .ZN(n7102) );
  NOR2_X1 U7584 ( .A1(P3_IR_REG_12__SCAN_IN), .A2(P3_IR_REG_10__SCAN_IN), .ZN(
        n6856) );
  NOR2_X1 U7585 ( .A1(P3_IR_REG_7__SCAN_IN), .A2(P3_IR_REG_9__SCAN_IN), .ZN(
        n6857) );
  NOR2_X1 U7586 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n7480) );
  NOR2_X1 U7587 ( .A1(P3_IR_REG_16__SCAN_IN), .A2(P3_IR_REG_13__SCAN_IN), .ZN(
        n6855) );
  INV_X1 U7588 ( .A(P3_IR_REG_20__SCAN_IN), .ZN(n8630) );
  INV_X4 U7589 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  INV_X1 U7590 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n15349) );
  INV_X1 U7591 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n6754) );
  XOR2_X1 U7592 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(P3_ADDR_REG_2__SCAN_IN), .Z(
        n14297) );
  INV_X1 U7593 ( .A(P3_IR_REG_18__SCAN_IN), .ZN(n8595) );
  INV_X1 U7594 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n8200) );
  INV_X1 U7595 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n7073) );
  INV_X1 U7596 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n15356) );
  NOR2_X1 U7597 ( .A1(P3_IR_REG_2__SCAN_IN), .A2(P3_IR_REG_3__SCAN_IN), .ZN(
        n8594) );
  INV_X4 U7598 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X1 U7599 ( .A(P3_IR_REG_11__SCAN_IN), .ZN(n8825) );
  NOR2_X1 U7600 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), .ZN(
        n8192) );
  NOR2_X1 U7601 ( .A1(P3_IR_REG_15__SCAN_IN), .A2(P3_IR_REG_14__SCAN_IN), .ZN(
        n6852) );
  NOR2_X1 U7602 ( .A1(P3_IR_REG_6__SCAN_IN), .A2(P3_IR_REG_4__SCAN_IN), .ZN(
        n6853) );
  NAND2_X1 U7603 ( .A1(n10998), .A2(n7846), .ZN(n6712) );
  NAND2_X1 U7604 ( .A1(n13930), .A2(n13932), .ZN(n7014) );
  AOI21_X1 U7605 ( .B1(n10542), .B2(n10543), .A(n6598), .ZN(n10766) );
  NOR2_X2 U7606 ( .A1(n14003), .A2(n7077), .ZN(n13987) );
  AOI21_X2 U7607 ( .B1(n12779), .B2(n12780), .A(n11852), .ZN(n12770) );
  OR2_X1 U7608 ( .A1(n15427), .A2(P2_ADDR_REG_5__SCAN_IN), .ZN(n6800) );
  OAI21_X1 U7610 ( .B1(n11607), .B2(n11606), .A(n13890), .ZN(n14145) );
  NAND2_X1 U7611 ( .A1(n7014), .A2(n6616), .ZN(n13890) );
  NOR2_X2 U7612 ( .A1(n14086), .A2(n14209), .ZN(n7270) );
  NAND2_X1 U7613 ( .A1(n13919), .A2(n13892), .ZN(n6813) );
  INV_X4 U7614 ( .A(n8393), .ZN(n8310) );
  OR2_X4 U7615 ( .A1(n10357), .A2(n8551), .ZN(n13269) );
  OAI21_X2 U7616 ( .B1(n14335), .B2(n14334), .A(n14587), .ZN(n14593) );
  NAND2_X1 U7617 ( .A1(n7932), .A2(n6848), .ZN(n7298) );
  AND2_X1 U7618 ( .A1(n7609), .A2(n7931), .ZN(n6848) );
  NAND2_X1 U7619 ( .A1(n7002), .A2(n7000), .ZN(n7687) );
  AND2_X1 U7620 ( .A1(n7683), .A2(n7001), .ZN(n7000) );
  INV_X1 U7621 ( .A(n8041), .ZN(n7001) );
  NAND2_X1 U7622 ( .A1(n7673), .A2(n7672), .ZN(n7676) );
  NAND2_X1 U7623 ( .A1(n9724), .A2(n9473), .ZN(n8852) );
  AND2_X1 U7624 ( .A1(n9724), .A2(n7626), .ZN(n8717) );
  NAND2_X1 U7625 ( .A1(n10502), .A2(P1_DATAO_REG_18__SCAN_IN), .ZN(n7353) );
  INV_X1 U7626 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n7713) );
  INV_X1 U7627 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n7712) );
  NOR2_X1 U7628 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n7715) );
  OAI21_X1 U7629 ( .B1(n8127), .B2(n8126), .A(n7705), .ZN(n8142) );
  NAND2_X1 U7630 ( .A1(n9331), .A2(n9330), .ZN(n10500) );
  INV_X1 U7631 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n9330) );
  NAND2_X1 U7632 ( .A1(n7662), .A2(n8869), .ZN(n7665) );
  OR2_X1 U7633 ( .A1(n12652), .A2(n12912), .ZN(n6702) );
  INV_X1 U7634 ( .A(n11805), .ZN(n7522) );
  NAND2_X1 U7635 ( .A1(n13104), .A2(n6609), .ZN(n11866) );
  NAND2_X1 U7636 ( .A1(n8513), .A2(n8534), .ZN(n8581) );
  AND3_X1 U7637 ( .A1(n13550), .A2(n7400), .A3(n6914), .ZN(n13239) );
  NOR2_X1 U7638 ( .A1(n13457), .A2(n6915), .ZN(n6914) );
  INV_X1 U7639 ( .A(n6916), .ZN(n6915) );
  NAND2_X1 U7640 ( .A1(n13424), .A2(n7465), .ZN(n7464) );
  NAND2_X1 U7641 ( .A1(n7766), .A2(n7626), .ZN(n7791) );
  INV_X1 U7642 ( .A(n12361), .ZN(n11606) );
  INV_X1 U7643 ( .A(n8370), .ZN(n7566) );
  NAND2_X1 U7644 ( .A1(n8364), .A2(n6599), .ZN(n7567) );
  AND2_X1 U7645 ( .A1(n8383), .A2(n7583), .ZN(n7582) );
  NAND2_X1 U7646 ( .A1(n7586), .A2(n7584), .ZN(n7583) );
  NOR2_X1 U7647 ( .A1(n6612), .A2(n6699), .ZN(n7054) );
  NOR2_X1 U7648 ( .A1(n12244), .A2(n7057), .ZN(n7056) );
  NAND2_X1 U7649 ( .A1(n7576), .A2(n7575), .ZN(n8395) );
  AND2_X1 U7650 ( .A1(n7045), .A2(n6588), .ZN(n7044) );
  NAND2_X1 U7651 ( .A1(n7048), .A2(n7046), .ZN(n7045) );
  OAI21_X1 U7652 ( .B1(n12271), .B2(n12270), .A(n12269), .ZN(n12273) );
  INV_X1 U7653 ( .A(n8823), .ZN(n7365) );
  NOR2_X1 U7654 ( .A1(n6843), .A2(n6560), .ZN(n6840) );
  OAI21_X1 U7655 ( .B1(n9473), .B2(n9492), .A(n6777), .ZN(n7638) );
  NAND2_X1 U7656 ( .A1(n9473), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n6777) );
  NAND2_X1 U7657 ( .A1(n12492), .A2(n6889), .ZN(n6888) );
  INV_X1 U7658 ( .A(n8981), .ZN(n7427) );
  INV_X1 U7659 ( .A(n12492), .ZN(n6890) );
  NAND2_X1 U7660 ( .A1(n12732), .A2(n7159), .ZN(n7158) );
  INV_X1 U7661 ( .A(n12085), .ZN(n7159) );
  NOR2_X1 U7662 ( .A1(n11182), .A2(n7514), .ZN(n7513) );
  INV_X1 U7663 ( .A(n11179), .ZN(n7514) );
  OR2_X1 U7664 ( .A1(n12958), .A2(n12414), .ZN(n11953) );
  OR2_X1 U7665 ( .A1(n12964), .A2(n12504), .ZN(n12070) );
  INV_X1 U7666 ( .A(P3_IR_REG_22__SCAN_IN), .ZN(n8618) );
  NOR2_X1 U7667 ( .A1(n8265), .A2(n7191), .ZN(n7190) );
  INV_X1 U7668 ( .A(n7193), .ZN(n7191) );
  NOR2_X1 U7669 ( .A1(n8260), .A2(n7216), .ZN(n7215) );
  INV_X1 U7670 ( .A(n8257), .ZN(n7216) );
  NOR2_X1 U7671 ( .A1(n8255), .A2(n7199), .ZN(n7198) );
  INV_X1 U7672 ( .A(n7201), .ZN(n7199) );
  NOR2_X1 U7673 ( .A1(n10860), .A2(n14516), .ZN(n6913) );
  NOR2_X1 U7674 ( .A1(n13246), .A2(n7206), .ZN(n7205) );
  INV_X1 U7675 ( .A(n8273), .ZN(n7206) );
  INV_X1 U7676 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n7720) );
  INV_X1 U7677 ( .A(n7727), .ZN(n6900) );
  INV_X1 U7678 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n8194) );
  NAND2_X1 U7679 ( .A1(n11146), .A2(n11145), .ZN(n11255) );
  NOR2_X1 U7680 ( .A1(n14531), .A2(n7254), .ZN(n7253) );
  INV_X1 U7681 ( .A(n11661), .ZN(n7254) );
  XNOR2_X1 U7682 ( .A(n14743), .B(n10699), .ZN(n12347) );
  AND2_X1 U7683 ( .A1(n14698), .A2(n6770), .ZN(n12153) );
  NOR2_X1 U7684 ( .A1(n14698), .A2(n13779), .ZN(n12151) );
  NAND2_X1 U7685 ( .A1(n11313), .A2(n11312), .ZN(n11315) );
  NAND2_X1 U7686 ( .A1(n8479), .A2(n8478), .ZN(n8482) );
  NAND2_X1 U7687 ( .A1(n7707), .A2(n7706), .ZN(n8154) );
  OAI21_X1 U7688 ( .B1(n8142), .B2(n13021), .A(n8140), .ZN(n7707) );
  NAND2_X1 U7689 ( .A1(n8142), .A2(n13021), .ZN(n7706) );
  NAND2_X1 U7690 ( .A1(n7701), .A2(n7700), .ZN(n8127) );
  NOR2_X1 U7691 ( .A1(n9172), .A2(n9176), .ZN(n9190) );
  NAND2_X1 U7692 ( .A1(n8061), .A2(n7688), .ZN(n6847) );
  AND2_X1 U7693 ( .A1(n7680), .A2(n7679), .ZN(n8019) );
  INV_X1 U7694 ( .A(n7676), .ZN(n7007) );
  INV_X1 U7695 ( .A(n7669), .ZN(n7008) );
  INV_X1 U7696 ( .A(n7998), .ZN(n7009) );
  AND2_X1 U7697 ( .A1(n7669), .A2(n7668), .ZN(n7982) );
  NAND2_X1 U7698 ( .A1(n7654), .A2(n15403), .ZN(n7657) );
  INV_X1 U7699 ( .A(n7317), .ZN(n7011) );
  AND2_X1 U7700 ( .A1(n7316), .A2(n7652), .ZN(n7315) );
  NAND2_X1 U7701 ( .A1(n7861), .A2(n7641), .ZN(n7644) );
  NOR2_X2 U7702 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n9364) );
  OAI22_X1 U7703 ( .A1(n14309), .A2(n14308), .B1(P1_ADDR_REG_6__SCAN_IN), .B2(
        n15223), .ZN(n14264) );
  INV_X1 U7704 ( .A(n7434), .ZN(n6871) );
  AND2_X1 U7705 ( .A1(n7415), .A2(n7417), .ZN(n7414) );
  INV_X1 U7706 ( .A(n12431), .ZN(n7415) );
  NAND2_X1 U7707 ( .A1(n7419), .A2(n7418), .ZN(n7417) );
  INV_X1 U7708 ( .A(n8728), .ZN(n7419) );
  NAND2_X1 U7709 ( .A1(n11287), .A2(n6523), .ZN(n6875) );
  OR2_X1 U7710 ( .A1(n9068), .A2(n9067), .ZN(n9141) );
  INV_X1 U7711 ( .A(n14428), .ZN(n11419) );
  BUF_X1 U7712 ( .A(n8698), .Z(n11899) );
  NAND2_X1 U7713 ( .A1(n6701), .A2(n6700), .ZN(n6825) );
  INV_X1 U7714 ( .A(n9793), .ZN(n6700) );
  NOR2_X1 U7715 ( .A1(n14961), .A2(n15119), .ZN(n14960) );
  NOR2_X1 U7716 ( .A1(n8745), .A2(P3_IR_REG_5__SCAN_IN), .ZN(n8671) );
  OR2_X1 U7717 ( .A1(n12559), .A2(n12558), .ZN(n12560) );
  NAND2_X1 U7718 ( .A1(n12609), .A2(n6692), .ZN(n12610) );
  NAND2_X1 U7719 ( .A1(n6702), .A2(n6591), .ZN(n6742) );
  INV_X1 U7720 ( .A(n6743), .ZN(n12665) );
  AND2_X1 U7721 ( .A1(n12732), .A2(n12081), .ZN(n7160) );
  NAND2_X1 U7722 ( .A1(n12734), .A2(n11822), .ZN(n12719) );
  NAND2_X1 U7723 ( .A1(n11180), .A2(n7513), .ZN(n7512) );
  NAND2_X1 U7724 ( .A1(n15052), .A2(n12557), .ZN(n7150) );
  AND3_X1 U7725 ( .A1(n8708), .A2(n8707), .A3(n8706), .ZN(n10149) );
  NAND2_X1 U7726 ( .A1(n12734), .A2(n7488), .ZN(n12722) );
  NOR2_X1 U7727 ( .A1(n12720), .A2(n7489), .ZN(n7488) );
  INV_X1 U7728 ( .A(n11822), .ZN(n7489) );
  AOI21_X1 U7729 ( .B1(n6716), .B2(n6543), .A(n6559), .ZN(n7521) );
  AOI21_X1 U7730 ( .B1(n12849), .B2(n12052), .A(n7140), .ZN(n7139) );
  INV_X1 U7731 ( .A(n11956), .ZN(n7140) );
  NAND2_X1 U7732 ( .A1(n7143), .A2(n12047), .ZN(n11847) );
  NOR2_X1 U7733 ( .A1(n11406), .A2(n7145), .ZN(n7144) );
  INV_X1 U7734 ( .A(n12042), .ZN(n7145) );
  NAND2_X1 U7735 ( .A1(n11288), .A2(n6523), .ZN(n15099) );
  NAND2_X1 U7736 ( .A1(n6879), .A2(n6877), .ZN(n7433) );
  AND2_X1 U7737 ( .A1(n9096), .A2(n6878), .ZN(n6877) );
  INV_X1 U7738 ( .A(P3_D_REG_0__SCAN_IN), .ZN(n6878) );
  NAND2_X1 U7739 ( .A1(n13006), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8601) );
  NAND2_X1 U7740 ( .A1(n6585), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8602) );
  NAND2_X1 U7741 ( .A1(n11487), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n7357) );
  NAND2_X1 U7742 ( .A1(n9084), .A2(n8618), .ZN(n9098) );
  NAND2_X1 U7743 ( .A1(n7350), .A2(n7353), .ZN(n7349) );
  INV_X1 U7744 ( .A(n8935), .ZN(n7350) );
  AND2_X1 U7745 ( .A1(n14457), .A2(n9260), .ZN(n7394) );
  NAND2_X1 U7746 ( .A1(n11866), .A2(n11865), .ZN(n11869) );
  NOR2_X1 U7747 ( .A1(n9288), .A2(n14890), .ZN(n9963) );
  OR2_X1 U7748 ( .A1(n8581), .A2(n8523), .ZN(n8546) );
  OR2_X1 U7749 ( .A1(n11023), .A2(n11024), .ZN(n6959) );
  NAND2_X1 U7750 ( .A1(n8084), .A2(n6573), .ZN(n7458) );
  NAND2_X1 U7751 ( .A1(n6589), .A2(n8084), .ZN(n7457) );
  AND2_X1 U7752 ( .A1(n13394), .A2(n7463), .ZN(n7462) );
  NAND2_X1 U7753 ( .A1(n8566), .A2(n6547), .ZN(n7172) );
  XNOR2_X1 U7754 ( .A(n8553), .B(n11796), .ZN(n8228) );
  NAND2_X1 U7755 ( .A1(n7734), .A2(n7733), .ZN(n13457) );
  INV_X1 U7756 ( .A(n13248), .ZN(n7207) );
  AND2_X1 U7757 ( .A1(n13405), .A2(n14901), .ZN(n13519) );
  NAND2_X1 U7758 ( .A1(n7737), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7739) );
  NAND2_X1 U7759 ( .A1(n7727), .A2(n7467), .ZN(n7737) );
  NAND2_X1 U7760 ( .A1(n8196), .A2(n8200), .ZN(n8204) );
  INV_X1 U7761 ( .A(n8199), .ZN(n8196) );
  OR2_X1 U7762 ( .A1(n7793), .A2(P2_IR_REG_3__SCAN_IN), .ZN(n7802) );
  AOI21_X1 U7763 ( .B1(n13780), .B2(n10452), .A(n9391), .ZN(n9894) );
  AND2_X1 U7764 ( .A1(n13740), .A2(n7235), .ZN(n7234) );
  NOR2_X1 U7765 ( .A1(n13721), .A2(n7236), .ZN(n7235) );
  NAND2_X1 U7766 ( .A1(n7246), .A2(n13660), .ZN(n7236) );
  OR2_X1 U7767 ( .A1(n6526), .A2(n9397), .ZN(n9399) );
  INV_X1 U7768 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n7616) );
  XNOR2_X1 U7769 ( .A(n14153), .B(n11621), .ZN(n13932) );
  OR2_X1 U7770 ( .A1(n14165), .A2(n11619), .ZN(n11620) );
  AOI21_X1 U7771 ( .B1(n7528), .B2(n7531), .A(n7525), .ZN(n7524) );
  INV_X1 U7772 ( .A(n13952), .ZN(n7525) );
  XNOR2_X1 U7773 ( .A(n14159), .B(n11583), .ZN(n13952) );
  NAND2_X1 U7774 ( .A1(n6769), .A2(n6545), .ZN(n6788) );
  INV_X1 U7775 ( .A(n12353), .ZN(n11312) );
  INV_X1 U7776 ( .A(n14029), .ZN(n14192) );
  NOR2_X1 U7777 ( .A1(n14747), .A2(n9357), .ZN(n14220) );
  INV_X1 U7778 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n9332) );
  NAND2_X1 U7779 ( .A1(n7002), .A2(n7683), .ZN(n8042) );
  OAI21_X1 U7780 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(n14276), .A(n14275), .ZN(
        n14286) );
  OAI21_X1 U7781 ( .B1(n14400), .B2(n14401), .A(P2_ADDR_REG_17__SCAN_IN), .ZN(
        n7023) );
  NAND2_X1 U7782 ( .A1(n6703), .A2(n12587), .ZN(n12562) );
  OR2_X1 U7783 ( .A1(n12560), .A2(n12582), .ZN(n6703) );
  NAND2_X1 U7784 ( .A1(n6947), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n6945) );
  INV_X1 U7785 ( .A(n6758), .ZN(n6757) );
  NAND2_X1 U7786 ( .A1(n13226), .A2(n14870), .ZN(n6759) );
  NAND2_X1 U7787 ( .A1(n7444), .A2(n8576), .ZN(n13244) );
  INV_X1 U7788 ( .A(n13243), .ZN(n7444) );
  AOI21_X1 U7789 ( .B1(n11626), .B2(n14694), .A(n11625), .ZN(n11627) );
  NAND2_X1 U7790 ( .A1(n7029), .A2(n7028), .ZN(n7026) );
  AOI21_X1 U7791 ( .B1(n12178), .B2(n12177), .A(n12176), .ZN(n12180) );
  NAND2_X1 U7792 ( .A1(n12170), .A2(n12169), .ZN(n12177) );
  NOR2_X1 U7793 ( .A1(n8345), .A2(n8342), .ZN(n6971) );
  INV_X1 U7794 ( .A(n8342), .ZN(n6972) );
  OAI22_X1 U7795 ( .A1(n12202), .A2(n7070), .B1(n12203), .B2(n7069), .ZN(
        n12208) );
  NOR2_X1 U7796 ( .A1(n12201), .A2(n12204), .ZN(n7070) );
  INV_X1 U7797 ( .A(n12201), .ZN(n7069) );
  NOR2_X1 U7798 ( .A1(n8364), .A2(n6599), .ZN(n7568) );
  OAI21_X1 U7799 ( .B1(n7567), .B2(n7566), .A(n7564), .ZN(n7563) );
  INV_X1 U7800 ( .A(n8368), .ZN(n7564) );
  NOR2_X1 U7801 ( .A1(n7568), .A2(n7566), .ZN(n7565) );
  INV_X1 U7802 ( .A(n12245), .ZN(n7057) );
  NAND2_X1 U7803 ( .A1(n6729), .A2(n7067), .ZN(n12220) );
  OR2_X1 U7804 ( .A1(n7068), .A2(n12216), .ZN(n7067) );
  NAND2_X1 U7805 ( .A1(n12244), .A2(n7057), .ZN(n7055) );
  OAI21_X1 U7806 ( .B1(n8377), .B2(n7586), .A(n6973), .ZN(n7612) );
  NOR2_X1 U7807 ( .A1(n8383), .A2(n6974), .ZN(n6973) );
  NAND2_X1 U7808 ( .A1(n7578), .A2(n7580), .ZN(n7577) );
  INV_X1 U7809 ( .A(n8388), .ZN(n7578) );
  AND2_X1 U7810 ( .A1(n8387), .A2(n8388), .ZN(n7579) );
  AND2_X1 U7811 ( .A1(n7058), .A2(n7049), .ZN(n7048) );
  NAND2_X1 U7812 ( .A1(n7600), .A2(n7597), .ZN(n8407) );
  NAND2_X1 U7813 ( .A1(n7599), .A2(n7598), .ZN(n7597) );
  INV_X1 U7814 ( .A(n8401), .ZN(n7599) );
  AND2_X1 U7815 ( .A1(n7042), .A2(n12265), .ZN(n7041) );
  NOR2_X1 U7816 ( .A1(n6578), .A2(n6552), .ZN(n6995) );
  NAND2_X1 U7817 ( .A1(n6644), .A2(n6558), .ZN(n6988) );
  AOI21_X1 U7818 ( .B1(n6643), .B2(n6996), .A(n6991), .ZN(n6990) );
  INV_X1 U7819 ( .A(n8434), .ZN(n7594) );
  NAND2_X1 U7820 ( .A1(n12285), .A2(n7061), .ZN(n7060) );
  INV_X1 U7821 ( .A(n12284), .ZN(n7061) );
  AND2_X1 U7822 ( .A1(n7338), .A2(n6654), .ZN(n7336) );
  INV_X1 U7823 ( .A(n7697), .ZN(n7017) );
  INV_X1 U7824 ( .A(n7692), .ZN(n7018) );
  NOR2_X1 U7825 ( .A1(n15037), .A2(n15061), .ZN(n11988) );
  INV_X1 U7826 ( .A(n6669), .ZN(n7363) );
  NAND2_X1 U7827 ( .A1(n6968), .A2(n6967), .ZN(n8469) );
  AND2_X1 U7828 ( .A1(n7571), .A2(n6626), .ZN(n6967) );
  NAND2_X1 U7829 ( .A1(n8472), .A2(n8474), .ZN(n7559) );
  NAND2_X1 U7830 ( .A1(n7570), .A2(n7569), .ZN(n8468) );
  AOI21_X1 U7831 ( .B1(n7573), .B2(n7571), .A(n6626), .ZN(n7569) );
  INV_X1 U7832 ( .A(n8474), .ZN(n7558) );
  AND2_X1 U7833 ( .A1(n6554), .A2(n7090), .ZN(n7088) );
  NAND2_X1 U7834 ( .A1(n6835), .A2(n7680), .ZN(n7681) );
  AOI21_X1 U7835 ( .B1(n7006), .B2(n7009), .A(n7005), .ZN(n7004) );
  NAND2_X1 U7836 ( .A1(n7677), .A2(n15158), .ZN(n7680) );
  AOI21_X1 U7837 ( .B1(n7665), .B2(n7964), .A(n7313), .ZN(n7311) );
  INV_X1 U7838 ( .A(n7982), .ZN(n7313) );
  AOI21_X1 U7839 ( .B1(n7645), .B2(n7320), .A(n6629), .ZN(n7319) );
  INV_X1 U7840 ( .A(n7643), .ZN(n7320) );
  OR2_X1 U7841 ( .A1(n9954), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n9586) );
  AOI21_X1 U7842 ( .B1(n7832), .B2(n7639), .A(n7844), .ZN(n7309) );
  INV_X1 U7843 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n9488) );
  NAND2_X1 U7844 ( .A1(n10041), .A2(n10149), .ZN(n11974) );
  INV_X1 U7845 ( .A(n7431), .ZN(n7430) );
  AOI21_X1 U7846 ( .B1(n7431), .B2(n10917), .A(n7429), .ZN(n7428) );
  NOR2_X1 U7847 ( .A1(n8809), .A2(n10918), .ZN(n7429) );
  AND2_X1 U7848 ( .A1(n12480), .A2(n9066), .ZN(n9143) );
  NOR2_X1 U7849 ( .A1(n12651), .A2(n7287), .ZN(n12679) );
  NOR2_X1 U7850 ( .A1(n12636), .A2(n12919), .ZN(n7287) );
  OR2_X1 U7851 ( .A1(n12671), .A2(n6747), .ZN(n6746) );
  NOR2_X1 U7852 ( .A1(n12680), .A2(n6748), .ZN(n6747) );
  INV_X1 U7853 ( .A(n12673), .ZN(n6748) );
  NAND2_X1 U7854 ( .A1(n11812), .A2(n7495), .ZN(n7494) );
  INV_X1 U7855 ( .A(n12780), .ZN(n7495) );
  NOR2_X1 U7856 ( .A1(n7131), .A2(n7134), .ZN(n7130) );
  INV_X1 U7857 ( .A(n11924), .ZN(n7131) );
  OR2_X1 U7858 ( .A1(n15053), .A2(n15046), .ZN(n11999) );
  NAND2_X1 U7859 ( .A1(n11973), .A2(n11974), .ZN(n10153) );
  OR2_X1 U7860 ( .A1(n12886), .A2(n15345), .ZN(n12084) );
  OR2_X1 U7861 ( .A1(n12940), .A2(n12735), .ZN(n12081) );
  NAND2_X1 U7862 ( .A1(n12491), .A2(n12784), .ZN(n11946) );
  NAND2_X1 U7863 ( .A1(n12947), .A2(n11811), .ZN(n11949) );
  INV_X1 U7864 ( .A(n7513), .ZN(n7508) );
  NAND4_X1 U7865 ( .A1(n7147), .A2(n8690), .A3(n8689), .A4(n7146), .ZN(n11969)
         );
  NOR2_X1 U7866 ( .A1(n6568), .A2(P3_IR_REG_19__SCAN_IN), .ZN(n7544) );
  INV_X1 U7867 ( .A(n8632), .ZN(n7545) );
  NAND2_X1 U7868 ( .A1(P2_DATAO_REG_23__SCAN_IN), .A2(n9028), .ZN(n9029) );
  NOR2_X1 U7869 ( .A1(n7334), .A2(n7331), .ZN(n7330) );
  INV_X1 U7870 ( .A(n8882), .ZN(n7331) );
  INV_X1 U7871 ( .A(n8884), .ZN(n7333) );
  INV_X1 U7872 ( .A(n7344), .ZN(n7343) );
  OAI21_X1 U7873 ( .B1(n8766), .B2(n7345), .A(n8774), .ZN(n7344) );
  INV_X1 U7874 ( .A(n8647), .ZN(n7345) );
  OR3_X1 U7875 ( .A1(n8777), .A2(P3_IR_REG_7__SCAN_IN), .A3(
        P3_IR_REG_8__SCAN_IN), .ZN(n8791) );
  NOR2_X1 U7876 ( .A1(n7326), .A2(n7323), .ZN(n7322) );
  INV_X1 U7877 ( .A(n8643), .ZN(n7325) );
  INV_X1 U7878 ( .A(n7378), .ZN(n7375) );
  INV_X1 U7879 ( .A(n8094), .ZN(n7456) );
  NAND2_X1 U7880 ( .A1(n10848), .A2(n8248), .ZN(n10899) );
  NOR2_X1 U7881 ( .A1(n10729), .A2(n7183), .ZN(n7182) );
  AND2_X1 U7882 ( .A1(n7186), .A2(n8241), .ZN(n7183) );
  OR2_X1 U7883 ( .A1(n10737), .A2(n10750), .ZN(n10550) );
  NOR2_X1 U7884 ( .A1(n8238), .A2(n8560), .ZN(n7437) );
  INV_X1 U7885 ( .A(n8264), .ZN(n7195) );
  AOI21_X1 U7886 ( .B1(n8264), .B2(n7194), .A(n6601), .ZN(n7193) );
  INV_X1 U7887 ( .A(n8263), .ZN(n7194) );
  NAND2_X1 U7888 ( .A1(n8237), .A2(n8236), .ZN(n10186) );
  NAND2_X1 U7889 ( .A1(n10558), .A2(n10557), .ZN(n10556) );
  INV_X1 U7890 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n7726) );
  INV_X1 U7891 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n7735) );
  NAND2_X1 U7892 ( .A1(n12313), .A2(n12314), .ZN(n7293) );
  XNOR2_X1 U7893 ( .A(n13891), .B(n13908), .ZN(n12361) );
  NAND2_X1 U7894 ( .A1(n13963), .A2(n11619), .ZN(n7535) );
  AND2_X1 U7895 ( .A1(n11046), .A2(n11002), .ZN(n12352) );
  INV_X1 U7896 ( .A(n14649), .ZN(n12187) );
  INV_X1 U7897 ( .A(n13957), .ZN(n13969) );
  NOR2_X1 U7898 ( .A1(n7537), .A2(n13969), .ZN(n7532) );
  NAND2_X1 U7899 ( .A1(n7534), .A2(n6571), .ZN(n7533) );
  AND2_X1 U7900 ( .A1(n14056), .A2(n11615), .ZN(n7097) );
  NAND2_X1 U7901 ( .A1(n8170), .A2(n7711), .ZN(n8479) );
  INV_X1 U7902 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n9341) );
  INV_X1 U7903 ( .A(n8073), .ZN(n7021) );
  NAND2_X1 U7904 ( .A1(n7687), .A2(n6681), .ZN(n8061) );
  NAND2_X1 U7905 ( .A1(n7689), .A2(n10609), .ZN(n8060) );
  AND2_X2 U7906 ( .A1(n7259), .A2(n7256), .ZN(n9331) );
  NAND2_X1 U7907 ( .A1(n7258), .A2(n9498), .ZN(n7257) );
  INV_X1 U7908 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n7258) );
  AND2_X1 U7909 ( .A1(n7676), .A2(n7675), .ZN(n7998) );
  NAND2_X1 U7910 ( .A1(n7665), .A2(n7663), .ZN(n7965) );
  NAND2_X1 U7911 ( .A1(n7648), .A2(SI_11_), .ZN(n7913) );
  INV_X1 U7912 ( .A(n14297), .ZN(n6739) );
  NOR2_X1 U7913 ( .A1(n14313), .A2(n14265), .ZN(n14266) );
  AND2_X1 U7914 ( .A1(n7603), .A2(n8840), .ZN(n7434) );
  NOR2_X1 U7915 ( .A1(n6871), .A2(n11389), .ZN(n6868) );
  NOR2_X1 U7916 ( .A1(n12418), .A2(n7432), .ZN(n7431) );
  INV_X1 U7917 ( .A(n8807), .ZN(n7432) );
  NAND2_X1 U7918 ( .A1(n7421), .A2(n7420), .ZN(n7416) );
  NAND2_X1 U7919 ( .A1(n11297), .A2(n12553), .ZN(n6874) );
  NAND2_X1 U7920 ( .A1(n6892), .A2(n12797), .ZN(n6891) );
  OR2_X1 U7921 ( .A1(n9019), .A2(n6675), .ZN(n6893) );
  INV_X1 U7922 ( .A(n9018), .ZN(n6892) );
  OAI22_X1 U7923 ( .A1(n7412), .A2(n9995), .B1(n8741), .B2(n7414), .ZN(n10109)
         );
  INV_X1 U7924 ( .A(n8741), .ZN(n7413) );
  AND2_X1 U7925 ( .A1(n8740), .A2(n15054), .ZN(n8741) );
  NAND2_X1 U7926 ( .A1(n8805), .A2(n8804), .ZN(n10914) );
  NAND2_X1 U7927 ( .A1(n6873), .A2(n6872), .ZN(n11387) );
  AND2_X1 U7928 ( .A1(n6874), .A2(n11389), .ZN(n6873) );
  AOI21_X1 U7929 ( .B1(n6544), .B2(n6890), .A(n6887), .ZN(n6886) );
  OAI21_X1 U7930 ( .B1(n12441), .B2(n6890), .A(n6544), .ZN(n12447) );
  OR2_X1 U7931 ( .A1(n12501), .A2(n12807), .ZN(n12499) );
  NAND2_X1 U7932 ( .A1(n6861), .A2(n6859), .ZN(n12510) );
  AOI21_X1 U7933 ( .B1(n6862), .B2(n6864), .A(n6860), .ZN(n6859) );
  INV_X1 U7934 ( .A(n8934), .ZN(n6860) );
  OR2_X1 U7935 ( .A1(n9145), .A2(n9144), .ZN(n12123) );
  NAND2_X1 U7936 ( .A1(n12126), .A2(n12120), .ZN(n12389) );
  NAND2_X1 U7937 ( .A1(n7411), .A2(n8880), .ZN(n12398) );
  INV_X1 U7938 ( .A(n12400), .ZN(n7411) );
  INV_X1 U7939 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n15376) );
  AND4_X1 U7940 ( .A1(n8950), .A2(n8949), .A3(n8948), .A4(n8947), .ZN(n11804)
         );
  OR2_X1 U7941 ( .A1(n9097), .A2(n11352), .ZN(n9195) );
  OR2_X1 U7942 ( .A1(n6525), .A2(n8688), .ZN(n8689) );
  NOR2_X1 U7943 ( .A1(n9786), .A2(n9785), .ZN(n10067) );
  INV_X1 U7944 ( .A(n14966), .ZN(n7104) );
  NOR2_X1 U7945 ( .A1(n14960), .A2(n10079), .ZN(n14981) );
  OR2_X1 U7946 ( .A1(n14981), .A2(n14980), .ZN(n6823) );
  NAND2_X1 U7947 ( .A1(n6740), .A2(n6676), .ZN(n7274) );
  NAND2_X1 U7948 ( .A1(n6820), .A2(n7272), .ZN(n12609) );
  NAND2_X1 U7949 ( .A1(n12621), .A2(n12620), .ZN(n12632) );
  NAND2_X1 U7950 ( .A1(n6715), .A2(n6714), .ZN(n7128) );
  INV_X1 U7951 ( .A(n12640), .ZN(n6714) );
  INV_X1 U7952 ( .A(n12668), .ZN(n7113) );
  OR2_X1 U7953 ( .A1(n9117), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n9149) );
  NAND2_X1 U7954 ( .A1(n9006), .A2(n9005), .ZN(n9035) );
  NOR2_X1 U7955 ( .A1(n11933), .A2(n7511), .ZN(n7510) );
  INV_X1 U7956 ( .A(n7515), .ZN(n7511) );
  NAND2_X1 U7957 ( .A1(n7512), .A2(n7515), .ZN(n11183) );
  NAND2_X1 U7958 ( .A1(n7165), .A2(n7164), .ZN(n14433) );
  NAND2_X1 U7959 ( .A1(n10814), .A2(n7485), .ZN(n10941) );
  AND2_X1 U7960 ( .A1(n12016), .A2(n10813), .ZN(n7485) );
  AND3_X1 U7961 ( .A1(n8781), .A2(n8780), .A3(n8779), .ZN(n10756) );
  INV_X1 U7962 ( .A(n12007), .ZN(n11928) );
  NOR2_X1 U7963 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n8749) );
  INV_X1 U7964 ( .A(n11969), .ZN(n10150) );
  NOR2_X1 U7965 ( .A1(n7553), .A2(n7552), .ZN(n7551) );
  NOR2_X1 U7966 ( .A1(n11844), .A2(n14418), .ZN(n7553) );
  NOR2_X1 U7967 ( .A1(n12736), .A2(n12864), .ZN(n7552) );
  OR2_X1 U7968 ( .A1(n11832), .A2(n11896), .ZN(n11835) );
  INV_X1 U7969 ( .A(n15345), .ZN(n12773) );
  AND2_X1 U7970 ( .A1(n12772), .A2(n11810), .ZN(n7496) );
  OR2_X1 U7971 ( .A1(n12781), .A2(n12780), .ZN(n12783) );
  AND2_X1 U7972 ( .A1(n12814), .A2(n6543), .ZN(n7520) );
  NAND2_X1 U7973 ( .A1(n7518), .A2(n6604), .ZN(n7517) );
  NAND2_X1 U7974 ( .A1(n12067), .A2(n12066), .ZN(n12814) );
  NAND2_X1 U7975 ( .A1(n7523), .A2(n12839), .ZN(n12834) );
  INV_X1 U7976 ( .A(n12836), .ZN(n7523) );
  AND2_X1 U7977 ( .A1(n11959), .A2(n11956), .ZN(n12849) );
  AND2_X1 U7978 ( .A1(n12048), .A2(n12047), .ZN(n12045) );
  INV_X1 U7979 ( .A(n12045), .ZN(n11406) );
  OR2_X1 U7980 ( .A1(n7162), .A2(n12030), .ZN(n7161) );
  NAND2_X1 U7981 ( .A1(n7163), .A2(n11933), .ZN(n7162) );
  AND3_X1 U7982 ( .A1(n8675), .A2(n8674), .A3(n8673), .ZN(n15086) );
  AND2_X1 U7983 ( .A1(n8654), .A2(n8651), .ZN(n7166) );
  NAND2_X1 U7984 ( .A1(n7546), .A2(n8595), .ZN(n7543) );
  NOR2_X1 U7985 ( .A1(P3_IR_REG_26__SCAN_IN), .A2(P3_IR_REG_19__SCAN_IN), .ZN(
        n7546) );
  INV_X1 U7986 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n8654) );
  AND2_X1 U7987 ( .A1(n6664), .A2(n8630), .ZN(n6895) );
  NOR2_X1 U7988 ( .A1(n8634), .A2(P3_IR_REG_21__SCAN_IN), .ZN(n9084) );
  NAND2_X1 U7989 ( .A1(n8984), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n6803) );
  NAND2_X1 U7990 ( .A1(n6683), .A2(n7353), .ZN(n7348) );
  INV_X1 U7991 ( .A(n7354), .ZN(n7351) );
  NAND2_X1 U7992 ( .A1(P2_DATAO_REG_17__SCAN_IN), .A2(n10179), .ZN(n7354) );
  NAND2_X1 U7993 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n7671), .ZN(n8913) );
  OR2_X1 U7994 ( .A1(P1_DATAO_REG_14__SCAN_IN), .A2(n9848), .ZN(n8882) );
  NAND2_X1 U7995 ( .A1(n8865), .A2(n8864), .ZN(n8883) );
  INV_X1 U7996 ( .A(n8822), .ZN(n7367) );
  XNOR2_X1 U7997 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(P2_DATAO_REG_8__SCAN_IN), 
        .ZN(n8774) );
  XNOR2_X1 U7998 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .ZN(n8766) );
  NAND2_X1 U7999 ( .A1(n8642), .A2(n8641), .ZN(n8677) );
  INV_X1 U8000 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n8640) );
  INV_X1 U8001 ( .A(n7103), .ZN(n6849) );
  AOI21_X1 U8002 ( .B1(n7387), .B2(n13038), .A(n7386), .ZN(n7385) );
  AND2_X1 U8003 ( .A1(n13068), .A2(n13064), .ZN(n7386) );
  INV_X1 U8004 ( .A(n6924), .ZN(n6921) );
  NAND2_X1 U8005 ( .A1(n6924), .A2(n7375), .ZN(n6923) );
  OR2_X1 U8006 ( .A1(n11114), .A2(n11115), .ZN(n11112) );
  INV_X1 U8007 ( .A(n9312), .ZN(n9244) );
  AOI21_X1 U8008 ( .B1(n7378), .B2(n7374), .A(n6633), .ZN(n7373) );
  INV_X1 U8009 ( .A(n9270), .ZN(n7374) );
  AND2_X1 U8010 ( .A1(n6925), .A2(n7373), .ZN(n6924) );
  INV_X1 U8011 ( .A(n13119), .ZN(n6925) );
  AOI21_X1 U8012 ( .B1(n7394), .B2(n11115), .A(n6637), .ZN(n7392) );
  INV_X1 U8013 ( .A(n8581), .ZN(n8542) );
  NAND2_X1 U8014 ( .A1(n6979), .A2(n6978), .ZN(n6977) );
  INV_X1 U8015 ( .A(n8496), .ZN(n6978) );
  NAND2_X1 U8016 ( .A1(n8498), .A2(n8497), .ZN(n6979) );
  NAND2_X1 U8017 ( .A1(n8500), .A2(n8501), .ZN(n6982) );
  AND2_X1 U8018 ( .A1(n8548), .A2(n6981), .ZN(n6980) );
  INV_X1 U8019 ( .A(n8499), .ZN(n6981) );
  OR2_X1 U8020 ( .A1(n8488), .A2(n9564), .ZN(n7765) );
  OR2_X1 U8021 ( .A1(n14803), .A2(n14802), .ZN(n6955) );
  NAND2_X1 U8022 ( .A1(n6955), .A2(n6954), .ZN(n6953) );
  NAND2_X1 U8023 ( .A1(n14806), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6954) );
  AND2_X1 U8024 ( .A1(n6953), .A2(n6952), .ZN(n14814) );
  INV_X1 U8025 ( .A(n14815), .ZN(n6952) );
  AND2_X1 U8026 ( .A1(n6959), .A2(n6958), .ZN(n11166) );
  OR2_X1 U8027 ( .A1(n11166), .A2(n11167), .ZN(n6957) );
  INV_X1 U8028 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n6830) );
  OR2_X1 U8029 ( .A1(n13474), .A2(n13294), .ZN(n7445) );
  NAND2_X1 U8030 ( .A1(n7448), .A2(n7447), .ZN(n7446) );
  INV_X1 U8031 ( .A(n13277), .ZN(n7448) );
  NOR2_X1 U8032 ( .A1(n8125), .A2(n7452), .ZN(n7451) );
  INV_X1 U8033 ( .A(n8558), .ZN(n7452) );
  INV_X1 U8034 ( .A(n8572), .ZN(n13342) );
  AOI21_X1 U8035 ( .B1(n7212), .B2(n7211), .A(n7210), .ZN(n7209) );
  NAND2_X1 U8036 ( .A1(n6764), .A2(n7212), .ZN(n7208) );
  INV_X1 U8037 ( .A(n7215), .ZN(n7211) );
  NOR2_X1 U8038 ( .A1(n13370), .A2(n7213), .ZN(n7212) );
  INV_X1 U8039 ( .A(n8259), .ZN(n7213) );
  NAND2_X1 U8040 ( .A1(n8258), .A2(n7215), .ZN(n7214) );
  INV_X1 U8041 ( .A(n8254), .ZN(n7203) );
  AOI21_X1 U8042 ( .B1(n8254), .B2(n7202), .A(n6614), .ZN(n7201) );
  INV_X1 U8043 ( .A(n8253), .ZN(n7202) );
  NAND2_X1 U8044 ( .A1(n7972), .A2(n7971), .ZN(n11233) );
  OR2_X1 U8045 ( .A1(n8567), .A2(n8249), .ZN(n7174) );
  OR2_X1 U8046 ( .A1(n9961), .A2(n8284), .ZN(n13538) );
  NAND2_X1 U8047 ( .A1(n10186), .A2(n8238), .ZN(n8240) );
  NOR2_X1 U8048 ( .A1(n10484), .A2(n6903), .ZN(n10738) );
  NAND2_X1 U8049 ( .A1(n10222), .A2(n10225), .ZN(n10221) );
  INV_X1 U8050 ( .A(n10240), .ZN(n7178) );
  INV_X1 U8051 ( .A(n13534), .ZN(n13407) );
  NAND2_X1 U8052 ( .A1(n8305), .A2(n10358), .ZN(n8559) );
  NAND2_X1 U8053 ( .A1(n8076), .A2(n8075), .ZN(n13359) );
  AND2_X1 U8054 ( .A1(n7724), .A2(n6651), .ZN(n6897) );
  AND2_X1 U8055 ( .A1(n7726), .A2(n7735), .ZN(n7467) );
  INV_X1 U8056 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n8197) );
  NAND2_X1 U8057 ( .A1(n7396), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7395) );
  INV_X1 U8058 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n8221) );
  NAND2_X1 U8059 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), 
        .ZN(n6984) );
  AND2_X1 U8060 ( .A1(n11210), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n11212) );
  NAND2_X1 U8061 ( .A1(n13709), .A2(n11724), .ZN(n13614) );
  NAND2_X1 U8062 ( .A1(n11255), .A2(n11254), .ZN(n11260) );
  AND2_X1 U8063 ( .A1(n7231), .A2(n13654), .ZN(n7230) );
  NAND2_X1 U8064 ( .A1(n7232), .A2(n13684), .ZN(n7231) );
  NAND2_X1 U8065 ( .A1(n7246), .A2(n7243), .ZN(n7242) );
  INV_X1 U8066 ( .A(n13670), .ZN(n7243) );
  NAND2_X1 U8067 ( .A1(n10450), .A2(n10449), .ZN(n10632) );
  OR2_X1 U8068 ( .A1(n11552), .A2(n15196), .ZN(n11554) );
  NOR2_X1 U8069 ( .A1(n10590), .A2(n7220), .ZN(n7219) );
  INV_X1 U8070 ( .A(n10634), .ZN(n7220) );
  NAND2_X1 U8071 ( .A1(n10442), .A2(n10446), .ZN(n10633) );
  INV_X1 U8072 ( .A(n7230), .ZN(n7229) );
  AOI21_X1 U8073 ( .B1(n7230), .B2(n7233), .A(n7228), .ZN(n7227) );
  INV_X1 U8074 ( .A(n11753), .ZN(n7228) );
  NAND2_X1 U8075 ( .A1(n11674), .A2(n11673), .ZN(n13745) );
  NOR2_X1 U8076 ( .A1(n6549), .A2(n6580), .ZN(n6798) );
  XNOR2_X1 U8077 ( .A(n13880), .B(n13877), .ZN(n12378) );
  AOI21_X1 U8078 ( .B1(P1_REG1_REG_2__SCAN_IN), .B2(n9598), .A(n9904), .ZN(
        n9601) );
  NAND2_X1 U8079 ( .A1(n13910), .A2(n7607), .ZN(n13918) );
  OR2_X1 U8080 ( .A1(n13909), .A2(n13908), .ZN(n7607) );
  OR2_X1 U8081 ( .A1(n13891), .A2(n13908), .ZN(n7015) );
  XNOR2_X1 U8082 ( .A(n14140), .B(n13913), .ZN(n13921) );
  NAND2_X1 U8083 ( .A1(n13890), .A2(n7012), .ZN(n13919) );
  NOR2_X1 U8084 ( .A1(n13921), .A2(n7013), .ZN(n7012) );
  INV_X1 U8085 ( .A(n7015), .ZN(n7013) );
  NOR2_X1 U8086 ( .A1(n13952), .A2(n7091), .ZN(n7090) );
  INV_X1 U8087 ( .A(n11620), .ZN(n7091) );
  NAND2_X1 U8088 ( .A1(n13942), .A2(n6602), .ZN(n13930) );
  OR2_X1 U8089 ( .A1(n7532), .A2(n7529), .ZN(n7528) );
  INV_X1 U8090 ( .A(n7535), .ZN(n7529) );
  NAND2_X1 U8092 ( .A1(n13997), .A2(n7076), .ZN(n6785) );
  INV_X1 U8093 ( .A(n13988), .ZN(n6787) );
  NAND2_X1 U8094 ( .A1(n12276), .A2(n7076), .ZN(n7075) );
  XOR2_X1 U8095 ( .A(n13759), .B(n13997), .Z(n13988) );
  INV_X1 U8096 ( .A(n14006), .ZN(n6761) );
  NAND2_X1 U8097 ( .A1(n11547), .A2(n11546), .ZN(n14031) );
  AND2_X1 U8098 ( .A1(n7501), .A2(n14048), .ZN(n7500) );
  INV_X1 U8099 ( .A(n12336), .ZN(n7505) );
  NOR2_X1 U8100 ( .A1(n11523), .A2(n10130), .ZN(n11540) );
  AOI21_X1 U8102 ( .B1(n14097), .B2(n11611), .A(n6582), .ZN(n14084) );
  AOI21_X1 U8103 ( .B1(n7082), .B2(n7084), .A(n6623), .ZN(n7080) );
  NAND2_X1 U8104 ( .A1(n10997), .A2(n7099), .ZN(n11047) );
  NOR2_X1 U8105 ( .A1(n11066), .A2(n7100), .ZN(n7099) );
  INV_X1 U8106 ( .A(n10996), .ZN(n7100) );
  AND2_X1 U8107 ( .A1(n14635), .A2(n10716), .ZN(n10890) );
  NAND2_X1 U8108 ( .A1(n10683), .A2(n10682), .ZN(n10868) );
  NAND2_X1 U8109 ( .A1(n6724), .A2(n6723), .ZN(n10876) );
  INV_X1 U8110 ( .A(n12346), .ZN(n6723) );
  OR2_X1 U8111 ( .A1(n11745), .A2(n10296), .ZN(n10525) );
  INV_X1 U8112 ( .A(n13880), .ZN(n14122) );
  NAND2_X1 U8113 ( .A1(n11585), .A2(n11584), .ZN(n14153) );
  NAND2_X1 U8114 ( .A1(n7003), .A2(n11475), .ZN(n14159) );
  NAND2_X1 U8115 ( .A1(n11474), .A2(n10677), .ZN(n7003) );
  NAND2_X1 U8116 ( .A1(n11513), .A2(n11512), .ZN(n14209) );
  NOR2_X1 U8117 ( .A1(n12247), .A2(n7484), .ZN(n7483) );
  INV_X1 U8118 ( .A(n11314), .ZN(n7484) );
  NAND2_X1 U8119 ( .A1(n12141), .A2(n12329), .ZN(n14694) );
  OR2_X1 U8120 ( .A1(n9402), .A2(n9477), .ZN(n9367) );
  OR2_X1 U8121 ( .A1(n10388), .A2(n9478), .ZN(n9368) );
  INV_X1 U8122 ( .A(n14742), .ZN(n14767) );
  AND2_X1 U8123 ( .A1(n9421), .A2(n9514), .ZN(n14221) );
  AND2_X1 U8124 ( .A1(n9331), .A2(n7538), .ZN(n9319) );
  AND2_X1 U8125 ( .A1(n7610), .A2(n7539), .ZN(n7538) );
  NOR2_X1 U8126 ( .A1(n7540), .A2(P1_IR_REG_28__SCAN_IN), .ZN(n7539) );
  INV_X1 U8127 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n9320) );
  NAND2_X1 U8128 ( .A1(n8168), .A2(n8167), .ZN(n8170) );
  NAND2_X1 U8129 ( .A1(n9331), .A2(n7610), .ZN(n9187) );
  NAND2_X1 U8130 ( .A1(n7541), .A2(n9341), .ZN(n7540) );
  INV_X1 U8131 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n7541) );
  XNOR2_X1 U8132 ( .A(n8154), .B(n8153), .ZN(n11595) );
  NOR2_X1 U8133 ( .A1(n9187), .A2(P1_IR_REG_26__SCAN_IN), .ZN(n9188) );
  XNOR2_X1 U8135 ( .A(n8127), .B(n8126), .ZN(n11474) );
  INV_X1 U8136 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n9177) );
  OR2_X1 U8137 ( .A1(n9193), .A2(P1_IR_REG_24__SCAN_IN), .ZN(n9183) );
  OAI21_X1 U8138 ( .B1(n8074), .B2(n7021), .A(n7692), .ZN(n8096) );
  XNOR2_X1 U8139 ( .A(n8096), .B(n8999), .ZN(n11570) );
  AND2_X1 U8140 ( .A1(n9354), .A2(n9335), .ZN(n11534) );
  NAND2_X1 U8141 ( .A1(n7967), .A2(n7665), .ZN(n7983) );
  NAND2_X1 U8142 ( .A1(n7934), .A2(n7657), .ZN(n7951) );
  NAND2_X1 U8143 ( .A1(n7644), .A2(n7643), .ZN(n7882) );
  XNOR2_X1 U8144 ( .A(n7845), .B(n7844), .ZN(n10678) );
  NAND2_X1 U8145 ( .A1(n7308), .A2(n7639), .ZN(n7845) );
  NAND2_X1 U8146 ( .A1(n7833), .A2(n7637), .ZN(n7308) );
  NAND2_X1 U8147 ( .A1(n7302), .A2(n6575), .ZN(n7303) );
  INV_X1 U8148 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n9164) );
  CLKBUF_X1 U8149 ( .A(n9364), .Z(n9403) );
  INV_X1 U8150 ( .A(n14293), .ZN(n6737) );
  NAND2_X1 U8151 ( .A1(n14376), .A2(n14375), .ZN(n7038) );
  OAI21_X1 U8152 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(n14271), .A(n14270), .ZN(
        n14287) );
  OAI21_X1 U8153 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(n14274), .A(n14273), .ZN(
        n14330) );
  INV_X1 U8154 ( .A(n14580), .ZN(n7028) );
  AOI22_X1 U8155 ( .A1(P3_ADDR_REG_13__SCAN_IN), .A2(n14279), .B1(n14286), 
        .B2(n14278), .ZN(n14332) );
  INV_X1 U8156 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n14412) );
  NAND2_X1 U8157 ( .A1(n8711), .A2(n8712), .ZN(n9853) );
  NAND2_X1 U8158 ( .A1(n10107), .A2(n6883), .ZN(n10274) );
  NAND2_X1 U8159 ( .A1(n8742), .A2(n6884), .ZN(n6883) );
  INV_X1 U8160 ( .A(n15037), .ZN(n6884) );
  INV_X1 U8161 ( .A(n12947), .ZN(n12491) );
  AND3_X1 U8162 ( .A1(n8994), .A2(n8993), .A3(n8992), .ZN(n12504) );
  NAND2_X1 U8163 ( .A1(n8943), .A2(n8942), .ZN(n12909) );
  NAND2_X1 U8164 ( .A1(n9107), .A2(n12868), .ZN(n12524) );
  OR2_X1 U8165 ( .A1(n6525), .A2(n8723), .ZN(n8724) );
  XNOR2_X1 U8166 ( .A(n8672), .B(P3_IR_REG_6__SCAN_IN), .ZN(n14986) );
  NAND2_X1 U8167 ( .A1(n6821), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n6822) );
  INV_X1 U8168 ( .A(n12562), .ZN(n6821) );
  NAND2_X1 U8169 ( .A1(n6749), .A2(n6816), .ZN(n6815) );
  NAND2_X1 U8170 ( .A1(n6742), .A2(n6741), .ZN(n12703) );
  INV_X1 U8171 ( .A(n12682), .ZN(n6741) );
  INV_X1 U8172 ( .A(n6742), .ZN(n12683) );
  INV_X1 U8173 ( .A(n7114), .ZN(n12669) );
  INV_X1 U8174 ( .A(n6828), .ZN(n6827) );
  AOI21_X1 U8175 ( .B1(n12686), .B2(n15015), .A(n12685), .ZN(n6828) );
  NAND2_X1 U8176 ( .A1(n12706), .A2(n15015), .ZN(n7278) );
  INV_X1 U8177 ( .A(n12697), .ZN(n6807) );
  INV_X1 U8178 ( .A(n12705), .ZN(n7277) );
  XNOR2_X1 U8179 ( .A(n7281), .B(n12704), .ZN(n7280) );
  NAND2_X1 U8180 ( .A1(n12703), .A2(n12702), .ZN(n7281) );
  XNOR2_X1 U8181 ( .A(n12718), .B(n12717), .ZN(n12874) );
  NAND2_X1 U8182 ( .A1(n7156), .A2(n7154), .ZN(n12718) );
  NOR2_X1 U8183 ( .A1(n7155), .A2(n12716), .ZN(n7154) );
  AND2_X1 U8184 ( .A1(n12725), .A2(n12724), .ZN(n12875) );
  NAND2_X1 U8185 ( .A1(n9017), .A2(n9016), .ZN(n12789) );
  NAND2_X1 U8186 ( .A1(n8902), .A2(n8901), .ZN(n12918) );
  NAND2_X1 U8187 ( .A1(n8888), .A2(n8887), .ZN(n12922) );
  NAND2_X1 U8188 ( .A1(n11826), .A2(n11825), .ZN(n12932) );
  AND2_X2 U8189 ( .A1(n9943), .A2(n9942), .ZN(n15131) );
  AND2_X1 U8190 ( .A1(n7551), .A2(n15110), .ZN(n7549) );
  INV_X1 U8191 ( .A(n7549), .ZN(n7548) );
  OAI21_X1 U8192 ( .B1(n12874), .B2(n12889), .A(n12875), .ZN(n12931) );
  NAND2_X1 U8193 ( .A1(n12932), .A2(n12988), .ZN(n7169) );
  NAND2_X1 U8194 ( .A1(n9001), .A2(n9000), .ZN(n12958) );
  NAND2_X1 U8195 ( .A1(n8958), .A2(n8957), .ZN(n12979) );
  AND2_X1 U8196 ( .A1(n15110), .A2(n14441), .ZN(n12988) );
  AND2_X1 U8197 ( .A1(n9072), .A2(n9071), .ZN(n13001) );
  OR2_X1 U8198 ( .A1(n11870), .A2(n6672), .ZN(n7369) );
  NAND2_X1 U8199 ( .A1(n8047), .A2(n8046), .ZN(n13516) );
  NOR2_X1 U8200 ( .A1(n7383), .A2(n14474), .ZN(n7381) );
  AND2_X1 U8201 ( .A1(n7385), .A2(n7388), .ZN(n7383) );
  NAND2_X1 U8202 ( .A1(n7385), .A2(n7389), .ZN(n7384) );
  OR2_X1 U8203 ( .A1(n7390), .A2(n13038), .ZN(n7389) );
  INV_X1 U8204 ( .A(n13068), .ZN(n7390) );
  OR2_X1 U8205 ( .A1(n13034), .A2(n13035), .ZN(n6935) );
  NAND2_X1 U8206 ( .A1(n13104), .A2(n9287), .ZN(n9295) );
  NAND2_X1 U8207 ( .A1(n7939), .A2(n7938), .ZN(n14516) );
  NAND2_X1 U8208 ( .A1(n7377), .A2(n7376), .ZN(n14476) );
  INV_X1 U8209 ( .A(n14472), .ZN(n7376) );
  INV_X1 U8210 ( .A(n14473), .ZN(n7377) );
  AND2_X1 U8211 ( .A1(n11435), .A2(n7379), .ZN(n7378) );
  NAND2_X1 U8212 ( .A1(n14472), .A2(n9270), .ZN(n7379) );
  NAND2_X1 U8213 ( .A1(n14473), .A2(n9270), .ZN(n7372) );
  NAND2_X1 U8214 ( .A1(n8027), .A2(n8026), .ZN(n14498) );
  NAND2_X1 U8215 ( .A1(n8065), .A2(n8064), .ZN(n13511) );
  NAND2_X1 U8216 ( .A1(n8033), .A2(n8032), .ZN(n13521) );
  NAND2_X1 U8217 ( .A1(n9297), .A2(n14877), .ZN(n14479) );
  NAND2_X1 U8218 ( .A1(n8556), .A2(n8554), .ZN(n8555) );
  INV_X1 U8219 ( .A(n11796), .ZN(n8589) );
  OR2_X1 U8220 ( .A1(n8488), .A2(n9545), .ZN(n7771) );
  OAI21_X1 U8221 ( .B1(n13167), .B2(n13178), .A(n9531), .ZN(n13183) );
  AOI21_X1 U8222 ( .B1(P2_REG1_REG_3__SCAN_IN), .B2(n13184), .A(n13174), .ZN(
        n9574) );
  AND2_X1 U8223 ( .A1(n11027), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n6962) );
  OAI21_X1 U8224 ( .B1(n14845), .B2(n14844), .A(n14843), .ZN(n14847) );
  XNOR2_X1 U8225 ( .A(n6570), .B(n6780), .ZN(n13226) );
  INV_X1 U8226 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n6780) );
  AND2_X1 U8227 ( .A1(n9542), .A2(n9550), .ZN(n14870) );
  AND2_X1 U8228 ( .A1(n6945), .A2(n6946), .ZN(n13225) );
  NAND2_X1 U8229 ( .A1(n6556), .A2(n13316), .ZN(n13450) );
  AOI21_X1 U8230 ( .B1(n13456), .B2(n13444), .A(n8294), .ZN(n8295) );
  NAND2_X1 U8231 ( .A1(n8114), .A2(n8113), .ZN(n13486) );
  AND2_X1 U8232 ( .A1(n8553), .A2(n14491), .ZN(n14883) );
  NAND3_X2 U8233 ( .A1(n7758), .A2(n7759), .A3(n7397), .ZN(n10824) );
  OR2_X1 U8234 ( .A1(n7791), .A2(n9474), .ZN(n7758) );
  OR2_X1 U8235 ( .A1(n7800), .A2(n9478), .ZN(n7397) );
  AND2_X1 U8236 ( .A1(n13450), .A2(n13452), .ZN(n13541) );
  OAI21_X1 U8237 ( .B1(n13463), .B2(n13519), .A(n7472), .ZN(n13548) );
  AND2_X1 U8238 ( .A1(n7204), .A2(n6655), .ZN(n7472) );
  NAND2_X1 U8239 ( .A1(n8217), .A2(n8216), .ZN(n14890) );
  NOR2_X1 U8240 ( .A1(n11348), .A2(n14249), .ZN(n7260) );
  OR3_X1 U8241 ( .A1(n13683), .A2(n13655), .A3(n13654), .ZN(n13656) );
  NAND2_X1 U8242 ( .A1(n7226), .A2(n7230), .ZN(n13657) );
  NAND2_X1 U8243 ( .A1(n13686), .A2(n7232), .ZN(n7226) );
  NAND2_X1 U8244 ( .A1(n14159), .A2(n14533), .ZN(n6795) );
  NAND2_X1 U8245 ( .A1(n11485), .A2(n11484), .ZN(n14165) );
  NAND2_X1 U8246 ( .A1(n9436), .A2(n9435), .ZN(n13727) );
  NAND2_X1 U8247 ( .A1(n9447), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14542) );
  INV_X1 U8248 ( .A(n13727), .ZN(n14535) );
  AND2_X1 U8249 ( .A1(n10294), .A2(n14221), .ZN(n14537) );
  OR2_X1 U8250 ( .A1(n11600), .A2(n9396), .ZN(n9400) );
  OR2_X1 U8251 ( .A1(n12325), .A2(n9597), .ZN(n9398) );
  OR2_X1 U8252 ( .A1(n11600), .A2(n9378), .ZN(n9381) );
  OR2_X1 U8253 ( .A1(n6539), .A2(n9387), .ZN(n9379) );
  NAND2_X1 U8254 ( .A1(n6733), .A2(n6732), .ZN(n9643) );
  NAND2_X1 U8255 ( .A1(n9652), .A2(n9596), .ZN(n6732) );
  OR2_X1 U8256 ( .A1(n9652), .A2(n9596), .ZN(n6733) );
  INV_X1 U8257 ( .A(n13869), .ZN(n6710) );
  OAI21_X1 U8258 ( .B1(n14624), .B2(n7616), .A(n13872), .ZN(n6709) );
  XOR2_X1 U8259 ( .A(n13921), .B(n13918), .Z(n14144) );
  AND2_X1 U8260 ( .A1(n6698), .A2(n13919), .ZN(n14141) );
  NAND2_X1 U8261 ( .A1(n13920), .A2(n13921), .ZN(n6698) );
  NAND2_X1 U8262 ( .A1(n13890), .A2(n7015), .ZN(n13920) );
  NAND2_X1 U8263 ( .A1(n11573), .A2(n10677), .ZN(n6831) );
  NAND2_X1 U8264 ( .A1(n11551), .A2(n11550), .ZN(n14029) );
  NAND2_X1 U8265 ( .A1(n11310), .A2(n11309), .ZN(n14534) );
  AND2_X1 U8266 ( .A1(n14146), .A2(n14148), .ZN(n6776) );
  NAND2_X1 U8267 ( .A1(n14386), .A2(P2_ADDR_REG_9__SCAN_IN), .ZN(n7033) );
  NAND2_X1 U8268 ( .A1(n14328), .A2(n14842), .ZN(n7030) );
  NAND2_X1 U8269 ( .A1(n6736), .A2(n6735), .ZN(n7025) );
  INV_X1 U8270 ( .A(n14597), .ZN(n6735) );
  AND3_X1 U8271 ( .A1(n12168), .A2(n12167), .A3(n12166), .ZN(n12169) );
  AOI21_X1 U8272 ( .B1(n7753), .B2(n8302), .A(n8308), .ZN(n8318) );
  NAND2_X1 U8273 ( .A1(n6584), .A2(n8353), .ZN(n8358) );
  INV_X1 U8274 ( .A(n12215), .ZN(n7068) );
  NAND2_X1 U8275 ( .A1(n7585), .A2(n7587), .ZN(n7584) );
  INV_X1 U8276 ( .A(n8376), .ZN(n7585) );
  INV_X1 U8277 ( .A(n7584), .ZN(n6974) );
  NAND2_X1 U8278 ( .A1(n7611), .A2(n8372), .ZN(n8377) );
  AND2_X1 U8279 ( .A1(n8375), .A2(n8376), .ZN(n7586) );
  NAND2_X1 U8280 ( .A1(n12220), .A2(n12221), .ZN(n12219) );
  AOI21_X1 U8281 ( .B1(n7579), .B2(n7577), .A(n6624), .ZN(n7575) );
  AND2_X1 U8282 ( .A1(n12255), .A2(n7051), .ZN(n7050) );
  NAND2_X1 U8283 ( .A1(n7054), .A2(n7052), .ZN(n7051) );
  INV_X1 U8284 ( .A(n7055), .ZN(n7052) );
  INV_X1 U8285 ( .A(n7054), .ZN(n7053) );
  INV_X1 U8286 ( .A(n7050), .ZN(n7046) );
  NAND2_X1 U8287 ( .A1(n6970), .A2(n6969), .ZN(n8396) );
  AND2_X1 U8288 ( .A1(n7577), .A2(n6624), .ZN(n6969) );
  INV_X1 U8289 ( .A(n8400), .ZN(n7598) );
  INV_X1 U8290 ( .A(n7048), .ZN(n7047) );
  AOI21_X1 U8291 ( .B1(n7591), .B2(n7590), .A(n6619), .ZN(n7589) );
  NAND2_X1 U8292 ( .A1(n8412), .A2(n8411), .ZN(n8416) );
  NAND2_X1 U8293 ( .A1(n6577), .A2(n7592), .ZN(n7590) );
  NOR2_X1 U8294 ( .A1(n6577), .A2(n7592), .ZN(n7591) );
  NOR2_X1 U8295 ( .A1(n8431), .A2(n6992), .ZN(n6991) );
  NAND2_X1 U8296 ( .A1(n6995), .A2(n6994), .ZN(n6992) );
  NAND2_X1 U8297 ( .A1(n6995), .A2(n6994), .ZN(n6993) );
  NAND2_X1 U8298 ( .A1(n7072), .A2(n12274), .ZN(n7071) );
  NAND2_X1 U8299 ( .A1(n7596), .A2(n7593), .ZN(n8442) );
  NAND2_X1 U8300 ( .A1(n7595), .A2(n7594), .ZN(n7593) );
  INV_X1 U8301 ( .A(n8435), .ZN(n7595) );
  NAND2_X1 U8302 ( .A1(n7063), .A2(n12284), .ZN(n7062) );
  INV_X1 U8303 ( .A(n12285), .ZN(n7063) );
  NAND2_X1 U8304 ( .A1(n11951), .A2(n12095), .ZN(n7337) );
  NAND2_X1 U8305 ( .A1(n7339), .A2(n6529), .ZN(n7338) );
  OAI21_X1 U8306 ( .B1(n12772), .B2(n11950), .A(n11949), .ZN(n7339) );
  NAND2_X1 U8307 ( .A1(n8450), .A2(n8451), .ZN(n7560) );
  NAND2_X1 U8308 ( .A1(n7572), .A2(n7574), .ZN(n7571) );
  INV_X1 U8309 ( .A(n8461), .ZN(n7572) );
  AND2_X1 U8310 ( .A1(n8460), .A2(n8461), .ZN(n7573) );
  INV_X1 U8311 ( .A(n12305), .ZN(n7297) );
  NOR2_X1 U8312 ( .A1(n12309), .A2(n12307), .ZN(n6843) );
  INV_X1 U8313 ( .A(n8019), .ZN(n7005) );
  INV_X1 U8314 ( .A(n7653), .ZN(n7318) );
  INV_X1 U8315 ( .A(n8968), .ZN(n6889) );
  NOR2_X1 U8316 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n7714) );
  INV_X1 U8317 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n7718) );
  INV_X1 U8318 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n7719) );
  AND2_X1 U8319 ( .A1(n7291), .A2(n6842), .ZN(n6841) );
  NAND2_X1 U8320 ( .A1(n12307), .A2(n12309), .ZN(n6842) );
  NAND2_X1 U8321 ( .A1(n12312), .A2(n7292), .ZN(n7291) );
  INV_X1 U8322 ( .A(n12314), .ZN(n7292) );
  AND3_X1 U8323 ( .A1(n9175), .A2(n9174), .A3(n9173), .ZN(n9180) );
  INV_X1 U8324 ( .A(n7020), .ZN(n7019) );
  AOI21_X1 U8325 ( .B1(n7020), .B2(n7018), .A(n7017), .ZN(n7016) );
  AOI21_X1 U8326 ( .B1(n7021), .B2(n7692), .A(n7694), .ZN(n7020) );
  AOI21_X1 U8327 ( .B1(n7609), .B2(n7301), .A(n7300), .ZN(n7299) );
  INV_X1 U8328 ( .A(n7657), .ZN(n7301) );
  INV_X1 U8329 ( .A(n7661), .ZN(n7300) );
  AND2_X1 U8330 ( .A1(n7319), .A2(n7318), .ZN(n7317) );
  NAND2_X1 U8331 ( .A1(n7317), .A2(n7860), .ZN(n7010) );
  OAI21_X1 U8332 ( .B1(n14301), .B2(P1_ADDR_REG_3__SCAN_IN), .A(n6630), .ZN(
        n6802) );
  INV_X1 U8333 ( .A(P3_ADDR_REG_4__SCAN_IN), .ZN(n14258) );
  NAND2_X1 U8334 ( .A1(n12499), .A2(n9013), .ZN(n9019) );
  NAND2_X1 U8335 ( .A1(n12082), .A2(n7359), .ZN(n7358) );
  AND2_X1 U8336 ( .A1(n12081), .A2(n12095), .ZN(n7359) );
  NAND2_X1 U8337 ( .A1(n7285), .A2(n7284), .ZN(n7283) );
  AND2_X1 U8338 ( .A1(n7116), .A2(n7115), .ZN(n9782) );
  AND2_X1 U8339 ( .A1(n6825), .A2(n6824), .ZN(n10078) );
  NAND2_X1 U8340 ( .A1(n14358), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n6824) );
  NAND2_X1 U8341 ( .A1(n6823), .A2(n6674), .ZN(n10082) );
  OR2_X1 U8342 ( .A1(n14975), .A2(n6551), .ZN(n7125) );
  OR2_X1 U8343 ( .A1(n10085), .A2(n10084), .ZN(n7271) );
  NAND2_X1 U8344 ( .A1(n6713), .A2(n6682), .ZN(n11087) );
  INV_X1 U8345 ( .A(n11127), .ZN(n7122) );
  XNOR2_X1 U8346 ( .A(n6746), .B(n12693), .ZN(n12674) );
  NAND2_X1 U8347 ( .A1(n14434), .A2(n11298), .ZN(n7515) );
  OR2_X1 U8348 ( .A1(n12932), .A2(n12736), .ZN(n12089) );
  NAND2_X1 U8349 ( .A1(n12814), .A2(n7519), .ZN(n7518) );
  INV_X1 U8350 ( .A(n7521), .ZN(n7519) );
  NOR2_X1 U8351 ( .A1(n7141), .A2(n7138), .ZN(n7137) );
  INV_X1 U8352 ( .A(n12849), .ZN(n7141) );
  OR2_X1 U8353 ( .A1(n12909), .A2(n11804), .ZN(n11958) );
  AND2_X1 U8354 ( .A1(n11963), .A2(n12055), .ZN(n12050) );
  NAND2_X1 U8355 ( .A1(n14432), .A2(n12030), .ZN(n7163) );
  INV_X1 U8356 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n7435) );
  AND2_X1 U8357 ( .A1(n10672), .A2(P1_DATAO_REG_19__SCAN_IN), .ZN(n6805) );
  INV_X1 U8358 ( .A(n8969), .ZN(n7346) );
  INV_X1 U8359 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n8843) );
  INV_X1 U8360 ( .A(n7362), .ZN(n7361) );
  AOI21_X1 U8361 ( .B1(n7364), .B2(n7363), .A(n6685), .ZN(n7362) );
  NOR2_X1 U8362 ( .A1(n8815), .A2(P3_IR_REG_10__SCAN_IN), .ZN(n8826) );
  NAND2_X1 U8363 ( .A1(n8696), .A2(n7102), .ZN(n7103) );
  NAND2_X1 U8364 ( .A1(n8473), .A2(n7558), .ZN(n7557) );
  INV_X1 U8365 ( .A(n7740), .ZN(n7170) );
  OR2_X1 U8366 ( .A1(n7740), .A2(n10822), .ZN(n7475) );
  NOR2_X1 U8367 ( .A1(n13469), .A2(n13474), .ZN(n6916) );
  INV_X1 U8368 ( .A(n8072), .ZN(n7459) );
  INV_X1 U8369 ( .A(n8262), .ZN(n7210) );
  NOR2_X1 U8370 ( .A1(n13425), .A2(n14498), .ZN(n7406) );
  INV_X1 U8371 ( .A(n10851), .ZN(n6810) );
  INV_X1 U8372 ( .A(n8241), .ZN(n7184) );
  INV_X1 U8373 ( .A(n8239), .ZN(n7187) );
  AND2_X1 U8374 ( .A1(n10484), .A2(n10731), .ZN(n8242) );
  INV_X1 U8375 ( .A(n8231), .ZN(n7177) );
  NAND2_X1 U8376 ( .A1(n13325), .A2(n13314), .ZN(n13317) );
  NAND2_X1 U8377 ( .A1(n6646), .A2(n8043), .ZN(n7396) );
  AND2_X1 U8378 ( .A1(n7717), .A2(n7716), .ZN(n7819) );
  AND2_X1 U8379 ( .A1(n13740), .A2(n13660), .ZN(n7244) );
  NOR2_X1 U8380 ( .A1(n11554), .A2(n13637), .ZN(n11561) );
  NAND2_X1 U8381 ( .A1(n13808), .A2(n13807), .ZN(n13809) );
  NAND2_X1 U8382 ( .A1(n6554), .A2(n6625), .ZN(n7087) );
  NAND2_X1 U8383 ( .A1(n6516), .A2(n6734), .ZN(n11630) );
  NOR2_X1 U8384 ( .A1(n7267), .A2(n14153), .ZN(n6734) );
  NAND2_X1 U8385 ( .A1(n13950), .A2(n7268), .ZN(n7267) );
  NOR2_X1 U8386 ( .A1(n14165), .A2(n13981), .ZN(n7268) );
  AND2_X1 U8387 ( .A1(n7083), .A2(n12353), .ZN(n7082) );
  OR2_X1 U8388 ( .A1(n12350), .A2(n7084), .ZN(n7083) );
  INV_X1 U8389 ( .A(n11197), .ZN(n7084) );
  OR2_X1 U8390 ( .A1(n7263), .A2(n12225), .ZN(n7262) );
  NAND2_X1 U8391 ( .A1(n14393), .A2(n14557), .ZN(n7263) );
  NAND2_X1 U8392 ( .A1(n7682), .A2(SI_18_), .ZN(n7683) );
  INV_X1 U8393 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n9170) );
  INV_X1 U8394 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n9169) );
  NAND2_X1 U8395 ( .A1(n7314), .A2(n7664), .ZN(n7967) );
  INV_X1 U8396 ( .A(n7965), .ZN(n7314) );
  AND2_X1 U8397 ( .A1(n7657), .A2(n7656), .ZN(n7931) );
  NAND2_X1 U8398 ( .A1(n7932), .A2(n7931), .ZN(n7934) );
  NOR2_X1 U8399 ( .A1(n9586), .A2(n9585), .ZN(n9693) );
  AOI21_X1 U8400 ( .B1(n7309), .B2(n7310), .A(n6634), .ZN(n7306) );
  INV_X1 U8401 ( .A(n7639), .ZN(n7310) );
  OAI21_X1 U8402 ( .B1(n9475), .B2(P2_DATAO_REG_3__SCAN_IN), .A(n6814), .ZN(
        n7627) );
  OR2_X1 U8403 ( .A1(n7626), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n6814) );
  INV_X1 U8404 ( .A(P2_RD_REG_SCAN_IN), .ZN(n6997) );
  INV_X1 U8405 ( .A(P1_RD_REG_SCAN_IN), .ZN(n7615) );
  AOI21_X1 U8406 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(n14269), .A(n14268), .ZN(
        n14321) );
  AND2_X1 U8407 ( .A1(n12123), .A2(n12122), .ZN(n12388) );
  OR2_X1 U8408 ( .A1(n9019), .A2(n9018), .ZN(n6894) );
  INV_X1 U8409 ( .A(P3_REG3_REG_10__SCAN_IN), .ZN(n8611) );
  AND2_X1 U8410 ( .A1(n9140), .A2(n9064), .ZN(n9066) );
  INV_X1 U8411 ( .A(n6863), .ZN(n6862) );
  OAI21_X1 U8412 ( .B1(n6553), .B2(n6864), .A(n7601), .ZN(n6863) );
  INV_X1 U8413 ( .A(n8910), .ZN(n6864) );
  NOR2_X1 U8414 ( .A1(n8759), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n8796) );
  OR3_X1 U8415 ( .A1(n8831), .A2(P3_REG3_REG_12__SCAN_IN), .A3(
        P3_REG3_REG_11__SCAN_IN), .ZN(n8855) );
  NAND2_X1 U8416 ( .A1(n8710), .A2(n7482), .ZN(n8712) );
  AOI21_X1 U8417 ( .B1(n10274), .B2(n10273), .A(n6882), .ZN(n12521) );
  AND2_X1 U8418 ( .A1(n8757), .A2(n10111), .ZN(n6882) );
  NAND2_X1 U8419 ( .A1(n12521), .A2(n12520), .ZN(n12519) );
  OR2_X1 U8420 ( .A1(n8889), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n8903) );
  INV_X1 U8421 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n15380) );
  INV_X1 U8422 ( .A(P3_ADDR_REG_1__SCAN_IN), .ZN(n15350) );
  OR2_X1 U8423 ( .A1(n9809), .A2(n9808), .ZN(n7285) );
  XNOR2_X1 U8424 ( .A(n9782), .B(n14952), .ZN(n14942) );
  XNOR2_X1 U8425 ( .A(n7283), .B(n7282), .ZN(n14940) );
  XNOR2_X1 U8426 ( .A(n10078), .B(n14966), .ZN(n14961) );
  INV_X1 U8427 ( .A(n7105), .ZN(n10068) );
  NAND2_X1 U8428 ( .A1(n10072), .A2(n7125), .ZN(n14994) );
  INV_X1 U8429 ( .A(P3_IR_REG_6__SCAN_IN), .ZN(n8656) );
  INV_X1 U8430 ( .A(n7271), .ZN(n10652) );
  OAI22_X1 U8431 ( .A1(n11093), .A2(n11092), .B1(n11091), .B2(n11090), .ZN(
        n15012) );
  NAND2_X1 U8432 ( .A1(n7123), .A2(n11096), .ZN(n7121) );
  INV_X1 U8433 ( .A(n11087), .ZN(n7123) );
  INV_X1 U8434 ( .A(n11126), .ZN(n7118) );
  INV_X1 U8435 ( .A(n11125), .ZN(n7119) );
  NAND2_X1 U8436 ( .A1(n7107), .A2(n7108), .ZN(n12572) );
  INV_X1 U8437 ( .A(n12582), .ZN(n7109) );
  OR2_X1 U8438 ( .A1(n8885), .A2(P3_IR_REG_14__SCAN_IN), .ZN(n8899) );
  INV_X1 U8439 ( .A(n12618), .ZN(n6816) );
  NAND2_X1 U8440 ( .A1(n12589), .A2(n6818), .ZN(n6817) );
  AND2_X1 U8441 ( .A1(n12632), .A2(n6749), .ZN(n6806) );
  NAND2_X1 U8442 ( .A1(n14384), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n7127) );
  INV_X1 U8443 ( .A(n6746), .ZN(n12696) );
  OR2_X1 U8444 ( .A1(n13011), .A2(n11896), .ZN(n11898) );
  INV_X1 U8445 ( .A(n7158), .ZN(n7155) );
  INV_X1 U8446 ( .A(n12717), .ZN(n12720) );
  NAND2_X1 U8447 ( .A1(n12747), .A2(n12081), .ZN(n7157) );
  INV_X1 U8448 ( .A(n9054), .ZN(n9053) );
  OR2_X1 U8449 ( .A1(n7496), .A2(n7493), .ZN(n7492) );
  INV_X1 U8450 ( .A(n11812), .ZN(n7493) );
  INV_X1 U8451 ( .A(n12757), .ZN(n12760) );
  NAND2_X1 U8452 ( .A1(n12760), .A2(n12759), .ZN(n12758) );
  AND2_X1 U8453 ( .A1(n12084), .A2(n12080), .ZN(n12757) );
  OR2_X1 U8454 ( .A1(n8974), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n8990) );
  OR2_X1 U8455 ( .A1(n8959), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n8974) );
  NAND2_X1 U8456 ( .A1(n8944), .A2(n12513), .ZN(n8959) );
  AND2_X1 U8457 ( .A1(n8926), .A2(n8925), .ZN(n8944) );
  NOR2_X1 U8458 ( .A1(n8903), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n8926) );
  INV_X1 U8459 ( .A(n12549), .ZN(n12865) );
  INV_X1 U8460 ( .A(P3_REG3_REG_14__SCAN_IN), .ZN(n12403) );
  NAND2_X1 U8461 ( .A1(n8873), .A2(n12403), .ZN(n8889) );
  NOR2_X1 U8462 ( .A1(n8855), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n8873) );
  NAND2_X1 U8463 ( .A1(n8798), .A2(n8611), .ZN(n8831) );
  AOI21_X1 U8464 ( .B1(n12003), .B2(n7133), .A(n12005), .ZN(n7132) );
  INV_X1 U8465 ( .A(n12001), .ZN(n7133) );
  NOR2_X1 U8466 ( .A1(n11928), .A2(n7487), .ZN(n7486) );
  INV_X1 U8467 ( .A(n10614), .ZN(n7487) );
  NAND2_X1 U8468 ( .A1(n10615), .A2(n10614), .ZN(n10616) );
  NAND2_X1 U8469 ( .A1(n10035), .A2(n11973), .ZN(n10094) );
  INV_X1 U8470 ( .A(n10611), .ZN(n9937) );
  NAND2_X1 U8471 ( .A1(n11821), .A2(n11820), .ZN(n12118) );
  AND2_X1 U8472 ( .A1(n12081), .A2(n12085), .ZN(n12748) );
  INV_X1 U8473 ( .A(n12803), .ZN(n12805) );
  AND2_X1 U8474 ( .A1(n12070), .A2(n12071), .ZN(n12803) );
  AND2_X1 U8475 ( .A1(n8972), .A2(n8971), .ZN(n11807) );
  NAND2_X1 U8476 ( .A1(n6717), .A2(n6716), .ZN(n12842) );
  INV_X1 U8477 ( .A(n15099), .ZN(n14441) );
  AOI21_X1 U8478 ( .B1(n7510), .B2(n7508), .A(n6613), .ZN(n7507) );
  INV_X1 U8479 ( .A(n7510), .ZN(n7509) );
  OR2_X1 U8480 ( .A1(n9861), .A2(n9092), .ZN(n9930) );
  AND2_X1 U8481 ( .A1(n9723), .A2(P3_STATE_REG_SCAN_IN), .ZN(n9856) );
  AND2_X1 U8482 ( .A1(n15197), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n6804) );
  NOR2_X1 U8483 ( .A1(n8625), .A2(n8624), .ZN(n9096) );
  INV_X1 U8484 ( .A(n8653), .ZN(n8624) );
  INV_X1 U8485 ( .A(n9014), .ZN(n7355) );
  AOI21_X1 U8486 ( .B1(n7333), .B2(n8895), .A(n6686), .ZN(n7332) );
  AND2_X1 U8487 ( .A1(n8845), .A2(n8844), .ZN(n8850) );
  AND2_X1 U8488 ( .A1(n8826), .A2(n8825), .ZN(n8845) );
  OR2_X1 U8489 ( .A1(n8791), .A2(P3_IR_REG_9__SCAN_IN), .ZN(n8815) );
  XNOR2_X1 U8490 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .ZN(n8810) );
  AOI21_X1 U8491 ( .B1(n7343), .B2(n7345), .A(n6641), .ZN(n7341) );
  XNOR2_X1 U8492 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(P2_DATAO_REG_9__SCAN_IN), 
        .ZN(n8789) );
  AOI21_X1 U8493 ( .B1(n7325), .B2(n8743), .A(n6642), .ZN(n7324) );
  INV_X1 U8494 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n8847) );
  NAND2_X1 U8495 ( .A1(n8637), .A2(n8636), .ZN(n8716) );
  INV_X1 U8496 ( .A(n10343), .ZN(n6928) );
  INV_X1 U8497 ( .A(n9224), .ZN(n6929) );
  OR2_X1 U8498 ( .A1(n7922), .A2(n7921), .ZN(n7941) );
  NAND2_X1 U8499 ( .A1(n7988), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8009) );
  OR2_X1 U8500 ( .A1(n8009), .A2(n8008), .ZN(n8015) );
  INV_X1 U8501 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n7823) );
  OR2_X1 U8502 ( .A1(n7370), .A2(n6576), .ZN(n7368) );
  OR2_X1 U8503 ( .A1(n13089), .A2(n6672), .ZN(n6941) );
  NAND2_X1 U8504 ( .A1(n6936), .A2(n6939), .ZN(n6938) );
  INV_X1 U8505 ( .A(n13089), .ZN(n6939) );
  INV_X1 U8506 ( .A(n7368), .ZN(n6936) );
  NOR2_X1 U8507 ( .A1(n8116), .A2(n8115), .ZN(n8132) );
  NOR2_X1 U8508 ( .A1(n7941), .A2(n7940), .ZN(n7973) );
  NOR2_X1 U8509 ( .A1(n8015), .A2(n11432), .ZN(n8034) );
  OR2_X1 U8510 ( .A1(n14473), .A2(n7375), .ZN(n6926) );
  NAND2_X1 U8511 ( .A1(n10353), .A2(n7391), .ZN(n10266) );
  NAND2_X1 U8512 ( .A1(n7769), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n7770) );
  MUX2_X1 U8513 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n15291), .S(n13162), .Z(
        n13169) );
  AND2_X1 U8514 ( .A1(n13176), .A2(n13177), .ZN(n13174) );
  OAI21_X1 U8515 ( .B1(n9661), .B2(n9660), .A(n9659), .ZN(n9658) );
  AOI21_X1 U8516 ( .B1(n11026), .B2(P2_REG2_REG_10__SCAN_IN), .A(n11025), .ZN(
        n14830) );
  AND2_X1 U8517 ( .A1(n14830), .A2(n14831), .ZN(n14845) );
  OR2_X1 U8518 ( .A1(n7984), .A2(P2_IR_REG_14__SCAN_IN), .ZN(n8000) );
  AND2_X1 U8519 ( .A1(n6957), .A2(n6956), .ZN(n11454) );
  NAND2_X1 U8520 ( .A1(n11452), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n6956) );
  OR2_X1 U8521 ( .A1(n14864), .A2(n7990), .ZN(n14861) );
  NAND2_X1 U8522 ( .A1(n6779), .A2(n6778), .ZN(n13215) );
  NOR2_X1 U8523 ( .A1(n13213), .A2(n13214), .ZN(n13221) );
  NOR2_X1 U8524 ( .A1(n13264), .A2(n7443), .ZN(n7442) );
  INV_X1 U8525 ( .A(n7445), .ZN(n7443) );
  NAND2_X1 U8526 ( .A1(n7400), .A2(n7401), .ZN(n13278) );
  INV_X1 U8527 ( .A(n7400), .ZN(n13300) );
  AOI21_X1 U8528 ( .B1(n7451), .B2(n7455), .A(n6557), .ZN(n7450) );
  INV_X1 U8529 ( .A(n7451), .ZN(n7449) );
  AOI21_X1 U8530 ( .B1(n7190), .B2(n7195), .A(n6636), .ZN(n7188) );
  NAND2_X1 U8531 ( .A1(n6906), .A2(n6905), .ZN(n13347) );
  OR2_X1 U8532 ( .A1(n8077), .A2(n7743), .ZN(n8088) );
  NAND2_X1 U8533 ( .A1(n7407), .A2(n7404), .ZN(n13374) );
  NAND2_X1 U8534 ( .A1(n7406), .A2(n7405), .ZN(n13409) );
  AOI21_X1 U8535 ( .B1(n7198), .B2(n7203), .A(n6635), .ZN(n7196) );
  INV_X1 U8536 ( .A(n7406), .ZN(n13426) );
  NAND2_X1 U8537 ( .A1(n13532), .A2(n8253), .ZN(n11336) );
  INV_X1 U8538 ( .A(n8569), .ZN(n13529) );
  AND2_X1 U8539 ( .A1(n7403), .A2(n6912), .ZN(n6910) );
  NOR2_X1 U8540 ( .A1(n11233), .A2(n13441), .ZN(n6912) );
  NAND2_X1 U8541 ( .A1(n6913), .A2(n6911), .ZN(n11230) );
  AND2_X1 U8542 ( .A1(n7403), .A2(n11079), .ZN(n6911) );
  NAND2_X1 U8543 ( .A1(n7403), .A2(n7402), .ZN(n10906) );
  XNOR2_X1 U8544 ( .A(n10860), .B(n10769), .ZN(n10851) );
  NOR2_X1 U8545 ( .A1(n7887), .A2(n7886), .ZN(n7899) );
  INV_X1 U8546 ( .A(n8563), .ZN(n10543) );
  OR2_X1 U8547 ( .A1(n7852), .A2(n7851), .ZN(n7873) );
  OR2_X1 U8548 ( .A1(n7873), .A2(n7872), .ZN(n7887) );
  NAND2_X1 U8549 ( .A1(n7181), .A2(n8241), .ZN(n10730) );
  NAND2_X1 U8550 ( .A1(n8240), .A2(n7185), .ZN(n7181) );
  INV_X1 U8551 ( .A(n7186), .ZN(n7185) );
  AOI21_X1 U8552 ( .B1(n10185), .B2(n7439), .A(n6621), .ZN(n7438) );
  INV_X1 U8553 ( .A(n7831), .ZN(n7439) );
  NOR2_X1 U8554 ( .A1(n10479), .A2(n10487), .ZN(n6901) );
  NAND2_X1 U8555 ( .A1(n6902), .A2(n6904), .ZN(n10223) );
  NOR2_X1 U8556 ( .A1(n10236), .A2(n10474), .ZN(n10252) );
  INV_X1 U8557 ( .A(n13538), .ZN(n13402) );
  NAND2_X1 U8558 ( .A1(n8484), .A2(n8483), .ZN(n13232) );
  AND2_X1 U8559 ( .A1(n13331), .A2(n13407), .ZN(n13493) );
  NAND2_X1 U8560 ( .A1(n7192), .A2(n7193), .ZN(n13330) );
  OR2_X1 U8561 ( .A1(n13353), .A2(n7195), .ZN(n7192) );
  CLKBUF_X1 U8562 ( .A(n8298), .Z(n14923) );
  INV_X1 U8563 ( .A(n7730), .ZN(n7731) );
  NAND2_X1 U8564 ( .A1(n6900), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7729) );
  NAND2_X1 U8565 ( .A1(n8195), .A2(n8194), .ZN(n8199) );
  OR2_X1 U8566 ( .A1(n7896), .A2(P2_IR_REG_9__SCAN_IN), .ZN(n7916) );
  OR2_X1 U8567 ( .A1(n7936), .A2(P2_IR_REG_6__SCAN_IN), .ZN(n7862) );
  INV_X1 U8568 ( .A(n11562), .ZN(n11578) );
  AND2_X1 U8569 ( .A1(n10984), .A2(n10973), .ZN(n7255) );
  NAND2_X1 U8570 ( .A1(n6745), .A2(n7244), .ZN(n13671) );
  OR2_X1 U8571 ( .A1(n11053), .A2(n11052), .ZN(n11203) );
  NOR2_X1 U8572 ( .A1(n11203), .A2(n11202), .ZN(n11210) );
  NAND2_X1 U8573 ( .A1(n6549), .A2(n6580), .ZN(n7252) );
  AND2_X1 U8574 ( .A1(n6837), .A2(n6836), .ZN(n12379) );
  NAND2_X1 U8575 ( .A1(n12333), .A2(n6838), .ZN(n6836) );
  AND3_X1 U8576 ( .A1(n11559), .A2(n11558), .A3(n11557), .ZN(n13627) );
  AND4_X1 U8577 ( .A1(n11508), .A2(n11507), .A3(n11506), .A4(n11505), .ZN(
        n13746) );
  AOI21_X1 U8578 ( .B1(n9627), .B2(P1_REG1_REG_4__SCAN_IN), .A(n9913), .ZN(
        n9681) );
  AOI21_X1 U8579 ( .B1(P1_REG1_REG_7__SCAN_IN), .B2(n10679), .A(n9821), .ZN(
        n9823) );
  NAND2_X1 U8580 ( .A1(n10791), .A2(n6760), .ZN(n10794) );
  OR2_X1 U8581 ( .A1(n11194), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n6760) );
  AOI21_X1 U8582 ( .B1(n13789), .B2(P1_REG1_REG_13__SCAN_IN), .A(n13788), .ZN(
        n13790) );
  AND2_X1 U8583 ( .A1(n13846), .A2(n13845), .ZN(n13853) );
  NOR2_X1 U8584 ( .A1(n13895), .A2(n13887), .ZN(n13882) );
  NAND2_X1 U8585 ( .A1(n12311), .A2(n12310), .ZN(n13896) );
  NAND2_X1 U8586 ( .A1(n13922), .A2(n14133), .ZN(n13895) );
  INV_X1 U8587 ( .A(n11577), .ZN(n11477) );
  NOR2_X1 U8588 ( .A1(n13992), .A2(n7266), .ZN(n13962) );
  INV_X1 U8589 ( .A(n7268), .ZN(n7266) );
  AOI21_X1 U8590 ( .B1(n13974), .B2(n13976), .A(n6722), .ZN(n13956) );
  AND2_X1 U8591 ( .A1(n13981), .A2(n11618), .ZN(n6722) );
  NOR2_X1 U8592 ( .A1(n14013), .A2(n7078), .ZN(n7077) );
  OAI21_X1 U8593 ( .B1(n14067), .B2(n7096), .A(n7094), .ZN(n14037) );
  AOI21_X1 U8594 ( .B1(n7097), .B2(n7095), .A(n6622), .ZN(n7094) );
  INV_X1 U8595 ( .A(n7097), .ZN(n7096) );
  INV_X1 U8596 ( .A(n11613), .ZN(n7095) );
  OR2_X1 U8597 ( .A1(n11503), .A2(n15369), .ZN(n11523) );
  NOR3_X1 U8598 ( .A1(n11062), .A2(n12225), .A3(n12235), .ZN(n11245) );
  NAND2_X1 U8599 ( .A1(n11047), .A2(n11046), .ZN(n11191) );
  NOR2_X1 U8600 ( .A1(n11062), .A2(n12225), .ZN(n11247) );
  XNOR2_X1 U8601 ( .A(n12225), .B(n11270), .ZN(n12355) );
  OR2_X1 U8602 ( .A1(n10705), .A2(n9747), .ZN(n10877) );
  NOR2_X1 U8603 ( .A1(n10877), .A2(n15304), .ZN(n11005) );
  NAND2_X1 U8604 ( .A1(n10875), .A2(n10694), .ZN(n12346) );
  NAND2_X1 U8605 ( .A1(n6536), .A2(n7261), .ZN(n14636) );
  NAND2_X1 U8606 ( .A1(n6706), .A2(n10299), .ZN(n14653) );
  NAND2_X2 U8607 ( .A1(n6772), .A2(n12143), .ZN(n14663) );
  INV_X1 U8608 ( .A(n9434), .ZN(n6772) );
  INV_X1 U8609 ( .A(n12151), .ZN(n7085) );
  CLKBUF_X1 U8610 ( .A(n12341), .Z(n6726) );
  NAND2_X1 U8611 ( .A1(n6773), .A2(n12144), .ZN(n9434) );
  INV_X1 U8612 ( .A(n13887), .ZN(n14130) );
  NAND2_X1 U8613 ( .A1(n7533), .A2(n7536), .ZN(n13968) );
  NAND2_X1 U8614 ( .A1(n7098), .A2(n7097), .ZN(n14055) );
  NAND2_X1 U8615 ( .A1(n14067), .A2(n11613), .ZN(n7098) );
  NAND2_X1 U8616 ( .A1(n11315), .A2(n11314), .ZN(n11316) );
  INV_X1 U8617 ( .A(n10298), .ZN(n14706) );
  NAND2_X1 U8618 ( .A1(n10526), .A2(n13868), .ZN(n14691) );
  OR2_X1 U8619 ( .A1(n6796), .A2(n14679), .ZN(n14747) );
  AND2_X1 U8620 ( .A1(n14691), .A2(n14747), .ZN(n14724) );
  XNOR2_X1 U8621 ( .A(n8505), .B(n8502), .ZN(n12315) );
  XNOR2_X1 U8622 ( .A(n8479), .B(n8478), .ZN(n12385) );
  XNOR2_X1 U8623 ( .A(n8142), .B(n8141), .ZN(n13593) );
  INV_X1 U8624 ( .A(n12144), .ZN(n14251) );
  XNOR2_X1 U8625 ( .A(n8063), .B(n8062), .ZN(n11548) );
  OAI21_X1 U8626 ( .B1(n7670), .B2(n7009), .A(n7006), .ZN(n8020) );
  INV_X1 U8627 ( .A(n9331), .ZN(n9172) );
  NAND2_X1 U8628 ( .A1(n7670), .A2(n7669), .ZN(n7999) );
  OR2_X1 U8629 ( .A1(n9490), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n9954) );
  OR2_X1 U8630 ( .A1(n9696), .A2(P1_IR_REG_12__SCAN_IN), .ZN(n9846) );
  XNOR2_X1 U8631 ( .A(n7915), .B(n7914), .ZN(n11048) );
  XNOR2_X1 U8632 ( .A(n7861), .B(n7860), .ZN(n10684) );
  XNOR2_X1 U8633 ( .A(n7833), .B(n7832), .ZN(n10400) );
  NAND2_X1 U8634 ( .A1(n9386), .A2(n7304), .ZN(n7754) );
  NAND2_X1 U8635 ( .A1(n7305), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n7304) );
  INV_X1 U8636 ( .A(n8693), .ZN(n7305) );
  NAND2_X1 U8637 ( .A1(n15349), .A2(P3_ADDR_REG_1__SCAN_IN), .ZN(n7036) );
  NAND2_X1 U8638 ( .A1(n6768), .A2(n14303), .ZN(n14306) );
  NOR2_X1 U8639 ( .A1(n14263), .A2(n14262), .ZN(n14309) );
  NOR2_X1 U8640 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n14304), .ZN(n14262) );
  XNOR2_X1 U8641 ( .A(P3_ADDR_REG_7__SCAN_IN), .B(n14264), .ZN(n14313) );
  NOR2_X1 U8642 ( .A1(n14318), .A2(n14319), .ZN(n14322) );
  AOI21_X1 U8643 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(n15030), .A(n14272), .ZN(
        n14327) );
  NOR2_X1 U8644 ( .A1(n14288), .A2(n14287), .ZN(n14272) );
  OAI21_X1 U8645 ( .B1(P3_ADDR_REG_14__SCAN_IN), .B2(n14281), .A(n14280), .ZN(
        n14336) );
  NAND2_X1 U8646 ( .A1(n12519), .A2(n6880), .ZN(n10583) );
  NAND2_X1 U8647 ( .A1(n6881), .A2(n15036), .ZN(n6880) );
  INV_X1 U8648 ( .A(n8758), .ZN(n6881) );
  AOI21_X1 U8649 ( .B1(n11297), .B2(n6869), .A(n6868), .ZN(n6867) );
  NOR2_X1 U8650 ( .A1(n6871), .A2(n11298), .ZN(n6869) );
  AND2_X1 U8651 ( .A1(n9012), .A2(n9011), .ZN(n12414) );
  NAND2_X1 U8652 ( .A1(n10914), .A2(n7431), .ZN(n12420) );
  NAND2_X1 U8653 ( .A1(n10914), .A2(n8807), .ZN(n12419) );
  NAND2_X1 U8654 ( .A1(n7416), .A2(n7417), .ZN(n12430) );
  AND2_X1 U8655 ( .A1(n7416), .A2(n7414), .ZN(n12429) );
  NAND2_X1 U8656 ( .A1(n12509), .A2(n8953), .ZN(n12440) );
  NOR2_X1 U8657 ( .A1(n9853), .A2(n6865), .ZN(n9851) );
  NAND2_X1 U8658 ( .A1(n6866), .A2(n10152), .ZN(n6865) );
  NAND2_X1 U8659 ( .A1(n10035), .A2(n8989), .ZN(n6866) );
  NAND2_X1 U8660 ( .A1(n8982), .A2(n8981), .ZN(n12449) );
  NAND2_X1 U8661 ( .A1(n12493), .A2(n12492), .ZN(n8982) );
  AND2_X1 U8662 ( .A1(n6872), .A2(n6874), .ZN(n11388) );
  OAI21_X1 U8663 ( .B1(n7409), .B2(n6864), .A(n6862), .ZN(n12474) );
  AND2_X1 U8664 ( .A1(n12126), .A2(n12480), .ZN(n12482) );
  NAND2_X1 U8665 ( .A1(n12441), .A2(n8968), .ZN(n12493) );
  NAND2_X1 U8666 ( .A1(n11387), .A2(n8840), .ZN(n11417) );
  NOR2_X1 U8667 ( .A1(n9002), .A2(n6887), .ZN(n7426) );
  INV_X1 U8668 ( .A(n12484), .ZN(n12535) );
  INV_X1 U8669 ( .A(n9144), .ZN(n7425) );
  NAND2_X1 U8670 ( .A1(n12398), .A2(n8881), .ZN(n12531) );
  INV_X1 U8671 ( .A(n12507), .ZN(n12533) );
  NAND2_X1 U8672 ( .A1(n9857), .A2(n12116), .ZN(n12540) );
  NAND2_X1 U8673 ( .A1(n9155), .A2(n9154), .ZN(n12750) );
  INV_X1 U8674 ( .A(n12735), .ZN(n12761) );
  INV_X1 U8675 ( .A(n12414), .ZN(n12807) );
  OR2_X1 U8676 ( .A1(n9195), .A2(n13002), .ZN(n12548) );
  NAND2_X1 U8677 ( .A1(n10144), .A2(P3_REG0_REG_4__SCAN_IN), .ZN(n8684) );
  OR2_X1 U8678 ( .A1(n6525), .A2(n8735), .ZN(n8736) );
  OR2_X1 U8679 ( .A1(n8946), .A2(n8699), .ZN(n8700) );
  INV_X1 U8680 ( .A(P3_ADDR_REG_0__SCAN_IN), .ZN(n14938) );
  INV_X1 U8681 ( .A(P3_ADDR_REG_3__SCAN_IN), .ZN(n14956) );
  INV_X1 U8682 ( .A(n6825), .ZN(n10077) );
  INV_X1 U8683 ( .A(P3_ADDR_REG_6__SCAN_IN), .ZN(n15223) );
  INV_X1 U8684 ( .A(n6823), .ZN(n14979) );
  NOR2_X1 U8685 ( .A1(n10642), .A2(n10643), .ZN(n11085) );
  NAND2_X1 U8686 ( .A1(n7274), .A2(n11119), .ZN(n11103) );
  AND3_X1 U8687 ( .A1(n7121), .A2(n7118), .A3(P3_REG2_REG_11__SCAN_IN), .ZN(
        n11125) );
  NAND2_X1 U8688 ( .A1(n7121), .A2(n7118), .ZN(n11089) );
  AND2_X1 U8689 ( .A1(n7275), .A2(n11119), .ZN(n11123) );
  INV_X1 U8690 ( .A(n12609), .ZN(n12608) );
  OR2_X1 U8691 ( .A1(n12585), .A2(n12584), .ZN(n12621) );
  XNOR2_X1 U8692 ( .A(n12632), .B(n6749), .ZN(n12623) );
  NOR2_X1 U8693 ( .A1(n12623), .A2(n12622), .ZN(n12631) );
  OR2_X1 U8694 ( .A1(n12612), .A2(n15387), .ZN(n7288) );
  OR2_X1 U8695 ( .A1(n12630), .A2(n15387), .ZN(n7286) );
  INV_X1 U8696 ( .A(n6702), .ZN(n12681) );
  INV_X1 U8697 ( .A(n12692), .ZN(n7111) );
  NAND2_X1 U8698 ( .A1(n7512), .A2(n7510), .ZN(n11280) );
  NAND2_X1 U8699 ( .A1(n14433), .A2(n12030), .ZN(n11282) );
  NAND2_X1 U8700 ( .A1(n11180), .A2(n11179), .ZN(n14426) );
  OR2_X1 U8701 ( .A1(n9872), .A2(n11287), .ZN(n11177) );
  NAND2_X1 U8702 ( .A1(n7135), .A2(n12001), .ZN(n10623) );
  NAND2_X1 U8703 ( .A1(n10464), .A2(n11924), .ZN(n7135) );
  NAND2_X1 U8704 ( .A1(n9934), .A2(n9106), .ZN(n12868) );
  AND2_X1 U8705 ( .A1(n7151), .A2(n7150), .ZN(n10155) );
  NAND2_X1 U8706 ( .A1(n7550), .A2(n7551), .ZN(n12709) );
  AND2_X1 U8707 ( .A1(n15131), .A2(n14441), .ZN(n12913) );
  NAND2_X1 U8708 ( .A1(n7328), .A2(n9032), .ZN(n12947) );
  NAND2_X1 U8709 ( .A1(n11275), .A2(n11913), .ZN(n7328) );
  NAND2_X1 U8710 ( .A1(n12783), .A2(n7496), .ZN(n12771) );
  INV_X1 U8711 ( .A(n12789), .ZN(n12952) );
  NAND2_X1 U8712 ( .A1(n8988), .A2(n8987), .ZN(n12964) );
  INV_X1 U8713 ( .A(n11807), .ZN(n12970) );
  NAND2_X1 U8714 ( .A1(n7516), .A2(n7521), .ZN(n12815) );
  NAND2_X1 U8715 ( .A1(n12836), .A2(n6543), .ZN(n7516) );
  NAND2_X1 U8716 ( .A1(n12834), .A2(n11805), .ZN(n12824) );
  NAND2_X1 U8717 ( .A1(n8924), .A2(n8923), .ZN(n12987) );
  NAND2_X1 U8718 ( .A1(n7142), .A2(n12056), .ZN(n12848) );
  NAND2_X1 U8719 ( .A1(n12859), .A2(n12860), .ZN(n7142) );
  NAND2_X1 U8720 ( .A1(n8872), .A2(n8871), .ZN(n12408) );
  NAND2_X1 U8721 ( .A1(n11362), .A2(n12042), .ZN(n11405) );
  NAND2_X1 U8722 ( .A1(n8854), .A2(n8853), .ZN(n11420) );
  NAND2_X1 U8723 ( .A1(n9724), .A2(n8695), .ZN(n6718) );
  INV_X1 U8724 ( .A(P3_IR_REG_29__SCAN_IN), .ZN(n8600) );
  INV_X1 U8725 ( .A(n8604), .ZN(n11466) );
  XNOR2_X1 U8726 ( .A(n8621), .B(n8620), .ZN(n11352) );
  OAI21_X1 U8727 ( .B1(n9100), .B2(P3_IR_REG_24__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8621) );
  XNOR2_X1 U8728 ( .A(n9047), .B(P2_DATAO_REG_24__SCAN_IN), .ZN(n11275) );
  XNOR2_X1 U8729 ( .A(n8619), .B(P3_IR_REG_24__SCAN_IN), .ZN(n8626) );
  NAND2_X1 U8730 ( .A1(n9100), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8619) );
  INV_X1 U8731 ( .A(n7356), .ZN(n9015) );
  NAND2_X1 U8732 ( .A1(n9087), .A2(n9098), .ZN(n11288) );
  INV_X1 U8733 ( .A(SI_20_), .ZN(n10609) );
  NAND2_X1 U8734 ( .A1(n7347), .A2(n7348), .ZN(n8970) );
  NAND2_X1 U8735 ( .A1(n7352), .A2(n7354), .ZN(n8955) );
  OR2_X1 U8736 ( .A1(n8936), .A2(n8935), .ZN(n7352) );
  INV_X1 U8737 ( .A(SI_15_), .ZN(n9705) );
  NAND2_X1 U8738 ( .A1(n7335), .A2(n8884), .ZN(n8896) );
  NAND2_X1 U8739 ( .A1(n8883), .A2(n8882), .ZN(n7335) );
  NAND2_X1 U8740 ( .A1(n7366), .A2(n8823), .ZN(n8841) );
  NAND2_X1 U8741 ( .A1(n7367), .A2(n6669), .ZN(n7366) );
  INV_X1 U8742 ( .A(SI_12_), .ZN(n15403) );
  INV_X1 U8743 ( .A(SI_10_), .ZN(n14369) );
  INV_X1 U8744 ( .A(n10648), .ZN(n11090) );
  NAND2_X1 U8745 ( .A1(n7342), .A2(n8647), .ZN(n8776) );
  NAND2_X1 U8746 ( .A1(n8767), .A2(n8766), .ZN(n7342) );
  NAND2_X1 U8747 ( .A1(n7327), .A2(n8643), .ZN(n8744) );
  NAND2_X1 U8748 ( .A1(n8677), .A2(n8676), .ZN(n7327) );
  NAND2_X1 U8749 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(P3_IR_REG_31__SCAN_IN), .ZN(
        n6826) );
  INV_X1 U8750 ( .A(n13038), .ZN(n6934) );
  NAND2_X1 U8751 ( .A1(n13469), .A2(n14479), .ZN(n13044) );
  NAND2_X1 U8752 ( .A1(n11112), .A2(n7394), .ZN(n14456) );
  AND2_X1 U8753 ( .A1(n9963), .A2(n9303), .ZN(n13131) );
  NAND2_X1 U8754 ( .A1(n9250), .A2(n10929), .ZN(n10935) );
  NAND2_X1 U8755 ( .A1(n6931), .A2(n10343), .ZN(n10353) );
  NAND2_X1 U8756 ( .A1(n6940), .A2(n6938), .ZN(n13088) );
  AOI21_X1 U8757 ( .B1(n6640), .B2(n6923), .A(n6561), .ZN(n6919) );
  NAND2_X1 U8758 ( .A1(n6920), .A2(n6922), .ZN(n13101) );
  NAND2_X1 U8759 ( .A1(n14473), .A2(n6924), .ZN(n6920) );
  NAND2_X1 U8760 ( .A1(n6926), .A2(n7373), .ZN(n13120) );
  NAND2_X1 U8761 ( .A1(n10353), .A2(n9218), .ZN(n10268) );
  INV_X1 U8762 ( .A(n8547), .ZN(n6975) );
  OR2_X1 U8763 ( .A1(n8162), .A2(n7760), .ZN(n7764) );
  OR2_X1 U8764 ( .A1(n8176), .A2(n7761), .ZN(n7763) );
  MUX2_X1 U8765 ( .A(n9545), .B(P2_REG1_REG_2__SCAN_IN), .S(n13162), .Z(n13166) );
  AOI21_X1 U8766 ( .B1(n13183), .B2(n9576), .A(n9575), .ZN(n9661) );
  NOR2_X1 U8767 ( .A1(n9876), .A2(n6671), .ZN(n14803) );
  INV_X1 U8768 ( .A(n6955), .ZN(n14801) );
  INV_X1 U8769 ( .A(n6953), .ZN(n14816) );
  NOR2_X1 U8770 ( .A1(n10170), .A2(n10169), .ZN(n11025) );
  AND2_X1 U8771 ( .A1(n11026), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n6963) );
  NOR2_X1 U8772 ( .A1(n6691), .A2(n6961), .ZN(n6960) );
  NOR2_X1 U8773 ( .A1(n14855), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n6961) );
  INV_X1 U8774 ( .A(n6959), .ZN(n11164) );
  AOI211_X1 U8775 ( .C1(n13438), .C2(n11031), .A(n11030), .B(n11032), .ZN(
        n11159) );
  XOR2_X1 U8776 ( .A(n11452), .B(n11443), .Z(n11445) );
  INV_X1 U8777 ( .A(n6957), .ZN(n11451) );
  OAI211_X1 U8778 ( .C1(n13202), .C2(n13200), .A(n13199), .B(n13198), .ZN(
        n13210) );
  AND2_X1 U8779 ( .A1(n11450), .A2(n11449), .ZN(n13202) );
  AND2_X1 U8780 ( .A1(n7204), .A2(n7207), .ZN(n13462) );
  NAND2_X1 U8781 ( .A1(n7446), .A2(n7445), .ZN(n13265) );
  NAND2_X1 U8782 ( .A1(n7446), .A2(n7442), .ZN(n13467) );
  NAND2_X1 U8783 ( .A1(n8129), .A2(n8128), .ZN(n13478) );
  NAND2_X1 U8784 ( .A1(n7453), .A2(n7451), .ZN(n13309) );
  NAND2_X1 U8785 ( .A1(n13340), .A2(n7454), .ZN(n7453) );
  NAND2_X1 U8786 ( .A1(n13340), .A2(n8094), .ZN(n13322) );
  NAND2_X1 U8787 ( .A1(n13353), .A2(n8263), .ZN(n13337) );
  NAND2_X1 U8788 ( .A1(n7460), .A2(n8072), .ZN(n13365) );
  NAND2_X1 U8789 ( .A1(n7461), .A2(n6573), .ZN(n7460) );
  NAND2_X1 U8790 ( .A1(n7214), .A2(n8259), .ZN(n13369) );
  NAND2_X1 U8791 ( .A1(n8258), .A2(n8257), .ZN(n13388) );
  NAND2_X1 U8792 ( .A1(n7464), .A2(n7463), .ZN(n13398) );
  NAND2_X1 U8793 ( .A1(n7200), .A2(n7201), .ZN(n13420) );
  OR2_X1 U8794 ( .A1(n13532), .A2(n7203), .ZN(n7200) );
  NAND2_X1 U8795 ( .A1(n7987), .A2(n7986), .ZN(n14489) );
  NAND2_X1 U8796 ( .A1(n7171), .A2(n6547), .ZN(n11227) );
  NAND2_X1 U8797 ( .A1(n10901), .A2(n8249), .ZN(n11076) );
  NAND2_X1 U8798 ( .A1(n8240), .A2(n8239), .ZN(n10202) );
  NAND2_X1 U8799 ( .A1(n10182), .A2(n10185), .ZN(n10181) );
  NAND2_X1 U8800 ( .A1(n10221), .A2(n7831), .ZN(n10182) );
  NAND2_X1 U8801 ( .A1(n7175), .A2(n8231), .ZN(n10255) );
  OR2_X1 U8802 ( .A1(n7178), .A2(n10232), .ZN(n7175) );
  INV_X1 U8803 ( .A(n13444), .ZN(n13432) );
  INV_X1 U8804 ( .A(n13414), .ZN(n13440) );
  INV_X1 U8805 ( .A(n13393), .ZN(n13442) );
  INV_X1 U8806 ( .A(n13232), .ZN(n13546) );
  OR2_X1 U8807 ( .A1(n13460), .A2(n13519), .ZN(n6725) );
  NAND2_X1 U8808 ( .A1(n7885), .A2(n7884), .ZN(n10750) );
  INV_X1 U8809 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n13576) );
  AND2_X1 U8810 ( .A1(n7467), .A2(n7738), .ZN(n7466) );
  OAI21_X1 U8811 ( .B1(n8204), .B2(P2_IR_REG_25__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8206) );
  INV_X1 U8812 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n11427) );
  XNOR2_X1 U8813 ( .A(n8198), .B(n8197), .ZN(n11426) );
  NAND2_X1 U8814 ( .A1(n8223), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8225) );
  OAI21_X1 U8815 ( .B1(n6535), .B2(n7728), .A(n6638), .ZN(n8223) );
  INV_X1 U8816 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n11045) );
  AND2_X1 U8817 ( .A1(n6984), .A2(n15356), .ZN(n6983) );
  INV_X1 U8818 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n9701) );
  INV_X1 U8819 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n9700) );
  AND2_X1 U8820 ( .A1(n7869), .A2(n7896), .ZN(n14819) );
  INV_X1 U8821 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n9496) );
  INV_X1 U8822 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n9494) );
  AND2_X1 U8823 ( .A1(n7794), .A2(n7802), .ZN(n13184) );
  INV_X1 U8824 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n9493) );
  INV_X1 U8825 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n9474) );
  NAND2_X1 U8826 ( .A1(n6950), .A2(n7757), .ZN(n14791) );
  AOI22_X1 U8827 ( .A1(n7728), .A2(n6951), .B1(P2_IR_REG_31__SCAN_IN), .B2(
        n6548), .ZN(n6950) );
  INV_X1 U8828 ( .A(n13981), .ZN(n14171) );
  NAND2_X1 U8829 ( .A1(n11262), .A2(n11261), .ZN(n11376) );
  NAND2_X1 U8830 ( .A1(n9986), .A2(n9417), .ZN(n9439) );
  NAND2_X1 U8831 ( .A1(n11537), .A2(n11536), .ZN(n14197) );
  NAND2_X1 U8832 ( .A1(n10974), .A2(n10973), .ZN(n10987) );
  AND2_X1 U8833 ( .A1(n9392), .A2(n9896), .ZN(n10014) );
  AND2_X1 U8834 ( .A1(n7221), .A2(n10632), .ZN(n10592) );
  NAND2_X1 U8835 ( .A1(n10633), .A2(n10634), .ZN(n7221) );
  NAND2_X1 U8836 ( .A1(n7241), .A2(n7242), .ZN(n13673) );
  NAND2_X1 U8837 ( .A1(n11376), .A2(n11375), .ZN(n11378) );
  NAND2_X1 U8838 ( .A1(n7245), .A2(n7240), .ZN(n7237) );
  INV_X1 U8839 ( .A(n10590), .ZN(n7222) );
  AND2_X1 U8840 ( .A1(n7224), .A2(n13731), .ZN(n7223) );
  NAND2_X1 U8841 ( .A1(n7227), .A2(n7229), .ZN(n7224) );
  OAI21_X1 U8842 ( .B1(n13686), .B2(n7229), .A(n7227), .ZN(n13730) );
  OAI21_X1 U8843 ( .B1(n12376), .B2(n12375), .A(n6627), .ZN(n7066) );
  NOR3_X1 U8844 ( .A1(n12379), .A2(n12378), .A3(n12377), .ZN(n12380) );
  OR2_X1 U8845 ( .A1(n11530), .A2(n11529), .ZN(n13763) );
  INV_X1 U8846 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n9984) );
  AND4_X1 U8847 ( .A1(n9752), .A2(n9751), .A3(n9750), .A4(n9749), .ZN(n13663)
         );
  INV_X1 U8848 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n9763) );
  AND4_X1 U8849 ( .A1(n9762), .A2(n9761), .A3(n9760), .A4(n9759), .ZN(n12186)
         );
  OR2_X1 U8850 ( .A1(n11600), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n9328) );
  AOI21_X1 U8851 ( .B1(P1_REG1_REG_3__SCAN_IN), .B2(n9630), .A(n9626), .ZN(
        n9915) );
  AOI21_X1 U8852 ( .B1(n10401), .B2(P1_REG1_REG_6__SCAN_IN), .A(n9706), .ZN(
        n9708) );
  AOI21_X1 U8853 ( .B1(n10999), .B2(P1_REG1_REG_10__SCAN_IN), .A(n10021), .ZN(
        n10023) );
  NAND2_X1 U8854 ( .A1(n10320), .A2(n10319), .ZN(n10791) );
  NAND2_X1 U8855 ( .A1(n13824), .A2(n13825), .ZN(n13846) );
  XNOR2_X1 U8856 ( .A(n13853), .B(n13852), .ZN(n13849) );
  NAND2_X1 U8857 ( .A1(n11597), .A2(n11596), .ZN(n13891) );
  AND2_X1 U8858 ( .A1(n7014), .A2(n6586), .ZN(n11607) );
  NAND2_X1 U8859 ( .A1(n7089), .A2(n7092), .ZN(n13931) );
  NAND2_X1 U8860 ( .A1(n6765), .A2(n7090), .ZN(n7089) );
  NAND2_X1 U8861 ( .A1(n6765), .A2(n11620), .ZN(n13953) );
  NAND2_X1 U8862 ( .A1(n7534), .A2(n7530), .ZN(n7527) );
  INV_X1 U8863 ( .A(n6788), .ZN(n13985) );
  INV_X1 U8864 ( .A(n6769), .ZN(n14009) );
  NAND2_X1 U8865 ( .A1(n7506), .A2(n12336), .ZN(n14054) );
  OR2_X1 U8866 ( .A1(n6750), .A2(n12335), .ZN(n7506) );
  NAND2_X1 U8867 ( .A1(n7081), .A2(n11197), .ZN(n11306) );
  NAND2_X1 U8868 ( .A1(n6763), .A2(n12350), .ZN(n7081) );
  NAND2_X1 U8869 ( .A1(n11200), .A2(n11199), .ZN(n13706) );
  NAND2_X1 U8870 ( .A1(n10997), .A2(n10996), .ZN(n11003) );
  NAND2_X1 U8871 ( .A1(n10681), .A2(n10680), .ZN(n14743) );
  INV_X1 U8872 ( .A(n14117), .ZN(n14669) );
  INV_X1 U8873 ( .A(n14673), .ZN(n14659) );
  INV_X1 U8874 ( .A(n14089), .ZN(n14662) );
  INV_X1 U8875 ( .A(n14095), .ZN(n14676) );
  INV_X1 U8876 ( .A(n14052), .ZN(n14675) );
  AND2_X1 U8877 ( .A1(n14220), .A2(n9448), .ZN(n14673) );
  AND2_X2 U8878 ( .A1(n14223), .A2(n14127), .ZN(n14788) );
  NAND2_X1 U8879 ( .A1(n14142), .A2(n6791), .ZN(n14227) );
  OR2_X1 U8880 ( .A1(n14194), .A2(n14193), .ZN(n14237) );
  OR2_X1 U8881 ( .A1(n9319), .A2(n9318), .ZN(n9321) );
  NAND2_X1 U8882 ( .A1(n8170), .A2(n8169), .ZN(n13584) );
  INV_X1 U8883 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n9338) );
  CLKBUF_X1 U8884 ( .A(n9599), .Z(n13875) );
  NAND2_X1 U8885 ( .A1(n9340), .A2(n9189), .ZN(n14249) );
  INV_X1 U8886 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n15197) );
  INV_X1 U8887 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n15212) );
  NAND2_X1 U8888 ( .A1(n9184), .A2(n9183), .ZN(n11348) );
  CLKBUF_X1 U8889 ( .A(n14251), .Z(n6796) );
  INV_X1 U8890 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n11487) );
  INV_X1 U8891 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n10672) );
  INV_X1 U8892 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n10502) );
  INV_X1 U8893 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n9848) );
  INV_X1 U8894 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n9623) );
  INV_X1 U8895 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n15379) );
  INV_X1 U8896 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n9509) );
  INV_X1 U8897 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n9505) );
  INV_X1 U8898 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n9165) );
  INV_X1 U8899 ( .A(n7303), .ZN(n7775) );
  MUX2_X1 U8900 ( .A(n9318), .B(n9404), .S(P1_IR_REG_2__SCAN_IN), .Z(n9405) );
  NAND2_X1 U8901 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n9363) );
  NAND2_X1 U8902 ( .A1(n6738), .A2(n14296), .ZN(n14350) );
  INV_X1 U8903 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n7039) );
  XNOR2_X1 U8904 ( .A(n14312), .B(n7037), .ZN(n15430) );
  XNOR2_X1 U8905 ( .A(n14322), .B(n7034), .ZN(n14386) );
  INV_X1 U8906 ( .A(n14323), .ZN(n7034) );
  OAI21_X1 U8907 ( .B1(n7029), .B2(n7028), .A(n14859), .ZN(n7027) );
  AND2_X1 U8908 ( .A1(n6767), .A2(n7025), .ZN(n14400) );
  NAND2_X1 U8909 ( .A1(n7024), .A2(n14598), .ZN(n6767) );
  NAND2_X1 U8910 ( .A1(n14596), .A2(n14597), .ZN(n7024) );
  NAND2_X1 U8911 ( .A1(n14400), .A2(n14401), .ZN(n14399) );
  OAI21_X1 U8912 ( .B1(P3_U3897), .B2(n7149), .A(n7148), .ZN(P3_U3491) );
  INV_X1 U8913 ( .A(P3_DATAO_REG_0__SCAN_IN), .ZN(n7149) );
  INV_X1 U8914 ( .A(n6822), .ZN(n12588) );
  AOI21_X1 U8915 ( .B1(n6829), .B2(n7279), .A(n6827), .ZN(n12687) );
  NAND2_X1 U8916 ( .A1(n12703), .A2(n12684), .ZN(n6829) );
  AOI21_X1 U8917 ( .B1(n7280), .B2(n7279), .A(n7276), .ZN(n12707) );
  AOI21_X1 U8918 ( .B1(n7549), .B2(n15043), .A(n6566), .ZN(n7547) );
  AOI21_X1 U8919 ( .B1(n12931), .B2(n15110), .A(n7167), .ZN(n12933) );
  NAND2_X1 U8920 ( .A1(n7169), .A2(n7168), .ZN(n7167) );
  NAND2_X1 U8921 ( .A1(n15109), .A2(P3_REG0_REG_28__SCAN_IN), .ZN(n7168) );
  INV_X1 U8922 ( .A(n7369), .ZN(n13025) );
  NAND2_X1 U8923 ( .A1(n7384), .A2(n14462), .ZN(n7382) );
  NAND2_X1 U8924 ( .A1(n7372), .A2(n7378), .ZN(n11441) );
  NOR2_X1 U8925 ( .A1(n6945), .A2(n13224), .ZN(n13223) );
  AOI21_X1 U8926 ( .B1(n6944), .B2(n14491), .A(n6943), .ZN(n6942) );
  INV_X1 U8927 ( .A(n13226), .ZN(n13228) );
  INV_X1 U8928 ( .A(n8296), .ZN(n8297) );
  OAI21_X1 U8929 ( .B1(n13459), .B2(n13419), .A(n8295), .ZN(n8296) );
  OAI21_X1 U8930 ( .B1(n13541), .B2(n14930), .A(n7398), .ZN(P2_U3530) );
  AOI21_X1 U8931 ( .B1(n13235), .B2(n13465), .A(n7399), .ZN(n7398) );
  NOR2_X1 U8932 ( .A1(n14929), .A2(n13451), .ZN(n7399) );
  NAND2_X1 U8933 ( .A1(n7471), .A2(n7469), .ZN(P2_U3527) );
  AOI21_X1 U8934 ( .B1(n13464), .B2(n13465), .A(n7470), .ZN(n7469) );
  NAND2_X1 U8935 ( .A1(n13548), .A2(n14929), .ZN(n7471) );
  NOR2_X1 U8936 ( .A1(n14929), .A2(n15378), .ZN(n7470) );
  OAI21_X1 U8937 ( .B1(n13541), .B2(n14924), .A(n6907), .ZN(P2_U3498) );
  AOI21_X1 U8938 ( .B1(n13235), .B2(n6909), .A(n6908), .ZN(n6907) );
  NOR2_X1 U8939 ( .A1(n14925), .A2(n13542), .ZN(n6908) );
  OAI21_X1 U8940 ( .B1(n13548), .B2(n14924), .A(n6753), .ZN(n13549) );
  NAND2_X1 U8941 ( .A1(n14924), .A2(n15135), .ZN(n6753) );
  NAND2_X1 U8942 ( .A1(n11662), .A2(n11661), .ZN(n14532) );
  NAND2_X1 U8943 ( .A1(n6795), .A2(n6794), .ZN(n6793) );
  INV_X1 U8944 ( .A(n13659), .ZN(n6794) );
  NAND2_X1 U8945 ( .A1(n6711), .A2(n6708), .ZN(P1_U3262) );
  OR2_X1 U8946 ( .A1(n13870), .A2(n13868), .ZN(n6711) );
  AOI21_X1 U8947 ( .B1(n6710), .B2(n13868), .A(n6709), .ZN(n6708) );
  NAND2_X1 U8948 ( .A1(n14772), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n6774) );
  INV_X1 U8949 ( .A(n7029), .ZN(n14581) );
  INV_X1 U8950 ( .A(n7026), .ZN(n14579) );
  INV_X1 U8951 ( .A(n7025), .ZN(n14595) );
  NOR2_X1 U8952 ( .A1(n14407), .A2(n14406), .ZN(n14417) );
  NOR2_X1 U8953 ( .A1(n11806), .A2(n7522), .ZN(n6543) );
  AND2_X1 U8954 ( .A1(n14250), .A2(n11572), .ZN(n12276) );
  AND2_X1 U8955 ( .A1(n6639), .A2(n6888), .ZN(n6544) );
  OR2_X1 U8956 ( .A1(n14013), .A2(n13760), .ZN(n6545) );
  NAND2_X4 U8957 ( .A1(n7433), .A2(n6562), .ZN(n8709) );
  OAI21_X1 U8958 ( .B1(n15008), .B2(n11102), .A(n11131), .ZN(n11119) );
  INV_X1 U8959 ( .A(n12247), .ZN(n6699) );
  AND3_X1 U8960 ( .A1(n6894), .A2(n11948), .A3(n12479), .ZN(n6546) );
  AND2_X1 U8961 ( .A1(n7174), .A2(n8250), .ZN(n6547) );
  AND2_X1 U8962 ( .A1(n15330), .A2(P2_IR_REG_1__SCAN_IN), .ZN(n6548) );
  AND2_X1 U8963 ( .A1(n11668), .A2(n11667), .ZN(n6549) );
  AND2_X1 U8964 ( .A1(n7315), .A2(n7010), .ZN(n6550) );
  NAND2_X1 U8965 ( .A1(n15004), .A2(n7124), .ZN(n6551) );
  NAND2_X1 U8966 ( .A1(n12560), .A2(n12582), .ZN(n12587) );
  XNOR2_X1 U8967 ( .A(n12118), .B(n12750), .ZN(n12732) );
  INV_X1 U8968 ( .A(n12732), .ZN(n7490) );
  AND2_X1 U8969 ( .A1(n8424), .A2(n8423), .ZN(n6552) );
  AND2_X1 U8970 ( .A1(n12532), .A2(n6615), .ZN(n6553) );
  OR2_X1 U8971 ( .A1(n14153), .A2(n11621), .ZN(n6554) );
  AND2_X1 U8972 ( .A1(n13469), .A2(n13141), .ZN(n6555) );
  NAND2_X1 U8973 ( .A1(n11489), .A2(n11488), .ZN(n14013) );
  XOR2_X1 U8974 ( .A(n13238), .B(n13235), .Z(n6556) );
  AND2_X1 U8975 ( .A1(n13486), .A2(n13295), .ZN(n6557) );
  OR2_X1 U8976 ( .A1(n8430), .A2(n6989), .ZN(n6558) );
  NOR2_X1 U8977 ( .A1(n12979), .A2(n12838), .ZN(n6559) );
  AND2_X1 U8978 ( .A1(n7296), .A2(n12305), .ZN(n6560) );
  INV_X1 U8979 ( .A(n13235), .ZN(n13543) );
  AND2_X1 U8980 ( .A1(n13098), .A2(n9282), .ZN(n6561) );
  AND3_X1 U8981 ( .A1(n6876), .A2(n8627), .A3(n6875), .ZN(n6562) );
  AND2_X1 U8982 ( .A1(n14153), .A2(n11621), .ZN(n6563) );
  AND2_X1 U8983 ( .A1(n7299), .A2(SI_14_), .ZN(n6564) );
  XNOR2_X1 U8984 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .ZN(n8743) );
  INV_X1 U8985 ( .A(n8743), .ZN(n7326) );
  INV_X1 U8986 ( .A(n8996), .ZN(n6887) );
  AND2_X1 U8987 ( .A1(n7122), .A2(P3_REG2_REG_11__SCAN_IN), .ZN(n6565) );
  XNOR2_X1 U8988 ( .A(n12214), .B(n10995), .ZN(n12348) );
  INV_X1 U8989 ( .A(n12348), .ZN(n7101) );
  AND2_X1 U8990 ( .A1(n15109), .A2(n12925), .ZN(n6566) );
  INV_X1 U8991 ( .A(n14431), .ZN(n7165) );
  AND2_X1 U8992 ( .A1(n12383), .A2(n12384), .ZN(n6567) );
  NAND4_X1 U8993 ( .A1(n8598), .A2(n8599), .A3(n8630), .A4(n8597), .ZN(n6568)
         );
  AND2_X1 U8994 ( .A1(n11415), .A2(n12552), .ZN(n6569) );
  OR2_X1 U8995 ( .A1(n13222), .A2(n13221), .ZN(n6570) );
  INV_X1 U8996 ( .A(n7881), .ZN(n7645) );
  XNOR2_X1 U8997 ( .A(n7646), .B(SI_9_), .ZN(n7881) );
  INV_X1 U8998 ( .A(n8567), .ZN(n11075) );
  NAND2_X1 U8999 ( .A1(n9364), .A2(n9164), .ZN(n9343) );
  OR2_X1 U9000 ( .A1(n13981), .A2(n13758), .ZN(n6571) );
  INV_X1 U9001 ( .A(n8578), .ZN(n8275) );
  OR2_X1 U9002 ( .A1(n11630), .A2(n13891), .ZN(n6572) );
  OR2_X1 U9003 ( .A1(n13511), .A2(n13355), .ZN(n6573) );
  INV_X1 U9004 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n8043) );
  AND2_X1 U9005 ( .A1(n9437), .A2(n9417), .ZN(n6574) );
  INV_X1 U9006 ( .A(n8576), .ZN(n13246) );
  OR2_X1 U9007 ( .A1(n7621), .A2(n9466), .ZN(n6575) );
  NAND2_X1 U9008 ( .A1(n11196), .A2(n11195), .ZN(n12235) );
  XOR2_X1 U9009 ( .A(n13326), .B(n13024), .Z(n6576) );
  AND2_X1 U9010 ( .A1(n8414), .A2(n8413), .ZN(n6577) );
  NAND2_X1 U9011 ( .A1(n8426), .A2(n8425), .ZN(n6578) );
  AND2_X1 U9012 ( .A1(n8468), .A2(n8467), .ZN(n6579) );
  XOR2_X1 U9013 ( .A(n11671), .B(n11775), .Z(n6580) );
  AND2_X1 U9014 ( .A1(n7157), .A2(n12085), .ZN(n6581) );
  NOR2_X1 U9015 ( .A1(n9497), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n9479) );
  NAND2_X1 U9016 ( .A1(n14883), .A2(n11796), .ZN(n8393) );
  NOR2_X1 U9017 ( .A1(n11610), .A2(n14082), .ZN(n6582) );
  NOR2_X1 U9018 ( .A1(n14204), .A2(n13763), .ZN(n6583) );
  OR2_X1 U9019 ( .A1(n8351), .A2(n8350), .ZN(n6584) );
  NAND3_X1 U9020 ( .A1(n7542), .A2(n8596), .A3(n7166), .ZN(n6585) );
  INV_X1 U9021 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n15262) );
  INV_X1 U9022 ( .A(n10149), .ZN(n7481) );
  NAND2_X1 U9023 ( .A1(n14153), .A2(n13755), .ZN(n6586) );
  INV_X1 U9024 ( .A(n12332), .ZN(n6838) );
  AOI21_X1 U9025 ( .B1(n7998), .B2(n7008), .A(n7007), .ZN(n7006) );
  INV_X1 U9026 ( .A(n7006), .ZN(n6833) );
  OR3_X1 U9027 ( .A1(n12772), .A2(n12079), .A3(n12078), .ZN(n6587) );
  AND3_X1 U9028 ( .A1(n14056), .A2(n12261), .A3(n12260), .ZN(n6588) );
  BUF_X2 U9029 ( .A(n12173), .Z(n12328) );
  MUX2_X2 U9030 ( .A(n6773), .B(n12142), .S(n12326), .Z(n12179) );
  OR2_X1 U9031 ( .A1(n13364), .A2(n7459), .ZN(n6589) );
  AND2_X1 U9032 ( .A1(n14358), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n6590) );
  OR2_X1 U9033 ( .A1(n12680), .A2(n12679), .ZN(n6591) );
  NAND2_X1 U9034 ( .A1(n9019), .A2(n9018), .ZN(n12479) );
  OR3_X1 U9035 ( .A1(P3_IR_REG_2__SCAN_IN), .A2(P3_IR_REG_1__SCAN_IN), .A3(
        P3_IR_REG_0__SCAN_IN), .ZN(n6592) );
  OR2_X1 U9036 ( .A1(n13992), .A2(n13981), .ZN(n6593) );
  OR2_X1 U9037 ( .A1(n11572), .A2(n9652), .ZN(n6594) );
  AND2_X1 U9038 ( .A1(n14362), .A2(n15113), .ZN(n6595) );
  OR2_X1 U9039 ( .A1(n14306), .A2(n14305), .ZN(n6596) );
  INV_X1 U9040 ( .A(n13721), .ZN(n7245) );
  AND2_X1 U9041 ( .A1(n12374), .A2(n12383), .ZN(n6597) );
  AND2_X1 U9042 ( .A1(n10750), .A2(n13153), .ZN(n6598) );
  INV_X1 U9043 ( .A(n10860), .ZN(n7402) );
  INV_X1 U9044 ( .A(n7233), .ZN(n7232) );
  OAI21_X1 U9045 ( .B1(n13684), .B2(n13685), .A(n11742), .ZN(n7233) );
  NAND2_X1 U9046 ( .A1(n7955), .A2(n7954), .ZN(n13441) );
  AND2_X1 U9047 ( .A1(n8362), .A2(n8361), .ZN(n6599) );
  NOR2_X1 U9048 ( .A1(n8842), .A2(n7365), .ZN(n7364) );
  AND2_X1 U9049 ( .A1(n11816), .A2(n11815), .ZN(n6600) );
  AND2_X1 U9050 ( .A1(n13346), .A2(n9304), .ZN(n6601) );
  NAND2_X1 U9051 ( .A1(n6578), .A2(n6552), .ZN(n6994) );
  INV_X1 U9052 ( .A(n6994), .ZN(n6989) );
  OAI211_X1 U9053 ( .C1(n12562), .C2(n6819), .A(n6817), .B(n6815), .ZN(n12629)
         );
  INV_X1 U9054 ( .A(n7964), .ZN(n7664) );
  INV_X1 U9055 ( .A(n15004), .ZN(n10081) );
  OR2_X1 U9056 ( .A1(n13950), .A2(n11583), .ZN(n6602) );
  AND2_X1 U9057 ( .A1(n7453), .A2(n8558), .ZN(n6603) );
  OR2_X1 U9058 ( .A1(n11807), .A2(n12453), .ZN(n6604) );
  NAND2_X1 U9059 ( .A1(n13441), .A2(n13149), .ZN(n6605) );
  AND2_X1 U9060 ( .A1(n6946), .A2(n6947), .ZN(n6606) );
  AND2_X1 U9061 ( .A1(n7101), .A2(n10875), .ZN(n6607) );
  INV_X1 U9062 ( .A(n8151), .ZN(n7447) );
  INV_X1 U9063 ( .A(n12275), .ZN(n7072) );
  AND2_X1 U9064 ( .A1(n7214), .A2(n7212), .ZN(n6608) );
  AND2_X1 U9065 ( .A1(n10624), .A2(n8771), .ZN(n12003) );
  INV_X1 U9066 ( .A(n7531), .ZN(n7530) );
  NAND2_X1 U9067 ( .A1(n7535), .A2(n6571), .ZN(n7531) );
  INV_X1 U9068 ( .A(n7265), .ZN(n13944) );
  NOR2_X1 U9069 ( .A1(n13992), .A2(n7267), .ZN(n7265) );
  AND2_X1 U9070 ( .A1(n9293), .A2(n9287), .ZN(n6609) );
  AND2_X1 U9071 ( .A1(n7490), .A2(n11815), .ZN(n6610) );
  AND2_X1 U9072 ( .A1(n8232), .A2(n13050), .ZN(n6611) );
  AND2_X1 U9073 ( .A1(n7056), .A2(n7055), .ZN(n6612) );
  AND2_X1 U9074 ( .A1(n11279), .A2(n14428), .ZN(n6613) );
  INV_X1 U9075 ( .A(n7093), .ZN(n7092) );
  INV_X1 U9076 ( .A(n7455), .ZN(n7454) );
  OR2_X1 U9077 ( .A1(n8110), .A2(n7456), .ZN(n7455) );
  AND2_X1 U9078 ( .A1(n14480), .A2(n13537), .ZN(n6614) );
  OR2_X1 U9079 ( .A1(n8880), .A2(n7410), .ZN(n6615) );
  AND2_X1 U9080 ( .A1(n11606), .A2(n6586), .ZN(n6616) );
  OR2_X1 U9081 ( .A1(n8327), .A2(n8328), .ZN(n6617) );
  INV_X1 U9082 ( .A(n7537), .ZN(n7536) );
  NOR2_X1 U9083 ( .A1(n14171), .A2(n11618), .ZN(n7537) );
  AND2_X1 U9084 ( .A1(n12036), .A2(n12037), .ZN(n11933) );
  OR2_X1 U9085 ( .A1(n11869), .A2(n11868), .ZN(n6618) );
  AND2_X1 U9086 ( .A1(n8418), .A2(n8417), .ZN(n6619) );
  AND2_X1 U9087 ( .A1(n7533), .A2(n7532), .ZN(n6620) );
  NOR2_X1 U9088 ( .A1(n10487), .A2(n13156), .ZN(n6621) );
  NOR2_X1 U9089 ( .A1(n14204), .A2(n13626), .ZN(n6622) );
  NOR2_X1 U9090 ( .A1(n13706), .A2(n11307), .ZN(n6623) );
  INV_X1 U9091 ( .A(n7240), .ZN(n7239) );
  NAND2_X1 U9092 ( .A1(n7242), .A2(n11688), .ZN(n7240) );
  AND2_X1 U9093 ( .A1(n8391), .A2(n8390), .ZN(n6624) );
  OR2_X1 U9094 ( .A1(n6563), .A2(n7093), .ZN(n6625) );
  AND2_X1 U9095 ( .A1(n8464), .A2(n8463), .ZN(n6626) );
  AND2_X1 U9096 ( .A1(n12373), .A2(n6597), .ZN(n6627) );
  AND2_X1 U9097 ( .A1(n13894), .A2(n13895), .ZN(n14135) );
  AND2_X1 U9098 ( .A1(n7161), .A2(n12037), .ZN(n6628) );
  AND2_X1 U9099 ( .A1(n7646), .A2(SI_9_), .ZN(n6629) );
  OR2_X1 U9100 ( .A1(n14256), .A2(n14956), .ZN(n6630) );
  AND2_X1 U9101 ( .A1(n7590), .A2(n6619), .ZN(n6631) );
  NOR2_X1 U9102 ( .A1(n12124), .A2(n12388), .ZN(n6632) );
  AND2_X1 U9103 ( .A1(n9274), .A2(n9273), .ZN(n6633) );
  AND2_X1 U9104 ( .A1(n7640), .A2(SI_7_), .ZN(n6634) );
  NOR2_X1 U9105 ( .A1(n14498), .A2(n14468), .ZN(n6635) );
  NOR2_X1 U9106 ( .A1(n13326), .A2(n13086), .ZN(n6636) );
  AND2_X1 U9107 ( .A1(n9263), .A2(n9262), .ZN(n6637) );
  AND2_X1 U9108 ( .A1(n7395), .A2(n8222), .ZN(n6638) );
  INV_X1 U9109 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n9492) );
  INV_X1 U9110 ( .A(n12839), .ZN(n6716) );
  NOR2_X1 U9111 ( .A1(n12450), .A2(n7427), .ZN(n6639) );
  AND2_X1 U9112 ( .A1(n6921), .A2(n9280), .ZN(n6640) );
  AND2_X1 U9113 ( .A1(n9509), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n6641) );
  AND2_X1 U9114 ( .A1(n9763), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n6642) );
  NAND2_X1 U9115 ( .A1(n8431), .A2(n6993), .ZN(n6643) );
  INV_X1 U9116 ( .A(n12276), .ZN(n13997) );
  OR2_X1 U9117 ( .A1(n8431), .A2(n6989), .ZN(n6644) );
  AND2_X1 U9118 ( .A1(n13528), .A2(n7979), .ZN(n8566) );
  OR2_X1 U9119 ( .A1(n13911), .A2(n13913), .ZN(n6645) );
  AND2_X1 U9120 ( .A1(n15356), .A2(n8221), .ZN(n6646) );
  INV_X1 U9121 ( .A(n9357), .ZN(n6773) );
  AND2_X1 U9122 ( .A1(n8618), .A2(n7435), .ZN(n6647) );
  INV_X1 U9123 ( .A(n12235), .ZN(n14393) );
  INV_X1 U9124 ( .A(n7249), .ZN(n7248) );
  NAND2_X1 U9125 ( .A1(n7250), .A2(n11375), .ZN(n7249) );
  NAND2_X1 U9126 ( .A1(n8434), .A2(n8435), .ZN(n6648) );
  OR2_X1 U9127 ( .A1(n14135), .A2(n14134), .ZN(n6649) );
  OR2_X1 U9128 ( .A1(n12680), .A2(n12665), .ZN(n6650) );
  AND3_X1 U9129 ( .A1(n7725), .A2(n8192), .A3(n8197), .ZN(n6651) );
  AND2_X1 U9130 ( .A1(n11690), .A2(n11691), .ZN(n6652) );
  INV_X1 U9131 ( .A(n8460), .ZN(n7574) );
  INV_X1 U9132 ( .A(n8387), .ZN(n7580) );
  AND2_X1 U9133 ( .A1(n7253), .A2(n6580), .ZN(n6653) );
  AND2_X1 U9134 ( .A1(n7337), .A2(n12757), .ZN(n6654) );
  AND2_X1 U9135 ( .A1(n13461), .A2(n7207), .ZN(n6655) );
  INV_X1 U9136 ( .A(n10070), .ZN(n7124) );
  AND2_X1 U9137 ( .A1(n7545), .A2(n7544), .ZN(n6656) );
  AND2_X1 U9138 ( .A1(n6648), .A2(n6990), .ZN(n6657) );
  AND2_X1 U9139 ( .A1(n12783), .A2(n11810), .ZN(n6658) );
  AND2_X1 U9140 ( .A1(n6822), .A2(n12587), .ZN(n6659) );
  OR2_X1 U9141 ( .A1(n7072), .A2(n12274), .ZN(n6660) );
  AND2_X1 U9142 ( .A1(n14147), .A2(n6776), .ZN(n6661) );
  AND2_X1 U9143 ( .A1(n7369), .A2(n7368), .ZN(n6662) );
  AND2_X1 U9144 ( .A1(n7288), .A2(n12611), .ZN(n6663) );
  AND2_X1 U9145 ( .A1(n6647), .A2(n6896), .ZN(n6664) );
  NAND2_X1 U9146 ( .A1(n7068), .A2(n12216), .ZN(n6665) );
  INV_X1 U9147 ( .A(n7388), .ZN(n7387) );
  OR2_X1 U9148 ( .A1(n13068), .A2(n13064), .ZN(n7388) );
  INV_X1 U9149 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n8651) );
  INV_X1 U9150 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n7738) );
  NAND2_X1 U9151 ( .A1(n8401), .A2(n8400), .ZN(n6666) );
  INV_X1 U9152 ( .A(n6918), .ZN(n6922) );
  NAND2_X1 U9153 ( .A1(n6923), .A2(n9280), .ZN(n6918) );
  NAND2_X1 U9154 ( .A1(n7561), .A2(n8448), .ZN(n6667) );
  AND2_X2 U9155 ( .A1(n13901), .A2(n14659), .ZN(n14674) );
  INV_X1 U9156 ( .A(n8162), .ZN(n7808) );
  INV_X1 U9157 ( .A(n12860), .ZN(n7138) );
  INV_X1 U9158 ( .A(n13346), .ZN(n6905) );
  AND2_X1 U9159 ( .A1(n7433), .A2(n8627), .ZN(n9069) );
  INV_X1 U9160 ( .A(P3_IR_REG_21__SCAN_IN), .ZN(n6896) );
  NAND2_X1 U9161 ( .A1(n6879), .A2(n9096), .ZN(n9070) );
  INV_X1 U9162 ( .A(n13759), .ZN(n7076) );
  NAND2_X1 U9163 ( .A1(n7409), .A2(n6553), .ZN(n12458) );
  AND2_X1 U9164 ( .A1(n6926), .A2(n6924), .ZN(n6668) );
  OR2_X1 U9165 ( .A1(P2_DATAO_REG_11__SCAN_IN), .A2(n9700), .ZN(n6669) );
  INV_X1 U9166 ( .A(SI_14_), .ZN(n8869) );
  NAND2_X1 U9167 ( .A1(n11376), .A2(n7248), .ZN(n11649) );
  INV_X1 U9168 ( .A(n13760), .ZN(n7078) );
  NAND2_X1 U9169 ( .A1(n7259), .A2(n9479), .ZN(n9952) );
  INV_X1 U9170 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n10178) );
  OR2_X1 U9171 ( .A1(n10651), .A2(n10073), .ZN(n6670) );
  NAND2_X1 U9172 ( .A1(n8144), .A2(n8143), .ZN(n13474) );
  INV_X1 U9173 ( .A(n13474), .ZN(n7401) );
  AND2_X1 U9174 ( .A1(n9884), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6671) );
  OR2_X1 U9175 ( .A1(n13086), .A2(n13316), .ZN(n6672) );
  XNOR2_X1 U9176 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .ZN(n8676) );
  INV_X1 U9177 ( .A(n8676), .ZN(n7323) );
  OR2_X1 U9178 ( .A1(n10651), .A2(n15125), .ZN(n6673) );
  AOI21_X1 U9179 ( .B1(n7504), .B2(n12335), .A(n6583), .ZN(n7503) );
  OR2_X1 U9180 ( .A1(n14986), .A2(n15121), .ZN(n6674) );
  AND2_X1 U9181 ( .A1(n9018), .A2(n11948), .ZN(n6675) );
  AND2_X1 U9182 ( .A1(n11096), .A2(n7273), .ZN(n6676) );
  INV_X1 U9183 ( .A(n8596), .ZN(n8938) );
  AND2_X1 U9184 ( .A1(n7241), .A2(n7239), .ZN(n6677) );
  INV_X1 U9185 ( .A(n7404), .ZN(n13382) );
  NOR2_X1 U9186 ( .A1(n13409), .A2(n13516), .ZN(n7404) );
  INV_X1 U9187 ( .A(n6906), .ZN(n13358) );
  NOR2_X1 U9188 ( .A1(n13374), .A2(n13359), .ZN(n6906) );
  AND2_X1 U9189 ( .A1(n7348), .A2(n7346), .ZN(n6678) );
  INV_X1 U9190 ( .A(n11096), .ZN(n11131) );
  AND2_X1 U9191 ( .A1(n7119), .A2(n7118), .ZN(n6679) );
  INV_X1 U9192 ( .A(n7270), .ZN(n14070) );
  NAND2_X1 U9193 ( .A1(n14083), .A2(n14082), .ZN(n6680) );
  AND2_X1 U9194 ( .A1(n7686), .A2(SI_20_), .ZN(n6681) );
  NAND2_X1 U9195 ( .A1(n14374), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n6682) );
  NOR2_X1 U9196 ( .A1(n7173), .A2(n7172), .ZN(n8251) );
  INV_X1 U9197 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n10179) );
  OR2_X1 U9198 ( .A1(n8954), .A2(n7351), .ZN(n6683) );
  AND2_X1 U9199 ( .A1(n7098), .A2(n11615), .ZN(n6684) );
  AND2_X1 U9200 ( .A1(n9589), .A2(P1_DATAO_REG_12__SCAN_IN), .ZN(n6685) );
  AND2_X1 U9201 ( .A1(n8897), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n6686) );
  INV_X1 U9202 ( .A(n11102), .ZN(n7273) );
  NAND2_X1 U9203 ( .A1(n12458), .A2(n8910), .ZN(n12457) );
  NOR2_X1 U9204 ( .A1(n8023), .A2(P2_IR_REG_18__SCAN_IN), .ZN(n6986) );
  INV_X1 U9205 ( .A(n6986), .ZN(n6985) );
  AND4_X1 U9206 ( .A1(n7715), .A2(n7714), .A3(n7713), .A4(n7712), .ZN(n7935)
         );
  INV_X1 U9207 ( .A(n8881), .ZN(n7410) );
  AND2_X1 U9208 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n6687) );
  AND2_X1 U9209 ( .A1(n11112), .A2(n9260), .ZN(n6688) );
  AND2_X1 U9210 ( .A1(n8965), .A2(n8953), .ZN(n6689) );
  AND2_X1 U9211 ( .A1(n13044), .A2(n13043), .ZN(n6690) );
  INV_X1 U9212 ( .A(n15018), .ZN(n7279) );
  INV_X1 U9213 ( .A(n13573), .ZN(n6909) );
  INV_X1 U9214 ( .A(n8895), .ZN(n7334) );
  INV_X1 U9215 ( .A(n6527), .ZN(n11044) );
  INV_X1 U9216 ( .A(n12636), .ZN(n14384) );
  INV_X2 U9217 ( .A(n14924), .ZN(n14925) );
  AND2_X1 U9218 ( .A1(n14855), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n6691) );
  INV_X1 U9219 ( .A(n15110), .ZN(n15109) );
  AND2_X1 U9220 ( .A1(n12618), .A2(n12626), .ZN(n6692) );
  INV_X1 U9221 ( .A(n13521), .ZN(n7405) );
  INV_X1 U9222 ( .A(n14204), .ZN(n7269) );
  AND2_X1 U9223 ( .A1(n14929), .A2(n14899), .ZN(n13465) );
  INV_X1 U9224 ( .A(n13511), .ZN(n7407) );
  OR2_X1 U9225 ( .A1(n11062), .A2(n7262), .ZN(n6693) );
  NAND2_X1 U9226 ( .A1(n9025), .A2(n9024), .ZN(n12797) );
  AND2_X1 U9227 ( .A1(n10876), .A2(n10875), .ZN(n6694) );
  INV_X1 U9228 ( .A(n6902), .ZN(n10560) );
  INV_X1 U9229 ( .A(n12590), .ZN(n7272) );
  INV_X1 U9230 ( .A(n7403), .ZN(n10857) );
  AND2_X1 U9231 ( .A1(n10814), .A2(n10813), .ZN(n6695) );
  AND2_X1 U9232 ( .A1(n6913), .A2(n7403), .ZN(n6696) );
  NOR2_X1 U9233 ( .A1(n9855), .A2(n7152), .ZN(n6697) );
  INV_X1 U9234 ( .A(n10479), .ZN(n6904) );
  INV_X1 U9235 ( .A(n12194), .ZN(n7261) );
  CLKBUF_X2 U9236 ( .A(n13779), .Z(n6770) );
  AND2_X1 U9237 ( .A1(n11968), .A2(n9937), .ZN(n12110) );
  INV_X1 U9238 ( .A(n12110), .ZN(n6876) );
  INV_X1 U9239 ( .A(n12557), .ZN(n7418) );
  INV_X1 U9240 ( .A(n14432), .ZN(n7164) );
  INV_X1 U9241 ( .A(n13877), .ZN(n12371) );
  NAND2_X1 U9242 ( .A1(n6901), .A2(n6902), .ZN(n6903) );
  XNOR2_X1 U9243 ( .A(n7074), .B(n7073), .ZN(n12144) );
  INV_X1 U9244 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n6951) );
  INV_X1 U9245 ( .A(n14952), .ZN(n7282) );
  INV_X1 U9246 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n7037) );
  NAND2_X1 U9247 ( .A1(n11165), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n6958) );
  AOI21_X1 U9248 ( .B1(P2_REG2_REG_13__SCAN_IN), .B2(n11165), .A(n11159), .ZN(
        n11443) );
  OR2_X1 U9249 ( .A1(n14498), .A2(n13400), .ZN(n7465) );
  NAND2_X1 U9250 ( .A1(n14498), .A2(n13400), .ZN(n7463) );
  NAND2_X2 U9251 ( .A1(n6533), .A2(P3_U3151), .ZN(n14368) );
  AOI21_X1 U9252 ( .B1(n12619), .B2(n12604), .A(n12626), .ZN(n12638) );
  NOR2_X1 U9253 ( .A1(n12590), .A2(n12626), .ZN(n6818) );
  OR3_X1 U9254 ( .A1(n12590), .A2(n12561), .A3(n12626), .ZN(n6819) );
  INV_X1 U9255 ( .A(n12626), .ZN(n6749) );
  NAND2_X2 U9256 ( .A1(n9599), .A2(n9450), .ZN(n11572) );
  OR2_X2 U9257 ( .A1(n14031), .A2(n14030), .ZN(n14189) );
  NAND2_X1 U9258 ( .A1(n7044), .A2(n7047), .ZN(n7042) );
  NAND2_X1 U9259 ( .A1(n7050), .A2(n7053), .ZN(n7049) );
  OAI21_X1 U9260 ( .B1(n12333), .B2(n6838), .A(n12334), .ZN(n6837) );
  NOR2_X1 U9261 ( .A1(n14940), .A2(n15115), .ZN(n14939) );
  NAND2_X1 U9262 ( .A1(n10653), .A2(n11090), .ZN(n11099) );
  NOR2_X1 U9263 ( .A1(n11123), .A2(n11122), .ZN(n12559) );
  AOI21_X1 U9264 ( .B1(n9814), .B2(P3_REG1_REG_2__SCAN_IN), .A(n6595), .ZN(
        n9808) );
  NOR2_X1 U9265 ( .A1(n15010), .A2(n15009), .ZN(n15008) );
  INV_X1 U9266 ( .A(n9794), .ZN(n6701) );
  NOR2_X1 U9267 ( .A1(n14995), .A2(n10083), .ZN(n10085) );
  NAND2_X1 U9268 ( .A1(n10974), .A2(n7255), .ZN(n11146) );
  NAND2_X1 U9269 ( .A1(n13642), .A2(n11653), .ZN(n13700) );
  NAND2_X1 U9270 ( .A1(n13603), .A2(n13604), .ZN(n13602) );
  NAND2_X2 U9271 ( .A1(n6799), .A2(n6798), .ZN(n13740) );
  NAND2_X1 U9272 ( .A1(n7225), .A2(n7223), .ZN(n13729) );
  NAND2_X1 U9273 ( .A1(n9394), .A2(n9393), .ZN(n10011) );
  XNOR2_X2 U9274 ( .A(n9334), .B(P1_IR_REG_21__SCAN_IN), .ZN(n9357) );
  NAND2_X1 U9275 ( .A1(n10970), .A2(n10969), .ZN(n10974) );
  NOR2_X1 U9276 ( .A1(n11101), .A2(n11100), .ZN(n15010) );
  NOR2_X1 U9277 ( .A1(n14996), .A2(n15123), .ZN(n14995) );
  NAND2_X1 U9278 ( .A1(n7217), .A2(n6797), .ZN(n10957) );
  NAND2_X1 U9279 ( .A1(n7238), .A2(n7237), .ZN(n13720) );
  OAI22_X1 U9280 ( .A1(n12612), .A2(n7286), .B1(n12611), .B2(n12630), .ZN(
        n12651) );
  NAND2_X1 U9281 ( .A1(n6949), .A2(n6948), .ZN(n6947) );
  NAND2_X1 U9282 ( .A1(n14852), .A2(n6960), .ZN(n14850) );
  NOR2_X1 U9283 ( .A1(n14829), .A2(n14828), .ZN(n14827) );
  NAND2_X1 U9284 ( .A1(n9881), .A2(n9880), .ZN(n10164) );
  NOR2_X1 U9285 ( .A1(n9657), .A2(n9656), .ZN(n9655) );
  OAI21_X1 U9286 ( .B1(n13190), .B2(n14509), .A(n13189), .ZN(n13192) );
  INV_X1 U9287 ( .A(n13224), .ZN(n6946) );
  NAND2_X1 U9288 ( .A1(n6759), .A2(n6757), .ZN(n6944) );
  NOR2_X1 U9289 ( .A1(n14827), .A2(n6962), .ZN(n14852) );
  NOR2_X1 U9290 ( .A1(n11021), .A2(n6963), .ZN(n14829) );
  OAI21_X1 U9291 ( .B1(n13227), .B2(n14863), .A(n14834), .ZN(n6758) );
  NAND3_X1 U9292 ( .A1(n7125), .A2(n10071), .A3(P3_REG2_REG_7__SCAN_IN), .ZN(
        n7126) );
  NOR2_X1 U9293 ( .A1(n12572), .A2(n12571), .ZN(n12593) );
  NAND2_X1 U9294 ( .A1(n10641), .A2(n11090), .ZN(n11084) );
  INV_X1 U9295 ( .A(n10640), .ZN(n6704) );
  NOR2_X2 U9296 ( .A1(n14977), .A2(n14976), .ZN(n14975) );
  NAND2_X1 U9297 ( .A1(n8646), .A2(n8645), .ZN(n8767) );
  NAND2_X1 U9298 ( .A1(n6587), .A2(n7336), .ZN(n12083) );
  INV_X1 U9299 ( .A(n15020), .ZN(n6713) );
  AOI21_X1 U9300 ( .B1(n12094), .B2(n12088), .A(n12717), .ZN(n12093) );
  OAI22_X2 U9301 ( .A1(n14642), .A2(n10392), .B1(n12186), .B2(n14649), .ZN(
        n10698) );
  NAND2_X1 U9302 ( .A1(n14035), .A2(n11616), .ZN(n14020) );
  NAND2_X1 U9303 ( .A1(n10309), .A2(n12172), .ZN(n10383) );
  NAND2_X1 U9304 ( .A1(n13956), .A2(n13969), .ZN(n13960) );
  NAND2_X1 U9305 ( .A1(n14626), .A2(n10700), .ZN(n10701) );
  NAND2_X1 U9306 ( .A1(n6762), .A2(n6761), .ZN(n6769) );
  NAND2_X1 U9307 ( .A1(n10675), .A2(n10697), .ZN(n6705) );
  NAND2_X1 U9308 ( .A1(n10662), .A2(n12340), .ZN(n6706) );
  NAND2_X2 U9309 ( .A1(n6786), .A2(n6785), .ZN(n13975) );
  XNOR2_X1 U9310 ( .A(n13779), .B(n14698), .ZN(n12341) );
  NAND2_X1 U9311 ( .A1(n6731), .A2(n11220), .ZN(n11238) );
  NAND2_X1 U9312 ( .A1(n10297), .A2(n12165), .ZN(n10662) );
  NAND2_X1 U9313 ( .A1(n7478), .A2(n10422), .ZN(n14640) );
  NAND2_X1 U9314 ( .A1(n6707), .A2(n11068), .ZN(n11219) );
  NAND2_X1 U9315 ( .A1(n11510), .A2(n11509), .ZN(n14076) );
  NAND2_X1 U9316 ( .A1(n11067), .A2(n11066), .ZN(n6707) );
  NAND2_X1 U9317 ( .A1(n13822), .A2(n13823), .ZN(n13824) );
  NAND2_X1 U9318 ( .A1(n11622), .A2(n12361), .ZN(n13910) );
  NAND2_X1 U9319 ( .A1(n7079), .A2(n7080), .ZN(n11608) );
  NOR2_X1 U9320 ( .A1(n13811), .A2(n13812), .ZN(n13821) );
  NAND3_X1 U9321 ( .A1(n13459), .A2(n6725), .A3(n13458), .ZN(n13547) );
  NOR2_X2 U9322 ( .A1(n12650), .A2(n12854), .ZN(n12666) );
  NOR2_X1 U9323 ( .A1(n15293), .A2(n12607), .ZN(n12637) );
  NOR2_X1 U9324 ( .A1(n12593), .A2(n6520), .ZN(n12595) );
  MUX2_X1 U9325 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n14227), .S(n14788), .Z(
        P1_U3556) );
  INV_X1 U9326 ( .A(n12639), .ZN(n6715) );
  NAND2_X1 U9327 ( .A1(n6744), .A2(n6650), .ZN(n7114) );
  INV_X1 U9328 ( .A(n10701), .ZN(n6724) );
  INV_X1 U9329 ( .A(n12840), .ZN(n6717) );
  AOI21_X1 U9330 ( .B1(n11854), .B2(n12770), .A(n11853), .ZN(n12756) );
  NAND2_X1 U9331 ( .A1(n10095), .A2(n11977), .ZN(n10361) );
  NAND2_X1 U9332 ( .A1(n11848), .A2(n12055), .ZN(n12859) );
  NAND2_X1 U9333 ( .A1(n10366), .A2(n11999), .ZN(n10464) );
  NAND3_X1 U9334 ( .A1(n8596), .A2(n7542), .A3(n8654), .ZN(n8650) );
  OAI21_X1 U9335 ( .B1(n9724), .B2(P3_IR_REG_0__SCAN_IN), .A(n6718), .ZN(n9947) );
  INV_X1 U9336 ( .A(n14698), .ZN(n12163) );
  NAND2_X1 U9337 ( .A1(n6719), .A2(n14698), .ZN(n12165) );
  AND3_X4 U9338 ( .A1(n9368), .A2(n9367), .A3(n6594), .ZN(n14698) );
  INV_X1 U9339 ( .A(n13779), .ZN(n6719) );
  XNOR2_X1 U9340 ( .A(n9415), .B(n9414), .ZN(n9988) );
  NAND2_X1 U9341 ( .A1(n11662), .A2(n7253), .ZN(n6799) );
  NOR2_X1 U9342 ( .A1(n13720), .A2(n6652), .ZN(n13625) );
  OAI21_X1 U9343 ( .B1(n10698), .B2(n10697), .A(n10696), .ZN(n14627) );
  INV_X1 U9344 ( .A(n6792), .ZN(n6791) );
  NAND2_X1 U9345 ( .A1(n6721), .A2(n11192), .ZN(n11240) );
  NAND2_X1 U9346 ( .A1(n7086), .A2(n7087), .ZN(n11622) );
  NAND2_X1 U9347 ( .A1(n11191), .A2(n11190), .ZN(n6721) );
  NAND2_X1 U9348 ( .A1(n13918), .A2(n13912), .ZN(n6730) );
  NAND2_X1 U9349 ( .A1(n10386), .A2(n10385), .ZN(n14642) );
  NAND2_X1 U9350 ( .A1(n8059), .A2(n8058), .ZN(n13368) );
  NAND2_X1 U9351 ( .A1(n7997), .A2(n7996), .ZN(n11341) );
  NAND2_X1 U9352 ( .A1(n7930), .A2(n7929), .ZN(n10897) );
  NAND2_X1 U9353 ( .A1(n7963), .A2(n7962), .ZN(n11226) );
  NAND2_X1 U9354 ( .A1(n10198), .A2(n7859), .ZN(n10728) );
  NAND2_X2 U9355 ( .A1(n6537), .A2(n7740), .ZN(n8162) );
  INV_X1 U9356 ( .A(n11629), .ZN(n14149) );
  NAND2_X1 U9357 ( .A1(n14149), .A2(n6661), .ZN(n14228) );
  OAI21_X1 U9358 ( .B1(n11628), .B2(n14691), .A(n11627), .ZN(n11629) );
  XNOR2_X2 U9359 ( .A(n9317), .B(P1_IR_REG_30__SCAN_IN), .ZN(n9323) );
  OR2_X1 U9360 ( .A1(n7311), .A2(n6833), .ZN(n6834) );
  NAND2_X1 U9361 ( .A1(n7698), .A2(n8111), .ZN(n7701) );
  NAND3_X1 U9362 ( .A1(n12283), .A2(n6727), .A3(n7060), .ZN(n7059) );
  NAND2_X1 U9363 ( .A1(n12278), .A2(n12277), .ZN(n6727) );
  NAND2_X1 U9364 ( .A1(n6728), .A2(n7071), .ZN(n12280) );
  NAND3_X1 U9365 ( .A1(n12273), .A2(n12272), .A3(n6660), .ZN(n6728) );
  NAND2_X1 U9366 ( .A1(n8911), .A2(n8912), .ZN(n8914) );
  NAND2_X1 U9367 ( .A1(n7329), .A2(n7332), .ZN(n8911) );
  NAND2_X1 U9368 ( .A1(n8639), .A2(n8638), .ZN(n8731) );
  NAND2_X1 U9369 ( .A1(n7321), .A2(n7324), .ZN(n8669) );
  XNOR2_X1 U9370 ( .A(n11944), .B(n12700), .ZN(n12106) );
  NAND2_X1 U9371 ( .A1(n12208), .A2(n12209), .ZN(n12207) );
  NOR2_X1 U9372 ( .A1(n7289), .A2(n7066), .ZN(n7065) );
  NAND3_X1 U9373 ( .A1(n12213), .A2(n12212), .A3(n6665), .ZN(n6729) );
  NAND2_X1 U9374 ( .A1(n12140), .A2(n12141), .ZN(n12326) );
  AOI21_X2 U9375 ( .B1(n14136), .B2(n14694), .A(n6649), .ZN(n7022) );
  NAND2_X1 U9376 ( .A1(n6730), .A2(n6645), .ZN(n13915) );
  NAND2_X1 U9377 ( .A1(n10307), .A2(n12166), .ZN(n14655) );
  NAND2_X1 U9378 ( .A1(n11219), .A2(n12355), .ZN(n6731) );
  INV_X1 U9379 ( .A(n14145), .ZN(n11628) );
  AOI21_X1 U9380 ( .B1(P1_REG1_REG_1__SCAN_IN), .B2(n9604), .A(n9642), .ZN(
        n9906) );
  OR2_X1 U9381 ( .A1(n10666), .A2(n14706), .ZN(n14665) );
  NAND2_X1 U9382 ( .A1(n7270), .A2(n7269), .ZN(n14058) );
  NAND2_X1 U9383 ( .A1(n14646), .A2(n12187), .ZN(n14647) );
  NAND2_X1 U9384 ( .A1(n14040), .A2(n14192), .ZN(n14026) );
  NOR2_X2 U9385 ( .A1(n14107), .A2(n14115), .ZN(n14108) );
  OAI21_X1 U9386 ( .B1(n14144), .B2(n14737), .A(n14143), .ZN(n6792) );
  NOR2_X1 U9387 ( .A1(n14388), .A2(n14389), .ZN(n14387) );
  NOR2_X1 U9388 ( .A1(n14585), .A2(n14584), .ZN(n14583) );
  INV_X1 U9389 ( .A(n14596), .ZN(n6736) );
  NAND2_X1 U9390 ( .A1(n15436), .A2(n15437), .ZN(n6738) );
  NOR2_X1 U9391 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n14385), .ZN(n14318) );
  OAI21_X1 U9392 ( .B1(n14593), .B2(n14592), .A(P2_ADDR_REG_15__SCAN_IN), .ZN(
        n6801) );
  NAND2_X1 U9393 ( .A1(n14591), .A2(n6801), .ZN(n14596) );
  XOR2_X1 U9394 ( .A(n12679), .B(n12672), .Z(n12652) );
  INV_X1 U9395 ( .A(n15008), .ZN(n6740) );
  NOR2_X1 U9396 ( .A1(n14942), .A2(n14943), .ZN(n14941) );
  INV_X1 U9397 ( .A(n11124), .ZN(n11126) );
  NOR2_X1 U9398 ( .A1(n15022), .A2(n15021), .ZN(n15020) );
  INV_X1 U9399 ( .A(n12568), .ZN(n12569) );
  INV_X1 U9400 ( .A(n12666), .ZN(n6744) );
  XNOR2_X1 U9401 ( .A(n7112), .B(n7111), .ZN(n12708) );
  OAI21_X1 U9402 ( .B1(n14975), .B2(n10070), .A(n10081), .ZN(n10071) );
  OAI21_X1 U9403 ( .B1(n6931), .B2(n6930), .A(n6927), .ZN(n9229) );
  INV_X1 U9404 ( .A(n9311), .ZN(n9245) );
  NAND2_X1 U9405 ( .A1(n9283), .A2(n13097), .ZN(n13104) );
  NAND2_X1 U9406 ( .A1(n12690), .A2(n12689), .ZN(n7112) );
  NAND2_X1 U9407 ( .A1(n6937), .A2(n13075), .ZN(n13074) );
  NAND2_X1 U9408 ( .A1(n7393), .A2(n7392), .ZN(n9267) );
  NAND2_X1 U9409 ( .A1(n8596), .A2(n7542), .ZN(n8653) );
  NAND2_X1 U9410 ( .A1(n7278), .A2(n7277), .ZN(n7276) );
  NOR2_X1 U9411 ( .A1(n12631), .A2(n6806), .ZN(n12634) );
  AOI22_X1 U9412 ( .A1(n14984), .A2(n14983), .B1(n14986), .B2(n10065), .ZN(
        n15003) );
  AOI21_X1 U9413 ( .B1(n12655), .B2(n14384), .A(n12654), .ZN(n12657) );
  NOR2_X1 U9414 ( .A1(n11135), .A2(n11136), .ZN(n12563) );
  NOR2_X1 U9415 ( .A1(n12694), .A2(n6809), .ZN(n6808) );
  BUF_X4 U9416 ( .A(n8852), .Z(n9031) );
  OAI22_X1 U9417 ( .A1(n11906), .A2(n11940), .B1(n14422), .B2(n12546), .ZN(
        n11921) );
  INV_X1 U9418 ( .A(n14254), .ZN(n14294) );
  INV_X1 U9419 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n6752) );
  NOR2_X1 U9420 ( .A1(P2_ADDR_REG_18__SCAN_IN), .A2(n14403), .ZN(n14407) );
  NAND2_X1 U9421 ( .A1(n13354), .A2(n13364), .ZN(n13353) );
  NAND2_X1 U9422 ( .A1(n7197), .A2(n7196), .ZN(n13395) );
  INV_X1 U9423 ( .A(n10899), .ZN(n6755) );
  NAND2_X1 U9424 ( .A1(n8252), .A2(n8569), .ZN(n13532) );
  OR2_X4 U9425 ( .A1(n6538), .A2(n7740), .ZN(n8176) );
  INV_X1 U9426 ( .A(n6764), .ZN(n8258) );
  NOR2_X1 U9427 ( .A1(n14291), .A2(P1_ADDR_REG_4__SCAN_IN), .ZN(n14259) );
  XNOR2_X1 U9428 ( .A(n7627), .B(SI_3_), .ZN(n7789) );
  OAI21_X2 U9429 ( .B1(n13340), .B2(n7449), .A(n7450), .ZN(n13290) );
  NAND2_X1 U9430 ( .A1(n13291), .A2(n8268), .ZN(n13283) );
  OR2_X2 U9431 ( .A1(n13306), .A2(n13310), .ZN(n8267) );
  NAND2_X2 U9432 ( .A1(n6755), .A2(n8564), .ZN(n10901) );
  NAND4_X2 U9433 ( .A1(n9456), .A2(n9455), .A3(n9454), .A4(n9453), .ZN(n13775)
         );
  NOR2_X2 U9434 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n9168) );
  OAI21_X1 U9435 ( .B1(n8154), .B2(n13017), .A(n8152), .ZN(n7709) );
  NAND2_X1 U9436 ( .A1(n7298), .A2(n7299), .ZN(n7662) );
  NAND2_X1 U9437 ( .A1(n8813), .A2(n8812), .ZN(n8822) );
  NAND2_X1 U9438 ( .A1(n8704), .A2(n8705), .ZN(n8637) );
  AOI21_X2 U9439 ( .B1(n9047), .B2(n11483), .A(n9046), .ZN(n9134) );
  NAND2_X1 U9440 ( .A1(n8677), .A2(n7322), .ZN(n7321) );
  INV_X1 U9441 ( .A(n14007), .ZN(n6762) );
  NOR2_X1 U9442 ( .A1(n14809), .A2(n14808), .ZN(n14807) );
  NOR2_X1 U9443 ( .A1(n14822), .A2(n14821), .ZN(n14820) );
  NAND2_X1 U9444 ( .A1(n11974), .A2(n10150), .ZN(n10035) );
  OAI21_X2 U9445 ( .B1(n12090), .B2(n12733), .A(n12089), .ZN(n11906) );
  NAND2_X1 U9446 ( .A1(n7114), .A2(n7113), .ZN(n12690) );
  NAND2_X1 U9447 ( .A1(n10362), .A2(n11987), .ZN(n15060) );
  NOR2_X2 U9448 ( .A1(n13395), .A2(n8256), .ZN(n6764) );
  AOI21_X2 U9449 ( .B1(n8289), .B2(n13407), .A(n8288), .ZN(n13459) );
  NAND2_X1 U9450 ( .A1(n8245), .A2(n8244), .ZN(n10768) );
  NAND2_X1 U9451 ( .A1(n9475), .A2(n9474), .ZN(n6766) );
  NAND2_X1 U9452 ( .A1(n7189), .A2(n7188), .ZN(n13306) );
  NAND2_X1 U9453 ( .A1(n6811), .A2(n6810), .ZN(n10848) );
  NAND2_X1 U9454 ( .A1(n15426), .A2(n15425), .ZN(n6768) );
  NOR2_X2 U9455 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n9167) );
  AND3_X2 U9456 ( .A1(n6783), .A2(n7935), .A3(n6897), .ZN(n7727) );
  NAND2_X1 U9457 ( .A1(n8271), .A2(n8270), .ZN(n13261) );
  INV_X1 U9458 ( .A(n10850), .ZN(n6811) );
  NAND2_X1 U9459 ( .A1(n7176), .A2(n6771), .ZN(n10564) );
  NAND3_X1 U9460 ( .A1(n14412), .A2(n6997), .A3(P2_ADDR_REG_19__SCAN_IN), .ZN(
        n7614) );
  NAND2_X1 U9461 ( .A1(n7625), .A2(n7624), .ZN(n7790) );
  NAND3_X1 U9462 ( .A1(n10240), .A2(n10239), .A3(n10254), .ZN(n6771) );
  NAND2_X1 U9463 ( .A1(n12792), .A2(n11952), .ZN(n11851) );
  NAND2_X1 U9464 ( .A1(n11850), .A2(n12070), .ZN(n12792) );
  NAND2_X1 U9465 ( .A1(n10464), .A2(n7130), .ZN(n7129) );
  AOI21_X2 U9466 ( .B1(n6581), .B2(n7490), .A(n12733), .ZN(n12740) );
  NAND2_X1 U9467 ( .A1(n13623), .A2(n11699), .ZN(n13693) );
  NAND2_X1 U9468 ( .A1(n10633), .A2(n7219), .ZN(n7217) );
  NAND2_X1 U9469 ( .A1(n13710), .A2(n13711), .ZN(n13709) );
  NAND2_X1 U9470 ( .A1(n7497), .A2(n7500), .ZN(n11547) );
  NAND2_X1 U9471 ( .A1(n14080), .A2(n11610), .ZN(n11510) );
  NAND2_X1 U9472 ( .A1(n6788), .A2(n6787), .ZN(n6786) );
  NAND2_X1 U9473 ( .A1(n14189), .A2(n11560), .ZN(n14007) );
  NAND2_X1 U9474 ( .A1(n6775), .A2(n6774), .ZN(P1_U3523) );
  NAND2_X1 U9475 ( .A1(n14228), .A2(n14774), .ZN(n6775) );
  NAND2_X1 U9476 ( .A1(n10082), .A2(n10081), .ZN(n10080) );
  NAND2_X1 U9477 ( .A1(n6784), .A2(n11016), .ZN(n11067) );
  NOR2_X1 U9478 ( .A1(n10654), .A2(n15127), .ZN(n11100) );
  XNOR2_X1 U9479 ( .A(n7699), .B(SI_24_), .ZN(n8112) );
  INV_X1 U9480 ( .A(n8112), .ZN(n7698) );
  NOR2_X1 U9481 ( .A1(n14939), .A2(n9792), .ZN(n9794) );
  XNOR2_X1 U9482 ( .A(n8183), .B(n8275), .ZN(n13460) );
  OAI21_X2 U9483 ( .B1(n13368), .B2(n7458), .A(n7457), .ZN(n13341) );
  OAI21_X2 U9484 ( .B1(n11341), .B2(n11340), .A(n8014), .ZN(n13424) );
  NOR2_X1 U9485 ( .A1(n13215), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n13222) );
  NAND2_X1 U9486 ( .A1(n13213), .A2(n13214), .ZN(n6778) );
  INV_X1 U9487 ( .A(n13221), .ZN(n6779) );
  OAI21_X1 U9488 ( .B1(n13230), .B2(n14491), .A(n6942), .ZN(P2_U3233) );
  INV_X1 U9489 ( .A(n6899), .ZN(n6783) );
  XNOR2_X2 U9490 ( .A(n8309), .B(n10218), .ZN(n10209) );
  NOR2_X1 U9491 ( .A1(n11085), .A2(n11086), .ZN(n15022) );
  NAND2_X1 U9492 ( .A1(n7129), .A2(n7132), .ZN(n10810) );
  OR2_X2 U9493 ( .A1(n11361), .A2(n11360), .ZN(n11362) );
  OR2_X2 U9494 ( .A1(n15054), .A2(n15075), .ZN(n11987) );
  NAND2_X1 U9495 ( .A1(n11847), .A2(n12050), .ZN(n11848) );
  NAND2_X1 U9496 ( .A1(n10811), .A2(n12013), .ZN(n10937) );
  INV_X1 U9497 ( .A(n11857), .ZN(n6781) );
  INV_X1 U9498 ( .A(n11858), .ZN(n6782) );
  NAND2_X1 U9499 ( .A1(n6782), .A2(n6781), .ZN(P3_U3488) );
  NAND2_X1 U9500 ( .A1(n11173), .A2(n11172), .ZN(n11175) );
  NAND3_X1 U9501 ( .A1(n7819), .A2(n7722), .A3(n7723), .ZN(n6899) );
  NAND2_X1 U9502 ( .A1(n7436), .A2(n7438), .ZN(n10199) );
  INV_X1 U9503 ( .A(n11073), .ZN(n7961) );
  NOR2_X2 U9504 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n9166) );
  NAND2_X1 U9505 ( .A1(n11015), .A2(n12348), .ZN(n6784) );
  INV_X1 U9506 ( .A(n6789), .ZN(P1_U3524) );
  AOI21_X1 U9507 ( .B1(n14227), .B2(n14774), .A(n6790), .ZN(n6789) );
  NOR2_X1 U9508 ( .A1(n14774), .A2(n15240), .ZN(n6790) );
  OR2_X1 U9509 ( .A1(n13658), .A2(n6793), .ZN(P1_U3225) );
  AOI21_X1 U9510 ( .B1(n10452), .B2(n6770), .A(n9372), .ZN(n9374) );
  NAND2_X1 U9511 ( .A1(n7218), .A2(n7222), .ZN(n6797) );
  NAND2_X1 U9512 ( .A1(n9333), .A2(n9336), .ZN(n9350) );
  INV_X1 U9513 ( .A(n14575), .ZN(n7031) );
  INV_X1 U9514 ( .A(n7035), .ZN(n14298) );
  NOR2_X1 U9515 ( .A1(n9045), .A2(n15386), .ZN(n9046) );
  INV_X1 U9516 ( .A(n12709), .ZN(n12926) );
  NAND2_X1 U9517 ( .A1(n8811), .A2(n8810), .ZN(n8813) );
  XNOR2_X1 U9518 ( .A(n11893), .B(n11892), .ZN(n11832) );
  INV_X1 U9519 ( .A(n11856), .ZN(n7555) );
  NAND2_X1 U9520 ( .A1(n7554), .A2(n15056), .ZN(n7550) );
  XNOR2_X1 U9521 ( .A(n6808), .B(n6807), .ZN(n12706) );
  AND2_X1 U9522 ( .A1(n12696), .A2(n12695), .ZN(n6809) );
  NAND3_X1 U9523 ( .A1(n7180), .A2(n7179), .A3(n8243), .ZN(n10544) );
  NOR2_X1 U9524 ( .A1(n10901), .A2(n8567), .ZN(n7173) );
  NAND2_X2 U9525 ( .A1(n11572), .A2(n7626), .ZN(n10388) );
  OAI211_X2 U9526 ( .C1(n11572), .C2(n10306), .A(n10305), .B(n10304), .ZN(
        n14720) );
  OAI21_X1 U9527 ( .B1(n14137), .B2(n14724), .A(n7022), .ZN(n14226) );
  NOR2_X1 U9528 ( .A1(n9789), .A2(n9790), .ZN(n9809) );
  OAI21_X1 U9529 ( .B1(n12561), .B2(n12562), .A(n12587), .ZN(n6820) );
  NAND2_X1 U9530 ( .A1(n7271), .A2(n6673), .ZN(n10653) );
  NAND3_X1 U9531 ( .A1(n6830), .A2(n7615), .A3(P3_ADDR_REG_19__SCAN_IN), .ZN(
        n7617) );
  OAI21_X1 U9532 ( .B1(n14874), .B2(n6830), .A(n13231), .ZN(n6943) );
  NAND2_X1 U9533 ( .A1(n7312), .A2(n7311), .ZN(n7670) );
  OAI211_X1 U9534 ( .C1(n7312), .C2(n6833), .A(n6834), .B(n7004), .ZN(n6835)
         );
  NAND2_X1 U9535 ( .A1(n6839), .A2(n6841), .ZN(n7290) );
  NAND2_X1 U9536 ( .A1(n7294), .A2(n6840), .ZN(n6839) );
  NAND2_X1 U9537 ( .A1(n6844), .A2(n7040), .ZN(n12299) );
  NAND2_X1 U9538 ( .A1(n6845), .A2(n12292), .ZN(n6844) );
  NAND2_X1 U9539 ( .A1(n6846), .A2(n12293), .ZN(n6845) );
  NAND2_X1 U9540 ( .A1(n12296), .A2(n12295), .ZN(n6846) );
  NOR2_X1 U9541 ( .A1(n6854), .A2(n6851), .ZN(n6850) );
  NAND4_X1 U9542 ( .A1(n6852), .A2(n6853), .A3(n8593), .A4(n8825), .ZN(n6851)
         );
  NAND4_X1 U9543 ( .A1(n6858), .A2(n6857), .A3(n6856), .A4(n6855), .ZN(n6854)
         );
  NOR2_X1 U9544 ( .A1(P3_IR_REG_5__SCAN_IN), .A2(P3_IR_REG_8__SCAN_IN), .ZN(
        n6858) );
  NAND2_X1 U9545 ( .A1(n7409), .A2(n6862), .ZN(n6861) );
  AOI21_X1 U9546 ( .B1(n11296), .B2(n7434), .A(n6569), .ZN(n6870) );
  INV_X1 U9547 ( .A(n11296), .ZN(n6872) );
  NAND2_X1 U9548 ( .A1(n8622), .A2(n11352), .ZN(n6879) );
  NAND2_X1 U9549 ( .A1(n12441), .A2(n6544), .ZN(n6885) );
  NAND2_X1 U9550 ( .A1(n6885), .A2(n6886), .ZN(n9003) );
  NAND2_X1 U9551 ( .A1(n6894), .A2(n12479), .ZN(n12411) );
  NAND2_X1 U9552 ( .A1(n8628), .A2(n8630), .ZN(n8634) );
  NAND2_X1 U9553 ( .A1(n8628), .A2(n6895), .ZN(n9100) );
  OR2_X2 U9554 ( .A1(n6899), .A2(n6898), .ZN(n8023) );
  INV_X1 U9555 ( .A(n7935), .ZN(n6898) );
  INV_X1 U9556 ( .A(n6903), .ZN(n10200) );
  NOR2_X2 U9557 ( .A1(n13347), .A2(n13326), .ZN(n13325) );
  NAND2_X1 U9558 ( .A1(n6913), .A2(n6910), .ZN(n13527) );
  AND2_X1 U9559 ( .A1(n7400), .A2(n6916), .ZN(n13272) );
  NAND3_X1 U9560 ( .A1(n13550), .A2(n7400), .A3(n6916), .ZN(n13255) );
  OAI21_X1 U9561 ( .B1(n6918), .B2(n14473), .A(n6919), .ZN(n9283) );
  AOI21_X1 U9562 ( .B1(n7391), .B2(n6928), .A(n6929), .ZN(n6927) );
  NAND2_X1 U9563 ( .A1(n11890), .A2(n9214), .ZN(n6931) );
  INV_X1 U9564 ( .A(n7391), .ZN(n6930) );
  NAND2_X1 U9565 ( .A1(n6932), .A2(n6690), .ZN(P2_U3186) );
  NAND2_X1 U9566 ( .A1(n6933), .A2(n14462), .ZN(n6932) );
  XNOR2_X1 U9567 ( .A(n13039), .B(n6934), .ZN(n6933) );
  NAND2_X1 U9568 ( .A1(n13133), .A2(n6935), .ZN(n13039) );
  NAND3_X1 U9569 ( .A1(n6940), .A2(n13027), .A3(n6938), .ZN(n6937) );
  INV_X1 U9570 ( .A(n13214), .ZN(n6948) );
  INV_X1 U9571 ( .A(n13207), .ZN(n6949) );
  MUX2_X1 U9572 ( .A(P2_REG1_REG_1__SCAN_IN), .B(n9544), .S(n14791), .Z(n14790) );
  NAND2_X1 U9573 ( .A1(n6965), .A2(n6964), .ZN(n8457) );
  INV_X1 U9574 ( .A(n8454), .ZN(n6964) );
  NAND2_X1 U9575 ( .A1(n8456), .A2(n8455), .ZN(n6965) );
  NAND2_X1 U9576 ( .A1(n6966), .A2(n7560), .ZN(n8456) );
  NAND3_X1 U9577 ( .A1(n8446), .A2(n6667), .A3(n8445), .ZN(n6966) );
  OR2_X1 U9578 ( .A1(n8389), .A2(n7579), .ZN(n6970) );
  OAI22_X1 U9579 ( .A1(n8343), .A2(n6971), .B1(n8344), .B2(n6972), .ZN(n8351)
         );
  AOI21_X1 U9580 ( .B1(n8351), .B2(n8350), .A(n8349), .ZN(n8352) );
  OAI21_X1 U9581 ( .B1(n8416), .B2(n7591), .A(n6631), .ZN(n7602) );
  NAND3_X1 U9582 ( .A1(n6982), .A2(n6980), .A3(n6977), .ZN(n6976) );
  OAI21_X1 U9583 ( .B1(n6535), .B2(n7728), .A(n6983), .ZN(n8219) );
  NAND2_X1 U9584 ( .A1(n8427), .A2(n6988), .ZN(n6987) );
  NAND2_X1 U9585 ( .A1(n6987), .A2(n6657), .ZN(n7596) );
  INV_X1 U9586 ( .A(n8430), .ZN(n6996) );
  NAND2_X1 U9587 ( .A1(n7816), .A2(n7634), .ZN(n6998) );
  NAND2_X1 U9588 ( .A1(n7799), .A2(n7798), .ZN(n6999) );
  XNOR2_X2 U9589 ( .A(n7681), .B(SI_18_), .ZN(n8030) );
  NAND3_X1 U9590 ( .A1(n12296), .A2(n12295), .A3(n12294), .ZN(n7040) );
  NAND2_X1 U9591 ( .A1(n7043), .A2(n7041), .ZN(n12268) );
  NAND2_X1 U9592 ( .A1(n12246), .A2(n7044), .ZN(n7043) );
  INV_X1 U9593 ( .A(n12254), .ZN(n7058) );
  NAND2_X1 U9594 ( .A1(n7059), .A2(n7062), .ZN(n12288) );
  AOI21_X1 U9595 ( .B1(n7064), .B2(n7065), .A(n6567), .ZN(P1_U3242) );
  INV_X1 U9596 ( .A(n12380), .ZN(n7064) );
  MUX2_X1 U9597 ( .A(n12162), .B(n12161), .S(n12179), .Z(n12170) );
  NAND2_X1 U9598 ( .A1(n11240), .A2(n7082), .ZN(n7079) );
  OAI21_X2 U9599 ( .B1(n12153), .B2(n12339), .A(n7085), .ZN(n10663) );
  NAND2_X1 U9600 ( .A1(n13960), .A2(n7088), .ZN(n7086) );
  NOR2_X1 U9601 ( .A1(n13950), .A2(n13756), .ZN(n7093) );
  NAND2_X1 U9602 ( .A1(n7103), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8719) );
  NAND2_X1 U9603 ( .A1(n12569), .A2(n12570), .ZN(n7110) );
  NAND2_X1 U9604 ( .A1(n12569), .A2(n7106), .ZN(n7108) );
  AND2_X1 U9605 ( .A1(n7109), .A2(n12570), .ZN(n7106) );
  INV_X1 U9606 ( .A(n7116), .ZN(n9803) );
  NAND2_X1 U9607 ( .A1(n14362), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n7115) );
  NOR2_X1 U9608 ( .A1(n9780), .A2(n9781), .ZN(n9805) );
  NAND2_X1 U9609 ( .A1(n11126), .A2(n7122), .ZN(n7117) );
  NAND2_X1 U9610 ( .A1(n7120), .A2(n7117), .ZN(n12568) );
  NAND3_X1 U9611 ( .A1(n7121), .A2(n11124), .A3(n6565), .ZN(n7120) );
  INV_X1 U9612 ( .A(n7126), .ZN(n14993) );
  INV_X1 U9613 ( .A(n7128), .ZN(n12649) );
  NOR2_X1 U9614 ( .A1(n12637), .A2(n12638), .ZN(n12639) );
  NAND2_X1 U9615 ( .A1(n12859), .A2(n7137), .ZN(n7136) );
  NAND2_X1 U9616 ( .A1(n7136), .A2(n7139), .ZN(n12840) );
  NAND2_X1 U9617 ( .A1(n11362), .A2(n7144), .ZN(n7143) );
  INV_X1 U9618 ( .A(n9947), .ZN(n7146) );
  NAND3_X1 U9619 ( .A1(n7147), .A2(n8689), .A3(n8690), .ZN(n7153) );
  AND2_X1 U9620 ( .A1(n8691), .A2(n8692), .ZN(n7147) );
  NAND2_X1 U9621 ( .A1(n7153), .A2(n9949), .ZN(n10152) );
  NAND2_X1 U9622 ( .A1(n7153), .A2(n9947), .ZN(n11966) );
  NAND2_X1 U9623 ( .A1(P3_U3897), .A2(n7153), .ZN(n7148) );
  NAND2_X1 U9624 ( .A1(n15038), .A2(n7153), .ZN(n7151) );
  AND2_X1 U9625 ( .A1(n12525), .A2(n7153), .ZN(n7152) );
  NAND4_X1 U9626 ( .A1(n7542), .A2(n8596), .A3(n7166), .A4(n8600), .ZN(n13006)
         );
  NAND2_X2 U9627 ( .A1(n7170), .A2(n6538), .ZN(n8488) );
  NAND3_X1 U9628 ( .A1(n7170), .A2(n6538), .A3(P2_REG1_REG_1__SCAN_IN), .ZN(
        n7473) );
  INV_X1 U9629 ( .A(n7173), .ZN(n7171) );
  AOI21_X1 U9630 ( .B1(n7177), .B2(n10254), .A(n6611), .ZN(n7176) );
  NAND2_X1 U9631 ( .A1(n7182), .A2(n7184), .ZN(n7179) );
  NAND2_X1 U9632 ( .A1(n7182), .A2(n8240), .ZN(n7180) );
  OR2_X1 U9633 ( .A1(n8242), .A2(n7187), .ZN(n7186) );
  NAND2_X1 U9634 ( .A1(n13353), .A2(n7190), .ZN(n7189) );
  NAND2_X1 U9635 ( .A1(n13532), .A2(n7198), .ZN(n7197) );
  NAND2_X1 U9636 ( .A1(n13250), .A2(n13249), .ZN(n7204) );
  NAND2_X1 U9637 ( .A1(n8274), .A2(n8273), .ZN(n13247) );
  OAI22_X2 U9638 ( .A1(n10210), .A2(n10209), .B1(n10218), .B2(n7753), .ZN(
        n10240) );
  INV_X1 U9639 ( .A(n8251), .ZN(n13530) );
  NOR2_X1 U9640 ( .A1(n12595), .A2(n12594), .ZN(n12603) );
  XNOR2_X1 U9641 ( .A(n8276), .B(n8275), .ZN(n8289) );
  OAI21_X1 U9642 ( .B1(n7475), .B2(n6538), .A(n7473), .ZN(n7474) );
  NAND2_X1 U9643 ( .A1(n7614), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n7619) );
  NAND2_X2 U9644 ( .A1(n7836), .A2(n7835), .ZN(n10487) );
  NAND2_X1 U9645 ( .A1(n10957), .A2(n10956), .ZN(n10959) );
  NAND2_X1 U9646 ( .A1(n10632), .A2(n10591), .ZN(n7218) );
  NAND2_X1 U9647 ( .A1(n13686), .A2(n7227), .ZN(n7225) );
  AOI21_X1 U9648 ( .B1(n13686), .B2(n13685), .A(n13684), .ZN(n13683) );
  NAND2_X1 U9649 ( .A1(n13745), .A2(n7234), .ZN(n7238) );
  NAND3_X1 U9650 ( .A1(n6745), .A2(n7244), .A3(n7246), .ZN(n7241) );
  INV_X1 U9651 ( .A(n13669), .ZN(n7246) );
  OAI211_X2 U9652 ( .C1(n11262), .C2(n7249), .A(n7247), .B(n11648), .ZN(n13642) );
  OR2_X2 U9653 ( .A1(n11261), .A2(n7249), .ZN(n7247) );
  INV_X1 U9654 ( .A(n11379), .ZN(n7250) );
  NAND2_X1 U9655 ( .A1(n11662), .A2(n6653), .ZN(n7251) );
  NAND2_X1 U9656 ( .A1(n7251), .A2(n7252), .ZN(n13742) );
  NOR2_X1 U9657 ( .A1(n9497), .A2(n7257), .ZN(n7256) );
  NOR2_X2 U9658 ( .A1(n9953), .A2(n9171), .ZN(n7259) );
  INV_X4 U9659 ( .A(n11702), .ZN(n11778) );
  NAND2_X2 U9660 ( .A1(n9443), .A2(n12159), .ZN(n11702) );
  NOR2_X2 U9661 ( .A1(n14636), .A2(n14743), .ZN(n14635) );
  NOR2_X1 U9662 ( .A1(n14666), .A2(n14720), .ZN(n14646) );
  INV_X1 U9663 ( .A(n7264), .ZN(n14107) );
  NOR2_X2 U9664 ( .A1(n14058), .A2(n14197), .ZN(n14040) );
  NAND3_X1 U9665 ( .A1(n7274), .A2(P3_REG1_REG_11__SCAN_IN), .A3(n11119), .ZN(
        n7275) );
  INV_X1 U9666 ( .A(n7275), .ZN(n11120) );
  INV_X1 U9667 ( .A(n7285), .ZN(n9807) );
  INV_X1 U9668 ( .A(n7283), .ZN(n9791) );
  NAND2_X1 U9669 ( .A1(n14362), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n7284) );
  INV_X1 U9670 ( .A(n7288), .ZN(n12628) );
  NAND2_X1 U9671 ( .A1(n7290), .A2(n7293), .ZN(n12333) );
  NAND3_X1 U9672 ( .A1(n12304), .A2(n12303), .A3(n7295), .ZN(n7294) );
  NAND2_X1 U9673 ( .A1(n12306), .A2(n7297), .ZN(n7295) );
  INV_X1 U9674 ( .A(n12306), .ZN(n7296) );
  NAND2_X1 U9675 ( .A1(n7298), .A2(n6564), .ZN(n7663) );
  NAND2_X1 U9676 ( .A1(n7303), .A2(n7622), .ZN(n7625) );
  NAND2_X1 U9677 ( .A1(n7754), .A2(n7755), .ZN(n7302) );
  XNOR2_X1 U9678 ( .A(n7621), .B(SI_1_), .ZN(n7755) );
  NAND2_X1 U9679 ( .A1(n7833), .A2(n7309), .ZN(n7307) );
  NAND2_X1 U9680 ( .A1(n7965), .A2(n7665), .ZN(n7312) );
  NAND3_X1 U9681 ( .A1(n7319), .A2(n7881), .A3(n7318), .ZN(n7316) );
  NAND2_X1 U9682 ( .A1(n7687), .A2(n7686), .ZN(n7689) );
  NAND2_X1 U9683 ( .A1(n8883), .A2(n7330), .ZN(n7329) );
  NAND2_X1 U9684 ( .A1(n8767), .A2(n7343), .ZN(n7340) );
  NAND2_X1 U9685 ( .A1(n7340), .A2(n7341), .ZN(n8790) );
  OAI22_X2 U9686 ( .A1(n7356), .A2(n7355), .B1(P1_DATAO_REG_22__SCAN_IN), .B2(
        n15376), .ZN(n9027) );
  NAND3_X1 U9687 ( .A1(n7360), .A2(n7358), .A3(n12732), .ZN(n12094) );
  NAND3_X1 U9688 ( .A1(n12086), .A2(n6529), .A3(n12085), .ZN(n7360) );
  NAND2_X1 U9689 ( .A1(n13039), .A2(n7381), .ZN(n7380) );
  OAI211_X1 U9690 ( .C1(n13039), .C2(n7382), .A(n7380), .B(n13073), .ZN(
        P2_U3192) );
  AND2_X1 U9691 ( .A1(n9223), .A2(n9218), .ZN(n7391) );
  NAND2_X1 U9692 ( .A1(n11114), .A2(n7394), .ZN(n7393) );
  NAND2_X1 U9693 ( .A1(n10218), .A2(n10358), .ZN(n10236) );
  INV_X2 U9694 ( .A(n10824), .ZN(n10218) );
  NOR2_X2 U9695 ( .A1(n13317), .A2(n13478), .ZN(n7400) );
  XNOR2_X2 U9696 ( .A(n7408), .B(n7735), .ZN(n8278) );
  AND2_X2 U9697 ( .A1(n7727), .A2(n7726), .ZN(n7730) );
  NAND2_X1 U9698 ( .A1(n12400), .A2(n8881), .ZN(n7409) );
  NAND2_X1 U9699 ( .A1(n7421), .A2(n7413), .ZN(n7412) );
  OR2_X1 U9700 ( .A1(n9851), .A2(n8713), .ZN(n7421) );
  INV_X1 U9701 ( .A(n7421), .ZN(n9994) );
  INV_X1 U9702 ( .A(n9995), .ZN(n7420) );
  NAND2_X1 U9703 ( .A1(n7422), .A2(n12533), .ZN(n9162) );
  NAND3_X1 U9704 ( .A1(n7423), .A2(n12123), .A3(n12389), .ZN(n7422) );
  NAND2_X1 U9705 ( .A1(n9142), .A2(n7424), .ZN(n7423) );
  NOR2_X1 U9706 ( .A1(n7425), .A2(n9146), .ZN(n7424) );
  NAND2_X1 U9707 ( .A1(n12126), .A2(n9143), .ZN(n9142) );
  NAND2_X1 U9708 ( .A1(n12447), .A2(n7426), .ZN(n9004) );
  NAND2_X1 U9709 ( .A1(n12509), .A2(n6689), .ZN(n12441) );
  OAI21_X1 U9710 ( .B1(n8805), .B2(n7430), .A(n7428), .ZN(n8821) );
  XNOR2_X1 U9711 ( .A(n8709), .B(n10149), .ZN(n8710) );
  NAND2_X1 U9712 ( .A1(n10222), .A2(n7437), .ZN(n7436) );
  INV_X1 U9713 ( .A(n13368), .ZN(n7461) );
  NAND2_X1 U9714 ( .A1(n7727), .A2(n7466), .ZN(n7468) );
  AOI21_X1 U9715 ( .B1(n7808), .B2(P2_REG0_REG_1__SCAN_IN), .A(n7474), .ZN(
        n7476) );
  INV_X1 U9716 ( .A(n6537), .ZN(n7741) );
  NAND2_X1 U9717 ( .A1(n7752), .A2(n7476), .ZN(n8309) );
  NAND2_X1 U9718 ( .A1(n14640), .A2(n14641), .ZN(n7477) );
  NAND2_X1 U9719 ( .A1(n10421), .A2(n10420), .ZN(n7478) );
  NAND2_X1 U9720 ( .A1(n11238), .A2(n11239), .ZN(n7479) );
  NAND2_X1 U9721 ( .A1(n9364), .A2(n7480), .ZN(n9497) );
  NAND4_X2 U9722 ( .A1(n8702), .A2(n8700), .A3(n8703), .A4(n8701), .ZN(n10041)
         );
  INV_X1 U9723 ( .A(n10153), .ZN(n11965) );
  OR2_X1 U9724 ( .A1(n12781), .A2(n7494), .ZN(n7491) );
  NAND2_X1 U9725 ( .A1(n7491), .A2(n7492), .ZN(n12759) );
  INV_X1 U9726 ( .A(n7503), .ZN(n7498) );
  NOR2_X1 U9727 ( .A1(n11531), .A2(n7505), .ZN(n7504) );
  NAND2_X1 U9728 ( .A1(n7499), .A2(n7503), .ZN(n14049) );
  NAND2_X1 U9729 ( .A1(n6750), .A2(n7504), .ZN(n7499) );
  NAND2_X1 U9730 ( .A1(n7503), .A2(n7502), .ZN(n7501) );
  INV_X1 U9731 ( .A(n7504), .ZN(n7502) );
  OAI21_X1 U9732 ( .B1(n11180), .B2(n7509), .A(n7507), .ZN(n11356) );
  AOI21_X1 U9733 ( .B1(n12836), .B2(n7520), .A(n7517), .ZN(n12806) );
  NAND2_X1 U9734 ( .A1(n13975), .A2(n7528), .ZN(n7526) );
  INV_X1 U9735 ( .A(n13975), .ZN(n7534) );
  NAND2_X1 U9736 ( .A1(n7527), .A2(n7528), .ZN(n13943) );
  NAND2_X1 U9737 ( .A1(n8596), .A2(n8595), .ZN(n8632) );
  OAI21_X1 U9738 ( .B1(n7554), .B2(n7548), .A(n7547), .ZN(n12929) );
  XNOR2_X1 U9739 ( .A(n11836), .B(n7555), .ZN(n7554) );
  NAND2_X1 U9740 ( .A1(n8469), .A2(n7559), .ZN(n7556) );
  INV_X1 U9741 ( .A(n8450), .ZN(n7561) );
  INV_X1 U9742 ( .A(n8365), .ZN(n7562) );
  OAI21_X1 U9743 ( .B1(n8365), .B2(n7568), .A(n7567), .ZN(n8371) );
  AOI21_X1 U9744 ( .B1(n7562), .B2(n7565), .A(n7563), .ZN(n8369) );
  NAND2_X1 U9745 ( .A1(n8462), .A2(n7571), .ZN(n7570) );
  NAND2_X1 U9746 ( .A1(n8389), .A2(n7577), .ZN(n7576) );
  NAND2_X1 U9747 ( .A1(n8377), .A2(n7584), .ZN(n7581) );
  NAND2_X1 U9748 ( .A1(n7581), .A2(n7582), .ZN(n8382) );
  INV_X1 U9749 ( .A(n8375), .ZN(n7587) );
  NAND2_X1 U9750 ( .A1(n8416), .A2(n7590), .ZN(n7588) );
  NAND2_X1 U9751 ( .A1(n7588), .A2(n7589), .ZN(n8421) );
  INV_X1 U9752 ( .A(n8415), .ZN(n7592) );
  NAND3_X1 U9753 ( .A1(n8397), .A2(n6666), .A3(n8396), .ZN(n7600) );
  NAND2_X1 U9754 ( .A1(n9245), .A2(n9244), .ZN(n9310) );
  NAND2_X1 U9755 ( .A1(n8649), .A2(n8648), .ZN(n8811) );
  NAND2_X1 U9756 ( .A1(n8790), .A2(n8789), .ZN(n8649) );
  NAND2_X1 U9757 ( .A1(n12243), .A2(n12242), .ZN(n12246) );
  XNOR2_X1 U9758 ( .A(n9267), .B(n9265), .ZN(n11329) );
  OR2_X1 U9759 ( .A1(P2_DATAO_REG_13__SCAN_IN), .A2(n8863), .ZN(n8864) );
  OR2_X1 U9760 ( .A1(n9116), .A2(n12670), .ZN(n9730) );
  INV_X1 U9761 ( .A(n12457), .ZN(n12473) );
  NAND2_X1 U9762 ( .A1(n9027), .A2(n9026), .ZN(n9030) );
  NAND2_X1 U9763 ( .A1(n7961), .A2(n6605), .ZN(n7963) );
  OR2_X2 U9764 ( .A1(n13778), .A2(n10298), .ZN(n12166) );
  NAND2_X1 U9765 ( .A1(n7617), .A2(n7616), .ZN(n7618) );
  XNOR2_X2 U9766 ( .A(n8719), .B(n8718), .ZN(n14362) );
  NOR2_X1 U9767 ( .A1(n12471), .A2(n12472), .ZN(n7601) );
  OR2_X1 U9768 ( .A1(n11415), .A2(n12552), .ZN(n7603) );
  INV_X1 U9769 ( .A(n13419), .ZN(n14884) );
  AND2_X1 U9770 ( .A1(n8550), .A2(n14491), .ZN(n7604) );
  AND2_X1 U9771 ( .A1(n6531), .A2(n14491), .ZN(n14876) );
  AND2_X1 U9772 ( .A1(n12958), .A2(n12807), .ZN(n7605) );
  OR2_X1 U9773 ( .A1(n13460), .A2(n13393), .ZN(n7606) );
  OR2_X1 U9774 ( .A1(n12728), .A2(n12736), .ZN(n7608) );
  INV_X1 U9775 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n10009) );
  INV_X1 U9776 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n7671) );
  AND2_X1 U9777 ( .A1(n7661), .A2(n7660), .ZN(n7609) );
  INV_X1 U9778 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n7851) );
  AND2_X1 U9779 ( .A1(n9180), .A2(n9179), .ZN(n7610) );
  OR2_X1 U9780 ( .A1(n8371), .A2(n8370), .ZN(n7611) );
  INV_X1 U9781 ( .A(n14674), .ZN(n14113) );
  NAND2_X1 U9782 ( .A1(n9351), .A2(n9332), .ZN(n9335) );
  OR2_X1 U9783 ( .A1(n8456), .A2(n8455), .ZN(n7613) );
  AND2_X1 U9784 ( .A1(n10824), .A2(n8310), .ZN(n8308) );
  AOI21_X1 U9785 ( .B1(n14491), .B2(n11796), .A(n9196), .ZN(n8312) );
  OAI21_X1 U9786 ( .B1(n12191), .B2(n12190), .A(n12189), .ZN(n12193) );
  OR2_X1 U9787 ( .A1(n12198), .A2(n12197), .ZN(n12199) );
  INV_X1 U9788 ( .A(P3_IR_REG_24__SCAN_IN), .ZN(n8597) );
  INV_X1 U9789 ( .A(P3_IR_REG_17__SCAN_IN), .ZN(n8593) );
  INV_X1 U9790 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n9028) );
  INV_X1 U9791 ( .A(n14140), .ZN(n13911) );
  INV_X1 U9792 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n8897) );
  INV_X1 U9793 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n7886) );
  NAND2_X1 U9794 ( .A1(n13911), .A2(n13913), .ZN(n13912) );
  INV_X1 U9795 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n10406) );
  INV_X1 U9796 ( .A(SI_16_), .ZN(n7672) );
  NAND2_X1 U9797 ( .A1(n9053), .A2(n9052), .ZN(n9117) );
  INV_X1 U9798 ( .A(n12028), .ZN(n11172) );
  NAND2_X1 U9799 ( .A1(n10375), .A2(n10374), .ZN(n10466) );
  OR2_X1 U9800 ( .A1(n9070), .A2(n9082), .ZN(n9860) );
  INV_X1 U9801 ( .A(n10269), .ZN(n9223) );
  INV_X1 U9802 ( .A(n9296), .ZN(n9293) );
  INV_X1 U9803 ( .A(n8131), .ZN(n8145) );
  NAND2_X1 U9804 ( .A1(n8048), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8077) );
  INV_X1 U9805 ( .A(n6531), .ZN(n8551) );
  NOR2_X1 U9806 ( .A1(n8305), .A2(n10358), .ZN(n8311) );
  NAND2_X1 U9807 ( .A1(n13139), .A2(n13233), .ZN(n8286) );
  OR2_X1 U9808 ( .A1(n9303), .A2(n9961), .ZN(n10191) );
  INV_X1 U9809 ( .A(n9440), .ZN(n9437) );
  INV_X1 U9810 ( .A(n10014), .ZN(n9393) );
  NAND2_X1 U9811 ( .A1(n11212), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n11503) );
  INV_X1 U9812 ( .A(n11476), .ZN(n11468) );
  INV_X1 U9813 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n15304) );
  OR2_X1 U9814 ( .A1(n10407), .A2(n10406), .ZN(n10705) );
  NAND2_X1 U9815 ( .A1(n7666), .A2(n9705), .ZN(n7669) );
  NOR2_X1 U9816 ( .A1(n14290), .A2(n14289), .ZN(n14268) );
  INV_X1 U9817 ( .A(n12439), .ZN(n8965) );
  AND2_X1 U9818 ( .A1(n9061), .A2(n9060), .ZN(n15345) );
  AND2_X1 U9819 ( .A1(n8796), .A2(n8605), .ZN(n8798) );
  OR2_X1 U9820 ( .A1(n8751), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n8759) );
  INV_X1 U9821 ( .A(n12525), .ZN(n12537) );
  INV_X1 U9822 ( .A(n6525), .ZN(n10144) );
  INV_X1 U9823 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n10275) );
  OR2_X1 U9824 ( .A1(n10142), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n12712) );
  OR2_X1 U9825 ( .A1(n9035), .A2(n9034), .ZN(n9054) );
  NOR2_X1 U9826 ( .A1(n8990), .A2(P3_REG3_REG_21__SCAN_IN), .ZN(n9006) );
  INV_X1 U9827 ( .A(n12550), .ZN(n12863) );
  INV_X1 U9828 ( .A(n12551), .ZN(n12538) );
  OR2_X1 U9829 ( .A1(n12555), .A2(n10756), .ZN(n12013) );
  OR2_X1 U9830 ( .A1(n15036), .A2(n15086), .ZN(n12001) );
  INV_X1 U9831 ( .A(n13001), .ZN(n9939) );
  INV_X1 U9832 ( .A(n11990), .ZN(n15035) );
  AOI21_X1 U9833 ( .B1(n10040), .B2(n10039), .A(n10038), .ZN(n15039) );
  INV_X1 U9834 ( .A(n9271), .ZN(n13024) );
  OR2_X1 U9835 ( .A1(n14474), .A2(n13316), .ZN(n13124) );
  NOR2_X1 U9836 ( .A1(n8088), .A2(n15194), .ZN(n8103) );
  AND2_X1 U9837 ( .A1(n8034), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8048) );
  INV_X1 U9838 ( .A(n8575), .ZN(n13292) );
  INV_X1 U9839 ( .A(n8564), .ZN(n10898) );
  NAND2_X1 U9840 ( .A1(n14884), .A2(n14488), .ZN(n13414) );
  INV_X1 U9841 ( .A(n8566), .ZN(n11228) );
  AND2_X1 U9842 ( .A1(n8489), .A2(n8277), .ZN(n13534) );
  AOI21_X1 U9843 ( .B1(n8209), .B2(n8208), .A(n14886), .ZN(n10194) );
  INV_X1 U9844 ( .A(n14678), .ZN(n13732) );
  INV_X1 U9845 ( .A(n11572), .ZN(n11533) );
  NAND2_X1 U9846 ( .A1(n11696), .A2(n11698), .ZN(n11699) );
  INV_X1 U9847 ( .A(n14159), .ZN(n13950) );
  INV_X1 U9848 ( .A(n12358), .ZN(n14030) );
  OR2_X1 U9849 ( .A1(n14674), .A2(n10314), .ZN(n14089) );
  INV_X1 U9850 ( .A(n12352), .ZN(n11066) );
  INV_X1 U9851 ( .A(n12344), .ZN(n10697) );
  AND2_X1 U9852 ( .A1(n9443), .A2(n9516), .ZN(n9448) );
  OAI21_X1 U9853 ( .B1(n12767), .B2(n12544), .A(n9129), .ZN(n9130) );
  AND2_X1 U9854 ( .A1(n9126), .A2(n15038), .ZN(n12525) );
  INV_X1 U9855 ( .A(n11288), .ZN(n12114) );
  AND2_X1 U9856 ( .A1(n9123), .A2(n9122), .ZN(n12735) );
  INV_X1 U9857 ( .A(n12701), .ZN(n15013) );
  AND2_X1 U9858 ( .A1(n9738), .A2(n9726), .ZN(n9729) );
  AND2_X1 U9859 ( .A1(P3_U3897), .A2(n9116), .ZN(n15015) );
  INV_X1 U9860 ( .A(n12868), .ZN(n15058) );
  AND3_X1 U9861 ( .A1(n9863), .A2(n9862), .A3(n9861), .ZN(n9943) );
  INV_X1 U9862 ( .A(n14422), .ZN(n14440) );
  INV_X1 U9863 ( .A(n12050), .ZN(n11935) );
  INV_X1 U9864 ( .A(n12889), .ZN(n15094) );
  INV_X1 U9865 ( .A(n9722), .ZN(n9934) );
  OR3_X1 U9866 ( .A1(n13597), .A2(n11426), .A3(n11349), .ZN(n9163) );
  AND2_X1 U9867 ( .A1(n7973), .A2(n7742), .ZN(n7988) );
  AND2_X1 U9868 ( .A1(n9963), .A2(n9292), .ZN(n14462) );
  OR2_X1 U9869 ( .A1(n9551), .A2(n9550), .ZN(n14863) );
  INV_X1 U9870 ( .A(n14834), .ZN(n14868) );
  INV_X1 U9871 ( .A(n14863), .ZN(n14853) );
  AND2_X1 U9872 ( .A1(n9291), .A2(n8284), .ZN(n13401) );
  AND2_X1 U9873 ( .A1(n14884), .A2(n13229), .ZN(n13444) );
  AND2_X1 U9874 ( .A1(n9290), .A2(n9289), .ZN(n14899) );
  INV_X1 U9875 ( .A(n13519), .ZN(n14515) );
  OR2_X1 U9876 ( .A1(n8207), .A2(n13597), .ZN(n14886) );
  INV_X1 U9877 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n8205) );
  AND2_X1 U9878 ( .A1(n7820), .A2(n7936), .ZN(n9667) );
  AND2_X1 U9879 ( .A1(n13601), .A2(n14742), .ZN(n14533) );
  OR2_X1 U9880 ( .A1(n14606), .A2(n9602), .ZN(n14619) );
  INV_X1 U9881 ( .A(n14619), .ZN(n13866) );
  OR2_X1 U9882 ( .A1(n14606), .A2(n14601), .ZN(n13847) );
  INV_X1 U9883 ( .A(n14663), .ZN(n14109) );
  INV_X1 U9884 ( .A(n14056), .ZN(n14053) );
  AND2_X1 U9885 ( .A1(n14221), .A2(n14126), .ZN(n14127) );
  INV_X1 U9886 ( .A(n14694), .ZN(n14737) );
  INV_X1 U9887 ( .A(n14724), .ZN(n14771) );
  AND2_X1 U9888 ( .A1(n14125), .A2(n14124), .ZN(n14223) );
  INV_X1 U9889 ( .A(n9448), .ZN(n9595) );
  INV_X1 U9890 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n9336) );
  AND2_X1 U9891 ( .A1(n9697), .A2(n9696), .ZN(n11049) );
  AND2_X1 U9892 ( .A1(n9738), .A2(n9737), .ZN(n15001) );
  INV_X1 U9893 ( .A(n9130), .ZN(n9131) );
  NAND2_X1 U9894 ( .A1(n9102), .A2(n9934), .ZN(n12507) );
  INV_X1 U9895 ( .A(n9160), .ZN(n9161) );
  AOI21_X1 U9896 ( .B1(n12726), .B2(n8697), .A(n10147), .ZN(n12736) );
  INV_X1 U9897 ( .A(P3_ADDR_REG_5__SCAN_IN), .ZN(n14974) );
  OR2_X1 U9898 ( .A1(n9731), .A2(n9730), .ZN(n15023) );
  AND2_X1 U9899 ( .A1(n10821), .A2(n10625), .ZN(n12873) );
  INV_X1 U9900 ( .A(n15131), .ZN(n15129) );
  INV_X1 U9901 ( .A(n12118), .ZN(n12937) );
  AND3_X1 U9902 ( .A1(n14446), .A2(n14445), .A3(n14444), .ZN(n14454) );
  AND3_X1 U9903 ( .A1(n15098), .A2(n15097), .A3(n15096), .ZN(n15126) );
  AND2_X2 U9904 ( .A1(n9935), .A2(n9934), .ZN(n15110) );
  NAND2_X1 U9905 ( .A1(n9070), .A2(n9856), .ZN(n11891) );
  INV_X1 U9906 ( .A(SI_17_), .ZN(n15158) );
  INV_X1 U9907 ( .A(SI_13_), .ZN(n9527) );
  INV_X2 U9908 ( .A(n14462), .ZN(n14474) );
  OR2_X1 U9909 ( .A1(n7978), .A2(n7977), .ZN(n13148) );
  INV_X1 U9910 ( .A(n14870), .ZN(n14836) );
  INV_X1 U9911 ( .A(n14789), .ZN(n14874) );
  AND2_X1 U9912 ( .A1(n10905), .A2(n10904), .ZN(n14522) );
  NAND2_X1 U9913 ( .A1(n14884), .A2(n14495), .ZN(n13393) );
  INV_X1 U9914 ( .A(n13465), .ZN(n13540) );
  INV_X2 U9915 ( .A(n14929), .ZN(n14930) );
  NAND2_X1 U9916 ( .A1(n14925), .A2(n14899), .ZN(n13573) );
  AND2_X1 U9917 ( .A1(n14522), .A2(n14521), .ZN(n14530) );
  OR2_X1 U9918 ( .A1(n10354), .A2(n10195), .ZN(n14924) );
  NAND2_X1 U9919 ( .A1(n14891), .A2(n14886), .ZN(n14887) );
  OR2_X1 U9920 ( .A1(n9536), .A2(n8214), .ZN(n14893) );
  XNOR2_X1 U9921 ( .A(n8206), .B(n8205), .ZN(n13597) );
  INV_X1 U9922 ( .A(n14491), .ZN(n13229) );
  INV_X1 U9923 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n9591) );
  INV_X1 U9924 ( .A(n14013), .ZN(n14183) );
  OR2_X1 U9925 ( .A1(n11544), .A2(n11543), .ZN(n13762) );
  OR2_X1 U9926 ( .A1(n14606), .A2(n9899), .ZN(n13862) );
  OR2_X1 U9927 ( .A1(n14674), .A2(n11534), .ZN(n14117) );
  OR2_X1 U9928 ( .A1(n14674), .A2(n10525), .ZN(n14095) );
  INV_X1 U9929 ( .A(n14788), .ZN(n14786) );
  INV_X1 U9930 ( .A(n14774), .ZN(n14772) );
  AND2_X2 U9931 ( .A1(n14223), .A2(n14222), .ZN(n14774) );
  INV_X1 U9932 ( .A(n9433), .ZN(n9516) );
  INV_X1 U9933 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n9589) );
  INV_X2 U9934 ( .A(n12548), .ZN(P3_U3897) );
  AND2_X1 U9935 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9537), .ZN(P2_U3947) );
  NAND2_X1 U9936 ( .A1(n7606), .A2(n8297), .ZN(P2_U3236) );
  NOR2_X1 U9937 ( .A1(n9443), .A2(n9433), .ZN(P1_U4016) );
  INV_X1 U9938 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n9477) );
  NAND2_X1 U9939 ( .A1(n9475), .A2(SI_0_), .ZN(n8693) );
  AND2_X1 U9940 ( .A1(P2_DATAO_REG_0__SCAN_IN), .A2(SI_0_), .ZN(n7620) );
  NAND2_X1 U9941 ( .A1(n7626), .A2(n7620), .ZN(n9386) );
  INV_X1 U9942 ( .A(SI_1_), .ZN(n9466) );
  MUX2_X1 U9943 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(P1_DATAO_REG_2__SCAN_IN), 
        .S(n9475), .Z(n7623) );
  XNOR2_X1 U9944 ( .A(n7623), .B(SI_2_), .ZN(n7774) );
  INV_X1 U9945 ( .A(n7774), .ZN(n7622) );
  NAND2_X1 U9946 ( .A1(n7623), .A2(SI_2_), .ZN(n7624) );
  INV_X1 U9947 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n9476) );
  NAND2_X1 U9948 ( .A1(n7790), .A2(n7789), .ZN(n7630) );
  INV_X1 U9949 ( .A(n7627), .ZN(n7628) );
  NAND2_X1 U9950 ( .A1(n7628), .A2(SI_3_), .ZN(n7629) );
  NAND2_X1 U9951 ( .A1(n7630), .A2(n7629), .ZN(n7799) );
  INV_X1 U9952 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n10302) );
  MUX2_X1 U9953 ( .A(n10302), .B(n9494), .S(n6533), .Z(n7631) );
  XNOR2_X1 U9954 ( .A(n7631), .B(SI_4_), .ZN(n7798) );
  INV_X1 U9955 ( .A(n7631), .ZN(n7632) );
  NAND2_X1 U9956 ( .A1(n7632), .A2(SI_4_), .ZN(n7633) );
  MUX2_X1 U9957 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(P1_DATAO_REG_5__SCAN_IN), 
        .S(n9473), .Z(n7635) );
  XNOR2_X1 U9958 ( .A(n7635), .B(SI_5_), .ZN(n7815) );
  INV_X1 U9959 ( .A(n7815), .ZN(n7634) );
  NAND2_X1 U9960 ( .A1(n7635), .A2(SI_5_), .ZN(n7636) );
  XNOR2_X1 U9961 ( .A(n7638), .B(SI_6_), .ZN(n7832) );
  INV_X1 U9962 ( .A(n7832), .ZN(n7637) );
  NAND2_X1 U9963 ( .A1(n7638), .A2(SI_6_), .ZN(n7639) );
  MUX2_X1 U9964 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(P1_DATAO_REG_7__SCAN_IN), 
        .S(n9473), .Z(n7640) );
  XNOR2_X1 U9965 ( .A(n7640), .B(SI_7_), .ZN(n7844) );
  MUX2_X1 U9966 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(P1_DATAO_REG_8__SCAN_IN), 
        .S(n6533), .Z(n7642) );
  XNOR2_X1 U9967 ( .A(n7642), .B(SI_8_), .ZN(n7860) );
  INV_X1 U9968 ( .A(n7860), .ZN(n7641) );
  NAND2_X1 U9969 ( .A1(n7642), .A2(SI_8_), .ZN(n7643) );
  MUX2_X1 U9970 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(P1_DATAO_REG_9__SCAN_IN), 
        .S(n9475), .Z(n7646) );
  MUX2_X1 U9971 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(P1_DATAO_REG_10__SCAN_IN), 
        .S(n9473), .Z(n7909) );
  INV_X1 U9972 ( .A(n7909), .ZN(n7647) );
  MUX2_X1 U9973 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(P1_DATAO_REG_11__SCAN_IN), 
        .S(n9473), .Z(n7648) );
  OAI21_X1 U9974 ( .B1(n7647), .B2(n14369), .A(n7913), .ZN(n7653) );
  NOR2_X1 U9975 ( .A1(n7909), .A2(SI_10_), .ZN(n7651) );
  INV_X1 U9976 ( .A(n7648), .ZN(n7649) );
  INV_X1 U9977 ( .A(SI_11_), .ZN(n9483) );
  NAND2_X1 U9978 ( .A1(n7649), .A2(n9483), .ZN(n7912) );
  INV_X1 U9979 ( .A(n7912), .ZN(n7650) );
  AOI21_X1 U9980 ( .B1(n7651), .B2(n7913), .A(n7650), .ZN(n7652) );
  MUX2_X1 U9981 ( .A(n9589), .B(n9591), .S(n9473), .Z(n7654) );
  INV_X1 U9982 ( .A(n7654), .ZN(n7655) );
  NAND2_X1 U9983 ( .A1(n7655), .A2(SI_12_), .ZN(n7656) );
  MUX2_X1 U9984 ( .A(n8843), .B(n9701), .S(n9473), .Z(n7658) );
  NAND2_X1 U9985 ( .A1(n7658), .A2(n9527), .ZN(n7661) );
  INV_X1 U9986 ( .A(n7658), .ZN(n7659) );
  NAND2_X1 U9987 ( .A1(n7659), .A2(SI_13_), .ZN(n7660) );
  MUX2_X1 U9988 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(P1_DATAO_REG_14__SCAN_IN), 
        .S(n9473), .Z(n7964) );
  MUX2_X1 U9989 ( .A(n8897), .B(n9984), .S(n9473), .Z(n7666) );
  INV_X1 U9990 ( .A(n7666), .ZN(n7667) );
  NAND2_X1 U9991 ( .A1(n7667), .A2(SI_15_), .ZN(n7668) );
  MUX2_X1 U9992 ( .A(n7671), .B(n10009), .S(n9473), .Z(n7673) );
  INV_X1 U9993 ( .A(n7673), .ZN(n7674) );
  NAND2_X1 U9994 ( .A1(n7674), .A2(SI_16_), .ZN(n7675) );
  MUX2_X1 U9995 ( .A(n10178), .B(n10179), .S(n9473), .Z(n7677) );
  INV_X1 U9996 ( .A(n7677), .ZN(n7678) );
  NAND2_X1 U9997 ( .A1(n7678), .A2(SI_17_), .ZN(n7679) );
  MUX2_X1 U9998 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(P1_DATAO_REG_18__SCAN_IN), 
        .S(n9473), .Z(n8028) );
  INV_X1 U9999 ( .A(n7681), .ZN(n7682) );
  MUX2_X1 U10000 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(P1_DATAO_REG_19__SCAN_IN), 
        .S(n9473), .Z(n7684) );
  XNOR2_X1 U10001 ( .A(n7684), .B(SI_19_), .ZN(n8041) );
  INV_X1 U10002 ( .A(n7684), .ZN(n7685) );
  INV_X1 U10003 ( .A(SI_19_), .ZN(n10001) );
  NAND2_X1 U10004 ( .A1(n7685), .A2(n10001), .ZN(n7686) );
  MUX2_X1 U10005 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(P1_DATAO_REG_20__SCAN_IN), 
        .S(n9473), .Z(n8062) );
  INV_X1 U10006 ( .A(n8062), .ZN(n7688) );
  MUX2_X1 U10007 ( .A(n11487), .B(n11045), .S(n9473), .Z(n7690) );
  XNOR2_X1 U10008 ( .A(n7690), .B(SI_21_), .ZN(n8073) );
  INV_X1 U10009 ( .A(n7690), .ZN(n7691) );
  NAND2_X1 U10010 ( .A1(n7691), .A2(SI_21_), .ZN(n7692) );
  MUX2_X1 U10011 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(P1_DATAO_REG_22__SCAN_IN), 
        .S(n9473), .Z(n8095) );
  MUX2_X1 U10012 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(P1_DATAO_REG_23__SCAN_IN), 
        .S(n6533), .Z(n8099) );
  INV_X1 U10013 ( .A(n8099), .ZN(n7693) );
  INV_X1 U10014 ( .A(SI_23_), .ZN(n11042) );
  NAND2_X1 U10015 ( .A1(n7693), .A2(n11042), .ZN(n7695) );
  OAI21_X1 U10016 ( .B1(SI_22_), .B2(n8095), .A(n7695), .ZN(n7694) );
  INV_X1 U10017 ( .A(n8095), .ZN(n8085) );
  INV_X1 U10018 ( .A(SI_22_), .ZN(n8999) );
  NOR2_X1 U10019 ( .A1(n8085), .A2(n8999), .ZN(n7696) );
  AOI22_X1 U10020 ( .A1(n7696), .A2(n7695), .B1(n8099), .B2(SI_23_), .ZN(n7697) );
  MUX2_X1 U10021 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(P1_DATAO_REG_24__SCAN_IN), 
        .S(n6533), .Z(n8111) );
  NAND2_X1 U10022 ( .A1(n7699), .A2(SI_24_), .ZN(n7700) );
  MUX2_X1 U10023 ( .A(n15212), .B(n11427), .S(n9473), .Z(n7702) );
  INV_X1 U10024 ( .A(SI_25_), .ZN(n11353) );
  NAND2_X1 U10025 ( .A1(n7702), .A2(n11353), .ZN(n7705) );
  INV_X1 U10026 ( .A(n7702), .ZN(n7703) );
  NAND2_X1 U10027 ( .A1(n7703), .A2(SI_25_), .ZN(n7704) );
  NAND2_X1 U10028 ( .A1(n7705), .A2(n7704), .ZN(n8126) );
  INV_X1 U10029 ( .A(SI_26_), .ZN(n13021) );
  INV_X1 U10030 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n13595) );
  MUX2_X1 U10031 ( .A(n15197), .B(n13595), .S(n9473), .Z(n8140) );
  INV_X1 U10032 ( .A(SI_27_), .ZN(n13017) );
  INV_X1 U10033 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n11817) );
  INV_X1 U10034 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n15253) );
  MUX2_X1 U10035 ( .A(n11817), .B(n15253), .S(n9473), .Z(n8152) );
  NAND2_X1 U10036 ( .A1(n8154), .A2(n13017), .ZN(n7708) );
  NAND2_X1 U10037 ( .A1(n7709), .A2(n7708), .ZN(n8168) );
  INV_X1 U10038 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n11772) );
  INV_X1 U10039 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n13587) );
  MUX2_X1 U10040 ( .A(n11772), .B(n13587), .S(n9473), .Z(n7710) );
  XNOR2_X1 U10041 ( .A(n7710), .B(SI_28_), .ZN(n8167) );
  INV_X1 U10042 ( .A(SI_28_), .ZN(n13015) );
  NAND2_X1 U10043 ( .A1(n7710), .A2(n13015), .ZN(n7711) );
  INV_X1 U10044 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n12386) );
  INV_X1 U10045 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n13581) );
  MUX2_X1 U10046 ( .A(n12386), .B(n13581), .S(n6533), .Z(n8480) );
  XNOR2_X1 U10047 ( .A(n8480), .B(SI_29_), .ZN(n8478) );
  NOR2_X1 U10048 ( .A1(P2_IR_REG_4__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), .ZN(
        n7717) );
  NOR2_X1 U10049 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n7716) );
  NOR2_X1 U10050 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P2_IR_REG_13__SCAN_IN), 
        .ZN(n7721) );
  NOR2_X1 U10051 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_26__SCAN_IN), 
        .ZN(n7725) );
  NAND2_X2 U10052 ( .A1(n8278), .A2(n9541), .ZN(n7766) );
  INV_X2 U10053 ( .A(n7800), .ZN(n7846) );
  NAND2_X1 U10054 ( .A1(n12385), .A2(n7846), .ZN(n7734) );
  OR2_X1 U10055 ( .A1(n8509), .A2(n13581), .ZN(n7733) );
  XNOR2_X2 U10056 ( .A(n7739), .B(n7738), .ZN(n7740) );
  INV_X2 U10057 ( .A(n8130), .ZN(n8485) );
  NAND2_X1 U10058 ( .A1(n8485), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n7751) );
  NAND2_X1 U10059 ( .A1(n7769), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n7750) );
  NAND2_X1 U10060 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n7824) );
  NOR2_X1 U10061 ( .A1(n7824), .A2(n7823), .ZN(n7837) );
  NAND2_X1 U10062 ( .A1(n7837), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n7852) );
  INV_X1 U10063 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n7872) );
  NAND2_X1 U10064 ( .A1(n7899), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n7922) );
  INV_X1 U10065 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n7921) );
  INV_X1 U10066 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n7940) );
  AND2_X1 U10067 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(P2_REG3_REG_14__SCAN_IN), 
        .ZN(n7742) );
  INV_X1 U10068 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n8008) );
  INV_X1 U10069 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n11432) );
  NAND2_X1 U10070 ( .A1(P2_REG3_REG_21__SCAN_IN), .A2(P2_REG3_REG_20__SCAN_IN), 
        .ZN(n7743) );
  INV_X1 U10071 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n15194) );
  NAND2_X1 U10072 ( .A1(n8103), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n8116) );
  INV_X1 U10073 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n8115) );
  NAND2_X1 U10074 ( .A1(n8132), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n8131) );
  NAND2_X1 U10075 ( .A1(P2_REG3_REG_26__SCAN_IN), .A2(n8145), .ZN(n8159) );
  INV_X1 U10076 ( .A(n8159), .ZN(n7744) );
  NAND2_X1 U10077 ( .A1(n7744), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n8174) );
  INV_X1 U10078 ( .A(n8174), .ZN(n7745) );
  NAND2_X1 U10079 ( .A1(n7745), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n8290) );
  OR2_X1 U10080 ( .A1(n8176), .A2(n8290), .ZN(n7749) );
  INV_X1 U10081 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n7747) );
  OR2_X1 U10082 ( .A1(n8488), .A2(n7747), .ZN(n7748) );
  NAND4_X1 U10083 ( .A1(n7751), .A2(n7750), .A3(n7749), .A4(n7748), .ZN(n13140) );
  XNOR2_X1 U10084 ( .A(n13457), .B(n13140), .ZN(n8578) );
  INV_X1 U10085 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n9528) );
  OR2_X1 U10086 ( .A1(n8130), .A2(n9528), .ZN(n7752) );
  INV_X1 U10087 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n10822) );
  INV_X1 U10088 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n9544) );
  CLKBUF_X2 U10089 ( .A(n8309), .Z(n7753) );
  XNOR2_X1 U10090 ( .A(n7754), .B(n7755), .ZN(n9478) );
  INV_X1 U10091 ( .A(n7756), .ZN(n7757) );
  OR2_X1 U10092 ( .A1(n7766), .A2(n14791), .ZN(n7759) );
  INV_X1 U10093 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n9564) );
  INV_X1 U10094 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n7760) );
  INV_X1 U10095 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n7761) );
  INV_X1 U10096 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n9565) );
  OR2_X1 U10097 ( .A1(n8130), .A2(n9565), .ZN(n7762) );
  INV_X1 U10098 ( .A(n15330), .ZN(n14794) );
  XNOR2_X1 U10099 ( .A(n8693), .B(n15262), .ZN(n13599) );
  MUX2_X1 U10100 ( .A(n14794), .B(n13599), .S(n9535), .Z(n10358) );
  INV_X1 U10101 ( .A(n10358), .ZN(n9960) );
  NAND2_X1 U10102 ( .A1(n8305), .A2(n9960), .ZN(n10208) );
  NAND2_X1 U10103 ( .A1(n10209), .A2(n10208), .ZN(n10207) );
  INV_X1 U10104 ( .A(n7753), .ZN(n7767) );
  NAND2_X1 U10105 ( .A1(n7767), .A2(n10218), .ZN(n7768) );
  NAND2_X1 U10106 ( .A1(n10207), .A2(n7768), .ZN(n10233) );
  NAND2_X1 U10107 ( .A1(n8485), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n7773) );
  INV_X1 U10108 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n13161) );
  OR2_X1 U10109 ( .A1(n8176), .A2(n13161), .ZN(n7772) );
  INV_X1 U10110 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n9545) );
  XNOR2_X1 U10111 ( .A(n7775), .B(n7774), .ZN(n9503) );
  NOR2_X1 U10112 ( .A1(n9503), .A2(n7800), .ZN(n7781) );
  NOR2_X1 U10113 ( .A1(n7756), .A2(n7728), .ZN(n7776) );
  MUX2_X1 U10114 ( .A(n7728), .B(n7776), .S(P2_IR_REG_2__SCAN_IN), .Z(n7777)
         );
  INV_X1 U10115 ( .A(n7777), .ZN(n7779) );
  INV_X1 U10116 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n7778) );
  NAND2_X1 U10117 ( .A1(n7756), .A2(n7778), .ZN(n7793) );
  OAI22_X1 U10118 ( .A1(n7791), .A2(n9493), .B1(n9535), .B2(n13162), .ZN(n7780) );
  OR2_X2 U10119 ( .A1(n7781), .A2(n7780), .ZN(n10474) );
  INV_X1 U10120 ( .A(n10474), .ZN(n10839) );
  NAND2_X1 U10121 ( .A1(n10233), .A2(n10232), .ZN(n10235) );
  INV_X1 U10122 ( .A(n8301), .ZN(n8230) );
  NAND2_X1 U10123 ( .A1(n8230), .A2(n10839), .ZN(n7782) );
  NAND2_X1 U10124 ( .A1(n10235), .A2(n7782), .ZN(n10251) );
  NAND2_X1 U10125 ( .A1(n8485), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n7788) );
  OR2_X1 U10126 ( .A1(n8176), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n7787) );
  INV_X1 U10127 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n7783) );
  OR2_X1 U10128 ( .A1(n8162), .A2(n7783), .ZN(n7786) );
  INV_X1 U10129 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n7784) );
  OR2_X1 U10130 ( .A1(n8488), .A2(n7784), .ZN(n7785) );
  NAND4_X2 U10131 ( .A1(n7788), .A2(n7785), .A3(n7786), .A4(n7787), .ZN(n13159) );
  XNOR2_X1 U10132 ( .A(n7789), .B(n7790), .ZN(n9487) );
  OR2_X1 U10133 ( .A1(n9487), .A2(n7800), .ZN(n7796) );
  INV_X2 U10134 ( .A(n7791), .ZN(n8045) );
  NAND2_X1 U10135 ( .A1(n7793), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7792) );
  MUX2_X1 U10136 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7792), .S(
        P2_IR_REG_3__SCAN_IN), .Z(n7794) );
  NAND2_X2 U10137 ( .A1(n7796), .A2(n7795), .ZN(n13050) );
  INV_X1 U10138 ( .A(n10254), .ZN(n10250) );
  NAND2_X1 U10139 ( .A1(n10251), .A2(n10250), .ZN(n10249) );
  INV_X1 U10140 ( .A(n13050), .ZN(n10831) );
  INV_X1 U10141 ( .A(n13159), .ZN(n8232) );
  NAND2_X1 U10142 ( .A1(n10831), .A2(n8232), .ZN(n7797) );
  NAND2_X1 U10143 ( .A1(n10249), .A2(n7797), .ZN(n10558) );
  XNOR2_X1 U10144 ( .A(n7799), .B(n7798), .ZN(n10303) );
  OR2_X1 U10145 ( .A1(n10303), .A2(n7800), .ZN(n7807) );
  NAND2_X1 U10146 ( .A1(n7802), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7801) );
  MUX2_X1 U10147 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7801), .S(
        P2_IR_REG_4__SCAN_IN), .Z(n7805) );
  INV_X1 U10148 ( .A(n7802), .ZN(n7804) );
  INV_X1 U10149 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n7803) );
  NAND2_X1 U10150 ( .A1(n7804), .A2(n7803), .ZN(n7817) );
  NAND2_X1 U10151 ( .A1(n7805), .A2(n7817), .ZN(n9579) );
  INV_X1 U10152 ( .A(n9579), .ZN(n9547) );
  AOI22_X1 U10153 ( .A1(n8045), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n8044), .B2(
        n9547), .ZN(n7806) );
  NAND2_X1 U10154 ( .A1(n7807), .A2(n7806), .ZN(n14898) );
  NAND2_X1 U10156 ( .A1(n8157), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n7813) );
  INV_X1 U10157 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n10567) );
  OR2_X1 U10158 ( .A1(n8130), .A2(n10567), .ZN(n7812) );
  OAI21_X1 U10159 ( .B1(P2_REG3_REG_4__SCAN_IN), .B2(P2_REG3_REG_3__SCAN_IN), 
        .A(n7824), .ZN(n11883) );
  OR2_X1 U10160 ( .A1(n8176), .A2(n11883), .ZN(n7811) );
  INV_X1 U10161 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n7809) );
  OR2_X1 U10162 ( .A1(n8162), .A2(n7809), .ZN(n7810) );
  NAND4_X1 U10163 ( .A1(n7813), .A2(n7812), .A3(n7811), .A4(n7810), .ZN(n13158) );
  XNOR2_X1 U10164 ( .A(n14898), .B(n13158), .ZN(n10563) );
  INV_X1 U10165 ( .A(n10563), .ZN(n10557) );
  INV_X1 U10166 ( .A(n14898), .ZN(n11884) );
  INV_X1 U10167 ( .A(n13158), .ZN(n8341) );
  NAND2_X1 U10168 ( .A1(n11884), .A2(n8341), .ZN(n7814) );
  NAND2_X1 U10169 ( .A1(n10556), .A2(n7814), .ZN(n10222) );
  XNOR2_X1 U10170 ( .A(n7816), .B(n7815), .ZN(n10389) );
  NAND2_X1 U10171 ( .A1(n10389), .A2(n7846), .ZN(n7822) );
  NAND2_X1 U10172 ( .A1(n7817), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7818) );
  MUX2_X1 U10173 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7818), .S(
        P2_IR_REG_5__SCAN_IN), .Z(n7820) );
  NAND2_X1 U10174 ( .A1(n7819), .A2(n7756), .ZN(n7936) );
  AOI22_X1 U10175 ( .A1(n8045), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n8044), .B2(
        n9667), .ZN(n7821) );
  NAND2_X1 U10176 ( .A1(n8157), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n7830) );
  INV_X1 U10178 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n9532) );
  OR2_X1 U10179 ( .A1(n8130), .A2(n9532), .ZN(n7829) );
  AND2_X1 U10180 ( .A1(n7824), .A2(n7823), .ZN(n7825) );
  OR2_X1 U10181 ( .A1(n7825), .A2(n7837), .ZN(n10506) );
  OR2_X1 U10182 ( .A1(n8176), .A2(n10506), .ZN(n7828) );
  INV_X1 U10183 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n7826) );
  OR2_X1 U10184 ( .A1(n8162), .A2(n7826), .ZN(n7827) );
  NAND4_X1 U10185 ( .A1(n7830), .A2(n7829), .A3(n7828), .A4(n7827), .ZN(n13157) );
  XNOR2_X1 U10186 ( .A(n10479), .B(n13157), .ZN(n8560) );
  INV_X1 U10187 ( .A(n8560), .ZN(n10225) );
  OR2_X1 U10188 ( .A1(n10479), .A2(n13157), .ZN(n7831) );
  NAND2_X1 U10189 ( .A1(n10400), .A2(n7846), .ZN(n7836) );
  NAND2_X1 U10190 ( .A1(n7936), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7834) );
  XNOR2_X1 U10191 ( .A(n7834), .B(P2_IR_REG_6__SCAN_IN), .ZN(n9884) );
  AOI22_X1 U10192 ( .A1(n8045), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n8044), .B2(
        n9884), .ZN(n7835) );
  NAND2_X1 U10193 ( .A1(n8157), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n7843) );
  INV_X1 U10194 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n10517) );
  OR2_X1 U10195 ( .A1(n8130), .A2(n10517), .ZN(n7842) );
  OR2_X1 U10196 ( .A1(n7837), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n7838) );
  NAND2_X1 U10197 ( .A1(n7852), .A2(n7838), .ZN(n10518) );
  OR2_X1 U10198 ( .A1(n8176), .A2(n10518), .ZN(n7841) );
  INV_X1 U10199 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n7839) );
  OR2_X1 U10200 ( .A1(n8162), .A2(n7839), .ZN(n7840) );
  NAND4_X1 U10201 ( .A1(n7843), .A2(n7842), .A3(n7841), .A4(n7840), .ZN(n13156) );
  INV_X1 U10202 ( .A(n13156), .ZN(n10120) );
  XNOR2_X1 U10203 ( .A(n10487), .B(n10120), .ZN(n10185) );
  NAND2_X1 U10204 ( .A1(n10678), .A2(n7846), .ZN(n7849) );
  NAND2_X1 U10205 ( .A1(n7862), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7847) );
  XNOR2_X1 U10206 ( .A(n7847), .B(P2_IR_REG_7__SCAN_IN), .ZN(n14806) );
  AOI22_X1 U10207 ( .A1(n8045), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n8044), .B2(
        n14806), .ZN(n7848) );
  NAND2_X1 U10208 ( .A1(n7849), .A2(n7848), .ZN(n10484) );
  NAND2_X1 U10209 ( .A1(n8157), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n7858) );
  INV_X1 U10210 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n7850) );
  OR2_X1 U10211 ( .A1(n8130), .A2(n7850), .ZN(n7857) );
  NAND2_X1 U10212 ( .A1(n7852), .A2(n7851), .ZN(n7853) );
  NAND2_X1 U10213 ( .A1(n7873), .A2(n7853), .ZN(n10493) );
  OR2_X1 U10214 ( .A1(n8176), .A2(n10493), .ZN(n7856) );
  INV_X1 U10215 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n7854) );
  OR2_X1 U10216 ( .A1(n8162), .A2(n7854), .ZN(n7855) );
  NAND4_X1 U10217 ( .A1(n7858), .A2(n7857), .A3(n7856), .A4(n7855), .ZN(n13155) );
  INV_X1 U10218 ( .A(n13155), .ZN(n10731) );
  XNOR2_X1 U10219 ( .A(n10484), .B(n10731), .ZN(n10201) );
  NAND2_X1 U10220 ( .A1(n10199), .A2(n10201), .ZN(n10198) );
  OR2_X1 U10221 ( .A1(n10484), .A2(n13155), .ZN(n7859) );
  NAND2_X1 U10222 ( .A1(n10684), .A2(n7846), .ZN(n7871) );
  INV_X1 U10223 ( .A(n7862), .ZN(n7864) );
  INV_X1 U10224 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n7863) );
  NAND2_X1 U10225 ( .A1(n7864), .A2(n7863), .ZN(n7866) );
  NAND2_X1 U10226 ( .A1(n7866), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7865) );
  MUX2_X1 U10227 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7865), .S(
        P2_IR_REG_8__SCAN_IN), .Z(n7869) );
  INV_X1 U10228 ( .A(n7866), .ZN(n7868) );
  INV_X1 U10229 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n7867) );
  NAND2_X1 U10230 ( .A1(n7868), .A2(n7867), .ZN(n7896) );
  AOI22_X1 U10231 ( .A1(n8045), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n8044), .B2(
        n14819), .ZN(n7870) );
  NAND2_X1 U10232 ( .A1(n7871), .A2(n7870), .ZN(n10741) );
  NAND2_X1 U10233 ( .A1(n8157), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n7879) );
  INV_X1 U10234 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n10736) );
  OR2_X1 U10235 ( .A1(n8130), .A2(n10736), .ZN(n7878) );
  NAND2_X1 U10236 ( .A1(n7873), .A2(n7872), .ZN(n7874) );
  NAND2_X1 U10237 ( .A1(n7887), .A2(n7874), .ZN(n10735) );
  OR2_X1 U10238 ( .A1(n8176), .A2(n10735), .ZN(n7877) );
  INV_X1 U10239 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n7875) );
  OR2_X1 U10240 ( .A1(n8162), .A2(n7875), .ZN(n7876) );
  NAND4_X1 U10241 ( .A1(n7879), .A2(n7878), .A3(n7877), .A4(n7876), .ZN(n13154) );
  INV_X1 U10242 ( .A(n13154), .ZN(n10546) );
  XNOR2_X1 U10243 ( .A(n10741), .B(n10546), .ZN(n10729) );
  INV_X1 U10244 ( .A(n10729), .ZN(n10727) );
  NAND2_X1 U10245 ( .A1(n10741), .A2(n13154), .ZN(n7880) );
  XNOR2_X1 U10246 ( .A(n7882), .B(n7881), .ZN(n10871) );
  NAND2_X1 U10247 ( .A1(n10871), .A2(n7846), .ZN(n7885) );
  NAND2_X1 U10248 ( .A1(n7896), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7883) );
  XNOR2_X1 U10249 ( .A(n7883), .B(P2_IR_REG_9__SCAN_IN), .ZN(n10168) );
  AOI22_X1 U10250 ( .A1(n8045), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n8044), .B2(
        n10168), .ZN(n7884) );
  NAND2_X1 U10251 ( .A1(n8485), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n7894) );
  INV_X1 U10252 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n9879) );
  OR2_X1 U10253 ( .A1(n8488), .A2(n9879), .ZN(n7893) );
  INV_X1 U10254 ( .A(n7899), .ZN(n7889) );
  NAND2_X1 U10255 ( .A1(n7887), .A2(n7886), .ZN(n7888) );
  NAND2_X1 U10256 ( .A1(n7889), .A2(n7888), .ZN(n10572) );
  OR2_X1 U10257 ( .A1(n8176), .A2(n10572), .ZN(n7892) );
  INV_X1 U10258 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n7890) );
  OR2_X1 U10259 ( .A1(n8162), .A2(n7890), .ZN(n7891) );
  NAND4_X1 U10260 ( .A1(n7894), .A2(n7893), .A3(n7892), .A4(n7891), .ZN(n13153) );
  XNOR2_X1 U10261 ( .A(n10750), .B(n13153), .ZN(n8563) );
  XNOR2_X1 U10262 ( .A(n7895), .B(n7909), .ZN(n7907) );
  XNOR2_X1 U10263 ( .A(n7907), .B(SI_10_), .ZN(n10998) );
  NAND2_X1 U10264 ( .A1(n7916), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7897) );
  XNOR2_X1 U10265 ( .A(n7897), .B(P2_IR_REG_10__SCAN_IN), .ZN(n11026) );
  AOI22_X1 U10266 ( .A1(n8045), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n8044), 
        .B2(n11026), .ZN(n7898) );
  NAND2_X1 U10267 ( .A1(n8157), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n7905) );
  INV_X1 U10268 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n10775) );
  OR2_X1 U10269 ( .A1(n8130), .A2(n10775), .ZN(n7904) );
  OR2_X1 U10270 ( .A1(n7899), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n7900) );
  NAND2_X1 U10271 ( .A1(n7922), .A2(n7900), .ZN(n10774) );
  OR2_X1 U10272 ( .A1(n8176), .A2(n10774), .ZN(n7903) );
  INV_X1 U10273 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n7901) );
  OR2_X1 U10274 ( .A1(n8162), .A2(n7901), .ZN(n7902) );
  NAND4_X1 U10275 ( .A1(n7905), .A2(n7904), .A3(n7903), .A4(n7902), .ZN(n13152) );
  INV_X1 U10276 ( .A(n13152), .ZN(n10545) );
  XNOR2_X1 U10277 ( .A(n10779), .B(n10545), .ZN(n10765) );
  INV_X1 U10278 ( .A(n10765), .ZN(n10767) );
  NAND2_X1 U10279 ( .A1(n10766), .A2(n10765), .ZN(n10764) );
  OR2_X1 U10280 ( .A1(n10779), .A2(n13152), .ZN(n7906) );
  NAND2_X1 U10281 ( .A1(n10764), .A2(n7906), .ZN(n10847) );
  INV_X1 U10282 ( .A(n7907), .ZN(n7908) );
  NAND2_X1 U10283 ( .A1(n7908), .A2(SI_10_), .ZN(n7911) );
  NAND2_X1 U10284 ( .A1(n7895), .A2(n7909), .ZN(n7910) );
  NAND2_X1 U10285 ( .A1(n7911), .A2(n7910), .ZN(n7915) );
  NAND2_X1 U10286 ( .A1(n7913), .A2(n7912), .ZN(n7914) );
  NAND2_X1 U10287 ( .A1(n11048), .A2(n7846), .ZN(n7919) );
  OAI21_X1 U10288 ( .B1(n7916), .B2(P2_IR_REG_10__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n7917) );
  XNOR2_X1 U10289 ( .A(n7917), .B(P2_IR_REG_11__SCAN_IN), .ZN(n11027) );
  AOI22_X1 U10290 ( .A1(n8045), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n11027), 
        .B2(n8044), .ZN(n7918) );
  NAND2_X2 U10291 ( .A1(n7919), .A2(n7918), .ZN(n10860) );
  NAND2_X1 U10292 ( .A1(n8485), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n7927) );
  INV_X1 U10293 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n7920) );
  OR2_X1 U10294 ( .A1(n8162), .A2(n7920), .ZN(n7926) );
  NAND2_X1 U10295 ( .A1(n7922), .A2(n7921), .ZN(n7923) );
  NAND2_X1 U10296 ( .A1(n7941), .A2(n7923), .ZN(n10855) );
  OR2_X1 U10297 ( .A1(n8176), .A2(n10855), .ZN(n7925) );
  INV_X1 U10298 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n11022) );
  OR2_X1 U10299 ( .A1(n8488), .A2(n11022), .ZN(n7924) );
  NAND4_X1 U10300 ( .A1(n7927), .A2(n7926), .A3(n7925), .A4(n7924), .ZN(n13151) );
  NAND2_X1 U10301 ( .A1(n10860), .A2(n13151), .ZN(n7928) );
  NAND2_X1 U10302 ( .A1(n10847), .A2(n7928), .ZN(n7930) );
  OR2_X1 U10303 ( .A1(n10860), .A2(n13151), .ZN(n7929) );
  OR2_X1 U10304 ( .A1(n7932), .A2(n7931), .ZN(n7933) );
  NAND2_X1 U10305 ( .A1(n7934), .A2(n7933), .ZN(n11193) );
  NAND2_X1 U10306 ( .A1(n11193), .A2(n7846), .ZN(n7939) );
  OR2_X1 U10307 ( .A1(n7936), .A2(n6898), .ZN(n7952) );
  NAND2_X1 U10308 ( .A1(n7952), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7937) );
  XNOR2_X1 U10309 ( .A(n7937), .B(P2_IR_REG_12__SCAN_IN), .ZN(n14855) );
  AOI22_X1 U10310 ( .A1(n8045), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n8044), 
        .B2(n14855), .ZN(n7938) );
  NAND2_X1 U10311 ( .A1(n8157), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n7948) );
  INV_X1 U10312 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n11029) );
  OR2_X1 U10313 ( .A1(n8130), .A2(n11029), .ZN(n7947) );
  INV_X1 U10314 ( .A(n7973), .ZN(n7943) );
  NAND2_X1 U10315 ( .A1(n7941), .A2(n7940), .ZN(n7942) );
  NAND2_X1 U10316 ( .A1(n7943), .A2(n7942), .ZN(n10927) );
  OR2_X1 U10317 ( .A1(n8176), .A2(n10927), .ZN(n7946) );
  INV_X1 U10318 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n7944) );
  OR2_X1 U10319 ( .A1(n8162), .A2(n7944), .ZN(n7945) );
  NAND4_X1 U10320 ( .A1(n7948), .A2(n7947), .A3(n7946), .A4(n7945), .ZN(n13150) );
  NOR2_X1 U10321 ( .A1(n14516), .A2(n13150), .ZN(n7949) );
  NAND2_X1 U10322 ( .A1(n14516), .A2(n13150), .ZN(n7950) );
  XNOR2_X1 U10323 ( .A(n7951), .B(n7609), .ZN(n11198) );
  NAND2_X1 U10324 ( .A1(n11198), .A2(n7846), .ZN(n7955) );
  NOR2_X1 U10325 ( .A1(n7952), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n7969) );
  OR2_X1 U10326 ( .A1(n7969), .A2(n7728), .ZN(n7953) );
  XNOR2_X1 U10327 ( .A(n7953), .B(P2_IR_REG_13__SCAN_IN), .ZN(n11165) );
  AOI22_X1 U10328 ( .A1(n8045), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n8044), 
        .B2(n11165), .ZN(n7954) );
  XNOR2_X1 U10329 ( .A(n7973), .B(P2_REG3_REG_13__SCAN_IN), .ZN(n13437) );
  OR2_X1 U10330 ( .A1(n13437), .A2(n8176), .ZN(n7960) );
  INV_X1 U10331 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n13438) );
  OR2_X1 U10332 ( .A1(n8130), .A2(n13438), .ZN(n7959) );
  INV_X1 U10333 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n7956) );
  OR2_X1 U10334 ( .A1(n8162), .A2(n7956), .ZN(n7958) );
  INV_X1 U10335 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n11019) );
  OR2_X1 U10336 ( .A1(n8488), .A2(n11019), .ZN(n7957) );
  NAND4_X1 U10337 ( .A1(n7960), .A2(n7959), .A3(n7958), .A4(n7957), .ZN(n13149) );
  OR2_X1 U10338 ( .A1(n13441), .A2(n13149), .ZN(n7962) );
  NAND2_X1 U10339 ( .A1(n7965), .A2(n7964), .ZN(n7966) );
  NAND2_X1 U10340 ( .A1(n7967), .A2(n7966), .ZN(n11308) );
  NAND2_X1 U10341 ( .A1(n11308), .A2(n7846), .ZN(n7972) );
  INV_X1 U10342 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n7968) );
  NAND2_X1 U10343 ( .A1(n7969), .A2(n7968), .ZN(n7984) );
  NAND2_X1 U10344 ( .A1(n7984), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7970) );
  XNOR2_X1 U10345 ( .A(n7970), .B(P2_IR_REG_14__SCAN_IN), .ZN(n11452) );
  AOI22_X1 U10346 ( .A1(n8045), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n8044), 
        .B2(n11452), .ZN(n7971) );
  AOI21_X1 U10347 ( .B1(n7973), .B2(P2_REG3_REG_13__SCAN_IN), .A(
        P2_REG3_REG_14__SCAN_IN), .ZN(n7974) );
  OR2_X1 U10348 ( .A1(n7988), .A2(n7974), .ZN(n14466) );
  NAND2_X1 U10349 ( .A1(n8485), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n7975) );
  OAI21_X1 U10350 ( .B1(n14466), .B2(n8176), .A(n7975), .ZN(n7978) );
  INV_X1 U10351 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n11162) );
  NAND2_X1 U10352 ( .A1(n7769), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n7976) );
  OAI21_X1 U10353 ( .B1(n8488), .B2(n11162), .A(n7976), .ZN(n7977) );
  INV_X1 U10354 ( .A(n13148), .ZN(n13535) );
  NAND2_X1 U10355 ( .A1(n11233), .A2(n13535), .ZN(n13528) );
  OR2_X1 U10356 ( .A1(n11233), .A2(n13535), .ZN(n7979) );
  NAND2_X1 U10357 ( .A1(n11226), .A2(n11228), .ZN(n7981) );
  OR2_X1 U10358 ( .A1(n11233), .A2(n13148), .ZN(n7980) );
  NAND2_X1 U10359 ( .A1(n7981), .A2(n7980), .ZN(n13525) );
  XNOR2_X1 U10360 ( .A(n7983), .B(n7982), .ZN(n11494) );
  NAND2_X1 U10361 ( .A1(n11494), .A2(n7846), .ZN(n7987) );
  NAND2_X1 U10362 ( .A1(n8000), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7985) );
  XNOR2_X1 U10363 ( .A(n7985), .B(P2_IR_REG_15__SCAN_IN), .ZN(n14867) );
  AOI22_X1 U10364 ( .A1(n8045), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n8044), 
        .B2(n14867), .ZN(n7986) );
  OR2_X1 U10365 ( .A1(n7988), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n7989) );
  NAND2_X1 U10366 ( .A1(n8009), .A2(n7989), .ZN(n14485) );
  INV_X1 U10367 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n7990) );
  OR2_X1 U10368 ( .A1(n8488), .A2(n7990), .ZN(n7993) );
  INV_X1 U10369 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n7991) );
  OR2_X1 U10370 ( .A1(n8130), .A2(n7991), .ZN(n7992) );
  AND2_X1 U10371 ( .A1(n7993), .A2(n7992), .ZN(n7995) );
  NAND2_X1 U10372 ( .A1(n7769), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n7994) );
  OAI211_X1 U10373 ( .C1(n14485), .C2(n8176), .A(n7995), .B(n7994), .ZN(n13147) );
  XNOR2_X1 U10374 ( .A(n14489), .B(n13147), .ZN(n8569) );
  NAND2_X1 U10375 ( .A1(n13525), .A2(n13529), .ZN(n7997) );
  OR2_X1 U10376 ( .A1(n14489), .A2(n13147), .ZN(n7996) );
  XNOR2_X1 U10377 ( .A(n7999), .B(n7998), .ZN(n11499) );
  NAND2_X1 U10378 ( .A1(n11499), .A2(n7846), .ZN(n8007) );
  INV_X1 U10379 ( .A(n8000), .ZN(n8002) );
  INV_X1 U10380 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n8001) );
  NAND2_X1 U10381 ( .A1(n8002), .A2(n8001), .ZN(n8004) );
  NAND2_X1 U10382 ( .A1(n8004), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8003) );
  MUX2_X1 U10383 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8003), .S(
        P2_IR_REG_16__SCAN_IN), .Z(n8005) );
  OR2_X1 U10384 ( .A1(n8004), .A2(P2_IR_REG_16__SCAN_IN), .ZN(n8021) );
  AND2_X1 U10385 ( .A1(n8005), .A2(n8021), .ZN(n11455) );
  AOI22_X1 U10386 ( .A1(n11455), .A2(n8044), .B1(n8045), .B2(
        P1_DATAO_REG_16__SCAN_IN), .ZN(n8006) );
  NAND2_X1 U10387 ( .A1(n8009), .A2(n8008), .ZN(n8010) );
  NAND2_X1 U10388 ( .A1(n8015), .A2(n8010), .ZN(n14483) );
  AOI22_X1 U10389 ( .A1(n8157), .A2(P2_REG1_REG_16__SCAN_IN), .B1(n7769), .B2(
        P2_REG0_REG_16__SCAN_IN), .ZN(n8012) );
  NAND2_X1 U10390 ( .A1(n8485), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n8011) );
  OAI211_X1 U10391 ( .C1(n14483), .C2(n8176), .A(n8012), .B(n8011), .ZN(n13146) );
  NAND2_X1 U10392 ( .A1(n14480), .A2(n13146), .ZN(n8014) );
  OR2_X1 U10393 ( .A1(n14480), .A2(n13146), .ZN(n8013) );
  NAND2_X1 U10394 ( .A1(n8014), .A2(n8013), .ZN(n11340) );
  AND2_X1 U10395 ( .A1(n8015), .A2(n11432), .ZN(n8016) );
  OR2_X1 U10396 ( .A1(n8016), .A2(n8034), .ZN(n13428) );
  AOI22_X1 U10397 ( .A1(n8157), .A2(P2_REG1_REG_17__SCAN_IN), .B1(n8485), .B2(
        P2_REG2_REG_17__SCAN_IN), .ZN(n8018) );
  NAND2_X1 U10398 ( .A1(n7769), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n8017) );
  OAI211_X1 U10399 ( .C1(n13428), .C2(n8176), .A(n8018), .B(n8017), .ZN(n13400) );
  XNOR2_X1 U10400 ( .A(n8020), .B(n8019), .ZN(n11511) );
  NAND2_X1 U10401 ( .A1(n11511), .A2(n7846), .ZN(n8027) );
  NAND2_X1 U10402 ( .A1(n8021), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8022) );
  MUX2_X1 U10403 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8022), .S(
        P2_IR_REG_17__SCAN_IN), .Z(n8024) );
  NAND2_X1 U10404 ( .A1(n8024), .A2(n8023), .ZN(n13211) );
  OAI22_X1 U10405 ( .A1(n13211), .A2(n9535), .B1(n8509), .B2(n10179), .ZN(
        n8025) );
  INV_X1 U10406 ( .A(n8025), .ZN(n8026) );
  INV_X1 U10407 ( .A(n8028), .ZN(n8029) );
  XNOR2_X1 U10408 ( .A(n8030), .B(n8029), .ZN(n11520) );
  NAND2_X1 U10409 ( .A1(n11520), .A2(n7846), .ZN(n8033) );
  NAND2_X1 U10410 ( .A1(n8023), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8031) );
  XNOR2_X1 U10411 ( .A(n8031), .B(P2_IR_REG_18__SCAN_IN), .ZN(n13214) );
  AOI22_X1 U10412 ( .A1(n8045), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n8044), 
        .B2(n13214), .ZN(n8032) );
  NOR2_X1 U10413 ( .A1(n8034), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8035) );
  OR2_X1 U10414 ( .A1(n8048), .A2(n8035), .ZN(n13411) );
  INV_X1 U10415 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n13208) );
  NAND2_X1 U10416 ( .A1(n7769), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n8037) );
  NAND2_X1 U10417 ( .A1(n8485), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n8036) );
  OAI211_X1 U10418 ( .C1(n8488), .C2(n13208), .A(n8037), .B(n8036), .ZN(n8038)
         );
  INV_X1 U10419 ( .A(n8038), .ZN(n8039) );
  OAI21_X1 U10420 ( .B1(n13411), .B2(n8176), .A(n8039), .ZN(n13145) );
  INV_X1 U10421 ( .A(n13145), .ZN(n13054) );
  XNOR2_X1 U10422 ( .A(n13521), .B(n13054), .ZN(n13394) );
  INV_X1 U10423 ( .A(n13394), .ZN(n13399) );
  OR2_X1 U10424 ( .A1(n13521), .A2(n13145), .ZN(n8040) );
  NAND2_X1 U10425 ( .A1(n13396), .A2(n8040), .ZN(n13381) );
  XNOR2_X1 U10426 ( .A(n8042), .B(n8041), .ZN(n11532) );
  NAND2_X1 U10427 ( .A1(n11532), .A2(n7846), .ZN(n8047) );
  XNOR2_X2 U10428 ( .A(n8218), .B(P2_IR_REG_19__SCAN_IN), .ZN(n14491) );
  AOI22_X1 U10429 ( .A1(n8045), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n8044), 
        .B2(n14491), .ZN(n8046) );
  OR2_X1 U10430 ( .A1(n8048), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8049) );
  AND2_X1 U10431 ( .A1(n8077), .A2(n8049), .ZN(n13383) );
  INV_X1 U10432 ( .A(n8176), .ZN(n8050) );
  NAND2_X1 U10433 ( .A1(n13383), .A2(n8050), .ZN(n8056) );
  INV_X1 U10434 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n8053) );
  NAND2_X1 U10435 ( .A1(n7769), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n8052) );
  NAND2_X1 U10436 ( .A1(n8485), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n8051) );
  OAI211_X1 U10437 ( .C1(n8488), .C2(n8053), .A(n8052), .B(n8051), .ZN(n8054)
         );
  INV_X1 U10438 ( .A(n8054), .ZN(n8055) );
  NAND2_X1 U10439 ( .A1(n8056), .A2(n8055), .ZN(n13403) );
  NAND2_X1 U10440 ( .A1(n13516), .A2(n13403), .ZN(n8057) );
  NAND2_X1 U10441 ( .A1(n13381), .A2(n8057), .ZN(n8059) );
  OR2_X1 U10442 ( .A1(n13516), .A2(n13403), .ZN(n8058) );
  NAND2_X1 U10443 ( .A1(n8061), .A2(n8060), .ZN(n8063) );
  NAND2_X1 U10444 ( .A1(n11548), .A2(n7846), .ZN(n8065) );
  INV_X1 U10445 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n11072) );
  OR2_X1 U10446 ( .A1(n8509), .A2(n11072), .ZN(n8064) );
  XNOR2_X1 U10447 ( .A(n8077), .B(P2_REG3_REG_20__SCAN_IN), .ZN(n13376) );
  NAND2_X1 U10448 ( .A1(n13376), .A2(n8050), .ZN(n8071) );
  INV_X1 U10449 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n8068) );
  NAND2_X1 U10450 ( .A1(n7769), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n8067) );
  NAND2_X1 U10451 ( .A1(n8485), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n8066) );
  OAI211_X1 U10452 ( .C1(n8488), .C2(n8068), .A(n8067), .B(n8066), .ZN(n8069)
         );
  INV_X1 U10453 ( .A(n8069), .ZN(n8070) );
  NAND2_X1 U10454 ( .A1(n8071), .A2(n8070), .ZN(n13355) );
  NAND2_X1 U10455 ( .A1(n13511), .A2(n13355), .ZN(n8072) );
  XNOR2_X1 U10456 ( .A(n8074), .B(n8073), .ZN(n11486) );
  NAND2_X1 U10457 ( .A1(n11486), .A2(n7846), .ZN(n8076) );
  OR2_X1 U10458 ( .A1(n8509), .A2(n11045), .ZN(n8075) );
  INV_X1 U10459 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n13093) );
  INV_X1 U10460 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n15385) );
  OAI21_X1 U10461 ( .B1(n8077), .B2(n13093), .A(n15385), .ZN(n8078) );
  NAND2_X1 U10462 ( .A1(n8078), .A2(n8088), .ZN(n13360) );
  OR2_X1 U10463 ( .A1(n13360), .A2(n8176), .ZN(n8083) );
  INV_X1 U10464 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n13361) );
  NAND2_X1 U10465 ( .A1(n8157), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n8080) );
  NAND2_X1 U10466 ( .A1(n7769), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n8079) );
  OAI211_X1 U10467 ( .C1(n8130), .C2(n13361), .A(n8080), .B(n8079), .ZN(n8081)
         );
  INV_X1 U10468 ( .A(n8081), .ZN(n8082) );
  NAND2_X1 U10469 ( .A1(n8083), .A2(n8082), .ZN(n13144) );
  XNOR2_X1 U10470 ( .A(n13359), .B(n13144), .ZN(n13364) );
  OR2_X1 U10471 ( .A1(n13359), .A2(n13144), .ZN(n8084) );
  XNOR2_X1 U10472 ( .A(n11570), .B(n8085), .ZN(n11795) );
  NAND2_X1 U10473 ( .A1(n11795), .A2(n7846), .ZN(n8087) );
  INV_X1 U10474 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n11798) );
  OR2_X1 U10475 ( .A1(n8509), .A2(n11798), .ZN(n8086) );
  NAND2_X2 U10476 ( .A1(n8087), .A2(n8086), .ZN(n13346) );
  AND2_X1 U10477 ( .A1(n8088), .A2(n15194), .ZN(n8089) );
  OR2_X1 U10478 ( .A1(n8089), .A2(n8103), .ZN(n13343) );
  INV_X1 U10479 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n13501) );
  NAND2_X1 U10480 ( .A1(n7769), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n8091) );
  NAND2_X1 U10481 ( .A1(n8485), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n8090) );
  OAI211_X1 U10482 ( .C1(n8488), .C2(n13501), .A(n8091), .B(n8090), .ZN(n8092)
         );
  INV_X1 U10483 ( .A(n8092), .ZN(n8093) );
  OAI21_X1 U10484 ( .B1(n13343), .B2(n8176), .A(n8093), .ZN(n13356) );
  XNOR2_X1 U10485 ( .A(n13346), .B(n13356), .ZN(n8572) );
  NAND2_X1 U10486 ( .A1(n13346), .A2(n13356), .ZN(n8094) );
  NAND2_X1 U10487 ( .A1(n11570), .A2(n8095), .ZN(n8098) );
  NAND2_X1 U10488 ( .A1(n8096), .A2(SI_22_), .ZN(n8097) );
  XNOR2_X1 U10489 ( .A(n8099), .B(SI_23_), .ZN(n8100) );
  NAND2_X1 U10490 ( .A1(n11573), .A2(n7846), .ZN(n8102) );
  OR2_X1 U10491 ( .A1(n8509), .A2(n9028), .ZN(n8101) );
  NAND2_X2 U10492 ( .A1(n8102), .A2(n8101), .ZN(n13326) );
  OR2_X1 U10493 ( .A1(n8103), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n8104) );
  NAND2_X1 U10494 ( .A1(n8116), .A2(n8104), .ZN(n13328) );
  OR2_X1 U10495 ( .A1(n13328), .A2(n8176), .ZN(n8109) );
  INV_X1 U10496 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n13495) );
  NAND2_X1 U10497 ( .A1(n8485), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n8106) );
  NAND2_X1 U10498 ( .A1(n7808), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n8105) );
  OAI211_X1 U10499 ( .C1(n8488), .C2(n13495), .A(n8106), .B(n8105), .ZN(n8107)
         );
  INV_X1 U10500 ( .A(n8107), .ZN(n8108) );
  NAND2_X1 U10501 ( .A1(n8109), .A2(n8108), .ZN(n13143) );
  NAND2_X1 U10502 ( .A1(n13326), .A2(n13143), .ZN(n8557) );
  INV_X1 U10503 ( .A(n8557), .ZN(n8110) );
  OR2_X1 U10504 ( .A1(n13326), .A2(n13143), .ZN(n8558) );
  XNOR2_X1 U10505 ( .A(n8112), .B(n8111), .ZN(n11482) );
  NAND2_X1 U10506 ( .A1(n11482), .A2(n7846), .ZN(n8114) );
  INV_X1 U10507 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n15386) );
  OR2_X1 U10508 ( .A1(n8509), .A2(n15386), .ZN(n8113) );
  NAND2_X1 U10509 ( .A1(n8116), .A2(n8115), .ZN(n8118) );
  INV_X1 U10510 ( .A(n8132), .ZN(n8117) );
  NAND2_X1 U10511 ( .A1(n8118), .A2(n8117), .ZN(n13311) );
  OR2_X1 U10512 ( .A1(n13311), .A2(n8176), .ZN(n8124) );
  INV_X1 U10513 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n8121) );
  NAND2_X1 U10514 ( .A1(n8485), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n8120) );
  NAND2_X1 U10515 ( .A1(n7769), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n8119) );
  OAI211_X1 U10516 ( .C1(n8121), .C2(n8488), .A(n8120), .B(n8119), .ZN(n8122)
         );
  INV_X1 U10517 ( .A(n8122), .ZN(n8123) );
  NAND2_X1 U10518 ( .A1(n8124), .A2(n8123), .ZN(n13295) );
  INV_X1 U10519 ( .A(n13295), .ZN(n13081) );
  XNOR2_X1 U10520 ( .A(n13486), .B(n13081), .ZN(n13310) );
  INV_X1 U10521 ( .A(n13310), .ZN(n8125) );
  NAND2_X1 U10522 ( .A1(n11474), .A2(n7846), .ZN(n8129) );
  OR2_X1 U10523 ( .A1(n8509), .A2(n11427), .ZN(n8128) );
  NAND2_X1 U10524 ( .A1(n8157), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n8136) );
  INV_X1 U10525 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n13298) );
  OR2_X1 U10526 ( .A1(n8130), .A2(n13298), .ZN(n8135) );
  OAI21_X1 U10527 ( .B1(P2_REG3_REG_25__SCAN_IN), .B2(n8132), .A(n8131), .ZN(
        n13297) );
  OR2_X1 U10528 ( .A1(n8176), .A2(n13297), .ZN(n8134) );
  INV_X1 U10529 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n15409) );
  OR2_X1 U10530 ( .A1(n8162), .A2(n15409), .ZN(n8133) );
  NAND4_X1 U10531 ( .A1(n8136), .A2(n8135), .A3(n8134), .A4(n8133), .ZN(n13142) );
  OR2_X1 U10532 ( .A1(n13478), .A2(n13142), .ZN(n8137) );
  NAND2_X1 U10533 ( .A1(n13290), .A2(n8137), .ZN(n8139) );
  NAND2_X1 U10534 ( .A1(n13478), .A2(n13142), .ZN(n8138) );
  XNOR2_X1 U10535 ( .A(n8140), .B(SI_26_), .ZN(n8141) );
  NAND2_X1 U10536 ( .A1(n13593), .A2(n7846), .ZN(n8144) );
  OR2_X1 U10537 ( .A1(n8509), .A2(n13595), .ZN(n8143) );
  NAND2_X1 U10538 ( .A1(n8485), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n8150) );
  INV_X1 U10539 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n15329) );
  OR2_X1 U10540 ( .A1(n8488), .A2(n15329), .ZN(n8149) );
  OAI21_X1 U10541 ( .B1(P2_REG3_REG_26__SCAN_IN), .B2(n8145), .A(n8159), .ZN(
        n13280) );
  OR2_X1 U10542 ( .A1(n8176), .A2(n13280), .ZN(n8148) );
  INV_X1 U10543 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n8146) );
  OR2_X1 U10544 ( .A1(n8162), .A2(n8146), .ZN(n8147) );
  NAND4_X1 U10545 ( .A1(n8150), .A2(n8149), .A3(n8148), .A4(n8147), .ZN(n13294) );
  AND2_X1 U10546 ( .A1(n13474), .A2(n13294), .ZN(n8151) );
  XNOR2_X1 U10547 ( .A(n8152), .B(SI_27_), .ZN(n8153) );
  NAND2_X1 U10548 ( .A1(n11595), .A2(n7846), .ZN(n8156) );
  OR2_X1 U10549 ( .A1(n8509), .A2(n15253), .ZN(n8155) );
  NAND2_X1 U10550 ( .A1(n8157), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n8166) );
  INV_X1 U10551 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n13267) );
  OR2_X1 U10552 ( .A1(n8130), .A2(n13267), .ZN(n8165) );
  INV_X1 U10553 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n8158) );
  NAND2_X1 U10554 ( .A1(n8159), .A2(n8158), .ZN(n8160) );
  NAND2_X1 U10555 ( .A1(n8174), .A2(n8160), .ZN(n13266) );
  OR2_X1 U10556 ( .A1(n8176), .A2(n13266), .ZN(n8164) );
  INV_X1 U10557 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n8161) );
  OR2_X1 U10558 ( .A1(n8162), .A2(n8161), .ZN(n8163) );
  NAND4_X1 U10559 ( .A1(n8166), .A2(n8165), .A3(n8164), .A4(n8163), .ZN(n13141) );
  XNOR2_X1 U10560 ( .A(n13469), .B(n13141), .ZN(n13264) );
  OR2_X1 U10561 ( .A1(n8168), .A2(n8167), .ZN(n8169) );
  NAND2_X1 U10562 ( .A1(n13584), .A2(n7846), .ZN(n8172) );
  OR2_X1 U10563 ( .A1(n8509), .A2(n13587), .ZN(n8171) );
  NAND2_X1 U10564 ( .A1(n8485), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n8180) );
  INV_X1 U10565 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n15378) );
  OR2_X1 U10566 ( .A1(n8488), .A2(n15378), .ZN(n8179) );
  INV_X1 U10567 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n8173) );
  NAND2_X1 U10568 ( .A1(n8174), .A2(n8173), .ZN(n8175) );
  NAND2_X1 U10569 ( .A1(n8290), .A2(n8175), .ZN(n13251) );
  OR2_X1 U10570 ( .A1(n8176), .A2(n13251), .ZN(n8178) );
  INV_X1 U10571 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n15135) );
  OR2_X1 U10572 ( .A1(n8162), .A2(n15135), .ZN(n8177) );
  NAND4_X1 U10573 ( .A1(n8180), .A2(n8179), .A3(n8178), .A4(n8177), .ZN(n13065) );
  NAND2_X1 U10574 ( .A1(n13464), .A2(n13065), .ZN(n8182) );
  OR2_X1 U10575 ( .A1(n13464), .A2(n13065), .ZN(n8181) );
  NAND2_X1 U10576 ( .A1(n8182), .A2(n8181), .ZN(n8576) );
  NAND2_X1 U10577 ( .A1(n13245), .A2(n8182), .ZN(n8183) );
  NOR4_X1 U10578 ( .A1(P2_D_REG_13__SCAN_IN), .A2(P2_D_REG_15__SCAN_IN), .A3(
        P2_D_REG_16__SCAN_IN), .A4(P2_D_REG_17__SCAN_IN), .ZN(n8187) );
  NOR4_X1 U10579 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_9__SCAN_IN), .A3(
        P2_D_REG_10__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n8186) );
  NOR4_X1 U10580 ( .A1(P2_D_REG_23__SCAN_IN), .A2(P2_D_REG_24__SCAN_IN), .A3(
        P2_D_REG_25__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n8185) );
  NOR4_X1 U10581 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_20__SCAN_IN), .A3(
        P2_D_REG_21__SCAN_IN), .A4(P2_D_REG_22__SCAN_IN), .ZN(n8184) );
  AND4_X1 U10582 ( .A1(n8187), .A2(n8186), .A3(n8185), .A4(n8184), .ZN(n8209)
         );
  NOR2_X1 U10583 ( .A1(P2_D_REG_6__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .ZN(
        n15352) );
  NOR4_X1 U10584 ( .A1(P2_D_REG_27__SCAN_IN), .A2(P2_D_REG_28__SCAN_IN), .A3(
        P2_D_REG_2__SCAN_IN), .A4(P2_D_REG_19__SCAN_IN), .ZN(n8190) );
  NOR4_X1 U10585 ( .A1(P2_D_REG_3__SCAN_IN), .A2(P2_D_REG_4__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_7__SCAN_IN), .ZN(n8189) );
  NOR4_X1 U10586 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_8__SCAN_IN), .A3(
        P2_D_REG_14__SCAN_IN), .A4(P2_D_REG_29__SCAN_IN), .ZN(n8188) );
  AND4_X1 U10587 ( .A1(n15352), .A2(n8190), .A3(n8189), .A4(n8188), .ZN(n8208)
         );
  NOR2_X1 U10588 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_22__SCAN_IN), 
        .ZN(n8191) );
  AND2_X1 U10589 ( .A1(n8192), .A2(n8191), .ZN(n8193) );
  NAND2_X1 U10590 ( .A1(n6986), .A2(n8193), .ZN(n8212) );
  INV_X1 U10591 ( .A(n8212), .ZN(n8195) );
  NAND2_X1 U10592 ( .A1(n8204), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8198) );
  NAND2_X1 U10593 ( .A1(n8199), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8201) );
  MUX2_X1 U10594 ( .A(n8201), .B(P2_IR_REG_31__SCAN_IN), .S(n8200), .Z(n8202)
         );
  NAND2_X1 U10595 ( .A1(n8202), .A2(n8204), .ZN(n11349) );
  INV_X1 U10596 ( .A(P2_B_REG_SCAN_IN), .ZN(n15296) );
  XOR2_X1 U10597 ( .A(n11349), .B(n15296), .Z(n8203) );
  AND2_X1 U10598 ( .A1(n11426), .A2(n8203), .ZN(n8207) );
  OR2_X1 U10599 ( .A1(n14886), .A2(P2_D_REG_1__SCAN_IN), .ZN(n8211) );
  NAND2_X1 U10600 ( .A1(n13597), .A2(n11426), .ZN(n8210) );
  NAND2_X1 U10601 ( .A1(n8211), .A2(n8210), .ZN(n10190) );
  INV_X1 U10602 ( .A(n10190), .ZN(n9298) );
  NAND2_X1 U10603 ( .A1(n8212), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8213) );
  XNOR2_X1 U10604 ( .A(n8213), .B(P2_IR_REG_23__SCAN_IN), .ZN(n9536) );
  NAND2_X1 U10605 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9163), .ZN(n8214) );
  INV_X1 U10606 ( .A(n14893), .ZN(n14891) );
  NAND2_X1 U10607 ( .A1(n9298), .A2(n14891), .ZN(n8215) );
  OR2_X1 U10608 ( .A1(n10194), .A2(n8215), .ZN(n9288) );
  OR2_X1 U10609 ( .A1(n14886), .A2(P2_D_REG_0__SCAN_IN), .ZN(n8217) );
  NAND2_X1 U10610 ( .A1(n13597), .A2(n11349), .ZN(n8216) );
  NAND2_X1 U10611 ( .A1(n6531), .A2(n13229), .ZN(n9289) );
  INV_X1 U10612 ( .A(n9289), .ZN(n9303) );
  INV_X1 U10613 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n8222) );
  INV_X1 U10614 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n8224) );
  NAND2_X1 U10615 ( .A1(n8589), .A2(n6527), .ZN(n9961) );
  NAND2_X1 U10616 ( .A1(n14890), .A2(n10191), .ZN(n8226) );
  NAND2_X1 U10617 ( .A1(n14923), .A2(n11044), .ZN(n10192) );
  OR2_X2 U10618 ( .A1(n10192), .A2(n14893), .ZN(n14877) );
  OAI21_X4 U10619 ( .B1(n9288), .B2(n8226), .A(n14877), .ZN(n13429) );
  NAND2_X2 U10620 ( .A1(n8228), .A2(n13229), .ZN(n13405) );
  INV_X1 U10621 ( .A(n14883), .ZN(n8229) );
  NAND2_X1 U10622 ( .A1(n13405), .A2(n8229), .ZN(n14495) );
  INV_X1 U10623 ( .A(n13065), .ZN(n13040) );
  INV_X1 U10624 ( .A(n8311), .ZN(n10210) );
  INV_X1 U10625 ( .A(n10232), .ZN(n10239) );
  NAND2_X1 U10626 ( .A1(n8230), .A2(n10474), .ZN(n8231) );
  NAND2_X1 U10627 ( .A1(n10564), .A2(n10563), .ZN(n8234) );
  NAND2_X1 U10628 ( .A1(n14898), .A2(n8341), .ZN(n8233) );
  NAND2_X1 U10629 ( .A1(n8234), .A2(n8233), .ZN(n10226) );
  NAND2_X1 U10630 ( .A1(n10226), .A2(n8560), .ZN(n8237) );
  INV_X1 U10631 ( .A(n13157), .ZN(n8235) );
  NAND2_X1 U10632 ( .A1(n10479), .A2(n8235), .ZN(n8236) );
  INV_X1 U10633 ( .A(n10185), .ZN(n8238) );
  NAND2_X1 U10634 ( .A1(n10487), .A2(n10120), .ZN(n8239) );
  OR2_X1 U10635 ( .A1(n10484), .A2(n10731), .ZN(n8241) );
  OR2_X1 U10636 ( .A1(n10741), .A2(n10546), .ZN(n8243) );
  NAND2_X1 U10637 ( .A1(n10544), .A2(n8563), .ZN(n8245) );
  INV_X1 U10638 ( .A(n13153), .ZN(n10770) );
  OR2_X1 U10639 ( .A1(n10750), .A2(n10770), .ZN(n8244) );
  NAND2_X1 U10640 ( .A1(n10768), .A2(n10767), .ZN(n8247) );
  OR2_X1 U10641 ( .A1(n10779), .A2(n10545), .ZN(n8246) );
  NAND2_X1 U10642 ( .A1(n8247), .A2(n8246), .ZN(n10850) );
  INV_X1 U10643 ( .A(n13151), .ZN(n10769) );
  NAND2_X1 U10644 ( .A1(n10860), .A2(n10769), .ZN(n8248) );
  XNOR2_X1 U10645 ( .A(n14516), .B(n13150), .ZN(n8564) );
  INV_X1 U10646 ( .A(n13150), .ZN(n11078) );
  OR2_X1 U10647 ( .A1(n14516), .A2(n11078), .ZN(n8249) );
  INV_X1 U10648 ( .A(n13149), .ZN(n14459) );
  XNOR2_X1 U10649 ( .A(n13441), .B(n14459), .ZN(n8567) );
  OR2_X1 U10650 ( .A1(n13441), .A2(n14459), .ZN(n8250) );
  NAND2_X1 U10651 ( .A1(n13530), .A2(n13528), .ZN(n8252) );
  INV_X1 U10652 ( .A(n13147), .ZN(n14471) );
  NAND2_X1 U10653 ( .A1(n14489), .A2(n14471), .ZN(n8253) );
  INV_X1 U10654 ( .A(n13146), .ZN(n13537) );
  OR2_X1 U10655 ( .A1(n14480), .A2(n13537), .ZN(n8254) );
  INV_X1 U10656 ( .A(n13400), .ZN(n14468) );
  AND2_X1 U10657 ( .A1(n14498), .A2(n14468), .ZN(n8255) );
  NOR2_X1 U10658 ( .A1(n13521), .A2(n13054), .ZN(n8256) );
  NAND2_X1 U10659 ( .A1(n13521), .A2(n13054), .ZN(n8257) );
  INV_X1 U10660 ( .A(n13403), .ZN(n13372) );
  AND2_X1 U10661 ( .A1(n13516), .A2(n13372), .ZN(n8260) );
  OR2_X1 U10662 ( .A1(n13516), .A2(n13372), .ZN(n8259) );
  INV_X1 U10663 ( .A(n13355), .ZN(n9305) );
  NAND2_X1 U10664 ( .A1(n13511), .A2(n9305), .ZN(n8262) );
  OR2_X1 U10665 ( .A1(n13511), .A2(n9305), .ZN(n8261) );
  NAND2_X1 U10666 ( .A1(n8262), .A2(n8261), .ZN(n13370) );
  INV_X1 U10667 ( .A(n13144), .ZN(n13373) );
  NAND2_X1 U10668 ( .A1(n13359), .A2(n13373), .ZN(n8263) );
  INV_X1 U10669 ( .A(n13356), .ZN(n9304) );
  OR2_X1 U10670 ( .A1(n13346), .A2(n9304), .ZN(n8264) );
  INV_X1 U10671 ( .A(n13143), .ZN(n13086) );
  AND2_X1 U10672 ( .A1(n13326), .A2(n13086), .ZN(n8265) );
  NAND2_X1 U10673 ( .A1(n13486), .A2(n13081), .ZN(n8266) );
  INV_X1 U10674 ( .A(n13142), .ZN(n13125) );
  XNOR2_X1 U10675 ( .A(n13478), .B(n13125), .ZN(n8575) );
  NAND2_X1 U10676 ( .A1(n13293), .A2(n13292), .ZN(n13291) );
  NAND2_X1 U10677 ( .A1(n13478), .A2(n13125), .ZN(n8268) );
  INV_X1 U10678 ( .A(n13294), .ZN(n13080) );
  OR2_X1 U10679 ( .A1(n13474), .A2(n13080), .ZN(n8269) );
  NAND2_X1 U10680 ( .A1(n13283), .A2(n8269), .ZN(n8271) );
  NAND2_X1 U10681 ( .A1(n13474), .A2(n13080), .ZN(n8270) );
  NAND2_X1 U10682 ( .A1(n13261), .A2(n13264), .ZN(n8274) );
  INV_X1 U10683 ( .A(n13141), .ZN(n8272) );
  NAND2_X1 U10684 ( .A1(n13469), .A2(n8272), .ZN(n8273) );
  OAI21_X1 U10685 ( .B1(n13040), .B2(n13464), .A(n13249), .ZN(n8276) );
  NAND2_X1 U10686 ( .A1(n8589), .A2(n14491), .ZN(n8489) );
  NAND2_X1 U10687 ( .A1(n8551), .A2(n8549), .ZN(n8277) );
  INV_X1 U10688 ( .A(n9961), .ZN(n9291) );
  INV_X1 U10689 ( .A(n8278), .ZN(n8284) );
  NAND2_X1 U10690 ( .A1(n13065), .A2(n13401), .ZN(n8287) );
  INV_X1 U10691 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n13454) );
  OR2_X1 U10692 ( .A1(n8488), .A2(n13454), .ZN(n8283) );
  INV_X1 U10693 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n8279) );
  OR2_X1 U10694 ( .A1(n8130), .A2(n8279), .ZN(n8282) );
  INV_X1 U10695 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n15402) );
  OR2_X1 U10696 ( .A1(n8162), .A2(n15402), .ZN(n8281) );
  AND3_X1 U10697 ( .A1(n8283), .A2(n8282), .A3(n8281), .ZN(n8491) );
  INV_X1 U10698 ( .A(n8491), .ZN(n13139) );
  NOR2_X1 U10699 ( .A1(n9541), .A2(n15296), .ZN(n8285) );
  NOR2_X1 U10700 ( .A1(n13538), .A2(n8285), .ZN(n13233) );
  NAND2_X1 U10701 ( .A1(n8287), .A2(n8286), .ZN(n8288) );
  INV_X1 U10702 ( .A(n13464), .ZN(n13550) );
  INV_X1 U10703 ( .A(n14480), .ZN(n14505) );
  INV_X1 U10704 ( .A(n10741), .ZN(n14909) );
  AND2_X1 U10705 ( .A1(n10252), .A2(n10831), .ZN(n10559) );
  INV_X1 U10706 ( .A(n10484), .ZN(n10492) );
  NAND2_X1 U10707 ( .A1(n14909), .A2(n10738), .ZN(n10737) );
  INV_X1 U10708 ( .A(n13441), .ZN(n11079) );
  NOR2_X1 U10709 ( .A1(n14489), .A2(n13527), .ZN(n13526) );
  NAND2_X1 U10710 ( .A1(n14505), .A2(n13526), .ZN(n13425) );
  INV_X1 U10711 ( .A(n13486), .ZN(n13314) );
  NAND2_X1 U10712 ( .A1(n11796), .A2(n11044), .ZN(n10357) );
  AOI211_X1 U10713 ( .C1(n13457), .C2(n13255), .A(n13269), .B(n13239), .ZN(
        n13456) );
  INV_X1 U10714 ( .A(n13457), .ZN(n8293) );
  NOR2_X1 U10715 ( .A1(n10357), .A2(n6531), .ZN(n14488) );
  INV_X1 U10716 ( .A(n8290), .ZN(n8291) );
  INV_X1 U10717 ( .A(n14877), .ZN(n14487) );
  AOI22_X1 U10718 ( .A1(n13419), .A2(P2_REG2_REG_29__SCAN_IN), .B1(n8291), 
        .B2(n14487), .ZN(n8292) );
  OAI21_X1 U10719 ( .B1(n8293), .B2(n13414), .A(n8292), .ZN(n8294) );
  NAND2_X1 U10720 ( .A1(n13474), .A2(n8517), .ZN(n8300) );
  NAND2_X1 U10721 ( .A1(n8298), .A2(n6527), .ZN(n8302) );
  NAND2_X1 U10722 ( .A1(n13294), .A2(n6534), .ZN(n8299) );
  NAND2_X1 U10723 ( .A1(n8300), .A2(n8299), .ZN(n8497) );
  INV_X1 U10724 ( .A(n8497), .ZN(n8501) );
  AOI22_X1 U10725 ( .A1(n8301), .A2(n8302), .B1(n10474), .B2(n8310), .ZN(n8327) );
  NAND2_X1 U10726 ( .A1(n8301), .A2(n8310), .ZN(n8304) );
  NAND2_X1 U10727 ( .A1(n10474), .A2(n8302), .ZN(n8303) );
  NAND2_X1 U10728 ( .A1(n8304), .A2(n8303), .ZN(n8328) );
  INV_X1 U10729 ( .A(n8559), .ZN(n9962) );
  NAND2_X1 U10730 ( .A1(n9962), .A2(n8348), .ZN(n8316) );
  NAND2_X1 U10731 ( .A1(n8309), .A2(n8310), .ZN(n8307) );
  NAND2_X1 U10732 ( .A1(n10824), .A2(n8302), .ZN(n8306) );
  NAND2_X1 U10733 ( .A1(n8307), .A2(n8306), .ZN(n8317) );
  NAND2_X1 U10734 ( .A1(n8317), .A2(n8318), .ZN(n8315) );
  NAND2_X1 U10735 ( .A1(n8311), .A2(n8439), .ZN(n8314) );
  INV_X1 U10736 ( .A(n8553), .ZN(n9196) );
  NAND2_X1 U10737 ( .A1(n8559), .A2(n8312), .ZN(n8313) );
  NAND4_X1 U10738 ( .A1(n8316), .A2(n8315), .A3(n8314), .A4(n8313), .ZN(n8322)
         );
  INV_X1 U10739 ( .A(n8317), .ZN(n8320) );
  INV_X1 U10740 ( .A(n8318), .ZN(n8319) );
  NAND2_X1 U10741 ( .A1(n8320), .A2(n8319), .ZN(n8321) );
  NAND3_X1 U10742 ( .A1(n6617), .A2(n8322), .A3(n8321), .ZN(n8331) );
  NAND2_X1 U10743 ( .A1(n13050), .A2(n8310), .ZN(n8324) );
  NAND2_X1 U10744 ( .A1(n13159), .A2(n8302), .ZN(n8323) );
  AND2_X1 U10745 ( .A1(n8324), .A2(n8323), .ZN(n8333) );
  NAND2_X1 U10746 ( .A1(n13050), .A2(n8302), .ZN(n8326) );
  NAND2_X1 U10747 ( .A1(n13159), .A2(n8310), .ZN(n8325) );
  NAND2_X1 U10748 ( .A1(n8326), .A2(n8325), .ZN(n8332) );
  NAND2_X1 U10749 ( .A1(n8333), .A2(n8332), .ZN(n8330) );
  NAND2_X1 U10750 ( .A1(n8327), .A2(n8328), .ZN(n8329) );
  NAND3_X1 U10751 ( .A1(n8331), .A2(n8330), .A3(n8329), .ZN(n8337) );
  INV_X1 U10752 ( .A(n8332), .ZN(n8335) );
  INV_X1 U10753 ( .A(n8333), .ZN(n8334) );
  NAND2_X1 U10754 ( .A1(n8335), .A2(n8334), .ZN(n8336) );
  NAND2_X1 U10755 ( .A1(n8337), .A2(n8336), .ZN(n8343) );
  NAND2_X1 U10756 ( .A1(n14898), .A2(n8310), .ZN(n8339) );
  NAND2_X1 U10757 ( .A1(n13158), .A2(n8302), .ZN(n8338) );
  NAND2_X1 U10758 ( .A1(n8339), .A2(n8338), .ZN(n8344) );
  NAND2_X1 U10759 ( .A1(n14898), .A2(n6534), .ZN(n8340) );
  OAI21_X1 U10760 ( .B1(n8341), .B2(n8439), .A(n8340), .ZN(n8342) );
  INV_X1 U10761 ( .A(n8344), .ZN(n8345) );
  NAND2_X1 U10762 ( .A1(n10479), .A2(n8302), .ZN(n8347) );
  NAND2_X1 U10763 ( .A1(n13157), .A2(n8517), .ZN(n8346) );
  NAND2_X1 U10764 ( .A1(n8347), .A2(n8346), .ZN(n8350) );
  AOI22_X1 U10765 ( .A1(n10479), .A2(n8517), .B1(n13157), .B2(n6534), .ZN(
        n8349) );
  INV_X1 U10766 ( .A(n8352), .ZN(n8353) );
  NAND2_X1 U10767 ( .A1(n10487), .A2(n8517), .ZN(n8355) );
  NAND2_X1 U10768 ( .A1(n13156), .A2(n8302), .ZN(n8354) );
  NAND2_X1 U10769 ( .A1(n8355), .A2(n8354), .ZN(n8357) );
  AOI22_X1 U10770 ( .A1(n10487), .A2(n6534), .B1(n8517), .B2(n13156), .ZN(
        n8356) );
  AOI21_X1 U10771 ( .B1(n8358), .B2(n8357), .A(n8356), .ZN(n8360) );
  NOR2_X1 U10772 ( .A1(n8358), .A2(n8357), .ZN(n8359) );
  NAND2_X1 U10773 ( .A1(n10484), .A2(n6534), .ZN(n8362) );
  NAND2_X1 U10774 ( .A1(n13155), .A2(n8517), .ZN(n8361) );
  NAND2_X1 U10775 ( .A1(n10484), .A2(n8517), .ZN(n8363) );
  OAI21_X1 U10776 ( .B1(n10731), .B2(n8348), .A(n8363), .ZN(n8364) );
  NAND2_X1 U10777 ( .A1(n10741), .A2(n8517), .ZN(n8367) );
  NAND2_X1 U10778 ( .A1(n13154), .A2(n6534), .ZN(n8366) );
  NAND2_X1 U10779 ( .A1(n8367), .A2(n8366), .ZN(n8370) );
  AOI22_X1 U10780 ( .A1(n10741), .A2(n8302), .B1(n8517), .B2(n13154), .ZN(
        n8368) );
  INV_X1 U10781 ( .A(n8369), .ZN(n8372) );
  NAND2_X1 U10782 ( .A1(n10750), .A2(n6534), .ZN(n8374) );
  NAND2_X1 U10783 ( .A1(n13153), .A2(n8310), .ZN(n8373) );
  NAND2_X1 U10784 ( .A1(n8374), .A2(n8373), .ZN(n8376) );
  AOI22_X1 U10785 ( .A1(n10750), .A2(n8517), .B1(n13153), .B2(n6534), .ZN(
        n8375) );
  NAND2_X1 U10786 ( .A1(n10779), .A2(n8517), .ZN(n8379) );
  NAND2_X1 U10787 ( .A1(n13152), .A2(n6534), .ZN(n8378) );
  NAND2_X1 U10788 ( .A1(n8379), .A2(n8378), .ZN(n8383) );
  NAND2_X1 U10789 ( .A1(n10779), .A2(n6534), .ZN(n8380) );
  OAI21_X1 U10790 ( .B1(n10545), .B2(n8439), .A(n8380), .ZN(n8381) );
  NAND2_X1 U10791 ( .A1(n8382), .A2(n8381), .ZN(n8384) );
  NAND2_X1 U10792 ( .A1(n8384), .A2(n7612), .ZN(n8389) );
  NAND2_X1 U10793 ( .A1(n10860), .A2(n6534), .ZN(n8386) );
  NAND2_X1 U10794 ( .A1(n13151), .A2(n8517), .ZN(n8385) );
  NAND2_X1 U10795 ( .A1(n8386), .A2(n8385), .ZN(n8388) );
  AOI22_X1 U10796 ( .A1(n10860), .A2(n8310), .B1(n13151), .B2(n6534), .ZN(
        n8387) );
  NAND2_X1 U10797 ( .A1(n14516), .A2(n8517), .ZN(n8391) );
  NAND2_X1 U10798 ( .A1(n13150), .A2(n6534), .ZN(n8390) );
  NAND2_X1 U10799 ( .A1(n14516), .A2(n6534), .ZN(n8392) );
  OAI21_X1 U10800 ( .B1(n11078), .B2(n8393), .A(n8392), .ZN(n8394) );
  NAND2_X1 U10801 ( .A1(n8395), .A2(n8394), .ZN(n8397) );
  NAND2_X1 U10802 ( .A1(n13441), .A2(n6534), .ZN(n8399) );
  NAND2_X1 U10803 ( .A1(n13149), .A2(n8517), .ZN(n8398) );
  NAND2_X1 U10804 ( .A1(n8399), .A2(n8398), .ZN(n8401) );
  AOI22_X1 U10805 ( .A1(n13441), .A2(n8310), .B1(n13149), .B2(n6534), .ZN(
        n8400) );
  NAND2_X1 U10806 ( .A1(n11233), .A2(n8517), .ZN(n8403) );
  NAND2_X1 U10807 ( .A1(n13148), .A2(n6534), .ZN(n8402) );
  NAND2_X1 U10808 ( .A1(n8403), .A2(n8402), .ZN(n8408) );
  NAND2_X1 U10809 ( .A1(n8407), .A2(n8408), .ZN(n8406) );
  NAND2_X1 U10810 ( .A1(n11233), .A2(n6534), .ZN(n8404) );
  OAI21_X1 U10811 ( .B1(n13535), .B2(n8439), .A(n8404), .ZN(n8405) );
  NAND2_X1 U10812 ( .A1(n8406), .A2(n8405), .ZN(n8412) );
  INV_X1 U10813 ( .A(n8407), .ZN(n8410) );
  INV_X1 U10814 ( .A(n8408), .ZN(n8409) );
  NAND2_X1 U10815 ( .A1(n8410), .A2(n8409), .ZN(n8411) );
  NAND2_X1 U10816 ( .A1(n14489), .A2(n6534), .ZN(n8414) );
  NAND2_X1 U10817 ( .A1(n13147), .A2(n8310), .ZN(n8413) );
  AOI22_X1 U10818 ( .A1(n14489), .A2(n8310), .B1(n13147), .B2(n6534), .ZN(
        n8415) );
  NAND2_X1 U10819 ( .A1(n14480), .A2(n8310), .ZN(n8418) );
  NAND2_X1 U10820 ( .A1(n13146), .A2(n6534), .ZN(n8417) );
  AOI22_X1 U10821 ( .A1(n14480), .A2(n6534), .B1(n8310), .B2(n13146), .ZN(
        n8419) );
  INV_X1 U10822 ( .A(n8419), .ZN(n8420) );
  NAND2_X1 U10823 ( .A1(n8421), .A2(n8420), .ZN(n8422) );
  NAND2_X1 U10824 ( .A1(n8422), .A2(n7602), .ZN(n8427) );
  NAND2_X1 U10825 ( .A1(n14498), .A2(n6534), .ZN(n8424) );
  NAND2_X1 U10826 ( .A1(n13400), .A2(n8517), .ZN(n8423) );
  NAND2_X1 U10827 ( .A1(n14498), .A2(n8310), .ZN(n8426) );
  NAND2_X1 U10828 ( .A1(n13400), .A2(n6534), .ZN(n8425) );
  NAND2_X1 U10829 ( .A1(n13521), .A2(n8310), .ZN(n8429) );
  NAND2_X1 U10830 ( .A1(n13145), .A2(n6534), .ZN(n8428) );
  NAND2_X1 U10831 ( .A1(n8429), .A2(n8428), .ZN(n8431) );
  AOI22_X1 U10832 ( .A1(n13521), .A2(n6534), .B1(n8310), .B2(n13145), .ZN(
        n8430) );
  NAND2_X1 U10833 ( .A1(n13516), .A2(n6534), .ZN(n8433) );
  NAND2_X1 U10834 ( .A1(n13403), .A2(n8517), .ZN(n8432) );
  NAND2_X1 U10835 ( .A1(n8433), .A2(n8432), .ZN(n8435) );
  AOI22_X1 U10836 ( .A1(n13516), .A2(n8517), .B1(n13403), .B2(n6534), .ZN(
        n8434) );
  AND2_X1 U10837 ( .A1(n13355), .A2(n6534), .ZN(n8436) );
  AOI21_X1 U10838 ( .B1(n13511), .B2(n8310), .A(n8436), .ZN(n8443) );
  INV_X1 U10839 ( .A(n8443), .ZN(n8437) );
  NAND2_X1 U10840 ( .A1(n8442), .A2(n8437), .ZN(n8441) );
  NAND2_X1 U10841 ( .A1(n13511), .A2(n6534), .ZN(n8438) );
  OAI21_X1 U10842 ( .B1(n9305), .B2(n8439), .A(n8438), .ZN(n8440) );
  NAND2_X1 U10843 ( .A1(n8441), .A2(n8440), .ZN(n8446) );
  INV_X1 U10844 ( .A(n8442), .ZN(n8444) );
  NAND2_X1 U10845 ( .A1(n8444), .A2(n8443), .ZN(n8445) );
  AND2_X1 U10846 ( .A1(n13144), .A2(n8517), .ZN(n8447) );
  AOI21_X1 U10847 ( .B1(n13359), .B2(n6534), .A(n8447), .ZN(n8451) );
  INV_X1 U10848 ( .A(n8451), .ZN(n8448) );
  NAND2_X1 U10849 ( .A1(n13359), .A2(n8517), .ZN(n8449) );
  OAI21_X1 U10850 ( .B1(n13373), .B2(n8348), .A(n8449), .ZN(n8450) );
  NAND2_X1 U10851 ( .A1(n13346), .A2(n8517), .ZN(n8453) );
  NAND2_X1 U10852 ( .A1(n13356), .A2(n6534), .ZN(n8452) );
  NAND2_X1 U10853 ( .A1(n8453), .A2(n8452), .ZN(n8455) );
  AOI22_X1 U10854 ( .A1(n13346), .A2(n6534), .B1(n8310), .B2(n13356), .ZN(
        n8454) );
  NAND2_X1 U10855 ( .A1(n8457), .A2(n7613), .ZN(n8462) );
  NAND2_X1 U10856 ( .A1(n13326), .A2(n6534), .ZN(n8459) );
  NAND2_X1 U10857 ( .A1(n13143), .A2(n8517), .ZN(n8458) );
  NAND2_X1 U10858 ( .A1(n8459), .A2(n8458), .ZN(n8461) );
  AOI22_X1 U10859 ( .A1(n13326), .A2(n8310), .B1(n13143), .B2(n6534), .ZN(
        n8460) );
  NAND2_X1 U10860 ( .A1(n13486), .A2(n8517), .ZN(n8464) );
  NAND2_X1 U10861 ( .A1(n13295), .A2(n6534), .ZN(n8463) );
  NAND2_X1 U10862 ( .A1(n13486), .A2(n6534), .ZN(n8466) );
  NAND2_X1 U10863 ( .A1(n13295), .A2(n8310), .ZN(n8465) );
  NAND2_X1 U10864 ( .A1(n8466), .A2(n8465), .ZN(n8467) );
  NAND2_X1 U10865 ( .A1(n13478), .A2(n6534), .ZN(n8471) );
  NAND2_X1 U10866 ( .A1(n13142), .A2(n8517), .ZN(n8470) );
  NAND2_X1 U10867 ( .A1(n8471), .A2(n8470), .ZN(n8474) );
  AOI22_X1 U10868 ( .A1(n13478), .A2(n8310), .B1(n13142), .B2(n6534), .ZN(
        n8472) );
  INV_X1 U10869 ( .A(n8472), .ZN(n8473) );
  INV_X1 U10870 ( .A(n8498), .ZN(n8500) );
  AND2_X1 U10871 ( .A1(n13141), .A2(n8310), .ZN(n8475) );
  AOI21_X1 U10872 ( .B1(n13469), .B2(n6534), .A(n8475), .ZN(n8527) );
  NAND2_X1 U10873 ( .A1(n13469), .A2(n8310), .ZN(n8477) );
  NAND2_X1 U10874 ( .A1(n13141), .A2(n6534), .ZN(n8476) );
  NAND2_X1 U10875 ( .A1(n8477), .A2(n8476), .ZN(n8526) );
  INV_X1 U10876 ( .A(SI_29_), .ZN(n11833) );
  NAND2_X1 U10877 ( .A1(n8480), .A2(n11833), .ZN(n8481) );
  INV_X1 U10878 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n12316) );
  INV_X1 U10879 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n11636) );
  MUX2_X1 U10880 ( .A(n12316), .B(n11636), .S(n9473), .Z(n8503) );
  XNOR2_X1 U10881 ( .A(n8503), .B(SI_30_), .ZN(n8502) );
  NAND2_X1 U10882 ( .A1(n12315), .A2(n7846), .ZN(n8484) );
  OR2_X1 U10883 ( .A1(n8509), .A2(n11636), .ZN(n8483) );
  INV_X1 U10884 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n13451) );
  NAND2_X1 U10885 ( .A1(n8485), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n8487) );
  NAND2_X1 U10886 ( .A1(n7808), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n8486) );
  OAI211_X1 U10887 ( .C1(n8488), .C2(n13451), .A(n8487), .B(n8486), .ZN(n13234) );
  OAI211_X1 U10888 ( .C1(n8489), .C2(n8551), .A(n6527), .B(n9289), .ZN(n8490)
         );
  AOI21_X1 U10889 ( .B1(n13234), .B2(n6534), .A(n8490), .ZN(n8492) );
  NOR2_X1 U10890 ( .A1(n8492), .A2(n8491), .ZN(n8493) );
  AOI21_X1 U10891 ( .B1(n13232), .B2(n8517), .A(n8493), .ZN(n8539) );
  NAND2_X1 U10892 ( .A1(n13232), .A2(n6534), .ZN(n8495) );
  NAND2_X1 U10893 ( .A1(n13139), .A2(n8310), .ZN(n8494) );
  NAND2_X1 U10894 ( .A1(n8495), .A2(n8494), .ZN(n8538) );
  NAND2_X1 U10895 ( .A1(n8539), .A2(n8538), .ZN(n8541) );
  OAI21_X1 U10896 ( .B1(n8527), .B2(n8526), .A(n8541), .ZN(n8499) );
  AOI22_X1 U10897 ( .A1(n13474), .A2(n6534), .B1(n8517), .B2(n13294), .ZN(
        n8496) );
  INV_X1 U10898 ( .A(n8502), .ZN(n8504) );
  INV_X1 U10899 ( .A(SI_30_), .ZN(n13010) );
  MUX2_X1 U10900 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n9473), .Z(n8506) );
  XNOR2_X1 U10901 ( .A(n8506), .B(SI_31_), .ZN(n8507) );
  XNOR2_X2 U10902 ( .A(n8508), .B(n8507), .ZN(n13575) );
  NAND2_X1 U10903 ( .A1(n13575), .A2(n7846), .ZN(n8511) );
  INV_X1 U10904 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n13577) );
  OR2_X1 U10905 ( .A1(n8509), .A2(n13577), .ZN(n8510) );
  NAND2_X2 U10906 ( .A1(n8511), .A2(n8510), .ZN(n13235) );
  INV_X1 U10907 ( .A(n13234), .ZN(n8512) );
  NAND2_X1 U10908 ( .A1(n13235), .A2(n8512), .ZN(n8534) );
  OR2_X1 U10909 ( .A1(n13235), .A2(n8512), .ZN(n8513) );
  NAND2_X1 U10910 ( .A1(n13457), .A2(n6534), .ZN(n8515) );
  NAND2_X1 U10911 ( .A1(n13140), .A2(n8310), .ZN(n8514) );
  NAND2_X1 U10912 ( .A1(n8515), .A2(n8514), .ZN(n8536) );
  INV_X1 U10913 ( .A(n8536), .ZN(n8522) );
  AND2_X1 U10914 ( .A1(n13140), .A2(n6534), .ZN(n8516) );
  AOI21_X1 U10915 ( .B1(n13457), .B2(n8517), .A(n8516), .ZN(n8537) );
  INV_X1 U10916 ( .A(n8537), .ZN(n8521) );
  AND2_X1 U10917 ( .A1(n13065), .A2(n8517), .ZN(n8518) );
  AOI21_X1 U10918 ( .B1(n13464), .B2(n6534), .A(n8518), .ZN(n8525) );
  NAND2_X1 U10919 ( .A1(n13464), .A2(n8310), .ZN(n8520) );
  NAND2_X1 U10920 ( .A1(n13065), .A2(n6534), .ZN(n8519) );
  NAND2_X1 U10921 ( .A1(n8520), .A2(n8519), .ZN(n8524) );
  OAI22_X1 U10922 ( .A1(n8522), .A2(n8521), .B1(n8525), .B2(n8524), .ZN(n8523)
         );
  INV_X1 U10923 ( .A(n8546), .ZN(n8548) );
  INV_X1 U10924 ( .A(n8524), .ZN(n8531) );
  INV_X1 U10925 ( .A(n8525), .ZN(n8530) );
  INV_X1 U10926 ( .A(n8526), .ZN(n8529) );
  INV_X1 U10927 ( .A(n8527), .ZN(n8528) );
  OAI22_X1 U10928 ( .A1(n8531), .A2(n8530), .B1(n8529), .B2(n8528), .ZN(n8532)
         );
  NAND2_X1 U10929 ( .A1(n8541), .A2(n8532), .ZN(n8545) );
  NAND2_X1 U10930 ( .A1(n13234), .A2(n8348), .ZN(n8533) );
  OAI22_X1 U10931 ( .A1(n8534), .A2(n8310), .B1(n13235), .B2(n8533), .ZN(n8535) );
  INV_X1 U10932 ( .A(n8535), .ZN(n8544) );
  OAI22_X1 U10933 ( .A1(n8539), .A2(n8538), .B1(n8537), .B2(n8536), .ZN(n8540)
         );
  NAND3_X1 U10934 ( .A1(n8542), .A2(n8541), .A3(n8540), .ZN(n8543) );
  OAI211_X1 U10935 ( .C1(n8546), .C2(n8545), .A(n8544), .B(n8543), .ZN(n8547)
         );
  MUX2_X1 U10936 ( .A(n8589), .B(n8549), .S(n8551), .Z(n8550) );
  AOI21_X1 U10937 ( .B1(n11044), .B2(n8551), .A(n14491), .ZN(n8552) );
  AOI21_X1 U10938 ( .B1(n8553), .B2(n11796), .A(n8552), .ZN(n8554) );
  AND2_X1 U10939 ( .A1(n9536), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8584) );
  INV_X1 U10940 ( .A(n8584), .ZN(n11327) );
  OAI211_X1 U10941 ( .C1(n8556), .C2(n7604), .A(n8555), .B(n8584), .ZN(n8592)
         );
  NAND2_X1 U10942 ( .A1(n8556), .A2(n6531), .ZN(n8585) );
  XOR2_X1 U10943 ( .A(n13139), .B(n13232), .Z(n8580) );
  XOR2_X1 U10944 ( .A(n13294), .B(n13474), .Z(n13284) );
  NAND2_X1 U10945 ( .A1(n8558), .A2(n8557), .ZN(n13329) );
  XNOR2_X1 U10946 ( .A(n13516), .B(n13372), .ZN(n13387) );
  XNOR2_X1 U10947 ( .A(n14498), .B(n13400), .ZN(n13423) );
  NAND2_X1 U10948 ( .A1(n10210), .A2(n8559), .ZN(n14882) );
  NOR4_X1 U10949 ( .A1(n10232), .A2(n14882), .A3(n10209), .A4(n6531), .ZN(
        n8561) );
  NAND4_X1 U10950 ( .A1(n10563), .A2(n8561), .A3(n8560), .A4(n10254), .ZN(
        n8562) );
  NOR4_X1 U10951 ( .A1(n10729), .A2(n10201), .A3(n8562), .A4(n10185), .ZN(
        n8565) );
  NAND4_X1 U10952 ( .A1(n8566), .A2(n8565), .A3(n8564), .A4(n8563), .ZN(n8568)
         );
  NOR4_X1 U10953 ( .A1(n8568), .A2(n10765), .A3(n8567), .A4(n10851), .ZN(n8570) );
  NAND4_X1 U10954 ( .A1(n13423), .A2(n8570), .A3(n11340), .A4(n8569), .ZN(
        n8571) );
  NOR4_X1 U10955 ( .A1(n13370), .A2(n13394), .A3(n13387), .A4(n8571), .ZN(
        n8573) );
  NAND4_X1 U10956 ( .A1(n13329), .A2(n8573), .A3(n8572), .A4(n13364), .ZN(
        n8574) );
  NOR4_X1 U10957 ( .A1(n13284), .A2(n13310), .A3(n8575), .A4(n8574), .ZN(n8577) );
  NAND4_X1 U10958 ( .A1(n8578), .A2(n8577), .A3(n8576), .A4(n13264), .ZN(n8579) );
  NOR3_X1 U10959 ( .A1(n8581), .A2(n8580), .A3(n8579), .ZN(n8582) );
  XOR2_X1 U10960 ( .A(n14491), .B(n8582), .Z(n8583) );
  NAND4_X1 U10961 ( .A1(n8585), .A2(n8584), .A3(n8583), .A4(n11044), .ZN(n8591) );
  INV_X1 U10962 ( .A(n9536), .ZN(n8586) );
  AND2_X1 U10963 ( .A1(n8586), .A2(n9163), .ZN(n8587) );
  AND2_X1 U10964 ( .A1(n10191), .A2(n8587), .ZN(n9301) );
  NOR2_X1 U10965 ( .A1(n9541), .A2(P2_U3088), .ZN(n13589) );
  NAND3_X1 U10966 ( .A1(n9301), .A2(n13401), .A3(n13589), .ZN(n8588) );
  OAI211_X1 U10967 ( .C1(n8589), .C2(n11327), .A(n8588), .B(P2_B_REG_SCAN_IN), 
        .ZN(n8590) );
  NAND3_X1 U10968 ( .A1(n8592), .A2(n8591), .A3(n8590), .ZN(P2_U3328) );
  INV_X2 U10969 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  NOR2_X1 U10970 ( .A1(P3_IR_REG_23__SCAN_IN), .A2(P3_IR_REG_25__SCAN_IN), 
        .ZN(n8599) );
  NOR2_X1 U10971 ( .A1(P3_IR_REG_22__SCAN_IN), .A2(P3_IR_REG_21__SCAN_IN), 
        .ZN(n8598) );
  NAND2_X1 U10972 ( .A1(n6542), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n8610) );
  NAND2_X1 U10973 ( .A1(n11899), .A2(P3_REG2_REG_11__SCAN_IN), .ZN(n8609) );
  NAND2_X1 U10974 ( .A1(n8749), .A2(n10275), .ZN(n8751) );
  NOR2_X1 U10975 ( .A1(P3_REG3_REG_9__SCAN_IN), .A2(P3_REG3_REG_8__SCAN_IN), 
        .ZN(n8605) );
  XNOR2_X1 U10976 ( .A(n8831), .B(P3_REG3_REG_11__SCAN_IN), .ZN(n14430) );
  NAND2_X1 U10977 ( .A1(n8697), .A2(n14430), .ZN(n8608) );
  INV_X1 U10978 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n8606) );
  OR2_X1 U10979 ( .A1(n6525), .A2(n8606), .ZN(n8607) );
  NAND4_X1 U10980 ( .A1(n8610), .A2(n8609), .A3(n8608), .A4(n8607), .ZN(n12553) );
  NAND2_X1 U10981 ( .A1(n8698), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n8617) );
  NAND2_X1 U10982 ( .A1(n6542), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n8616) );
  OR2_X1 U10983 ( .A1(n8798), .A2(n8611), .ZN(n8612) );
  NAND2_X1 U10984 ( .A1(n8831), .A2(n8612), .ZN(n12424) );
  NAND2_X1 U10985 ( .A1(n8697), .A2(n12424), .ZN(n8615) );
  INV_X1 U10986 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n8613) );
  OR2_X1 U10987 ( .A1(n6525), .A2(n8613), .ZN(n8614) );
  NAND4_X1 U10988 ( .A1(n8617), .A2(n8616), .A3(n8615), .A4(n8614), .ZN(n14427) );
  INV_X1 U10989 ( .A(n14427), .ZN(n10918) );
  INV_X1 U10990 ( .A(P3_B_REG_SCAN_IN), .ZN(n11837) );
  XNOR2_X1 U10991 ( .A(n8626), .B(n11837), .ZN(n8622) );
  INV_X1 U10992 ( .A(P3_IR_REG_25__SCAN_IN), .ZN(n8620) );
  NOR2_X1 U10993 ( .A1(n6656), .A2(n8847), .ZN(n8623) );
  MUX2_X1 U10994 ( .A(n8847), .B(n8623), .S(P3_IR_REG_26__SCAN_IN), .Z(n8625)
         );
  OR2_X1 U10995 ( .A1(n8626), .A2(n9096), .ZN(n8627) );
  INV_X1 U10996 ( .A(n8628), .ZN(n8629) );
  NAND2_X1 U10997 ( .A1(n8629), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8631) );
  XNOR2_X1 U10998 ( .A(n8631), .B(n8630), .ZN(n10611) );
  NAND2_X1 U10999 ( .A1(n8632), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8633) );
  XNOR2_X2 U11000 ( .A(n8633), .B(P3_IR_REG_19__SCAN_IN), .ZN(n12691) );
  NAND2_X1 U11001 ( .A1(n10611), .A2(n12691), .ZN(n12104) );
  INV_X1 U11002 ( .A(n12104), .ZN(n11287) );
  NAND2_X1 U11003 ( .A1(n8634), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8635) );
  XNOR2_X1 U11004 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .ZN(n8705) );
  NAND2_X1 U11005 ( .A1(n9474), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n8636) );
  XNOR2_X1 U11006 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .ZN(n8714) );
  NAND2_X1 U11007 ( .A1(n8716), .A2(n8714), .ZN(n8639) );
  NAND2_X1 U11008 ( .A1(n9493), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n8638) );
  XNOR2_X1 U11009 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .ZN(n8729) );
  NAND2_X1 U11010 ( .A1(n8731), .A2(n8729), .ZN(n8642) );
  NAND2_X1 U11011 ( .A1(n8640), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n8641) );
  NAND2_X1 U11012 ( .A1(n9494), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n8643) );
  NAND2_X1 U11013 ( .A1(n9492), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n8645) );
  NAND2_X1 U11014 ( .A1(n9505), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n8647) );
  NAND2_X1 U11015 ( .A1(n15379), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n8648) );
  XNOR2_X1 U11016 ( .A(n8811), .B(n8810), .ZN(n14371) );
  NAND2_X1 U11017 ( .A1(n8650), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8652) );
  XNOR2_X2 U11018 ( .A(n8652), .B(n8651), .ZN(n9116) );
  NAND2_X1 U11019 ( .A1(n14371), .A2(n11913), .ZN(n8661) );
  NAND2_X1 U11020 ( .A1(n8678), .A2(n8679), .ZN(n8745) );
  NAND2_X1 U11021 ( .A1(n8671), .A2(n8656), .ZN(n8777) );
  NAND2_X1 U11022 ( .A1(n8815), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8658) );
  INV_X1 U11023 ( .A(P3_IR_REG_10__SCAN_IN), .ZN(n8657) );
  XNOR2_X1 U11024 ( .A(n8658), .B(n8657), .ZN(n14374) );
  INV_X1 U11025 ( .A(n14374), .ZN(n15014) );
  OAI22_X1 U11026 ( .A1(n9031), .A2(SI_10_), .B1(n15014), .B2(n9724), .ZN(
        n8659) );
  INV_X1 U11027 ( .A(n8659), .ZN(n8660) );
  NAND2_X1 U11028 ( .A1(n8661), .A2(n8660), .ZN(n10946) );
  INV_X1 U11029 ( .A(n10946), .ZN(n12423) );
  XNOR2_X1 U11030 ( .A(n8709), .B(n12423), .ZN(n8808) );
  INV_X1 U11031 ( .A(n8808), .ZN(n8809) );
  NAND2_X1 U11032 ( .A1(n8698), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n8667) );
  NAND2_X1 U11033 ( .A1(n8751), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n8662) );
  NAND2_X1 U11034 ( .A1(n8759), .A2(n8662), .ZN(n12526) );
  NAND2_X1 U11035 ( .A1(n8697), .A2(n12526), .ZN(n8666) );
  NAND2_X1 U11036 ( .A1(n6542), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n8665) );
  INV_X1 U11037 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n8663) );
  OR2_X1 U11038 ( .A1(n6525), .A2(n8663), .ZN(n8664) );
  NAND4_X1 U11039 ( .A1(n8667), .A2(n8666), .A3(n8665), .A4(n8664), .ZN(n15036) );
  INV_X1 U11040 ( .A(n15036), .ZN(n10585) );
  XNOR2_X1 U11041 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .ZN(n8668) );
  XNOR2_X1 U11042 ( .A(n8669), .B(n8668), .ZN(n14352) );
  NAND2_X1 U11043 ( .A1(n11913), .A2(n14352), .ZN(n8675) );
  INV_X1 U11044 ( .A(SI_6_), .ZN(n8670) );
  OR2_X1 U11045 ( .A1(n9031), .A2(n8670), .ZN(n8674) );
  OR2_X1 U11046 ( .A1(n8671), .A2(n8847), .ZN(n8672) );
  INV_X1 U11047 ( .A(n14986), .ZN(n14354) );
  OR2_X1 U11048 ( .A1(n9724), .A2(n14354), .ZN(n8673) );
  XNOR2_X1 U11049 ( .A(n8709), .B(n15086), .ZN(n8758) );
  XNOR2_X1 U11050 ( .A(n8677), .B(n7323), .ZN(n14355) );
  NAND2_X1 U11051 ( .A1(n8717), .A2(n14355), .ZN(n8682) );
  OR2_X1 U11052 ( .A1(n8678), .A2(n8847), .ZN(n8680) );
  XNOR2_X1 U11053 ( .A(n8680), .B(n8679), .ZN(n14358) );
  INV_X1 U11054 ( .A(n14358), .ZN(n10056) );
  OR2_X1 U11055 ( .A1(n9724), .A2(n10056), .ZN(n8681) );
  OAI211_X1 U11056 ( .C1(n9031), .C2(SI_4_), .A(n8682), .B(n8681), .ZN(n15061)
         );
  XNOR2_X1 U11057 ( .A(n8709), .B(n15061), .ZN(n8742) );
  NAND2_X1 U11058 ( .A1(n8698), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n8687) );
  OR2_X1 U11059 ( .A1(n6687), .A2(n8749), .ZN(n15057) );
  NAND2_X1 U11060 ( .A1(n8697), .A2(n15057), .ZN(n8686) );
  NAND2_X1 U11061 ( .A1(n6542), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n8685) );
  INV_X1 U11062 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n8683) );
  NAND2_X1 U11063 ( .A1(n8697), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n8692) );
  NAND2_X1 U11064 ( .A1(n6541), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n8691) );
  NAND2_X1 U11065 ( .A1(n8698), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n8690) );
  INV_X1 U11066 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n8688) );
  INV_X1 U11067 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n8696) );
  INV_X1 U11068 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n9383) );
  AND2_X1 U11069 ( .A1(n9383), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n15357) );
  NOR2_X1 U11070 ( .A1(n8704), .A2(n15357), .ZN(n8694) );
  OAI21_X1 U11071 ( .B1(n9473), .B2(n8694), .A(n8693), .ZN(n13023) );
  INV_X1 U11072 ( .A(n13023), .ZN(n8695) );
  NAND2_X1 U11073 ( .A1(n8697), .A2(P3_REG3_REG_1__SCAN_IN), .ZN(n8703) );
  NAND2_X1 U11074 ( .A1(n8698), .A2(P3_REG2_REG_1__SCAN_IN), .ZN(n8702) );
  NAND2_X1 U11075 ( .A1(n6541), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n8701) );
  INV_X1 U11076 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n8699) );
  XNOR2_X1 U11077 ( .A(n8705), .B(n8704), .ZN(n9464) );
  NAND2_X1 U11078 ( .A1(n8717), .A2(n9464), .ZN(n8708) );
  OR2_X1 U11079 ( .A1(n8852), .A2(n9466), .ZN(n8707) );
  OR2_X1 U11080 ( .A1(n9724), .A2(n6532), .ZN(n8706) );
  NAND3_X1 U11081 ( .A1(n8709), .A2(n7481), .A3(n10041), .ZN(n8711) );
  INV_X1 U11082 ( .A(n9947), .ZN(n9949) );
  INV_X1 U11083 ( .A(n8712), .ZN(n8713) );
  INV_X1 U11084 ( .A(n8714), .ZN(n8715) );
  XNOR2_X1 U11085 ( .A(n8716), .B(n8715), .ZN(n14359) );
  NAND2_X1 U11086 ( .A1(n8717), .A2(n14359), .ZN(n8722) );
  OR2_X1 U11087 ( .A1(n8852), .A2(SI_2_), .ZN(n8721) );
  INV_X1 U11088 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n8718) );
  OR2_X1 U11089 ( .A1(n9724), .A2(n9814), .ZN(n8720) );
  XNOR2_X1 U11090 ( .A(n8709), .B(n10096), .ZN(n8728) );
  NAND2_X1 U11091 ( .A1(n8698), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n8727) );
  NAND2_X1 U11092 ( .A1(n8697), .A2(P3_REG3_REG_2__SCAN_IN), .ZN(n8726) );
  NAND2_X1 U11093 ( .A1(n6541), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n8725) );
  INV_X1 U11094 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n8723) );
  XNOR2_X1 U11095 ( .A(n8728), .B(n12557), .ZN(n9995) );
  INV_X1 U11096 ( .A(n8729), .ZN(n8730) );
  XNOR2_X1 U11097 ( .A(n8731), .B(n8730), .ZN(n9463) );
  NAND2_X1 U11098 ( .A1(n8717), .A2(n9463), .ZN(n8734) );
  NAND2_X1 U11099 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(n6592), .ZN(n8732) );
  OR2_X1 U11100 ( .A1(n9724), .A2(n14952), .ZN(n8733) );
  OAI211_X1 U11101 ( .C1(n9031), .C2(SI_3_), .A(n8734), .B(n8733), .ZN(n15075)
         );
  INV_X1 U11102 ( .A(n15075), .ZN(n12433) );
  XNOR2_X1 U11103 ( .A(n8709), .B(n12433), .ZN(n8740) );
  INV_X1 U11104 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n12434) );
  NAND2_X1 U11105 ( .A1(n8697), .A2(n12434), .ZN(n8739) );
  NAND2_X1 U11106 ( .A1(n8698), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n8738) );
  NAND2_X1 U11107 ( .A1(n6542), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n8737) );
  INV_X1 U11108 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n8735) );
  XNOR2_X1 U11109 ( .A(n8740), .B(n15054), .ZN(n12431) );
  XNOR2_X1 U11110 ( .A(n8742), .B(n15037), .ZN(n10108) );
  NAND2_X1 U11111 ( .A1(n10109), .A2(n10108), .ZN(n10107) );
  XNOR2_X1 U11112 ( .A(n8744), .B(n7326), .ZN(n9470) );
  NAND2_X1 U11113 ( .A1(n11913), .A2(n9470), .ZN(n8748) );
  NAND2_X1 U11114 ( .A1(n8745), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8746) );
  OR2_X1 U11115 ( .A1(n9724), .A2(n14966), .ZN(n8747) );
  OAI211_X1 U11116 ( .C1(n9031), .C2(SI_5_), .A(n8748), .B(n8747), .ZN(n15046)
         );
  XNOR2_X1 U11117 ( .A(n8709), .B(n15046), .ZN(n8757) );
  NAND2_X1 U11118 ( .A1(n6542), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n8756) );
  NAND2_X1 U11119 ( .A1(n8698), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n8755) );
  OR2_X1 U11120 ( .A1(n8749), .A2(n10275), .ZN(n8750) );
  NAND2_X1 U11121 ( .A1(n8751), .A2(n8750), .ZN(n15047) );
  NAND2_X1 U11122 ( .A1(n8697), .A2(n15047), .ZN(n8754) );
  INV_X1 U11123 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n8752) );
  OR2_X1 U11124 ( .A1(n6525), .A2(n8752), .ZN(n8753) );
  NAND4_X1 U11125 ( .A1(n8756), .A2(n8755), .A3(n8754), .A4(n8753), .ZN(n15053) );
  XNOR2_X1 U11126 ( .A(n8757), .B(n15053), .ZN(n10273) );
  INV_X1 U11127 ( .A(n15053), .ZN(n10111) );
  XNOR2_X1 U11128 ( .A(n8758), .B(n15036), .ZN(n12520) );
  NAND2_X1 U11129 ( .A1(n6542), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n8765) );
  NAND2_X1 U11130 ( .A1(n8698), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n8764) );
  AND2_X1 U11131 ( .A1(n8759), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n8760) );
  OR2_X1 U11132 ( .A1(n8760), .A2(n8796), .ZN(n10470) );
  NAND2_X1 U11133 ( .A1(n8697), .A2(n10470), .ZN(n8763) );
  INV_X1 U11134 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n8761) );
  OR2_X1 U11135 ( .A1(n6525), .A2(n8761), .ZN(n8762) );
  NAND4_X1 U11136 ( .A1(n8765), .A2(n8764), .A3(n8763), .A4(n8762), .ZN(n12556) );
  XNOR2_X1 U11137 ( .A(n8767), .B(n8766), .ZN(n9467) );
  NAND2_X1 U11138 ( .A1(n11913), .A2(n9467), .ZN(n8770) );
  NAND2_X1 U11139 ( .A1(n8777), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8768) );
  XNOR2_X1 U11140 ( .A(n8768), .B(P3_IR_REG_7__SCAN_IN), .ZN(n15004) );
  OR2_X1 U11141 ( .A1(n9724), .A2(n15004), .ZN(n8769) );
  OAI211_X1 U11142 ( .C1(n9031), .C2(SI_7_), .A(n8770), .B(n8769), .ZN(n10584)
         );
  INV_X1 U11143 ( .A(n12005), .ZN(n10624) );
  AND2_X1 U11144 ( .A1(n12556), .A2(n10584), .ZN(n12006) );
  INV_X1 U11145 ( .A(n12006), .ZN(n8771) );
  XNOR2_X1 U11146 ( .A(n12003), .B(n8989), .ZN(n10582) );
  NAND2_X1 U11147 ( .A1(n10583), .A2(n10582), .ZN(n10581) );
  INV_X1 U11148 ( .A(n10582), .ZN(n8772) );
  INV_X1 U11149 ( .A(n12556), .ZN(n10758) );
  NAND2_X1 U11150 ( .A1(n8772), .A2(n12556), .ZN(n8773) );
  NAND2_X1 U11151 ( .A1(n10581), .A2(n8773), .ZN(n10755) );
  INV_X1 U11152 ( .A(n8774), .ZN(n8775) );
  XNOR2_X1 U11153 ( .A(n8776), .B(n8775), .ZN(n14365) );
  NAND2_X1 U11154 ( .A1(n11913), .A2(n14365), .ZN(n8781) );
  INV_X1 U11155 ( .A(SI_8_), .ZN(n14363) );
  OR2_X1 U11156 ( .A1(n9031), .A2(n14363), .ZN(n8780) );
  OAI21_X1 U11157 ( .B1(n8777), .B2(P3_IR_REG_7__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8778) );
  XNOR2_X1 U11158 ( .A(n8778), .B(P3_IR_REG_8__SCAN_IN), .ZN(n10651) );
  INV_X1 U11159 ( .A(n10651), .ZN(n14367) );
  OR2_X1 U11160 ( .A1(n9724), .A2(n14367), .ZN(n8779) );
  XNOR2_X1 U11161 ( .A(n8709), .B(n10756), .ZN(n8787) );
  NAND2_X1 U11162 ( .A1(n8698), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n8786) );
  NAND2_X1 U11163 ( .A1(n6542), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n8785) );
  INV_X1 U11164 ( .A(P3_REG3_REG_8__SCAN_IN), .ZN(n10086) );
  XNOR2_X1 U11165 ( .A(n8796), .B(n10086), .ZN(n10621) );
  NAND2_X1 U11166 ( .A1(n8697), .A2(n10621), .ZN(n8784) );
  INV_X1 U11167 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n8782) );
  OR2_X1 U11168 ( .A1(n6525), .A2(n8782), .ZN(n8783) );
  NAND4_X1 U11169 ( .A1(n8786), .A2(n8785), .A3(n8784), .A4(n8783), .ZN(n12555) );
  XNOR2_X1 U11170 ( .A(n8787), .B(n12555), .ZN(n10754) );
  NAND2_X1 U11171 ( .A1(n10755), .A2(n10754), .ZN(n10753) );
  INV_X1 U11172 ( .A(n12555), .ZN(n10919) );
  OR2_X1 U11173 ( .A1(n8787), .A2(n10919), .ZN(n8788) );
  NAND2_X1 U11174 ( .A1(n10753), .A2(n8788), .ZN(n10916) );
  INV_X1 U11175 ( .A(n10916), .ZN(n8805) );
  XNOR2_X1 U11176 ( .A(n8790), .B(n8789), .ZN(n9471) );
  NAND2_X1 U11177 ( .A1(n9471), .A2(n11913), .ZN(n8795) );
  NAND2_X1 U11178 ( .A1(n8791), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8792) );
  MUX2_X1 U11179 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8792), .S(
        P3_IR_REG_9__SCAN_IN), .Z(n8793) );
  AND2_X1 U11180 ( .A1(n8793), .A2(n8815), .ZN(n10648) );
  OR2_X1 U11181 ( .A1(n9724), .A2(n10648), .ZN(n8794) );
  OAI211_X1 U11182 ( .C1(SI_9_), .C2(n9031), .A(n8795), .B(n8794), .ZN(n15100)
         );
  INV_X1 U11183 ( .A(n15100), .ZN(n10939) );
  XNOR2_X1 U11184 ( .A(n8709), .B(n10939), .ZN(n8806) );
  NAND2_X1 U11185 ( .A1(n6542), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n8803) );
  NAND2_X1 U11186 ( .A1(n8698), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n8802) );
  INV_X1 U11187 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n10649) );
  AOI21_X1 U11188 ( .B1(n8796), .B2(n10086), .A(n10649), .ZN(n8797) );
  OR2_X1 U11189 ( .A1(n8798), .A2(n8797), .ZN(n10922) );
  NAND2_X1 U11190 ( .A1(n8697), .A2(n10922), .ZN(n8801) );
  INV_X1 U11191 ( .A(P3_REG0_REG_9__SCAN_IN), .ZN(n8799) );
  OR2_X1 U11192 ( .A1(n6525), .A2(n8799), .ZN(n8800) );
  NAND4_X1 U11193 ( .A1(n8803), .A2(n8802), .A3(n8801), .A4(n8800), .ZN(n12554) );
  XNOR2_X1 U11194 ( .A(n8806), .B(n12554), .ZN(n10917) );
  INV_X1 U11195 ( .A(n10917), .ZN(n8804) );
  OR2_X1 U11196 ( .A1(n8806), .A2(n12554), .ZN(n8807) );
  XNOR2_X1 U11197 ( .A(n8808), .B(n14427), .ZN(n12418) );
  NAND2_X1 U11198 ( .A1(n9623), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n8812) );
  XNOR2_X1 U11199 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .ZN(n8814) );
  XNOR2_X1 U11200 ( .A(n8822), .B(n8814), .ZN(n9482) );
  NAND2_X1 U11201 ( .A1(n9482), .A2(n11913), .ZN(n8819) );
  OR2_X1 U11202 ( .A1(n8826), .A2(n8847), .ZN(n8816) );
  XNOR2_X1 U11203 ( .A(n8816), .B(P3_IR_REG_11__SCAN_IN), .ZN(n11096) );
  OAI22_X1 U11204 ( .A1(n9031), .A2(SI_11_), .B1(n11096), .B2(n9724), .ZN(
        n8817) );
  INV_X1 U11205 ( .A(n8817), .ZN(n8818) );
  NAND2_X1 U11206 ( .A1(n8819), .A2(n8818), .ZN(n14434) );
  INV_X1 U11207 ( .A(n14434), .ZN(n11181) );
  XNOR2_X1 U11208 ( .A(n11181), .B(n8709), .ZN(n8820) );
  AND2_X1 U11209 ( .A1(n8821), .A2(n8820), .ZN(n11296) );
  NAND2_X1 U11210 ( .A1(n9700), .A2(P2_DATAO_REG_11__SCAN_IN), .ZN(n8823) );
  XNOR2_X1 U11211 ( .A(n9589), .B(P1_DATAO_REG_12__SCAN_IN), .ZN(n8842) );
  INV_X1 U11212 ( .A(n8842), .ZN(n8824) );
  XNOR2_X1 U11213 ( .A(n8841), .B(n8824), .ZN(n9507) );
  NAND2_X1 U11214 ( .A1(n9507), .A2(n11913), .ZN(n8830) );
  OR2_X1 U11215 ( .A1(n8845), .A2(n8847), .ZN(n8827) );
  INV_X1 U11216 ( .A(P3_IR_REG_12__SCAN_IN), .ZN(n8844) );
  XNOR2_X1 U11217 ( .A(n8827), .B(n8844), .ZN(n12564) );
  OAI22_X1 U11218 ( .A1(n9031), .A2(n15403), .B1(n12564), .B2(n9724), .ZN(
        n8828) );
  INV_X1 U11219 ( .A(n8828), .ZN(n8829) );
  NAND2_X1 U11220 ( .A1(n8830), .A2(n8829), .ZN(n11279) );
  XNOR2_X1 U11221 ( .A(n11279), .B(n8709), .ZN(n8838) );
  NAND2_X1 U11222 ( .A1(n6542), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n8837) );
  NAND2_X1 U11223 ( .A1(n11899), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n8836) );
  OAI21_X1 U11224 ( .B1(n8831), .B2(P3_REG3_REG_11__SCAN_IN), .A(
        P3_REG3_REG_12__SCAN_IN), .ZN(n8832) );
  NAND2_X1 U11225 ( .A1(n8832), .A2(n8855), .ZN(n11395) );
  NAND2_X1 U11226 ( .A1(n8697), .A2(n11395), .ZN(n8835) );
  INV_X1 U11227 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n8833) );
  OR2_X1 U11228 ( .A1(n6525), .A2(n8833), .ZN(n8834) );
  NAND4_X1 U11229 ( .A1(n8837), .A2(n8836), .A3(n8835), .A4(n8834), .ZN(n14428) );
  XNOR2_X1 U11230 ( .A(n8838), .B(n11419), .ZN(n11389) );
  INV_X1 U11231 ( .A(n8838), .ZN(n8839) );
  NAND2_X1 U11232 ( .A1(n8839), .A2(n11419), .ZN(n8840) );
  XNOR2_X1 U11233 ( .A(n8863), .B(n8843), .ZN(n8862) );
  XNOR2_X1 U11234 ( .A(n8862), .B(P1_DATAO_REG_13__SCAN_IN), .ZN(n9526) );
  NAND2_X1 U11235 ( .A1(n9526), .A2(n11913), .ZN(n8854) );
  NOR2_X1 U11236 ( .A1(n8850), .A2(n8847), .ZN(n8846) );
  MUX2_X1 U11237 ( .A(n8847), .B(n8846), .S(P3_IR_REG_13__SCAN_IN), .Z(n8848)
         );
  INV_X1 U11238 ( .A(n8848), .ZN(n8851) );
  INV_X1 U11239 ( .A(P3_IR_REG_13__SCAN_IN), .ZN(n8849) );
  NAND2_X1 U11240 ( .A1(n8850), .A2(n8849), .ZN(n8885) );
  NAND2_X1 U11241 ( .A1(n8851), .A2(n8885), .ZN(n12582) );
  INV_X1 U11242 ( .A(n9724), .ZN(n8922) );
  INV_X1 U11243 ( .A(n9031), .ZN(n8900) );
  AOI22_X1 U11244 ( .A1(n12582), .A2(n8922), .B1(n8900), .B2(n9527), .ZN(n8853) );
  XOR2_X1 U11245 ( .A(n8709), .B(n11420), .Z(n11415) );
  NAND2_X1 U11246 ( .A1(n8698), .A2(P3_REG2_REG_13__SCAN_IN), .ZN(n8861) );
  NAND2_X1 U11247 ( .A1(n6542), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n8860) );
  INV_X1 U11248 ( .A(n8873), .ZN(n8857) );
  NAND2_X1 U11249 ( .A1(n8855), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n8856) );
  NAND2_X1 U11250 ( .A1(n8857), .A2(n8856), .ZN(n11423) );
  NAND2_X1 U11251 ( .A1(n8697), .A2(n11423), .ZN(n8859) );
  INV_X1 U11252 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n11291) );
  OR2_X1 U11253 ( .A1(n6525), .A2(n11291), .ZN(n8858) );
  NAND4_X1 U11254 ( .A1(n8861), .A2(n8860), .A3(n8859), .A4(n8858), .ZN(n12552) );
  NAND2_X1 U11255 ( .A1(n8862), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n8865) );
  XNOR2_X1 U11256 ( .A(n9848), .B(P1_DATAO_REG_14__SCAN_IN), .ZN(n8866) );
  XNOR2_X1 U11257 ( .A(n8883), .B(n8866), .ZN(n14377) );
  NAND2_X1 U11258 ( .A1(n14377), .A2(n11913), .ZN(n8872) );
  NAND2_X1 U11259 ( .A1(n8885), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8868) );
  INV_X1 U11260 ( .A(P3_IR_REG_14__SCAN_IN), .ZN(n8867) );
  XNOR2_X1 U11261 ( .A(n8868), .B(n8867), .ZN(n14379) );
  OAI22_X1 U11262 ( .A1(n14379), .A2(n9724), .B1(n8869), .B2(n9031), .ZN(n8870) );
  INV_X1 U11263 ( .A(n8870), .ZN(n8871) );
  XNOR2_X1 U11264 ( .A(n12408), .B(n8989), .ZN(n8879) );
  NAND2_X1 U11265 ( .A1(n11899), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n8878) );
  OR2_X1 U11266 ( .A1(n8873), .A2(n12403), .ZN(n8874) );
  NAND2_X1 U11267 ( .A1(n8889), .A2(n8874), .ZN(n12402) );
  NAND2_X1 U11268 ( .A1(n8697), .A2(n12402), .ZN(n8877) );
  NAND2_X1 U11269 ( .A1(n6542), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n8876) );
  INV_X1 U11270 ( .A(P3_REG0_REG_14__SCAN_IN), .ZN(n15160) );
  OR2_X1 U11271 ( .A1(n6525), .A2(n15160), .ZN(n8875) );
  NAND4_X1 U11272 ( .A1(n8878), .A2(n8877), .A3(n8876), .A4(n8875), .ZN(n12551) );
  NAND2_X1 U11273 ( .A1(n8879), .A2(n12538), .ZN(n8881) );
  OAI21_X1 U11274 ( .B1(n8879), .B2(n12538), .A(n8881), .ZN(n12401) );
  INV_X1 U11275 ( .A(n12401), .ZN(n8880) );
  NAND2_X1 U11276 ( .A1(n9848), .A2(P1_DATAO_REG_14__SCAN_IN), .ZN(n8884) );
  XNOR2_X1 U11277 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .ZN(n8895) );
  XNOR2_X1 U11278 ( .A(n8896), .B(n7334), .ZN(n9703) );
  NAND2_X1 U11279 ( .A1(n9703), .A2(n11913), .ZN(n8888) );
  NAND2_X1 U11280 ( .A1(n8899), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8886) );
  XNOR2_X1 U11281 ( .A(n8886), .B(P3_IR_REG_15__SCAN_IN), .ZN(n12626) );
  AOI22_X1 U11282 ( .A1(n12626), .A2(n8922), .B1(SI_15_), .B2(n8900), .ZN(
        n8887) );
  XNOR2_X1 U11283 ( .A(n12922), .B(n8709), .ZN(n8909) );
  NAND2_X1 U11284 ( .A1(n11899), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n8894) );
  NAND2_X1 U11285 ( .A1(n6542), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n8893) );
  NAND2_X1 U11286 ( .A1(n8889), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n8890) );
  NAND2_X1 U11287 ( .A1(n8903), .A2(n8890), .ZN(n12541) );
  NAND2_X1 U11288 ( .A1(n8697), .A2(n12541), .ZN(n8892) );
  INV_X1 U11289 ( .A(P3_REG0_REG_15__SCAN_IN), .ZN(n12997) );
  OR2_X1 U11290 ( .A1(n6525), .A2(n12997), .ZN(n8891) );
  NAND4_X1 U11291 ( .A1(n8894), .A2(n8893), .A3(n8892), .A4(n8891), .ZN(n12550) );
  XNOR2_X1 U11292 ( .A(n8909), .B(n12863), .ZN(n12532) );
  XNOR2_X1 U11293 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(P2_DATAO_REG_16__SCAN_IN), 
        .ZN(n8912) );
  INV_X1 U11294 ( .A(n8912), .ZN(n8898) );
  XNOR2_X1 U11295 ( .A(n8911), .B(n8898), .ZN(n14382) );
  NAND2_X1 U11296 ( .A1(n14382), .A2(n11913), .ZN(n8902) );
  OAI21_X1 U11297 ( .B1(n8899), .B2(P3_IR_REG_15__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8918) );
  XNOR2_X1 U11298 ( .A(n8918), .B(P3_IR_REG_16__SCAN_IN), .ZN(n12636) );
  AOI22_X1 U11299 ( .A1(n12636), .A2(n8922), .B1(SI_16_), .B2(n8900), .ZN(
        n8901) );
  XNOR2_X1 U11300 ( .A(n12918), .B(n8709), .ZN(n8933) );
  NAND2_X1 U11301 ( .A1(n11899), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n8908) );
  NAND2_X1 U11302 ( .A1(n6542), .A2(P3_REG1_REG_16__SCAN_IN), .ZN(n8907) );
  AND2_X1 U11303 ( .A1(n8903), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n8904) );
  OR2_X1 U11304 ( .A1(n8904), .A2(n8926), .ZN(n12867) );
  NAND2_X1 U11305 ( .A1(n8697), .A2(n12867), .ZN(n8906) );
  INV_X1 U11306 ( .A(P3_REG0_REG_16__SCAN_IN), .ZN(n15276) );
  OR2_X1 U11307 ( .A1(n6525), .A2(n15276), .ZN(n8905) );
  NAND4_X1 U11308 ( .A1(n8908), .A2(n8907), .A3(n8906), .A4(n8905), .ZN(n12851) );
  XNOR2_X1 U11309 ( .A(n8933), .B(n12851), .ZN(n12459) );
  NOR2_X1 U11310 ( .A1(n8909), .A2(n12550), .ZN(n12460) );
  NOR2_X1 U11311 ( .A1(n12459), .A2(n12460), .ZN(n8910) );
  AOI22_X1 U11312 ( .A1(P2_DATAO_REG_17__SCAN_IN), .A2(n10179), .B1(
        P1_DATAO_REG_17__SCAN_IN), .B2(n10178), .ZN(n8915) );
  INV_X1 U11313 ( .A(n8915), .ZN(n8916) );
  XNOR2_X1 U11314 ( .A(n8936), .B(n8916), .ZN(n9926) );
  NAND2_X1 U11315 ( .A1(n9926), .A2(n11913), .ZN(n8924) );
  INV_X1 U11316 ( .A(P3_IR_REG_16__SCAN_IN), .ZN(n8917) );
  NAND2_X1 U11317 ( .A1(n8918), .A2(n8917), .ZN(n8919) );
  NAND2_X1 U11318 ( .A1(n8919), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8920) );
  XNOR2_X1 U11319 ( .A(n8920), .B(P3_IR_REG_17__SCAN_IN), .ZN(n12680) );
  NOR2_X1 U11320 ( .A1(n9031), .A2(n15158), .ZN(n8921) );
  AOI21_X1 U11321 ( .B1(n12680), .B2(n8922), .A(n8921), .ZN(n8923) );
  XNOR2_X1 U11322 ( .A(n12987), .B(n8989), .ZN(n8932) );
  NAND2_X1 U11323 ( .A1(n11899), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n8931) );
  INV_X1 U11324 ( .A(P3_REG3_REG_17__SCAN_IN), .ZN(n8925) );
  NOR2_X1 U11325 ( .A1(n8926), .A2(n8925), .ZN(n8927) );
  OR2_X1 U11326 ( .A1(n8944), .A2(n8927), .ZN(n12855) );
  NAND2_X1 U11327 ( .A1(n8697), .A2(n12855), .ZN(n8930) );
  NAND2_X1 U11328 ( .A1(n6542), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n8929) );
  INV_X1 U11329 ( .A(P3_REG0_REG_17__SCAN_IN), .ZN(n12986) );
  OR2_X1 U11330 ( .A1(n6525), .A2(n12986), .ZN(n8928) );
  NAND4_X1 U11331 ( .A1(n8931), .A2(n8930), .A3(n8929), .A4(n8928), .ZN(n12549) );
  NAND2_X1 U11332 ( .A1(n8932), .A2(n12865), .ZN(n8934) );
  OAI21_X1 U11333 ( .B1(n8932), .B2(n12865), .A(n8934), .ZN(n12471) );
  AND2_X1 U11334 ( .A1(n8933), .A2(n12851), .ZN(n12472) );
  NOR2_X1 U11335 ( .A1(P2_DATAO_REG_17__SCAN_IN), .A2(n10179), .ZN(n8935) );
  INV_X1 U11336 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n10503) );
  AOI22_X1 U11337 ( .A1(P2_DATAO_REG_18__SCAN_IN), .A2(
        P1_DATAO_REG_18__SCAN_IN), .B1(n10503), .B2(n10502), .ZN(n8954) );
  INV_X1 U11338 ( .A(n8954), .ZN(n8937) );
  XNOR2_X1 U11339 ( .A(n8955), .B(n8937), .ZN(n9981) );
  NAND2_X1 U11340 ( .A1(n9981), .A2(n11913), .ZN(n8943) );
  INV_X1 U11341 ( .A(SI_18_), .ZN(n9983) );
  NAND2_X1 U11342 ( .A1(n8938), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8939) );
  MUX2_X1 U11343 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8939), .S(
        P3_IR_REG_18__SCAN_IN), .Z(n8940) );
  NAND2_X1 U11344 ( .A1(n8940), .A2(n8632), .ZN(n12693) );
  OAI22_X1 U11345 ( .A1(n9031), .A2(n9983), .B1(n9724), .B2(n12693), .ZN(n8941) );
  INV_X1 U11346 ( .A(n8941), .ZN(n8942) );
  XNOR2_X1 U11347 ( .A(n12909), .B(n8709), .ZN(n8951) );
  INV_X1 U11348 ( .A(P3_REG3_REG_18__SCAN_IN), .ZN(n12513) );
  OR2_X1 U11349 ( .A1(n8944), .A2(n12513), .ZN(n8945) );
  NAND2_X1 U11350 ( .A1(n8959), .A2(n8945), .ZN(n12843) );
  NAND2_X1 U11351 ( .A1(n12843), .A2(n8697), .ZN(n8950) );
  NAND2_X1 U11352 ( .A1(n6542), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n8949) );
  NAND2_X1 U11353 ( .A1(n11899), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n8948) );
  INV_X1 U11354 ( .A(P3_REG0_REG_18__SCAN_IN), .ZN(n12982) );
  OR2_X1 U11355 ( .A1(n6525), .A2(n12982), .ZN(n8947) );
  XNOR2_X1 U11356 ( .A(n8951), .B(n11804), .ZN(n12511) );
  NAND2_X1 U11357 ( .A1(n12510), .A2(n12511), .ZN(n12509) );
  INV_X1 U11358 ( .A(n8951), .ZN(n8952) );
  NAND2_X1 U11359 ( .A1(n8952), .A2(n11804), .ZN(n8953) );
  INV_X1 U11360 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n10674) );
  AOI22_X1 U11361 ( .A1(P2_DATAO_REG_19__SCAN_IN), .A2(
        P1_DATAO_REG_19__SCAN_IN), .B1(n10674), .B2(n10672), .ZN(n8969) );
  XNOR2_X1 U11362 ( .A(n8970), .B(n8969), .ZN(n10002) );
  NAND2_X1 U11363 ( .A1(n10002), .A2(n11913), .ZN(n8958) );
  OAI22_X1 U11364 ( .A1(n9031), .A2(SI_19_), .B1(n12691), .B2(n9724), .ZN(
        n8956) );
  INV_X1 U11365 ( .A(n8956), .ZN(n8957) );
  XNOR2_X1 U11366 ( .A(n12979), .B(n8709), .ZN(n8966) );
  INV_X1 U11367 ( .A(P3_REG0_REG_19__SCAN_IN), .ZN(n12975) );
  NAND2_X1 U11368 ( .A1(n8959), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n8960) );
  NAND2_X1 U11369 ( .A1(n8974), .A2(n8960), .ZN(n12829) );
  NAND2_X1 U11370 ( .A1(n12829), .A2(n8697), .ZN(n8964) );
  NAND2_X1 U11371 ( .A1(n6542), .A2(P3_REG1_REG_19__SCAN_IN), .ZN(n8962) );
  NAND2_X1 U11372 ( .A1(n11899), .A2(P3_REG2_REG_19__SCAN_IN), .ZN(n8961) );
  AND2_X1 U11373 ( .A1(n8962), .A2(n8961), .ZN(n8963) );
  OAI211_X1 U11374 ( .C1(n6525), .C2(n12975), .A(n8964), .B(n8963), .ZN(n12816) );
  INV_X1 U11375 ( .A(n12816), .ZN(n12838) );
  XNOR2_X1 U11376 ( .A(n8966), .B(n12838), .ZN(n12439) );
  INV_X1 U11377 ( .A(n8966), .ZN(n8967) );
  NAND2_X1 U11378 ( .A1(n8967), .A2(n12816), .ZN(n8968) );
  XNOR2_X1 U11379 ( .A(n8984), .B(P2_DATAO_REG_20__SCAN_IN), .ZN(n10608) );
  NAND2_X1 U11380 ( .A1(n10608), .A2(n11913), .ZN(n8972) );
  OR2_X1 U11381 ( .A1(n9031), .A2(n10609), .ZN(n8971) );
  XNOR2_X1 U11382 ( .A(n11807), .B(n8709), .ZN(n8979) );
  INV_X1 U11383 ( .A(n6542), .ZN(n8978) );
  INV_X1 U11384 ( .A(P3_REG1_REG_20__SCAN_IN), .ZN(n12901) );
  NAND2_X1 U11385 ( .A1(n8974), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n8975) );
  NAND2_X1 U11386 ( .A1(n8990), .A2(n8975), .ZN(n12820) );
  NAND2_X1 U11387 ( .A1(n12820), .A2(n8697), .ZN(n8977) );
  AOI22_X1 U11388 ( .A1(n10144), .A2(P3_REG0_REG_20__SCAN_IN), .B1(n11899), 
        .B2(P3_REG2_REG_20__SCAN_IN), .ZN(n8976) );
  OAI211_X1 U11389 ( .C1(n8978), .C2(n12901), .A(n8977), .B(n8976), .ZN(n12826) );
  XNOR2_X1 U11390 ( .A(n8979), .B(n12826), .ZN(n12492) );
  INV_X1 U11391 ( .A(n8979), .ZN(n8980) );
  NAND2_X1 U11392 ( .A1(n8980), .A2(n12826), .ZN(n8981) );
  NAND2_X1 U11393 ( .A1(n8983), .A2(n11072), .ZN(n8985) );
  AOI22_X1 U11394 ( .A1(P2_DATAO_REG_21__SCAN_IN), .A2(
        P1_DATAO_REG_21__SCAN_IN), .B1(n11045), .B2(n11487), .ZN(n8998) );
  INV_X1 U11395 ( .A(n8998), .ZN(n8986) );
  XNOR2_X1 U11396 ( .A(n8997), .B(n8986), .ZN(n10723) );
  NAND2_X1 U11397 ( .A1(n10723), .A2(n11913), .ZN(n8988) );
  INV_X1 U11398 ( .A(SI_21_), .ZN(n10725) );
  OR2_X1 U11399 ( .A1(n9031), .A2(n10725), .ZN(n8987) );
  XNOR2_X1 U11400 ( .A(n12964), .B(n8989), .ZN(n8995) );
  AND2_X1 U11401 ( .A1(n8990), .A2(P3_REG3_REG_21__SCAN_IN), .ZN(n8991) );
  OR2_X1 U11402 ( .A1(n8991), .A2(n9006), .ZN(n12810) );
  NAND2_X1 U11403 ( .A1(n12810), .A2(n8697), .ZN(n8994) );
  AOI22_X1 U11404 ( .A1(n6542), .A2(P3_REG1_REG_21__SCAN_IN), .B1(n11899), 
        .B2(P3_REG2_REG_21__SCAN_IN), .ZN(n8993) );
  INV_X1 U11405 ( .A(P3_REG0_REG_21__SCAN_IN), .ZN(n12963) );
  OR2_X1 U11406 ( .A1(n6525), .A2(n12963), .ZN(n8992) );
  NAND2_X1 U11407 ( .A1(n8995), .A2(n12504), .ZN(n8996) );
  OAI21_X1 U11408 ( .B1(n8995), .B2(n12504), .A(n8996), .ZN(n12450) );
  AOI22_X1 U11409 ( .A1(P2_DATAO_REG_22__SCAN_IN), .A2(n11798), .B1(
        P1_DATAO_REG_22__SCAN_IN), .B2(n15376), .ZN(n9014) );
  XNOR2_X1 U11410 ( .A(n9015), .B(n9014), .ZN(n10866) );
  NAND2_X1 U11411 ( .A1(n10866), .A2(n11913), .ZN(n9001) );
  OR2_X1 U11412 ( .A1(n9031), .A2(n8999), .ZN(n9000) );
  XOR2_X1 U11413 ( .A(n8709), .B(n12958), .Z(n9002) );
  NAND2_X1 U11414 ( .A1(n9003), .A2(n9002), .ZN(n9013) );
  NAND2_X1 U11415 ( .A1(n9013), .A2(n9004), .ZN(n12501) );
  INV_X1 U11416 ( .A(P3_REG3_REG_22__SCAN_IN), .ZN(n9005) );
  OR2_X1 U11417 ( .A1(n9006), .A2(n9005), .ZN(n9007) );
  NAND2_X1 U11418 ( .A1(n9035), .A2(n9007), .ZN(n12800) );
  NAND2_X1 U11419 ( .A1(n12800), .A2(n8697), .ZN(n9012) );
  INV_X1 U11420 ( .A(P3_REG0_REG_22__SCAN_IN), .ZN(n12957) );
  NAND2_X1 U11421 ( .A1(n6542), .A2(P3_REG1_REG_22__SCAN_IN), .ZN(n9009) );
  NAND2_X1 U11422 ( .A1(n11899), .A2(P3_REG2_REG_22__SCAN_IN), .ZN(n9008) );
  OAI211_X1 U11423 ( .C1(n12957), .C2(n6525), .A(n9009), .B(n9008), .ZN(n9010)
         );
  INV_X1 U11424 ( .A(n9010), .ZN(n9011) );
  INV_X1 U11425 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n11574) );
  AOI22_X1 U11426 ( .A1(P2_DATAO_REG_23__SCAN_IN), .A2(n9028), .B1(
        P1_DATAO_REG_23__SCAN_IN), .B2(n11574), .ZN(n9026) );
  XNOR2_X1 U11427 ( .A(n9026), .B(n9027), .ZN(n11040) );
  NAND2_X1 U11428 ( .A1(n11040), .A2(n11913), .ZN(n9017) );
  OR2_X1 U11429 ( .A1(n9031), .A2(n11042), .ZN(n9016) );
  XNOR2_X1 U11430 ( .A(n12952), .B(n8709), .ZN(n9018) );
  XNOR2_X1 U11431 ( .A(n9035), .B(P3_REG3_REG_23__SCAN_IN), .ZN(n12788) );
  NAND2_X1 U11432 ( .A1(n12788), .A2(n8697), .ZN(n9025) );
  INV_X1 U11433 ( .A(P3_REG0_REG_23__SCAN_IN), .ZN(n9022) );
  NAND2_X1 U11434 ( .A1(n6542), .A2(P3_REG1_REG_23__SCAN_IN), .ZN(n9021) );
  NAND2_X1 U11435 ( .A1(n11899), .A2(P3_REG2_REG_23__SCAN_IN), .ZN(n9020) );
  OAI211_X1 U11436 ( .C1(n9022), .C2(n6525), .A(n9021), .B(n9020), .ZN(n9023)
         );
  INV_X1 U11437 ( .A(n9023), .ZN(n9024) );
  INV_X1 U11438 ( .A(SI_24_), .ZN(n11277) );
  OR2_X1 U11439 ( .A1(n9031), .A2(n11277), .ZN(n9032) );
  XNOR2_X1 U11440 ( .A(n12491), .B(n8709), .ZN(n9042) );
  OAI21_X1 U11441 ( .B1(n9035), .B2(P3_REG3_REG_23__SCAN_IN), .A(
        P3_REG3_REG_24__SCAN_IN), .ZN(n9036) );
  INV_X1 U11442 ( .A(P3_REG3_REG_24__SCAN_IN), .ZN(n15172) );
  INV_X1 U11443 ( .A(P3_REG3_REG_23__SCAN_IN), .ZN(n9033) );
  NAND2_X1 U11444 ( .A1(n15172), .A2(n9033), .ZN(n9034) );
  NAND2_X1 U11445 ( .A1(n9036), .A2(n9054), .ZN(n12776) );
  NAND2_X1 U11446 ( .A1(n12776), .A2(n8697), .ZN(n9041) );
  INV_X1 U11447 ( .A(P3_REG0_REG_24__SCAN_IN), .ZN(n12946) );
  NAND2_X1 U11448 ( .A1(n6542), .A2(P3_REG1_REG_24__SCAN_IN), .ZN(n9038) );
  NAND2_X1 U11449 ( .A1(n11899), .A2(P3_REG2_REG_24__SCAN_IN), .ZN(n9037) );
  OAI211_X1 U11450 ( .C1(n12946), .C2(n6525), .A(n9038), .B(n9037), .ZN(n9039)
         );
  INV_X1 U11451 ( .A(n9039), .ZN(n9040) );
  NAND2_X1 U11452 ( .A1(n9041), .A2(n9040), .ZN(n12784) );
  INV_X1 U11453 ( .A(n12784), .ZN(n11811) );
  NAND2_X1 U11454 ( .A1(n9042), .A2(n11811), .ZN(n9067) );
  INV_X1 U11455 ( .A(n9042), .ZN(n9043) );
  NAND2_X1 U11456 ( .A1(n9043), .A2(n12784), .ZN(n9044) );
  AND2_X1 U11457 ( .A1(n9067), .A2(n9044), .ZN(n12480) );
  INV_X1 U11458 ( .A(n9067), .ZN(n9065) );
  INV_X1 U11459 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n11483) );
  AOI22_X1 U11460 ( .A1(P2_DATAO_REG_25__SCAN_IN), .A2(
        P1_DATAO_REG_25__SCAN_IN), .B1(n11427), .B2(n15212), .ZN(n9048) );
  INV_X1 U11461 ( .A(n9048), .ZN(n9049) );
  XNOR2_X1 U11462 ( .A(n9134), .B(n9049), .ZN(n11351) );
  NAND2_X1 U11463 ( .A1(n11351), .A2(n11913), .ZN(n9051) );
  OR2_X1 U11464 ( .A1(n9031), .A2(n11353), .ZN(n9050) );
  XNOR2_X1 U11465 ( .A(n12886), .B(n8989), .ZN(n9062) );
  INV_X1 U11466 ( .A(P3_REG3_REG_25__SCAN_IN), .ZN(n9052) );
  NAND2_X1 U11467 ( .A1(n9054), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n9055) );
  NAND2_X1 U11468 ( .A1(n9117), .A2(n9055), .ZN(n12764) );
  NAND2_X1 U11469 ( .A1(n12764), .A2(n8697), .ZN(n9061) );
  INV_X1 U11470 ( .A(P3_REG0_REG_25__SCAN_IN), .ZN(n9058) );
  NAND2_X1 U11471 ( .A1(n6542), .A2(P3_REG1_REG_25__SCAN_IN), .ZN(n9057) );
  NAND2_X1 U11472 ( .A1(n11899), .A2(P3_REG2_REG_25__SCAN_IN), .ZN(n9056) );
  OAI211_X1 U11473 ( .C1(n9058), .C2(n6525), .A(n9057), .B(n9056), .ZN(n9059)
         );
  INV_X1 U11474 ( .A(n9059), .ZN(n9060) );
  NAND2_X1 U11475 ( .A1(n9062), .A2(n15345), .ZN(n9140) );
  INV_X1 U11476 ( .A(n9062), .ZN(n9063) );
  NAND2_X1 U11477 ( .A1(n9063), .A2(n12773), .ZN(n9064) );
  NOR3_X1 U11478 ( .A1(n12482), .A2(n9065), .A3(n9066), .ZN(n9104) );
  INV_X1 U11479 ( .A(n9066), .ZN(n9068) );
  NAND2_X1 U11480 ( .A1(n9142), .A2(n9141), .ZN(n9103) );
  OR2_X1 U11481 ( .A1(n9070), .A2(P3_D_REG_1__SCAN_IN), .ZN(n9072) );
  INV_X1 U11482 ( .A(n9096), .ZN(n13020) );
  NAND2_X1 U11483 ( .A1(n11352), .A2(n13020), .ZN(n9071) );
  NAND2_X1 U11484 ( .A1(n9069), .A2(n13001), .ZN(n9863) );
  INV_X1 U11485 ( .A(n9863), .ZN(n9083) );
  NOR4_X1 U11486 ( .A1(P3_D_REG_19__SCAN_IN), .A2(P3_D_REG_12__SCAN_IN), .A3(
        P3_D_REG_10__SCAN_IN), .A4(P3_D_REG_26__SCAN_IN), .ZN(n15363) );
  NOR2_X1 U11487 ( .A1(P3_D_REG_8__SCAN_IN), .A2(P3_D_REG_7__SCAN_IN), .ZN(
        n9075) );
  NOR4_X1 U11488 ( .A1(P3_D_REG_20__SCAN_IN), .A2(P3_D_REG_22__SCAN_IN), .A3(
        P3_D_REG_25__SCAN_IN), .A4(P3_D_REG_18__SCAN_IN), .ZN(n9074) );
  NOR4_X1 U11489 ( .A1(P3_D_REG_14__SCAN_IN), .A2(P3_D_REG_21__SCAN_IN), .A3(
        P3_D_REG_2__SCAN_IN), .A4(P3_D_REG_17__SCAN_IN), .ZN(n9073) );
  NAND4_X1 U11490 ( .A1(n15363), .A2(n9075), .A3(n9074), .A4(n9073), .ZN(n9081) );
  NOR4_X1 U11491 ( .A1(P3_D_REG_31__SCAN_IN), .A2(P3_D_REG_11__SCAN_IN), .A3(
        P3_D_REG_16__SCAN_IN), .A4(P3_D_REG_15__SCAN_IN), .ZN(n9079) );
  NOR4_X1 U11492 ( .A1(P3_D_REG_27__SCAN_IN), .A2(P3_D_REG_24__SCAN_IN), .A3(
        P3_D_REG_29__SCAN_IN), .A4(P3_D_REG_9__SCAN_IN), .ZN(n9078) );
  NOR4_X1 U11493 ( .A1(P3_D_REG_23__SCAN_IN), .A2(P3_D_REG_4__SCAN_IN), .A3(
        P3_D_REG_3__SCAN_IN), .A4(P3_D_REG_5__SCAN_IN), .ZN(n9077) );
  NOR4_X1 U11494 ( .A1(P3_D_REG_30__SCAN_IN), .A2(P3_D_REG_13__SCAN_IN), .A3(
        P3_D_REG_6__SCAN_IN), .A4(P3_D_REG_28__SCAN_IN), .ZN(n9076) );
  NAND4_X1 U11495 ( .A1(n9079), .A2(n9078), .A3(n9077), .A4(n9076), .ZN(n9080)
         );
  NOR2_X1 U11496 ( .A1(n9081), .A2(n9080), .ZN(n9082) );
  NAND2_X1 U11497 ( .A1(n9083), .A2(n9860), .ZN(n9933) );
  INV_X1 U11498 ( .A(n9084), .ZN(n9085) );
  NAND2_X1 U11499 ( .A1(n9085), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9086) );
  MUX2_X1 U11500 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9086), .S(
        P3_IR_REG_22__SCAN_IN), .Z(n9087) );
  OAI21_X1 U11501 ( .B1(n11288), .B2(n9937), .A(n12691), .ZN(n9088) );
  NAND2_X1 U11502 ( .A1(n9088), .A2(n6523), .ZN(n9090) );
  OAI21_X1 U11503 ( .B1(n11968), .B2(n9937), .A(n11288), .ZN(n9089) );
  NAND2_X1 U11504 ( .A1(n9090), .A2(n9089), .ZN(n10040) );
  NAND2_X1 U11505 ( .A1(n10040), .A2(n15099), .ZN(n9095) );
  INV_X1 U11506 ( .A(n9069), .ZN(n9091) );
  NAND2_X1 U11507 ( .A1(n9091), .A2(n9939), .ZN(n9861) );
  INV_X1 U11508 ( .A(n9860), .ZN(n9092) );
  NAND2_X1 U11509 ( .A1(n12114), .A2(n12691), .ZN(n10045) );
  INV_X1 U11510 ( .A(n10045), .ZN(n9094) );
  NAND2_X1 U11511 ( .A1(n6523), .A2(n9937), .ZN(n12107) );
  INV_X1 U11512 ( .A(n12107), .ZN(n9093) );
  NAND2_X1 U11513 ( .A1(n9094), .A2(n9093), .ZN(n9929) );
  OAI22_X1 U11514 ( .A1(n9933), .A2(n9095), .B1(n9930), .B2(n9929), .ZN(n9102)
         );
  NAND2_X1 U11515 ( .A1(n8626), .A2(n9096), .ZN(n9097) );
  NAND2_X1 U11516 ( .A1(n9098), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9099) );
  MUX2_X1 U11517 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9099), .S(
        P3_IR_REG_23__SCAN_IN), .Z(n9101) );
  NAND2_X1 U11518 ( .A1(n9101), .A2(n9100), .ZN(n9723) );
  NAND2_X1 U11519 ( .A1(n9195), .A2(n9856), .ZN(n9722) );
  OAI21_X1 U11520 ( .B1(n9104), .B2(n9103), .A(n12533), .ZN(n9132) );
  INV_X1 U11521 ( .A(n12886), .ZN(n12767) );
  NAND2_X1 U11522 ( .A1(n9934), .A2(n14441), .ZN(n9105) );
  OR2_X1 U11523 ( .A1(n9933), .A2(n9105), .ZN(n9107) );
  NOR2_X1 U11524 ( .A1(n15099), .A2(n12104), .ZN(n9106) );
  INV_X1 U11525 ( .A(n12524), .ZN(n12544) );
  NAND2_X1 U11526 ( .A1(n9933), .A2(n10040), .ZN(n9111) );
  INV_X1 U11527 ( .A(n9929), .ZN(n9109) );
  INV_X1 U11528 ( .A(n12691), .ZN(n12700) );
  NAND2_X1 U11529 ( .A1(n10611), .A2(n12700), .ZN(n12103) );
  NAND2_X1 U11530 ( .A1(n6529), .A2(n12103), .ZN(n9865) );
  NAND2_X1 U11531 ( .A1(n9195), .A2(n9865), .ZN(n9108) );
  AOI21_X1 U11532 ( .B1(n9930), .B2(n9109), .A(n9108), .ZN(n9110) );
  NAND2_X1 U11533 ( .A1(n9111), .A2(n9110), .ZN(n9113) );
  INV_X1 U11534 ( .A(n12103), .ZN(n10036) );
  NAND2_X1 U11535 ( .A1(n6529), .A2(n10036), .ZN(n9928) );
  NOR2_X1 U11536 ( .A1(n9722), .A2(n9928), .ZN(n12112) );
  AND2_X1 U11537 ( .A1(n9930), .A2(n12112), .ZN(n9112) );
  AOI21_X1 U11538 ( .B1(n9113), .B2(P3_STATE_REG_SCAN_IN), .A(n9112), .ZN(
        n9857) );
  INV_X1 U11539 ( .A(n9723), .ZN(n9114) );
  NAND2_X1 U11540 ( .A1(n9114), .A2(P3_STATE_REG_SCAN_IN), .ZN(n12116) );
  NAND2_X1 U11541 ( .A1(n9934), .A2(n10036), .ZN(n9115) );
  NOR2_X1 U11542 ( .A1(n9930), .A2(n9115), .ZN(n9126) );
  AND2_X1 U11543 ( .A1(n9724), .A2(n9730), .ZN(n9124) );
  AND2_X2 U11544 ( .A1(n9124), .A2(n6529), .ZN(n15038) );
  NAND2_X1 U11545 ( .A1(n9117), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n9118) );
  NAND2_X1 U11546 ( .A1(n9149), .A2(n9118), .ZN(n12753) );
  NAND2_X1 U11547 ( .A1(n12753), .A2(n8697), .ZN(n9123) );
  INV_X1 U11548 ( .A(P3_REG0_REG_26__SCAN_IN), .ZN(n12939) );
  NAND2_X1 U11549 ( .A1(n11899), .A2(P3_REG2_REG_26__SCAN_IN), .ZN(n9120) );
  NAND2_X1 U11550 ( .A1(n6542), .A2(P3_REG1_REG_26__SCAN_IN), .ZN(n9119) );
  OAI211_X1 U11551 ( .C1(n6525), .C2(n12939), .A(n9120), .B(n9119), .ZN(n9121)
         );
  INV_X1 U11552 ( .A(n9121), .ZN(n9122) );
  INV_X1 U11553 ( .A(n9124), .ZN(n9125) );
  AND2_X2 U11554 ( .A1(n9125), .A2(n6529), .ZN(n15052) );
  NAND2_X1 U11555 ( .A1(n9126), .A2(n15052), .ZN(n12484) );
  AOI22_X1 U11556 ( .A1(n12761), .A2(n12535), .B1(P3_REG3_REG_25__SCAN_IN), 
        .B2(P3_U3151), .ZN(n9127) );
  OAI21_X1 U11557 ( .B1(n11811), .B2(n12537), .A(n9127), .ZN(n9128) );
  AOI21_X1 U11558 ( .B1(n12764), .B2(n12540), .A(n9128), .ZN(n9129) );
  NAND2_X1 U11559 ( .A1(n9132), .A2(n9131), .ZN(P3_U3165) );
  NOR2_X1 U11560 ( .A1(P1_DATAO_REG_25__SCAN_IN), .A2(n15212), .ZN(n9133) );
  AOI22_X1 U11561 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(n13595), .B1(
        P1_DATAO_REG_26__SCAN_IN), .B2(n15197), .ZN(n9135) );
  INV_X1 U11562 ( .A(n9135), .ZN(n9136) );
  XNOR2_X1 U11563 ( .A(n11463), .B(n9136), .ZN(n13019) );
  NAND2_X1 U11564 ( .A1(n13019), .A2(n11913), .ZN(n9138) );
  OR2_X1 U11565 ( .A1(n9031), .A2(n13021), .ZN(n9137) );
  XNOR2_X1 U11566 ( .A(n12940), .B(n8709), .ZN(n9139) );
  NOR2_X1 U11567 ( .A1(n9139), .A2(n12761), .ZN(n12121) );
  AOI21_X1 U11568 ( .B1(n12761), .B2(n9139), .A(n12121), .ZN(n9146) );
  AND2_X1 U11569 ( .A1(n9141), .A2(n9140), .ZN(n9144) );
  AND2_X1 U11570 ( .A1(n9143), .A2(n9146), .ZN(n12120) );
  INV_X1 U11571 ( .A(n9146), .ZN(n9145) );
  INV_X1 U11572 ( .A(n12940), .ZN(n9159) );
  INV_X1 U11573 ( .A(n9149), .ZN(n9148) );
  INV_X1 U11574 ( .A(P3_REG3_REG_27__SCAN_IN), .ZN(n9147) );
  NAND2_X1 U11575 ( .A1(n9148), .A2(n9147), .ZN(n10142) );
  NAND2_X1 U11576 ( .A1(n9149), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n9150) );
  NAND2_X1 U11577 ( .A1(n10142), .A2(n9150), .ZN(n12741) );
  NAND2_X1 U11578 ( .A1(n12741), .A2(n8697), .ZN(n9155) );
  INV_X1 U11579 ( .A(P3_REG0_REG_27__SCAN_IN), .ZN(n12935) );
  NAND2_X1 U11580 ( .A1(n6542), .A2(P3_REG1_REG_27__SCAN_IN), .ZN(n9152) );
  NAND2_X1 U11581 ( .A1(n11899), .A2(P3_REG2_REG_27__SCAN_IN), .ZN(n9151) );
  OAI211_X1 U11582 ( .C1(n12935), .C2(n6525), .A(n9152), .B(n9151), .ZN(n9153)
         );
  INV_X1 U11583 ( .A(n9153), .ZN(n9154) );
  INV_X1 U11584 ( .A(n12750), .ZN(n11845) );
  AOI22_X1 U11585 ( .A1(n12773), .A2(n12525), .B1(P3_REG3_REG_26__SCAN_IN), 
        .B2(P3_U3151), .ZN(n9156) );
  OAI21_X1 U11586 ( .B1(n11845), .B2(n12484), .A(n9156), .ZN(n9157) );
  AOI21_X1 U11587 ( .B1(n12753), .B2(n12540), .A(n9157), .ZN(n9158) );
  OAI21_X1 U11588 ( .B1(n9159), .B2(n12544), .A(n9158), .ZN(n9160) );
  NAND2_X1 U11589 ( .A1(n9162), .A2(n9161), .ZN(P3_U3180) );
  NOR2_X1 U11590 ( .A1(n9536), .A2(n9163), .ZN(n9537) );
  NAND4_X1 U11591 ( .A1(n9584), .A2(n9168), .A3(n9167), .A4(n9166), .ZN(n9953)
         );
  NAND3_X1 U11592 ( .A1(n9488), .A2(n9170), .A3(n9169), .ZN(n9171) );
  NOR2_X1 U11593 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), 
        .ZN(n9175) );
  NOR2_X1 U11594 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), 
        .ZN(n9174) );
  NOR2_X1 U11595 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_20__SCAN_IN), 
        .ZN(n9173) );
  INV_X1 U11596 ( .A(n9180), .ZN(n9176) );
  NAND2_X1 U11597 ( .A1(n9190), .A2(n9177), .ZN(n9193) );
  NAND2_X1 U11598 ( .A1(n9183), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9178) );
  MUX2_X1 U11599 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9178), .S(
        P1_IR_REG_25__SCAN_IN), .Z(n9181) );
  NOR3_X1 U11600 ( .A1(P1_IR_REG_23__SCAN_IN), .A2(P1_IR_REG_24__SCAN_IN), 
        .A3(P1_IR_REG_25__SCAN_IN), .ZN(n9179) );
  NAND2_X1 U11601 ( .A1(n9193), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9182) );
  MUX2_X1 U11602 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9182), .S(
        P1_IR_REG_24__SCAN_IN), .Z(n9184) );
  NAND2_X1 U11603 ( .A1(n9185), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9186) );
  MUX2_X1 U11604 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9186), .S(
        P1_IR_REG_26__SCAN_IN), .Z(n9189) );
  INV_X1 U11605 ( .A(n9188), .ZN(n9340) );
  INV_X1 U11606 ( .A(n9190), .ZN(n9191) );
  NAND2_X1 U11607 ( .A1(n9191), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9192) );
  MUX2_X1 U11608 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9192), .S(
        P1_IR_REG_23__SCAN_IN), .Z(n9194) );
  NAND2_X1 U11609 ( .A1(n9194), .A2(n9193), .ZN(n9592) );
  NAND2_X1 U11610 ( .A1(n9592), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9433) );
  INV_X1 U11611 ( .A(n9856), .ZN(n13002) );
  NAND2_X1 U11612 ( .A1(n13405), .A2(n9196), .ZN(n9197) );
  XNOR2_X1 U11613 ( .A(n13359), .B(n9271), .ZN(n11861) );
  NAND2_X1 U11614 ( .A1(n13144), .A2(n13269), .ZN(n11862) );
  XNOR2_X1 U11615 ( .A(n11861), .B(n11862), .ZN(n9296) );
  NAND2_X1 U11616 ( .A1(n7753), .A2(n13269), .ZN(n9199) );
  XNOR2_X1 U11617 ( .A(n9197), .B(n10824), .ZN(n10428) );
  XNOR2_X1 U11618 ( .A(n9199), .B(n10428), .ZN(n10337) );
  INV_X1 U11619 ( .A(n10208), .ZN(n10336) );
  AND2_X1 U11620 ( .A1(n9271), .A2(n10358), .ZN(n10335) );
  AOI21_X1 U11621 ( .B1(n10336), .B2(n13269), .A(n10335), .ZN(n9198) );
  NAND2_X1 U11622 ( .A1(n10337), .A2(n9198), .ZN(n10429) );
  INV_X1 U11623 ( .A(n10428), .ZN(n9200) );
  NAND2_X1 U11624 ( .A1(n9200), .A2(n9199), .ZN(n9201) );
  NAND2_X1 U11625 ( .A1(n10429), .A2(n9201), .ZN(n9202) );
  XNOR2_X1 U11626 ( .A(n10474), .B(n9197), .ZN(n9203) );
  NAND2_X1 U11627 ( .A1(n8301), .A2(n13269), .ZN(n9204) );
  XNOR2_X1 U11628 ( .A(n9203), .B(n9204), .ZN(n10430) );
  NAND2_X1 U11629 ( .A1(n9202), .A2(n10430), .ZN(n10436) );
  INV_X1 U11630 ( .A(n9203), .ZN(n9205) );
  NAND2_X1 U11631 ( .A1(n9205), .A2(n9204), .ZN(n9206) );
  NAND2_X1 U11632 ( .A1(n10436), .A2(n9206), .ZN(n13046) );
  XNOR2_X1 U11633 ( .A(n13050), .B(n9239), .ZN(n11879) );
  AND2_X1 U11634 ( .A1(n13159), .A2(n13269), .ZN(n9207) );
  NAND2_X1 U11635 ( .A1(n11879), .A2(n9207), .ZN(n9211) );
  INV_X1 U11636 ( .A(n11879), .ZN(n9209) );
  INV_X1 U11637 ( .A(n9207), .ZN(n9208) );
  NAND2_X1 U11638 ( .A1(n9209), .A2(n9208), .ZN(n9210) );
  NAND2_X1 U11639 ( .A1(n9211), .A2(n9210), .ZN(n13045) );
  OR2_X1 U11640 ( .A1(n13046), .A2(n13045), .ZN(n13047) );
  XNOR2_X1 U11641 ( .A(n14898), .B(n9239), .ZN(n10342) );
  NAND2_X1 U11642 ( .A1(n13158), .A2(n13269), .ZN(n9212) );
  XNOR2_X1 U11643 ( .A(n10342), .B(n9212), .ZN(n11878) );
  NAND3_X1 U11644 ( .A1(n13047), .A2(n11878), .A3(n9211), .ZN(n11890) );
  INV_X1 U11645 ( .A(n10342), .ZN(n9213) );
  NAND2_X1 U11646 ( .A1(n9213), .A2(n9212), .ZN(n9214) );
  XNOR2_X1 U11647 ( .A(n10479), .B(n9239), .ZN(n9215) );
  NAND2_X1 U11648 ( .A1(n13157), .A2(n13269), .ZN(n9216) );
  XNOR2_X1 U11649 ( .A(n9215), .B(n9216), .ZN(n10343) );
  INV_X1 U11650 ( .A(n9215), .ZN(n9217) );
  NAND2_X1 U11651 ( .A1(n9217), .A2(n9216), .ZN(n9218) );
  XNOR2_X1 U11652 ( .A(n10487), .B(n9239), .ZN(n9219) );
  AND2_X1 U11653 ( .A1(n13156), .A2(n13269), .ZN(n9220) );
  NAND2_X1 U11654 ( .A1(n9219), .A2(n9220), .ZN(n9224) );
  INV_X1 U11655 ( .A(n9219), .ZN(n10121) );
  INV_X1 U11656 ( .A(n9220), .ZN(n9221) );
  NAND2_X1 U11657 ( .A1(n10121), .A2(n9221), .ZN(n9222) );
  NAND2_X1 U11658 ( .A1(n9224), .A2(n9222), .ZN(n10269) );
  XNOR2_X1 U11659 ( .A(n10484), .B(n9239), .ZN(n9225) );
  AND2_X1 U11660 ( .A1(n13155), .A2(n13269), .ZN(n9226) );
  NAND2_X1 U11661 ( .A1(n9225), .A2(n9226), .ZN(n9230) );
  INV_X1 U11662 ( .A(n9225), .ZN(n10287) );
  INV_X1 U11663 ( .A(n9226), .ZN(n9227) );
  NAND2_X1 U11664 ( .A1(n10287), .A2(n9227), .ZN(n9228) );
  AND2_X1 U11665 ( .A1(n9230), .A2(n9228), .ZN(n10118) );
  NAND2_X1 U11666 ( .A1(n9229), .A2(n10118), .ZN(n10281) );
  XNOR2_X1 U11667 ( .A(n10741), .B(n9239), .ZN(n10573) );
  NAND2_X1 U11668 ( .A1(n13154), .A2(n13269), .ZN(n9231) );
  XNOR2_X1 U11669 ( .A(n10573), .B(n9231), .ZN(n10288) );
  NAND3_X1 U11670 ( .A1(n10281), .A2(n10288), .A3(n9230), .ZN(n10282) );
  INV_X1 U11671 ( .A(n10573), .ZN(n9232) );
  NAND2_X1 U11672 ( .A1(n9232), .A2(n9231), .ZN(n9233) );
  NAND2_X1 U11673 ( .A1(n10282), .A2(n9233), .ZN(n9234) );
  XNOR2_X1 U11674 ( .A(n10750), .B(n9239), .ZN(n9235) );
  NAND2_X1 U11675 ( .A1(n13153), .A2(n13269), .ZN(n9236) );
  XNOR2_X1 U11676 ( .A(n9235), .B(n9236), .ZN(n10574) );
  NAND2_X1 U11677 ( .A1(n9234), .A2(n10574), .ZN(n10580) );
  INV_X1 U11678 ( .A(n9235), .ZN(n9237) );
  NAND2_X1 U11679 ( .A1(n9237), .A2(n9236), .ZN(n9238) );
  NAND2_X1 U11680 ( .A1(n10580), .A2(n9238), .ZN(n9311) );
  XNOR2_X1 U11681 ( .A(n10779), .B(n9239), .ZN(n9240) );
  AND2_X1 U11682 ( .A1(n13152), .A2(n13269), .ZN(n9241) );
  NAND2_X1 U11683 ( .A1(n9240), .A2(n9241), .ZN(n9246) );
  INV_X1 U11684 ( .A(n9240), .ZN(n10804) );
  INV_X1 U11685 ( .A(n9241), .ZN(n9242) );
  NAND2_X1 U11686 ( .A1(n10804), .A2(n9242), .ZN(n9243) );
  NAND2_X1 U11687 ( .A1(n9246), .A2(n9243), .ZN(n9312) );
  XNOR2_X1 U11688 ( .A(n10860), .B(n13024), .ZN(n10928) );
  NAND2_X1 U11689 ( .A1(n13151), .A2(n13269), .ZN(n9247) );
  XNOR2_X1 U11690 ( .A(n10928), .B(n9247), .ZN(n10805) );
  NAND3_X1 U11691 ( .A1(n9310), .A2(n10805), .A3(n9246), .ZN(n10799) );
  INV_X1 U11692 ( .A(n10928), .ZN(n9248) );
  NAND2_X1 U11693 ( .A1(n9248), .A2(n9247), .ZN(n9249) );
  NAND2_X1 U11694 ( .A1(n10799), .A2(n9249), .ZN(n9250) );
  XNOR2_X1 U11695 ( .A(n14516), .B(n13024), .ZN(n9251) );
  NAND2_X1 U11696 ( .A1(n13150), .A2(n13269), .ZN(n9252) );
  XNOR2_X1 U11697 ( .A(n9251), .B(n9252), .ZN(n10929) );
  INV_X1 U11698 ( .A(n9251), .ZN(n9253) );
  NAND2_X1 U11699 ( .A1(n9253), .A2(n9252), .ZN(n9254) );
  NAND2_X1 U11700 ( .A1(n10935), .A2(n9254), .ZN(n11114) );
  XNOR2_X1 U11701 ( .A(n13441), .B(n13024), .ZN(n9255) );
  AND2_X1 U11702 ( .A1(n13149), .A2(n13269), .ZN(n9256) );
  NAND2_X1 U11703 ( .A1(n9255), .A2(n9256), .ZN(n9260) );
  INV_X1 U11704 ( .A(n9255), .ZN(n9258) );
  INV_X1 U11705 ( .A(n9256), .ZN(n9257) );
  NAND2_X1 U11706 ( .A1(n9258), .A2(n9257), .ZN(n9259) );
  NAND2_X1 U11707 ( .A1(n9260), .A2(n9259), .ZN(n11115) );
  XNOR2_X1 U11708 ( .A(n11233), .B(n13024), .ZN(n9261) );
  NAND2_X1 U11709 ( .A1(n13148), .A2(n13269), .ZN(n9262) );
  XNOR2_X1 U11710 ( .A(n9261), .B(n9262), .ZN(n14457) );
  INV_X1 U11711 ( .A(n9261), .ZN(n9263) );
  XNOR2_X1 U11712 ( .A(n14489), .B(n13024), .ZN(n9265) );
  AND2_X1 U11713 ( .A1(n13147), .A2(n13269), .ZN(n9264) );
  NAND2_X1 U11714 ( .A1(n11329), .A2(n9264), .ZN(n11330) );
  INV_X1 U11715 ( .A(n9265), .ZN(n9266) );
  OR2_X1 U11716 ( .A1(n9267), .A2(n9266), .ZN(n9268) );
  XNOR2_X1 U11717 ( .A(n14480), .B(n9271), .ZN(n11436) );
  NAND2_X1 U11718 ( .A1(n13146), .A2(n13269), .ZN(n9269) );
  XNOR2_X1 U11719 ( .A(n11436), .B(n9269), .ZN(n14472) );
  NAND2_X1 U11720 ( .A1(n11436), .A2(n9269), .ZN(n9270) );
  XNOR2_X1 U11721 ( .A(n14498), .B(n13024), .ZN(n9272) );
  NAND2_X1 U11722 ( .A1(n13400), .A2(n13269), .ZN(n9273) );
  XNOR2_X1 U11723 ( .A(n9272), .B(n9273), .ZN(n11435) );
  INV_X1 U11724 ( .A(n9272), .ZN(n9274) );
  XNOR2_X1 U11725 ( .A(n13521), .B(n13024), .ZN(n9275) );
  AND2_X1 U11726 ( .A1(n13145), .A2(n13269), .ZN(n9276) );
  NAND2_X1 U11727 ( .A1(n9275), .A2(n9276), .ZN(n9279) );
  INV_X1 U11728 ( .A(n9275), .ZN(n13055) );
  INV_X1 U11729 ( .A(n9276), .ZN(n9277) );
  NAND2_X1 U11730 ( .A1(n13055), .A2(n9277), .ZN(n9278) );
  NAND2_X1 U11731 ( .A1(n9279), .A2(n9278), .ZN(n13119) );
  XNOR2_X1 U11732 ( .A(n13516), .B(n13024), .ZN(n9281) );
  NAND2_X1 U11733 ( .A1(n13403), .A2(n13269), .ZN(n9282) );
  XNOR2_X1 U11734 ( .A(n9281), .B(n9282), .ZN(n13061) );
  AND2_X1 U11735 ( .A1(n13061), .A2(n9279), .ZN(n9280) );
  INV_X1 U11736 ( .A(n9281), .ZN(n13098) );
  XNOR2_X1 U11737 ( .A(n13511), .B(n13024), .ZN(n9284) );
  NAND2_X1 U11738 ( .A1(n13355), .A2(n13269), .ZN(n9285) );
  XNOR2_X1 U11739 ( .A(n9284), .B(n9285), .ZN(n13097) );
  INV_X1 U11740 ( .A(n9284), .ZN(n9286) );
  NAND2_X1 U11741 ( .A1(n9286), .A2(n9285), .ZN(n9287) );
  INV_X1 U11742 ( .A(n10357), .ZN(n9290) );
  NOR2_X1 U11743 ( .A1(n14899), .A2(n9291), .ZN(n9292) );
  INV_X1 U11744 ( .A(n11866), .ZN(n9294) );
  AOI211_X1 U11745 ( .C1(n9296), .C2(n9295), .A(n14474), .B(n9294), .ZN(n9309)
         );
  INV_X1 U11746 ( .A(n13359), .ZN(n13567) );
  NAND2_X1 U11747 ( .A1(n9963), .A2(n14488), .ZN(n9297) );
  INV_X1 U11748 ( .A(n14479), .ZN(n14458) );
  NOR2_X1 U11749 ( .A1(n13567), .A2(n14458), .ZN(n9308) );
  INV_X1 U11750 ( .A(n14890), .ZN(n10195) );
  NAND2_X1 U11751 ( .A1(n10195), .A2(n9298), .ZN(n9299) );
  OR2_X1 U11752 ( .A1(n10194), .A2(n9299), .ZN(n9300) );
  NAND2_X1 U11753 ( .A1(n9300), .A2(n10192), .ZN(n9302) );
  NAND2_X1 U11754 ( .A1(n9302), .A2(n9301), .ZN(n9958) );
  OAI22_X1 U11755 ( .A1(n14467), .A2(n13360), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n15385), .ZN(n9307) );
  NAND2_X1 U11756 ( .A1(n13131), .A2(n13401), .ZN(n14470) );
  NAND2_X1 U11757 ( .A1(n13131), .A2(n13402), .ZN(n14469) );
  OAI22_X1 U11758 ( .A1(n9305), .A2(n14470), .B1(n14469), .B2(n9304), .ZN(
        n9306) );
  OR4_X1 U11759 ( .A1(n9309), .A2(n9308), .A3(n9307), .A4(n9306), .ZN(P2_U3195) );
  INV_X1 U11760 ( .A(n9310), .ZN(n10801) );
  AOI211_X1 U11761 ( .C1(n9312), .C2(n9311), .A(n14474), .B(n10801), .ZN(n9316) );
  INV_X1 U11762 ( .A(n10779), .ZN(n14914) );
  NOR2_X1 U11763 ( .A1(n14914), .A2(n14458), .ZN(n9315) );
  INV_X1 U11764 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n15210) );
  OAI22_X1 U11765 ( .A1(n14467), .A2(n10774), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n15210), .ZN(n9314) );
  OAI22_X1 U11766 ( .A1(n10770), .A2(n14470), .B1(n14469), .B2(n10769), .ZN(
        n9313) );
  OR4_X1 U11767 ( .A1(n9316), .A2(n9315), .A3(n9314), .A4(n9313), .ZN(P2_U3189) );
  NAND2_X1 U11768 ( .A1(n9319), .A2(n9320), .ZN(n14242) );
  INV_X1 U11769 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n9318) );
  XNOR2_X2 U11770 ( .A(n9321), .B(n9320), .ZN(n12387) );
  INV_X2 U11771 ( .A(n6540), .ZN(n11783) );
  NAND2_X1 U11772 ( .A1(n11783), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n9329) );
  NAND2_X4 U11773 ( .A1(n9323), .A2(n9322), .ZN(n11600) );
  INV_X1 U11774 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n14660) );
  OR2_X1 U11775 ( .A1(n6526), .A2(n14660), .ZN(n9327) );
  INV_X1 U11776 ( .A(n12321), .ZN(n9325) );
  INV_X1 U11777 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n9324) );
  OR2_X1 U11778 ( .A1(n9325), .A2(n9324), .ZN(n9326) );
  INV_X1 U11779 ( .A(n9335), .ZN(n9333) );
  NAND2_X1 U11780 ( .A1(n9350), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9334) );
  NAND2_X1 U11781 ( .A1(n9335), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9337) );
  INV_X1 U11782 ( .A(n12159), .ZN(n10295) );
  AND2_X2 U11783 ( .A1(n10295), .A2(n9443), .ZN(n10439) );
  INV_X1 U11784 ( .A(n11701), .ZN(n9413) );
  NAND2_X1 U11785 ( .A1(n13776), .A2(n9413), .ZN(n9349) );
  XNOR2_X2 U11786 ( .A(n9339), .B(n9338), .ZN(n9450) );
  OR2_X1 U11787 ( .A1(n10388), .A2(n9487), .ZN(n9347) );
  OR2_X1 U11788 ( .A1(n12317), .A2(n9476), .ZN(n9346) );
  NAND2_X1 U11789 ( .A1(n9343), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9344) );
  XNOR2_X1 U11790 ( .A(n9344), .B(n9165), .ZN(n9625) );
  OR2_X1 U11791 ( .A1(n11572), .A2(n9625), .ZN(n9345) );
  AND3_X2 U11792 ( .A1(n9347), .A2(n9346), .A3(n9345), .ZN(n14714) );
  OR2_X1 U11793 ( .A1(n14714), .A2(n11702), .ZN(n9348) );
  NAND2_X1 U11794 ( .A1(n9349), .A2(n9348), .ZN(n9356) );
  INV_X1 U11795 ( .A(n9351), .ZN(n9352) );
  NAND2_X1 U11796 ( .A1(n9352), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9353) );
  MUX2_X1 U11797 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9353), .S(
        P1_IR_REG_19__SCAN_IN), .Z(n9354) );
  NAND2_X1 U11798 ( .A1(n14251), .A2(n13868), .ZN(n9355) );
  AND2_X2 U11799 ( .A1(n9355), .A2(n12159), .ZN(n11745) );
  XNOR2_X1 U11800 ( .A(n9356), .B(n11745), .ZN(n10438) );
  AND2_X2 U11801 ( .A1(n14663), .A2(n11778), .ZN(n10452) );
  INV_X1 U11802 ( .A(n14714), .ZN(n14664) );
  AOI22_X1 U11803 ( .A1(n13776), .A2(n10452), .B1(n14664), .B2(n9413), .ZN(
        n10437) );
  XNOR2_X1 U11804 ( .A(n10438), .B(n10437), .ZN(n9440) );
  NAND2_X1 U11805 ( .A1(n12321), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n9362) );
  INV_X1 U11806 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n10529) );
  OR2_X1 U11807 ( .A1(n11600), .A2(n10529), .ZN(n9361) );
  INV_X1 U11808 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n9358) );
  INV_X1 U11809 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n9596) );
  NAND2_X1 U11810 ( .A1(n6770), .A2(n10439), .ZN(n9370) );
  MUX2_X1 U11811 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9363), .S(
        P1_IR_REG_1__SCAN_IN), .Z(n9366) );
  INV_X1 U11812 ( .A(n9403), .ZN(n9365) );
  NAND2_X1 U11813 ( .A1(n12163), .A2(n11778), .ZN(n9369) );
  NAND2_X1 U11814 ( .A1(n9370), .A2(n9369), .ZN(n9371) );
  XNOR2_X1 U11815 ( .A(n9371), .B(n11745), .ZN(n9373) );
  AND2_X1 U11816 ( .A1(n10439), .A2(n12163), .ZN(n9372) );
  NAND2_X1 U11817 ( .A1(n9373), .A2(n9374), .ZN(n9395) );
  INV_X1 U11818 ( .A(n9373), .ZN(n9376) );
  INV_X1 U11819 ( .A(n9374), .ZN(n9375) );
  NAND2_X1 U11820 ( .A1(n9376), .A2(n9375), .ZN(n9377) );
  NAND2_X1 U11821 ( .A1(n9395), .A2(n9377), .ZN(n10013) );
  INV_X1 U11822 ( .A(n10013), .ZN(n9394) );
  NAND2_X1 U11823 ( .A1(n12321), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n9382) );
  INV_X1 U11824 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n9378) );
  INV_X1 U11825 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n9603) );
  OR2_X1 U11826 ( .A1(n6526), .A2(n9603), .ZN(n9380) );
  INV_X1 U11827 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n9387) );
  NAND2_X1 U11828 ( .A1(n13780), .A2(n10439), .ZN(n9390) );
  INV_X1 U11829 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n14602) );
  INV_X1 U11830 ( .A(SI_0_), .ZN(n9384) );
  OAI21_X1 U11831 ( .B1(n9473), .B2(n9384), .A(n9383), .ZN(n9385) );
  NAND2_X1 U11832 ( .A1(n9386), .A2(n9385), .ZN(n14252) );
  MUX2_X1 U11833 ( .A(n14602), .B(n14252), .S(n11572), .Z(n14677) );
  OAI22_X1 U11834 ( .A1(n14677), .A2(n11702), .B1(n9443), .B2(n9387), .ZN(
        n9388) );
  INV_X1 U11835 ( .A(n9388), .ZN(n9389) );
  NAND2_X1 U11836 ( .A1(n9390), .A2(n9389), .ZN(n9893) );
  OR2_X1 U11837 ( .A1(n9893), .A2(n11745), .ZN(n9392) );
  OAI22_X1 U11838 ( .A1(n14677), .A2(n11701), .B1(n9443), .B2(n14602), .ZN(
        n9391) );
  NAND2_X1 U11839 ( .A1(n9893), .A2(n9894), .ZN(n9896) );
  NAND2_X1 U11840 ( .A1(n10011), .A2(n9395), .ZN(n9987) );
  NAND2_X1 U11841 ( .A1(n12321), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n9401) );
  INV_X1 U11842 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n9396) );
  INV_X1 U11843 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n9397) );
  INV_X1 U11844 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n9597) );
  NAND2_X1 U11845 ( .A1(n13778), .A2(n9413), .ZN(n9411) );
  OR2_X1 U11846 ( .A1(n10388), .A2(n9503), .ZN(n9409) );
  INV_X1 U11847 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n9502) );
  OR2_X1 U11848 ( .A1(n9402), .A2(n9502), .ZN(n9408) );
  NOR2_X1 U11849 ( .A1(n9403), .A2(n9318), .ZN(n9404) );
  INV_X1 U11850 ( .A(n9405), .ZN(n9406) );
  NAND2_X1 U11851 ( .A1(n9406), .A2(n9343), .ZN(n9909) );
  OR2_X1 U11852 ( .A1(n11572), .A2(n9909), .ZN(n9407) );
  AND3_X2 U11853 ( .A1(n9409), .A2(n9408), .A3(n9407), .ZN(n10298) );
  OR2_X1 U11854 ( .A1(n10298), .A2(n11702), .ZN(n9410) );
  NAND2_X1 U11855 ( .A1(n9411), .A2(n9410), .ZN(n9412) );
  XNOR2_X1 U11856 ( .A(n9412), .B(n11775), .ZN(n9414) );
  AOI22_X1 U11857 ( .A1(n13778), .A2(n10452), .B1(n14706), .B2(n9413), .ZN(
        n9415) );
  INV_X1 U11858 ( .A(n9414), .ZN(n9416) );
  NAND2_X1 U11859 ( .A1(n9416), .A2(n9415), .ZN(n9417) );
  INV_X1 U11860 ( .A(P1_B_REG_SCAN_IN), .ZN(n15224) );
  NOR2_X1 U11861 ( .A1(n11428), .A2(n15224), .ZN(n9418) );
  MUX2_X1 U11862 ( .A(n15224), .B(n9418), .S(n11348), .Z(n9419) );
  NOR2_X1 U11863 ( .A1(n9419), .A2(n14249), .ZN(n9513) );
  INV_X1 U11864 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n9420) );
  NAND2_X1 U11865 ( .A1(n9513), .A2(n9420), .ZN(n9421) );
  NAND2_X1 U11866 ( .A1(n11348), .A2(n14249), .ZN(n9514) );
  INV_X1 U11867 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n9518) );
  INV_X1 U11868 ( .A(n14249), .ZN(n9422) );
  NOR2_X1 U11869 ( .A1(n11428), .A2(n9422), .ZN(n9517) );
  AOI21_X1 U11870 ( .B1(n9513), .B2(n9518), .A(n9517), .ZN(n14123) );
  NOR2_X1 U11871 ( .A1(P1_D_REG_7__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .ZN(
        n9426) );
  NOR4_X1 U11872 ( .A1(P1_D_REG_28__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_29__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n9425) );
  NOR4_X1 U11873 ( .A1(P1_D_REG_5__SCAN_IN), .A2(P1_D_REG_6__SCAN_IN), .A3(
        P1_D_REG_9__SCAN_IN), .A4(P1_D_REG_10__SCAN_IN), .ZN(n9424) );
  NOR4_X1 U11874 ( .A1(P1_D_REG_8__SCAN_IN), .A2(P1_D_REG_2__SCAN_IN), .A3(
        P1_D_REG_3__SCAN_IN), .A4(P1_D_REG_4__SCAN_IN), .ZN(n9423) );
  NAND4_X1 U11875 ( .A1(n9426), .A2(n9425), .A3(n9424), .A4(n9423), .ZN(n9432)
         );
  NOR4_X1 U11876 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_16__SCAN_IN), .A3(
        P1_D_REG_17__SCAN_IN), .A4(P1_D_REG_18__SCAN_IN), .ZN(n9430) );
  NOR4_X1 U11877 ( .A1(P1_D_REG_13__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_14__SCAN_IN), .ZN(n9429) );
  NOR4_X1 U11878 ( .A1(P1_D_REG_23__SCAN_IN), .A2(P1_D_REG_25__SCAN_IN), .A3(
        P1_D_REG_26__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n9428) );
  NOR4_X1 U11879 ( .A1(P1_D_REG_19__SCAN_IN), .A2(P1_D_REG_20__SCAN_IN), .A3(
        P1_D_REG_21__SCAN_IN), .A4(P1_D_REG_22__SCAN_IN), .ZN(n9427) );
  NAND4_X1 U11880 ( .A1(n9430), .A2(n9429), .A3(n9428), .A4(n9427), .ZN(n9431)
         );
  OAI21_X1 U11881 ( .B1(n9432), .B2(n9431), .A(n9513), .ZN(n9458) );
  NAND3_X1 U11882 ( .A1(n14221), .A2(n14123), .A3(n9458), .ZN(n9441) );
  OR2_X1 U11883 ( .A1(n9441), .A2(n9595), .ZN(n9449) );
  INV_X1 U11884 ( .A(n9449), .ZN(n9436) );
  INV_X1 U11885 ( .A(n12143), .ZN(n12142) );
  NAND2_X1 U11886 ( .A1(n6773), .A2(n12142), .ZN(n12375) );
  OR2_X1 U11887 ( .A1(n12375), .A2(n6796), .ZN(n10314) );
  OAI21_X2 U11888 ( .B1(n9434), .B2(n13868), .A(n10314), .ZN(n14742) );
  NAND2_X1 U11889 ( .A1(n6796), .A2(n9357), .ZN(n12146) );
  INV_X1 U11890 ( .A(n12146), .ZN(n9451) );
  NOR2_X1 U11891 ( .A1(n14742), .A2(n9451), .ZN(n9435) );
  INV_X1 U11892 ( .A(n10450), .ZN(n9438) );
  AOI211_X1 U11893 ( .C1(n9440), .C2(n9439), .A(n13727), .B(n9438), .ZN(n9461)
         );
  NAND2_X1 U11894 ( .A1(n12143), .A2(n11534), .ZN(n14679) );
  INV_X1 U11895 ( .A(n14220), .ZN(n14126) );
  NAND2_X1 U11896 ( .A1(n9441), .A2(n14126), .ZN(n9446) );
  AND2_X1 U11897 ( .A1(n12143), .A2(n13868), .ZN(n9442) );
  OR2_X1 U11898 ( .A1(n12146), .A2(n9442), .ZN(n9990) );
  AND2_X1 U11899 ( .A1(n9443), .A2(n9592), .ZN(n9444) );
  NAND2_X1 U11900 ( .A1(n9990), .A2(n9444), .ZN(n9457) );
  INV_X1 U11901 ( .A(n9457), .ZN(n9445) );
  NAND2_X1 U11902 ( .A1(n9446), .A2(n9445), .ZN(n9447) );
  INV_X1 U11903 ( .A(n14542), .ZN(n13717) );
  MUX2_X1 U11904 ( .A(n13717), .B(P1_U3086), .S(P1_REG3_REG_3__SCAN_IN), .Z(
        n9460) );
  NAND2_X1 U11905 ( .A1(n9449), .A2(n14659), .ZN(n13601) );
  INV_X1 U11906 ( .A(n14533), .ZN(n13753) );
  INV_X1 U11907 ( .A(n9450), .ZN(n9899) );
  AND2_X2 U11908 ( .A1(n9451), .A2(n9899), .ZN(n13897) );
  NAND2_X1 U11909 ( .A1(n11783), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n9456) );
  INV_X1 U11910 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n9452) );
  OR2_X1 U11911 ( .A1(n11784), .A2(n9452), .ZN(n9455) );
  NAND2_X1 U11912 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n9756) );
  OAI21_X1 U11913 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(n9756), .ZN(n10631) );
  OR2_X1 U11914 ( .A1(n11600), .A2(n10631), .ZN(n9454) );
  INV_X1 U11915 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n10313) );
  OR2_X1 U11916 ( .A1(n6526), .A2(n10313), .ZN(n9453) );
  OR2_X1 U11917 ( .A1(n12146), .A2(n9899), .ZN(n14678) );
  AOI22_X1 U11918 ( .A1(n13897), .A2(n13778), .B1(n13775), .B2(n13732), .ZN(
        n14656) );
  NOR2_X1 U11919 ( .A1(n9457), .A2(P1_U3086), .ZN(n12381) );
  AND2_X1 U11920 ( .A1(n12381), .A2(n9458), .ZN(n14124) );
  AND2_X1 U11921 ( .A1(n14124), .A2(n14123), .ZN(n10294) );
  INV_X1 U11922 ( .A(n14537), .ZN(n13715) );
  OAI22_X1 U11923 ( .A1(n13753), .A2(n14714), .B1(n14656), .B2(n13715), .ZN(
        n9459) );
  OR3_X1 U11924 ( .A1(n9461), .A2(n9460), .A3(n9459), .ZN(P1_U3218) );
  NOR2_X1 U11925 ( .A1(n9473), .A2(P3_STATE_REG_SCAN_IN), .ZN(n14381) );
  INV_X1 U11926 ( .A(n14381), .ZN(n14370) );
  INV_X1 U11927 ( .A(SI_3_), .ZN(n9462) );
  OAI222_X1 U11928 ( .A1(P3_U3151), .A2(n7282), .B1(n14370), .B2(n9463), .C1(
        n9462), .C2(n14368), .ZN(P3_U3292) );
  INV_X1 U11929 ( .A(n9464), .ZN(n9465) );
  OAI222_X1 U11930 ( .A1(P3_U3151), .A2(n6532), .B1(n14368), .B2(n9466), .C1(
        n14370), .C2(n9465), .ZN(P3_U3294) );
  INV_X1 U11931 ( .A(SI_7_), .ZN(n9468) );
  OAI222_X1 U11932 ( .A1(P3_U3151), .A2(n10081), .B1(n14368), .B2(n9468), .C1(
        n14370), .C2(n9467), .ZN(P3_U3288) );
  INV_X1 U11933 ( .A(n14368), .ZN(n14380) );
  AOI22_X1 U11934 ( .A1(n14966), .A2(P3_STATE_REG_SCAN_IN), .B1(SI_5_), .B2(
        n14380), .ZN(n9469) );
  OAI21_X1 U11935 ( .B1(n9470), .B2(n14370), .A(n9469), .ZN(P3_U3290) );
  INV_X1 U11936 ( .A(SI_9_), .ZN(n9472) );
  OAI222_X1 U11937 ( .A1(P3_U3151), .A2(n11090), .B1(n14368), .B2(n9472), .C1(
        n14370), .C2(n9471), .ZN(P3_U3286) );
  NAND2_X1 U11938 ( .A1(n7626), .A2(P2_U3088), .ZN(n13594) );
  AND2_X1 U11939 ( .A1(n9473), .A2(P2_U3088), .ZN(n13583) );
  INV_X2 U11940 ( .A(n13583), .ZN(n13596) );
  OAI222_X1 U11941 ( .A1(n13594), .A2(n9474), .B1(n13596), .B2(n9478), .C1(
        P2_U3088), .C2(n14791), .ZN(P2_U3326) );
  AND2_X1 U11942 ( .A1(n7626), .A2(P1_U3086), .ZN(n11325) );
  INV_X2 U11943 ( .A(n11325), .ZN(n11860) );
  OAI222_X1 U11944 ( .A1(n9625), .A2(P1_U3086), .B1(n11860), .B2(n9487), .C1(
        n9476), .C2(n14247), .ZN(P1_U3352) );
  OAI222_X1 U11945 ( .A1(n9652), .A2(P1_U3086), .B1(n11860), .B2(n9478), .C1(
        n9477), .C2(n14247), .ZN(P1_U3354) );
  OR2_X1 U11946 ( .A1(n9479), .A2(n9318), .ZN(n9480) );
  XNOR2_X1 U11947 ( .A(n9480), .B(P1_IR_REG_5__SCAN_IN), .ZN(n10387) );
  INV_X1 U11948 ( .A(n10387), .ZN(n9692) );
  INV_X1 U11949 ( .A(n10389), .ZN(n9485) );
  INV_X1 U11950 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n9481) );
  OAI222_X1 U11951 ( .A1(n9692), .A2(P1_U3086), .B1(n11860), .B2(n9485), .C1(
        n9481), .C2(n14247), .ZN(P1_U3350) );
  OAI222_X1 U11952 ( .A1(P3_U3151), .A2(n11131), .B1(n14368), .B2(n9483), .C1(
        n14370), .C2(n9482), .ZN(P3_U3284) );
  INV_X1 U11953 ( .A(n13594), .ZN(n13590) );
  AOI22_X1 U11954 ( .A1(n9667), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_5__SCAN_IN), .B2(n13590), .ZN(n9484) );
  OAI21_X1 U11955 ( .B1(n9485), .B2(n13596), .A(n9484), .ZN(P2_U3322) );
  AOI22_X1 U11956 ( .A1(n13184), .A2(P2_STATE_REG_SCAN_IN), .B1(n13590), .B2(
        P1_DATAO_REG_3__SCAN_IN), .ZN(n9486) );
  OAI21_X1 U11957 ( .B1(n9487), .B2(n13596), .A(n9486), .ZN(P2_U3324) );
  NAND2_X1 U11958 ( .A1(n9479), .A2(n9488), .ZN(n9490) );
  NAND2_X1 U11959 ( .A1(n9490), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9489) );
  MUX2_X1 U11960 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9489), .S(
        P1_IR_REG_6__SCAN_IN), .Z(n9491) );
  AND2_X1 U11961 ( .A1(n9491), .A2(n9954), .ZN(n10401) );
  INV_X1 U11962 ( .A(n10401), .ZN(n9710) );
  INV_X1 U11963 ( .A(n10400), .ZN(n9495) );
  OAI222_X1 U11964 ( .A1(n9710), .A2(P1_U3086), .B1(n11860), .B2(n9495), .C1(
        n9492), .C2(n14247), .ZN(P1_U3349) );
  INV_X1 U11965 ( .A(n13590), .ZN(n13588) );
  OAI222_X1 U11966 ( .A1(n13588), .A2(n9493), .B1(n13596), .B2(n9503), .C1(
        P2_U3088), .C2(n13162), .ZN(P2_U3325) );
  OAI222_X1 U11967 ( .A1(n13588), .A2(n9494), .B1(n13596), .B2(n10303), .C1(
        P2_U3088), .C2(n9579), .ZN(P2_U3323) );
  INV_X1 U11968 ( .A(n9884), .ZN(n9558) );
  OAI222_X1 U11969 ( .A1(n13588), .A2(n9496), .B1(n13596), .B2(n9495), .C1(
        P2_U3088), .C2(n9558), .ZN(P2_U3321) );
  NAND2_X1 U11970 ( .A1(n9497), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9499) );
  INV_X1 U11971 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n9498) );
  XNOR2_X1 U11972 ( .A(n9499), .B(n9498), .ZN(n10306) );
  OAI222_X1 U11973 ( .A1(n14247), .A2(n10302), .B1(n11860), .B2(n10303), .C1(
        n10306), .C2(P1_U3086), .ZN(P1_U3351) );
  INV_X1 U11974 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n9501) );
  INV_X1 U11975 ( .A(n10678), .ZN(n9506) );
  INV_X1 U11976 ( .A(n14806), .ZN(n9500) );
  OAI222_X1 U11977 ( .A1(n13588), .A2(n9501), .B1(n13596), .B2(n9506), .C1(
        P2_U3088), .C2(n9500), .ZN(P2_U3320) );
  OAI222_X1 U11978 ( .A1(n9909), .A2(P1_U3086), .B1(n11860), .B2(n9503), .C1(
        n9502), .C2(n14247), .ZN(P1_U3353) );
  NAND2_X1 U11979 ( .A1(n9954), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9504) );
  XNOR2_X1 U11980 ( .A(n9504), .B(P1_IR_REG_7__SCAN_IN), .ZN(n10679) );
  INV_X1 U11981 ( .A(n10679), .ZN(n9717) );
  OAI222_X1 U11982 ( .A1(n9717), .A2(P1_U3086), .B1(n11860), .B2(n9506), .C1(
        n9505), .C2(n14247), .ZN(P1_U3348) );
  INV_X1 U11983 ( .A(n9507), .ZN(n9508) );
  OAI222_X1 U11984 ( .A1(n12564), .A2(P3_U3151), .B1(n14370), .B2(n9508), .C1(
        n15403), .C2(n14368), .ZN(P3_U3283) );
  NAND2_X1 U11985 ( .A1(n9586), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9522) );
  XNOR2_X1 U11986 ( .A(n9522), .B(n6751), .ZN(n10685) );
  INV_X1 U11987 ( .A(n10685), .ZN(n9833) );
  INV_X1 U11988 ( .A(n10684), .ZN(n9511) );
  OAI222_X1 U11989 ( .A1(n9833), .A2(P1_U3086), .B1(n11860), .B2(n9511), .C1(
        n9509), .C2(n14247), .ZN(P1_U3347) );
  INV_X1 U11990 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n9512) );
  INV_X1 U11991 ( .A(n14819), .ZN(n9510) );
  OAI222_X1 U11992 ( .A1(n13588), .A2(n9512), .B1(n13596), .B2(n9511), .C1(
        P2_U3088), .C2(n9510), .ZN(P2_U3319) );
  OR2_X1 U11993 ( .A1(n9513), .A2(n9595), .ZN(n14685) );
  INV_X1 U11994 ( .A(n9514), .ZN(n9515) );
  AOI22_X1 U11995 ( .A1(n14685), .A2(n9420), .B1(n9515), .B2(n9516), .ZN(
        P1_U3445) );
  AOI22_X1 U11996 ( .A1(n14685), .A2(n9518), .B1(n9517), .B2(n9516), .ZN(
        P1_U3446) );
  INV_X1 U11997 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n9520) );
  INV_X1 U11998 ( .A(n10871), .ZN(n9524) );
  INV_X1 U11999 ( .A(n10168), .ZN(n9519) );
  OAI222_X1 U12000 ( .A1(n13588), .A2(n9520), .B1(n13596), .B2(n9524), .C1(
        P2_U3088), .C2(n9519), .ZN(P2_U3318) );
  INV_X1 U12001 ( .A(n6751), .ZN(n9521) );
  NAND2_X1 U12002 ( .A1(n9522), .A2(n9521), .ZN(n9523) );
  NAND2_X1 U12003 ( .A1(n9523), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9619) );
  XNOR2_X1 U12004 ( .A(n9619), .B(P1_IR_REG_9__SCAN_IN), .ZN(n10872) );
  INV_X1 U12005 ( .A(n10872), .ZN(n9841) );
  OAI222_X1 U12006 ( .A1(n14247), .A2(n15379), .B1(n11860), .B2(n9524), .C1(
        n9841), .C2(P1_U3086), .ZN(P1_U3346) );
  INV_X1 U12007 ( .A(n11891), .ZN(n9525) );
  INV_X1 U12008 ( .A(P3_D_REG_21__SCAN_IN), .ZN(n15167) );
  NOR2_X1 U12009 ( .A1(n9525), .A2(n15167), .ZN(P3_U3244) );
  INV_X1 U12010 ( .A(P3_D_REG_12__SCAN_IN), .ZN(n15207) );
  NOR2_X1 U12011 ( .A1(n9525), .A2(n15207), .ZN(P3_U3253) );
  INV_X1 U12012 ( .A(P3_D_REG_26__SCAN_IN), .ZN(n15281) );
  NOR2_X1 U12013 ( .A1(n9525), .A2(n15281), .ZN(P3_U3239) );
  INV_X1 U12014 ( .A(P3_D_REG_19__SCAN_IN), .ZN(n15155) );
  NOR2_X1 U12015 ( .A1(n9525), .A2(n15155), .ZN(P3_U3246) );
  INV_X1 U12016 ( .A(P3_D_REG_10__SCAN_IN), .ZN(n15261) );
  NOR2_X1 U12017 ( .A1(n9525), .A2(n15261), .ZN(P3_U3255) );
  INV_X1 U12018 ( .A(P3_D_REG_2__SCAN_IN), .ZN(n15396) );
  NOR2_X1 U12019 ( .A1(n9525), .A2(n15396), .ZN(P3_U3263) );
  INV_X1 U12020 ( .A(P3_D_REG_14__SCAN_IN), .ZN(n15136) );
  NOR2_X1 U12021 ( .A1(n9525), .A2(n15136), .ZN(P3_U3251) );
  OAI222_X1 U12022 ( .A1(P3_U3151), .A2(n12582), .B1(n14368), .B2(n9527), .C1(
        n14370), .C2(n9526), .ZN(P3_U3282) );
  MUX2_X1 U12023 ( .A(n9528), .B(P2_REG2_REG_1__SCAN_IN), .S(n14791), .Z(
        n14796) );
  NAND3_X1 U12024 ( .A1(n14796), .A2(P2_REG2_REG_0__SCAN_IN), .A3(n15330), 
        .ZN(n14795) );
  INV_X1 U12025 ( .A(n14791), .ZN(n9529) );
  NAND2_X1 U12026 ( .A1(n9529), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n13168) );
  INV_X1 U12027 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n15291) );
  AOI21_X1 U12028 ( .B1(n14795), .B2(n13168), .A(n13169), .ZN(n13167) );
  NOR2_X1 U12029 ( .A1(n13162), .A2(n15291), .ZN(n13178) );
  INV_X1 U12030 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n9530) );
  MUX2_X1 U12031 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n9530), .S(n13184), .Z(n9531) );
  NAND2_X1 U12032 ( .A1(n13184), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n9576) );
  MUX2_X1 U12033 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n10567), .S(n9579), .Z(n9575) );
  NOR2_X1 U12034 ( .A1(n9579), .A2(n10567), .ZN(n9660) );
  MUX2_X1 U12035 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n9532), .S(n9667), .Z(n9659)
         );
  NAND2_X1 U12036 ( .A1(n9667), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n9534) );
  MUX2_X1 U12037 ( .A(n10517), .B(P2_REG2_REG_6__SCAN_IN), .S(n9884), .Z(n9533) );
  AOI21_X1 U12038 ( .B1(n9658), .B2(n9534), .A(n9533), .ZN(n9883) );
  NAND3_X1 U12039 ( .A1(n9658), .A2(n9534), .A3(n9533), .ZN(n9543) );
  OAI21_X1 U12040 ( .B1(n9961), .B2(n9536), .A(n9535), .ZN(n9539) );
  INV_X1 U12041 ( .A(n9537), .ZN(n9538) );
  AND2_X1 U12042 ( .A1(n9539), .A2(n9538), .ZN(n9555) );
  INV_X1 U12043 ( .A(n9555), .ZN(n9557) );
  OR2_X1 U12044 ( .A1(n8278), .A2(P2_U3088), .ZN(n13585) );
  INV_X1 U12045 ( .A(n13585), .ZN(n9540) );
  NAND2_X1 U12046 ( .A1(n9557), .A2(n9540), .ZN(n9551) );
  INV_X1 U12047 ( .A(n9551), .ZN(n9542) );
  INV_X1 U12048 ( .A(n9541), .ZN(n9550) );
  NAND2_X1 U12049 ( .A1(n9543), .A2(n14870), .ZN(n9563) );
  NAND2_X1 U12050 ( .A1(n15330), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n15358) );
  NAND2_X1 U12051 ( .A1(n13166), .A2(n13165), .ZN(n13164) );
  OAI21_X1 U12052 ( .B1(n9545), .B2(n13162), .A(n13164), .ZN(n13176) );
  MUX2_X1 U12053 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n7784), .S(n13184), .Z(
        n13177) );
  INV_X1 U12054 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n9546) );
  MUX2_X1 U12055 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n9546), .S(n9579), .Z(n9573)
         );
  NOR2_X1 U12056 ( .A1(n9574), .A2(n9573), .ZN(n9572) );
  AOI21_X1 U12057 ( .B1(n9547), .B2(P2_REG1_REG_4__SCAN_IN), .A(n9572), .ZN(
        n9657) );
  INV_X1 U12058 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n9548) );
  MUX2_X1 U12059 ( .A(n9548), .B(P2_REG1_REG_5__SCAN_IN), .S(n9667), .Z(n9656)
         );
  AOI21_X1 U12060 ( .B1(P2_REG1_REG_5__SCAN_IN), .B2(n9667), .A(n9655), .ZN(
        n9553) );
  INV_X1 U12061 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n9549) );
  MUX2_X1 U12062 ( .A(n9549), .B(P2_REG1_REG_6__SCAN_IN), .S(n9884), .Z(n9552)
         );
  NOR2_X1 U12063 ( .A1(n9553), .A2(n9552), .ZN(n9876) );
  AOI211_X1 U12064 ( .C1(n9553), .C2(n9552), .A(n14863), .B(n9876), .ZN(n9554)
         );
  INV_X1 U12065 ( .A(n9554), .ZN(n9562) );
  AND2_X1 U12066 ( .A1(n9555), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14789) );
  NAND2_X1 U12067 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3088), .ZN(n10264) );
  INV_X1 U12068 ( .A(n10264), .ZN(n9560) );
  AND2_X1 U12069 ( .A1(n8278), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9556) );
  NAND2_X1 U12070 ( .A1(n9557), .A2(n9556), .ZN(n14834) );
  NOR2_X1 U12071 ( .A1(n14834), .A2(n9558), .ZN(n9559) );
  AOI211_X1 U12072 ( .C1(P2_ADDR_REG_6__SCAN_IN), .C2(n14789), .A(n9560), .B(
        n9559), .ZN(n9561) );
  OAI211_X1 U12073 ( .C1(n9883), .C2(n9563), .A(n9562), .B(n9561), .ZN(
        P2_U3220) );
  OAI22_X1 U12074 ( .A1(n14836), .A2(n9565), .B1(n9564), .B2(n14863), .ZN(
        n9568) );
  NAND2_X1 U12075 ( .A1(n14870), .A2(n9565), .ZN(n9566) );
  OAI211_X1 U12076 ( .C1(P2_REG1_REG_0__SCAN_IN), .C2(n14863), .A(n9566), .B(
        n14834), .ZN(n9567) );
  MUX2_X1 U12077 ( .A(n9568), .B(n9567), .S(n15330), .Z(n9571) );
  INV_X1 U12078 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n9569) );
  OAI22_X1 U12079 ( .A1(n14874), .A2(n9569), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7761), .ZN(n9570) );
  OR2_X1 U12080 ( .A1(n9571), .A2(n9570), .ZN(P2_U3214) );
  AOI211_X1 U12081 ( .C1(n9574), .C2(n9573), .A(n14863), .B(n9572), .ZN(n9582)
         );
  AND3_X1 U12082 ( .A1(n13183), .A2(n9576), .A3(n9575), .ZN(n9577) );
  NOR3_X1 U12083 ( .A1(n14836), .A2(n9661), .A3(n9577), .ZN(n9581) );
  NAND2_X1 U12084 ( .A1(n14789), .A2(P2_ADDR_REG_4__SCAN_IN), .ZN(n9578) );
  NAND2_X1 U12085 ( .A1(P2_U3088), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n11881) );
  OAI211_X1 U12086 ( .C1(n14834), .C2(n9579), .A(n9578), .B(n11881), .ZN(n9580) );
  OR3_X1 U12087 ( .A1(n9582), .A2(n9581), .A3(n9580), .ZN(P2_U3218) );
  INV_X1 U12088 ( .A(n11193), .ZN(n9590) );
  INV_X1 U12089 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n9583) );
  NAND2_X1 U12090 ( .A1(n9584), .A2(n9583), .ZN(n9585) );
  INV_X1 U12091 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n9587) );
  NAND2_X1 U12092 ( .A1(n9693), .A2(n9587), .ZN(n9696) );
  NAND2_X1 U12093 ( .A1(n9696), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9588) );
  XNOR2_X1 U12094 ( .A(n9588), .B(P1_IR_REG_12__SCAN_IN), .ZN(n11194) );
  INV_X1 U12095 ( .A(n11194), .ZN(n10323) );
  OAI222_X1 U12096 ( .A1(n14247), .A2(n9589), .B1(n11860), .B2(n9590), .C1(
        n10323), .C2(P1_U3086), .ZN(P1_U3343) );
  INV_X1 U12097 ( .A(n14855), .ZN(n14849) );
  OAI222_X1 U12098 ( .A1(n13594), .A2(n9591), .B1(n13596), .B2(n9590), .C1(
        P2_U3088), .C2(n14849), .ZN(P2_U3315) );
  INV_X1 U12099 ( .A(n9592), .ZN(n9594) );
  OR2_X1 U12100 ( .A1(n12146), .A2(n9594), .ZN(n9593) );
  AND2_X1 U12101 ( .A1(n11572), .A2(n9593), .ZN(n9611) );
  NAND2_X1 U12102 ( .A1(n9594), .A2(P1_STATE_REG_SCAN_IN), .ZN(n12384) );
  NAND2_X1 U12103 ( .A1(n9595), .A2(n12384), .ZN(n9612) );
  NAND2_X1 U12104 ( .A1(n9611), .A2(n9612), .ZN(n14606) );
  INV_X1 U12105 ( .A(n9909), .ZN(n9598) );
  INV_X1 U12106 ( .A(n9652), .ZN(n9604) );
  NOR3_X1 U12107 ( .A1(n9643), .A2(n9387), .A3(n14602), .ZN(n9642) );
  MUX2_X1 U12108 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n9597), .S(n9909), .Z(n9905)
         );
  NOR2_X1 U12109 ( .A1(n9906), .A2(n9905), .ZN(n9904) );
  XOR2_X1 U12110 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n9625), .Z(n9600) );
  NOR2_X1 U12111 ( .A1(n9601), .A2(n9600), .ZN(n9626) );
  INV_X1 U12112 ( .A(n13875), .ZN(n14601) );
  AOI211_X1 U12113 ( .C1(n9601), .C2(n9600), .A(n9626), .B(n13847), .ZN(n9610)
         );
  OR2_X1 U12114 ( .A1(n9450), .A2(n13875), .ZN(n9602) );
  MUX2_X1 U12115 ( .A(P1_REG2_REG_1__SCAN_IN), .B(n9358), .S(n9652), .Z(n9646)
         );
  NOR3_X1 U12116 ( .A1(n9646), .A2(n14602), .A3(n9603), .ZN(n9645) );
  AOI21_X1 U12117 ( .B1(n9604), .B2(P1_REG2_REG_1__SCAN_IN), .A(n9645), .ZN(
        n9903) );
  MUX2_X1 U12118 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n9397), .S(n9909), .Z(n9902)
         );
  NOR2_X1 U12119 ( .A1(n9903), .A2(n9902), .ZN(n9901) );
  NOR2_X1 U12120 ( .A1(n9909), .A2(n9397), .ZN(n9606) );
  MUX2_X1 U12121 ( .A(n14660), .B(P1_REG2_REG_3__SCAN_IN), .S(n9625), .Z(n9605) );
  OAI21_X1 U12122 ( .B1(n9901), .B2(n9606), .A(n9605), .ZN(n9918) );
  INV_X1 U12123 ( .A(n9918), .ZN(n9608) );
  NOR3_X1 U12124 ( .A1(n9901), .A2(n9606), .A3(n9605), .ZN(n9607) );
  NOR3_X1 U12125 ( .A1(n14619), .A2(n9608), .A3(n9607), .ZN(n9609) );
  NOR2_X1 U12126 ( .A1(n9610), .A2(n9609), .ZN(n9615) );
  INV_X1 U12127 ( .A(n9611), .ZN(n9613) );
  AND2_X1 U12128 ( .A1(n9613), .A2(n9612), .ZN(n14604) );
  AOI22_X1 U12129 ( .A1(n14604), .A2(P1_ADDR_REG_3__SCAN_IN), .B1(
        P1_REG3_REG_3__SCAN_IN), .B2(P1_U3086), .ZN(n9614) );
  OAI211_X1 U12130 ( .C1(n9625), .C2(n13862), .A(n9615), .B(n9614), .ZN(
        P1_U3246) );
  INV_X1 U12131 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n9617) );
  INV_X1 U12132 ( .A(n10998), .ZN(n9622) );
  INV_X1 U12133 ( .A(n11026), .ZN(n9616) );
  OAI222_X1 U12134 ( .A1(n13588), .A2(n9617), .B1(n13596), .B2(n9622), .C1(
        P2_U3088), .C2(n9616), .ZN(P2_U3317) );
  INV_X1 U12135 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n9618) );
  NAND2_X1 U12136 ( .A1(n9619), .A2(n9618), .ZN(n9620) );
  NAND2_X1 U12137 ( .A1(n9620), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9621) );
  XNOR2_X1 U12138 ( .A(n9621), .B(P1_IR_REG_10__SCAN_IN), .ZN(n10999) );
  INV_X1 U12139 ( .A(n10999), .ZN(n10024) );
  OAI222_X1 U12140 ( .A1(n14247), .A2(n9623), .B1(n11860), .B2(n9622), .C1(
        n10024), .C2(P1_U3086), .ZN(P1_U3345) );
  INV_X1 U12141 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n9624) );
  MUX2_X1 U12142 ( .A(n9624), .B(P1_REG1_REG_6__SCAN_IN), .S(n10401), .Z(n9629) );
  INV_X1 U12143 ( .A(n10306), .ZN(n9627) );
  INV_X1 U12144 ( .A(n9625), .ZN(n9630) );
  XOR2_X1 U12145 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n10306), .Z(n9914) );
  NOR2_X1 U12146 ( .A1(n9915), .A2(n9914), .ZN(n9913) );
  INV_X1 U12147 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n9754) );
  MUX2_X1 U12148 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n9754), .S(n10387), .Z(n9680) );
  NAND2_X1 U12149 ( .A1(n9681), .A2(n9680), .ZN(n9679) );
  OAI21_X1 U12150 ( .B1(n10387), .B2(P1_REG1_REG_5__SCAN_IN), .A(n9679), .ZN(
        n9628) );
  NOR2_X1 U12151 ( .A1(n9628), .A2(n9629), .ZN(n9706) );
  AOI211_X1 U12152 ( .C1(n9629), .C2(n9628), .A(n13847), .B(n9706), .ZN(n9635)
         );
  NAND2_X1 U12153 ( .A1(n9630), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n9917) );
  MUX2_X1 U12154 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n10313), .S(n10306), .Z(
        n9916) );
  AOI21_X1 U12155 ( .B1(n9918), .B2(n9917), .A(n9916), .ZN(n9920) );
  NOR2_X1 U12156 ( .A1(n10306), .A2(n10313), .ZN(n9684) );
  INV_X1 U12157 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n9758) );
  MUX2_X1 U12158 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n9758), .S(n10387), .Z(n9683) );
  OAI21_X1 U12159 ( .B1(n9920), .B2(n9684), .A(n9683), .ZN(n9682) );
  NAND2_X1 U12160 ( .A1(n10387), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n9632) );
  INV_X1 U12161 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n9709) );
  MUX2_X1 U12162 ( .A(n9709), .B(P1_REG2_REG_6__SCAN_IN), .S(n10401), .Z(n9631) );
  AOI21_X1 U12163 ( .B1(n9682), .B2(n9632), .A(n9631), .ZN(n9713) );
  AND3_X1 U12164 ( .A1(n9682), .A2(n9632), .A3(n9631), .ZN(n9633) );
  NOR3_X1 U12165 ( .A1(n9713), .A2(n14619), .A3(n9633), .ZN(n9634) );
  NOR2_X1 U12166 ( .A1(n9635), .A2(n9634), .ZN(n9638) );
  AND2_X1 U12167 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n9636) );
  AOI21_X1 U12168 ( .B1(n14604), .B2(P1_ADDR_REG_6__SCAN_IN), .A(n9636), .ZN(
        n9637) );
  OAI211_X1 U12169 ( .C1(n9710), .C2(n13862), .A(n9638), .B(n9637), .ZN(
        P1_U3249) );
  CLKBUF_X2 U12170 ( .A(P1_U4016), .Z(n13777) );
  NOR2_X1 U12171 ( .A1(n14604), .A2(n13777), .ZN(P1_U3085) );
  INV_X1 U12172 ( .A(P3_DATAO_REG_6__SCAN_IN), .ZN(n15237) );
  NAND2_X1 U12173 ( .A1(n15036), .A2(P3_U3897), .ZN(n9639) );
  OAI21_X1 U12174 ( .B1(P3_U3897), .B2(n15237), .A(n9639), .ZN(P3_U3497) );
  INV_X1 U12175 ( .A(P3_DATAO_REG_4__SCAN_IN), .ZN(n15306) );
  NAND2_X1 U12176 ( .A1(n15037), .A2(P3_U3897), .ZN(n9640) );
  OAI21_X1 U12177 ( .B1(P3_U3897), .B2(n15306), .A(n9640), .ZN(P3_U3495) );
  INV_X1 U12178 ( .A(P3_DATAO_REG_12__SCAN_IN), .ZN(n15244) );
  NAND2_X1 U12179 ( .A1(n14428), .A2(P3_U3897), .ZN(n9641) );
  OAI21_X1 U12180 ( .B1(P3_U3897), .B2(n15244), .A(n9641), .ZN(P3_U3503) );
  NAND2_X1 U12181 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n9644) );
  AOI211_X1 U12182 ( .C1(n9644), .C2(n9643), .A(n9642), .B(n13847), .ZN(n9649)
         );
  NOR2_X1 U12183 ( .A1(n14602), .A2(n9603), .ZN(n9897) );
  INV_X1 U12184 ( .A(n9897), .ZN(n9647) );
  AOI211_X1 U12185 ( .C1(n9647), .C2(n9646), .A(n9645), .B(n14619), .ZN(n9648)
         );
  NOR2_X1 U12186 ( .A1(n9649), .A2(n9648), .ZN(n9651) );
  AOI22_X1 U12187 ( .A1(n14604), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n9650) );
  OAI211_X1 U12188 ( .C1(n9652), .C2(n13862), .A(n9651), .B(n9650), .ZN(
        P1_U3244) );
  INV_X1 U12189 ( .A(P3_DATAO_REG_1__SCAN_IN), .ZN(n9654) );
  NAND2_X1 U12190 ( .A1(n10041), .A2(P3_U3897), .ZN(n9653) );
  OAI21_X1 U12191 ( .B1(P3_U3897), .B2(n9654), .A(n9653), .ZN(P3_U3492) );
  INV_X1 U12192 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n9670) );
  AOI211_X1 U12193 ( .C1(n9657), .C2(n9656), .A(n14863), .B(n9655), .ZN(n9665)
         );
  INV_X1 U12194 ( .A(n9658), .ZN(n9663) );
  NOR3_X1 U12195 ( .A1(n9661), .A2(n9660), .A3(n9659), .ZN(n9662) );
  NOR3_X1 U12196 ( .A1(n9663), .A2(n14836), .A3(n9662), .ZN(n9664) );
  NOR2_X1 U12197 ( .A1(n9665), .A2(n9664), .ZN(n9669) );
  AND2_X1 U12198 ( .A1(P2_U3088), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n9666) );
  AOI21_X1 U12199 ( .B1(n14868), .B2(n9667), .A(n9666), .ZN(n9668) );
  OAI211_X1 U12200 ( .C1(n14874), .C2(n9670), .A(n9669), .B(n9668), .ZN(
        P2_U3219) );
  INV_X1 U12201 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n9671) );
  OR2_X1 U12202 ( .A1(n6540), .A2(n9671), .ZN(n9675) );
  INV_X1 U12203 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n13874) );
  OR2_X1 U12204 ( .A1(n6526), .A2(n13874), .ZN(n9674) );
  INV_X1 U12205 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n9672) );
  OR2_X1 U12206 ( .A1(n11784), .A2(n9672), .ZN(n9673) );
  AND3_X1 U12207 ( .A1(n9675), .A2(n9674), .A3(n9673), .ZN(n13877) );
  NAND2_X1 U12208 ( .A1(n12371), .A2(P1_U4016), .ZN(n9676) );
  OAI21_X1 U12209 ( .B1(n13777), .B2(n13577), .A(n9676), .ZN(P1_U3591) );
  INV_X1 U12210 ( .A(n11198), .ZN(n9702) );
  NAND2_X1 U12211 ( .A1(n9846), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9677) );
  XNOR2_X1 U12212 ( .A(n9677), .B(n6756), .ZN(n13789) );
  INV_X1 U12213 ( .A(n14247), .ZN(n14244) );
  AOI22_X1 U12214 ( .A1(n13789), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n14244), .ZN(n9678) );
  OAI21_X1 U12215 ( .B1(n9702), .B2(n11860), .A(n9678), .ZN(P1_U3342) );
  OAI21_X1 U12216 ( .B1(n9681), .B2(n9680), .A(n9679), .ZN(n9688) );
  INV_X1 U12217 ( .A(n13847), .ZN(n14614) );
  INV_X1 U12218 ( .A(n9682), .ZN(n9686) );
  NOR3_X1 U12219 ( .A1(n9920), .A2(n9684), .A3(n9683), .ZN(n9685) );
  NOR3_X1 U12220 ( .A1(n14619), .A2(n9686), .A3(n9685), .ZN(n9687) );
  AOI21_X1 U12221 ( .B1(n9688), .B2(n14614), .A(n9687), .ZN(n9691) );
  NAND2_X1 U12222 ( .A1(P1_U3086), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n10460) );
  INV_X1 U12223 ( .A(n10460), .ZN(n9689) );
  AOI21_X1 U12224 ( .B1(n14604), .B2(P1_ADDR_REG_5__SCAN_IN), .A(n9689), .ZN(
        n9690) );
  OAI211_X1 U12225 ( .C1(n9692), .C2(n13862), .A(n9691), .B(n9690), .ZN(
        P1_U3248) );
  INV_X1 U12226 ( .A(n9693), .ZN(n9694) );
  NAND2_X1 U12227 ( .A1(n9694), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9695) );
  MUX2_X1 U12228 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9695), .S(
        P1_IR_REG_11__SCAN_IN), .Z(n9697) );
  INV_X1 U12229 ( .A(n11049), .ZN(n10322) );
  INV_X1 U12230 ( .A(n11048), .ZN(n9699) );
  INV_X1 U12231 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n9698) );
  OAI222_X1 U12232 ( .A1(n10322), .A2(P1_U3086), .B1(n11860), .B2(n9699), .C1(
        n9698), .C2(n14247), .ZN(P1_U3344) );
  INV_X1 U12233 ( .A(n11027), .ZN(n14835) );
  OAI222_X1 U12234 ( .A1(n13594), .A2(n9700), .B1(n13596), .B2(n9699), .C1(
        P2_U3088), .C2(n14835), .ZN(P2_U3316) );
  INV_X1 U12235 ( .A(n11165), .ZN(n11031) );
  OAI222_X1 U12236 ( .A1(P2_U3088), .A2(n11031), .B1(n13596), .B2(n9702), .C1(
        n9701), .C2(n13588), .ZN(P2_U3314) );
  INV_X1 U12237 ( .A(n9703), .ZN(n9704) );
  OAI222_X1 U12238 ( .A1(P3_U3151), .A2(n6749), .B1(n14368), .B2(n9705), .C1(
        n14370), .C2(n9704), .ZN(P3_U3280) );
  INV_X1 U12239 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n10409) );
  MUX2_X1 U12240 ( .A(n10409), .B(P1_REG1_REG_7__SCAN_IN), .S(n10679), .Z(
        n9707) );
  NOR2_X1 U12241 ( .A1(n9708), .A2(n9707), .ZN(n9821) );
  AOI211_X1 U12242 ( .C1(n9708), .C2(n9707), .A(n13847), .B(n9821), .ZN(n9720)
         );
  NOR2_X1 U12243 ( .A1(n9710), .A2(n9709), .ZN(n9712) );
  INV_X1 U12244 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n10405) );
  MUX2_X1 U12245 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n10405), .S(n10679), .Z(
        n9711) );
  OAI21_X1 U12246 ( .B1(n9713), .B2(n9712), .A(n9711), .ZN(n9819) );
  INV_X1 U12247 ( .A(n9819), .ZN(n9715) );
  NOR3_X1 U12248 ( .A1(n9713), .A2(n9712), .A3(n9711), .ZN(n9714) );
  NOR3_X1 U12249 ( .A1(n9715), .A2(n9714), .A3(n14619), .ZN(n9719) );
  NAND2_X1 U12250 ( .A1(n14604), .A2(P1_ADDR_REG_7__SCAN_IN), .ZN(n9716) );
  NAND2_X1 U12251 ( .A1(P1_U3086), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n10955) );
  OAI211_X1 U12252 ( .C1(n13862), .C2(n9717), .A(n9716), .B(n10955), .ZN(n9718) );
  OR3_X1 U12253 ( .A1(n9720), .A2(n9719), .A3(n9718), .ZN(P1_U3250) );
  INV_X1 U12254 ( .A(n15015), .ZN(n14948) );
  INV_X1 U12255 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n9873) );
  INV_X1 U12256 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n9945) );
  MUX2_X1 U12257 ( .A(n9873), .B(n9945), .S(n12670), .Z(n14932) );
  AND2_X1 U12258 ( .A1(n14932), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n14935) );
  MUX2_X1 U12259 ( .A(P3_REG2_REG_1__SCAN_IN), .B(P3_REG1_REG_1__SCAN_IN), .S(
        n9721), .Z(n9766) );
  INV_X1 U12260 ( .A(n6532), .ZN(n9767) );
  XNOR2_X1 U12261 ( .A(n9766), .B(n9767), .ZN(n9765) );
  XOR2_X1 U12262 ( .A(n14935), .B(n9765), .Z(n9745) );
  NAND2_X1 U12263 ( .A1(n9722), .A2(n12116), .ZN(n9738) );
  NAND2_X1 U12264 ( .A1(n6529), .A2(n9723), .ZN(n9725) );
  NAND2_X1 U12265 ( .A1(n9725), .A2(n9724), .ZN(n9737) );
  INV_X1 U12266 ( .A(n9737), .ZN(n9726) );
  INV_X1 U12267 ( .A(n9729), .ZN(n9731) );
  INV_X1 U12268 ( .A(n9116), .ZN(n12111) );
  MUX2_X1 U12269 ( .A(n9731), .B(n12548), .S(n12111), .Z(n12701) );
  NOR2_X1 U12270 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(n9945), .ZN(n9728) );
  NOR3_X1 U12271 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), .A3(
        n9945), .ZN(n9790) );
  INV_X1 U12272 ( .A(n9790), .ZN(n9727) );
  OAI21_X1 U12273 ( .B1(n6532), .B2(n9728), .A(n9727), .ZN(n9788) );
  XNOR2_X1 U12274 ( .A(n9788), .B(P3_REG1_REG_1__SCAN_IN), .ZN(n9742) );
  NAND2_X1 U12275 ( .A1(n9729), .A2(n12670), .ZN(n15018) );
  INV_X1 U12276 ( .A(n15023), .ZN(n9736) );
  NOR2_X1 U12277 ( .A1(n9873), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n9733) );
  INV_X1 U12278 ( .A(n9781), .ZN(n9732) );
  OAI21_X1 U12279 ( .B1(n6532), .B2(n9733), .A(n9732), .ZN(n9779) );
  INV_X1 U12280 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n10159) );
  XNOR2_X1 U12281 ( .A(n9779), .B(n10159), .ZN(n9735) );
  NAND2_X1 U12282 ( .A1(n9736), .A2(n9735), .ZN(n9741) );
  INV_X1 U12283 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n10158) );
  NOR2_X1 U12284 ( .A1(n10158), .A2(P3_STATE_REG_SCAN_IN), .ZN(n9739) );
  AOI21_X1 U12285 ( .B1(n15001), .B2(P3_ADDR_REG_1__SCAN_IN), .A(n9739), .ZN(
        n9740) );
  OAI211_X1 U12286 ( .C1(n9742), .C2(n15018), .A(n9741), .B(n9740), .ZN(n9743)
         );
  AOI21_X1 U12287 ( .B1(n9767), .B2(n15013), .A(n9743), .ZN(n9744) );
  OAI21_X1 U12288 ( .B1(n14948), .B2(n9745), .A(n9744), .ZN(P3_U3183) );
  NAND2_X1 U12289 ( .A1(n11783), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n9752) );
  INV_X1 U12290 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n9746) );
  OR2_X1 U12291 ( .A1(n11784), .A2(n9746), .ZN(n9751) );
  INV_X1 U12292 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n9755) );
  NOR2_X1 U12293 ( .A1(n9756), .A2(n9755), .ZN(n10394) );
  NAND2_X1 U12294 ( .A1(n10394), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n10407) );
  NAND2_X1 U12295 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_REG3_REG_8__SCAN_IN), 
        .ZN(n9747) );
  NAND2_X1 U12296 ( .A1(n11005), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n11053) );
  INV_X1 U12297 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n11052) );
  INV_X1 U12298 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n11202) );
  OR2_X1 U12299 ( .A1(n11212), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9748) );
  NAND2_X1 U12300 ( .A1(n11503), .A2(n9748), .ZN(n14111) );
  OR2_X1 U12301 ( .A1(n11600), .A2(n14111), .ZN(n9750) );
  INV_X1 U12302 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n14112) );
  OR2_X1 U12303 ( .A1(n6526), .A2(n14112), .ZN(n9749) );
  MUX2_X1 U12304 ( .A(n9984), .B(n13663), .S(n13777), .Z(n9753) );
  INV_X1 U12305 ( .A(n9753), .ZN(P1_U3575) );
  NAND2_X1 U12306 ( .A1(n12321), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n9762) );
  OR2_X1 U12307 ( .A1(n6539), .A2(n9754), .ZN(n9761) );
  AND2_X1 U12308 ( .A1(n9756), .A2(n9755), .ZN(n9757) );
  OR2_X1 U12309 ( .A1(n9757), .A2(n10394), .ZN(n14644) );
  OR2_X1 U12310 ( .A1(n11600), .A2(n14644), .ZN(n9760) );
  OR2_X1 U12311 ( .A1(n6526), .A2(n9758), .ZN(n9759) );
  MUX2_X1 U12312 ( .A(n9763), .B(n12186), .S(n13777), .Z(n9764) );
  INV_X1 U12313 ( .A(n9764), .ZN(P1_U3565) );
  MUX2_X1 U12314 ( .A(P3_REG2_REG_4__SCAN_IN), .B(P3_REG1_REG_4__SCAN_IN), .S(
        n12670), .Z(n10055) );
  XNOR2_X1 U12315 ( .A(n10055), .B(n10056), .ZN(n10053) );
  NAND2_X1 U12316 ( .A1(n9765), .A2(n14935), .ZN(n9770) );
  INV_X1 U12317 ( .A(n9766), .ZN(n9768) );
  NAND2_X1 U12318 ( .A1(n9768), .A2(n9767), .ZN(n9769) );
  NAND2_X1 U12319 ( .A1(n9770), .A2(n9769), .ZN(n9801) );
  MUX2_X1 U12320 ( .A(P3_REG2_REG_2__SCAN_IN), .B(P3_REG1_REG_2__SCAN_IN), .S(
        n12670), .Z(n9771) );
  XNOR2_X1 U12321 ( .A(n9771), .B(n9814), .ZN(n9802) );
  NAND2_X1 U12322 ( .A1(n9801), .A2(n9802), .ZN(n9774) );
  INV_X1 U12323 ( .A(n9771), .ZN(n9772) );
  NAND2_X1 U12324 ( .A1(n9772), .A2(n9814), .ZN(n9773) );
  NAND2_X1 U12325 ( .A1(n9774), .A2(n9773), .ZN(n14946) );
  MUX2_X1 U12326 ( .A(P3_REG2_REG_3__SCAN_IN), .B(P3_REG1_REG_3__SCAN_IN), .S(
        n12670), .Z(n9775) );
  XNOR2_X1 U12327 ( .A(n9775), .B(n14952), .ZN(n14947) );
  NAND2_X1 U12328 ( .A1(n14946), .A2(n14947), .ZN(n9778) );
  INV_X1 U12329 ( .A(n9775), .ZN(n9776) );
  NAND2_X1 U12330 ( .A1(n9776), .A2(n14952), .ZN(n9777) );
  NAND2_X1 U12331 ( .A1(n9778), .A2(n9777), .ZN(n10054) );
  XOR2_X1 U12332 ( .A(n10054), .B(n10053), .Z(n9800) );
  NOR2_X1 U12333 ( .A1(n9779), .A2(n10159), .ZN(n9780) );
  INV_X1 U12334 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n10051) );
  NOR2_X1 U12335 ( .A1(n14952), .A2(n9782), .ZN(n9783) );
  INV_X1 U12336 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n14943) );
  INV_X1 U12337 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n9784) );
  AOI22_X1 U12338 ( .A1(n10056), .A2(P3_REG2_REG_4__SCAN_IN), .B1(n9784), .B2(
        n14358), .ZN(n9785) );
  AOI21_X1 U12339 ( .B1(n9786), .B2(n9785), .A(n10067), .ZN(n9787) );
  NOR2_X1 U12340 ( .A1(n15023), .A2(n9787), .ZN(n9798) );
  INV_X1 U12341 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n15111) );
  NOR2_X1 U12342 ( .A1(n9788), .A2(n15111), .ZN(n9789) );
  INV_X1 U12343 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n15113) );
  NOR2_X1 U12344 ( .A1(n14952), .A2(n9791), .ZN(n9792) );
  INV_X1 U12345 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n15115) );
  INV_X1 U12346 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n15117) );
  AOI22_X1 U12347 ( .A1(n10056), .A2(P3_REG1_REG_4__SCAN_IN), .B1(n15117), 
        .B2(n14358), .ZN(n9793) );
  AOI21_X1 U12348 ( .B1(n9794), .B2(n9793), .A(n10077), .ZN(n9796) );
  AND2_X1 U12349 ( .A1(P3_U3151), .A2(P3_REG3_REG_4__SCAN_IN), .ZN(n10114) );
  AOI21_X1 U12350 ( .B1(n15001), .B2(P3_ADDR_REG_4__SCAN_IN), .A(n10114), .ZN(
        n9795) );
  OAI21_X1 U12351 ( .B1(n15018), .B2(n9796), .A(n9795), .ZN(n9797) );
  AOI211_X1 U12352 ( .C1(n15013), .C2(n10056), .A(n9798), .B(n9797), .ZN(n9799) );
  OAI21_X1 U12353 ( .B1(n9800), .B2(n14948), .A(n9799), .ZN(P3_U3186) );
  XOR2_X1 U12354 ( .A(n9801), .B(n9802), .Z(n9816) );
  AOI21_X1 U12355 ( .B1(n9805), .B2(n9804), .A(n9803), .ZN(n9806) );
  NOR2_X1 U12356 ( .A1(n15023), .A2(n9806), .ZN(n9813) );
  AOI21_X1 U12357 ( .B1(n9809), .B2(n9808), .A(n9807), .ZN(n9811) );
  AOI22_X1 U12358 ( .A1(n15001), .A2(P3_ADDR_REG_2__SCAN_IN), .B1(
        P3_REG3_REG_2__SCAN_IN), .B2(P3_U3151), .ZN(n9810) );
  OAI21_X1 U12359 ( .B1(n9811), .B2(n15018), .A(n9810), .ZN(n9812) );
  AOI211_X1 U12360 ( .C1(n15013), .C2(n9814), .A(n9813), .B(n9812), .ZN(n9815)
         );
  OAI21_X1 U12361 ( .B1(n9816), .B2(n14948), .A(n9815), .ZN(P3_U3184) );
  NAND2_X1 U12362 ( .A1(n10679), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n9818) );
  INV_X1 U12363 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n9832) );
  MUX2_X1 U12364 ( .A(n9832), .B(P1_REG2_REG_8__SCAN_IN), .S(n10685), .Z(n9817) );
  AOI21_X1 U12365 ( .B1(n9819), .B2(n9818), .A(n9817), .ZN(n9836) );
  NAND3_X1 U12366 ( .A1(n9819), .A2(n9818), .A3(n9817), .ZN(n9820) );
  NAND2_X1 U12367 ( .A1(n9820), .A2(n13866), .ZN(n9828) );
  INV_X1 U12368 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n10688) );
  MUX2_X1 U12369 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n10688), .S(n10685), .Z(
        n9822) );
  NAND2_X1 U12370 ( .A1(n9823), .A2(n9822), .ZN(n9829) );
  OAI21_X1 U12371 ( .B1(n9823), .B2(n9822), .A(n9829), .ZN(n9824) );
  NAND2_X1 U12372 ( .A1(n9824), .A2(n14614), .ZN(n9827) );
  INV_X1 U12373 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n15221) );
  NOR2_X1 U12374 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n15221), .ZN(n10988) );
  NOR2_X1 U12375 ( .A1(n13862), .A2(n9833), .ZN(n9825) );
  AOI211_X1 U12376 ( .C1(n14604), .C2(P1_ADDR_REG_8__SCAN_IN), .A(n10988), .B(
        n9825), .ZN(n9826) );
  OAI211_X1 U12377 ( .C1(n9836), .C2(n9828), .A(n9827), .B(n9826), .ZN(
        P1_U3251) );
  INV_X1 U12378 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n10707) );
  MUX2_X1 U12379 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n10707), .S(n10872), .Z(
        n9831) );
  OAI21_X1 U12380 ( .B1(P1_REG1_REG_8__SCAN_IN), .B2(n10685), .A(n9829), .ZN(
        n9830) );
  NAND2_X1 U12381 ( .A1(n9830), .A2(n9831), .ZN(n9968) );
  OAI21_X1 U12382 ( .B1(n9831), .B2(n9830), .A(n9968), .ZN(n9844) );
  NOR2_X1 U12383 ( .A1(n9833), .A2(n9832), .ZN(n9835) );
  INV_X1 U12384 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n10703) );
  MUX2_X1 U12385 ( .A(P1_REG2_REG_9__SCAN_IN), .B(n10703), .S(n10872), .Z(
        n9834) );
  OAI21_X1 U12386 ( .B1(n9836), .B2(n9835), .A(n9834), .ZN(n9974) );
  INV_X1 U12387 ( .A(n9974), .ZN(n9838) );
  NOR3_X1 U12388 ( .A1(n9836), .A2(n9835), .A3(n9834), .ZN(n9837) );
  NOR3_X1 U12389 ( .A1(n9838), .A2(n9837), .A3(n14619), .ZN(n9843) );
  NAND2_X1 U12390 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_U3086), .ZN(n11153) );
  INV_X1 U12391 ( .A(n11153), .ZN(n9839) );
  AOI21_X1 U12392 ( .B1(n14604), .B2(P1_ADDR_REG_9__SCAN_IN), .A(n9839), .ZN(
        n9840) );
  OAI21_X1 U12393 ( .B1(n9841), .B2(n13862), .A(n9840), .ZN(n9842) );
  AOI211_X1 U12394 ( .C1(n9844), .C2(n14614), .A(n9843), .B(n9842), .ZN(n9845)
         );
  INV_X1 U12395 ( .A(n9845), .ZN(P1_U3252) );
  INV_X1 U12396 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n15170) );
  INV_X1 U12397 ( .A(n11308), .ZN(n9849) );
  INV_X1 U12398 ( .A(n11452), .ZN(n11442) );
  OAI222_X1 U12399 ( .A1(n13594), .A2(n15170), .B1(n13596), .B2(n9849), .C1(
        P2_U3088), .C2(n11442), .ZN(P2_U3313) );
  OAI21_X1 U12400 ( .B1(n9846), .B2(n6756), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n9847) );
  XNOR2_X1 U12401 ( .A(n9847), .B(P1_IR_REG_14__SCAN_IN), .ZN(n13806) );
  INV_X1 U12402 ( .A(n13806), .ZN(n9850) );
  OAI222_X1 U12403 ( .A1(n9850), .A2(P1_U3086), .B1(n11860), .B2(n9849), .C1(
        n9848), .C2(n14247), .ZN(P1_U3341) );
  INV_X1 U12404 ( .A(n10152), .ZN(n9854) );
  NOR3_X1 U12405 ( .A1(n11965), .A2(n10150), .A3(n8709), .ZN(n9852) );
  AOI211_X1 U12406 ( .C1(n9854), .C2(n9853), .A(n9852), .B(n9851), .ZN(n9859)
         );
  OAI22_X1 U12407 ( .A1(n12544), .A2(n10149), .B1(n7418), .B2(n12484), .ZN(
        n9855) );
  NAND2_X1 U12408 ( .A1(n9857), .A2(n9856), .ZN(n9998) );
  NAND2_X1 U12409 ( .A1(n9998), .A2(P3_REG3_REG_1__SCAN_IN), .ZN(n9858) );
  OAI211_X1 U12410 ( .C1(n9859), .C2(n12507), .A(n6697), .B(n9858), .ZN(
        P3_U3162) );
  AND2_X1 U12411 ( .A1(n9860), .A2(n9934), .ZN(n9862) );
  NOR2_X1 U12412 ( .A1(n10611), .A2(n12691), .ZN(n9864) );
  NAND2_X1 U12413 ( .A1(n12114), .A2(n9864), .ZN(n10037) );
  NAND2_X1 U12414 ( .A1(n12095), .A2(n10037), .ZN(n9866) );
  AND2_X1 U12415 ( .A1(n9866), .A2(n9865), .ZN(n9941) );
  NAND2_X1 U12416 ( .A1(n13001), .A2(n9866), .ZN(n9867) );
  OAI21_X1 U12417 ( .B1(n13001), .B2(n9941), .A(n9867), .ZN(n9868) );
  INV_X1 U12418 ( .A(n9868), .ZN(n9869) );
  NAND2_X1 U12419 ( .A1(n9943), .A2(n9869), .ZN(n9872) );
  NOR2_X2 U12420 ( .A1(n11177), .A2(n15099), .ZN(n14423) );
  AOI22_X1 U12421 ( .A1(n14423), .A2(n9949), .B1(n15058), .B2(
        P3_REG3_REG_0__SCAN_IN), .ZN(n9875) );
  NAND2_X1 U12422 ( .A1(n11969), .A2(n11966), .ZN(n9948) );
  AND2_X1 U12423 ( .A1(n9928), .A2(n15099), .ZN(n9871) );
  AND2_X1 U12424 ( .A1(n10041), .A2(n15052), .ZN(n9870) );
  AOI21_X1 U12425 ( .B1(n9948), .B2(n9871), .A(n9870), .ZN(n9944) );
  MUX2_X1 U12426 ( .A(n9944), .B(n9873), .S(n15066), .Z(n9874) );
  NAND2_X1 U12427 ( .A1(n9875), .A2(n9874), .ZN(P3_U3233) );
  INV_X1 U12428 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n9877) );
  MUX2_X1 U12429 ( .A(n9877), .B(P2_REG1_REG_7__SCAN_IN), .S(n14806), .Z(
        n14802) );
  INV_X1 U12430 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n9878) );
  MUX2_X1 U12431 ( .A(n9878), .B(P2_REG1_REG_8__SCAN_IN), .S(n14819), .Z(
        n14815) );
  AOI21_X1 U12432 ( .B1(n14819), .B2(P2_REG1_REG_8__SCAN_IN), .A(n14814), .ZN(
        n9881) );
  MUX2_X1 U12433 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n9879), .S(n10168), .Z(n9880) );
  OAI21_X1 U12434 ( .B1(n9881), .B2(n9880), .A(n10164), .ZN(n9882) );
  NAND2_X1 U12435 ( .A1(n9882), .A2(n14853), .ZN(n9892) );
  AOI21_X1 U12436 ( .B1(n9884), .B2(P2_REG2_REG_6__SCAN_IN), .A(n9883), .ZN(
        n14809) );
  MUX2_X1 U12437 ( .A(n7850), .B(P2_REG2_REG_7__SCAN_IN), .S(n14806), .Z(
        n14808) );
  AOI21_X1 U12438 ( .B1(n14806), .B2(P2_REG2_REG_7__SCAN_IN), .A(n14807), .ZN(
        n14822) );
  MUX2_X1 U12439 ( .A(n10736), .B(P2_REG2_REG_8__SCAN_IN), .S(n14819), .Z(
        n14821) );
  AOI21_X1 U12440 ( .B1(n14819), .B2(P2_REG2_REG_8__SCAN_IN), .A(n14820), .ZN(
        n9887) );
  INV_X1 U12441 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n9885) );
  MUX2_X1 U12442 ( .A(P2_REG2_REG_9__SCAN_IN), .B(n9885), .S(n10168), .Z(n9886) );
  NAND2_X1 U12443 ( .A1(n9887), .A2(n9886), .ZN(n10167) );
  OAI21_X1 U12444 ( .B1(n9887), .B2(n9886), .A(n10167), .ZN(n9890) );
  INV_X1 U12445 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n15353) );
  NAND2_X1 U12446 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3088), .ZN(n10570) );
  NAND2_X1 U12447 ( .A1(n14868), .A2(n10168), .ZN(n9888) );
  OAI211_X1 U12448 ( .C1(n14874), .C2(n15353), .A(n10570), .B(n9888), .ZN(
        n9889) );
  AOI21_X1 U12449 ( .B1(n9890), .B2(n14870), .A(n9889), .ZN(n9891) );
  NAND2_X1 U12450 ( .A1(n9892), .A2(n9891), .ZN(P2_U3223) );
  OR2_X1 U12451 ( .A1(n9894), .A2(n9893), .ZN(n9895) );
  AND2_X1 U12452 ( .A1(n9896), .A2(n9895), .ZN(n10006) );
  MUX2_X1 U12453 ( .A(n10006), .B(n9897), .S(n14601), .Z(n9900) );
  AOI21_X1 U12454 ( .B1(n14601), .B2(n9603), .A(n9450), .ZN(n14600) );
  OAI21_X1 U12455 ( .B1(n14600), .B2(P1_IR_REG_0__SCAN_IN), .A(P1_U4016), .ZN(
        n9898) );
  AOI21_X1 U12456 ( .B1(n9900), .B2(n9899), .A(n9898), .ZN(n9925) );
  AOI211_X1 U12457 ( .C1(n9903), .C2(n9902), .A(n9901), .B(n14619), .ZN(n9912)
         );
  AOI211_X1 U12458 ( .C1(n9906), .C2(n9905), .A(n9904), .B(n13847), .ZN(n9911)
         );
  NAND2_X1 U12459 ( .A1(n14604), .A2(P1_ADDR_REG_2__SCAN_IN), .ZN(n9908) );
  NAND2_X1 U12460 ( .A1(P1_U3086), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n9907) );
  OAI211_X1 U12461 ( .C1(n13862), .C2(n9909), .A(n9908), .B(n9907), .ZN(n9910)
         );
  OR4_X1 U12462 ( .A1(n9925), .A2(n9912), .A3(n9911), .A4(n9910), .ZN(P1_U3245) );
  AOI211_X1 U12463 ( .C1(n9915), .C2(n9914), .A(n13847), .B(n9913), .ZN(n9924)
         );
  AND3_X1 U12464 ( .A1(n9918), .A2(n9917), .A3(n9916), .ZN(n9919) );
  NOR3_X1 U12465 ( .A1(n14619), .A2(n9920), .A3(n9919), .ZN(n9923) );
  NAND2_X1 U12466 ( .A1(n14604), .A2(P1_ADDR_REG_4__SCAN_IN), .ZN(n9921) );
  NAND2_X1 U12467 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n10630) );
  OAI211_X1 U12468 ( .C1(n13862), .C2(n10306), .A(n9921), .B(n10630), .ZN(
        n9922) );
  OR4_X1 U12469 ( .A1(n9925), .A2(n9924), .A3(n9923), .A4(n9922), .ZN(P1_U3247) );
  INV_X1 U12470 ( .A(n12680), .ZN(n12672) );
  INV_X1 U12471 ( .A(n9926), .ZN(n9927) );
  OAI222_X1 U12472 ( .A1(P3_U3151), .A2(n12672), .B1(n14368), .B2(n15158), 
        .C1(n14370), .C2(n9927), .ZN(P3_U3278) );
  AND2_X1 U12473 ( .A1(n9929), .A2(n9928), .ZN(n9932) );
  INV_X1 U12474 ( .A(n10040), .ZN(n9931) );
  OAI22_X1 U12475 ( .A1(n9933), .A2(n9932), .B1(n9931), .B2(n9930), .ZN(n9935)
         );
  INV_X1 U12476 ( .A(n12988), .ZN(n12980) );
  MUX2_X1 U12477 ( .A(n8688), .B(n9944), .S(n15110), .Z(n9936) );
  OAI21_X1 U12478 ( .B1(n12980), .B2(n9947), .A(n9936), .ZN(P3_U3390) );
  OAI22_X1 U12479 ( .A1(n15099), .A2(n9937), .B1(n12691), .B2(n11288), .ZN(
        n9938) );
  AOI21_X1 U12480 ( .B1(n9938), .B2(n12103), .A(n6529), .ZN(n9940) );
  MUX2_X1 U12481 ( .A(n9941), .B(n9940), .S(n9939), .Z(n9942) );
  INV_X1 U12482 ( .A(n12913), .ZN(n12907) );
  MUX2_X1 U12483 ( .A(n9945), .B(n9944), .S(n15131), .Z(n9946) );
  OAI21_X1 U12484 ( .B1(n12907), .B2(n9947), .A(n9946), .ZN(P3_U3459) );
  INV_X1 U12485 ( .A(n9948), .ZN(n11923) );
  NAND2_X1 U12486 ( .A1(n9998), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n9951) );
  AOI22_X1 U12487 ( .A1(n12535), .A2(n10041), .B1(n12524), .B2(n9949), .ZN(
        n9950) );
  OAI211_X1 U12488 ( .C1(n11923), .C2(n12507), .A(n9951), .B(n9950), .ZN(
        P3_U3172) );
  INV_X1 U12489 ( .A(n11494), .ZN(n9985) );
  OAI21_X1 U12490 ( .B1(n9954), .B2(n9953), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n9955) );
  MUX2_X1 U12491 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9955), .S(
        P1_IR_REG_15__SCAN_IN), .Z(n9956) );
  AND2_X1 U12492 ( .A1(n9952), .A2(n9956), .ZN(n14615) );
  AOI22_X1 U12493 ( .A1(n14615), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n14244), .ZN(n9957) );
  OAI21_X1 U12494 ( .B1(n9985), .B2(n11860), .A(n9957), .ZN(P1_U3340) );
  NOR2_X1 U12495 ( .A1(n9958), .A2(P2_U3088), .ZN(n10426) );
  OAI21_X1 U12496 ( .B1(n13269), .B2(n14474), .A(n14458), .ZN(n9959) );
  INV_X1 U12497 ( .A(n14469), .ZN(n13117) );
  AOI22_X1 U12498 ( .A1(n9960), .A2(n9959), .B1(n13117), .B2(n7753), .ZN(n9967) );
  NAND4_X1 U12499 ( .A1(n9963), .A2(n9962), .A3(n10357), .A4(n9961), .ZN(n9964) );
  OAI21_X1 U12500 ( .B1(n14474), .B2(n10210), .A(n9964), .ZN(n9965) );
  INV_X1 U12501 ( .A(n9965), .ZN(n9966) );
  OAI211_X1 U12502 ( .C1(n10426), .C2(n7761), .A(n9967), .B(n9966), .ZN(
        P2_U3204) );
  INV_X1 U12503 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n10880) );
  MUX2_X1 U12504 ( .A(n10880), .B(P1_REG1_REG_10__SCAN_IN), .S(n10999), .Z(
        n9970) );
  OAI21_X1 U12505 ( .B1(n10872), .B2(P1_REG1_REG_9__SCAN_IN), .A(n9968), .ZN(
        n9969) );
  NOR2_X1 U12506 ( .A1(n9969), .A2(n9970), .ZN(n10021) );
  AOI211_X1 U12507 ( .C1(n9970), .C2(n9969), .A(n13847), .B(n10021), .ZN(n9980) );
  NAND2_X1 U12508 ( .A1(n10872), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n9973) );
  INV_X1 U12509 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n9971) );
  MUX2_X1 U12510 ( .A(n9971), .B(P1_REG2_REG_10__SCAN_IN), .S(n10999), .Z(
        n9972) );
  AOI21_X1 U12511 ( .B1(n9974), .B2(n9973), .A(n9972), .ZN(n10027) );
  INV_X1 U12512 ( .A(n10027), .ZN(n9976) );
  NAND3_X1 U12513 ( .A1(n9974), .A2(n9973), .A3(n9972), .ZN(n9975) );
  NAND3_X1 U12514 ( .A1(n9976), .A2(n13866), .A3(n9975), .ZN(n9978) );
  NOR2_X1 U12515 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n15304), .ZN(n11266) );
  AOI21_X1 U12516 ( .B1(n14604), .B2(P1_ADDR_REG_10__SCAN_IN), .A(n11266), 
        .ZN(n9977) );
  OAI211_X1 U12517 ( .C1(n13862), .C2(n10024), .A(n9978), .B(n9977), .ZN(n9979) );
  OR2_X1 U12518 ( .A1(n9980), .A2(n9979), .ZN(P1_U3253) );
  INV_X1 U12519 ( .A(n9981), .ZN(n9982) );
  OAI222_X1 U12520 ( .A1(P3_U3151), .A2(n12693), .B1(n14368), .B2(n9983), .C1(
        n14370), .C2(n9982), .ZN(P3_U3277) );
  INV_X1 U12521 ( .A(n14867), .ZN(n11453) );
  OAI222_X1 U12522 ( .A1(P2_U3088), .A2(n11453), .B1(n13596), .B2(n9985), .C1(
        n9984), .C2(n13588), .ZN(P2_U3312) );
  OAI21_X1 U12523 ( .B1(n9988), .B2(n9987), .A(n9986), .ZN(n9989) );
  NAND2_X1 U12524 ( .A1(n9989), .A2(n14535), .ZN(n9993) );
  NAND2_X1 U12525 ( .A1(n13601), .A2(n9990), .ZN(n10018) );
  AOI22_X1 U12526 ( .A1(n13897), .A2(n6770), .B1(n13776), .B2(n13732), .ZN(
        n10664) );
  INV_X1 U12527 ( .A(n10664), .ZN(n9991) );
  AOI22_X1 U12528 ( .A1(n10018), .A2(P1_REG3_REG_2__SCAN_IN), .B1(n14537), 
        .B2(n9991), .ZN(n9992) );
  OAI211_X1 U12529 ( .C1(n10298), .C2(n13753), .A(n9993), .B(n9992), .ZN(
        P1_U3237) );
  XOR2_X1 U12530 ( .A(n9995), .B(n9994), .Z(n10000) );
  AOI22_X1 U12531 ( .A1(n12535), .A2(n15054), .B1(n12524), .B2(n10096), .ZN(
        n9996) );
  OAI21_X1 U12532 ( .B1(n7482), .B2(n12537), .A(n9996), .ZN(n9997) );
  AOI21_X1 U12533 ( .B1(P3_REG3_REG_2__SCAN_IN), .B2(n9998), .A(n9997), .ZN(
        n9999) );
  OAI21_X1 U12534 ( .B1(n10000), .B2(n12507), .A(n9999), .ZN(P3_U3177) );
  OAI222_X1 U12535 ( .A1(n14370), .A2(n10002), .B1(n14368), .B2(n10001), .C1(
        P3_U3151), .C2(n12700), .ZN(P3_U3276) );
  INV_X1 U12536 ( .A(n11499), .ZN(n10010) );
  NAND2_X1 U12537 ( .A1(n9952), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10003) );
  MUX2_X1 U12538 ( .A(P1_IR_REG_31__SCAN_IN), .B(n10003), .S(
        P1_IR_REG_16__SCAN_IN), .Z(n10004) );
  AND2_X1 U12539 ( .A1(n10004), .A2(n9172), .ZN(n13820) );
  AOI22_X1 U12540 ( .A1(n13820), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n14244), .ZN(n10005) );
  OAI21_X1 U12541 ( .B1(n10010), .B2(n11860), .A(n10005), .ZN(P1_U3339) );
  NAND2_X1 U12542 ( .A1(n14537), .A2(n13732), .ZN(n11269) );
  OAI22_X1 U12543 ( .A1(n11269), .A2(n6719), .B1(n13727), .B2(n10006), .ZN(
        n10007) );
  AOI21_X1 U12544 ( .B1(P1_REG3_REG_0__SCAN_IN), .B2(n10018), .A(n10007), .ZN(
        n10008) );
  OAI21_X1 U12545 ( .B1(n14677), .B2(n13753), .A(n10008), .ZN(P1_U3232) );
  INV_X1 U12546 ( .A(n11455), .ZN(n13190) );
  OAI222_X1 U12547 ( .A1(P2_U3088), .A2(n13190), .B1(n13596), .B2(n10010), 
        .C1(n10009), .C2(n13588), .ZN(P2_U3311) );
  INV_X1 U12548 ( .A(n10011), .ZN(n10012) );
  AOI21_X1 U12549 ( .B1(n10014), .B2(n10013), .A(n10012), .ZN(n10020) );
  NOR2_X1 U12550 ( .A1(n13753), .A2(n14698), .ZN(n10017) );
  INV_X1 U12551 ( .A(n13897), .ZN(n13674) );
  NOR2_X1 U12552 ( .A1(n13715), .A2(n13674), .ZN(n11267) );
  INV_X1 U12553 ( .A(n11267), .ZN(n10015) );
  INV_X1 U12554 ( .A(n13780), .ZN(n10539) );
  INV_X1 U12555 ( .A(n13778), .ZN(n10538) );
  OAI22_X1 U12556 ( .A1(n10015), .A2(n10539), .B1(n10538), .B2(n11269), .ZN(
        n10016) );
  AOI211_X1 U12557 ( .C1(P1_REG3_REG_1__SCAN_IN), .C2(n10018), .A(n10017), .B(
        n10016), .ZN(n10019) );
  OAI21_X1 U12558 ( .B1(n10020), .B2(n13727), .A(n10019), .ZN(P1_U3222) );
  INV_X1 U12559 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n11007) );
  MUX2_X1 U12560 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n11007), .S(n11049), .Z(
        n10022) );
  NAND2_X1 U12561 ( .A1(n10023), .A2(n10022), .ZN(n10318) );
  OAI21_X1 U12562 ( .B1(n10023), .B2(n10022), .A(n10318), .ZN(n10033) );
  NOR2_X1 U12563 ( .A1(n10024), .A2(n9971), .ZN(n10026) );
  INV_X1 U12564 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n11063) );
  MUX2_X1 U12565 ( .A(P1_REG2_REG_11__SCAN_IN), .B(n11063), .S(n11049), .Z(
        n10025) );
  OAI21_X1 U12566 ( .B1(n10027), .B2(n10026), .A(n10025), .ZN(n10321) );
  OR3_X1 U12567 ( .A1(n10027), .A2(n10026), .A3(n10025), .ZN(n10028) );
  NAND3_X1 U12568 ( .A1(n10321), .A2(n13866), .A3(n10028), .ZN(n10031) );
  NAND2_X1 U12569 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n11382)
         );
  INV_X1 U12570 ( .A(n11382), .ZN(n10029) );
  AOI21_X1 U12571 ( .B1(n14604), .B2(P1_ADDR_REG_11__SCAN_IN), .A(n10029), 
        .ZN(n10030) );
  OAI211_X1 U12572 ( .C1(n13862), .C2(n10322), .A(n10031), .B(n10030), .ZN(
        n10032) );
  AOI21_X1 U12573 ( .B1(n10033), .B2(n14614), .A(n10032), .ZN(n10034) );
  INV_X1 U12574 ( .A(n10034), .ZN(P1_U3254) );
  INV_X1 U12575 ( .A(n11975), .ZN(n10044) );
  XNOR2_X1 U12576 ( .A(n10094), .B(n10044), .ZN(n15070) );
  OR2_X1 U12577 ( .A1(n6523), .A2(n12104), .ZN(n15031) );
  OR2_X1 U12578 ( .A1(n15066), .A2(n15031), .ZN(n10821) );
  NAND2_X1 U12579 ( .A1(n10096), .A2(n14441), .ZN(n15071) );
  NOR2_X1 U12580 ( .A1(n15071), .A2(n11287), .ZN(n10049) );
  AND2_X1 U12581 ( .A1(n15099), .A2(n10036), .ZN(n10039) );
  INV_X1 U12582 ( .A(n10037), .ZN(n10038) );
  NAND2_X1 U12583 ( .A1(n10153), .A2(n10152), .ZN(n10151) );
  OR2_X1 U12584 ( .A1(n10041), .A2(n7481), .ZN(n10042) );
  NAND2_X1 U12585 ( .A1(n10151), .A2(n10042), .ZN(n10043) );
  NAND2_X1 U12586 ( .A1(n10043), .A2(n10044), .ZN(n10100) );
  OAI21_X1 U12587 ( .B1(n10044), .B2(n10043), .A(n10100), .ZN(n10047) );
  NAND2_X2 U12588 ( .A1(n10045), .A2(n6876), .ZN(n15056) );
  INV_X1 U12589 ( .A(n15038), .ZN(n12864) );
  INV_X1 U12590 ( .A(n15054), .ZN(n10112) );
  INV_X1 U12591 ( .A(n15052), .ZN(n12866) );
  OAI22_X1 U12592 ( .A1(n7482), .A2(n12864), .B1(n10112), .B2(n12866), .ZN(
        n10046) );
  AOI21_X1 U12593 ( .B1(n10047), .B2(n15056), .A(n10046), .ZN(n10048) );
  OAI21_X1 U12594 ( .B1(n15039), .B2(n15070), .A(n10048), .ZN(n15072) );
  AOI211_X1 U12595 ( .C1(n15058), .C2(P3_REG3_REG_2__SCAN_IN), .A(n10049), .B(
        n15072), .ZN(n10050) );
  INV_X2 U12596 ( .A(n15066), .ZN(n15049) );
  MUX2_X1 U12597 ( .A(n10051), .B(n10050), .S(n15049), .Z(n10052) );
  OAI21_X1 U12598 ( .B1(n15070), .B2(n10821), .A(n10052), .ZN(P3_U3231) );
  NAND2_X1 U12599 ( .A1(n10054), .A2(n10053), .ZN(n10059) );
  INV_X1 U12600 ( .A(n10055), .ZN(n10057) );
  NAND2_X1 U12601 ( .A1(n10057), .A2(n10056), .ZN(n10058) );
  NAND2_X1 U12602 ( .A1(n10059), .A2(n10058), .ZN(n14964) );
  MUX2_X1 U12603 ( .A(P3_REG2_REG_5__SCAN_IN), .B(P3_REG1_REG_5__SCAN_IN), .S(
        n12670), .Z(n10060) );
  XNOR2_X1 U12604 ( .A(n10060), .B(n14966), .ZN(n14963) );
  NAND2_X1 U12605 ( .A1(n14964), .A2(n14963), .ZN(n10063) );
  INV_X1 U12606 ( .A(n10060), .ZN(n10061) );
  NAND2_X1 U12607 ( .A1(n10061), .A2(n14966), .ZN(n10062) );
  NAND2_X1 U12608 ( .A1(n10063), .A2(n10062), .ZN(n14984) );
  MUX2_X1 U12609 ( .A(P3_REG2_REG_6__SCAN_IN), .B(P3_REG1_REG_6__SCAN_IN), .S(
        n12670), .Z(n10064) );
  XNOR2_X1 U12610 ( .A(n10064), .B(n14986), .ZN(n14983) );
  INV_X1 U12611 ( .A(n10064), .ZN(n10065) );
  MUX2_X1 U12612 ( .A(P3_REG2_REG_7__SCAN_IN), .B(P3_REG1_REG_7__SCAN_IN), .S(
        n12670), .Z(n10066) );
  XOR2_X1 U12613 ( .A(n15004), .B(n10066), .Z(n15002) );
  OAI22_X1 U12614 ( .A1(n15003), .A2(n15002), .B1(n10066), .B2(n10081), .ZN(
        n10647) );
  MUX2_X1 U12615 ( .A(P3_REG2_REG_8__SCAN_IN), .B(P3_REG1_REG_8__SCAN_IN), .S(
        n12670), .Z(n10644) );
  XNOR2_X1 U12616 ( .A(n10644), .B(n10651), .ZN(n10646) );
  XNOR2_X1 U12617 ( .A(n10647), .B(n10646), .ZN(n10092) );
  NOR2_X1 U12618 ( .A1(n14966), .A2(n10068), .ZN(n10069) );
  INV_X1 U12619 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n15156) );
  INV_X1 U12620 ( .A(P3_REG2_REG_6__SCAN_IN), .ZN(n15325) );
  AOI22_X1 U12621 ( .A1(n14986), .A2(P3_REG2_REG_6__SCAN_IN), .B1(n15325), 
        .B2(n14354), .ZN(n14976) );
  NOR2_X1 U12622 ( .A1(n14986), .A2(n15325), .ZN(n10070) );
  INV_X1 U12623 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n15316) );
  INV_X1 U12624 ( .A(P3_REG2_REG_8__SCAN_IN), .ZN(n10073) );
  AOI22_X1 U12625 ( .A1(n10651), .A2(P3_REG2_REG_8__SCAN_IN), .B1(n10073), 
        .B2(n14367), .ZN(n10074) );
  NOR2_X1 U12626 ( .A1(n10075), .A2(n10074), .ZN(n10640) );
  AOI21_X1 U12627 ( .B1(n10075), .B2(n10074), .A(n10640), .ZN(n10076) );
  NOR2_X1 U12628 ( .A1(n10076), .A2(n15023), .ZN(n10091) );
  NOR2_X1 U12629 ( .A1(n14966), .A2(n10078), .ZN(n10079) );
  INV_X1 U12630 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n15119) );
  INV_X1 U12631 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n15121) );
  AOI22_X1 U12632 ( .A1(n14986), .A2(P3_REG1_REG_6__SCAN_IN), .B1(n15121), 
        .B2(n14354), .ZN(n14980) );
  INV_X1 U12633 ( .A(n10080), .ZN(n10083) );
  INV_X1 U12634 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n15123) );
  OAI21_X1 U12635 ( .B1(n10082), .B2(n10081), .A(n10080), .ZN(n14996) );
  INV_X1 U12636 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n15125) );
  AOI22_X1 U12637 ( .A1(n10651), .A2(P3_REG1_REG_8__SCAN_IN), .B1(n15125), 
        .B2(n14367), .ZN(n10084) );
  AOI21_X1 U12638 ( .B1(n10085), .B2(n10084), .A(n10652), .ZN(n10089) );
  NOR2_X1 U12639 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10086), .ZN(n10760) );
  AOI21_X1 U12640 ( .B1(n15001), .B2(P3_ADDR_REG_8__SCAN_IN), .A(n10760), .ZN(
        n10088) );
  NAND2_X1 U12641 ( .A1(n15013), .A2(n10651), .ZN(n10087) );
  OAI211_X1 U12642 ( .C1(n10089), .C2(n15018), .A(n10088), .B(n10087), .ZN(
        n10090) );
  AOI211_X1 U12643 ( .C1(n15015), .C2(n10092), .A(n10091), .B(n10090), .ZN(
        n10093) );
  INV_X1 U12644 ( .A(n10093), .ZN(P3_U3190) );
  NAND2_X1 U12645 ( .A1(n15054), .A2(n15075), .ZN(n11985) );
  AND2_X2 U12646 ( .A1(n11987), .A2(n11985), .ZN(n11925) );
  NAND2_X1 U12647 ( .A1(n10094), .A2(n11975), .ZN(n10095) );
  INV_X1 U12648 ( .A(n10096), .ZN(n11982) );
  OR2_X1 U12649 ( .A1(n12557), .A2(n11982), .ZN(n11977) );
  XOR2_X1 U12650 ( .A(n11925), .B(n10361), .Z(n15076) );
  AOI22_X1 U12651 ( .A1(n15038), .A2(n12557), .B1(n15037), .B2(n15052), .ZN(
        n10103) );
  INV_X1 U12652 ( .A(n10100), .ZN(n10097) );
  NOR2_X1 U12653 ( .A1(n12557), .A2(n10096), .ZN(n10098) );
  OAI21_X1 U12654 ( .B1(n10097), .B2(n10098), .A(n11925), .ZN(n10101) );
  NOR2_X1 U12655 ( .A1(n11925), .A2(n10098), .ZN(n10099) );
  NAND2_X1 U12656 ( .A1(n10100), .A2(n10099), .ZN(n10368) );
  NAND3_X1 U12657 ( .A1(n10101), .A2(n15056), .A3(n10368), .ZN(n10102) );
  OAI211_X1 U12658 ( .C1(n15076), .C2(n15039), .A(n10103), .B(n10102), .ZN(
        n15078) );
  NAND2_X1 U12659 ( .A1(n15078), .A2(n15049), .ZN(n10106) );
  OAI22_X1 U12660 ( .A1(n15049), .A2(n14943), .B1(n12868), .B2(
        P3_REG3_REG_3__SCAN_IN), .ZN(n10104) );
  AOI21_X1 U12661 ( .B1(n12433), .B2(n14423), .A(n10104), .ZN(n10105) );
  OAI211_X1 U12662 ( .C1(n15076), .C2(n10821), .A(n10106), .B(n10105), .ZN(
        P3_U3230) );
  INV_X1 U12663 ( .A(n15057), .ZN(n10117) );
  INV_X1 U12664 ( .A(n12540), .ZN(n12486) );
  OAI21_X1 U12665 ( .B1(n10109), .B2(n10108), .A(n10107), .ZN(n10110) );
  NAND2_X1 U12666 ( .A1(n10110), .A2(n12533), .ZN(n10116) );
  INV_X1 U12667 ( .A(n15061), .ZN(n10369) );
  OAI22_X1 U12668 ( .A1(n12537), .A2(n10112), .B1(n10111), .B2(n12484), .ZN(
        n10113) );
  AOI211_X1 U12669 ( .C1(n10369), .C2(n12524), .A(n10114), .B(n10113), .ZN(
        n10115) );
  OAI211_X1 U12670 ( .C1(n10117), .C2(n12486), .A(n10116), .B(n10115), .ZN(
        P3_U3170) );
  INV_X1 U12671 ( .A(n10118), .ZN(n10119) );
  AOI21_X1 U12672 ( .B1(n10266), .B2(n10119), .A(n14474), .ZN(n10123) );
  NOR3_X1 U12673 ( .A1(n13124), .A2(n10121), .A3(n10120), .ZN(n10122) );
  OAI21_X1 U12674 ( .B1(n10123), .B2(n10122), .A(n10281), .ZN(n10129) );
  NAND2_X1 U12675 ( .A1(n13154), .A2(n13402), .ZN(n10125) );
  NAND2_X1 U12676 ( .A1(n13156), .A2(n13401), .ZN(n10124) );
  AND2_X1 U12677 ( .A1(n10125), .A2(n10124), .ZN(n10203) );
  INV_X1 U12678 ( .A(n10203), .ZN(n10127) );
  NOR2_X1 U12679 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7851), .ZN(n14805) );
  NOR2_X1 U12680 ( .A1(n14467), .A2(n10493), .ZN(n10126) );
  AOI211_X1 U12681 ( .C1(n13131), .C2(n10127), .A(n14805), .B(n10126), .ZN(
        n10128) );
  OAI211_X1 U12682 ( .C1(n10492), .C2(n14458), .A(n10129), .B(n10128), .ZN(
        P2_U3185) );
  NAND2_X1 U12683 ( .A1(n11783), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n10140) );
  INV_X1 U12684 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n15240) );
  OR2_X1 U12685 ( .A1(n11784), .A2(n15240), .ZN(n10139) );
  INV_X1 U12686 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n15369) );
  NAND2_X1 U12687 ( .A1(P1_REG3_REG_18__SCAN_IN), .A2(P1_REG3_REG_17__SCAN_IN), 
        .ZN(n10130) );
  NAND2_X1 U12688 ( .A1(n11540), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n11552) );
  INV_X1 U12689 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n15196) );
  INV_X1 U12690 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n13637) );
  NAND2_X1 U12691 ( .A1(n11561), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n11562) );
  NAND2_X1 U12692 ( .A1(n11578), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n11577) );
  NAND2_X1 U12693 ( .A1(n11477), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n11476) );
  NAND2_X1 U12694 ( .A1(P1_REG3_REG_25__SCAN_IN), .A2(n11468), .ZN(n11588) );
  INV_X1 U12695 ( .A(n11588), .ZN(n10131) );
  NAND2_X1 U12696 ( .A1(n10131), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n11599) );
  INV_X1 U12697 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n13607) );
  INV_X1 U12698 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n10132) );
  OAI21_X1 U12699 ( .B1(n11599), .B2(n13607), .A(n10132), .ZN(n10135) );
  INV_X1 U12700 ( .A(n11599), .ZN(n10134) );
  AND2_X1 U12701 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(P1_REG3_REG_28__SCAN_IN), 
        .ZN(n10133) );
  NAND2_X1 U12702 ( .A1(n10134), .A2(n10133), .ZN(n13900) );
  NAND2_X1 U12703 ( .A1(n10135), .A2(n13900), .ZN(n13923) );
  OR2_X1 U12704 ( .A1(n11600), .A2(n13923), .ZN(n10138) );
  INV_X1 U12705 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n10136) );
  OR2_X1 U12706 ( .A1(n6526), .A2(n10136), .ZN(n10137) );
  NAND4_X1 U12707 ( .A1(n10140), .A2(n10139), .A3(n10138), .A4(n10137), .ZN(
        n13913) );
  NAND2_X1 U12708 ( .A1(n13913), .A2(P1_U4016), .ZN(n10141) );
  OAI21_X1 U12709 ( .B1(n13777), .B2(n13587), .A(n10141), .ZN(P1_U3588) );
  NAND2_X1 U12710 ( .A1(n10142), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n10143) );
  NAND2_X1 U12711 ( .A1(n12712), .A2(n10143), .ZN(n12726) );
  INV_X1 U12712 ( .A(P3_REG1_REG_28__SCAN_IN), .ZN(n15404) );
  NAND2_X1 U12713 ( .A1(n11899), .A2(P3_REG2_REG_28__SCAN_IN), .ZN(n10146) );
  NAND2_X1 U12714 ( .A1(n10144), .A2(P3_REG0_REG_28__SCAN_IN), .ZN(n10145) );
  OAI211_X1 U12715 ( .C1(n15404), .C2(n8978), .A(n10146), .B(n10145), .ZN(
        n10147) );
  NAND2_X1 U12716 ( .A1(n12548), .A2(P3_DATAO_REG_28__SCAN_IN), .ZN(n10148) );
  OAI21_X1 U12717 ( .B1(n12736), .B2(n12548), .A(n10148), .ZN(P3_U3519) );
  NOR2_X1 U12718 ( .A1(n10149), .A2(n15099), .ZN(n15068) );
  XNOR2_X1 U12719 ( .A(n10150), .B(n11965), .ZN(n15069) );
  INV_X1 U12720 ( .A(n15069), .ZN(n10157) );
  OAI21_X1 U12721 ( .B1(n10153), .B2(n10152), .A(n10151), .ZN(n10154) );
  NAND2_X1 U12722 ( .A1(n10154), .A2(n15056), .ZN(n10156) );
  OAI211_X1 U12723 ( .C1(n10157), .C2(n15039), .A(n10156), .B(n10155), .ZN(
        n15067) );
  AOI21_X1 U12724 ( .B1(n15068), .B2(n12104), .A(n15067), .ZN(n10162) );
  INV_X1 U12725 ( .A(n10821), .ZN(n12744) );
  OAI22_X1 U12726 ( .A1(n15049), .A2(n10159), .B1(n10158), .B2(n12868), .ZN(
        n10160) );
  AOI21_X1 U12727 ( .B1(n12744), .B2(n15069), .A(n10160), .ZN(n10161) );
  OAI21_X1 U12728 ( .B1(n15066), .B2(n10162), .A(n10161), .ZN(P3_U3232) );
  INV_X1 U12729 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n10163) );
  MUX2_X1 U12730 ( .A(n10163), .B(P2_REG1_REG_10__SCAN_IN), .S(n11026), .Z(
        n10166) );
  OAI21_X1 U12731 ( .B1(n10168), .B2(P2_REG1_REG_9__SCAN_IN), .A(n10164), .ZN(
        n10165) );
  NOR2_X1 U12732 ( .A1(n10165), .A2(n10166), .ZN(n11021) );
  AOI211_X1 U12733 ( .C1(n10166), .C2(n10165), .A(n14863), .B(n11021), .ZN(
        n10176) );
  OAI21_X1 U12734 ( .B1(n10168), .B2(P2_REG2_REG_9__SCAN_IN), .A(n10167), .ZN(
        n10170) );
  MUX2_X1 U12735 ( .A(n10775), .B(P2_REG2_REG_10__SCAN_IN), .S(n11026), .Z(
        n10169) );
  AOI211_X1 U12736 ( .C1(n10170), .C2(n10169), .A(n14836), .B(n11025), .ZN(
        n10175) );
  INV_X1 U12737 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n10173) );
  NOR2_X1 U12738 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n15210), .ZN(n10171) );
  AOI21_X1 U12739 ( .B1(n14868), .B2(n11026), .A(n10171), .ZN(n10172) );
  OAI21_X1 U12740 ( .B1(n14874), .B2(n10173), .A(n10172), .ZN(n10174) );
  OR3_X1 U12741 ( .A1(n10176), .A2(n10175), .A3(n10174), .ZN(P2_U3224) );
  NAND2_X1 U12742 ( .A1(n9172), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10177) );
  XNOR2_X1 U12743 ( .A(n10177), .B(P1_IR_REG_17__SCAN_IN), .ZN(n13844) );
  INV_X1 U12744 ( .A(n13844), .ZN(n13838) );
  INV_X1 U12745 ( .A(n11511), .ZN(n10180) );
  OAI222_X1 U12746 ( .A1(P1_U3086), .A2(n13838), .B1(n11860), .B2(n10180), 
        .C1(n10178), .C2(n14247), .ZN(P1_U3338) );
  OAI222_X1 U12747 ( .A1(P2_U3088), .A2(n13211), .B1(n13596), .B2(n10180), 
        .C1(n10179), .C2(n13588), .ZN(P2_U3310) );
  INV_X1 U12748 ( .A(n14923), .ZN(n14901) );
  OAI21_X1 U12749 ( .B1(n10182), .B2(n10185), .A(n10181), .ZN(n10514) );
  NAND2_X1 U12750 ( .A1(n10223), .A2(n10487), .ZN(n10183) );
  NAND2_X1 U12751 ( .A1(n10183), .A2(n13316), .ZN(n10184) );
  NOR2_X1 U12752 ( .A1(n10200), .A2(n10184), .ZN(n10521) );
  XNOR2_X1 U12753 ( .A(n10186), .B(n10185), .ZN(n10189) );
  NAND2_X1 U12754 ( .A1(n13155), .A2(n13402), .ZN(n10188) );
  NAND2_X1 U12755 ( .A1(n13157), .A2(n13401), .ZN(n10187) );
  AND2_X1 U12756 ( .A1(n10188), .A2(n10187), .ZN(n10262) );
  OAI21_X1 U12757 ( .B1(n10189), .B2(n13534), .A(n10262), .ZN(n10515) );
  AOI211_X1 U12758 ( .C1(n14515), .C2(n10514), .A(n10521), .B(n10515), .ZN(
        n10489) );
  AND2_X1 U12759 ( .A1(n10190), .A2(n14891), .ZN(n14892) );
  NAND3_X1 U12760 ( .A1(n14892), .A2(n10192), .A3(n10191), .ZN(n10193) );
  OR2_X1 U12761 ( .A1(n10194), .A2(n10193), .ZN(n10354) );
  INV_X1 U12762 ( .A(n10487), .ZN(n10519) );
  OAI22_X1 U12763 ( .A1(n13573), .A2(n10519), .B1(n14925), .B2(n7839), .ZN(
        n10196) );
  INV_X1 U12764 ( .A(n10196), .ZN(n10197) );
  OAI21_X1 U12765 ( .B1(n10489), .B2(n14924), .A(n10197), .ZN(P2_U3448) );
  OAI21_X1 U12766 ( .B1(n10199), .B2(n10201), .A(n10198), .ZN(n10490) );
  AOI211_X1 U12767 ( .C1(n10484), .C2(n6903), .A(n13269), .B(n10738), .ZN(
        n10496) );
  XNOR2_X1 U12768 ( .A(n10202), .B(n10201), .ZN(n10204) );
  OAI21_X1 U12769 ( .B1(n10204), .B2(n13534), .A(n10203), .ZN(n10491) );
  AOI211_X1 U12770 ( .C1(n14515), .C2(n10490), .A(n10496), .B(n10491), .ZN(
        n10486) );
  OAI22_X1 U12771 ( .A1(n13573), .A2(n10492), .B1(n14925), .B2(n7854), .ZN(
        n10205) );
  INV_X1 U12772 ( .A(n10205), .ZN(n10206) );
  OAI21_X1 U12773 ( .B1(n10486), .B2(n14924), .A(n10206), .ZN(P2_U3451) );
  OAI21_X1 U12774 ( .B1(n10209), .B2(n10208), .A(n10207), .ZN(n10828) );
  INV_X1 U12775 ( .A(n13269), .ZN(n13316) );
  OAI211_X1 U12776 ( .C1(n10218), .C2(n10358), .A(n10236), .B(n13316), .ZN(
        n10826) );
  INV_X1 U12777 ( .A(n10826), .ZN(n10216) );
  XNOR2_X1 U12778 ( .A(n10210), .B(n10209), .ZN(n10214) );
  NAND2_X1 U12779 ( .A1(n8301), .A2(n13402), .ZN(n10212) );
  NAND2_X1 U12780 ( .A1(n8305), .A2(n13401), .ZN(n10211) );
  AND2_X1 U12781 ( .A1(n10212), .A2(n10211), .ZN(n10334) );
  INV_X1 U12782 ( .A(n10334), .ZN(n10213) );
  AOI21_X1 U12783 ( .B1(n10214), .B2(n13407), .A(n10213), .ZN(n10830) );
  INV_X1 U12784 ( .A(n10830), .ZN(n10215) );
  AOI211_X1 U12785 ( .C1(n14515), .C2(n10828), .A(n10216), .B(n10215), .ZN(
        n10483) );
  INV_X1 U12786 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n10217) );
  OAI22_X1 U12787 ( .A1(n13573), .A2(n10218), .B1(n14925), .B2(n10217), .ZN(
        n10219) );
  INV_X1 U12788 ( .A(n10219), .ZN(n10220) );
  OAI21_X1 U12789 ( .B1(n10483), .B2(n14924), .A(n10220), .ZN(P2_U3433) );
  OAI21_X1 U12790 ( .B1(n10222), .B2(n10225), .A(n10221), .ZN(n10505) );
  INV_X1 U12791 ( .A(n10223), .ZN(n10224) );
  AOI211_X1 U12792 ( .C1(n10479), .C2(n10560), .A(n13269), .B(n10224), .ZN(
        n10509) );
  XNOR2_X1 U12793 ( .A(n10226), .B(n10225), .ZN(n10229) );
  NAND2_X1 U12794 ( .A1(n13156), .A2(n13402), .ZN(n10228) );
  NAND2_X1 U12795 ( .A1(n13158), .A2(n13401), .ZN(n10227) );
  AND2_X1 U12796 ( .A1(n10228), .A2(n10227), .ZN(n10346) );
  OAI21_X1 U12797 ( .B1(n10229), .B2(n13534), .A(n10346), .ZN(n10510) );
  AOI211_X1 U12798 ( .C1(n14515), .C2(n10505), .A(n10509), .B(n10510), .ZN(
        n10481) );
  OAI22_X1 U12799 ( .A1(n13573), .A2(n6904), .B1(n14925), .B2(n7826), .ZN(
        n10230) );
  INV_X1 U12800 ( .A(n10230), .ZN(n10231) );
  OAI21_X1 U12801 ( .B1(n10481), .B2(n14924), .A(n10231), .ZN(P2_U3445) );
  OR2_X1 U12802 ( .A1(n10233), .A2(n10232), .ZN(n10234) );
  NAND2_X1 U12803 ( .A1(n10235), .A2(n10234), .ZN(n10843) );
  NAND2_X1 U12804 ( .A1(n10236), .A2(n10474), .ZN(n10237) );
  NAND2_X1 U12805 ( .A1(n10237), .A2(n13316), .ZN(n10238) );
  NOR2_X1 U12806 ( .A1(n10252), .A2(n10238), .ZN(n10842) );
  XNOR2_X1 U12807 ( .A(n10240), .B(n10239), .ZN(n10244) );
  NAND2_X1 U12808 ( .A1(n13159), .A2(n13402), .ZN(n10242) );
  NAND2_X1 U12809 ( .A1(n7753), .A2(n13401), .ZN(n10241) );
  AND2_X1 U12810 ( .A1(n10242), .A2(n10241), .ZN(n10427) );
  INV_X1 U12811 ( .A(n10427), .ZN(n10243) );
  AOI21_X1 U12812 ( .B1(n10244), .B2(n13407), .A(n10243), .ZN(n10846) );
  INV_X1 U12813 ( .A(n10846), .ZN(n10245) );
  AOI211_X1 U12814 ( .C1(n14515), .C2(n10843), .A(n10842), .B(n10245), .ZN(
        n10476) );
  INV_X1 U12815 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n10246) );
  OAI22_X1 U12816 ( .A1(n13573), .A2(n10839), .B1(n14925), .B2(n10246), .ZN(
        n10247) );
  INV_X1 U12817 ( .A(n10247), .ZN(n10248) );
  OAI21_X1 U12818 ( .B1(n10476), .B2(n14924), .A(n10248), .ZN(P2_U3436) );
  OAI21_X1 U12819 ( .B1(n10251), .B2(n10250), .A(n10249), .ZN(n10835) );
  OAI21_X1 U12820 ( .B1(n10252), .B2(n10831), .A(n13316), .ZN(n10253) );
  NOR2_X1 U12821 ( .A1(n10253), .A2(n10559), .ZN(n10834) );
  XNOR2_X1 U12822 ( .A(n10255), .B(n10254), .ZN(n10258) );
  NAND2_X1 U12823 ( .A1(n13158), .A2(n13402), .ZN(n10257) );
  NAND2_X1 U12824 ( .A1(n8301), .A2(n13401), .ZN(n10256) );
  NAND2_X1 U12825 ( .A1(n10257), .A2(n10256), .ZN(n13049) );
  AOI21_X1 U12826 ( .B1(n10258), .B2(n13407), .A(n13049), .ZN(n10838) );
  INV_X1 U12827 ( .A(n10838), .ZN(n10259) );
  AOI211_X1 U12828 ( .C1(n14515), .C2(n10835), .A(n10834), .B(n10259), .ZN(
        n10478) );
  OAI22_X1 U12829 ( .A1(n13573), .A2(n10831), .B1(n14925), .B2(n7783), .ZN(
        n10260) );
  INV_X1 U12830 ( .A(n10260), .ZN(n10261) );
  OAI21_X1 U12831 ( .B1(n10478), .B2(n14924), .A(n10261), .ZN(P2_U3439) );
  INV_X1 U12832 ( .A(n10262), .ZN(n10263) );
  NAND2_X1 U12833 ( .A1(n13131), .A2(n10263), .ZN(n10265) );
  OAI211_X1 U12834 ( .C1(n14467), .C2(n10518), .A(n10265), .B(n10264), .ZN(
        n10271) );
  INV_X1 U12835 ( .A(n10266), .ZN(n10267) );
  AOI211_X1 U12836 ( .C1(n10269), .C2(n10268), .A(n14474), .B(n10267), .ZN(
        n10270) );
  AOI211_X1 U12837 ( .C1(n10487), .C2(n14479), .A(n10271), .B(n10270), .ZN(
        n10272) );
  INV_X1 U12838 ( .A(n10272), .ZN(P2_U3211) );
  XOR2_X1 U12839 ( .A(n10274), .B(n10273), .Z(n10280) );
  INV_X1 U12840 ( .A(n15046), .ZN(n10372) );
  NOR2_X1 U12841 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10275), .ZN(n14971) );
  AOI21_X1 U12842 ( .B1(n12524), .B2(n10372), .A(n14971), .ZN(n10277) );
  NAND2_X1 U12843 ( .A1(n12525), .A2(n15037), .ZN(n10276) );
  OAI211_X1 U12844 ( .C1(n10585), .C2(n12484), .A(n10277), .B(n10276), .ZN(
        n10278) );
  AOI21_X1 U12845 ( .B1(n15047), .B2(n12540), .A(n10278), .ZN(n10279) );
  OAI21_X1 U12846 ( .B1(n10280), .B2(n12507), .A(n10279), .ZN(P3_U3167) );
  INV_X1 U12847 ( .A(n10281), .ZN(n10284) );
  INV_X1 U12848 ( .A(n10288), .ZN(n10283) );
  INV_X1 U12849 ( .A(n10282), .ZN(n10576) );
  AOI21_X1 U12850 ( .B1(n10284), .B2(n10283), .A(n10576), .ZN(n10292) );
  NAND2_X1 U12851 ( .A1(n13117), .A2(n13153), .ZN(n10285) );
  NAND2_X1 U12852 ( .A1(P2_U3088), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n14813) );
  OAI211_X1 U12853 ( .C1(n14467), .C2(n10735), .A(n10285), .B(n14813), .ZN(
        n10286) );
  AOI21_X1 U12854 ( .B1(n10741), .B2(n14479), .A(n10286), .ZN(n10291) );
  NOR3_X1 U12855 ( .A1(n10288), .A2(n10287), .A3(n13124), .ZN(n10289) );
  INV_X1 U12856 ( .A(n14470), .ZN(n13116) );
  OAI21_X1 U12857 ( .B1(n10289), .B2(n13116), .A(n13155), .ZN(n10290) );
  OAI211_X1 U12858 ( .C1(n10292), .C2(n14474), .A(n10291), .B(n10290), .ZN(
        P2_U3193) );
  INV_X1 U12859 ( .A(n14221), .ZN(n10293) );
  NAND2_X1 U12860 ( .A1(n10294), .A2(n10293), .ZN(n13901) );
  AND2_X1 U12861 ( .A1(n10295), .A2(n6796), .ZN(n10296) );
  INV_X1 U12862 ( .A(n14677), .ZN(n10530) );
  NAND2_X1 U12863 ( .A1(n12341), .A2(n10528), .ZN(n10297) );
  NAND2_X1 U12864 ( .A1(n13778), .A2(n10298), .ZN(n12167) );
  OR2_X1 U12865 ( .A1(n13778), .A2(n14706), .ZN(n10299) );
  NAND2_X1 U12866 ( .A1(n14653), .A2(n14654), .ZN(n10301) );
  OR2_X1 U12867 ( .A1(n13776), .A2(n14664), .ZN(n10300) );
  OR2_X1 U12868 ( .A1(n12317), .A2(n10302), .ZN(n10305) );
  OR2_X1 U12869 ( .A1(n10388), .A2(n10303), .ZN(n10304) );
  XNOR2_X2 U12870 ( .A(n13775), .B(n14720), .ZN(n12342) );
  XNOR2_X1 U12871 ( .A(n10421), .B(n12342), .ZN(n14723) );
  INV_X1 U12872 ( .A(n12340), .ZN(n10661) );
  NAND2_X1 U12873 ( .A1(n10663), .A2(n10661), .ZN(n10307) );
  INV_X1 U12874 ( .A(n14654), .ZN(n10308) );
  NAND2_X1 U12875 ( .A1(n14655), .A2(n10308), .ZN(n10309) );
  XNOR2_X1 U12876 ( .A(n10383), .B(n12342), .ZN(n10312) );
  NAND2_X1 U12877 ( .A1(n14251), .A2(n11534), .ZN(n12141) );
  NAND2_X1 U12878 ( .A1(n9357), .A2(n12142), .ZN(n12329) );
  OR2_X1 U12879 ( .A1(n12186), .A2(n14678), .ZN(n10311) );
  NAND2_X1 U12880 ( .A1(n13776), .A2(n13897), .ZN(n10310) );
  NAND2_X1 U12881 ( .A1(n10311), .A2(n10310), .ZN(n10628) );
  AOI21_X1 U12882 ( .B1(n10312), .B2(n14694), .A(n10628), .ZN(n14721) );
  MUX2_X1 U12883 ( .A(n10313), .B(n14721), .S(n14113), .Z(n10317) );
  NAND2_X1 U12884 ( .A1(n14698), .A2(n14677), .ZN(n10666) );
  AOI211_X1 U12885 ( .C1(n14720), .C2(n14666), .A(n14663), .B(n14646), .ZN(
        n14719) );
  INV_X1 U12886 ( .A(n14720), .ZN(n10384) );
  OAI22_X1 U12887 ( .A1(n14089), .A2(n10384), .B1(n10631), .B2(n14659), .ZN(
        n10315) );
  AOI21_X1 U12888 ( .B1(n14719), .B2(n14669), .A(n10315), .ZN(n10316) );
  OAI211_X1 U12889 ( .C1(n14095), .C2(n14723), .A(n10317), .B(n10316), .ZN(
        P1_U3289) );
  OAI21_X1 U12890 ( .B1(n11049), .B2(P1_REG1_REG_11__SCAN_IN), .A(n10318), 
        .ZN(n10320) );
  INV_X1 U12891 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n15368) );
  AOI22_X1 U12892 ( .A1(n11194), .A2(P1_REG1_REG_12__SCAN_IN), .B1(n15368), 
        .B2(n10323), .ZN(n10319) );
  OAI21_X1 U12893 ( .B1(n10320), .B2(n10319), .A(n10791), .ZN(n10331) );
  OAI21_X1 U12894 ( .B1(n11063), .B2(n10322), .A(n10321), .ZN(n10326) );
  INV_X1 U12895 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n10324) );
  AOI22_X1 U12896 ( .A1(n11194), .A2(n10324), .B1(P1_REG2_REG_12__SCAN_IN), 
        .B2(n10323), .ZN(n10325) );
  NOR2_X1 U12897 ( .A1(n10325), .A2(n10326), .ZN(n10783) );
  AOI21_X1 U12898 ( .B1(n10326), .B2(n10325), .A(n10783), .ZN(n10329) );
  AND2_X1 U12899 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n13647) );
  AOI21_X1 U12900 ( .B1(n14604), .B2(P1_ADDR_REG_12__SCAN_IN), .A(n13647), 
        .ZN(n10328) );
  INV_X1 U12901 ( .A(n13862), .ZN(n14616) );
  NAND2_X1 U12902 ( .A1(n14616), .A2(n11194), .ZN(n10327) );
  OAI211_X1 U12903 ( .C1(n10329), .C2(n14619), .A(n10328), .B(n10327), .ZN(
        n10330) );
  AOI21_X1 U12904 ( .B1(n10331), .B2(n14614), .A(n10330), .ZN(n10332) );
  INV_X1 U12905 ( .A(n10332), .ZN(P1_U3255) );
  NAND2_X1 U12906 ( .A1(n13065), .A2(P2_U3947), .ZN(n10333) );
  OAI21_X1 U12907 ( .B1(n11772), .B2(P2_U3947), .A(n10333), .ZN(P2_U3559) );
  INV_X1 U12908 ( .A(n13131), .ZN(n13110) );
  OAI22_X1 U12909 ( .A1(n13110), .A2(n10334), .B1(n10426), .B2(n10822), .ZN(
        n10340) );
  INV_X1 U12910 ( .A(n13124), .ZN(n13105) );
  AOI22_X1 U12911 ( .A1(n13105), .A2(n10336), .B1(n10335), .B2(n14462), .ZN(
        n10338) );
  NOR2_X1 U12912 ( .A1(n10338), .A2(n10337), .ZN(n10339) );
  AOI211_X1 U12913 ( .C1(n10824), .C2(n14479), .A(n10340), .B(n10339), .ZN(
        n10341) );
  OAI21_X1 U12914 ( .B1(n10429), .B2(n14474), .A(n10341), .ZN(P2_U3194) );
  AOI22_X1 U12915 ( .A1(n13105), .A2(n13158), .B1(n14462), .B2(n10342), .ZN(
        n10345) );
  INV_X1 U12916 ( .A(n11890), .ZN(n10344) );
  NOR3_X1 U12917 ( .A1(n10345), .A2(n10344), .A3(n10343), .ZN(n10351) );
  INV_X1 U12918 ( .A(n10346), .ZN(n10347) );
  AOI22_X1 U12919 ( .A1(n13131), .A2(n10347), .B1(P2_REG3_REG_5__SCAN_IN), 
        .B2(P2_U3088), .ZN(n10349) );
  NAND2_X1 U12920 ( .A1(n14479), .A2(n10479), .ZN(n10348) );
  OAI211_X1 U12921 ( .C1(n14467), .C2(n10506), .A(n10349), .B(n10348), .ZN(
        n10350) );
  NOR2_X1 U12922 ( .A1(n10351), .A2(n10350), .ZN(n10352) );
  OAI21_X1 U12923 ( .B1(n10353), .B2(n14474), .A(n10352), .ZN(P2_U3199) );
  NOR2_X4 U12924 ( .A1(n10354), .A2(n14890), .ZN(n14929) );
  NAND2_X1 U12925 ( .A1(n13405), .A2(n13534), .ZN(n10356) );
  AND2_X1 U12926 ( .A1(n7753), .A2(n13402), .ZN(n10355) );
  AOI21_X1 U12927 ( .B1(n14882), .B2(n10356), .A(n10355), .ZN(n14879) );
  NOR2_X1 U12928 ( .A1(n10358), .A2(n10357), .ZN(n14875) );
  AOI21_X1 U12929 ( .B1(n14882), .B2(n14923), .A(n14875), .ZN(n10359) );
  AND2_X1 U12930 ( .A1(n14879), .A2(n10359), .ZN(n14895) );
  NAND2_X1 U12931 ( .A1(n14930), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n10360) );
  OAI21_X1 U12932 ( .B1(n14930), .B2(n14895), .A(n10360), .ZN(P2_U3499) );
  NAND2_X1 U12933 ( .A1(n15036), .A2(n15086), .ZN(n12004) );
  NAND2_X1 U12934 ( .A1(n10361), .A2(n11925), .ZN(n10362) );
  INV_X1 U12935 ( .A(n11988), .ZN(n10364) );
  AND2_X1 U12936 ( .A1(n15037), .A2(n15061), .ZN(n11989) );
  INV_X1 U12937 ( .A(n11989), .ZN(n10363) );
  NAND2_X1 U12938 ( .A1(n15060), .A2(n15059), .ZN(n10365) );
  NAND2_X1 U12939 ( .A1(n10365), .A2(n10364), .ZN(n15032) );
  NAND2_X1 U12940 ( .A1(n15053), .A2(n15046), .ZN(n11995) );
  NAND2_X1 U12941 ( .A1(n11999), .A2(n11995), .ZN(n11990) );
  NAND2_X1 U12942 ( .A1(n15032), .A2(n15035), .ZN(n10366) );
  XOR2_X1 U12943 ( .A(n10464), .B(n11924), .Z(n15087) );
  AOI22_X1 U12944 ( .A1(n15052), .A2(n12556), .B1(n15053), .B2(n15038), .ZN(
        n10378) );
  NAND2_X1 U12945 ( .A1(n15054), .A2(n12433), .ZN(n10367) );
  NAND2_X1 U12946 ( .A1(n10368), .A2(n10367), .ZN(n15051) );
  INV_X1 U12947 ( .A(n15059), .ZN(n11926) );
  NAND2_X1 U12948 ( .A1(n15051), .A2(n11926), .ZN(n10371) );
  NAND2_X1 U12949 ( .A1(n15037), .A2(n10369), .ZN(n10370) );
  NAND2_X1 U12950 ( .A1(n10371), .A2(n10370), .ZN(n15034) );
  OR2_X1 U12951 ( .A1(n15034), .A2(n15035), .ZN(n10375) );
  INV_X1 U12952 ( .A(n10375), .ZN(n15033) );
  NOR2_X1 U12953 ( .A1(n15053), .A2(n10372), .ZN(n10373) );
  OAI21_X1 U12954 ( .B1(n15033), .B2(n10373), .A(n11924), .ZN(n10376) );
  NOR2_X1 U12955 ( .A1(n11924), .A2(n10373), .ZN(n10374) );
  NAND3_X1 U12956 ( .A1(n10376), .A2(n15056), .A3(n10466), .ZN(n10377) );
  OAI211_X1 U12957 ( .C1(n15087), .C2(n15039), .A(n10378), .B(n10377), .ZN(
        n15089) );
  NAND2_X1 U12958 ( .A1(n15089), .A2(n15049), .ZN(n10382) );
  INV_X1 U12959 ( .A(n15086), .ZN(n12523) );
  INV_X1 U12960 ( .A(n12526), .ZN(n10379) );
  OAI22_X1 U12961 ( .A1(n15049), .A2(n15325), .B1(n10379), .B2(n12868), .ZN(
        n10380) );
  AOI21_X1 U12962 ( .B1(n14423), .B2(n12523), .A(n10380), .ZN(n10381) );
  OAI211_X1 U12963 ( .C1(n15087), .C2(n10821), .A(n10382), .B(n10381), .ZN(
        P3_U3227) );
  NAND2_X1 U12964 ( .A1(n10383), .A2(n12342), .ZN(n10386) );
  OR2_X1 U12965 ( .A1(n13775), .A2(n10384), .ZN(n10385) );
  INV_X2 U12966 ( .A(n12317), .ZN(n11535) );
  AOI22_X1 U12967 ( .A1(n11535), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n11533), 
        .B2(n10387), .ZN(n10391) );
  INV_X2 U12968 ( .A(n10388), .ZN(n10677) );
  NAND2_X1 U12969 ( .A1(n10389), .A2(n10677), .ZN(n10390) );
  AND2_X1 U12970 ( .A1(n12186), .A2(n14649), .ZN(n10392) );
  NAND2_X1 U12971 ( .A1(n11783), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n10399) );
  INV_X1 U12972 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n10393) );
  OR2_X1 U12973 ( .A1(n11784), .A2(n10393), .ZN(n10398) );
  OR2_X1 U12974 ( .A1(n10394), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n10395) );
  NAND2_X1 U12975 ( .A1(n10407), .A2(n10395), .ZN(n10604) );
  OR2_X1 U12976 ( .A1(n11600), .A2(n10604), .ZN(n10397) );
  OR2_X1 U12977 ( .A1(n6526), .A2(n9709), .ZN(n10396) );
  NAND4_X1 U12978 ( .A1(n10399), .A2(n10398), .A3(n10397), .A4(n10396), .ZN(
        n13774) );
  NAND2_X1 U12979 ( .A1(n10400), .A2(n10677), .ZN(n10403) );
  AOI22_X1 U12980 ( .A1(n11535), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n11533), 
        .B2(n10401), .ZN(n10402) );
  NAND2_X1 U12981 ( .A1(n10403), .A2(n10402), .ZN(n12194) );
  XNOR2_X1 U12982 ( .A(n13774), .B(n12194), .ZN(n12344) );
  XNOR2_X1 U12983 ( .A(n10698), .B(n12344), .ZN(n14738) );
  OR2_X1 U12984 ( .A1(n14674), .A2(n14737), .ZN(n14052) );
  INV_X1 U12985 ( .A(n14636), .ZN(n10404) );
  AOI211_X1 U12986 ( .C1(n12194), .C2(n14647), .A(n14663), .B(n10404), .ZN(
        n14735) );
  NOR2_X1 U12987 ( .A1(n14089), .A2(n7261), .ZN(n10419) );
  OR2_X1 U12988 ( .A1(n12186), .A2(n13674), .ZN(n10415) );
  NAND2_X1 U12989 ( .A1(n12321), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n10413) );
  OR2_X1 U12990 ( .A1(n6526), .A2(n10405), .ZN(n10412) );
  NAND2_X1 U12991 ( .A1(n10407), .A2(n10406), .ZN(n10408) );
  NAND2_X1 U12992 ( .A1(n10705), .A2(n10408), .ZN(n14633) );
  OR2_X1 U12993 ( .A1(n11600), .A2(n14633), .ZN(n10411) );
  OR2_X1 U12994 ( .A1(n6540), .A2(n10409), .ZN(n10410) );
  NAND4_X1 U12995 ( .A1(n10413), .A2(n10412), .A3(n10411), .A4(n10410), .ZN(
        n13773) );
  NAND2_X1 U12996 ( .A1(n13773), .A2(n13732), .ZN(n10414) );
  NAND2_X1 U12997 ( .A1(n10415), .A2(n10414), .ZN(n14733) );
  INV_X1 U12998 ( .A(n14733), .ZN(n10416) );
  MUX2_X1 U12999 ( .A(n10416), .B(n9709), .S(n14674), .Z(n10417) );
  OAI21_X1 U13000 ( .B1(n14659), .B2(n10604), .A(n10417), .ZN(n10418) );
  AOI211_X1 U13001 ( .C1(n14735), .C2(n14669), .A(n10419), .B(n10418), .ZN(
        n10425) );
  INV_X1 U13002 ( .A(n12342), .ZN(n10420) );
  OR2_X1 U13003 ( .A1(n13775), .A2(n14720), .ZN(n10422) );
  INV_X1 U13004 ( .A(n12186), .ZN(n12188) );
  XNOR2_X1 U13005 ( .A(n12188), .B(n14649), .ZN(n12343) );
  INV_X1 U13006 ( .A(n12343), .ZN(n14641) );
  NAND2_X1 U13007 ( .A1(n12186), .A2(n12187), .ZN(n10423) );
  XNOR2_X1 U13008 ( .A(n10675), .B(n10697), .ZN(n14740) );
  NAND2_X1 U13009 ( .A1(n14740), .A2(n14676), .ZN(n10424) );
  OAI211_X1 U13010 ( .C1(n14738), .C2(n14052), .A(n10425), .B(n10424), .ZN(
        P1_U3287) );
  OAI22_X1 U13011 ( .A1(n13110), .A2(n10427), .B1(n10426), .B2(n13161), .ZN(
        n10434) );
  AOI22_X1 U13012 ( .A1(n13105), .A2(n7753), .B1(n14462), .B2(n10428), .ZN(
        n10432) );
  INV_X1 U13013 ( .A(n10429), .ZN(n10431) );
  NOR3_X1 U13014 ( .A1(n10432), .A2(n10431), .A3(n10430), .ZN(n10433) );
  AOI211_X1 U13015 ( .C1(n10474), .C2(n14479), .A(n10434), .B(n10433), .ZN(
        n10435) );
  OAI21_X1 U13016 ( .B1(n10436), .B2(n14474), .A(n10435), .ZN(P2_U3209) );
  OR2_X1 U13017 ( .A1(n10438), .A2(n10437), .ZN(n10448) );
  NAND2_X1 U13018 ( .A1(n10450), .A2(n10448), .ZN(n10442) );
  NAND2_X1 U13019 ( .A1(n13775), .A2(n6720), .ZN(n10441) );
  INV_X2 U13020 ( .A(n11701), .ZN(n11777) );
  NAND2_X1 U13021 ( .A1(n11777), .A2(n14720), .ZN(n10440) );
  NAND2_X1 U13022 ( .A1(n10441), .A2(n10440), .ZN(n10446) );
  NAND2_X1 U13023 ( .A1(n13775), .A2(n11777), .ZN(n10444) );
  NAND2_X1 U13024 ( .A1(n14720), .A2(n11778), .ZN(n10443) );
  NAND2_X1 U13025 ( .A1(n10444), .A2(n10443), .ZN(n10445) );
  XNOR2_X1 U13026 ( .A(n10445), .B(n11745), .ZN(n10634) );
  INV_X1 U13027 ( .A(n10446), .ZN(n10447) );
  AND2_X1 U13028 ( .A1(n10448), .A2(n10447), .ZN(n10449) );
  OAI22_X1 U13029 ( .A1(n12186), .A2(n11701), .B1(n12187), .B2(n11702), .ZN(
        n10451) );
  XNOR2_X1 U13030 ( .A(n10451), .B(n11775), .ZN(n10454) );
  OAI22_X1 U13031 ( .A1(n12186), .A2(n11700), .B1(n12187), .B2(n11701), .ZN(
        n10453) );
  OR2_X1 U13032 ( .A1(n10454), .A2(n10453), .ZN(n10591) );
  INV_X1 U13033 ( .A(n10591), .ZN(n10455) );
  AND2_X1 U13034 ( .A1(n10454), .A2(n10453), .ZN(n10590) );
  NOR2_X1 U13035 ( .A1(n10455), .A2(n10590), .ZN(n10456) );
  XNOR2_X1 U13036 ( .A(n10592), .B(n10456), .ZN(n10463) );
  AND2_X1 U13037 ( .A1(n14649), .A2(n14742), .ZN(n14728) );
  NAND2_X1 U13038 ( .A1(n13774), .A2(n13732), .ZN(n10458) );
  NAND2_X1 U13039 ( .A1(n13775), .A2(n13897), .ZN(n10457) );
  NAND2_X1 U13040 ( .A1(n10458), .A2(n10457), .ZN(n14726) );
  NAND2_X1 U13041 ( .A1(n14537), .A2(n14726), .ZN(n10459) );
  OAI211_X1 U13042 ( .C1(n14542), .C2(n14644), .A(n10460), .B(n10459), .ZN(
        n10461) );
  AOI21_X1 U13043 ( .B1(n14728), .B2(n13601), .A(n10461), .ZN(n10462) );
  OAI21_X1 U13044 ( .B1(n10463), .B2(n13727), .A(n10462), .ZN(P1_U3227) );
  XNOR2_X1 U13045 ( .A(n10623), .B(n7134), .ZN(n15091) );
  NAND2_X1 U13046 ( .A1(n15036), .A2(n12523), .ZN(n10465) );
  NAND2_X1 U13047 ( .A1(n10466), .A2(n10465), .ZN(n10612) );
  XNOR2_X1 U13048 ( .A(n10612), .B(n12003), .ZN(n10467) );
  NAND2_X1 U13049 ( .A1(n10467), .A2(n15056), .ZN(n10469) );
  AOI22_X1 U13050 ( .A1(n15038), .A2(n15036), .B1(n12555), .B2(n15052), .ZN(
        n10468) );
  OAI211_X1 U13051 ( .C1(n15091), .C2(n15039), .A(n10469), .B(n10468), .ZN(
        n15093) );
  NAND2_X1 U13052 ( .A1(n15093), .A2(n15049), .ZN(n10473) );
  OR2_X1 U13053 ( .A1(n10584), .A2(n15099), .ZN(n15090) );
  INV_X1 U13054 ( .A(n10470), .ZN(n10589) );
  OAI22_X1 U13055 ( .A1(n11177), .A2(n15090), .B1(n10589), .B2(n12868), .ZN(
        n10471) );
  AOI21_X1 U13056 ( .B1(n15066), .B2(P3_REG2_REG_7__SCAN_IN), .A(n10471), .ZN(
        n10472) );
  OAI211_X1 U13057 ( .C1(n15091), .C2(n10821), .A(n10473), .B(n10472), .ZN(
        P3_U3226) );
  AOI22_X1 U13058 ( .A1(n13465), .A2(n10474), .B1(n14930), .B2(
        P2_REG1_REG_2__SCAN_IN), .ZN(n10475) );
  OAI21_X1 U13059 ( .B1(n10476), .B2(n14930), .A(n10475), .ZN(P2_U3501) );
  AOI22_X1 U13060 ( .A1(n13465), .A2(n13050), .B1(n14930), .B2(
        P2_REG1_REG_3__SCAN_IN), .ZN(n10477) );
  OAI21_X1 U13061 ( .B1(n10478), .B2(n14930), .A(n10477), .ZN(P2_U3502) );
  AOI22_X1 U13062 ( .A1(n13465), .A2(n10479), .B1(n14930), .B2(
        P2_REG1_REG_5__SCAN_IN), .ZN(n10480) );
  OAI21_X1 U13063 ( .B1(n10481), .B2(n14930), .A(n10480), .ZN(P2_U3504) );
  AOI22_X1 U13064 ( .A1(n13465), .A2(n10824), .B1(n14930), .B2(
        P2_REG1_REG_1__SCAN_IN), .ZN(n10482) );
  OAI21_X1 U13065 ( .B1(n10483), .B2(n14930), .A(n10482), .ZN(P2_U3500) );
  AOI22_X1 U13066 ( .A1(n13465), .A2(n10484), .B1(n14930), .B2(
        P2_REG1_REG_7__SCAN_IN), .ZN(n10485) );
  OAI21_X1 U13067 ( .B1(n10486), .B2(n14930), .A(n10485), .ZN(P2_U3506) );
  AOI22_X1 U13068 ( .A1(n13465), .A2(n10487), .B1(n14930), .B2(
        P2_REG1_REG_6__SCAN_IN), .ZN(n10488) );
  OAI21_X1 U13069 ( .B1(n10489), .B2(n14930), .A(n10488), .ZN(P2_U3505) );
  INV_X1 U13070 ( .A(n10490), .ZN(n10499) );
  NAND2_X1 U13071 ( .A1(n10491), .A2(n13429), .ZN(n10498) );
  NOR2_X1 U13072 ( .A1(n13414), .A2(n10492), .ZN(n10495) );
  OAI22_X1 U13073 ( .A1(n14884), .A2(n7850), .B1(n10493), .B2(n14877), .ZN(
        n10494) );
  AOI211_X1 U13074 ( .C1(n10496), .C2(n13444), .A(n10495), .B(n10494), .ZN(
        n10497) );
  OAI211_X1 U13075 ( .C1(n10499), .C2(n13393), .A(n10498), .B(n10497), .ZN(
        P2_U3258) );
  NAND2_X1 U13076 ( .A1(n10500), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10501) );
  XNOR2_X1 U13077 ( .A(n10501), .B(P1_IR_REG_18__SCAN_IN), .ZN(n13858) );
  INV_X1 U13078 ( .A(n13858), .ZN(n13852) );
  INV_X1 U13079 ( .A(n11520), .ZN(n10504) );
  OAI222_X1 U13080 ( .A1(P1_U3086), .A2(n13852), .B1(n11860), .B2(n10504), 
        .C1(n10502), .C2(n14247), .ZN(P1_U3337) );
  OAI222_X1 U13081 ( .A1(P2_U3088), .A2(n6948), .B1(n13596), .B2(n10504), .C1(
        n10503), .C2(n13594), .ZN(P2_U3309) );
  INV_X1 U13082 ( .A(n10505), .ZN(n10513) );
  OAI22_X1 U13083 ( .A1(n14884), .A2(n9532), .B1(n10506), .B2(n14877), .ZN(
        n10508) );
  NOR2_X1 U13084 ( .A1(n13414), .A2(n6904), .ZN(n10507) );
  AOI211_X1 U13085 ( .C1(n10509), .C2(n13444), .A(n10508), .B(n10507), .ZN(
        n10512) );
  NAND2_X1 U13086 ( .A1(n10510), .A2(n13429), .ZN(n10511) );
  OAI211_X1 U13087 ( .C1(n13393), .C2(n10513), .A(n10512), .B(n10511), .ZN(
        P2_U3260) );
  INV_X1 U13088 ( .A(n10514), .ZN(n10524) );
  INV_X1 U13089 ( .A(n10515), .ZN(n10516) );
  MUX2_X1 U13090 ( .A(n10517), .B(n10516), .S(n14884), .Z(n10523) );
  OAI22_X1 U13091 ( .A1(n13414), .A2(n10519), .B1(n14877), .B2(n10518), .ZN(
        n10520) );
  AOI21_X1 U13092 ( .B1(n13444), .B2(n10521), .A(n10520), .ZN(n10522) );
  OAI211_X1 U13093 ( .C1(n13393), .C2(n10524), .A(n10523), .B(n10522), .ZN(
        P2_U3259) );
  OR2_X1 U13094 ( .A1(n12159), .A2(n13868), .ZN(n12147) );
  NOR2_X1 U13095 ( .A1(n14674), .A2(n12147), .ZN(n14670) );
  INV_X1 U13096 ( .A(n10525), .ZN(n10526) );
  NOR2_X1 U13097 ( .A1(n14674), .A2(n14691), .ZN(n10527) );
  OR2_X1 U13098 ( .A1(n14670), .A2(n10527), .ZN(n13970) );
  INV_X1 U13099 ( .A(n13970), .ZN(n14066) );
  XOR2_X1 U13100 ( .A(n6726), .B(n10528), .Z(n14690) );
  OAI22_X1 U13101 ( .A1(n14113), .A2(n9358), .B1(n10529), .B2(n14659), .ZN(
        n10537) );
  NAND2_X1 U13102 ( .A1(n10530), .A2(n12163), .ZN(n10531) );
  NAND2_X1 U13103 ( .A1(n10666), .A2(n10531), .ZN(n10533) );
  XNOR2_X1 U13104 ( .A(n10533), .B(n6770), .ZN(n14693) );
  NAND2_X1 U13105 ( .A1(n14675), .A2(n14693), .ZN(n10535) );
  OR2_X1 U13106 ( .A1(n6726), .A2(n10539), .ZN(n10532) );
  AOI21_X1 U13107 ( .B1(n10532), .B2(n14694), .A(n13897), .ZN(n14692) );
  INV_X1 U13108 ( .A(n10533), .ZN(n10534) );
  NAND2_X1 U13109 ( .A1(n10534), .A2(n14109), .ZN(n14696) );
  OAI22_X1 U13110 ( .A1(n10535), .A2(n14692), .B1(n14117), .B2(n14696), .ZN(
        n10536) );
  AOI211_X1 U13111 ( .C1(n14662), .C2(n12163), .A(n10537), .B(n10536), .ZN(
        n10541) );
  OAI22_X1 U13112 ( .A1(n14692), .A2(n10539), .B1(n10538), .B2(n14678), .ZN(
        n14699) );
  INV_X1 U13113 ( .A(n14674), .ZN(n14680) );
  NAND2_X1 U13114 ( .A1(n14699), .A2(n14680), .ZN(n10540) );
  OAI211_X1 U13115 ( .C1(n14066), .C2(n14690), .A(n10541), .B(n10540), .ZN(
        P1_U3292) );
  XNOR2_X1 U13116 ( .A(n10542), .B(n10543), .ZN(n10744) );
  NAND2_X1 U13117 ( .A1(n13429), .A2(n14883), .ZN(n13415) );
  XNOR2_X1 U13118 ( .A(n10544), .B(n10543), .ZN(n10548) );
  INV_X1 U13119 ( .A(n13401), .ZN(n13536) );
  OAI22_X1 U13120 ( .A1(n10546), .A2(n13536), .B1(n10545), .B2(n13538), .ZN(
        n10547) );
  AOI21_X1 U13121 ( .B1(n10548), .B2(n13407), .A(n10547), .ZN(n10549) );
  OAI21_X1 U13122 ( .B1(n10744), .B2(n13405), .A(n10549), .ZN(n10745) );
  NAND2_X1 U13123 ( .A1(n10745), .A2(n13429), .ZN(n10555) );
  INV_X1 U13124 ( .A(n10550), .ZN(n10776) );
  AOI211_X1 U13125 ( .C1(n10750), .C2(n10737), .A(n13269), .B(n10776), .ZN(
        n10746) );
  INV_X1 U13126 ( .A(n10750), .ZN(n10551) );
  NOR2_X1 U13127 ( .A1(n10551), .A2(n13414), .ZN(n10553) );
  OAI22_X1 U13128 ( .A1(n14884), .A2(n9885), .B1(n10572), .B2(n14877), .ZN(
        n10552) );
  AOI211_X1 U13129 ( .C1(n10746), .C2(n13444), .A(n10553), .B(n10552), .ZN(
        n10554) );
  OAI211_X1 U13130 ( .C1(n10744), .C2(n13415), .A(n10555), .B(n10554), .ZN(
        P2_U3256) );
  OAI21_X1 U13131 ( .B1(n10558), .B2(n10557), .A(n10556), .ZN(n14905) );
  INV_X1 U13132 ( .A(n14905), .ZN(n14902) );
  INV_X1 U13133 ( .A(n10559), .ZN(n10561) );
  AOI211_X1 U13134 ( .C1(n14898), .C2(n10561), .A(n13269), .B(n6902), .ZN(
        n14897) );
  OAI22_X1 U13135 ( .A1(n13414), .A2(n11884), .B1(n11883), .B2(n14877), .ZN(
        n10562) );
  AOI21_X1 U13136 ( .B1(n13444), .B2(n14897), .A(n10562), .ZN(n10569) );
  XNOR2_X1 U13137 ( .A(n10564), .B(n10563), .ZN(n10566) );
  AOI22_X1 U13138 ( .A1(n13401), .A2(n13159), .B1(n13157), .B2(n13402), .ZN(
        n11882) );
  INV_X1 U13139 ( .A(n11882), .ZN(n10565) );
  AOI21_X1 U13140 ( .B1(n10566), .B2(n13407), .A(n10565), .ZN(n14896) );
  MUX2_X1 U13141 ( .A(n10567), .B(n14896), .S(n14884), .Z(n10568) );
  OAI211_X1 U13142 ( .C1(n14902), .C2(n13393), .A(n10569), .B(n10568), .ZN(
        P2_U3261) );
  AOI22_X1 U13143 ( .A1(n13116), .A2(n13154), .B1(n13117), .B2(n13152), .ZN(
        n10571) );
  OAI211_X1 U13144 ( .C1(n10572), .C2(n14467), .A(n10571), .B(n10570), .ZN(
        n10578) );
  AOI22_X1 U13145 ( .A1(n13105), .A2(n13154), .B1(n14462), .B2(n10573), .ZN(
        n10575) );
  NOR3_X1 U13146 ( .A1(n10576), .A2(n10575), .A3(n10574), .ZN(n10577) );
  AOI211_X1 U13147 ( .C1(n10750), .C2(n14479), .A(n10578), .B(n10577), .ZN(
        n10579) );
  OAI21_X1 U13148 ( .B1(n10580), .B2(n14474), .A(n10579), .ZN(P2_U3203) );
  OAI211_X1 U13149 ( .C1(n10583), .C2(n10582), .A(n10581), .B(n12533), .ZN(
        n10588) );
  INV_X1 U13150 ( .A(n10584), .ZN(n10613) );
  INV_X1 U13151 ( .A(P3_REG3_REG_7__SCAN_IN), .ZN(n15354) );
  NOR2_X1 U13152 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15354), .ZN(n15000) );
  OAI22_X1 U13153 ( .A1(n12537), .A2(n10585), .B1(n10919), .B2(n12484), .ZN(
        n10586) );
  AOI211_X1 U13154 ( .C1(n10613), .C2(n12524), .A(n15000), .B(n10586), .ZN(
        n10587) );
  OAI211_X1 U13155 ( .C1(n10589), .C2(n12486), .A(n10588), .B(n10587), .ZN(
        P3_U3153) );
  NAND2_X1 U13156 ( .A1(n13774), .A2(n11777), .ZN(n10594) );
  NAND2_X1 U13157 ( .A1(n12194), .A2(n11778), .ZN(n10593) );
  NAND2_X1 U13158 ( .A1(n10594), .A2(n10593), .ZN(n10595) );
  XNOR2_X1 U13159 ( .A(n10595), .B(n11775), .ZN(n10601) );
  INV_X1 U13160 ( .A(n10601), .ZN(n10599) );
  NAND2_X1 U13161 ( .A1(n13774), .A2(n6720), .ZN(n10597) );
  NAND2_X1 U13162 ( .A1(n12194), .A2(n11777), .ZN(n10596) );
  NAND2_X1 U13163 ( .A1(n10597), .A2(n10596), .ZN(n10600) );
  INV_X1 U13164 ( .A(n10600), .ZN(n10598) );
  NAND2_X1 U13165 ( .A1(n10599), .A2(n10598), .ZN(n10958) );
  NAND2_X1 U13166 ( .A1(n10601), .A2(n10600), .ZN(n10956) );
  NAND2_X1 U13167 ( .A1(n10958), .A2(n10956), .ZN(n10602) );
  XNOR2_X1 U13168 ( .A(n10957), .B(n10602), .ZN(n10607) );
  NOR2_X1 U13169 ( .A1(n7261), .A2(n14767), .ZN(n14734) );
  AOI22_X1 U13170 ( .A1(n14537), .A2(n14733), .B1(P1_REG3_REG_6__SCAN_IN), 
        .B2(P1_U3086), .ZN(n10603) );
  OAI21_X1 U13171 ( .B1(n10604), .B2(n14542), .A(n10603), .ZN(n10605) );
  AOI21_X1 U13172 ( .B1(n14734), .B2(n13601), .A(n10605), .ZN(n10606) );
  OAI21_X1 U13173 ( .B1(n10607), .B2(n13727), .A(n10606), .ZN(P1_U3239) );
  INV_X1 U13174 ( .A(n10608), .ZN(n10610) );
  OAI222_X1 U13175 ( .A1(P3_U3151), .A2(n10611), .B1(n14370), .B2(n10610), 
        .C1(n10609), .C2(n14368), .ZN(P3_U3275) );
  NAND2_X1 U13176 ( .A1(n10612), .A2(n7134), .ZN(n10615) );
  NAND2_X1 U13177 ( .A1(n12556), .A2(n10613), .ZN(n10614) );
  NAND2_X1 U13178 ( .A1(n12555), .A2(n10756), .ZN(n12012) );
  NAND2_X1 U13179 ( .A1(n12013), .A2(n12012), .ZN(n12007) );
  NAND2_X1 U13180 ( .A1(n10616), .A2(n11928), .ZN(n10617) );
  NAND2_X1 U13181 ( .A1(n10814), .A2(n10617), .ZN(n10618) );
  NAND2_X1 U13182 ( .A1(n10618), .A2(n15056), .ZN(n10620) );
  AOI22_X1 U13183 ( .A1(n15038), .A2(n12556), .B1(n12554), .B2(n15052), .ZN(
        n10619) );
  AND2_X1 U13184 ( .A1(n10620), .A2(n10619), .ZN(n15098) );
  OR2_X1 U13185 ( .A1(n10756), .A2(n15099), .ZN(n15096) );
  INV_X1 U13186 ( .A(n10621), .ZN(n10763) );
  OAI22_X1 U13187 ( .A1(n11177), .A2(n15096), .B1(n10763), .B2(n12868), .ZN(
        n10622) );
  AOI21_X1 U13188 ( .B1(P3_REG2_REG_8__SCAN_IN), .B2(n15066), .A(n10622), .ZN(
        n10627) );
  XNOR2_X1 U13189 ( .A(n10810), .B(n11928), .ZN(n15095) );
  OR2_X1 U13190 ( .A1(n15066), .A2(n15039), .ZN(n10625) );
  INV_X1 U13191 ( .A(n12873), .ZN(n15063) );
  NAND2_X1 U13192 ( .A1(n15095), .A2(n15063), .ZN(n10626) );
  OAI211_X1 U13193 ( .C1(n15098), .C2(n15066), .A(n10627), .B(n10626), .ZN(
        P3_U3225) );
  NAND2_X1 U13194 ( .A1(n14537), .A2(n10628), .ZN(n10629) );
  OAI211_X1 U13195 ( .C1(n14542), .C2(n10631), .A(n10630), .B(n10629), .ZN(
        n10638) );
  NAND2_X1 U13196 ( .A1(n10633), .A2(n10632), .ZN(n10635) );
  XNOR2_X1 U13197 ( .A(n10635), .B(n10634), .ZN(n10636) );
  NOR2_X1 U13198 ( .A1(n10636), .A2(n13727), .ZN(n10637) );
  AOI211_X1 U13199 ( .C1(n14533), .C2(n14720), .A(n10638), .B(n10637), .ZN(
        n10639) );
  INV_X1 U13200 ( .A(n10639), .ZN(P1_U3230) );
  OAI21_X1 U13201 ( .B1(n10641), .B2(n11090), .A(n11084), .ZN(n10643) );
  INV_X1 U13202 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n10642) );
  AOI21_X1 U13203 ( .B1(n10643), .B2(n10642), .A(n11085), .ZN(n10660) );
  INV_X1 U13204 ( .A(n10644), .ZN(n10645) );
  AOI22_X1 U13205 ( .A1(n10647), .A2(n10646), .B1(n10651), .B2(n10645), .ZN(
        n11093) );
  MUX2_X1 U13206 ( .A(P3_REG2_REG_9__SCAN_IN), .B(P3_REG1_REG_9__SCAN_IN), .S(
        n12670), .Z(n11091) );
  XOR2_X1 U13207 ( .A(n10648), .B(n11091), .Z(n11092) );
  XNOR2_X1 U13208 ( .A(n11093), .B(n11092), .ZN(n10658) );
  NOR2_X1 U13209 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10649), .ZN(n10921) );
  AOI21_X1 U13210 ( .B1(n15001), .B2(P3_ADDR_REG_9__SCAN_IN), .A(n10921), .ZN(
        n10650) );
  OAI21_X1 U13211 ( .B1(n12701), .B2(n11090), .A(n10650), .ZN(n10657) );
  OAI21_X1 U13212 ( .B1(n10653), .B2(n11090), .A(n11099), .ZN(n10654) );
  INV_X1 U13213 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n15127) );
  AOI21_X1 U13214 ( .B1(n10654), .B2(n15127), .A(n11100), .ZN(n10655) );
  NOR2_X1 U13215 ( .A1(n10655), .A2(n15018), .ZN(n10656) );
  AOI211_X1 U13216 ( .C1(n15015), .C2(n10658), .A(n10657), .B(n10656), .ZN(
        n10659) );
  OAI21_X1 U13217 ( .B1(n10660), .B2(n15023), .A(n10659), .ZN(P3_U3191) );
  XNOR2_X1 U13218 ( .A(n10662), .B(n10661), .ZN(n14708) );
  XNOR2_X1 U13219 ( .A(n12340), .B(n10663), .ZN(n10665) );
  OAI21_X1 U13220 ( .B1(n10665), .B2(n14737), .A(n10664), .ZN(n14704) );
  AOI21_X1 U13221 ( .B1(n10666), .B2(n14706), .A(n14663), .ZN(n10667) );
  NAND2_X1 U13222 ( .A1(n10667), .A2(n14665), .ZN(n14703) );
  NAND2_X1 U13223 ( .A1(n14662), .A2(n14706), .ZN(n10669) );
  AOI22_X1 U13224 ( .A1(n14674), .A2(P1_REG2_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(n14673), .ZN(n10668) );
  OAI211_X1 U13225 ( .C1(n14703), .C2(n14117), .A(n10669), .B(n10668), .ZN(
        n10670) );
  AOI21_X1 U13226 ( .B1(n14680), .B2(n14704), .A(n10670), .ZN(n10671) );
  OAI21_X1 U13227 ( .B1(n14066), .B2(n14708), .A(n10671), .ZN(P1_U3291) );
  INV_X1 U13228 ( .A(n11532), .ZN(n10673) );
  OAI222_X1 U13229 ( .A1(n13868), .A2(P1_U3086), .B1(n11860), .B2(n10673), 
        .C1(n10672), .C2(n14247), .ZN(P1_U3336) );
  OAI222_X1 U13230 ( .A1(n13594), .A2(n10674), .B1(n13596), .B2(n10673), .C1(
        n13229), .C2(P2_U3088), .ZN(P2_U3308) );
  OR2_X1 U13231 ( .A1(n13774), .A2(n12194), .ZN(n10676) );
  NAND2_X1 U13232 ( .A1(n10678), .A2(n10677), .ZN(n10681) );
  AOI22_X1 U13233 ( .A1(n11535), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n11533), 
        .B2(n10679), .ZN(n10680) );
  INV_X1 U13234 ( .A(n13773), .ZN(n10699) );
  NAND2_X1 U13235 ( .A1(n14629), .A2(n12347), .ZN(n10683) );
  OR2_X1 U13236 ( .A1(n14743), .A2(n13773), .ZN(n10682) );
  NAND2_X1 U13237 ( .A1(n10684), .A2(n10677), .ZN(n10687) );
  AOI22_X1 U13238 ( .A1(n11535), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n11533), 
        .B2(n10685), .ZN(n10686) );
  NAND2_X1 U13239 ( .A1(n10687), .A2(n10686), .ZN(n12205) );
  NAND2_X1 U13240 ( .A1(n12321), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n10692) );
  OR2_X1 U13241 ( .A1(n6539), .A2(n10688), .ZN(n10691) );
  XNOR2_X1 U13242 ( .A(n10705), .B(n15221), .ZN(n10991) );
  OR2_X1 U13243 ( .A1(n11600), .A2(n10991), .ZN(n10690) );
  OR2_X1 U13244 ( .A1(n6526), .A2(n9832), .ZN(n10689) );
  NAND4_X1 U13245 ( .A1(n10692), .A2(n10691), .A3(n10690), .A4(n10689), .ZN(
        n13772) );
  INV_X1 U13246 ( .A(n13772), .ZN(n10693) );
  OR2_X1 U13247 ( .A1(n12205), .A2(n10693), .ZN(n10875) );
  NAND2_X1 U13248 ( .A1(n12205), .A2(n10693), .ZN(n10694) );
  XNOR2_X1 U13249 ( .A(n10868), .B(n12346), .ZN(n14750) );
  INV_X1 U13250 ( .A(n14750), .ZN(n10722) );
  INV_X1 U13251 ( .A(n13774), .ZN(n10695) );
  NAND2_X1 U13252 ( .A1(n10695), .A2(n12194), .ZN(n10696) );
  INV_X1 U13253 ( .A(n12347), .ZN(n14628) );
  NAND2_X1 U13254 ( .A1(n14627), .A2(n14628), .ZN(n14626) );
  NAND2_X1 U13255 ( .A1(n14743), .A2(n10699), .ZN(n10700) );
  NAND2_X1 U13256 ( .A1(n10701), .A2(n12346), .ZN(n10702) );
  NAND3_X1 U13257 ( .A1(n10876), .A2(n14694), .A3(n10702), .ZN(n10715) );
  NAND2_X1 U13258 ( .A1(n13773), .A2(n13897), .ZN(n10713) );
  NAND2_X1 U13259 ( .A1(n12321), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n10711) );
  OR2_X1 U13260 ( .A1(n6526), .A2(n10703), .ZN(n10710) );
  INV_X1 U13261 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n10704) );
  OAI21_X1 U13262 ( .B1(n10705), .B2(n15221), .A(n10704), .ZN(n10706) );
  NAND2_X1 U13263 ( .A1(n10706), .A2(n10877), .ZN(n11154) );
  OR2_X1 U13264 ( .A1(n11600), .A2(n11154), .ZN(n10709) );
  OR2_X1 U13265 ( .A1(n6540), .A2(n10707), .ZN(n10708) );
  NAND4_X1 U13266 ( .A1(n10711), .A2(n10710), .A3(n10709), .A4(n10708), .ZN(
        n13771) );
  NAND2_X1 U13267 ( .A1(n13771), .A2(n13732), .ZN(n10712) );
  NAND2_X1 U13268 ( .A1(n10713), .A2(n10712), .ZN(n10989) );
  INV_X1 U13269 ( .A(n10989), .ZN(n10714) );
  NAND2_X1 U13270 ( .A1(n10715), .A2(n10714), .ZN(n14756) );
  INV_X1 U13271 ( .A(n12205), .ZN(n10716) );
  OAI21_X1 U13272 ( .B1(n14635), .B2(n10716), .A(n14109), .ZN(n10717) );
  OR2_X1 U13273 ( .A1(n10717), .A2(n10890), .ZN(n14753) );
  OAI22_X1 U13274 ( .A1(n14113), .A2(n9832), .B1(n10991), .B2(n14659), .ZN(
        n10718) );
  AOI21_X1 U13275 ( .B1(n14662), .B2(n12205), .A(n10718), .ZN(n10719) );
  OAI21_X1 U13276 ( .B1(n14753), .B2(n14117), .A(n10719), .ZN(n10720) );
  AOI21_X1 U13277 ( .B1(n14756), .B2(n14113), .A(n10720), .ZN(n10721) );
  OAI21_X1 U13278 ( .B1(n10722), .B2(n14095), .A(n10721), .ZN(P1_U3285) );
  INV_X1 U13279 ( .A(n10723), .ZN(n10726) );
  OAI222_X1 U13280 ( .A1(n14370), .A2(n10726), .B1(n14368), .B2(n10725), .C1(
        P3_U3151), .C2(n6523), .ZN(P3_U3274) );
  XNOR2_X1 U13281 ( .A(n10728), .B(n10727), .ZN(n14907) );
  XNOR2_X1 U13282 ( .A(n10730), .B(n10729), .ZN(n10733) );
  OAI22_X1 U13283 ( .A1(n10731), .A2(n13536), .B1(n10770), .B2(n13538), .ZN(
        n10732) );
  AOI21_X1 U13284 ( .B1(n10733), .B2(n13407), .A(n10732), .ZN(n10734) );
  OAI21_X1 U13285 ( .B1(n14907), .B2(n13405), .A(n10734), .ZN(n14910) );
  NAND2_X1 U13286 ( .A1(n14910), .A2(n13429), .ZN(n10743) );
  OAI22_X1 U13287 ( .A1(n14884), .A2(n10736), .B1(n10735), .B2(n14877), .ZN(
        n10740) );
  OAI211_X1 U13288 ( .C1(n14909), .C2(n10738), .A(n13316), .B(n10737), .ZN(
        n14908) );
  NOR2_X1 U13289 ( .A1(n14908), .A2(n13432), .ZN(n10739) );
  AOI211_X1 U13290 ( .C1(n13440), .C2(n10741), .A(n10740), .B(n10739), .ZN(
        n10742) );
  OAI211_X1 U13291 ( .C1(n14907), .C2(n13415), .A(n10743), .B(n10742), .ZN(
        P2_U3257) );
  INV_X1 U13292 ( .A(n10744), .ZN(n10747) );
  AOI211_X1 U13293 ( .C1(n14923), .C2(n10747), .A(n10746), .B(n10745), .ZN(
        n10752) );
  NOR2_X1 U13294 ( .A1(n14925), .A2(n7890), .ZN(n10748) );
  AOI21_X1 U13295 ( .B1(n6909), .B2(n10750), .A(n10748), .ZN(n10749) );
  OAI21_X1 U13296 ( .B1(n10752), .B2(n14924), .A(n10749), .ZN(P2_U3457) );
  AOI22_X1 U13297 ( .A1(n13465), .A2(n10750), .B1(n14930), .B2(
        P2_REG1_REG_9__SCAN_IN), .ZN(n10751) );
  OAI21_X1 U13298 ( .B1(n10752), .B2(n14930), .A(n10751), .ZN(P2_U3508) );
  OAI211_X1 U13299 ( .C1(n10755), .C2(n10754), .A(n10753), .B(n12533), .ZN(
        n10762) );
  INV_X1 U13300 ( .A(n10756), .ZN(n10812) );
  INV_X1 U13301 ( .A(n12554), .ZN(n10757) );
  OAI22_X1 U13302 ( .A1(n12537), .A2(n10758), .B1(n10757), .B2(n12484), .ZN(
        n10759) );
  AOI211_X1 U13303 ( .C1(n10812), .C2(n12524), .A(n10760), .B(n10759), .ZN(
        n10761) );
  OAI211_X1 U13304 ( .C1(n12486), .C2(n10763), .A(n10762), .B(n10761), .ZN(
        P3_U3161) );
  OAI21_X1 U13305 ( .B1(n10766), .B2(n10765), .A(n10764), .ZN(n14917) );
  INV_X1 U13306 ( .A(n14917), .ZN(n10782) );
  XNOR2_X1 U13307 ( .A(n10767), .B(n10768), .ZN(n10773) );
  INV_X1 U13308 ( .A(n13405), .ZN(n14906) );
  OAI22_X1 U13309 ( .A1(n10770), .A2(n13536), .B1(n10769), .B2(n13538), .ZN(
        n10771) );
  AOI21_X1 U13310 ( .B1(n14917), .B2(n14906), .A(n10771), .ZN(n10772) );
  OAI21_X1 U13311 ( .B1(n13534), .B2(n10773), .A(n10772), .ZN(n14915) );
  NAND2_X1 U13312 ( .A1(n14915), .A2(n13429), .ZN(n10781) );
  OAI22_X1 U13313 ( .A1(n14884), .A2(n10775), .B1(n10774), .B2(n14877), .ZN(
        n10778) );
  OAI211_X1 U13314 ( .C1(n14914), .C2(n10776), .A(n13316), .B(n10857), .ZN(
        n14913) );
  NOR2_X1 U13315 ( .A1(n14913), .A2(n13432), .ZN(n10777) );
  AOI211_X1 U13316 ( .C1(n13440), .C2(n10779), .A(n10778), .B(n10777), .ZN(
        n10780) );
  OAI211_X1 U13317 ( .C1(n10782), .C2(n13415), .A(n10781), .B(n10780), .ZN(
        P2_U3255) );
  NOR2_X1 U13318 ( .A1(n11194), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n10784) );
  NOR2_X1 U13319 ( .A1(n10784), .A2(n10783), .ZN(n10788) );
  INV_X1 U13320 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n10785) );
  MUX2_X1 U13321 ( .A(n10785), .B(P1_REG2_REG_13__SCAN_IN), .S(n13789), .Z(
        n10786) );
  INV_X1 U13322 ( .A(n10786), .ZN(n10787) );
  NAND2_X1 U13323 ( .A1(n10787), .A2(n10788), .ZN(n13781) );
  OAI211_X1 U13324 ( .C1(n10788), .C2(n10787), .A(n13866), .B(n13781), .ZN(
        n10798) );
  NAND2_X1 U13325 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3086), .ZN(n13703)
         );
  INV_X1 U13326 ( .A(n13703), .ZN(n10789) );
  AOI21_X1 U13327 ( .B1(n14604), .B2(P1_ADDR_REG_13__SCAN_IN), .A(n10789), 
        .ZN(n10790) );
  INV_X1 U13328 ( .A(n10790), .ZN(n10796) );
  INV_X1 U13329 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n10792) );
  MUX2_X1 U13330 ( .A(n10792), .B(P1_REG1_REG_13__SCAN_IN), .S(n13789), .Z(
        n10793) );
  NOR2_X1 U13331 ( .A1(n10794), .A2(n10793), .ZN(n13788) );
  AOI211_X1 U13332 ( .C1(n10794), .C2(n10793), .A(n13788), .B(n13847), .ZN(
        n10795) );
  AOI211_X1 U13333 ( .C1(n14616), .C2(n13789), .A(n10796), .B(n10795), .ZN(
        n10797) );
  NAND2_X1 U13334 ( .A1(n10798), .A2(n10797), .ZN(P1_U3256) );
  INV_X1 U13335 ( .A(n10805), .ZN(n10800) );
  INV_X1 U13336 ( .A(n10799), .ZN(n10931) );
  AOI21_X1 U13337 ( .B1(n10801), .B2(n10800), .A(n10931), .ZN(n10809) );
  NAND2_X1 U13338 ( .A1(n13117), .A2(n13150), .ZN(n10802) );
  NAND2_X1 U13339 ( .A1(P2_REG3_REG_11__SCAN_IN), .A2(P2_U3088), .ZN(n14840)
         );
  OAI211_X1 U13340 ( .C1(n14467), .C2(n10855), .A(n10802), .B(n14840), .ZN(
        n10803) );
  AOI21_X1 U13341 ( .B1(n10860), .B2(n14479), .A(n10803), .ZN(n10808) );
  NOR3_X1 U13342 ( .A1(n10805), .A2(n10804), .A3(n13124), .ZN(n10806) );
  OAI21_X1 U13343 ( .B1(n10806), .B2(n13116), .A(n13152), .ZN(n10807) );
  OAI211_X1 U13344 ( .C1(n10809), .C2(n14474), .A(n10808), .B(n10807), .ZN(
        P2_U3208) );
  NAND2_X1 U13345 ( .A1(n10810), .A2(n11928), .ZN(n10811) );
  OR2_X1 U13346 ( .A1(n12554), .A2(n15100), .ZN(n10936) );
  NAND2_X1 U13347 ( .A1(n12554), .A2(n15100), .ZN(n12018) );
  NAND2_X1 U13348 ( .A1(n10936), .A2(n12018), .ZN(n12016) );
  XNOR2_X1 U13349 ( .A(n10937), .B(n12016), .ZN(n15102) );
  OR2_X1 U13350 ( .A1(n12555), .A2(n10812), .ZN(n10813) );
  INV_X1 U13351 ( .A(n12016), .ZN(n11929) );
  OAI211_X1 U13352 ( .C1(n6695), .C2(n12016), .A(n15056), .B(n10941), .ZN(
        n10816) );
  AOI22_X1 U13353 ( .A1(n15038), .A2(n12555), .B1(n14427), .B2(n15052), .ZN(
        n10815) );
  OAI211_X1 U13354 ( .C1(n15039), .C2(n15102), .A(n10816), .B(n10815), .ZN(
        n15104) );
  NAND2_X1 U13355 ( .A1(n15104), .A2(n15049), .ZN(n10820) );
  INV_X1 U13356 ( .A(n10922), .ZN(n10817) );
  OAI22_X1 U13357 ( .A1(n15049), .A2(n10642), .B1(n10817), .B2(n12868), .ZN(
        n10818) );
  AOI21_X1 U13358 ( .B1(n10939), .B2(n14423), .A(n10818), .ZN(n10819) );
  OAI211_X1 U13359 ( .C1(n15102), .C2(n10821), .A(n10820), .B(n10819), .ZN(
        P3_U3224) );
  OAI22_X1 U13360 ( .A1(n13429), .A2(n9528), .B1(n10822), .B2(n14877), .ZN(
        n10823) );
  AOI21_X1 U13361 ( .B1(n13440), .B2(n10824), .A(n10823), .ZN(n10825) );
  OAI21_X1 U13362 ( .B1(n13432), .B2(n10826), .A(n10825), .ZN(n10827) );
  AOI21_X1 U13363 ( .B1(n13442), .B2(n10828), .A(n10827), .ZN(n10829) );
  OAI21_X1 U13364 ( .B1(n13419), .B2(n10830), .A(n10829), .ZN(P2_U3264) );
  OAI22_X1 U13365 ( .A1(n13429), .A2(n9530), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        n14877), .ZN(n10833) );
  NOR2_X1 U13366 ( .A1(n13414), .A2(n10831), .ZN(n10832) );
  AOI211_X1 U13367 ( .C1(n10834), .C2(n13444), .A(n10833), .B(n10832), .ZN(
        n10837) );
  NAND2_X1 U13368 ( .A1(n13442), .A2(n10835), .ZN(n10836) );
  OAI211_X1 U13369 ( .C1(n13419), .C2(n10838), .A(n10837), .B(n10836), .ZN(
        P2_U3262) );
  OAI22_X1 U13370 ( .A1(n13429), .A2(n15291), .B1(n13161), .B2(n14877), .ZN(
        n10841) );
  NOR2_X1 U13371 ( .A1(n13414), .A2(n10839), .ZN(n10840) );
  AOI211_X1 U13372 ( .C1(n10842), .C2(n13444), .A(n10841), .B(n10840), .ZN(
        n10845) );
  NAND2_X1 U13373 ( .A1(n13442), .A2(n10843), .ZN(n10844) );
  OAI211_X1 U13374 ( .C1(n13419), .C2(n10846), .A(n10845), .B(n10844), .ZN(
        P2_U3263) );
  XNOR2_X1 U13375 ( .A(n10847), .B(n10851), .ZN(n14922) );
  INV_X1 U13376 ( .A(n14922), .ZN(n10863) );
  INV_X1 U13377 ( .A(n10848), .ZN(n10849) );
  AOI21_X1 U13378 ( .B1(n10851), .B2(n10850), .A(n10849), .ZN(n10854) );
  AOI22_X1 U13379 ( .A1(n13401), .A2(n13152), .B1(n13150), .B2(n13402), .ZN(
        n10853) );
  NAND2_X1 U13380 ( .A1(n14922), .A2(n14906), .ZN(n10852) );
  OAI211_X1 U13381 ( .C1(n10854), .C2(n13534), .A(n10853), .B(n10852), .ZN(
        n14920) );
  NAND2_X1 U13382 ( .A1(n14920), .A2(n13429), .ZN(n10862) );
  INV_X1 U13383 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n10856) );
  OAI22_X1 U13384 ( .A1(n13429), .A2(n10856), .B1(n10855), .B2(n14877), .ZN(
        n10859) );
  OAI211_X1 U13385 ( .C1(n7402), .C2(n7403), .A(n13316), .B(n10906), .ZN(
        n14918) );
  NOR2_X1 U13386 ( .A1(n14918), .A2(n13432), .ZN(n10858) );
  AOI211_X1 U13387 ( .C1(n13440), .C2(n10860), .A(n10859), .B(n10858), .ZN(
        n10861) );
  OAI211_X1 U13388 ( .C1(n10863), .C2(n13415), .A(n10862), .B(n10861), .ZN(
        P2_U3254) );
  NOR2_X1 U13389 ( .A1(n14368), .A2(SI_22_), .ZN(n10864) );
  AOI21_X1 U13390 ( .B1(n11288), .B2(P3_STATE_REG_SCAN_IN), .A(n10864), .ZN(
        n10865) );
  OAI21_X1 U13391 ( .B1(n10866), .B2(n14370), .A(n10865), .ZN(n10867) );
  INV_X1 U13392 ( .A(n10867), .ZN(P3_U3273) );
  NAND2_X1 U13393 ( .A1(n10868), .A2(n12346), .ZN(n10870) );
  OR2_X1 U13394 ( .A1(n12205), .A2(n13772), .ZN(n10869) );
  NAND2_X1 U13395 ( .A1(n10870), .A2(n10869), .ZN(n11015) );
  NAND2_X1 U13396 ( .A1(n10871), .A2(n10677), .ZN(n10874) );
  AOI22_X1 U13397 ( .A1(n11535), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n11533), 
        .B2(n10872), .ZN(n10873) );
  NAND2_X1 U13398 ( .A1(n10874), .A2(n10873), .ZN(n12214) );
  INV_X1 U13399 ( .A(n13771), .ZN(n10995) );
  XNOR2_X1 U13400 ( .A(n11015), .B(n7101), .ZN(n10889) );
  OAI21_X1 U13401 ( .B1(n6694), .B2(n7101), .A(n10997), .ZN(n10887) );
  NAND2_X1 U13402 ( .A1(n12321), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n10884) );
  OR2_X1 U13403 ( .A1(n6526), .A2(n9971), .ZN(n10883) );
  INV_X1 U13404 ( .A(n11005), .ZN(n10879) );
  NAND2_X1 U13405 ( .A1(n10877), .A2(n15304), .ZN(n10878) );
  NAND2_X1 U13406 ( .A1(n10879), .A2(n10878), .ZN(n11265) );
  OR2_X1 U13407 ( .A1(n11600), .A2(n11265), .ZN(n10882) );
  OR2_X1 U13408 ( .A1(n6539), .A2(n10880), .ZN(n10881) );
  NAND4_X1 U13409 ( .A1(n10884), .A2(n10883), .A3(n10882), .A4(n10881), .ZN(
        n13770) );
  NAND2_X1 U13410 ( .A1(n13770), .A2(n13732), .ZN(n10886) );
  NAND2_X1 U13411 ( .A1(n13772), .A2(n13897), .ZN(n10885) );
  NAND2_X1 U13412 ( .A1(n10886), .A2(n10885), .ZN(n11151) );
  AOI21_X1 U13413 ( .B1(n10887), .B2(n14694), .A(n11151), .ZN(n10888) );
  OAI21_X1 U13414 ( .B1(n14691), .B2(n10889), .A(n10888), .ZN(n14760) );
  INV_X1 U13415 ( .A(n14760), .ZN(n10896) );
  INV_X1 U13416 ( .A(n10889), .ZN(n14762) );
  INV_X1 U13417 ( .A(n12214), .ZN(n14759) );
  NAND2_X1 U13418 ( .A1(n10890), .A2(n14759), .ZN(n11061) );
  OAI211_X1 U13419 ( .C1(n10890), .C2(n14759), .A(n14109), .B(n11061), .ZN(
        n14758) );
  INV_X1 U13420 ( .A(n11154), .ZN(n10891) );
  AOI22_X1 U13421 ( .A1(n14674), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n10891), 
        .B2(n14673), .ZN(n10893) );
  NAND2_X1 U13422 ( .A1(n14662), .A2(n12214), .ZN(n10892) );
  OAI211_X1 U13423 ( .C1(n14758), .C2(n14117), .A(n10893), .B(n10892), .ZN(
        n10894) );
  AOI21_X1 U13424 ( .B1(n14762), .B2(n14670), .A(n10894), .ZN(n10895) );
  OAI21_X1 U13425 ( .B1(n10896), .B2(n14674), .A(n10895), .ZN(P1_U3284) );
  XNOR2_X1 U13426 ( .A(n10897), .B(n10898), .ZN(n14520) );
  NAND2_X1 U13427 ( .A1(n14520), .A2(n14906), .ZN(n10905) );
  NAND2_X1 U13428 ( .A1(n10899), .A2(n10898), .ZN(n10900) );
  NAND3_X1 U13429 ( .A1(n10901), .A2(n13407), .A3(n10900), .ZN(n10903) );
  AOI22_X1 U13430 ( .A1(n13401), .A2(n13151), .B1(n13149), .B2(n13402), .ZN(
        n10902) );
  AND2_X1 U13431 ( .A1(n10903), .A2(n10902), .ZN(n10904) );
  INV_X1 U13432 ( .A(n13415), .ZN(n10912) );
  NAND2_X1 U13433 ( .A1(n10906), .A2(n14516), .ZN(n10907) );
  NAND2_X1 U13434 ( .A1(n10907), .A2(n13316), .ZN(n10908) );
  OR2_X1 U13435 ( .A1(n10908), .A2(n6696), .ZN(n14517) );
  OAI22_X1 U13436 ( .A1(n13429), .A2(n11029), .B1(n10927), .B2(n14877), .ZN(
        n10909) );
  AOI21_X1 U13437 ( .B1(n14516), .B2(n13440), .A(n10909), .ZN(n10910) );
  OAI21_X1 U13438 ( .B1(n14517), .B2(n13432), .A(n10910), .ZN(n10911) );
  AOI21_X1 U13439 ( .B1(n14520), .B2(n10912), .A(n10911), .ZN(n10913) );
  OAI21_X1 U13440 ( .B1(n14522), .B2(n13419), .A(n10913), .ZN(P2_U3253) );
  INV_X1 U13441 ( .A(n10914), .ZN(n10915) );
  AOI21_X1 U13442 ( .B1(n10917), .B2(n10916), .A(n10915), .ZN(n10925) );
  OAI22_X1 U13443 ( .A1(n12537), .A2(n10919), .B1(n10918), .B2(n12484), .ZN(
        n10920) );
  AOI211_X1 U13444 ( .C1(n10939), .C2(n12524), .A(n10921), .B(n10920), .ZN(
        n10924) );
  NAND2_X1 U13445 ( .A1(n12540), .A2(n10922), .ZN(n10923) );
  OAI211_X1 U13446 ( .C1(n10925), .C2(n12507), .A(n10924), .B(n10923), .ZN(
        P3_U3171) );
  AOI22_X1 U13447 ( .A1(n13116), .A2(n13151), .B1(n13117), .B2(n13149), .ZN(
        n10926) );
  NAND2_X1 U13448 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3088), .ZN(n14857)
         );
  OAI211_X1 U13449 ( .C1(n10927), .C2(n14467), .A(n10926), .B(n14857), .ZN(
        n10933) );
  AOI22_X1 U13450 ( .A1(n10928), .A2(n14462), .B1(n13105), .B2(n13151), .ZN(
        n10930) );
  NOR3_X1 U13451 ( .A1(n10931), .A2(n10930), .A3(n10929), .ZN(n10932) );
  AOI211_X1 U13452 ( .C1(n14516), .C2(n14479), .A(n10933), .B(n10932), .ZN(
        n10934) );
  OAI21_X1 U13453 ( .B1(n10935), .B2(n14474), .A(n10934), .ZN(P2_U3196) );
  INV_X1 U13454 ( .A(n10936), .ZN(n12019) );
  NOR2_X1 U13455 ( .A1(n14427), .A2(n10946), .ZN(n12024) );
  INV_X1 U13456 ( .A(n12024), .ZN(n10938) );
  AND2_X1 U13457 ( .A1(n14427), .A2(n10946), .ZN(n12025) );
  INV_X1 U13458 ( .A(n12025), .ZN(n11174) );
  NAND2_X1 U13459 ( .A1(n10938), .A2(n11174), .ZN(n12028) );
  XNOR2_X1 U13460 ( .A(n11173), .B(n11172), .ZN(n10945) );
  NAND2_X1 U13461 ( .A1(n12554), .A2(n10939), .ZN(n10940) );
  NAND2_X1 U13462 ( .A1(n10941), .A2(n10940), .ZN(n11178) );
  XNOR2_X1 U13463 ( .A(n11178), .B(n11172), .ZN(n10942) );
  NAND2_X1 U13464 ( .A1(n10942), .A2(n15056), .ZN(n10944) );
  AOI22_X1 U13465 ( .A1(n15038), .A2(n12554), .B1(n12553), .B2(n15052), .ZN(
        n10943) );
  OAI211_X1 U13466 ( .C1(n15039), .C2(n10945), .A(n10944), .B(n10943), .ZN(
        n15105) );
  INV_X1 U13467 ( .A(n15105), .ZN(n10951) );
  INV_X1 U13468 ( .A(n10945), .ZN(n15107) );
  INV_X1 U13469 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n10948) );
  INV_X1 U13470 ( .A(n11177), .ZN(n15062) );
  NOR2_X1 U13471 ( .A1(n10946), .A2(n15099), .ZN(n15106) );
  AOI22_X1 U13472 ( .A1(n15062), .A2(n15106), .B1(n15058), .B2(n12424), .ZN(
        n10947) );
  OAI21_X1 U13473 ( .B1(n10948), .B2(n15049), .A(n10947), .ZN(n10949) );
  AOI21_X1 U13474 ( .B1(n15107), .B2(n12744), .A(n10949), .ZN(n10950) );
  OAI21_X1 U13475 ( .B1(n10951), .B2(n15066), .A(n10950), .ZN(P3_U3223) );
  NAND2_X1 U13476 ( .A1(n13772), .A2(n13732), .ZN(n10953) );
  NAND2_X1 U13477 ( .A1(n13774), .A2(n13897), .ZN(n10952) );
  NAND2_X1 U13478 ( .A1(n10953), .A2(n10952), .ZN(n14631) );
  NAND2_X1 U13479 ( .A1(n14537), .A2(n14631), .ZN(n10954) );
  OAI211_X1 U13480 ( .C1(n14542), .C2(n14633), .A(n10955), .B(n10954), .ZN(
        n10965) );
  NAND2_X1 U13481 ( .A1(n10959), .A2(n10958), .ZN(n10967) );
  NAND2_X1 U13482 ( .A1(n14743), .A2(n11778), .ZN(n10961) );
  NAND2_X1 U13483 ( .A1(n13773), .A2(n11777), .ZN(n10960) );
  NAND2_X1 U13484 ( .A1(n10961), .A2(n10960), .ZN(n10962) );
  XNOR2_X1 U13485 ( .A(n10962), .B(n11745), .ZN(n10972) );
  AOI22_X1 U13486 ( .A1(n14743), .A2(n11777), .B1(n6720), .B2(n13773), .ZN(
        n10971) );
  XNOR2_X1 U13487 ( .A(n10972), .B(n10971), .ZN(n10968) );
  XNOR2_X1 U13488 ( .A(n10967), .B(n10968), .ZN(n10963) );
  NOR2_X1 U13489 ( .A1(n10963), .A2(n13727), .ZN(n10964) );
  AOI211_X1 U13490 ( .C1(n14533), .C2(n14743), .A(n10965), .B(n10964), .ZN(
        n10966) );
  INV_X1 U13491 ( .A(n10966), .ZN(P1_U3213) );
  INV_X1 U13492 ( .A(n10967), .ZN(n10970) );
  INV_X1 U13493 ( .A(n10968), .ZN(n10969) );
  OR2_X1 U13494 ( .A1(n10972), .A2(n10971), .ZN(n10973) );
  NAND2_X1 U13495 ( .A1(n12205), .A2(n11778), .ZN(n10976) );
  NAND2_X1 U13496 ( .A1(n13772), .A2(n11777), .ZN(n10975) );
  NAND2_X1 U13497 ( .A1(n10976), .A2(n10975), .ZN(n10977) );
  XNOR2_X1 U13498 ( .A(n10977), .B(n11745), .ZN(n10979) );
  AND2_X1 U13499 ( .A1(n13772), .A2(n6720), .ZN(n10978) );
  AOI21_X1 U13500 ( .B1(n12205), .B2(n11777), .A(n10978), .ZN(n10980) );
  NAND2_X1 U13501 ( .A1(n10979), .A2(n10980), .ZN(n11145) );
  INV_X1 U13502 ( .A(n10979), .ZN(n10982) );
  INV_X1 U13503 ( .A(n10980), .ZN(n10981) );
  NAND2_X1 U13504 ( .A1(n10982), .A2(n10981), .ZN(n10983) );
  NAND2_X1 U13505 ( .A1(n11145), .A2(n10983), .ZN(n10986) );
  INV_X1 U13506 ( .A(n10986), .ZN(n10984) );
  INV_X1 U13507 ( .A(n11146), .ZN(n10985) );
  AOI21_X1 U13508 ( .B1(n10987), .B2(n10986), .A(n10985), .ZN(n10994) );
  AND2_X1 U13509 ( .A1(n12205), .A2(n14742), .ZN(n14751) );
  AOI21_X1 U13510 ( .B1(n14537), .B2(n10989), .A(n10988), .ZN(n10990) );
  OAI21_X1 U13511 ( .B1(n10991), .B2(n14542), .A(n10990), .ZN(n10992) );
  AOI21_X1 U13512 ( .B1(n14751), .B2(n13601), .A(n10992), .ZN(n10993) );
  OAI21_X1 U13513 ( .B1(n10994), .B2(n13727), .A(n10993), .ZN(P1_U3221) );
  INV_X1 U13514 ( .A(n11548), .ZN(n11071) );
  INV_X1 U13515 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n11549) );
  OAI222_X1 U13516 ( .A1(P1_U3086), .A2(n12143), .B1(n11860), .B2(n11071), 
        .C1(n11549), .C2(n14247), .ZN(P1_U3335) );
  NAND2_X1 U13517 ( .A1(n12214), .A2(n10995), .ZN(n10996) );
  NAND2_X1 U13518 ( .A1(n10998), .A2(n10677), .ZN(n11001) );
  AOI22_X1 U13519 ( .A1(n11535), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n11533), 
        .B2(n10999), .ZN(n11000) );
  NAND2_X2 U13520 ( .A1(n11001), .A2(n11000), .ZN(n12217) );
  INV_X1 U13521 ( .A(n13770), .ZN(n11059) );
  OR2_X1 U13522 ( .A1(n12217), .A2(n11059), .ZN(n11046) );
  NAND2_X1 U13523 ( .A1(n12217), .A2(n11059), .ZN(n11002) );
  AOI21_X1 U13524 ( .B1(n11003), .B2(n11066), .A(n14737), .ZN(n11004) );
  AOI22_X1 U13525 ( .A1(n11004), .A2(n11047), .B1(n13897), .B2(n13771), .ZN(
        n14766) );
  OAI22_X1 U13526 ( .A1(n14113), .A2(n9971), .B1(n11265), .B2(n14659), .ZN(
        n11014) );
  INV_X1 U13527 ( .A(n12217), .ZN(n14768) );
  XNOR2_X1 U13528 ( .A(n11061), .B(n14768), .ZN(n11012) );
  NAND2_X1 U13529 ( .A1(n12321), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n11011) );
  OR2_X1 U13530 ( .A1(n11005), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n11006) );
  NAND2_X1 U13531 ( .A1(n11053), .A2(n11006), .ZN(n11383) );
  OR2_X1 U13532 ( .A1(n11600), .A2(n11383), .ZN(n11010) );
  OR2_X1 U13533 ( .A1(n6526), .A2(n11063), .ZN(n11009) );
  OR2_X1 U13534 ( .A1(n6540), .A2(n11007), .ZN(n11008) );
  NAND4_X1 U13535 ( .A1(n11011), .A2(n11010), .A3(n11009), .A4(n11008), .ZN(
        n13769) );
  AOI22_X1 U13536 ( .A1(n11012), .A2(n14109), .B1(n13732), .B2(n13769), .ZN(
        n14765) );
  NOR2_X1 U13537 ( .A1(n14765), .A2(n14117), .ZN(n11013) );
  AOI211_X1 U13538 ( .C1(n14662), .C2(n12217), .A(n11014), .B(n11013), .ZN(
        n11018) );
  OR2_X1 U13539 ( .A1(n12214), .A2(n13771), .ZN(n11016) );
  XNOR2_X1 U13540 ( .A(n11067), .B(n11066), .ZN(n14770) );
  NAND2_X1 U13541 ( .A1(n14770), .A2(n14676), .ZN(n11017) );
  OAI211_X1 U13542 ( .C1(n14766), .C2(n14674), .A(n11018), .B(n11017), .ZN(
        P1_U3283) );
  NOR2_X1 U13543 ( .A1(n11165), .A2(n11019), .ZN(n11020) );
  AOI21_X1 U13544 ( .B1(n11019), .B2(n11165), .A(n11020), .ZN(n11024) );
  MUX2_X1 U13545 ( .A(n11022), .B(P2_REG1_REG_11__SCAN_IN), .S(n11027), .Z(
        n14828) );
  OAI21_X1 U13546 ( .B1(n14855), .B2(P2_REG1_REG_12__SCAN_IN), .A(n14850), 
        .ZN(n11023) );
  AOI211_X1 U13547 ( .C1(n11024), .C2(n11023), .A(n14863), .B(n11164), .ZN(
        n11039) );
  MUX2_X1 U13548 ( .A(n13438), .B(P2_REG2_REG_13__SCAN_IN), .S(n11165), .Z(
        n11033) );
  MUX2_X1 U13549 ( .A(P2_REG2_REG_11__SCAN_IN), .B(n10856), .S(n11027), .Z(
        n14831) );
  NOR2_X1 U13550 ( .A1(n11027), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n14844) );
  NAND2_X1 U13551 ( .A1(n14855), .A2(n11029), .ZN(n11028) );
  OAI21_X1 U13552 ( .B1(n14855), .B2(n11029), .A(n11028), .ZN(n14843) );
  OAI21_X1 U13553 ( .B1(n14855), .B2(P2_REG2_REG_12__SCAN_IN), .A(n14847), 
        .ZN(n11032) );
  NOR2_X1 U13554 ( .A1(n11031), .A2(n13438), .ZN(n11030) );
  AOI211_X1 U13555 ( .C1(n11033), .C2(n11032), .A(n14836), .B(n11159), .ZN(
        n11038) );
  INV_X1 U13556 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n11036) );
  NAND2_X1 U13557 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(P2_U3088), .ZN(n11110)
         );
  INV_X1 U13558 ( .A(n11110), .ZN(n11034) );
  AOI21_X1 U13559 ( .B1(n14868), .B2(n11165), .A(n11034), .ZN(n11035) );
  OAI21_X1 U13560 ( .B1(n14874), .B2(n11036), .A(n11035), .ZN(n11037) );
  OR3_X1 U13561 ( .A1(n11039), .A2(n11038), .A3(n11037), .ZN(P2_U3227) );
  NAND2_X1 U13562 ( .A1(n11040), .A2(n14381), .ZN(n11041) );
  OAI211_X1 U13563 ( .C1(n11042), .C2(n14368), .A(n11041), .B(n12116), .ZN(
        P3_U3272) );
  INV_X1 U13564 ( .A(n11486), .ZN(n11043) );
  OAI222_X1 U13565 ( .A1(P1_U3086), .A2(n6773), .B1(n11860), .B2(n11043), .C1(
        n11487), .C2(n14247), .ZN(P1_U3334) );
  OAI222_X1 U13566 ( .A1(n13594), .A2(n11045), .B1(P2_U3088), .B2(n11044), 
        .C1(n13596), .C2(n11043), .ZN(P2_U3306) );
  NAND2_X1 U13567 ( .A1(n11048), .A2(n10677), .ZN(n11051) );
  AOI22_X1 U13568 ( .A1(n11535), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n11533), 
        .B2(n11049), .ZN(n11050) );
  INV_X1 U13569 ( .A(n13769), .ZN(n11270) );
  XNOR2_X1 U13570 ( .A(n11191), .B(n12355), .ZN(n11060) );
  NAND2_X1 U13571 ( .A1(n12321), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n11058) );
  OR2_X1 U13572 ( .A1(n6526), .A2(n10324), .ZN(n11057) );
  NAND2_X1 U13573 ( .A1(n11053), .A2(n11052), .ZN(n11054) );
  NAND2_X1 U13574 ( .A1(n11203), .A2(n11054), .ZN(n13645) );
  OR2_X1 U13575 ( .A1(n11600), .A2(n13645), .ZN(n11056) );
  OR2_X1 U13576 ( .A1(n6539), .A2(n15368), .ZN(n11055) );
  NAND4_X1 U13577 ( .A1(n11058), .A2(n11057), .A3(n11056), .A4(n11055), .ZN(
        n13768) );
  INV_X1 U13578 ( .A(n13768), .ZN(n11217) );
  OAI22_X1 U13579 ( .A1(n11059), .A2(n13674), .B1(n11217), .B2(n14678), .ZN(
        n11380) );
  AOI21_X1 U13580 ( .B1(n11060), .B2(n14694), .A(n11380), .ZN(n14565) );
  OR2_X2 U13581 ( .A1(n11061), .A2(n12217), .ZN(n11062) );
  AOI211_X1 U13582 ( .C1(n12225), .C2(n11062), .A(n14663), .B(n11247), .ZN(
        n14562) );
  INV_X1 U13583 ( .A(n12225), .ZN(n14564) );
  NOR2_X1 U13584 ( .A1(n14564), .A2(n14089), .ZN(n11065) );
  OAI22_X1 U13585 ( .A1(n14113), .A2(n11063), .B1(n11383), .B2(n14659), .ZN(
        n11064) );
  AOI211_X1 U13586 ( .C1(n14562), .C2(n14669), .A(n11065), .B(n11064), .ZN(
        n11070) );
  OR2_X1 U13587 ( .A1(n12217), .A2(n13770), .ZN(n11068) );
  XNOR2_X1 U13588 ( .A(n11219), .B(n12355), .ZN(n14568) );
  NAND2_X1 U13589 ( .A1(n14568), .A2(n14676), .ZN(n11069) );
  OAI211_X1 U13590 ( .C1(n14565), .C2(n14674), .A(n11070), .B(n11069), .ZN(
        P1_U3282) );
  OAI222_X1 U13591 ( .A1(n13588), .A2(n11072), .B1(P2_U3088), .B2(n6531), .C1(
        n13596), .C2(n11071), .ZN(P2_U3307) );
  XNOR2_X1 U13592 ( .A(n11073), .B(n11075), .ZN(n13443) );
  OR2_X1 U13593 ( .A1(n6696), .A2(n11079), .ZN(n11074) );
  AND3_X1 U13594 ( .A1(n11230), .A2(n13316), .A3(n11074), .ZN(n13445) );
  XNOR2_X1 U13595 ( .A(n11076), .B(n11075), .ZN(n11077) );
  OAI222_X1 U13596 ( .A1(n13538), .A2(n13535), .B1(n13536), .B2(n11078), .C1(
        n11077), .C2(n13534), .ZN(n13436) );
  AOI211_X1 U13597 ( .C1(n14515), .C2(n13443), .A(n13445), .B(n13436), .ZN(
        n11083) );
  OAI22_X1 U13598 ( .A1(n11079), .A2(n13573), .B1(n14925), .B2(n7956), .ZN(
        n11080) );
  INV_X1 U13599 ( .A(n11080), .ZN(n11081) );
  OAI21_X1 U13600 ( .B1(n11083), .B2(n14924), .A(n11081), .ZN(P2_U3469) );
  AOI22_X1 U13601 ( .A1(n13441), .A2(n13465), .B1(n14930), .B2(
        P2_REG1_REG_13__SCAN_IN), .ZN(n11082) );
  OAI21_X1 U13602 ( .B1(n11083), .B2(n14930), .A(n11082), .ZN(P2_U3512) );
  INV_X1 U13603 ( .A(n11084), .ZN(n11086) );
  AOI22_X1 U13604 ( .A1(n15014), .A2(P3_REG2_REG_10__SCAN_IN), .B1(n10948), 
        .B2(n14374), .ZN(n15021) );
  NAND2_X1 U13605 ( .A1(n11087), .A2(n11131), .ZN(n11124) );
  INV_X1 U13606 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n11088) );
  AOI21_X1 U13607 ( .B1(n11089), .B2(n11088), .A(n11125), .ZN(n11109) );
  MUX2_X1 U13608 ( .A(P3_REG2_REG_10__SCAN_IN), .B(P3_REG1_REG_10__SCAN_IN), 
        .S(n12670), .Z(n11094) );
  XNOR2_X1 U13609 ( .A(n11094), .B(n15014), .ZN(n15011) );
  INV_X1 U13610 ( .A(n11094), .ZN(n11095) );
  AOI22_X1 U13611 ( .A1(n15012), .A2(n15011), .B1(n15014), .B2(n11095), .ZN(
        n11134) );
  MUX2_X1 U13612 ( .A(P3_REG2_REG_11__SCAN_IN), .B(P3_REG1_REG_11__SCAN_IN), 
        .S(n12670), .Z(n11132) );
  XOR2_X1 U13613 ( .A(n11096), .B(n11132), .Z(n11133) );
  XNOR2_X1 U13614 ( .A(n11134), .B(n11133), .ZN(n11107) );
  INV_X1 U13615 ( .A(P3_REG3_REG_11__SCAN_IN), .ZN(n11097) );
  NOR2_X1 U13616 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11097), .ZN(n11301) );
  AOI21_X1 U13617 ( .B1(n15001), .B2(P3_ADDR_REG_11__SCAN_IN), .A(n11301), 
        .ZN(n11098) );
  OAI21_X1 U13618 ( .B1(n12701), .B2(n11131), .A(n11098), .ZN(n11106) );
  INV_X1 U13619 ( .A(n11099), .ZN(n11101) );
  INV_X1 U13620 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n15269) );
  AOI22_X1 U13621 ( .A1(n15014), .A2(P3_REG1_REG_10__SCAN_IN), .B1(n15269), 
        .B2(n14374), .ZN(n15009) );
  AND2_X1 U13622 ( .A1(n14374), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n11102) );
  INV_X1 U13623 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n15377) );
  AOI21_X1 U13624 ( .B1(n11103), .B2(n15377), .A(n11120), .ZN(n11104) );
  NOR2_X1 U13625 ( .A1(n11104), .A2(n15018), .ZN(n11105) );
  AOI211_X1 U13626 ( .C1(n15015), .C2(n11107), .A(n11106), .B(n11105), .ZN(
        n11108) );
  OAI21_X1 U13627 ( .B1(n11109), .B2(n15023), .A(n11108), .ZN(P3_U3193) );
  AOI22_X1 U13628 ( .A1(n13116), .A2(n13150), .B1(n13117), .B2(n13148), .ZN(
        n11111) );
  OAI211_X1 U13629 ( .C1(n13437), .C2(n14467), .A(n11111), .B(n11110), .ZN(
        n11117) );
  INV_X1 U13630 ( .A(n11112), .ZN(n11113) );
  AOI211_X1 U13631 ( .C1(n11115), .C2(n11114), .A(n14474), .B(n11113), .ZN(
        n11116) );
  AOI211_X1 U13632 ( .C1(n13441), .C2(n14479), .A(n11117), .B(n11116), .ZN(
        n11118) );
  INV_X1 U13633 ( .A(n11118), .ZN(P2_U3206) );
  NAND2_X1 U13634 ( .A1(P3_REG1_REG_12__SCAN_IN), .A2(n12564), .ZN(n11121) );
  OAI21_X1 U13635 ( .B1(P3_REG1_REG_12__SCAN_IN), .B2(n12564), .A(n11121), 
        .ZN(n11122) );
  AOI21_X1 U13636 ( .B1(n11123), .B2(n11122), .A(n12559), .ZN(n11141) );
  INV_X1 U13637 ( .A(n12564), .ZN(n11139) );
  NAND2_X1 U13638 ( .A1(n12564), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n12570) );
  OAI21_X1 U13639 ( .B1(P3_REG2_REG_12__SCAN_IN), .B2(n12564), .A(n12570), 
        .ZN(n11127) );
  AOI21_X1 U13640 ( .B1(n11127), .B2(n6679), .A(n12568), .ZN(n11130) );
  INV_X1 U13641 ( .A(P3_REG3_REG_12__SCAN_IN), .ZN(n11128) );
  NOR2_X1 U13642 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11128), .ZN(n11391) );
  AOI21_X1 U13643 ( .B1(n15001), .B2(P3_ADDR_REG_12__SCAN_IN), .A(n11391), 
        .ZN(n11129) );
  OAI21_X1 U13644 ( .B1(n11130), .B2(n15023), .A(n11129), .ZN(n11138) );
  MUX2_X1 U13645 ( .A(P3_REG2_REG_12__SCAN_IN), .B(P3_REG1_REG_12__SCAN_IN), 
        .S(n12670), .Z(n12565) );
  XNOR2_X1 U13646 ( .A(n12564), .B(n12565), .ZN(n11136) );
  OAI22_X1 U13647 ( .A1(n11134), .A2(n11133), .B1(n11132), .B2(n11131), .ZN(
        n11135) );
  AOI211_X1 U13648 ( .C1(n11136), .C2(n11135), .A(n14948), .B(n12563), .ZN(
        n11137) );
  AOI211_X1 U13649 ( .C1(n15013), .C2(n11139), .A(n11138), .B(n11137), .ZN(
        n11140) );
  OAI21_X1 U13650 ( .B1(n11141), .B2(n15018), .A(n11140), .ZN(P3_U3194) );
  NAND2_X1 U13651 ( .A1(n12214), .A2(n11778), .ZN(n11143) );
  NAND2_X1 U13652 ( .A1(n13771), .A2(n11777), .ZN(n11142) );
  NAND2_X1 U13653 ( .A1(n11143), .A2(n11142), .ZN(n11144) );
  XNOR2_X1 U13654 ( .A(n11144), .B(n11745), .ZN(n11150) );
  NAND2_X1 U13655 ( .A1(n12214), .A2(n11777), .ZN(n11148) );
  NAND2_X1 U13656 ( .A1(n13771), .A2(n6720), .ZN(n11147) );
  NAND2_X1 U13657 ( .A1(n11148), .A2(n11147), .ZN(n11253) );
  XNOR2_X1 U13658 ( .A(n11255), .B(n11253), .ZN(n11149) );
  OAI21_X1 U13659 ( .B1(n11150), .B2(n11149), .A(n11262), .ZN(n11157) );
  NOR2_X1 U13660 ( .A1(n13753), .A2(n14759), .ZN(n11156) );
  NAND2_X1 U13661 ( .A1(n14537), .A2(n11151), .ZN(n11152) );
  OAI211_X1 U13662 ( .C1(n14542), .C2(n11154), .A(n11153), .B(n11152), .ZN(
        n11155) );
  AOI211_X1 U13663 ( .C1(n11157), .C2(n14535), .A(n11156), .B(n11155), .ZN(
        n11158) );
  INV_X1 U13664 ( .A(n11158), .ZN(P1_U3231) );
  INV_X1 U13665 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n11444) );
  XNOR2_X1 U13666 ( .A(n11445), .B(n11444), .ZN(n11171) );
  NAND2_X1 U13667 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3088), .ZN(n14464)
         );
  INV_X1 U13668 ( .A(n14464), .ZN(n11160) );
  AOI21_X1 U13669 ( .B1(n14868), .B2(n11452), .A(n11160), .ZN(n11161) );
  INV_X1 U13670 ( .A(n11161), .ZN(n11169) );
  NOR2_X1 U13671 ( .A1(n11452), .A2(n11162), .ZN(n11163) );
  AOI21_X1 U13672 ( .B1(n11452), .B2(n11162), .A(n11163), .ZN(n11167) );
  AOI211_X1 U13673 ( .C1(n11167), .C2(n11166), .A(n14863), .B(n11451), .ZN(
        n11168) );
  AOI211_X1 U13674 ( .C1(n14789), .C2(P2_ADDR_REG_14__SCAN_IN), .A(n11169), 
        .B(n11168), .ZN(n11170) );
  OAI21_X1 U13675 ( .B1(n11171), .B2(n14836), .A(n11170), .ZN(P2_U3228) );
  NAND2_X1 U13676 ( .A1(n11175), .A2(n11174), .ZN(n14431) );
  OR2_X1 U13677 ( .A1(n14434), .A2(n12553), .ZN(n12030) );
  NAND2_X1 U13678 ( .A1(n14434), .A2(n12553), .ZN(n12035) );
  NAND2_X1 U13679 ( .A1(n12030), .A2(n12035), .ZN(n14432) );
  INV_X1 U13680 ( .A(n11279), .ZN(n11398) );
  AND2_X1 U13681 ( .A1(n11398), .A2(n14428), .ZN(n12032) );
  INV_X1 U13682 ( .A(n12032), .ZN(n12036) );
  NAND2_X1 U13683 ( .A1(n11279), .A2(n11419), .ZN(n12037) );
  XNOR2_X1 U13684 ( .A(n11282), .B(n11933), .ZN(n14443) );
  NAND2_X1 U13685 ( .A1(n11279), .A2(n14441), .ZN(n14444) );
  AOI22_X1 U13686 ( .A1(n15066), .A2(P3_REG2_REG_12__SCAN_IN), .B1(n15058), 
        .B2(n11395), .ZN(n11176) );
  OAI21_X1 U13687 ( .B1(n11177), .B2(n14444), .A(n11176), .ZN(n11188) );
  NAND2_X1 U13688 ( .A1(n11178), .A2(n12028), .ZN(n11180) );
  NAND2_X1 U13689 ( .A1(n12423), .A2(n14427), .ZN(n11179) );
  INV_X1 U13690 ( .A(n12553), .ZN(n11298) );
  NOR2_X1 U13691 ( .A1(n14434), .A2(n11298), .ZN(n11182) );
  NAND2_X1 U13692 ( .A1(n11183), .A2(n11933), .ZN(n11184) );
  NAND3_X1 U13693 ( .A1(n11280), .A2(n15056), .A3(n11184), .ZN(n11186) );
  AOI22_X1 U13694 ( .A1(n15038), .A2(n12553), .B1(n12552), .B2(n15052), .ZN(
        n11185) );
  AND2_X1 U13695 ( .A1(n11186), .A2(n11185), .ZN(n14446) );
  NOR2_X1 U13696 ( .A1(n14446), .A2(n15066), .ZN(n11187) );
  AOI211_X1 U13697 ( .C1(n14443), .C2(n15063), .A(n11188), .B(n11187), .ZN(
        n11189) );
  INV_X1 U13698 ( .A(n11189), .ZN(P3_U3221) );
  INV_X1 U13699 ( .A(n12355), .ZN(n11190) );
  OR2_X1 U13700 ( .A1(n12225), .A2(n11270), .ZN(n11192) );
  NAND2_X1 U13701 ( .A1(n11193), .A2(n10677), .ZN(n11196) );
  AOI22_X1 U13702 ( .A1(n11535), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n11533), 
        .B2(n11194), .ZN(n11195) );
  XNOR2_X1 U13703 ( .A(n12235), .B(n13768), .ZN(n12350) );
  OR2_X1 U13704 ( .A1(n12235), .A2(n11217), .ZN(n11197) );
  NAND2_X1 U13705 ( .A1(n11198), .A2(n10677), .ZN(n11200) );
  AOI22_X1 U13706 ( .A1(n11535), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n11533), 
        .B2(n13789), .ZN(n11199) );
  NAND2_X1 U13707 ( .A1(n11783), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n11209) );
  INV_X1 U13708 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n11201) );
  OR2_X1 U13709 ( .A1(n11784), .A2(n11201), .ZN(n11208) );
  INV_X1 U13710 ( .A(n11210), .ZN(n11205) );
  NAND2_X1 U13711 ( .A1(n11203), .A2(n11202), .ZN(n11204) );
  NAND2_X1 U13712 ( .A1(n11205), .A2(n11204), .ZN(n13704) );
  OR2_X1 U13713 ( .A1(n11600), .A2(n13704), .ZN(n11207) );
  OR2_X1 U13714 ( .A1(n6526), .A2(n10785), .ZN(n11206) );
  NAND4_X1 U13715 ( .A1(n11209), .A2(n11208), .A3(n11207), .A4(n11206), .ZN(
        n13767) );
  XNOR2_X1 U13716 ( .A(n13706), .B(n13767), .ZN(n12353) );
  XNOR2_X1 U13717 ( .A(n11306), .B(n11312), .ZN(n11218) );
  NAND2_X1 U13718 ( .A1(n12321), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n11216) );
  INV_X1 U13719 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n13787) );
  OR2_X1 U13720 ( .A1(n6540), .A2(n13787), .ZN(n11215) );
  NOR2_X1 U13721 ( .A1(n11210), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n11211) );
  OR2_X1 U13722 ( .A1(n11212), .A2(n11211), .ZN(n14541) );
  OR2_X1 U13723 ( .A1(n11600), .A2(n14541), .ZN(n11214) );
  INV_X1 U13724 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n13783) );
  OR2_X1 U13725 ( .A1(n6526), .A2(n13783), .ZN(n11213) );
  NAND4_X1 U13726 ( .A1(n11216), .A2(n11215), .A3(n11214), .A4(n11213), .ZN(
        n13766) );
  INV_X1 U13727 ( .A(n13766), .ZN(n11609) );
  OAI22_X1 U13728 ( .A1(n11609), .A2(n14678), .B1(n11217), .B2(n13674), .ZN(
        n13701) );
  AOI21_X1 U13729 ( .B1(n11218), .B2(n14694), .A(n13701), .ZN(n14558) );
  OR2_X1 U13730 ( .A1(n12225), .A2(n13769), .ZN(n11220) );
  INV_X1 U13731 ( .A(n12350), .ZN(n11239) );
  OR2_X1 U13732 ( .A1(n12235), .A2(n13768), .ZN(n11221) );
  XNOR2_X1 U13733 ( .A(n11313), .B(n11312), .ZN(n14561) );
  INV_X1 U13734 ( .A(n13706), .ZN(n14557) );
  OAI211_X1 U13735 ( .C1(n11245), .C2(n14557), .A(n14109), .B(n6693), .ZN(
        n14556) );
  OAI22_X1 U13736 ( .A1(n14113), .A2(n10785), .B1(n13704), .B2(n14659), .ZN(
        n11222) );
  AOI21_X1 U13737 ( .B1(n13706), .B2(n14662), .A(n11222), .ZN(n11223) );
  OAI21_X1 U13738 ( .B1(n14556), .B2(n14117), .A(n11223), .ZN(n11224) );
  AOI21_X1 U13739 ( .B1(n14561), .B2(n14676), .A(n11224), .ZN(n11225) );
  OAI21_X1 U13740 ( .B1(n14558), .B2(n14674), .A(n11225), .ZN(P1_U3280) );
  XNOR2_X1 U13741 ( .A(n11226), .B(n11228), .ZN(n14514) );
  INV_X1 U13742 ( .A(n14514), .ZN(n11237) );
  AOI21_X1 U13743 ( .B1(n11228), .B2(n11227), .A(n8251), .ZN(n11229) );
  OAI222_X1 U13744 ( .A1(n13536), .A2(n14459), .B1(n13538), .B2(n14471), .C1(
        n13534), .C2(n11229), .ZN(n14512) );
  INV_X1 U13745 ( .A(n11230), .ZN(n11231) );
  INV_X1 U13746 ( .A(n11233), .ZN(n14511) );
  OAI211_X1 U13747 ( .C1(n11231), .C2(n14511), .A(n13316), .B(n13527), .ZN(
        n14510) );
  OAI22_X1 U13748 ( .A1(n13429), .A2(n11444), .B1(n14466), .B2(n14877), .ZN(
        n11232) );
  AOI21_X1 U13749 ( .B1(n11233), .B2(n13440), .A(n11232), .ZN(n11234) );
  OAI21_X1 U13750 ( .B1(n14510), .B2(n13432), .A(n11234), .ZN(n11235) );
  AOI21_X1 U13751 ( .B1(n14512), .B2(n13429), .A(n11235), .ZN(n11236) );
  OAI21_X1 U13752 ( .B1(n11237), .B2(n13393), .A(n11236), .ZN(P2_U3251) );
  XNOR2_X1 U13753 ( .A(n11238), .B(n12350), .ZN(n14391) );
  INV_X1 U13754 ( .A(n14670), .ZN(n11252) );
  XNOR2_X1 U13755 ( .A(n6763), .B(n11239), .ZN(n11243) );
  NAND2_X1 U13756 ( .A1(n13767), .A2(n13732), .ZN(n11242) );
  NAND2_X1 U13757 ( .A1(n13769), .A2(n13897), .ZN(n11241) );
  NAND2_X1 U13758 ( .A1(n11242), .A2(n11241), .ZN(n13648) );
  AOI21_X1 U13759 ( .B1(n11243), .B2(n14694), .A(n13648), .ZN(n11244) );
  OAI21_X1 U13760 ( .B1(n14691), .B2(n14391), .A(n11244), .ZN(n14394) );
  NAND2_X1 U13761 ( .A1(n14394), .A2(n14113), .ZN(n11251) );
  OAI22_X1 U13762 ( .A1(n14113), .A2(n10324), .B1(n13645), .B2(n14659), .ZN(
        n11249) );
  INV_X1 U13763 ( .A(n11245), .ZN(n11246) );
  OAI211_X1 U13764 ( .C1(n14393), .C2(n11247), .A(n11246), .B(n14109), .ZN(
        n14392) );
  NOR2_X1 U13765 ( .A1(n14392), .A2(n14117), .ZN(n11248) );
  AOI211_X1 U13766 ( .C1(n14662), .C2(n12235), .A(n11249), .B(n11248), .ZN(
        n11250) );
  OAI211_X1 U13767 ( .C1(n14391), .C2(n11252), .A(n11251), .B(n11250), .ZN(
        P1_U3281) );
  INV_X1 U13768 ( .A(n11253), .ZN(n11254) );
  AND2_X1 U13769 ( .A1(n11262), .A2(n11260), .ZN(n11264) );
  NAND2_X1 U13770 ( .A1(n12217), .A2(n11778), .ZN(n11257) );
  NAND2_X1 U13771 ( .A1(n13770), .A2(n11777), .ZN(n11256) );
  NAND2_X1 U13772 ( .A1(n11257), .A2(n11256), .ZN(n11258) );
  XNOR2_X1 U13773 ( .A(n11258), .B(n11775), .ZN(n11374) );
  AND2_X1 U13774 ( .A1(n13770), .A2(n6720), .ZN(n11259) );
  AOI21_X1 U13775 ( .B1(n12217), .B2(n11777), .A(n11259), .ZN(n11372) );
  XNOR2_X1 U13776 ( .A(n11374), .B(n11372), .ZN(n11263) );
  OAI211_X1 U13777 ( .C1(n11264), .C2(n11263), .A(n14535), .B(n11376), .ZN(
        n11274) );
  INV_X1 U13778 ( .A(n11265), .ZN(n11272) );
  AOI21_X1 U13779 ( .B1(n11267), .B2(n13771), .A(n11266), .ZN(n11268) );
  OAI21_X1 U13780 ( .B1(n11270), .B2(n11269), .A(n11268), .ZN(n11271) );
  AOI21_X1 U13781 ( .B1(n11272), .B2(n13717), .A(n11271), .ZN(n11273) );
  OAI211_X1 U13782 ( .C1(n14768), .C2(n13753), .A(n11274), .B(n11273), .ZN(
        P1_U3217) );
  INV_X1 U13783 ( .A(n11275), .ZN(n11278) );
  INV_X1 U13784 ( .A(n8626), .ZN(n11276) );
  OAI222_X1 U13785 ( .A1(n14370), .A2(n11278), .B1(n14368), .B2(n11277), .C1(
        P3_U3151), .C2(n11276), .ZN(P3_U3271) );
  OR2_X1 U13786 ( .A1(n11420), .A2(n12552), .ZN(n12043) );
  NAND2_X1 U13787 ( .A1(n11420), .A2(n12552), .ZN(n12042) );
  AND2_X1 U13788 ( .A1(n12043), .A2(n12042), .ZN(n12040) );
  XNOR2_X1 U13789 ( .A(n11356), .B(n12040), .ZN(n11281) );
  AOI222_X1 U13790 ( .A1(n15056), .A2(n11281), .B1(n12551), .B2(n15052), .C1(
        n14428), .C2(n15038), .ZN(n11295) );
  XNOR2_X1 U13791 ( .A(n11361), .B(n12040), .ZN(n11293) );
  INV_X1 U13792 ( .A(n14423), .ZN(n12766) );
  NOR2_X1 U13793 ( .A1(n11420), .A2(n12766), .ZN(n11285) );
  INV_X1 U13794 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n12571) );
  INV_X1 U13795 ( .A(n11423), .ZN(n11283) );
  OAI22_X1 U13796 ( .A1(n15049), .A2(n12571), .B1(n11283), .B2(n12868), .ZN(
        n11284) );
  AOI211_X1 U13797 ( .C1(n11293), .C2(n15063), .A(n11285), .B(n11284), .ZN(
        n11286) );
  OAI21_X1 U13798 ( .B1(n11295), .B2(n15066), .A(n11286), .ZN(P3_U3220) );
  NAND2_X1 U13799 ( .A1(n11288), .A2(n11287), .ZN(n15101) );
  AND2_X1 U13800 ( .A1(n15039), .A2(n15101), .ZN(n12889) );
  NAND2_X1 U13801 ( .A1(n15131), .A2(n15094), .ZN(n12924) );
  INV_X1 U13802 ( .A(n12924), .ZN(n12914) );
  INV_X1 U13803 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n12561) );
  OAI22_X1 U13804 ( .A1(n11420), .A2(n12907), .B1(n15131), .B2(n12561), .ZN(
        n11289) );
  AOI21_X1 U13805 ( .B1(n11293), .B2(n12914), .A(n11289), .ZN(n11290) );
  OAI21_X1 U13806 ( .B1(n11295), .B2(n15129), .A(n11290), .ZN(P3_U3472) );
  NAND2_X1 U13807 ( .A1(n15110), .A2(n15094), .ZN(n12999) );
  INV_X1 U13808 ( .A(n12999), .ZN(n12989) );
  OAI22_X1 U13809 ( .A1(n11420), .A2(n12980), .B1(n15110), .B2(n11291), .ZN(
        n11292) );
  AOI21_X1 U13810 ( .B1(n11293), .B2(n12989), .A(n11292), .ZN(n11294) );
  OAI21_X1 U13811 ( .B1(n11295), .B2(n15109), .A(n11294), .ZN(P3_U3429) );
  NAND2_X1 U13812 ( .A1(n6872), .A2(n11297), .ZN(n11299) );
  XNOR2_X1 U13813 ( .A(n11299), .B(n11298), .ZN(n11305) );
  NOR2_X1 U13814 ( .A1(n12484), .A2(n11419), .ZN(n11300) );
  AOI211_X1 U13815 ( .C1(n12525), .C2(n14427), .A(n11301), .B(n11300), .ZN(
        n11302) );
  OAI21_X1 U13816 ( .B1(n12544), .B2(n14434), .A(n11302), .ZN(n11303) );
  AOI21_X1 U13817 ( .B1(n14430), .B2(n12540), .A(n11303), .ZN(n11304) );
  OAI21_X1 U13818 ( .B1(n11305), .B2(n12507), .A(n11304), .ZN(P3_U3176) );
  INV_X1 U13819 ( .A(n13767), .ZN(n11307) );
  NAND2_X1 U13820 ( .A1(n11308), .A2(n10677), .ZN(n11310) );
  AOI22_X1 U13821 ( .A1(n11535), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n13806), 
        .B2(n11533), .ZN(n11309) );
  XNOR2_X1 U13822 ( .A(n14534), .B(n13766), .ZN(n12247) );
  XNOR2_X1 U13823 ( .A(n11608), .B(n6699), .ZN(n14555) );
  AOI21_X1 U13824 ( .B1(n6693), .B2(n14534), .A(n14663), .ZN(n11311) );
  NAND2_X1 U13825 ( .A1(n11311), .A2(n14107), .ZN(n14549) );
  OR2_X1 U13826 ( .A1(n13706), .A2(n13767), .ZN(n11314) );
  NAND2_X1 U13827 ( .A1(n11316), .A2(n12247), .ZN(n14551) );
  NAND3_X1 U13828 ( .A1(n14552), .A2(n14551), .A3(n14676), .ZN(n11322) );
  NOR2_X1 U13829 ( .A1(n14113), .A2(n13783), .ZN(n11320) );
  OR2_X1 U13830 ( .A1(n13663), .A2(n14678), .ZN(n11318) );
  NAND2_X1 U13831 ( .A1(n13767), .A2(n13897), .ZN(n11317) );
  NAND2_X1 U13832 ( .A1(n11318), .A2(n11317), .ZN(n14538) );
  INV_X1 U13833 ( .A(n14538), .ZN(n14548) );
  OAI22_X1 U13834 ( .A1(n14674), .A2(n14548), .B1(n14541), .B2(n14659), .ZN(
        n11319) );
  AOI211_X1 U13835 ( .C1(n14534), .C2(n14662), .A(n11320), .B(n11319), .ZN(
        n11321) );
  OAI211_X1 U13836 ( .C1(n14549), .C2(n14117), .A(n11322), .B(n11321), .ZN(
        n11323) );
  AOI21_X1 U13837 ( .B1(n14555), .B2(n14675), .A(n11323), .ZN(n11324) );
  INV_X1 U13838 ( .A(n11324), .ZN(P1_U3279) );
  NAND2_X1 U13839 ( .A1(n11573), .A2(n11325), .ZN(n11326) );
  OAI211_X1 U13840 ( .C1(n11574), .C2(n14247), .A(n11326), .B(n12384), .ZN(
        P1_U3332) );
  NAND2_X1 U13841 ( .A1(n11573), .A2(n13583), .ZN(n11328) );
  OAI211_X1 U13842 ( .C1(n9028), .C2(n13588), .A(n11328), .B(n11327), .ZN(
        P2_U3304) );
  AOI22_X1 U13843 ( .A1(n11329), .A2(n14462), .B1(n13105), .B2(n13147), .ZN(
        n11335) );
  INV_X1 U13844 ( .A(n11330), .ZN(n11334) );
  INV_X1 U13845 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n14860) );
  OAI22_X1 U13846 ( .A1(n14467), .A2(n14485), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14860), .ZN(n11332) );
  OAI22_X1 U13847 ( .A1(n13535), .A2(n14470), .B1(n14469), .B2(n13537), .ZN(
        n11331) );
  AOI211_X1 U13848 ( .C1(n14489), .C2(n14479), .A(n11332), .B(n11331), .ZN(
        n11333) );
  OAI21_X1 U13849 ( .B1(n11335), .B2(n11334), .A(n11333), .ZN(P2_U3213) );
  XNOR2_X1 U13850 ( .A(n11336), .B(n11340), .ZN(n11337) );
  NAND2_X1 U13851 ( .A1(n11337), .A2(n13407), .ZN(n11339) );
  AOI22_X1 U13852 ( .A1(n13400), .A2(n13402), .B1(n13401), .B2(n13147), .ZN(
        n11338) );
  NAND2_X1 U13853 ( .A1(n11339), .A2(n11338), .ZN(n14506) );
  INV_X1 U13854 ( .A(n14506), .ZN(n11347) );
  XOR2_X1 U13855 ( .A(n11341), .B(n11340), .Z(n14508) );
  OAI211_X1 U13856 ( .C1(n14505), .C2(n13526), .A(n13316), .B(n13425), .ZN(
        n14504) );
  INV_X1 U13857 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n11342) );
  OAI22_X1 U13858 ( .A1(n13429), .A2(n11342), .B1(n14483), .B2(n14877), .ZN(
        n11343) );
  AOI21_X1 U13859 ( .B1(n14480), .B2(n13440), .A(n11343), .ZN(n11344) );
  OAI21_X1 U13860 ( .B1(n14504), .B2(n13432), .A(n11344), .ZN(n11345) );
  AOI21_X1 U13861 ( .B1(n14508), .B2(n13442), .A(n11345), .ZN(n11346) );
  OAI21_X1 U13862 ( .B1(n13419), .B2(n11347), .A(n11346), .ZN(P2_U3249) );
  INV_X1 U13863 ( .A(n11482), .ZN(n11350) );
  OAI222_X1 U13864 ( .A1(n11348), .A2(P1_U3086), .B1(n11860), .B2(n11350), 
        .C1(n11483), .C2(n14247), .ZN(P1_U3331) );
  OAI222_X1 U13865 ( .A1(n13588), .A2(n15386), .B1(n13596), .B2(n11350), .C1(
        P2_U3088), .C2(n11349), .ZN(P2_U3303) );
  INV_X1 U13866 ( .A(n11351), .ZN(n11354) );
  OAI222_X1 U13867 ( .A1(n14370), .A2(n11354), .B1(n14368), .B2(n11353), .C1(
        P3_U3151), .C2(n11352), .ZN(P3_U3270) );
  INV_X1 U13868 ( .A(n12552), .ZN(n12406) );
  NAND2_X1 U13869 ( .A1(n11420), .A2(n12406), .ZN(n11355) );
  NAND2_X1 U13870 ( .A1(n11356), .A2(n11355), .ZN(n11358) );
  OR2_X1 U13871 ( .A1(n11420), .A2(n12406), .ZN(n11357) );
  NAND2_X1 U13872 ( .A1(n11358), .A2(n11357), .ZN(n11407) );
  OR2_X1 U13873 ( .A1(n12408), .A2(n12538), .ZN(n12048) );
  NAND2_X1 U13874 ( .A1(n12408), .A2(n12538), .ZN(n12047) );
  XNOR2_X1 U13875 ( .A(n11407), .B(n12045), .ZN(n11359) );
  AOI222_X1 U13876 ( .A1(n15056), .A2(n11359), .B1(n12552), .B2(n15038), .C1(
        n12550), .C2(n15052), .ZN(n11400) );
  MUX2_X1 U13877 ( .A(n15160), .B(n11400), .S(n15110), .Z(n11364) );
  INV_X1 U13878 ( .A(n12043), .ZN(n11360) );
  XNOR2_X1 U13879 ( .A(n11405), .B(n11406), .ZN(n11399) );
  AOI22_X1 U13880 ( .A1(n11399), .A2(n12989), .B1(n12988), .B2(n12408), .ZN(
        n11363) );
  NAND2_X1 U13881 ( .A1(n11364), .A2(n11363), .ZN(P3_U3432) );
  INV_X1 U13882 ( .A(P3_REG1_REG_14__SCAN_IN), .ZN(n11365) );
  MUX2_X1 U13883 ( .A(n11365), .B(n11400), .S(n15131), .Z(n11367) );
  AOI22_X1 U13884 ( .A1(n11399), .A2(n12914), .B1(n12913), .B2(n12408), .ZN(
        n11366) );
  NAND2_X1 U13885 ( .A1(n11367), .A2(n11366), .ZN(P3_U3473) );
  NAND2_X1 U13886 ( .A1(n12225), .A2(n11778), .ZN(n11369) );
  NAND2_X1 U13887 ( .A1(n13769), .A2(n11777), .ZN(n11368) );
  NAND2_X1 U13888 ( .A1(n11369), .A2(n11368), .ZN(n11370) );
  XNOR2_X1 U13889 ( .A(n11370), .B(n11745), .ZN(n11643) );
  AND2_X1 U13890 ( .A1(n13769), .A2(n6720), .ZN(n11371) );
  AOI21_X1 U13891 ( .B1(n12225), .B2(n11777), .A(n11371), .ZN(n11642) );
  XNOR2_X1 U13892 ( .A(n11643), .B(n11642), .ZN(n11379) );
  INV_X1 U13893 ( .A(n11372), .ZN(n11373) );
  NAND2_X1 U13894 ( .A1(n11374), .A2(n11373), .ZN(n11375) );
  INV_X1 U13895 ( .A(n11649), .ZN(n11377) );
  AOI21_X1 U13896 ( .B1(n11379), .B2(n11378), .A(n11377), .ZN(n11386) );
  NAND2_X1 U13897 ( .A1(n14537), .A2(n11380), .ZN(n11381) );
  OAI211_X1 U13898 ( .C1(n14542), .C2(n11383), .A(n11382), .B(n11381), .ZN(
        n11384) );
  AOI21_X1 U13899 ( .B1(n12225), .B2(n14533), .A(n11384), .ZN(n11385) );
  OAI21_X1 U13900 ( .B1(n11386), .B2(n13727), .A(n11385), .ZN(P1_U3236) );
  OAI21_X1 U13901 ( .B1(n11389), .B2(n11388), .A(n11387), .ZN(n11390) );
  NAND2_X1 U13902 ( .A1(n11390), .A2(n12533), .ZN(n11397) );
  NAND2_X1 U13903 ( .A1(n12525), .A2(n12553), .ZN(n11393) );
  INV_X1 U13904 ( .A(n11391), .ZN(n11392) );
  OAI211_X1 U13905 ( .C1(n12406), .C2(n12484), .A(n11393), .B(n11392), .ZN(
        n11394) );
  AOI21_X1 U13906 ( .B1(n12540), .B2(n11395), .A(n11394), .ZN(n11396) );
  OAI211_X1 U13907 ( .C1(n11398), .C2(n12544), .A(n11397), .B(n11396), .ZN(
        P3_U3164) );
  INV_X1 U13908 ( .A(n11399), .ZN(n11404) );
  INV_X1 U13909 ( .A(P3_REG2_REG_14__SCAN_IN), .ZN(n11401) );
  MUX2_X1 U13910 ( .A(n11401), .B(n11400), .S(n15049), .Z(n11403) );
  AOI22_X1 U13911 ( .A1(n12408), .A2(n14423), .B1(n15058), .B2(n12402), .ZN(
        n11402) );
  OAI211_X1 U13912 ( .C1(n12873), .C2(n11404), .A(n11403), .B(n11402), .ZN(
        P3_U3219) );
  OR2_X1 U13913 ( .A1(n12922), .A2(n12863), .ZN(n11963) );
  NAND2_X1 U13914 ( .A1(n12922), .A2(n12863), .ZN(n12055) );
  XNOR2_X1 U13915 ( .A(n11847), .B(n11935), .ZN(n13000) );
  INV_X1 U13916 ( .A(n12851), .ZN(n12470) );
  NAND2_X1 U13917 ( .A1(n11407), .A2(n11406), .ZN(n11409) );
  NAND2_X1 U13918 ( .A1(n12408), .A2(n12551), .ZN(n11408) );
  NAND2_X1 U13919 ( .A1(n11409), .A2(n11408), .ZN(n11799) );
  XNOR2_X1 U13920 ( .A(n11799), .B(n11935), .ZN(n11410) );
  INV_X1 U13921 ( .A(n15056), .ZN(n15043) );
  OAI222_X1 U13922 ( .A1(n12864), .A2(n12538), .B1(n12866), .B2(n12470), .C1(
        n11410), .C2(n15043), .ZN(n12921) );
  NAND2_X1 U13923 ( .A1(n12921), .A2(n15049), .ZN(n11414) );
  INV_X1 U13924 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n15293) );
  INV_X1 U13925 ( .A(n12541), .ZN(n11411) );
  OAI22_X1 U13926 ( .A1(n15049), .A2(n15293), .B1(n11411), .B2(n12868), .ZN(
        n11412) );
  AOI21_X1 U13927 ( .B1(n12922), .B2(n14423), .A(n11412), .ZN(n11413) );
  OAI211_X1 U13928 ( .C1(n12873), .C2(n13000), .A(n11414), .B(n11413), .ZN(
        P3_U3218) );
  XNOR2_X1 U13929 ( .A(n11415), .B(n12552), .ZN(n11416) );
  XNOR2_X1 U13930 ( .A(n11417), .B(n11416), .ZN(n11425) );
  AND2_X1 U13931 ( .A1(P3_U3151), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n12575) );
  AOI21_X1 U13932 ( .B1(n12535), .B2(n12551), .A(n12575), .ZN(n11418) );
  OAI21_X1 U13933 ( .B1(n11419), .B2(n12537), .A(n11418), .ZN(n11422) );
  NOR2_X1 U13934 ( .A1(n11420), .A2(n12544), .ZN(n11421) );
  AOI211_X1 U13935 ( .C1(n11423), .C2(n12540), .A(n11422), .B(n11421), .ZN(
        n11424) );
  OAI21_X1 U13936 ( .B1(n11425), .B2(n12507), .A(n11424), .ZN(P3_U3174) );
  INV_X1 U13937 ( .A(n11474), .ZN(n11429) );
  OAI222_X1 U13938 ( .A1(n13594), .A2(n11427), .B1(n13596), .B2(n11429), .C1(
        P2_U3088), .C2(n11426), .ZN(P2_U3302) );
  INV_X1 U13939 ( .A(n11428), .ZN(n11430) );
  OAI222_X1 U13940 ( .A1(n11430), .A2(P1_U3086), .B1(n11860), .B2(n11429), 
        .C1(n15212), .C2(n14247), .ZN(P1_U3330) );
  NOR2_X1 U13941 ( .A1(n14467), .A2(n13428), .ZN(n11434) );
  AND2_X1 U13942 ( .A1(n13146), .A2(n13401), .ZN(n11431) );
  AOI21_X1 U13943 ( .B1(n13145), .B2(n13402), .A(n11431), .ZN(n13421) );
  OAI22_X1 U13944 ( .A1(n13110), .A2(n13421), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n11432), .ZN(n11433) );
  AOI211_X1 U13945 ( .C1(n14498), .C2(n14479), .A(n11434), .B(n11433), .ZN(
        n11440) );
  INV_X1 U13946 ( .A(n11435), .ZN(n11438) );
  OAI22_X1 U13947 ( .A1(n11436), .A2(n14474), .B1(n13537), .B2(n13124), .ZN(
        n11437) );
  NAND3_X1 U13948 ( .A1(n14476), .A2(n11438), .A3(n11437), .ZN(n11439) );
  OAI211_X1 U13949 ( .C1(n11441), .C2(n14474), .A(n11440), .B(n11439), .ZN(
        P2_U3200) );
  OAI22_X1 U13950 ( .A1(n11445), .A2(n11444), .B1(n11443), .B2(n11442), .ZN(
        n11446) );
  NAND2_X1 U13951 ( .A1(n14867), .A2(n11446), .ZN(n11447) );
  XNOR2_X1 U13952 ( .A(n11446), .B(n11453), .ZN(n14871) );
  NAND2_X1 U13953 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n14871), .ZN(n14869) );
  NAND2_X1 U13954 ( .A1(n11447), .A2(n14869), .ZN(n11450) );
  NAND2_X1 U13955 ( .A1(n11455), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n13195) );
  OAI21_X1 U13956 ( .B1(n11455), .B2(P2_REG2_REG_16__SCAN_IN), .A(n13195), 
        .ZN(n11448) );
  INV_X1 U13957 ( .A(n11448), .ZN(n11449) );
  OAI21_X1 U13958 ( .B1(n11450), .B2(n11449), .A(n14870), .ZN(n11462) );
  XOR2_X1 U13959 ( .A(n14867), .B(n11454), .Z(n14864) );
  OAI21_X1 U13960 ( .B1(n11454), .B2(n11453), .A(n14861), .ZN(n11457) );
  INV_X1 U13961 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n14509) );
  MUX2_X1 U13962 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n14509), .S(n11455), .Z(
        n11456) );
  NAND2_X1 U13963 ( .A1(n11457), .A2(n11456), .ZN(n13189) );
  OAI211_X1 U13964 ( .C1(n11457), .C2(n11456), .A(n13189), .B(n14853), .ZN(
        n11461) );
  NAND2_X1 U13965 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(P2_U3088), .ZN(n14481)
         );
  INV_X1 U13966 ( .A(n14481), .ZN(n11459) );
  NOR2_X1 U13967 ( .A1(n14834), .A2(n13190), .ZN(n11458) );
  AOI211_X1 U13968 ( .C1(P2_ADDR_REG_16__SCAN_IN), .C2(n14789), .A(n11459), 
        .B(n11458), .ZN(n11460) );
  OAI211_X1 U13969 ( .C1(n13202), .C2(n11462), .A(n11461), .B(n11460), .ZN(
        P2_U3230) );
  NOR2_X1 U13970 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(n11817), .ZN(n11465) );
  NAND2_X1 U13971 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(n13595), .ZN(n11464) );
  AOI222_X1 U13972 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(n6517), .B1(
        P1_DATAO_REG_28__SCAN_IN), .B2(n11772), .C1(n11824), .C2(n11772), .ZN(
        n11893) );
  AOI22_X1 U13973 ( .A1(P2_DATAO_REG_29__SCAN_IN), .A2(
        P1_DATAO_REG_29__SCAN_IN), .B1(n13581), .B2(n12386), .ZN(n11892) );
  OAI222_X1 U13974 ( .A1(n14370), .A2(n11832), .B1(P3_U3151), .B2(n11466), 
        .C1(n11833), .C2(n14368), .ZN(P3_U3266) );
  INV_X1 U13975 ( .A(n11595), .ZN(n13592) );
  OAI222_X1 U13976 ( .A1(P1_U3086), .A2(n13875), .B1(n11860), .B2(n13592), 
        .C1(n11817), .C2(n14247), .ZN(P1_U3328) );
  NAND2_X1 U13977 ( .A1(n11783), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n11473) );
  INV_X1 U13978 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n11467) );
  OR2_X1 U13979 ( .A1(n11784), .A2(n11467), .ZN(n11472) );
  OAI21_X1 U13980 ( .B1(P1_REG3_REG_25__SCAN_IN), .B2(n11468), .A(n11588), 
        .ZN(n13946) );
  OR2_X1 U13981 ( .A1(n11600), .A2(n13946), .ZN(n11471) );
  INV_X1 U13982 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n11469) );
  OR2_X1 U13983 ( .A1(n6526), .A2(n11469), .ZN(n11470) );
  NAND4_X1 U13984 ( .A1(n11473), .A2(n11472), .A3(n11471), .A4(n11470), .ZN(
        n13756) );
  INV_X1 U13985 ( .A(n13756), .ZN(n11583) );
  OR2_X1 U13986 ( .A1(n12317), .A2(n15212), .ZN(n11475) );
  NAND2_X1 U13987 ( .A1(n12321), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n11481) );
  INV_X1 U13988 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n15308) );
  OR2_X1 U13989 ( .A1(n6540), .A2(n15308), .ZN(n11480) );
  OAI21_X1 U13990 ( .B1(P1_REG3_REG_24__SCAN_IN), .B2(n11477), .A(n11476), 
        .ZN(n13964) );
  OR2_X1 U13991 ( .A1(n11600), .A2(n13964), .ZN(n11479) );
  INV_X1 U13992 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n13965) );
  OR2_X1 U13993 ( .A1(n6526), .A2(n13965), .ZN(n11478) );
  NAND4_X1 U13994 ( .A1(n11481), .A2(n11480), .A3(n11479), .A4(n11478), .ZN(
        n13757) );
  INV_X1 U13995 ( .A(n13757), .ZN(n11619) );
  NAND2_X1 U13996 ( .A1(n11482), .A2(n10677), .ZN(n11485) );
  OR2_X1 U13997 ( .A1(n12317), .A2(n11483), .ZN(n11484) );
  INV_X1 U13998 ( .A(n14165), .ZN(n13963) );
  NAND2_X1 U13999 ( .A1(n11486), .A2(n10677), .ZN(n11489) );
  OR2_X1 U14000 ( .A1(n12317), .A2(n11487), .ZN(n11488) );
  AND2_X1 U14001 ( .A1(n11554), .A2(n13637), .ZN(n11490) );
  OR2_X1 U14002 ( .A1(n11561), .A2(n11490), .ZN(n13636) );
  AOI22_X1 U14003 ( .A1(n11783), .A2(P1_REG1_REG_21__SCAN_IN), .B1(n12321), 
        .B2(P1_REG0_REG_21__SCAN_IN), .ZN(n11492) );
  INV_X1 U14004 ( .A(n6526), .ZN(n12320) );
  NAND2_X1 U14005 ( .A1(n12320), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n11491) );
  OAI211_X1 U14006 ( .C1(n13636), .C2(n11600), .A(n11492), .B(n11491), .ZN(
        n13760) );
  NAND2_X1 U14007 ( .A1(n14534), .A2(n13766), .ZN(n11493) );
  NAND2_X1 U14008 ( .A1(n11494), .A2(n10677), .ZN(n11496) );
  AOI22_X1 U14009 ( .A1(n11535), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n11533), 
        .B2(n14615), .ZN(n11495) );
  OR2_X1 U14010 ( .A1(n14115), .A2(n13663), .ZN(n12252) );
  NAND2_X1 U14011 ( .A1(n14115), .A2(n13663), .ZN(n14082) );
  NAND2_X1 U14012 ( .A1(n12252), .A2(n14082), .ZN(n14105) );
  INV_X1 U14013 ( .A(n14105), .ZN(n14098) );
  OR2_X2 U14014 ( .A1(n14103), .A2(n14098), .ZN(n14104) );
  INV_X1 U14015 ( .A(n13663), .ZN(n11497) );
  OR2_X1 U14016 ( .A1(n14115), .A2(n11497), .ZN(n11498) );
  NAND2_X1 U14017 ( .A1(n11499), .A2(n10677), .ZN(n11501) );
  AOI22_X1 U14018 ( .A1(n11535), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n11533), 
        .B2(n13820), .ZN(n11500) );
  INV_X1 U14019 ( .A(n14215), .ZN(n12251) );
  NAND2_X1 U14020 ( .A1(n11783), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n11508) );
  INV_X1 U14021 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n11502) );
  OR2_X1 U14022 ( .A1(n11784), .A2(n11502), .ZN(n11507) );
  NAND2_X1 U14023 ( .A1(n11503), .A2(n15369), .ZN(n11504) );
  NAND2_X1 U14024 ( .A1(n11523), .A2(n11504), .ZN(n14088) );
  OR2_X1 U14025 ( .A1(n11600), .A2(n14088), .ZN(n11506) );
  INV_X1 U14026 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n13827) );
  OR2_X1 U14027 ( .A1(n6526), .A2(n13827), .ZN(n11505) );
  INV_X1 U14028 ( .A(n13746), .ZN(n13765) );
  XNOR2_X1 U14029 ( .A(n12251), .B(n13765), .ZN(n14085) );
  INV_X1 U14030 ( .A(n14085), .ZN(n11610) );
  NAND2_X1 U14031 ( .A1(n14215), .A2(n13746), .ZN(n11509) );
  NAND2_X1 U14032 ( .A1(n11511), .A2(n10677), .ZN(n11513) );
  AOI22_X1 U14033 ( .A1(n11535), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n11533), 
        .B2(n13844), .ZN(n11512) );
  NAND2_X1 U14034 ( .A1(n11783), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n11519) );
  INV_X1 U14035 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n11514) );
  XNOR2_X1 U14036 ( .A(n11523), .B(n11514), .ZN(n14071) );
  OR2_X1 U14037 ( .A1(n11600), .A2(n14071), .ZN(n11518) );
  INV_X1 U14038 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n11515) );
  OR2_X1 U14039 ( .A1(n11784), .A2(n11515), .ZN(n11517) );
  INV_X1 U14040 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n13831) );
  OR2_X1 U14041 ( .A1(n6526), .A2(n13831), .ZN(n11516) );
  NAND4_X1 U14042 ( .A1(n11519), .A2(n11518), .A3(n11517), .A4(n11516), .ZN(
        n13764) );
  NOR2_X1 U14043 ( .A1(n14209), .A2(n13764), .ZN(n12335) );
  NAND2_X1 U14044 ( .A1(n14209), .A2(n13764), .ZN(n12336) );
  NAND2_X1 U14045 ( .A1(n11520), .A2(n10677), .ZN(n11522) );
  AOI22_X1 U14046 ( .A1(n11535), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n11533), 
        .B2(n13858), .ZN(n11521) );
  INV_X1 U14047 ( .A(n11523), .ZN(n11524) );
  AOI21_X1 U14048 ( .B1(n11524), .B2(P1_REG3_REG_17__SCAN_IN), .A(
        P1_REG3_REG_18__SCAN_IN), .ZN(n11525) );
  OR2_X1 U14049 ( .A1(n11525), .A2(n11540), .ZN(n14060) );
  INV_X1 U14050 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n14061) );
  OR2_X1 U14051 ( .A1(n6526), .A2(n14061), .ZN(n11526) );
  OAI21_X1 U14052 ( .B1(n11600), .B2(n14060), .A(n11526), .ZN(n11530) );
  INV_X1 U14053 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n13848) );
  INV_X1 U14054 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n11527) );
  OR2_X1 U14055 ( .A1(n11784), .A2(n11527), .ZN(n11528) );
  OAI21_X1 U14056 ( .B1(n6539), .B2(n13848), .A(n11528), .ZN(n11529) );
  AND2_X1 U14057 ( .A1(n14204), .A2(n13763), .ZN(n11531) );
  NAND2_X1 U14058 ( .A1(n11532), .A2(n10677), .ZN(n11537) );
  AOI22_X1 U14059 ( .A1(n11535), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n11534), 
        .B2(n11533), .ZN(n11536) );
  INV_X1 U14060 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n11539) );
  NAND2_X1 U14061 ( .A1(n12321), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n11538) );
  OAI21_X1 U14062 ( .B1(n6540), .B2(n11539), .A(n11538), .ZN(n11544) );
  OR2_X1 U14063 ( .A1(n11540), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n11541) );
  NAND2_X1 U14064 ( .A1(n11552), .A2(n11541), .ZN(n14041) );
  NAND2_X1 U14065 ( .A1(n12320), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n11542) );
  OAI21_X1 U14066 ( .B1(n14041), .B2(n11600), .A(n11542), .ZN(n11543) );
  INV_X1 U14067 ( .A(n13762), .ZN(n11545) );
  OR2_X1 U14068 ( .A1(n14197), .A2(n11545), .ZN(n12266) );
  NAND2_X1 U14069 ( .A1(n14197), .A2(n11545), .ZN(n14019) );
  NAND2_X1 U14070 ( .A1(n12266), .A2(n14019), .ZN(n14048) );
  OR2_X1 U14071 ( .A1(n14197), .A2(n13762), .ZN(n11546) );
  NAND2_X1 U14072 ( .A1(n11548), .A2(n10677), .ZN(n11551) );
  OR2_X1 U14073 ( .A1(n12317), .A2(n11549), .ZN(n11550) );
  NAND2_X1 U14074 ( .A1(n11552), .A2(n15196), .ZN(n11553) );
  NAND2_X1 U14075 ( .A1(n11554), .A2(n11553), .ZN(n14024) );
  OR2_X1 U14076 ( .A1(n14024), .A2(n11600), .ZN(n11559) );
  NAND2_X1 U14077 ( .A1(n12321), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n11556) );
  NAND2_X1 U14078 ( .A1(n12320), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n11555) );
  AND2_X1 U14079 ( .A1(n11556), .A2(n11555), .ZN(n11558) );
  NAND2_X1 U14080 ( .A1(n11783), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n11557) );
  XNOR2_X1 U14081 ( .A(n14029), .B(n13627), .ZN(n12358) );
  OR2_X1 U14082 ( .A1(n14192), .A2(n13627), .ZN(n11560) );
  XNOR2_X1 U14083 ( .A(n14013), .B(n13760), .ZN(n14006) );
  OR2_X1 U14084 ( .A1(n11561), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n11563) );
  NAND2_X1 U14085 ( .A1(n11563), .A2(n11562), .ZN(n13713) );
  OR2_X1 U14086 ( .A1(n13713), .A2(n11600), .ZN(n11569) );
  INV_X1 U14087 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n11566) );
  NAND2_X1 U14088 ( .A1(n12320), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n11565) );
  NAND2_X1 U14089 ( .A1(n12321), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n11564) );
  OAI211_X1 U14090 ( .C1(n6539), .C2(n11566), .A(n11565), .B(n11564), .ZN(
        n11567) );
  INV_X1 U14091 ( .A(n11567), .ZN(n11568) );
  NAND2_X1 U14092 ( .A1(n11569), .A2(n11568), .ZN(n13759) );
  NAND2_X1 U14093 ( .A1(n11570), .A2(n7626), .ZN(n11571) );
  XNOR2_X1 U14094 ( .A(n11571), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n14250) );
  OR2_X1 U14095 ( .A1(n12317), .A2(n11574), .ZN(n11575) );
  NAND2_X1 U14096 ( .A1(n11783), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n11582) );
  INV_X1 U14097 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n11576) );
  OR2_X1 U14098 ( .A1(n11784), .A2(n11576), .ZN(n11581) );
  OAI21_X1 U14099 ( .B1(P1_REG3_REG_23__SCAN_IN), .B2(n11578), .A(n11577), 
        .ZN(n13978) );
  OR2_X1 U14100 ( .A1(n11600), .A2(n13978), .ZN(n11580) );
  INV_X1 U14101 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n13977) );
  OR2_X1 U14102 ( .A1(n6526), .A2(n13977), .ZN(n11579) );
  NAND4_X1 U14103 ( .A1(n11582), .A2(n11581), .A3(n11580), .A4(n11579), .ZN(
        n13758) );
  INV_X1 U14104 ( .A(n13758), .ZN(n11618) );
  XNOR2_X1 U14105 ( .A(n14165), .B(n11619), .ZN(n13957) );
  NAND2_X1 U14106 ( .A1(n13593), .A2(n10677), .ZN(n11585) );
  OR2_X1 U14107 ( .A1(n12317), .A2(n15197), .ZN(n11584) );
  NAND2_X1 U14108 ( .A1(n11783), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n11594) );
  INV_X1 U14109 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n11586) );
  OR2_X1 U14110 ( .A1(n11784), .A2(n11586), .ZN(n11593) );
  INV_X1 U14111 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n11587) );
  NAND2_X1 U14112 ( .A1(n11588), .A2(n11587), .ZN(n11589) );
  NAND2_X1 U14113 ( .A1(n11599), .A2(n11589), .ZN(n13934) );
  OR2_X1 U14114 ( .A1(n11600), .A2(n13934), .ZN(n11592) );
  INV_X1 U14115 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n11590) );
  OR2_X1 U14116 ( .A1(n6526), .A2(n11590), .ZN(n11591) );
  NAND4_X1 U14117 ( .A1(n11594), .A2(n11593), .A3(n11592), .A4(n11591), .ZN(
        n13755) );
  INV_X1 U14118 ( .A(n13755), .ZN(n11621) );
  NAND2_X1 U14119 ( .A1(n11595), .A2(n10677), .ZN(n11597) );
  OR2_X1 U14120 ( .A1(n12317), .A2(n11817), .ZN(n11596) );
  NAND2_X1 U14121 ( .A1(n11783), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n11605) );
  INV_X1 U14122 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n11598) );
  OR2_X1 U14123 ( .A1(n11784), .A2(n11598), .ZN(n11604) );
  XNOR2_X1 U14124 ( .A(n11599), .B(n13607), .ZN(n13606) );
  OR2_X1 U14125 ( .A1(n11600), .A2(n13606), .ZN(n11603) );
  INV_X1 U14126 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n11631) );
  OR2_X1 U14127 ( .A1(n6526), .A2(n11631), .ZN(n11602) );
  NAND4_X1 U14128 ( .A1(n11605), .A2(n11604), .A3(n11603), .A4(n11602), .ZN(
        n13908) );
  NAND2_X1 U14129 ( .A1(n11608), .A2(n12247), .ZN(n14097) );
  OR2_X1 U14130 ( .A1(n14534), .A2(n11609), .ZN(n14096) );
  AND2_X1 U14131 ( .A1(n14096), .A2(n12252), .ZN(n14081) );
  AND2_X1 U14132 ( .A1(n14081), .A2(n14085), .ZN(n11611) );
  OR2_X1 U14133 ( .A1(n14215), .A2(n13765), .ZN(n11612) );
  NAND2_X1 U14134 ( .A1(n14084), .A2(n11612), .ZN(n14067) );
  INV_X1 U14135 ( .A(n13764), .ZN(n11614) );
  OR2_X1 U14136 ( .A1(n14209), .A2(n11614), .ZN(n11613) );
  NAND2_X1 U14137 ( .A1(n14209), .A2(n11614), .ZN(n11615) );
  XNOR2_X1 U14138 ( .A(n14204), .B(n13763), .ZN(n14056) );
  INV_X1 U14139 ( .A(n13763), .ZN(n13626) );
  AND2_X1 U14140 ( .A1(n14030), .A2(n14019), .ZN(n11616) );
  INV_X1 U14141 ( .A(n13627), .ZN(n13761) );
  NAND2_X1 U14142 ( .A1(n14192), .A2(n13761), .ZN(n11617) );
  NAND2_X1 U14143 ( .A1(n14020), .A2(n11617), .ZN(n14001) );
  XNOR2_X1 U14144 ( .A(n13981), .B(n13758), .ZN(n13976) );
  INV_X1 U14145 ( .A(n14153), .ZN(n13938) );
  OAI21_X1 U14146 ( .B1(n11622), .B2(n12361), .A(n13910), .ZN(n11626) );
  NAND2_X1 U14147 ( .A1(n13913), .A2(n13732), .ZN(n11624) );
  NAND2_X1 U14148 ( .A1(n13755), .A2(n13897), .ZN(n11623) );
  AND2_X1 U14149 ( .A1(n11624), .A2(n11623), .ZN(n13608) );
  INV_X1 U14150 ( .A(n13608), .ZN(n11625) );
  INV_X1 U14151 ( .A(n13891), .ZN(n13909) );
  NAND2_X1 U14152 ( .A1(n14108), .A2(n14215), .ZN(n14086) );
  OR2_X2 U14153 ( .A1(n14026), .A2(n14013), .ZN(n14010) );
  INV_X1 U14154 ( .A(n11630), .ZN(n13933) );
  OAI211_X1 U14155 ( .C1(n13909), .C2(n13933), .A(n14109), .B(n6572), .ZN(
        n14146) );
  OAI22_X1 U14156 ( .A1(n14680), .A2(n11631), .B1(n13606), .B2(n14659), .ZN(
        n11632) );
  AOI21_X1 U14157 ( .B1(n13891), .B2(n14662), .A(n11632), .ZN(n11633) );
  OAI21_X1 U14158 ( .B1(n14146), .B2(n14117), .A(n11633), .ZN(n11634) );
  AOI21_X1 U14159 ( .B1(n14145), .B2(n14670), .A(n11634), .ZN(n11635) );
  OAI21_X1 U14160 ( .B1(n14149), .B2(n14674), .A(n11635), .ZN(P1_U3266) );
  INV_X1 U14161 ( .A(n12315), .ZN(n11638) );
  OAI222_X1 U14162 ( .A1(n13596), .A2(n11638), .B1(P2_U3088), .B2(n6538), .C1(
        n11636), .C2(n13594), .ZN(P2_U3297) );
  OAI222_X1 U14163 ( .A1(n11860), .A2(n11638), .B1(n11637), .B2(P1_U3086), 
        .C1(n12316), .C2(n14247), .ZN(P1_U3325) );
  AOI22_X1 U14164 ( .A1(n14204), .A2(n11777), .B1(n6720), .B2(n13763), .ZN(
        n11691) );
  NAND2_X1 U14165 ( .A1(n14204), .A2(n11778), .ZN(n11640) );
  NAND2_X1 U14166 ( .A1(n13763), .A2(n11777), .ZN(n11639) );
  NAND2_X1 U14167 ( .A1(n11640), .A2(n11639), .ZN(n11641) );
  XNOR2_X1 U14168 ( .A(n11641), .B(n11775), .ZN(n11689) );
  INV_X1 U14169 ( .A(n11689), .ZN(n11690) );
  NAND2_X1 U14170 ( .A1(n11643), .A2(n11642), .ZN(n13641) );
  NAND2_X1 U14171 ( .A1(n12235), .A2(n11778), .ZN(n11645) );
  NAND2_X1 U14172 ( .A1(n13768), .A2(n11777), .ZN(n11644) );
  NAND2_X1 U14173 ( .A1(n11645), .A2(n11644), .ZN(n11646) );
  XNOR2_X1 U14174 ( .A(n11646), .B(n11775), .ZN(n11652) );
  AND2_X1 U14175 ( .A1(n13768), .A2(n6720), .ZN(n11647) );
  AOI21_X1 U14176 ( .B1(n12235), .B2(n11777), .A(n11647), .ZN(n11650) );
  XNOR2_X1 U14177 ( .A(n11652), .B(n11650), .ZN(n13643) );
  AND2_X1 U14178 ( .A1(n13641), .A2(n13643), .ZN(n11648) );
  INV_X1 U14179 ( .A(n11650), .ZN(n11651) );
  NAND2_X1 U14180 ( .A1(n11652), .A2(n11651), .ZN(n11653) );
  NAND2_X1 U14181 ( .A1(n13706), .A2(n11778), .ZN(n11655) );
  NAND2_X1 U14182 ( .A1(n13767), .A2(n11777), .ZN(n11654) );
  NAND2_X1 U14183 ( .A1(n11655), .A2(n11654), .ZN(n11656) );
  XNOR2_X1 U14184 ( .A(n11656), .B(n11775), .ZN(n11660) );
  AND2_X1 U14185 ( .A1(n13767), .A2(n6720), .ZN(n11657) );
  AOI21_X1 U14186 ( .B1(n13706), .B2(n11777), .A(n11657), .ZN(n11658) );
  XNOR2_X1 U14187 ( .A(n11660), .B(n11658), .ZN(n13699) );
  INV_X1 U14188 ( .A(n11658), .ZN(n11659) );
  NAND2_X1 U14189 ( .A1(n11660), .A2(n11659), .ZN(n11661) );
  NAND2_X1 U14190 ( .A1(n14534), .A2(n11778), .ZN(n11664) );
  NAND2_X1 U14191 ( .A1(n13766), .A2(n11777), .ZN(n11663) );
  NAND2_X1 U14192 ( .A1(n11664), .A2(n11663), .ZN(n11665) );
  XNOR2_X1 U14193 ( .A(n11665), .B(n11745), .ZN(n11668) );
  AND2_X1 U14194 ( .A1(n13766), .A2(n6720), .ZN(n11666) );
  AOI21_X1 U14195 ( .B1(n14534), .B2(n11777), .A(n11666), .ZN(n11667) );
  XNOR2_X1 U14196 ( .A(n11668), .B(n11667), .ZN(n14531) );
  NAND2_X1 U14197 ( .A1(n14115), .A2(n11778), .ZN(n11670) );
  OR2_X1 U14198 ( .A1(n13663), .A2(n11701), .ZN(n11669) );
  NAND2_X1 U14199 ( .A1(n11670), .A2(n11669), .ZN(n11671) );
  INV_X1 U14200 ( .A(n13742), .ZN(n11674) );
  NOR2_X1 U14201 ( .A1(n13663), .A2(n11700), .ZN(n11672) );
  AOI21_X1 U14202 ( .B1(n14115), .B2(n11777), .A(n11672), .ZN(n13741) );
  INV_X1 U14203 ( .A(n13741), .ZN(n11673) );
  OAI22_X1 U14204 ( .A1(n14215), .A2(n11702), .B1(n13746), .B2(n11701), .ZN(
        n11675) );
  XNOR2_X1 U14205 ( .A(n11675), .B(n11775), .ZN(n11677) );
  OAI22_X1 U14206 ( .A1(n14215), .A2(n11701), .B1(n13746), .B2(n11700), .ZN(
        n11676) );
  OR2_X1 U14207 ( .A1(n11677), .A2(n11676), .ZN(n13670) );
  NAND2_X1 U14208 ( .A1(n11677), .A2(n11676), .ZN(n11678) );
  AND2_X1 U14209 ( .A1(n13670), .A2(n11678), .ZN(n13660) );
  NAND2_X1 U14210 ( .A1(n14209), .A2(n11778), .ZN(n11680) );
  NAND2_X1 U14211 ( .A1(n13764), .A2(n11777), .ZN(n11679) );
  NAND2_X1 U14212 ( .A1(n11680), .A2(n11679), .ZN(n11681) );
  XNOR2_X1 U14213 ( .A(n11681), .B(n11745), .ZN(n11683) );
  AND2_X1 U14214 ( .A1(n13764), .A2(n6720), .ZN(n11682) );
  AOI21_X1 U14215 ( .B1(n14209), .B2(n11777), .A(n11682), .ZN(n11684) );
  NAND2_X1 U14216 ( .A1(n11683), .A2(n11684), .ZN(n11688) );
  INV_X1 U14217 ( .A(n11683), .ZN(n11686) );
  INV_X1 U14218 ( .A(n11684), .ZN(n11685) );
  NAND2_X1 U14219 ( .A1(n11686), .A2(n11685), .ZN(n11687) );
  NAND2_X1 U14220 ( .A1(n11688), .A2(n11687), .ZN(n13669) );
  XOR2_X1 U14221 ( .A(n11691), .B(n11689), .Z(n13721) );
  NAND2_X1 U14222 ( .A1(n14197), .A2(n11778), .ZN(n11693) );
  NAND2_X1 U14223 ( .A1(n13762), .A2(n11777), .ZN(n11692) );
  NAND2_X1 U14224 ( .A1(n11693), .A2(n11692), .ZN(n11694) );
  XNOR2_X1 U14225 ( .A(n11694), .B(n11775), .ZN(n11696) );
  AND2_X1 U14226 ( .A1(n13762), .A2(n6720), .ZN(n11695) );
  AOI21_X1 U14227 ( .B1(n14197), .B2(n9413), .A(n11695), .ZN(n11697) );
  XNOR2_X1 U14228 ( .A(n11696), .B(n11697), .ZN(n13624) );
  INV_X1 U14229 ( .A(n11697), .ZN(n11698) );
  OAI22_X1 U14230 ( .A1(n14192), .A2(n11701), .B1(n13627), .B2(n11700), .ZN(
        n11704) );
  OAI22_X1 U14231 ( .A1(n14192), .A2(n11702), .B1(n13627), .B2(n11701), .ZN(
        n11703) );
  XNOR2_X1 U14232 ( .A(n11703), .B(n11775), .ZN(n11705) );
  XOR2_X1 U14233 ( .A(n11704), .B(n11705), .Z(n13692) );
  AND2_X1 U14234 ( .A1(n11705), .A2(n11704), .ZN(n11706) );
  NAND2_X1 U14235 ( .A1(n14013), .A2(n11778), .ZN(n11708) );
  NAND2_X1 U14236 ( .A1(n13760), .A2(n11777), .ZN(n11707) );
  NAND2_X1 U14237 ( .A1(n11708), .A2(n11707), .ZN(n11709) );
  XNOR2_X1 U14238 ( .A(n11709), .B(n11775), .ZN(n11713) );
  NAND2_X1 U14239 ( .A1(n14013), .A2(n11777), .ZN(n11711) );
  NAND2_X1 U14240 ( .A1(n13760), .A2(n6720), .ZN(n11710) );
  NAND2_X1 U14241 ( .A1(n11711), .A2(n11710), .ZN(n11712) );
  NOR2_X1 U14242 ( .A1(n11713), .A2(n11712), .ZN(n11714) );
  AOI21_X1 U14243 ( .B1(n11713), .B2(n11712), .A(n11714), .ZN(n13633) );
  NAND2_X1 U14244 ( .A1(n6518), .A2(n13633), .ZN(n13632) );
  INV_X1 U14245 ( .A(n11714), .ZN(n11715) );
  NAND2_X1 U14246 ( .A1(n13632), .A2(n11715), .ZN(n13710) );
  NAND2_X1 U14247 ( .A1(n12276), .A2(n11778), .ZN(n11717) );
  NAND2_X1 U14248 ( .A1(n13759), .A2(n10439), .ZN(n11716) );
  NAND2_X1 U14249 ( .A1(n11717), .A2(n11716), .ZN(n11718) );
  XNOR2_X1 U14250 ( .A(n11718), .B(n11775), .ZN(n11722) );
  NAND2_X1 U14251 ( .A1(n12276), .A2(n11777), .ZN(n11720) );
  NAND2_X1 U14252 ( .A1(n13759), .A2(n6720), .ZN(n11719) );
  NAND2_X1 U14253 ( .A1(n11720), .A2(n11719), .ZN(n11721) );
  NOR2_X1 U14254 ( .A1(n11722), .A2(n11721), .ZN(n11723) );
  AOI21_X1 U14255 ( .B1(n11722), .B2(n11721), .A(n11723), .ZN(n13711) );
  INV_X1 U14256 ( .A(n11723), .ZN(n11724) );
  NAND2_X1 U14257 ( .A1(n13981), .A2(n11778), .ZN(n11726) );
  NAND2_X1 U14258 ( .A1(n13758), .A2(n11777), .ZN(n11725) );
  NAND2_X1 U14259 ( .A1(n11726), .A2(n11725), .ZN(n11727) );
  XNOR2_X1 U14260 ( .A(n11727), .B(n11775), .ZN(n11731) );
  NAND2_X1 U14261 ( .A1(n13981), .A2(n11777), .ZN(n11729) );
  NAND2_X1 U14262 ( .A1(n13758), .A2(n6720), .ZN(n11728) );
  NAND2_X1 U14263 ( .A1(n11729), .A2(n11728), .ZN(n11730) );
  NOR2_X1 U14264 ( .A1(n11731), .A2(n11730), .ZN(n11732) );
  AOI21_X1 U14265 ( .B1(n11731), .B2(n11730), .A(n11732), .ZN(n13615) );
  NAND2_X2 U14266 ( .A1(n13614), .A2(n13615), .ZN(n13686) );
  INV_X1 U14267 ( .A(n11732), .ZN(n13685) );
  NAND2_X1 U14268 ( .A1(n14165), .A2(n11778), .ZN(n11734) );
  NAND2_X1 U14269 ( .A1(n13757), .A2(n11777), .ZN(n11733) );
  NAND2_X1 U14270 ( .A1(n11734), .A2(n11733), .ZN(n11735) );
  XNOR2_X1 U14271 ( .A(n11735), .B(n11745), .ZN(n11737) );
  AND2_X1 U14272 ( .A1(n13757), .A2(n6720), .ZN(n11736) );
  AOI21_X1 U14273 ( .B1(n14165), .B2(n11777), .A(n11736), .ZN(n11738) );
  NAND2_X1 U14274 ( .A1(n11737), .A2(n11738), .ZN(n11742) );
  INV_X1 U14275 ( .A(n11737), .ZN(n11740) );
  INV_X1 U14276 ( .A(n11738), .ZN(n11739) );
  NAND2_X1 U14277 ( .A1(n11740), .A2(n11739), .ZN(n11741) );
  NAND2_X1 U14278 ( .A1(n11742), .A2(n11741), .ZN(n13684) );
  INV_X1 U14279 ( .A(n11742), .ZN(n13655) );
  NAND2_X1 U14280 ( .A1(n14159), .A2(n11778), .ZN(n11744) );
  NAND2_X1 U14281 ( .A1(n13756), .A2(n11777), .ZN(n11743) );
  NAND2_X1 U14282 ( .A1(n11744), .A2(n11743), .ZN(n11746) );
  XNOR2_X1 U14283 ( .A(n11746), .B(n11745), .ZN(n11748) );
  AND2_X1 U14284 ( .A1(n13756), .A2(n6720), .ZN(n11747) );
  AOI21_X1 U14285 ( .B1(n14159), .B2(n10439), .A(n11747), .ZN(n11749) );
  NAND2_X1 U14286 ( .A1(n11748), .A2(n11749), .ZN(n11753) );
  INV_X1 U14287 ( .A(n11748), .ZN(n11751) );
  INV_X1 U14288 ( .A(n11749), .ZN(n11750) );
  NAND2_X1 U14289 ( .A1(n11751), .A2(n11750), .ZN(n11752) );
  AND2_X1 U14290 ( .A1(n11753), .A2(n11752), .ZN(n13654) );
  NAND2_X1 U14291 ( .A1(n14153), .A2(n11778), .ZN(n11755) );
  NAND2_X1 U14292 ( .A1(n13755), .A2(n11777), .ZN(n11754) );
  NAND2_X1 U14293 ( .A1(n11755), .A2(n11754), .ZN(n11756) );
  XNOR2_X1 U14294 ( .A(n11756), .B(n11775), .ZN(n11760) );
  NAND2_X1 U14295 ( .A1(n14153), .A2(n11777), .ZN(n11758) );
  NAND2_X1 U14296 ( .A1(n13755), .A2(n6720), .ZN(n11757) );
  NAND2_X1 U14297 ( .A1(n11758), .A2(n11757), .ZN(n11759) );
  NOR2_X1 U14298 ( .A1(n11760), .A2(n11759), .ZN(n11761) );
  AOI21_X1 U14299 ( .B1(n11760), .B2(n11759), .A(n11761), .ZN(n13731) );
  INV_X1 U14300 ( .A(n11761), .ZN(n11762) );
  NAND2_X1 U14301 ( .A1(n13729), .A2(n11762), .ZN(n13603) );
  NAND2_X1 U14302 ( .A1(n13891), .A2(n11778), .ZN(n11764) );
  NAND2_X1 U14303 ( .A1(n13908), .A2(n11777), .ZN(n11763) );
  NAND2_X1 U14304 ( .A1(n11764), .A2(n11763), .ZN(n11765) );
  XNOR2_X1 U14305 ( .A(n11765), .B(n11775), .ZN(n11769) );
  NAND2_X1 U14306 ( .A1(n13891), .A2(n10439), .ZN(n11767) );
  NAND2_X1 U14307 ( .A1(n13908), .A2(n6720), .ZN(n11766) );
  NAND2_X1 U14308 ( .A1(n11767), .A2(n11766), .ZN(n11768) );
  NOR2_X1 U14309 ( .A1(n11769), .A2(n11768), .ZN(n11770) );
  AOI21_X1 U14310 ( .B1(n11769), .B2(n11768), .A(n11770), .ZN(n13604) );
  INV_X1 U14311 ( .A(n11770), .ZN(n11771) );
  NAND2_X1 U14312 ( .A1(n13602), .A2(n11771), .ZN(n11782) );
  NAND2_X1 U14313 ( .A1(n13584), .A2(n10677), .ZN(n11774) );
  OR2_X1 U14314 ( .A1(n12317), .A2(n11772), .ZN(n11773) );
  AOI22_X1 U14315 ( .A1(n14140), .A2(n10439), .B1(n6720), .B2(n13913), .ZN(
        n11776) );
  XNOR2_X1 U14316 ( .A(n11776), .B(n11775), .ZN(n11780) );
  AOI22_X1 U14317 ( .A1(n14140), .A2(n11778), .B1(n11777), .B2(n13913), .ZN(
        n11779) );
  XNOR2_X1 U14318 ( .A(n11780), .B(n11779), .ZN(n11781) );
  XNOR2_X1 U14319 ( .A(n11782), .B(n11781), .ZN(n11794) );
  NAND2_X1 U14320 ( .A1(n11783), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n11788) );
  NAND2_X1 U14321 ( .A1(n12320), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n11787) );
  INV_X1 U14322 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n15270) );
  OR2_X1 U14323 ( .A1(n11784), .A2(n15270), .ZN(n11786) );
  OR2_X1 U14324 ( .A1(n11600), .A2(n13900), .ZN(n11785) );
  NAND4_X1 U14325 ( .A1(n11788), .A2(n11787), .A3(n11786), .A4(n11785), .ZN(
        n13754) );
  NAND2_X1 U14326 ( .A1(n13754), .A2(n13732), .ZN(n11790) );
  NAND2_X1 U14327 ( .A1(n13908), .A2(n13897), .ZN(n11789) );
  NAND2_X1 U14328 ( .A1(n11790), .A2(n11789), .ZN(n14139) );
  AOI22_X1 U14329 ( .A1(n14537), .A2(n14139), .B1(P1_REG3_REG_28__SCAN_IN), 
        .B2(P1_U3086), .ZN(n11791) );
  OAI21_X1 U14330 ( .B1(n13923), .B2(n14542), .A(n11791), .ZN(n11792) );
  AOI21_X1 U14331 ( .B1(n14140), .B2(n14533), .A(n11792), .ZN(n11793) );
  OAI21_X1 U14332 ( .B1(n11794), .B2(n13727), .A(n11793), .ZN(P1_U3220) );
  INV_X1 U14333 ( .A(n11795), .ZN(n11797) );
  OAI222_X1 U14334 ( .A1(n13594), .A2(n11798), .B1(n13596), .B2(n11797), .C1(
        n11796), .C2(P2_U3088), .ZN(P2_U3305) );
  NAND2_X1 U14335 ( .A1(n12886), .A2(n15345), .ZN(n12080) );
  NAND2_X1 U14336 ( .A1(n11799), .A2(n11935), .ZN(n11801) );
  NAND2_X1 U14337 ( .A1(n12922), .A2(n12550), .ZN(n11800) );
  NAND2_X1 U14338 ( .A1(n11801), .A2(n11800), .ZN(n12861) );
  AND2_X1 U14339 ( .A1(n12918), .A2(n12851), .ZN(n11802) );
  OR2_X1 U14340 ( .A1(n12987), .A2(n12865), .ZN(n11959) );
  NAND2_X1 U14341 ( .A1(n12987), .A2(n12865), .ZN(n11956) );
  NAND2_X1 U14342 ( .A1(n12987), .A2(n12549), .ZN(n11803) );
  NAND2_X1 U14343 ( .A1(n12909), .A2(n11804), .ZN(n11957) );
  NAND2_X1 U14344 ( .A1(n11958), .A2(n11957), .ZN(n12839) );
  INV_X1 U14345 ( .A(n11804), .ZN(n12852) );
  OR2_X1 U14346 ( .A1(n12909), .A2(n12852), .ZN(n11805) );
  AND2_X1 U14347 ( .A1(n12979), .A2(n12838), .ZN(n11806) );
  NAND2_X1 U14348 ( .A1(n11807), .A2(n12826), .ZN(n12067) );
  INV_X1 U14349 ( .A(n12826), .ZN(n12453) );
  NAND2_X1 U14350 ( .A1(n12970), .A2(n12453), .ZN(n12066) );
  NAND2_X1 U14351 ( .A1(n12964), .A2(n12504), .ZN(n12071) );
  NAND2_X1 U14352 ( .A1(n12806), .A2(n12805), .ZN(n12793) );
  INV_X1 U14353 ( .A(n12504), .ZN(n12817) );
  OR2_X1 U14354 ( .A1(n12964), .A2(n12817), .ZN(n12794) );
  OR2_X1 U14355 ( .A1(n12958), .A2(n12807), .ZN(n11808) );
  AND2_X1 U14356 ( .A1(n12794), .A2(n11808), .ZN(n11809) );
  XNOR2_X1 U14357 ( .A(n12789), .B(n12797), .ZN(n12780) );
  NAND2_X1 U14358 ( .A1(n12789), .A2(n12797), .ZN(n11810) );
  NAND2_X1 U14359 ( .A1(n12491), .A2(n11811), .ZN(n11812) );
  NAND2_X1 U14360 ( .A1(n12886), .A2(n12773), .ZN(n11813) );
  NAND2_X1 U14361 ( .A1(n12758), .A2(n11813), .ZN(n12749) );
  OR2_X1 U14362 ( .A1(n12940), .A2(n12761), .ZN(n11814) );
  NAND2_X1 U14363 ( .A1(n12749), .A2(n11814), .ZN(n11816) );
  NAND2_X1 U14364 ( .A1(n12940), .A2(n12761), .ZN(n11815) );
  AOI22_X1 U14365 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(n11817), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(n15253), .ZN(n11818) );
  XNOR2_X1 U14366 ( .A(n11819), .B(n11818), .ZN(n13016) );
  NAND2_X1 U14367 ( .A1(n13016), .A2(n11913), .ZN(n11821) );
  OR2_X1 U14368 ( .A1(n9031), .A2(n13017), .ZN(n11820) );
  OR2_X1 U14369 ( .A1(n12118), .A2(n12750), .ZN(n11822) );
  AOI22_X1 U14370 ( .A1(P2_DATAO_REG_28__SCAN_IN), .A2(
        P1_DATAO_REG_28__SCAN_IN), .B1(n13587), .B2(n11772), .ZN(n11823) );
  XNOR2_X1 U14371 ( .A(n6517), .B(n11823), .ZN(n13013) );
  NAND2_X1 U14372 ( .A1(n13013), .A2(n11913), .ZN(n11826) );
  OR2_X1 U14373 ( .A1(n9031), .A2(n13015), .ZN(n11825) );
  NAND2_X1 U14374 ( .A1(n12932), .A2(n12736), .ZN(n11846) );
  INV_X1 U14375 ( .A(n12932), .ZN(n12728) );
  NAND2_X1 U14376 ( .A1(n12722), .A2(n7608), .ZN(n11836) );
  INV_X1 U14377 ( .A(n12712), .ZN(n11827) );
  NAND2_X1 U14378 ( .A1(n11827), .A2(n8697), .ZN(n11905) );
  INV_X1 U14379 ( .A(P3_REG0_REG_29__SCAN_IN), .ZN(n12925) );
  NAND2_X1 U14380 ( .A1(n11899), .A2(P3_REG2_REG_29__SCAN_IN), .ZN(n11829) );
  NAND2_X1 U14381 ( .A1(n6542), .A2(P3_REG1_REG_29__SCAN_IN), .ZN(n11828) );
  OAI211_X1 U14382 ( .C1(n12925), .C2(n6525), .A(n11829), .B(n11828), .ZN(
        n11830) );
  INV_X1 U14383 ( .A(n11830), .ZN(n11831) );
  NAND2_X1 U14384 ( .A1(n11905), .A2(n11831), .ZN(n12723) );
  OR2_X1 U14385 ( .A1(n9031), .A2(n11833), .ZN(n11834) );
  NAND2_X1 U14386 ( .A1(n12723), .A2(n12711), .ZN(n12097) );
  NAND2_X1 U14387 ( .A1(n11907), .A2(n12097), .ZN(n11856) );
  OR2_X1 U14388 ( .A1(n9116), .A2(n11837), .ZN(n11838) );
  NAND2_X1 U14389 ( .A1(n15052), .A2(n11838), .ZN(n14418) );
  INV_X1 U14390 ( .A(P3_REG0_REG_30__SCAN_IN), .ZN(n11841) );
  NAND2_X1 U14391 ( .A1(n6542), .A2(P3_REG1_REG_30__SCAN_IN), .ZN(n11840) );
  NAND2_X1 U14392 ( .A1(n8698), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n11839) );
  OAI211_X1 U14393 ( .C1(n11841), .C2(n6525), .A(n11840), .B(n11839), .ZN(
        n11842) );
  INV_X1 U14394 ( .A(n11842), .ZN(n11843) );
  NAND2_X1 U14395 ( .A1(n11905), .A2(n11843), .ZN(n12547) );
  INV_X1 U14396 ( .A(n12547), .ZN(n11844) );
  MUX2_X1 U14397 ( .A(n12709), .B(P3_REG1_REG_29__SCAN_IN), .S(n15129), .Z(
        n11858) );
  NAND2_X1 U14398 ( .A1(n12118), .A2(n11845), .ZN(n12715) );
  NAND2_X1 U14399 ( .A1(n11846), .A2(n12715), .ZN(n12090) );
  INV_X1 U14400 ( .A(n12772), .ZN(n11854) );
  NAND2_X1 U14401 ( .A1(n12958), .A2(n12414), .ZN(n11952) );
  XNOR2_X1 U14402 ( .A(n12918), .B(n12851), .ZN(n12860) );
  AND2_X1 U14403 ( .A1(n12918), .A2(n12470), .ZN(n12052) );
  INV_X1 U14404 ( .A(n12052), .ZN(n12056) );
  NAND2_X1 U14405 ( .A1(n12979), .A2(n12816), .ZN(n12061) );
  INV_X1 U14406 ( .A(n12061), .ZN(n11849) );
  OR2_X1 U14407 ( .A1(n12979), .A2(n12816), .ZN(n12062) );
  NAND2_X1 U14408 ( .A1(n12804), .A2(n12071), .ZN(n11850) );
  NAND2_X1 U14409 ( .A1(n11851), .A2(n11953), .ZN(n12779) );
  NAND2_X1 U14410 ( .A1(n12952), .A2(n12797), .ZN(n11945) );
  INV_X1 U14411 ( .A(n11945), .ZN(n11852) );
  INV_X1 U14412 ( .A(n11949), .ZN(n11853) );
  NAND2_X1 U14413 ( .A1(n12080), .A2(n12756), .ZN(n11855) );
  NAND2_X1 U14414 ( .A1(n12940), .A2(n12735), .ZN(n12085) );
  XOR2_X1 U14415 ( .A(n11856), .B(n11906), .Z(n12930) );
  OAI22_X1 U14416 ( .A1(n12930), .A2(n12924), .B1(n12711), .B2(n12907), .ZN(
        n11857) );
  INV_X1 U14417 ( .A(n13584), .ZN(n11859) );
  OAI222_X1 U14418 ( .A1(n9450), .A2(P1_U3086), .B1(n11860), .B2(n11859), .C1(
        n14247), .C2(n11772), .ZN(P1_U3327) );
  INV_X1 U14419 ( .A(n11861), .ZN(n11864) );
  INV_X1 U14420 ( .A(n11862), .ZN(n11863) );
  NAND2_X1 U14421 ( .A1(n11864), .A2(n11863), .ZN(n11865) );
  XNOR2_X1 U14422 ( .A(n13346), .B(n9271), .ZN(n11867) );
  NAND2_X1 U14423 ( .A1(n13356), .A2(n13269), .ZN(n13106) );
  INV_X1 U14424 ( .A(n11867), .ZN(n11868) );
  INV_X1 U14425 ( .A(n11870), .ZN(n11871) );
  AOI22_X1 U14426 ( .A1(n11871), .A2(n14462), .B1(n13105), .B2(n13143), .ZN(
        n11877) );
  NAND2_X1 U14427 ( .A1(n13295), .A2(n13402), .ZN(n11873) );
  NAND2_X1 U14428 ( .A1(n13356), .A2(n13401), .ZN(n11872) );
  NAND2_X1 U14429 ( .A1(n11873), .A2(n11872), .ZN(n13491) );
  AOI22_X1 U14430 ( .A1(n13491), .A2(n13131), .B1(P2_REG3_REG_23__SCAN_IN), 
        .B2(P2_U3088), .ZN(n11874) );
  OAI21_X1 U14431 ( .B1(n13328), .B2(n14467), .A(n11874), .ZN(n11875) );
  AOI21_X1 U14432 ( .B1(n13326), .B2(n14479), .A(n11875), .ZN(n11876) );
  OAI21_X1 U14433 ( .B1(n13025), .B2(n11877), .A(n11876), .ZN(P2_U3188) );
  INV_X1 U14434 ( .A(n11878), .ZN(n11888) );
  NAND3_X1 U14435 ( .A1(n13105), .A2(n11879), .A3(n13159), .ZN(n11880) );
  OAI21_X1 U14436 ( .B1(n14474), .B2(n13047), .A(n11880), .ZN(n11887) );
  OAI21_X1 U14437 ( .B1(n13110), .B2(n11882), .A(n11881), .ZN(n11886) );
  OAI22_X1 U14438 ( .A1(n14458), .A2(n11884), .B1(n11883), .B2(n14467), .ZN(
        n11885) );
  AOI211_X1 U14439 ( .C1(n11888), .C2(n11887), .A(n11886), .B(n11885), .ZN(
        n11889) );
  OAI21_X1 U14440 ( .B1(n11890), .B2(n14474), .A(n11889), .ZN(P2_U3202) );
  AND2_X1 U14441 ( .A1(n11891), .A2(P3_D_REG_31__SCAN_IN), .ZN(P3_U3234) );
  AND2_X1 U14442 ( .A1(n11891), .A2(P3_D_REG_30__SCAN_IN), .ZN(P3_U3235) );
  AND2_X1 U14443 ( .A1(n11891), .A2(P3_D_REG_28__SCAN_IN), .ZN(P3_U3237) );
  AND2_X1 U14444 ( .A1(n11891), .A2(P3_D_REG_23__SCAN_IN), .ZN(P3_U3242) );
  AND2_X1 U14445 ( .A1(n11891), .A2(P3_D_REG_20__SCAN_IN), .ZN(P3_U3245) );
  AND2_X1 U14446 ( .A1(n11891), .A2(P3_D_REG_15__SCAN_IN), .ZN(P3_U3250) );
  AND2_X1 U14447 ( .A1(n11891), .A2(P3_D_REG_11__SCAN_IN), .ZN(P3_U3254) );
  AND2_X1 U14448 ( .A1(n11891), .A2(P3_D_REG_9__SCAN_IN), .ZN(P3_U3256) );
  AND2_X1 U14449 ( .A1(n11891), .A2(P3_D_REG_7__SCAN_IN), .ZN(P3_U3258) );
  AND2_X1 U14450 ( .A1(n11891), .A2(P3_D_REG_4__SCAN_IN), .ZN(P3_U3261) );
  AND2_X1 U14451 ( .A1(n11891), .A2(P3_D_REG_25__SCAN_IN), .ZN(P3_U3240) );
  AND2_X1 U14452 ( .A1(n11891), .A2(P3_D_REG_17__SCAN_IN), .ZN(P3_U3248) );
  AND2_X1 U14453 ( .A1(n11891), .A2(P3_D_REG_3__SCAN_IN), .ZN(P3_U3262) );
  AND2_X1 U14454 ( .A1(n11891), .A2(P3_D_REG_5__SCAN_IN), .ZN(P3_U3260) );
  AND2_X1 U14455 ( .A1(n11891), .A2(P3_D_REG_6__SCAN_IN), .ZN(P3_U3259) );
  AND2_X1 U14456 ( .A1(n11891), .A2(P3_D_REG_8__SCAN_IN), .ZN(P3_U3257) );
  AND2_X1 U14457 ( .A1(n11891), .A2(P3_D_REG_13__SCAN_IN), .ZN(P3_U3252) );
  AND2_X1 U14458 ( .A1(n11891), .A2(P3_D_REG_16__SCAN_IN), .ZN(P3_U3249) );
  AND2_X1 U14459 ( .A1(n11891), .A2(P3_D_REG_18__SCAN_IN), .ZN(P3_U3247) );
  AND2_X1 U14460 ( .A1(n11891), .A2(P3_D_REG_22__SCAN_IN), .ZN(P3_U3243) );
  AND2_X1 U14461 ( .A1(n11891), .A2(P3_D_REG_24__SCAN_IN), .ZN(P3_U3241) );
  AND2_X1 U14462 ( .A1(n11891), .A2(P3_D_REG_27__SCAN_IN), .ZN(P3_U3238) );
  AND2_X1 U14463 ( .A1(n11891), .A2(P3_D_REG_29__SCAN_IN), .ZN(P3_U3236) );
  INV_X1 U14464 ( .A(n12097), .ZN(n11940) );
  NAND2_X1 U14465 ( .A1(P1_DATAO_REG_30__SCAN_IN), .A2(n12316), .ZN(n11909) );
  OAI21_X1 U14466 ( .B1(n12316), .B2(P1_DATAO_REG_30__SCAN_IN), .A(n11909), 
        .ZN(n11895) );
  OAI22_X1 U14467 ( .A1(P2_DATAO_REG_29__SCAN_IN), .A2(n13581), .B1(n11893), 
        .B2(n11892), .ZN(n11908) );
  INV_X1 U14468 ( .A(n11908), .ZN(n11894) );
  XNOR2_X1 U14469 ( .A(n11895), .B(n11894), .ZN(n13011) );
  OR2_X1 U14470 ( .A1(n9031), .A2(n13010), .ZN(n11897) );
  INV_X1 U14471 ( .A(P3_REG0_REG_31__SCAN_IN), .ZN(n11902) );
  NAND2_X1 U14472 ( .A1(n6542), .A2(P3_REG1_REG_31__SCAN_IN), .ZN(n11901) );
  NAND2_X1 U14473 ( .A1(n11899), .A2(P3_REG2_REG_31__SCAN_IN), .ZN(n11900) );
  OAI211_X1 U14474 ( .C1(n11902), .C2(n6525), .A(n11901), .B(n11900), .ZN(
        n11903) );
  INV_X1 U14475 ( .A(n11903), .ZN(n11904) );
  AND2_X1 U14476 ( .A1(n11905), .A2(n11904), .ZN(n14419) );
  INV_X1 U14477 ( .A(n14419), .ZN(n12546) );
  INV_X1 U14478 ( .A(n12096), .ZN(n11916) );
  OAI21_X1 U14479 ( .B1(P1_DATAO_REG_30__SCAN_IN), .B2(n12316), .A(n11908), 
        .ZN(n11910) );
  NAND2_X1 U14480 ( .A1(n11910), .A2(n11909), .ZN(n11912) );
  INV_X1 U14481 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n12137) );
  AOI22_X1 U14482 ( .A1(P2_DATAO_REG_31__SCAN_IN), .A2(n13577), .B1(
        P1_DATAO_REG_31__SCAN_IN), .B2(n12137), .ZN(n11911) );
  XOR2_X1 U14483 ( .A(n11912), .B(n11911), .Z(n13008) );
  NAND2_X1 U14484 ( .A1(n13008), .A2(n11913), .ZN(n11915) );
  INV_X1 U14485 ( .A(SI_31_), .ZN(n13004) );
  OR2_X1 U14486 ( .A1(n9031), .A2(n13004), .ZN(n11914) );
  INV_X1 U14487 ( .A(n14437), .ZN(n11919) );
  NAND2_X1 U14488 ( .A1(n11919), .A2(n12546), .ZN(n12099) );
  INV_X1 U14489 ( .A(n11943), .ZN(n11920) );
  NAND2_X1 U14490 ( .A1(n14437), .A2(n14419), .ZN(n11918) );
  NAND2_X1 U14491 ( .A1(n12547), .A2(n14422), .ZN(n11917) );
  NAND2_X1 U14492 ( .A1(n11918), .A2(n11917), .ZN(n12100) );
  INV_X1 U14493 ( .A(n12100), .ZN(n11942) );
  OAI22_X1 U14494 ( .A1(n11921), .A2(n11920), .B1(n11942), .B2(n11919), .ZN(
        n11922) );
  XNOR2_X1 U14495 ( .A(n11922), .B(n12691), .ZN(n12109) );
  NAND2_X1 U14496 ( .A1(n11953), .A2(n11952), .ZN(n12795) );
  NAND4_X1 U14497 ( .A1(n11965), .A2(n11925), .A3(n11924), .A4(n11923), .ZN(
        n11927) );
  NOR4_X1 U14498 ( .A1(n11927), .A2(n7134), .A3(n11926), .A4(n11990), .ZN(
        n11930) );
  NAND4_X1 U14499 ( .A1(n11930), .A2(n11929), .A3(n11928), .A4(n11975), .ZN(
        n11931) );
  NOR3_X1 U14500 ( .A1(n11931), .A2(n12028), .A3(n14432), .ZN(n11932) );
  NAND4_X1 U14501 ( .A1(n12045), .A2(n11933), .A3(n12040), .A4(n11932), .ZN(
        n11934) );
  NOR4_X1 U14502 ( .A1(n12839), .A2(n7138), .A3(n11935), .A4(n11934), .ZN(
        n11936) );
  XNOR2_X1 U14503 ( .A(n12979), .B(n12838), .ZN(n12825) );
  NAND4_X1 U14504 ( .A1(n12849), .A2(n12803), .A3(n11936), .A4(n12825), .ZN(
        n11937) );
  NOR4_X1 U14505 ( .A1(n12772), .A2(n12814), .A3(n12795), .A4(n11937), .ZN(
        n11938) );
  NAND4_X1 U14506 ( .A1(n12757), .A2(n12780), .A3(n12748), .A4(n11938), .ZN(
        n11939) );
  NOR3_X1 U14507 ( .A1(n12717), .A2(n11940), .A3(n11939), .ZN(n11941) );
  NAND4_X1 U14508 ( .A1(n11943), .A2(n11942), .A3(n11941), .A4(n12732), .ZN(
        n11944) );
  NAND2_X1 U14509 ( .A1(n11946), .A2(n11945), .ZN(n11947) );
  AND2_X1 U14510 ( .A1(n11947), .A2(n11949), .ZN(n11951) );
  INV_X1 U14511 ( .A(n12797), .ZN(n11948) );
  NAND2_X1 U14512 ( .A1(n12789), .A2(n11948), .ZN(n11950) );
  INV_X1 U14513 ( .A(n11952), .ZN(n11955) );
  INV_X1 U14514 ( .A(n11953), .ZN(n11954) );
  MUX2_X1 U14515 ( .A(n11955), .B(n11954), .S(n6529), .Z(n12079) );
  OAI211_X1 U14516 ( .C1(n12839), .C2(n11956), .A(n12062), .B(n11957), .ZN(
        n11962) );
  INV_X1 U14517 ( .A(n11957), .ZN(n11960) );
  OAI211_X1 U14518 ( .C1(n11960), .C2(n11959), .A(n12061), .B(n11958), .ZN(
        n11961) );
  MUX2_X1 U14519 ( .A(n11962), .B(n11961), .S(n6529), .Z(n12065) );
  OAI21_X1 U14520 ( .B1(n12918), .B2(n12470), .A(n11963), .ZN(n11964) );
  NAND2_X1 U14521 ( .A1(n11964), .A2(n12095), .ZN(n12054) );
  NAND3_X1 U14522 ( .A1(n11965), .A2(n12114), .A3(n11966), .ZN(n11972) );
  OAI21_X1 U14523 ( .B1(n11966), .B2(n12114), .A(n11968), .ZN(n11967) );
  NAND2_X1 U14524 ( .A1(n11967), .A2(n11973), .ZN(n11971) );
  NOR2_X1 U14525 ( .A1(n11969), .A2(n11968), .ZN(n11970) );
  AOI21_X1 U14526 ( .B1(n11972), .B2(n11971), .A(n11970), .ZN(n11981) );
  MUX2_X1 U14527 ( .A(n11974), .B(n11973), .S(n6529), .Z(n11976) );
  NAND2_X1 U14528 ( .A1(n11976), .A2(n11975), .ZN(n11980) );
  NAND2_X1 U14529 ( .A1(n11987), .A2(n11977), .ZN(n11978) );
  NAND2_X1 U14530 ( .A1(n11978), .A2(n12095), .ZN(n11979) );
  OAI21_X1 U14531 ( .B1(n11981), .B2(n11980), .A(n11979), .ZN(n11986) );
  NAND2_X1 U14532 ( .A1(n12557), .A2(n11982), .ZN(n11983) );
  AOI21_X1 U14533 ( .B1(n11985), .B2(n11983), .A(n12095), .ZN(n11984) );
  AOI21_X1 U14534 ( .B1(n11986), .B2(n11985), .A(n11984), .ZN(n11994) );
  OAI21_X1 U14535 ( .B1(n12095), .B2(n11987), .A(n15059), .ZN(n11993) );
  MUX2_X1 U14536 ( .A(n11989), .B(n11988), .S(n12095), .Z(n11991) );
  NOR2_X1 U14537 ( .A1(n11991), .A2(n11990), .ZN(n11992) );
  OAI21_X1 U14538 ( .B1(n11994), .B2(n11993), .A(n11992), .ZN(n11998) );
  NAND2_X1 U14539 ( .A1(n12004), .A2(n11995), .ZN(n11996) );
  NAND2_X1 U14540 ( .A1(n11996), .A2(n12095), .ZN(n11997) );
  NAND2_X1 U14541 ( .A1(n11998), .A2(n11997), .ZN(n12002) );
  AOI21_X1 U14542 ( .B1(n12001), .B2(n11999), .A(n12095), .ZN(n12000) );
  AOI21_X1 U14543 ( .B1(n12002), .B2(n12001), .A(n12000), .ZN(n12011) );
  OAI21_X1 U14544 ( .B1(n12095), .B2(n12004), .A(n12003), .ZN(n12010) );
  MUX2_X1 U14545 ( .A(n12006), .B(n12005), .S(n6529), .Z(n12008) );
  NOR2_X1 U14546 ( .A1(n12008), .A2(n12007), .ZN(n12009) );
  OAI21_X1 U14547 ( .B1(n12011), .B2(n12010), .A(n12009), .ZN(n12023) );
  INV_X1 U14548 ( .A(n12012), .ZN(n12015) );
  INV_X1 U14549 ( .A(n12013), .ZN(n12014) );
  MUX2_X1 U14550 ( .A(n12015), .B(n12014), .S(n12095), .Z(n12017) );
  NOR2_X1 U14551 ( .A1(n12017), .A2(n12016), .ZN(n12022) );
  INV_X1 U14552 ( .A(n12018), .ZN(n12020) );
  MUX2_X1 U14553 ( .A(n12020), .B(n12019), .S(n6529), .Z(n12021) );
  AOI21_X1 U14554 ( .B1(n12023), .B2(n12022), .A(n12021), .ZN(n12029) );
  MUX2_X1 U14555 ( .A(n12025), .B(n12024), .S(n6529), .Z(n12026) );
  NOR2_X1 U14556 ( .A1(n14432), .A2(n12026), .ZN(n12027) );
  OAI21_X1 U14557 ( .B1(n12029), .B2(n12028), .A(n12027), .ZN(n12034) );
  NAND2_X1 U14558 ( .A1(n12037), .A2(n12030), .ZN(n12031) );
  NAND2_X1 U14559 ( .A1(n12031), .A2(n12095), .ZN(n12033) );
  AOI21_X1 U14560 ( .B1(n12034), .B2(n12033), .A(n12032), .ZN(n12039) );
  AOI21_X1 U14561 ( .B1(n12036), .B2(n12035), .A(n12095), .ZN(n12038) );
  OAI22_X1 U14562 ( .A1(n12039), .A2(n12038), .B1(n12095), .B2(n12037), .ZN(
        n12041) );
  NAND2_X1 U14563 ( .A1(n12041), .A2(n12040), .ZN(n12046) );
  MUX2_X1 U14564 ( .A(n12043), .B(n12042), .S(n12095), .Z(n12044) );
  NAND3_X1 U14565 ( .A1(n12046), .A2(n12045), .A3(n12044), .ZN(n12051) );
  MUX2_X1 U14566 ( .A(n12048), .B(n12047), .S(n12095), .Z(n12049) );
  NAND3_X1 U14567 ( .A1(n12051), .A2(n12050), .A3(n12049), .ZN(n12053) );
  AOI21_X1 U14568 ( .B1(n12054), .B2(n12053), .A(n12052), .ZN(n12059) );
  AOI21_X1 U14569 ( .B1(n12056), .B2(n12055), .A(n12095), .ZN(n12058) );
  NAND2_X1 U14570 ( .A1(n12851), .A2(n6529), .ZN(n12057) );
  OAI22_X1 U14571 ( .A1(n12059), .A2(n12058), .B1(n12918), .B2(n12057), .ZN(
        n12060) );
  AND3_X1 U14572 ( .A1(n6716), .A2(n12849), .A3(n12060), .ZN(n12064) );
  MUX2_X1 U14573 ( .A(n12062), .B(n12061), .S(n12095), .Z(n12063) );
  OAI21_X1 U14574 ( .B1(n12065), .B2(n12064), .A(n12063), .ZN(n12069) );
  MUX2_X1 U14575 ( .A(n12067), .B(n12066), .S(n12095), .Z(n12068) );
  OAI211_X1 U14576 ( .C1(n12814), .C2(n12069), .A(n12068), .B(n12803), .ZN(
        n12076) );
  INV_X1 U14577 ( .A(n12070), .ZN(n12073) );
  INV_X1 U14578 ( .A(n12071), .ZN(n12072) );
  MUX2_X1 U14579 ( .A(n12073), .B(n12072), .S(n6529), .Z(n12074) );
  INV_X1 U14580 ( .A(n12074), .ZN(n12075) );
  NAND2_X1 U14581 ( .A1(n12076), .A2(n12075), .ZN(n12077) );
  OAI21_X1 U14582 ( .B1(n12795), .B2(n12077), .A(n12780), .ZN(n12078) );
  NAND3_X1 U14583 ( .A1(n12748), .A2(n12080), .A3(n12083), .ZN(n12082) );
  NAND3_X1 U14584 ( .A1(n12748), .A2(n12084), .A3(n12083), .ZN(n12086) );
  NAND2_X1 U14585 ( .A1(n12937), .A2(n12750), .ZN(n12088) );
  INV_X1 U14586 ( .A(n12089), .ZN(n12092) );
  NOR2_X1 U14587 ( .A1(n12090), .A2(n12095), .ZN(n12091) );
  OAI33_X1 U14588 ( .A1(n12095), .A2(n12094), .A3(n12717), .B1(n12093), .B2(
        n12092), .B3(n12091), .ZN(n12098) );
  AOI21_X1 U14589 ( .B1(n12098), .B2(n12097), .A(n12096), .ZN(n12101) );
  OAI21_X1 U14590 ( .B1(n12101), .B2(n12100), .A(n12099), .ZN(n12102) );
  MUX2_X1 U14591 ( .A(n12104), .B(n12103), .S(n12102), .Z(n12105) );
  OAI21_X1 U14592 ( .B1(n12107), .B2(n12106), .A(n12105), .ZN(n12108) );
  AOI21_X1 U14593 ( .B1(n12110), .B2(n12109), .A(n12108), .ZN(n12117) );
  NAND3_X1 U14594 ( .A1(n12112), .A2(n12111), .A3(n12670), .ZN(n12113) );
  OAI211_X1 U14595 ( .C1(n12114), .C2(n12116), .A(n12113), .B(P3_B_REG_SCAN_IN), .ZN(n12115) );
  OAI21_X1 U14596 ( .B1(n12117), .B2(n12116), .A(n12115), .ZN(P3_U3296) );
  XNOR2_X1 U14597 ( .A(n12118), .B(n8709), .ZN(n12119) );
  NOR2_X1 U14598 ( .A1(n12119), .A2(n12750), .ZN(n12127) );
  AOI21_X1 U14599 ( .B1(n12750), .B2(n12119), .A(n12127), .ZN(n12392) );
  AND2_X1 U14600 ( .A1(n12120), .A2(n12392), .ZN(n12125) );
  INV_X1 U14601 ( .A(n12392), .ZN(n12124) );
  INV_X1 U14602 ( .A(n12121), .ZN(n12122) );
  INV_X1 U14603 ( .A(n12127), .ZN(n12128) );
  NAND2_X1 U14604 ( .A1(n12390), .A2(n12128), .ZN(n12130) );
  XNOR2_X1 U14605 ( .A(n12720), .B(n8709), .ZN(n12129) );
  XNOR2_X1 U14606 ( .A(n12130), .B(n12129), .ZN(n12136) );
  INV_X1 U14607 ( .A(n12723), .ZN(n12133) );
  AOI22_X1 U14608 ( .A1(n12750), .A2(n12525), .B1(P3_REG3_REG_28__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12132) );
  NAND2_X1 U14609 ( .A1(n12726), .A2(n12540), .ZN(n12131) );
  OAI211_X1 U14610 ( .C1(n12133), .C2(n12484), .A(n12132), .B(n12131), .ZN(
        n12134) );
  AOI21_X1 U14611 ( .B1(n12932), .B2(n12524), .A(n12134), .ZN(n12135) );
  OAI21_X1 U14612 ( .B1(n12136), .B2(n12507), .A(n12135), .ZN(P3_U3160) );
  NAND2_X1 U14613 ( .A1(n13575), .A2(n10677), .ZN(n12139) );
  OR2_X1 U14614 ( .A1(n12317), .A2(n12137), .ZN(n12138) );
  NAND2_X1 U14615 ( .A1(n12144), .A2(n13868), .ZN(n12140) );
  NOR2_X1 U14616 ( .A1(n13880), .A2(n12330), .ZN(n12370) );
  NAND2_X1 U14617 ( .A1(n12144), .A2(n12143), .ZN(n12145) );
  NAND2_X1 U14618 ( .A1(n12146), .A2(n12145), .ZN(n12148) );
  NAND2_X1 U14619 ( .A1(n12148), .A2(n12147), .ZN(n12377) );
  NAND2_X1 U14620 ( .A1(n12377), .A2(n12375), .ZN(n12366) );
  NAND2_X1 U14621 ( .A1(n13880), .A2(n12330), .ZN(n12368) );
  NOR2_X1 U14622 ( .A1(n12368), .A2(n12371), .ZN(n12149) );
  AOI211_X1 U14623 ( .C1(n12370), .C2(n12371), .A(n12366), .B(n12149), .ZN(
        n12150) );
  OR2_X1 U14624 ( .A1(n12167), .A2(n12179), .ZN(n12157) );
  NAND3_X1 U14625 ( .A1(n12151), .A2(n12179), .A3(n12167), .ZN(n12156) );
  INV_X1 U14626 ( .A(n12166), .ZN(n12152) );
  NAND2_X1 U14627 ( .A1(n12152), .A2(n12179), .ZN(n12155) );
  NAND3_X1 U14628 ( .A1(n12153), .A2(n12166), .A3(n12173), .ZN(n12154) );
  NAND4_X1 U14629 ( .A1(n12157), .A2(n12156), .A3(n12155), .A4(n12154), .ZN(
        n12158) );
  NOR2_X1 U14630 ( .A1(n12158), .A2(n14654), .ZN(n12178) );
  NAND2_X1 U14631 ( .A1(n12339), .A2(n12159), .ZN(n12160) );
  NAND2_X1 U14632 ( .A1(n13780), .A2(n14677), .ZN(n12338) );
  NAND2_X1 U14633 ( .A1(n12160), .A2(n12338), .ZN(n12162) );
  INV_X1 U14634 ( .A(n12339), .ZN(n12161) );
  NAND2_X1 U14635 ( .A1(n6770), .A2(n12163), .ZN(n12164) );
  NAND2_X1 U14636 ( .A1(n12165), .A2(n12164), .ZN(n12168) );
  INV_X1 U14637 ( .A(n12171), .ZN(n12175) );
  INV_X1 U14638 ( .A(n12172), .ZN(n12174) );
  MUX2_X1 U14639 ( .A(n12175), .B(n12174), .S(n12173), .Z(n12176) );
  MUX2_X1 U14640 ( .A(n13775), .B(n14720), .S(n12179), .Z(n12181) );
  NAND2_X1 U14641 ( .A1(n12180), .A2(n12181), .ZN(n12185) );
  MUX2_X1 U14642 ( .A(n14720), .B(n13775), .S(n12179), .Z(n12184) );
  INV_X1 U14643 ( .A(n12180), .ZN(n12183) );
  INV_X1 U14644 ( .A(n12181), .ZN(n12182) );
  MUX2_X1 U14645 ( .A(n12187), .B(n12186), .S(n12179), .Z(n12190) );
  MUX2_X1 U14646 ( .A(n12188), .B(n14649), .S(n12179), .Z(n12189) );
  NAND2_X1 U14647 ( .A1(n12191), .A2(n12190), .ZN(n12192) );
  NAND2_X1 U14648 ( .A1(n12193), .A2(n12192), .ZN(n12198) );
  MUX2_X1 U14649 ( .A(n13774), .B(n12194), .S(n12179), .Z(n12197) );
  NAND2_X1 U14650 ( .A1(n12198), .A2(n12197), .ZN(n12196) );
  MUX2_X1 U14651 ( .A(n12194), .B(n13774), .S(n12330), .Z(n12195) );
  NAND2_X1 U14652 ( .A1(n12196), .A2(n12195), .ZN(n12200) );
  NAND2_X1 U14653 ( .A1(n12200), .A2(n12199), .ZN(n12202) );
  MUX2_X1 U14654 ( .A(n13773), .B(n14743), .S(n12328), .Z(n12203) );
  MUX2_X1 U14655 ( .A(n13773), .B(n14743), .S(n12330), .Z(n12201) );
  INV_X1 U14656 ( .A(n12203), .ZN(n12204) );
  MUX2_X1 U14657 ( .A(n13772), .B(n12205), .S(n12330), .Z(n12209) );
  MUX2_X1 U14658 ( .A(n13772), .B(n12205), .S(n12328), .Z(n12206) );
  NAND2_X1 U14659 ( .A1(n12207), .A2(n12206), .ZN(n12213) );
  INV_X1 U14660 ( .A(n12208), .ZN(n12211) );
  INV_X1 U14661 ( .A(n12209), .ZN(n12210) );
  NAND2_X1 U14662 ( .A1(n12211), .A2(n12210), .ZN(n12212) );
  MUX2_X1 U14663 ( .A(n13771), .B(n12214), .S(n12328), .Z(n12216) );
  MUX2_X1 U14664 ( .A(n13771), .B(n12214), .S(n12330), .Z(n12215) );
  MUX2_X1 U14665 ( .A(n13770), .B(n12217), .S(n12330), .Z(n12221) );
  MUX2_X1 U14666 ( .A(n13770), .B(n12217), .S(n12328), .Z(n12218) );
  NAND2_X1 U14667 ( .A1(n12219), .A2(n12218), .ZN(n12232) );
  INV_X1 U14668 ( .A(n12220), .ZN(n12223) );
  INV_X1 U14669 ( .A(n12221), .ZN(n12222) );
  NAND2_X1 U14670 ( .A1(n12223), .A2(n12222), .ZN(n12229) );
  NAND2_X1 U14671 ( .A1(n12232), .A2(n12229), .ZN(n12224) );
  MUX2_X1 U14672 ( .A(n13769), .B(n12225), .S(n12328), .Z(n12228) );
  NAND2_X1 U14673 ( .A1(n12224), .A2(n12228), .ZN(n12227) );
  MUX2_X1 U14674 ( .A(n13769), .B(n12225), .S(n12330), .Z(n12226) );
  NAND2_X1 U14675 ( .A1(n12227), .A2(n12226), .ZN(n12234) );
  INV_X1 U14676 ( .A(n12228), .ZN(n12230) );
  AND2_X1 U14677 ( .A1(n12230), .A2(n12229), .ZN(n12231) );
  NAND2_X1 U14678 ( .A1(n12232), .A2(n12231), .ZN(n12233) );
  NAND2_X1 U14679 ( .A1(n12234), .A2(n12233), .ZN(n12238) );
  MUX2_X1 U14680 ( .A(n13768), .B(n12235), .S(n12330), .Z(n12239) );
  NAND2_X1 U14681 ( .A1(n12238), .A2(n12239), .ZN(n12237) );
  MUX2_X1 U14682 ( .A(n13768), .B(n12235), .S(n12328), .Z(n12236) );
  NAND2_X1 U14683 ( .A1(n12237), .A2(n12236), .ZN(n12243) );
  INV_X1 U14684 ( .A(n12238), .ZN(n12241) );
  INV_X1 U14685 ( .A(n12239), .ZN(n12240) );
  NAND2_X1 U14686 ( .A1(n12241), .A2(n12240), .ZN(n12242) );
  MUX2_X1 U14687 ( .A(n13767), .B(n13706), .S(n12328), .Z(n12245) );
  MUX2_X1 U14688 ( .A(n13767), .B(n13706), .S(n12330), .Z(n12244) );
  INV_X1 U14689 ( .A(n14534), .ZN(n14550) );
  OAI21_X1 U14690 ( .B1(n14550), .B2(n13766), .A(n14082), .ZN(n12249) );
  NAND2_X1 U14691 ( .A1(n12252), .A2(n14096), .ZN(n12248) );
  MUX2_X1 U14692 ( .A(n12249), .B(n12248), .S(n12328), .Z(n12250) );
  INV_X1 U14693 ( .A(n12250), .ZN(n12255) );
  MUX2_X1 U14694 ( .A(n13746), .B(n14215), .S(n12328), .Z(n12257) );
  MUX2_X1 U14695 ( .A(n13765), .B(n12251), .S(n12330), .Z(n12256) );
  MUX2_X1 U14696 ( .A(n13764), .B(n14209), .S(n12330), .Z(n12259) );
  OR2_X1 U14697 ( .A1(n12259), .A2(n12335), .ZN(n12258) );
  MUX2_X1 U14698 ( .A(n14082), .B(n12252), .S(n12330), .Z(n12253) );
  OAI211_X1 U14699 ( .C1(n12257), .C2(n12256), .A(n12258), .B(n12253), .ZN(
        n12254) );
  NAND3_X1 U14700 ( .A1(n12258), .A2(n12257), .A3(n12256), .ZN(n12261) );
  NAND2_X1 U14701 ( .A1(n12259), .A2(n12336), .ZN(n12260) );
  AND2_X1 U14702 ( .A1(n12330), .A2(n13763), .ZN(n12263) );
  NOR2_X1 U14703 ( .A1(n12330), .A2(n13763), .ZN(n12262) );
  MUX2_X1 U14704 ( .A(n12263), .B(n12262), .S(n14204), .Z(n12264) );
  NOR2_X1 U14705 ( .A1(n14048), .A2(n12264), .ZN(n12265) );
  MUX2_X1 U14706 ( .A(n14019), .B(n12266), .S(n12328), .Z(n12267) );
  NAND2_X1 U14707 ( .A1(n12268), .A2(n12267), .ZN(n12271) );
  MUX2_X1 U14708 ( .A(n13627), .B(n14192), .S(n12328), .Z(n12270) );
  MUX2_X1 U14709 ( .A(n13761), .B(n14029), .S(n12330), .Z(n12269) );
  NAND2_X1 U14710 ( .A1(n12271), .A2(n12270), .ZN(n12272) );
  MUX2_X1 U14711 ( .A(n13760), .B(n14013), .S(n12330), .Z(n12275) );
  MUX2_X1 U14712 ( .A(n13760), .B(n14013), .S(n12328), .Z(n12274) );
  INV_X1 U14713 ( .A(n12280), .ZN(n12278) );
  MUX2_X1 U14714 ( .A(n13759), .B(n12276), .S(n12328), .Z(n12279) );
  INV_X1 U14715 ( .A(n12279), .ZN(n12277) );
  NAND2_X1 U14716 ( .A1(n12280), .A2(n12279), .ZN(n12282) );
  MUX2_X1 U14717 ( .A(n13759), .B(n12276), .S(n12330), .Z(n12281) );
  NAND2_X1 U14718 ( .A1(n12282), .A2(n12281), .ZN(n12283) );
  MUX2_X1 U14719 ( .A(n13758), .B(n13981), .S(n12330), .Z(n12285) );
  MUX2_X1 U14720 ( .A(n13758), .B(n13981), .S(n12328), .Z(n12284) );
  MUX2_X1 U14721 ( .A(n13757), .B(n14165), .S(n12328), .Z(n12289) );
  NAND2_X1 U14722 ( .A1(n12288), .A2(n12289), .ZN(n12287) );
  MUX2_X1 U14723 ( .A(n13757), .B(n14165), .S(n12330), .Z(n12286) );
  NAND2_X1 U14724 ( .A1(n12287), .A2(n12286), .ZN(n12296) );
  INV_X1 U14725 ( .A(n12288), .ZN(n12291) );
  INV_X1 U14726 ( .A(n12289), .ZN(n12290) );
  NAND2_X1 U14727 ( .A1(n12291), .A2(n12290), .ZN(n12295) );
  MUX2_X1 U14728 ( .A(n13756), .B(n14159), .S(n12330), .Z(n12293) );
  MUX2_X1 U14729 ( .A(n13756), .B(n14159), .S(n12328), .Z(n12292) );
  INV_X1 U14730 ( .A(n12293), .ZN(n12294) );
  MUX2_X1 U14731 ( .A(n13755), .B(n14153), .S(n12328), .Z(n12300) );
  NAND2_X1 U14732 ( .A1(n12299), .A2(n12300), .ZN(n12298) );
  MUX2_X1 U14733 ( .A(n13755), .B(n14153), .S(n12330), .Z(n12297) );
  NAND2_X1 U14734 ( .A1(n12298), .A2(n12297), .ZN(n12304) );
  INV_X1 U14735 ( .A(n12299), .ZN(n12302) );
  INV_X1 U14736 ( .A(n12300), .ZN(n12301) );
  NAND2_X1 U14737 ( .A1(n12302), .A2(n12301), .ZN(n12303) );
  MUX2_X1 U14738 ( .A(n13908), .B(n13891), .S(n12330), .Z(n12306) );
  MUX2_X1 U14739 ( .A(n13908), .B(n13891), .S(n12328), .Z(n12305) );
  MUX2_X1 U14740 ( .A(n13913), .B(n14140), .S(n12328), .Z(n12308) );
  MUX2_X1 U14741 ( .A(n13913), .B(n14140), .S(n12330), .Z(n12307) );
  INV_X1 U14742 ( .A(n12308), .ZN(n12309) );
  NAND2_X1 U14743 ( .A1(n12385), .A2(n10677), .ZN(n12311) );
  OR2_X1 U14744 ( .A1(n12317), .A2(n12386), .ZN(n12310) );
  MUX2_X1 U14745 ( .A(n13754), .B(n13896), .S(n12330), .Z(n12312) );
  MUX2_X1 U14746 ( .A(n13754), .B(n13896), .S(n12328), .Z(n12314) );
  INV_X1 U14747 ( .A(n12312), .ZN(n12313) );
  NAND2_X1 U14748 ( .A1(n12315), .A2(n10677), .ZN(n12319) );
  OR2_X1 U14749 ( .A1(n12317), .A2(n12316), .ZN(n12318) );
  INV_X1 U14750 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n12324) );
  NAND2_X1 U14751 ( .A1(n12320), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n12323) );
  NAND2_X1 U14752 ( .A1(n12321), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n12322) );
  OAI211_X1 U14753 ( .C1(n6539), .C2(n12324), .A(n12323), .B(n12322), .ZN(
        n13899) );
  OAI22_X1 U14754 ( .A1(n12328), .A2(n13877), .B1(n9357), .B2(n12326), .ZN(
        n12327) );
  AOI22_X1 U14755 ( .A1(n13887), .A2(n12328), .B1(n13899), .B2(n12327), .ZN(
        n12332) );
  OAI21_X1 U14756 ( .B1(n12371), .B2(n12329), .A(n13899), .ZN(n12331) );
  MUX2_X1 U14757 ( .A(n12331), .B(n14130), .S(n12330), .Z(n12334) );
  XNOR2_X1 U14758 ( .A(n14130), .B(n13899), .ZN(n12364) );
  XNOR2_X1 U14759 ( .A(n13896), .B(n13754), .ZN(n13914) );
  INV_X1 U14760 ( .A(n12335), .ZN(n12337) );
  NAND2_X1 U14761 ( .A1(n12337), .A2(n12336), .ZN(n14075) );
  NAND2_X1 U14762 ( .A1(n12339), .A2(n12338), .ZN(n14688) );
  NOR4_X1 U14763 ( .A1(n6726), .A2(n14654), .A3(n12340), .A4(n14688), .ZN(
        n12345) );
  NAND4_X1 U14764 ( .A1(n12345), .A2(n12344), .A3(n12343), .A4(n12342), .ZN(
        n12349) );
  NOR4_X1 U14765 ( .A1(n12349), .A2(n12348), .A3(n12347), .A4(n12346), .ZN(
        n12351) );
  NAND4_X1 U14766 ( .A1(n12353), .A2(n12352), .A3(n12351), .A4(n12350), .ZN(
        n12354) );
  NOR4_X1 U14767 ( .A1(n14105), .A2(n6699), .A3(n12355), .A4(n12354), .ZN(
        n12356) );
  NAND3_X1 U14768 ( .A1(n14075), .A2(n12356), .A3(n14085), .ZN(n12357) );
  NOR4_X1 U14769 ( .A1(n12358), .A2(n14053), .A3(n14048), .A4(n12357), .ZN(
        n12359) );
  NAND4_X1 U14770 ( .A1(n13988), .A2(n13976), .A3(n12359), .A4(n14006), .ZN(
        n12360) );
  NOR4_X1 U14771 ( .A1(n13932), .A2(n13952), .A3(n13957), .A4(n12360), .ZN(
        n12362) );
  NAND4_X1 U14772 ( .A1(n13914), .A2(n12362), .A3(n13921), .A4(n12361), .ZN(
        n12363) );
  NOR3_X1 U14773 ( .A1(n12378), .A2(n12364), .A3(n12363), .ZN(n12365) );
  XOR2_X1 U14774 ( .A(n13868), .B(n12365), .Z(n12376) );
  NOR3_X1 U14775 ( .A1(n14122), .A2(n12371), .A3(n12366), .ZN(n12369) );
  NOR3_X1 U14776 ( .A1(n12368), .A2(n12371), .A3(n12377), .ZN(n12367) );
  AOI21_X1 U14777 ( .B1(n12369), .B2(n12368), .A(n12367), .ZN(n12374) );
  XOR2_X1 U14778 ( .A(n12377), .B(n12370), .Z(n12372) );
  NAND4_X1 U14779 ( .A1(n12372), .A2(n14122), .A3(n12371), .A4(n12375), .ZN(
        n12373) );
  NAND3_X1 U14780 ( .A1(n12381), .A2(n14601), .A3(n13897), .ZN(n12382) );
  OAI211_X1 U14781 ( .C1(n6796), .C2(n12384), .A(n12382), .B(P1_B_REG_SCAN_IN), 
        .ZN(n12383) );
  INV_X1 U14782 ( .A(n12385), .ZN(n13582) );
  OAI222_X1 U14783 ( .A1(n11860), .A2(n13582), .B1(n12387), .B2(P1_U3086), 
        .C1(n12386), .C2(n14247), .ZN(P1_U3326) );
  NAND2_X1 U14784 ( .A1(n12389), .A2(n12388), .ZN(n12391) );
  OAI21_X1 U14785 ( .B1(n12392), .B2(n12391), .A(n12390), .ZN(n12393) );
  NAND2_X1 U14786 ( .A1(n12393), .A2(n12533), .ZN(n12397) );
  AOI22_X1 U14787 ( .A1(n12761), .A2(n12525), .B1(P3_REG3_REG_27__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12394) );
  OAI21_X1 U14788 ( .B1(n12736), .B2(n12484), .A(n12394), .ZN(n12395) );
  AOI21_X1 U14789 ( .B1(n12741), .B2(n12540), .A(n12395), .ZN(n12396) );
  OAI211_X1 U14790 ( .C1(n12937), .C2(n12544), .A(n12397), .B(n12396), .ZN(
        P3_U3154) );
  INV_X1 U14791 ( .A(n12398), .ZN(n12399) );
  AOI21_X1 U14792 ( .B1(n12401), .B2(n12400), .A(n12399), .ZN(n12410) );
  NAND2_X1 U14793 ( .A1(n12540), .A2(n12402), .ZN(n12405) );
  NOR2_X1 U14794 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n12403), .ZN(n12597) );
  AOI21_X1 U14795 ( .B1(n12535), .B2(n12550), .A(n12597), .ZN(n12404) );
  OAI211_X1 U14796 ( .C1(n12406), .C2(n12537), .A(n12405), .B(n12404), .ZN(
        n12407) );
  AOI21_X1 U14797 ( .B1(n12408), .B2(n12524), .A(n12407), .ZN(n12409) );
  OAI21_X1 U14798 ( .B1(n12410), .B2(n12507), .A(n12409), .ZN(P3_U3155) );
  AOI21_X1 U14799 ( .B1(n12797), .B2(n12411), .A(n6546), .ZN(n12417) );
  NAND2_X1 U14800 ( .A1(n12540), .A2(n12788), .ZN(n12413) );
  AOI22_X1 U14801 ( .A1(n12784), .A2(n12535), .B1(P3_REG3_REG_23__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12412) );
  OAI211_X1 U14802 ( .C1(n12414), .C2(n12537), .A(n12413), .B(n12412), .ZN(
        n12415) );
  AOI21_X1 U14803 ( .B1(n12789), .B2(n12524), .A(n12415), .ZN(n12416) );
  OAI21_X1 U14804 ( .B1(n12417), .B2(n12507), .A(n12416), .ZN(P3_U3156) );
  AOI21_X1 U14805 ( .B1(n12419), .B2(n12418), .A(n12507), .ZN(n12421) );
  NAND2_X1 U14806 ( .A1(n12421), .A2(n12420), .ZN(n12428) );
  NAND2_X1 U14807 ( .A1(P3_REG3_REG_10__SCAN_IN), .A2(P3_U3151), .ZN(n15027)
         );
  INV_X1 U14808 ( .A(n15027), .ZN(n12422) );
  AOI21_X1 U14809 ( .B1(n12524), .B2(n12423), .A(n12422), .ZN(n12427) );
  AOI22_X1 U14810 ( .A1(n12535), .A2(n12553), .B1(n12525), .B2(n12554), .ZN(
        n12426) );
  NAND2_X1 U14811 ( .A1(n12540), .A2(n12424), .ZN(n12425) );
  NAND4_X1 U14812 ( .A1(n12428), .A2(n12427), .A3(n12426), .A4(n12425), .ZN(
        P3_U3157) );
  AOI211_X1 U14813 ( .C1(n12431), .C2(n12430), .A(n12507), .B(n12429), .ZN(
        n12432) );
  INV_X1 U14814 ( .A(n12432), .ZN(n12438) );
  NOR2_X1 U14815 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n12434), .ZN(n14953) );
  AOI21_X1 U14816 ( .B1(n12524), .B2(n12433), .A(n14953), .ZN(n12437) );
  AOI22_X1 U14817 ( .A1(n12535), .A2(n15037), .B1(n12525), .B2(n12557), .ZN(
        n12436) );
  NAND2_X1 U14818 ( .A1(n12540), .A2(n12434), .ZN(n12435) );
  NAND4_X1 U14819 ( .A1(n12438), .A2(n12437), .A3(n12436), .A4(n12435), .ZN(
        P3_U3158) );
  AOI21_X1 U14820 ( .B1(n12440), .B2(n12439), .A(n12507), .ZN(n12442) );
  NAND2_X1 U14821 ( .A1(n12442), .A2(n12441), .ZN(n12446) );
  NAND2_X1 U14822 ( .A1(n12525), .A2(n12852), .ZN(n12443) );
  NAND2_X1 U14823 ( .A1(P3_U3151), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n12699)
         );
  OAI211_X1 U14824 ( .C1(n12453), .C2(n12484), .A(n12443), .B(n12699), .ZN(
        n12444) );
  AOI21_X1 U14825 ( .B1(n12540), .B2(n12829), .A(n12444), .ZN(n12445) );
  OAI211_X1 U14826 ( .C1(n12544), .C2(n12979), .A(n12446), .B(n12445), .ZN(
        P3_U3159) );
  INV_X1 U14827 ( .A(n12447), .ZN(n12448) );
  AOI21_X1 U14828 ( .B1(n12450), .B2(n12449), .A(n12448), .ZN(n12456) );
  NAND2_X1 U14829 ( .A1(n12540), .A2(n12810), .ZN(n12452) );
  AOI22_X1 U14830 ( .A1(n12807), .A2(n12535), .B1(P3_REG3_REG_21__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12451) );
  OAI211_X1 U14831 ( .C1(n12453), .C2(n12537), .A(n12452), .B(n12451), .ZN(
        n12454) );
  AOI21_X1 U14832 ( .B1(n12964), .B2(n12524), .A(n12454), .ZN(n12455) );
  OAI21_X1 U14833 ( .B1(n12456), .B2(n12507), .A(n12455), .ZN(P3_U3163) );
  INV_X1 U14834 ( .A(n12918), .ZN(n12467) );
  INV_X1 U14835 ( .A(n12458), .ZN(n12461) );
  OAI21_X1 U14836 ( .B1(n12461), .B2(n12460), .A(n12459), .ZN(n12462) );
  NAND3_X1 U14837 ( .A1(n12457), .A2(n12462), .A3(n12533), .ZN(n12466) );
  NAND2_X1 U14838 ( .A1(n12525), .A2(n12550), .ZN(n12463) );
  NAND2_X1 U14839 ( .A1(P3_U3151), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n12642)
         );
  OAI211_X1 U14840 ( .C1(n12865), .C2(n12484), .A(n12463), .B(n12642), .ZN(
        n12464) );
  AOI21_X1 U14841 ( .B1(n12540), .B2(n12867), .A(n12464), .ZN(n12465) );
  OAI211_X1 U14842 ( .C1(n12467), .C2(n12544), .A(n12466), .B(n12465), .ZN(
        P3_U3166) );
  NAND2_X1 U14843 ( .A1(n12540), .A2(n12855), .ZN(n12469) );
  AND2_X1 U14844 ( .A1(P3_U3151), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n12658) );
  AOI21_X1 U14845 ( .B1(n12535), .B2(n12852), .A(n12658), .ZN(n12468) );
  OAI211_X1 U14846 ( .C1(n12470), .C2(n12537), .A(n12469), .B(n12468), .ZN(
        n12477) );
  OAI21_X1 U14847 ( .B1(n12473), .B2(n12472), .A(n12471), .ZN(n12475) );
  AOI21_X1 U14848 ( .B1(n12475), .B2(n12474), .A(n12507), .ZN(n12476) );
  AOI211_X1 U14849 ( .C1(n12987), .C2(n12524), .A(n12477), .B(n12476), .ZN(
        n12478) );
  INV_X1 U14850 ( .A(n12478), .ZN(P3_U3168) );
  INV_X1 U14851 ( .A(n12479), .ZN(n12481) );
  NOR3_X1 U14852 ( .A1(n6546), .A2(n12481), .A3(n12480), .ZN(n12483) );
  OAI21_X1 U14853 ( .B1(n12483), .B2(n12482), .A(n12533), .ZN(n12490) );
  OAI22_X1 U14854 ( .A1(n15345), .A2(n12484), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n15172), .ZN(n12488) );
  INV_X1 U14855 ( .A(n12776), .ZN(n12485) );
  NOR2_X1 U14856 ( .A1(n12486), .A2(n12485), .ZN(n12487) );
  AOI211_X1 U14857 ( .C1(n12525), .C2(n12797), .A(n12488), .B(n12487), .ZN(
        n12489) );
  OAI211_X1 U14858 ( .C1(n12491), .C2(n12544), .A(n12490), .B(n12489), .ZN(
        P3_U3169) );
  XNOR2_X1 U14859 ( .A(n12493), .B(n12492), .ZN(n12498) );
  NAND2_X1 U14860 ( .A1(n12540), .A2(n12820), .ZN(n12495) );
  AOI22_X1 U14861 ( .A1(n12535), .A2(n12817), .B1(P3_REG3_REG_20__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12494) );
  OAI211_X1 U14862 ( .C1(n12838), .C2(n12537), .A(n12495), .B(n12494), .ZN(
        n12496) );
  AOI21_X1 U14863 ( .B1(n12970), .B2(n12524), .A(n12496), .ZN(n12497) );
  OAI21_X1 U14864 ( .B1(n12498), .B2(n12507), .A(n12497), .ZN(P3_U3173) );
  INV_X1 U14865 ( .A(n12499), .ZN(n12500) );
  AOI21_X1 U14866 ( .B1(n12807), .B2(n12501), .A(n12500), .ZN(n12508) );
  NAND2_X1 U14867 ( .A1(n12540), .A2(n12800), .ZN(n12503) );
  AOI22_X1 U14868 ( .A1(n12797), .A2(n12535), .B1(P3_REG3_REG_22__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12502) );
  OAI211_X1 U14869 ( .C1(n12504), .C2(n12537), .A(n12503), .B(n12502), .ZN(
        n12505) );
  AOI21_X1 U14870 ( .B1(n12958), .B2(n12524), .A(n12505), .ZN(n12506) );
  OAI21_X1 U14871 ( .B1(n12508), .B2(n12507), .A(n12506), .ZN(P3_U3175) );
  INV_X1 U14872 ( .A(n12909), .ZN(n12518) );
  OAI21_X1 U14873 ( .B1(n12511), .B2(n12510), .A(n12509), .ZN(n12512) );
  NAND2_X1 U14874 ( .A1(n12512), .A2(n12533), .ZN(n12517) );
  NOR2_X1 U14875 ( .A1(n12513), .A2(P3_STATE_REG_SCAN_IN), .ZN(n12677) );
  AOI21_X1 U14876 ( .B1(n12535), .B2(n12816), .A(n12677), .ZN(n12514) );
  OAI21_X1 U14877 ( .B1(n12865), .B2(n12537), .A(n12514), .ZN(n12515) );
  AOI21_X1 U14878 ( .B1(n12843), .B2(n12540), .A(n12515), .ZN(n12516) );
  OAI211_X1 U14879 ( .C1(n12518), .C2(n12544), .A(n12517), .B(n12516), .ZN(
        P3_U3178) );
  OAI211_X1 U14880 ( .C1(n12521), .C2(n12520), .A(n12519), .B(n12533), .ZN(
        n12530) );
  NAND2_X1 U14881 ( .A1(P3_REG3_REG_6__SCAN_IN), .A2(P3_U3151), .ZN(n14991) );
  INV_X1 U14882 ( .A(n14991), .ZN(n12522) );
  AOI21_X1 U14883 ( .B1(n12524), .B2(n12523), .A(n12522), .ZN(n12529) );
  AOI22_X1 U14884 ( .A1(n12535), .A2(n12556), .B1(n12525), .B2(n15053), .ZN(
        n12528) );
  NAND2_X1 U14885 ( .A1(n12540), .A2(n12526), .ZN(n12527) );
  NAND4_X1 U14886 ( .A1(n12530), .A2(n12529), .A3(n12528), .A4(n12527), .ZN(
        P3_U3179) );
  INV_X1 U14887 ( .A(n12922), .ZN(n12545) );
  OAI21_X1 U14888 ( .B1(n12532), .B2(n12531), .A(n12458), .ZN(n12534) );
  NAND2_X1 U14889 ( .A1(n12534), .A2(n12533), .ZN(n12543) );
  INV_X1 U14890 ( .A(P3_REG3_REG_15__SCAN_IN), .ZN(n15355) );
  NOR2_X1 U14891 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15355), .ZN(n12615) );
  AOI21_X1 U14892 ( .B1(n12535), .B2(n12851), .A(n12615), .ZN(n12536) );
  OAI21_X1 U14893 ( .B1(n12538), .B2(n12537), .A(n12536), .ZN(n12539) );
  AOI21_X1 U14894 ( .B1(n12541), .B2(n12540), .A(n12539), .ZN(n12542) );
  OAI211_X1 U14895 ( .C1(n12545), .C2(n12544), .A(n12543), .B(n12542), .ZN(
        P3_U3181) );
  MUX2_X1 U14896 ( .A(P3_DATAO_REG_31__SCAN_IN), .B(n12546), .S(P3_U3897), .Z(
        P3_U3522) );
  MUX2_X1 U14897 ( .A(n12547), .B(P3_DATAO_REG_30__SCAN_IN), .S(n12548), .Z(
        P3_U3521) );
  MUX2_X1 U14898 ( .A(n12723), .B(P3_DATAO_REG_29__SCAN_IN), .S(n12548), .Z(
        P3_U3520) );
  MUX2_X1 U14899 ( .A(P3_DATAO_REG_27__SCAN_IN), .B(n12750), .S(P3_U3897), .Z(
        P3_U3518) );
  MUX2_X1 U14900 ( .A(P3_DATAO_REG_26__SCAN_IN), .B(n12761), .S(P3_U3897), .Z(
        P3_U3517) );
  MUX2_X1 U14901 ( .A(P3_DATAO_REG_24__SCAN_IN), .B(n12784), .S(P3_U3897), .Z(
        P3_U3515) );
  MUX2_X1 U14902 ( .A(n12797), .B(P3_DATAO_REG_23__SCAN_IN), .S(n12548), .Z(
        P3_U3514) );
  MUX2_X1 U14903 ( .A(n12807), .B(P3_DATAO_REG_22__SCAN_IN), .S(n12548), .Z(
        P3_U3513) );
  MUX2_X1 U14904 ( .A(n12817), .B(P3_DATAO_REG_21__SCAN_IN), .S(n12548), .Z(
        P3_U3512) );
  MUX2_X1 U14905 ( .A(n12826), .B(P3_DATAO_REG_20__SCAN_IN), .S(n12548), .Z(
        P3_U3511) );
  MUX2_X1 U14906 ( .A(P3_DATAO_REG_19__SCAN_IN), .B(n12816), .S(P3_U3897), .Z(
        P3_U3510) );
  MUX2_X1 U14907 ( .A(n12852), .B(P3_DATAO_REG_18__SCAN_IN), .S(n12548), .Z(
        P3_U3509) );
  MUX2_X1 U14908 ( .A(P3_DATAO_REG_17__SCAN_IN), .B(n12549), .S(P3_U3897), .Z(
        P3_U3508) );
  MUX2_X1 U14909 ( .A(P3_DATAO_REG_16__SCAN_IN), .B(n12851), .S(P3_U3897), .Z(
        P3_U3507) );
  MUX2_X1 U14910 ( .A(P3_DATAO_REG_15__SCAN_IN), .B(n12550), .S(P3_U3897), .Z(
        P3_U3506) );
  MUX2_X1 U14911 ( .A(P3_DATAO_REG_14__SCAN_IN), .B(n12551), .S(P3_U3897), .Z(
        P3_U3505) );
  MUX2_X1 U14912 ( .A(P3_DATAO_REG_13__SCAN_IN), .B(n12552), .S(P3_U3897), .Z(
        P3_U3504) );
  MUX2_X1 U14913 ( .A(P3_DATAO_REG_11__SCAN_IN), .B(n12553), .S(P3_U3897), .Z(
        P3_U3502) );
  MUX2_X1 U14914 ( .A(P3_DATAO_REG_10__SCAN_IN), .B(n14427), .S(P3_U3897), .Z(
        P3_U3501) );
  MUX2_X1 U14915 ( .A(P3_DATAO_REG_9__SCAN_IN), .B(n12554), .S(P3_U3897), .Z(
        P3_U3500) );
  MUX2_X1 U14916 ( .A(P3_DATAO_REG_8__SCAN_IN), .B(n12555), .S(P3_U3897), .Z(
        P3_U3499) );
  MUX2_X1 U14917 ( .A(P3_DATAO_REG_7__SCAN_IN), .B(n12556), .S(P3_U3897), .Z(
        P3_U3498) );
  MUX2_X1 U14918 ( .A(P3_DATAO_REG_5__SCAN_IN), .B(n15053), .S(P3_U3897), .Z(
        P3_U3496) );
  MUX2_X1 U14919 ( .A(P3_DATAO_REG_3__SCAN_IN), .B(n15054), .S(P3_U3897), .Z(
        P3_U3494) );
  MUX2_X1 U14920 ( .A(P3_DATAO_REG_2__SCAN_IN), .B(n12557), .S(P3_U3897), .Z(
        P3_U3493) );
  AND2_X1 U14921 ( .A1(n12564), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n12558) );
  AOI21_X1 U14922 ( .B1(n12562), .B2(n12561), .A(n12588), .ZN(n12580) );
  AOI21_X1 U14923 ( .B1(n12565), .B2(n12564), .A(n12563), .ZN(n12567) );
  MUX2_X1 U14924 ( .A(P3_REG2_REG_13__SCAN_IN), .B(P3_REG1_REG_13__SCAN_IN), 
        .S(n12670), .Z(n12583) );
  XOR2_X1 U14925 ( .A(n12583), .B(n12582), .Z(n12566) );
  NAND2_X1 U14926 ( .A1(n12567), .A2(n12566), .ZN(n12581) );
  OAI21_X1 U14927 ( .B1(n12567), .B2(n12566), .A(n12581), .ZN(n12578) );
  AOI21_X1 U14928 ( .B1(n12572), .B2(n12571), .A(n12593), .ZN(n12573) );
  NOR2_X1 U14929 ( .A1(n12573), .A2(n15023), .ZN(n12574) );
  AOI211_X1 U14930 ( .C1(n15001), .C2(P3_ADDR_REG_13__SCAN_IN), .A(n12575), 
        .B(n12574), .ZN(n12576) );
  OAI21_X1 U14931 ( .B1(n12582), .B2(n12701), .A(n12576), .ZN(n12577) );
  AOI21_X1 U14932 ( .B1(n12578), .B2(n15015), .A(n12577), .ZN(n12579) );
  OAI21_X1 U14933 ( .B1(n12580), .B2(n15018), .A(n12579), .ZN(P3_U3195) );
  OAI21_X1 U14934 ( .B1(n12583), .B2(n12582), .A(n12581), .ZN(n12585) );
  NAND2_X1 U14935 ( .A1(n14379), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n12619) );
  OAI21_X1 U14936 ( .B1(P3_REG2_REG_14__SCAN_IN), .B2(n14379), .A(n12619), 
        .ZN(n12594) );
  NAND2_X1 U14937 ( .A1(n14379), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n12618) );
  OAI21_X1 U14938 ( .B1(n14379), .B2(P3_REG1_REG_14__SCAN_IN), .A(n12618), 
        .ZN(n12590) );
  MUX2_X1 U14939 ( .A(n12594), .B(n12590), .S(n12670), .Z(n12584) );
  AOI21_X1 U14940 ( .B1(n12585), .B2(n12584), .A(n14948), .ZN(n12586) );
  NAND2_X1 U14941 ( .A1(n12586), .A2(n12621), .ZN(n12602) );
  INV_X1 U14942 ( .A(n12587), .ZN(n12589) );
  AOI21_X1 U14943 ( .B1(n12590), .B2(n6659), .A(n12608), .ZN(n12591) );
  NOR2_X1 U14944 ( .A1(n12591), .A2(n15018), .ZN(n12600) );
  INV_X1 U14945 ( .A(n15001), .ZN(n15029) );
  INV_X1 U14946 ( .A(P3_ADDR_REG_14__SCAN_IN), .ZN(n12592) );
  NOR2_X1 U14947 ( .A1(n15029), .A2(n12592), .ZN(n12599) );
  AOI21_X1 U14948 ( .B1(n12595), .B2(n12594), .A(n12603), .ZN(n12596) );
  NOR2_X1 U14949 ( .A1(n15023), .A2(n12596), .ZN(n12598) );
  NOR4_X1 U14950 ( .A1(n12600), .A2(n12599), .A3(n12598), .A4(n12597), .ZN(
        n12601) );
  OAI211_X1 U14951 ( .C1(n12701), .C2(n14379), .A(n12602), .B(n12601), .ZN(
        P3_U3196) );
  INV_X1 U14952 ( .A(n12603), .ZN(n12604) );
  INV_X1 U14953 ( .A(n12638), .ZN(n12606) );
  NAND3_X1 U14954 ( .A1(n12619), .A2(n12626), .A3(n12604), .ZN(n12605) );
  NAND2_X1 U14955 ( .A1(n12606), .A2(n12605), .ZN(n12607) );
  AOI21_X1 U14956 ( .B1(n12607), .B2(n15293), .A(n12637), .ZN(n12617) );
  INV_X1 U14957 ( .A(n12629), .ZN(n12611) );
  NAND2_X1 U14958 ( .A1(n12611), .A2(n12610), .ZN(n12612) );
  INV_X1 U14959 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n15387) );
  AOI21_X1 U14960 ( .B1(n12612), .B2(n15387), .A(n12628), .ZN(n12613) );
  NOR2_X1 U14961 ( .A1(n12613), .A2(n15018), .ZN(n12614) );
  AOI211_X1 U14962 ( .C1(n15001), .C2(P3_ADDR_REG_15__SCAN_IN), .A(n12615), 
        .B(n12614), .ZN(n12616) );
  OAI21_X1 U14963 ( .B1(n12617), .B2(n15023), .A(n12616), .ZN(n12625) );
  MUX2_X1 U14964 ( .A(n12619), .B(n12618), .S(n12670), .Z(n12620) );
  MUX2_X1 U14965 ( .A(n15293), .B(n15387), .S(n12670), .Z(n12622) );
  AOI211_X1 U14966 ( .C1(n12623), .C2(n12622), .A(n14948), .B(n12631), .ZN(
        n12624) );
  AOI211_X1 U14967 ( .C1(n15013), .C2(n12626), .A(n12625), .B(n12624), .ZN(
        n12627) );
  INV_X1 U14968 ( .A(n12627), .ZN(P3_U3197) );
  INV_X1 U14969 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n12919) );
  AOI22_X1 U14970 ( .A1(P3_REG1_REG_16__SCAN_IN), .A2(n12636), .B1(n14384), 
        .B2(n12919), .ZN(n12630) );
  AOI21_X1 U14971 ( .B1(n6663), .B2(n12630), .A(n12651), .ZN(n12648) );
  MUX2_X1 U14972 ( .A(P3_REG2_REG_16__SCAN_IN), .B(P3_REG1_REG_16__SCAN_IN), 
        .S(n12670), .Z(n12655) );
  XNOR2_X1 U14973 ( .A(n14384), .B(n12655), .ZN(n12633) );
  NOR2_X1 U14974 ( .A1(n12634), .A2(n12633), .ZN(n12654) );
  AOI211_X1 U14975 ( .C1(n12634), .C2(n12633), .A(n14948), .B(n12654), .ZN(
        n12646) );
  INV_X1 U14976 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n12635) );
  AOI22_X1 U14977 ( .A1(P3_REG2_REG_16__SCAN_IN), .A2(n12636), .B1(n14384), 
        .B2(n12635), .ZN(n12640) );
  AOI21_X1 U14978 ( .B1(n12640), .B2(n12639), .A(n12649), .ZN(n12641) );
  NOR2_X1 U14979 ( .A1(n12641), .A2(n15023), .ZN(n12645) );
  NOR2_X1 U14980 ( .A1(n12701), .A2(n14384), .ZN(n12644) );
  INV_X1 U14981 ( .A(P3_ADDR_REG_16__SCAN_IN), .ZN(n14338) );
  OAI21_X1 U14982 ( .B1(n15029), .B2(n14338), .A(n12642), .ZN(n12643) );
  NOR4_X1 U14983 ( .A1(n12646), .A2(n12645), .A3(n12644), .A4(n12643), .ZN(
        n12647) );
  OAI21_X1 U14984 ( .B1(n12648), .B2(n15018), .A(n12647), .ZN(P3_U3198) );
  INV_X1 U14985 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n12854) );
  AOI21_X1 U14986 ( .B1(n12650), .B2(n12854), .A(n12666), .ZN(n12664) );
  INV_X1 U14987 ( .A(P3_REG1_REG_17__SCAN_IN), .ZN(n12912) );
  AOI21_X1 U14988 ( .B1(n12912), .B2(n12652), .A(n12681), .ZN(n12653) );
  NOR2_X1 U14989 ( .A1(n12653), .A2(n15018), .ZN(n12662) );
  MUX2_X1 U14990 ( .A(P3_REG2_REG_17__SCAN_IN), .B(P3_REG1_REG_17__SCAN_IN), 
        .S(n12670), .Z(n12673) );
  XNOR2_X1 U14991 ( .A(n12672), .B(n12673), .ZN(n12656) );
  NOR2_X1 U14992 ( .A1(n12657), .A2(n12656), .ZN(n12671) );
  AOI211_X1 U14993 ( .C1(n12657), .C2(n12656), .A(n14948), .B(n12671), .ZN(
        n12661) );
  AOI21_X1 U14994 ( .B1(n15001), .B2(P3_ADDR_REG_17__SCAN_IN), .A(n12658), 
        .ZN(n12659) );
  OAI21_X1 U14995 ( .B1(n12701), .B2(n12672), .A(n12659), .ZN(n12660) );
  NOR3_X1 U14996 ( .A1(n12662), .A2(n12661), .A3(n12660), .ZN(n12663) );
  OAI21_X1 U14997 ( .B1(n12664), .B2(n15023), .A(n12663), .ZN(P3_U3199) );
  NAND2_X1 U14998 ( .A1(n12693), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n12689) );
  OAI21_X1 U14999 ( .B1(n12693), .B2(P3_REG2_REG_18__SCAN_IN), .A(n12689), 
        .ZN(n12668) );
  INV_X1 U15000 ( .A(n12690), .ZN(n12667) );
  AOI21_X1 U15001 ( .B1(n12669), .B2(n12668), .A(n12667), .ZN(n12688) );
  MUX2_X1 U15002 ( .A(P3_REG2_REG_18__SCAN_IN), .B(P3_REG1_REG_18__SCAN_IN), 
        .S(n12670), .Z(n12675) );
  NOR2_X1 U15003 ( .A1(n12674), .A2(n12675), .ZN(n12694) );
  AOI21_X1 U15004 ( .B1(n12675), .B2(n12674), .A(n12694), .ZN(n12676) );
  INV_X1 U15005 ( .A(n12676), .ZN(n12686) );
  AOI21_X1 U15006 ( .B1(n15001), .B2(P3_ADDR_REG_18__SCAN_IN), .A(n12677), 
        .ZN(n12678) );
  OAI21_X1 U15007 ( .B1(n12701), .B2(n12693), .A(n12678), .ZN(n12685) );
  NAND2_X1 U15008 ( .A1(n12693), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n12702) );
  OAI21_X1 U15009 ( .B1(n12693), .B2(P3_REG1_REG_18__SCAN_IN), .A(n12702), 
        .ZN(n12682) );
  NAND2_X1 U15010 ( .A1(n12683), .A2(n12682), .ZN(n12684) );
  OAI21_X1 U15011 ( .B1(n12688), .B2(n15023), .A(n12687), .ZN(P3_U3200) );
  XNOR2_X1 U15012 ( .A(n12691), .B(P3_REG2_REG_19__SCAN_IN), .ZN(n12692) );
  XNOR2_X1 U15013 ( .A(n12691), .B(P3_REG1_REG_19__SCAN_IN), .ZN(n12704) );
  MUX2_X1 U15014 ( .A(n12692), .B(n12704), .S(n12670), .Z(n12697) );
  INV_X1 U15015 ( .A(n12693), .ZN(n12695) );
  NAND2_X1 U15016 ( .A1(n15001), .A2(P3_ADDR_REG_19__SCAN_IN), .ZN(n12698) );
  OAI211_X1 U15017 ( .C1(n12701), .C2(n12700), .A(n12699), .B(n12698), .ZN(
        n12705) );
  OAI21_X1 U15018 ( .B1(n12708), .B2(n15023), .A(n12707), .ZN(P3_U3201) );
  INV_X1 U15019 ( .A(P3_REG2_REG_29__SCAN_IN), .ZN(n12710) );
  INV_X1 U15020 ( .A(n12711), .ZN(n12927) );
  NOR2_X1 U15021 ( .A1(n12712), .A2(n12868), .ZN(n14420) );
  AOI21_X1 U15022 ( .B1(n14423), .B2(n12927), .A(n14420), .ZN(n12713) );
  OAI211_X1 U15023 ( .C1(n12930), .C2(n12873), .A(n12714), .B(n12713), .ZN(
        P3_U3204) );
  INV_X1 U15024 ( .A(n12715), .ZN(n12716) );
  NAND2_X1 U15025 ( .A1(n12720), .A2(n12719), .ZN(n12721) );
  NAND3_X1 U15026 ( .A1(n12722), .A2(n15056), .A3(n12721), .ZN(n12725) );
  AOI22_X1 U15027 ( .A1(n12723), .A2(n15052), .B1(n15038), .B2(n12750), .ZN(
        n12724) );
  INV_X1 U15028 ( .A(n12875), .ZN(n12730) );
  AOI22_X1 U15029 ( .A1(n12726), .A2(n15058), .B1(n15066), .B2(
        P3_REG2_REG_28__SCAN_IN), .ZN(n12727) );
  OAI21_X1 U15030 ( .B1(n12728), .B2(n12766), .A(n12727), .ZN(n12729) );
  AOI21_X1 U15031 ( .B1(n12730), .B2(n15049), .A(n12729), .ZN(n12731) );
  OAI21_X1 U15032 ( .B1(n12873), .B2(n12874), .A(n12731), .ZN(P3_U3205) );
  OAI21_X1 U15033 ( .B1(n6600), .B2(n7490), .A(n12734), .ZN(n12738) );
  OAI22_X1 U15034 ( .A1(n12736), .A2(n12866), .B1(n12735), .B2(n12864), .ZN(
        n12737) );
  AOI21_X1 U15035 ( .B1(n12738), .B2(n15056), .A(n12737), .ZN(n12739) );
  OAI21_X1 U15036 ( .B1(n12740), .B2(n15039), .A(n12739), .ZN(n12878) );
  INV_X1 U15037 ( .A(n12878), .ZN(n12746) );
  INV_X1 U15038 ( .A(n12740), .ZN(n12879) );
  AOI22_X1 U15039 ( .A1(n12741), .A2(n15058), .B1(n15066), .B2(
        P3_REG2_REG_27__SCAN_IN), .ZN(n12742) );
  OAI21_X1 U15040 ( .B1(n12937), .B2(n12766), .A(n12742), .ZN(n12743) );
  AOI21_X1 U15041 ( .B1(n12879), .B2(n12744), .A(n12743), .ZN(n12745) );
  OAI21_X1 U15042 ( .B1(n12746), .B2(n15066), .A(n12745), .ZN(P3_U3206) );
  XOR2_X1 U15043 ( .A(n12747), .B(n12748), .Z(n12943) );
  INV_X1 U15044 ( .A(P3_REG2_REG_26__SCAN_IN), .ZN(n12752) );
  XNOR2_X1 U15045 ( .A(n12749), .B(n12748), .ZN(n12751) );
  AOI222_X1 U15046 ( .A1(n15056), .A2(n12751), .B1(n12750), .B2(n15052), .C1(
        n12773), .C2(n15038), .ZN(n12938) );
  MUX2_X1 U15047 ( .A(n12752), .B(n12938), .S(n15049), .Z(n12755) );
  AOI22_X1 U15048 ( .A1(n12940), .A2(n14423), .B1(n15058), .B2(n12753), .ZN(
        n12754) );
  OAI211_X1 U15049 ( .C1(n12873), .C2(n12943), .A(n12755), .B(n12754), .ZN(
        P3_U3207) );
  XNOR2_X1 U15050 ( .A(n12757), .B(n12756), .ZN(n12888) );
  OAI211_X1 U15051 ( .C1(n12760), .C2(n12759), .A(n12758), .B(n15056), .ZN(
        n12763) );
  AOI22_X1 U15052 ( .A1(n12761), .A2(n15052), .B1(n15038), .B2(n12784), .ZN(
        n12762) );
  NAND2_X1 U15053 ( .A1(n12763), .A2(n12762), .ZN(n12885) );
  AOI22_X1 U15054 ( .A1(n15066), .A2(P3_REG2_REG_25__SCAN_IN), .B1(n12764), 
        .B2(n15058), .ZN(n12765) );
  OAI21_X1 U15055 ( .B1(n12767), .B2(n12766), .A(n12765), .ZN(n12768) );
  AOI21_X1 U15056 ( .B1(n12885), .B2(n15049), .A(n12768), .ZN(n12769) );
  OAI21_X1 U15057 ( .B1(n12873), .B2(n12888), .A(n12769), .ZN(P3_U3208) );
  XNOR2_X1 U15058 ( .A(n12772), .B(n12770), .ZN(n12950) );
  INV_X1 U15059 ( .A(P3_REG2_REG_24__SCAN_IN), .ZN(n12775) );
  OAI21_X1 U15060 ( .B1(n6658), .B2(n12772), .A(n12771), .ZN(n12774) );
  AOI222_X1 U15061 ( .A1(n15056), .A2(n12774), .B1(n12773), .B2(n15052), .C1(
        n12797), .C2(n15038), .ZN(n12945) );
  MUX2_X1 U15062 ( .A(n12775), .B(n12945), .S(n15049), .Z(n12778) );
  AOI22_X1 U15063 ( .A1(n12947), .A2(n14423), .B1(n15058), .B2(n12776), .ZN(
        n12777) );
  OAI211_X1 U15064 ( .C1(n12873), .C2(n12950), .A(n12778), .B(n12777), .ZN(
        P3_U3209) );
  XNOR2_X1 U15065 ( .A(n12779), .B(n12780), .ZN(n12953) );
  NAND2_X1 U15066 ( .A1(n12781), .A2(n12780), .ZN(n12782) );
  NAND3_X1 U15067 ( .A1(n12783), .A2(n15056), .A3(n12782), .ZN(n12786) );
  AOI22_X1 U15068 ( .A1(n15052), .A2(n12784), .B1(n12807), .B2(n15038), .ZN(
        n12785) );
  NAND2_X1 U15069 ( .A1(n12786), .A2(n12785), .ZN(n12951) );
  MUX2_X1 U15070 ( .A(P3_REG2_REG_23__SCAN_IN), .B(n12951), .S(n15049), .Z(
        n12787) );
  INV_X1 U15071 ( .A(n12787), .ZN(n12791) );
  AOI22_X1 U15072 ( .A1(n12789), .A2(n14423), .B1(n15058), .B2(n12788), .ZN(
        n12790) );
  OAI211_X1 U15073 ( .C1(n12873), .C2(n12953), .A(n12791), .B(n12790), .ZN(
        P3_U3210) );
  XOR2_X1 U15074 ( .A(n12792), .B(n12795), .Z(n12961) );
  INV_X1 U15075 ( .A(P3_REG2_REG_22__SCAN_IN), .ZN(n12799) );
  NAND2_X1 U15076 ( .A1(n12793), .A2(n12794), .ZN(n12796) );
  XNOR2_X1 U15077 ( .A(n12796), .B(n12795), .ZN(n12798) );
  AOI222_X1 U15078 ( .A1(n15056), .A2(n12798), .B1(n12817), .B2(n15038), .C1(
        n12797), .C2(n15052), .ZN(n12956) );
  MUX2_X1 U15079 ( .A(n12799), .B(n12956), .S(n15049), .Z(n12802) );
  AOI22_X1 U15080 ( .A1(n12958), .A2(n14423), .B1(n15058), .B2(n12800), .ZN(
        n12801) );
  OAI211_X1 U15081 ( .C1(n12873), .C2(n12961), .A(n12802), .B(n12801), .ZN(
        P3_U3211) );
  XNOR2_X1 U15082 ( .A(n12804), .B(n12803), .ZN(n12967) );
  INV_X1 U15083 ( .A(P3_REG2_REG_21__SCAN_IN), .ZN(n12809) );
  OAI21_X1 U15084 ( .B1(n12806), .B2(n12805), .A(n12793), .ZN(n12808) );
  AOI222_X1 U15085 ( .A1(n15056), .A2(n12808), .B1(n12826), .B2(n15038), .C1(
        n12807), .C2(n15052), .ZN(n12962) );
  MUX2_X1 U15086 ( .A(n12809), .B(n12962), .S(n15049), .Z(n12812) );
  AOI22_X1 U15087 ( .A1(n12964), .A2(n14423), .B1(n15058), .B2(n12810), .ZN(
        n12811) );
  OAI211_X1 U15088 ( .C1(n12873), .C2(n12967), .A(n12812), .B(n12811), .ZN(
        P3_U3212) );
  XNOR2_X1 U15089 ( .A(n12814), .B(n12813), .ZN(n12973) );
  INV_X1 U15090 ( .A(P3_REG2_REG_20__SCAN_IN), .ZN(n12819) );
  XOR2_X1 U15091 ( .A(n12815), .B(n12814), .Z(n12818) );
  AOI222_X1 U15092 ( .A1(n15056), .A2(n12818), .B1(n12817), .B2(n15052), .C1(
        n12816), .C2(n15038), .ZN(n12968) );
  MUX2_X1 U15093 ( .A(n12819), .B(n12968), .S(n15049), .Z(n12822) );
  AOI22_X1 U15094 ( .A1(n12970), .A2(n14423), .B1(n15058), .B2(n12820), .ZN(
        n12821) );
  OAI211_X1 U15095 ( .C1(n12873), .C2(n12973), .A(n12822), .B(n12821), .ZN(
        P3_U3213) );
  XOR2_X1 U15096 ( .A(n12825), .B(n12823), .Z(n12976) );
  INV_X1 U15097 ( .A(n12976), .ZN(n12833) );
  INV_X1 U15098 ( .A(P3_REG2_REG_19__SCAN_IN), .ZN(n12828) );
  XOR2_X1 U15099 ( .A(n12825), .B(n12824), .Z(n12827) );
  AOI222_X1 U15100 ( .A1(n15056), .A2(n12827), .B1(n12852), .B2(n15038), .C1(
        n12826), .C2(n15052), .ZN(n12974) );
  MUX2_X1 U15101 ( .A(n12828), .B(n12974), .S(n15049), .Z(n12832) );
  INV_X1 U15102 ( .A(n12979), .ZN(n12830) );
  AOI22_X1 U15103 ( .A1(n12830), .A2(n14423), .B1(n15058), .B2(n12829), .ZN(
        n12831) );
  OAI211_X1 U15104 ( .C1(n12873), .C2(n12833), .A(n12832), .B(n12831), .ZN(
        P3_U3214) );
  INV_X1 U15105 ( .A(n12834), .ZN(n12835) );
  AOI21_X1 U15106 ( .B1(n6716), .B2(n12836), .A(n12835), .ZN(n12837) );
  OAI222_X1 U15107 ( .A1(n12866), .A2(n12838), .B1(n12864), .B2(n12865), .C1(
        n15043), .C2(n12837), .ZN(n12908) );
  NAND2_X1 U15108 ( .A1(n12840), .A2(n12839), .ZN(n12841) );
  NAND2_X1 U15109 ( .A1(n12842), .A2(n12841), .ZN(n12984) );
  AOI22_X1 U15110 ( .A1(n15066), .A2(P3_REG2_REG_18__SCAN_IN), .B1(n15058), 
        .B2(n12843), .ZN(n12845) );
  NAND2_X1 U15111 ( .A1(n12909), .A2(n14423), .ZN(n12844) );
  OAI211_X1 U15112 ( .C1(n12984), .C2(n12873), .A(n12845), .B(n12844), .ZN(
        n12846) );
  AOI21_X1 U15113 ( .B1(n12908), .B2(n15049), .A(n12846), .ZN(n12847) );
  INV_X1 U15114 ( .A(n12847), .ZN(P3_U3215) );
  XNOR2_X1 U15115 ( .A(n12848), .B(n12849), .ZN(n12990) );
  INV_X1 U15116 ( .A(n12990), .ZN(n12858) );
  XOR2_X1 U15117 ( .A(n12850), .B(n12849), .Z(n12853) );
  AOI222_X1 U15118 ( .A1(n15056), .A2(n12853), .B1(n12852), .B2(n15052), .C1(
        n12851), .C2(n15038), .ZN(n12985) );
  MUX2_X1 U15119 ( .A(n12854), .B(n12985), .S(n15049), .Z(n12857) );
  AOI22_X1 U15120 ( .A1(n12987), .A2(n14423), .B1(n15058), .B2(n12855), .ZN(
        n12856) );
  OAI211_X1 U15121 ( .C1(n12873), .C2(n12858), .A(n12857), .B(n12856), .ZN(
        P3_U3216) );
  XOR2_X1 U15122 ( .A(n12859), .B(n12860), .Z(n12995) );
  XOR2_X1 U15123 ( .A(n12861), .B(n12860), .Z(n12862) );
  OAI222_X1 U15124 ( .A1(n12866), .A2(n12865), .B1(n12864), .B2(n12863), .C1(
        n15043), .C2(n12862), .ZN(n12917) );
  NAND2_X1 U15125 ( .A1(n12917), .A2(n15049), .ZN(n12872) );
  INV_X1 U15126 ( .A(n12867), .ZN(n12869) );
  OAI22_X1 U15127 ( .A1(n15049), .A2(n12635), .B1(n12869), .B2(n12868), .ZN(
        n12870) );
  AOI21_X1 U15128 ( .B1(n12918), .B2(n14423), .A(n12870), .ZN(n12871) );
  OAI211_X1 U15129 ( .C1(n12873), .C2(n12995), .A(n12872), .B(n12871), .ZN(
        P3_U3217) );
  AOI21_X1 U15130 ( .B1(n12913), .B2(n12932), .A(n12876), .ZN(n12877) );
  INV_X1 U15131 ( .A(n12877), .ZN(P3_U3487) );
  INV_X1 U15132 ( .A(P3_REG1_REG_27__SCAN_IN), .ZN(n12880) );
  INV_X1 U15133 ( .A(n15101), .ZN(n15108) );
  AOI21_X1 U15134 ( .B1(n15108), .B2(n12879), .A(n12878), .ZN(n12934) );
  MUX2_X1 U15135 ( .A(n12880), .B(n12934), .S(n15131), .Z(n12881) );
  OAI21_X1 U15136 ( .B1(n12937), .B2(n12907), .A(n12881), .ZN(P3_U3486) );
  INV_X1 U15137 ( .A(P3_REG1_REG_26__SCAN_IN), .ZN(n12882) );
  MUX2_X1 U15138 ( .A(n12882), .B(n12938), .S(n15131), .Z(n12884) );
  NAND2_X1 U15139 ( .A1(n12940), .A2(n12913), .ZN(n12883) );
  OAI211_X1 U15140 ( .C1(n12943), .C2(n12924), .A(n12884), .B(n12883), .ZN(
        P3_U3485) );
  AOI21_X1 U15141 ( .B1(n14441), .B2(n12886), .A(n12885), .ZN(n12887) );
  OAI21_X1 U15142 ( .B1(n12889), .B2(n12888), .A(n12887), .ZN(n12944) );
  MUX2_X1 U15143 ( .A(P3_REG1_REG_25__SCAN_IN), .B(n12944), .S(n15131), .Z(
        P3_U3484) );
  INV_X1 U15144 ( .A(P3_REG1_REG_24__SCAN_IN), .ZN(n12890) );
  MUX2_X1 U15145 ( .A(n12890), .B(n12945), .S(n15131), .Z(n12892) );
  NAND2_X1 U15146 ( .A1(n12947), .A2(n12913), .ZN(n12891) );
  OAI211_X1 U15147 ( .C1(n12950), .C2(n12924), .A(n12892), .B(n12891), .ZN(
        P3_U3483) );
  MUX2_X1 U15148 ( .A(P3_REG1_REG_23__SCAN_IN), .B(n12951), .S(n15131), .Z(
        n12894) );
  OAI22_X1 U15149 ( .A1(n12953), .A2(n12924), .B1(n12952), .B2(n12907), .ZN(
        n12893) );
  OR2_X1 U15150 ( .A1(n12894), .A2(n12893), .ZN(P3_U3482) );
  INV_X1 U15151 ( .A(P3_REG1_REG_22__SCAN_IN), .ZN(n12895) );
  MUX2_X1 U15152 ( .A(n12895), .B(n12956), .S(n15131), .Z(n12897) );
  NAND2_X1 U15153 ( .A1(n12958), .A2(n12913), .ZN(n12896) );
  OAI211_X1 U15154 ( .C1(n12961), .C2(n12924), .A(n12897), .B(n12896), .ZN(
        P3_U3481) );
  INV_X1 U15155 ( .A(P3_REG1_REG_21__SCAN_IN), .ZN(n12898) );
  MUX2_X1 U15156 ( .A(n12898), .B(n12962), .S(n15131), .Z(n12900) );
  NAND2_X1 U15157 ( .A1(n12964), .A2(n12913), .ZN(n12899) );
  OAI211_X1 U15158 ( .C1(n12967), .C2(n12924), .A(n12900), .B(n12899), .ZN(
        P3_U3480) );
  MUX2_X1 U15159 ( .A(n12901), .B(n12968), .S(n15131), .Z(n12903) );
  NAND2_X1 U15160 ( .A1(n12970), .A2(n12913), .ZN(n12902) );
  OAI211_X1 U15161 ( .C1(n12924), .C2(n12973), .A(n12903), .B(n12902), .ZN(
        P3_U3479) );
  INV_X1 U15162 ( .A(P3_REG1_REG_19__SCAN_IN), .ZN(n12904) );
  MUX2_X1 U15163 ( .A(n12904), .B(n12974), .S(n15131), .Z(n12906) );
  NAND2_X1 U15164 ( .A1(n12976), .A2(n12914), .ZN(n12905) );
  OAI211_X1 U15165 ( .C1(n12907), .C2(n12979), .A(n12906), .B(n12905), .ZN(
        P3_U3478) );
  INV_X1 U15166 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n12910) );
  AOI21_X1 U15167 ( .B1(n14441), .B2(n12909), .A(n12908), .ZN(n12981) );
  MUX2_X1 U15168 ( .A(n12910), .B(n12981), .S(n15131), .Z(n12911) );
  OAI21_X1 U15169 ( .B1(n12924), .B2(n12984), .A(n12911), .ZN(P3_U3477) );
  MUX2_X1 U15170 ( .A(n12912), .B(n12985), .S(n15131), .Z(n12916) );
  AOI22_X1 U15171 ( .A1(n12990), .A2(n12914), .B1(n12913), .B2(n12987), .ZN(
        n12915) );
  NAND2_X1 U15172 ( .A1(n12916), .A2(n12915), .ZN(P3_U3476) );
  AOI21_X1 U15173 ( .B1(n14441), .B2(n12918), .A(n12917), .ZN(n12993) );
  MUX2_X1 U15174 ( .A(n12919), .B(n12993), .S(n15131), .Z(n12920) );
  OAI21_X1 U15175 ( .B1(n12995), .B2(n12924), .A(n12920), .ZN(P3_U3475) );
  AOI21_X1 U15176 ( .B1(n14441), .B2(n12922), .A(n12921), .ZN(n12996) );
  MUX2_X1 U15177 ( .A(n15387), .B(n12996), .S(n15131), .Z(n12923) );
  OAI21_X1 U15178 ( .B1(n12924), .B2(n13000), .A(n12923), .ZN(P3_U3474) );
  NAND2_X1 U15179 ( .A1(n12988), .A2(n12927), .ZN(n12928) );
  OAI211_X1 U15180 ( .C1(n12930), .C2(n12999), .A(n12929), .B(n12928), .ZN(
        P3_U3456) );
  INV_X1 U15181 ( .A(n12933), .ZN(P3_U3455) );
  MUX2_X1 U15182 ( .A(n12935), .B(n12934), .S(n15110), .Z(n12936) );
  OAI21_X1 U15183 ( .B1(n12937), .B2(n12980), .A(n12936), .ZN(P3_U3454) );
  MUX2_X1 U15184 ( .A(n12939), .B(n12938), .S(n15110), .Z(n12942) );
  NAND2_X1 U15185 ( .A1(n12940), .A2(n12988), .ZN(n12941) );
  OAI211_X1 U15186 ( .C1(n12943), .C2(n12999), .A(n12942), .B(n12941), .ZN(
        P3_U3453) );
  MUX2_X1 U15187 ( .A(P3_REG0_REG_25__SCAN_IN), .B(n12944), .S(n15110), .Z(
        P3_U3452) );
  MUX2_X1 U15188 ( .A(n12946), .B(n12945), .S(n15110), .Z(n12949) );
  NAND2_X1 U15189 ( .A1(n12947), .A2(n12988), .ZN(n12948) );
  OAI211_X1 U15190 ( .C1(n12950), .C2(n12999), .A(n12949), .B(n12948), .ZN(
        P3_U3451) );
  MUX2_X1 U15191 ( .A(P3_REG0_REG_23__SCAN_IN), .B(n12951), .S(n15110), .Z(
        n12955) );
  OAI22_X1 U15192 ( .A1(n12953), .A2(n12999), .B1(n12952), .B2(n12980), .ZN(
        n12954) );
  OR2_X1 U15193 ( .A1(n12955), .A2(n12954), .ZN(P3_U3450) );
  MUX2_X1 U15194 ( .A(n12957), .B(n12956), .S(n15110), .Z(n12960) );
  NAND2_X1 U15195 ( .A1(n12958), .A2(n12988), .ZN(n12959) );
  OAI211_X1 U15196 ( .C1(n12961), .C2(n12999), .A(n12960), .B(n12959), .ZN(
        P3_U3449) );
  MUX2_X1 U15197 ( .A(n12963), .B(n12962), .S(n15110), .Z(n12966) );
  NAND2_X1 U15198 ( .A1(n12964), .A2(n12988), .ZN(n12965) );
  OAI211_X1 U15199 ( .C1(n12967), .C2(n12999), .A(n12966), .B(n12965), .ZN(
        P3_U3448) );
  INV_X1 U15200 ( .A(P3_REG0_REG_20__SCAN_IN), .ZN(n12969) );
  MUX2_X1 U15201 ( .A(n12969), .B(n12968), .S(n15110), .Z(n12972) );
  NAND2_X1 U15202 ( .A1(n12970), .A2(n12988), .ZN(n12971) );
  OAI211_X1 U15203 ( .C1(n12973), .C2(n12999), .A(n12972), .B(n12971), .ZN(
        P3_U3447) );
  MUX2_X1 U15204 ( .A(n12975), .B(n12974), .S(n15110), .Z(n12978) );
  NAND2_X1 U15205 ( .A1(n12976), .A2(n12989), .ZN(n12977) );
  OAI211_X1 U15206 ( .C1(n12980), .C2(n12979), .A(n12978), .B(n12977), .ZN(
        P3_U3446) );
  MUX2_X1 U15207 ( .A(n12982), .B(n12981), .S(n15110), .Z(n12983) );
  OAI21_X1 U15208 ( .B1(n12984), .B2(n12999), .A(n12983), .ZN(P3_U3444) );
  MUX2_X1 U15209 ( .A(n12986), .B(n12985), .S(n15110), .Z(n12992) );
  AOI22_X1 U15210 ( .A1(n12990), .A2(n12989), .B1(n12988), .B2(n12987), .ZN(
        n12991) );
  NAND2_X1 U15211 ( .A1(n12992), .A2(n12991), .ZN(P3_U3441) );
  MUX2_X1 U15212 ( .A(n15276), .B(n12993), .S(n15110), .Z(n12994) );
  OAI21_X1 U15213 ( .B1(n12995), .B2(n12999), .A(n12994), .ZN(P3_U3438) );
  MUX2_X1 U15214 ( .A(n12997), .B(n12996), .S(n15110), .Z(n12998) );
  OAI21_X1 U15215 ( .B1(n13000), .B2(n12999), .A(n12998), .ZN(P3_U3435) );
  MUX2_X1 U15216 ( .A(n13001), .B(P3_D_REG_1__SCAN_IN), .S(n13002), .Z(
        P3_U3377) );
  MUX2_X1 U15217 ( .A(n9069), .B(P3_D_REG_0__SCAN_IN), .S(n13002), .Z(P3_U3376) );
  INV_X1 U15218 ( .A(P3_IR_REG_30__SCAN_IN), .ZN(n13003) );
  NAND3_X1 U15219 ( .A1(n13003), .A2(P3_IR_REG_31__SCAN_IN), .A3(
        P3_STATE_REG_SCAN_IN), .ZN(n13005) );
  OAI22_X1 U15220 ( .A1(n13006), .A2(n13005), .B1(n13004), .B2(n14368), .ZN(
        n13007) );
  AOI21_X1 U15221 ( .B1(n13008), .B2(n14381), .A(n13007), .ZN(n13009) );
  INV_X1 U15222 ( .A(n13009), .ZN(P3_U3264) );
  OAI222_X1 U15223 ( .A1(P3_U3151), .A2(n13012), .B1(n14370), .B2(n13011), 
        .C1(n13010), .C2(n14368), .ZN(P3_U3265) );
  INV_X1 U15224 ( .A(n13013), .ZN(n13014) );
  OAI222_X1 U15225 ( .A1(n14368), .A2(n13015), .B1(n14370), .B2(n13014), .C1(
        n9116), .C2(P3_U3151), .ZN(P3_U3267) );
  INV_X1 U15226 ( .A(n13016), .ZN(n13018) );
  OAI222_X1 U15227 ( .A1(P3_U3151), .A2(n12670), .B1(n14370), .B2(n13018), 
        .C1(n13017), .C2(n14368), .ZN(P3_U3268) );
  INV_X1 U15228 ( .A(n13019), .ZN(n13022) );
  OAI222_X1 U15229 ( .A1(n14370), .A2(n13022), .B1(n14368), .B2(n13021), .C1(
        P3_U3151), .C2(n13020), .ZN(P3_U3269) );
  MUX2_X1 U15230 ( .A(n13023), .B(P3_IR_REG_0__SCAN_IN), .S(
        P3_STATE_REG_SCAN_IN), .Z(P3_U3295) );
  NAND2_X1 U15231 ( .A1(n13294), .A2(n13269), .ZN(n13032) );
  INV_X1 U15232 ( .A(n13032), .ZN(n13035) );
  XNOR2_X1 U15233 ( .A(n13474), .B(n13024), .ZN(n13034) );
  XNOR2_X1 U15234 ( .A(n13486), .B(n13024), .ZN(n13076) );
  AND2_X1 U15235 ( .A1(n13295), .A2(n13269), .ZN(n13026) );
  NAND2_X1 U15236 ( .A1(n13076), .A2(n13026), .ZN(n13027) );
  OAI21_X1 U15237 ( .B1(n13076), .B2(n13026), .A(n13027), .ZN(n13089) );
  XNOR2_X1 U15238 ( .A(n13478), .B(n13024), .ZN(n13028) );
  AND2_X1 U15239 ( .A1(n13142), .A2(n13269), .ZN(n13029) );
  NAND2_X1 U15240 ( .A1(n13028), .A2(n13029), .ZN(n13033) );
  INV_X1 U15241 ( .A(n13028), .ZN(n13126) );
  INV_X1 U15242 ( .A(n13029), .ZN(n13030) );
  NAND2_X1 U15243 ( .A1(n13126), .A2(n13030), .ZN(n13031) );
  AND2_X1 U15244 ( .A1(n13033), .A2(n13031), .ZN(n13075) );
  XNOR2_X1 U15245 ( .A(n13034), .B(n13032), .ZN(n13137) );
  NAND3_X1 U15246 ( .A1(n13074), .A2(n13033), .A3(n13137), .ZN(n13133) );
  XNOR2_X1 U15247 ( .A(n13469), .B(n13024), .ZN(n13037) );
  AND2_X1 U15248 ( .A1(n13141), .A2(n13269), .ZN(n13036) );
  NAND2_X1 U15249 ( .A1(n13037), .A2(n13036), .ZN(n13063) );
  OAI21_X1 U15250 ( .B1(n13037), .B2(n13036), .A(n13063), .ZN(n13038) );
  OAI22_X1 U15251 ( .A1(n13040), .A2(n13538), .B1(n13080), .B2(n13536), .ZN(
        n13262) );
  AOI22_X1 U15252 ( .A1(n13131), .A2(n13262), .B1(P2_REG3_REG_27__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13041) );
  OAI21_X1 U15253 ( .B1(n13266), .B2(n14467), .A(n13041), .ZN(n13042) );
  INV_X1 U15254 ( .A(n13042), .ZN(n13043) );
  AOI21_X1 U15255 ( .B1(n13046), .B2(n13045), .A(n14474), .ZN(n13048) );
  NAND2_X1 U15256 ( .A1(n13048), .A2(n13047), .ZN(n13053) );
  AOI22_X1 U15257 ( .A1(n13050), .A2(n14479), .B1(n13131), .B2(n13049), .ZN(
        n13052) );
  MUX2_X1 U15258 ( .A(n14467), .B(P2_STATE_REG_SCAN_IN), .S(
        P2_REG3_REG_3__SCAN_IN), .Z(n13051) );
  NAND3_X1 U15259 ( .A1(n13053), .A2(n13052), .A3(n13051), .ZN(P2_U3190) );
  NOR3_X1 U15260 ( .A1(n13055), .A2(n13054), .A3(n13124), .ZN(n13056) );
  AOI21_X1 U15261 ( .B1(n6668), .B2(n14462), .A(n13056), .ZN(n13062) );
  AOI22_X1 U15262 ( .A1(n13355), .A2(n13402), .B1(n13401), .B2(n13145), .ZN(
        n13389) );
  NAND2_X1 U15263 ( .A1(P2_U3088), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n13231)
         );
  INV_X1 U15264 ( .A(n14467), .ZN(n13112) );
  NAND2_X1 U15265 ( .A1(n13112), .A2(n13383), .ZN(n13057) );
  OAI211_X1 U15266 ( .C1(n13110), .C2(n13389), .A(n13231), .B(n13057), .ZN(
        n13059) );
  NOR2_X1 U15267 ( .A1(n13101), .A2(n14474), .ZN(n13058) );
  AOI211_X1 U15268 ( .C1(n13516), .C2(n14479), .A(n13059), .B(n13058), .ZN(
        n13060) );
  OAI21_X1 U15269 ( .B1(n13062), .B2(n13061), .A(n13060), .ZN(P2_U3191) );
  INV_X1 U15270 ( .A(n13063), .ZN(n13064) );
  NAND2_X1 U15271 ( .A1(n13065), .A2(n13269), .ZN(n13066) );
  XOR2_X1 U15272 ( .A(n13024), .B(n13066), .Z(n13067) );
  XNOR2_X1 U15273 ( .A(n13464), .B(n13067), .ZN(n13068) );
  NAND2_X1 U15274 ( .A1(n13140), .A2(n13402), .ZN(n13070) );
  NAND2_X1 U15275 ( .A1(n13141), .A2(n13401), .ZN(n13069) );
  NAND2_X1 U15276 ( .A1(n13070), .A2(n13069), .ZN(n13248) );
  AOI22_X1 U15277 ( .A1(n13131), .A2(n13248), .B1(P2_REG3_REG_28__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13071) );
  OAI21_X1 U15278 ( .B1(n13251), .B2(n14467), .A(n13071), .ZN(n13072) );
  AOI21_X1 U15279 ( .B1(n13464), .B2(n14479), .A(n13072), .ZN(n13073) );
  INV_X1 U15280 ( .A(n13074), .ZN(n13128) );
  OR2_X1 U15281 ( .A1(n13088), .A2(n13075), .ZN(n13078) );
  NOR2_X1 U15282 ( .A1(n13081), .A2(n13124), .ZN(n13077) );
  AOI22_X1 U15283 ( .A1(n13078), .A2(n14462), .B1(n13077), .B2(n13076), .ZN(
        n13085) );
  INV_X1 U15284 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n13079) );
  OAI22_X1 U15285 ( .A1(n14467), .A2(n13297), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13079), .ZN(n13083) );
  OAI22_X1 U15286 ( .A1(n13081), .A2(n14470), .B1(n14469), .B2(n13080), .ZN(
        n13082) );
  AOI211_X1 U15287 ( .C1(n13478), .C2(n14479), .A(n13083), .B(n13082), .ZN(
        n13084) );
  OAI21_X1 U15288 ( .B1(n13128), .B2(n13085), .A(n13084), .ZN(P2_U3197) );
  OAI22_X1 U15289 ( .A1(n13086), .A2(n13536), .B1(n13125), .B2(n13538), .ZN(
        n13307) );
  AOI22_X1 U15290 ( .A1(n13307), .A2(n13131), .B1(P2_REG3_REG_24__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13087) );
  OAI21_X1 U15291 ( .B1(n13311), .B2(n14467), .A(n13087), .ZN(n13091) );
  AOI211_X1 U15292 ( .C1(n6662), .C2(n13089), .A(n14474), .B(n13088), .ZN(
        n13090) );
  AOI211_X1 U15293 ( .C1(n13486), .C2(n14479), .A(n13091), .B(n13090), .ZN(
        n13092) );
  INV_X1 U15294 ( .A(n13092), .ZN(P2_U3201) );
  INV_X1 U15295 ( .A(n13376), .ZN(n13094) );
  OAI22_X1 U15296 ( .A1(n14467), .A2(n13094), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13093), .ZN(n13096) );
  OAI22_X1 U15297 ( .A1(n13372), .A2(n14470), .B1(n14469), .B2(n13373), .ZN(
        n13095) );
  AOI211_X1 U15298 ( .C1(n13511), .C2(n14479), .A(n13096), .B(n13095), .ZN(
        n13103) );
  INV_X1 U15299 ( .A(n13097), .ZN(n13100) );
  OAI22_X1 U15300 ( .A1(n13098), .A2(n14474), .B1(n13372), .B2(n13124), .ZN(
        n13099) );
  NAND3_X1 U15301 ( .A1(n13101), .A2(n13100), .A3(n13099), .ZN(n13102) );
  OAI211_X1 U15302 ( .C1(n13104), .C2(n14474), .A(n13103), .B(n13102), .ZN(
        P2_U3205) );
  NAND2_X1 U15303 ( .A1(n13105), .A2(n13356), .ZN(n13109) );
  NAND2_X1 U15304 ( .A1(n14462), .A2(n13106), .ZN(n13108) );
  MUX2_X1 U15305 ( .A(n13109), .B(n13108), .S(n13107), .Z(n13115) );
  INV_X1 U15306 ( .A(n13343), .ZN(n13113) );
  AOI22_X1 U15307 ( .A1(n13143), .A2(n13402), .B1(n13401), .B2(n13144), .ZN(
        n13338) );
  OAI22_X1 U15308 ( .A1(n13338), .A2(n13110), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n15194), .ZN(n13111) );
  AOI21_X1 U15309 ( .B1(n13113), .B2(n13112), .A(n13111), .ZN(n13114) );
  OAI211_X1 U15310 ( .C1(n6905), .C2(n14458), .A(n13115), .B(n13114), .ZN(
        P2_U3207) );
  AOI22_X1 U15311 ( .A1(n13117), .A2(n13403), .B1(n13116), .B2(n13400), .ZN(
        n13118) );
  NAND2_X1 U15312 ( .A1(P2_U3088), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n13209)
         );
  OAI211_X1 U15313 ( .C1(n14467), .C2(n13411), .A(n13118), .B(n13209), .ZN(
        n13122) );
  AOI211_X1 U15314 ( .C1(n13120), .C2(n13119), .A(n14474), .B(n6668), .ZN(
        n13121) );
  AOI211_X1 U15315 ( .C1(n13521), .C2(n14479), .A(n13122), .B(n13121), .ZN(
        n13123) );
  INV_X1 U15316 ( .A(n13123), .ZN(P2_U3210) );
  NOR3_X1 U15317 ( .A1(n13126), .A2(n13125), .A3(n13124), .ZN(n13127) );
  AOI21_X1 U15318 ( .B1(n13128), .B2(n14462), .A(n13127), .ZN(n13138) );
  NAND2_X1 U15319 ( .A1(n13142), .A2(n13401), .ZN(n13130) );
  NAND2_X1 U15320 ( .A1(n13141), .A2(n13402), .ZN(n13129) );
  NAND2_X1 U15321 ( .A1(n13130), .A2(n13129), .ZN(n13285) );
  AOI22_X1 U15322 ( .A1(n13131), .A2(n13285), .B1(P2_REG3_REG_26__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13132) );
  OAI21_X1 U15323 ( .B1(n13280), .B2(n14467), .A(n13132), .ZN(n13135) );
  NOR2_X1 U15324 ( .A1(n13133), .A2(n14474), .ZN(n13134) );
  OAI21_X1 U15325 ( .B1(n13138), .B2(n13137), .A(n13136), .ZN(P2_U3212) );
  INV_X2 U15326 ( .A(P2_U3947), .ZN(n13160) );
  MUX2_X1 U15327 ( .A(n13234), .B(P2_DATAO_REG_31__SCAN_IN), .S(n13160), .Z(
        P2_U3562) );
  MUX2_X1 U15328 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n13139), .S(P2_U3947), .Z(
        P2_U3561) );
  MUX2_X1 U15329 ( .A(n13140), .B(P2_DATAO_REG_29__SCAN_IN), .S(n13160), .Z(
        P2_U3560) );
  MUX2_X1 U15330 ( .A(n13141), .B(P2_DATAO_REG_27__SCAN_IN), .S(n13160), .Z(
        P2_U3558) );
  MUX2_X1 U15331 ( .A(n13294), .B(P2_DATAO_REG_26__SCAN_IN), .S(n13160), .Z(
        P2_U3557) );
  MUX2_X1 U15332 ( .A(n13142), .B(P2_DATAO_REG_25__SCAN_IN), .S(n13160), .Z(
        P2_U3556) );
  MUX2_X1 U15333 ( .A(n13295), .B(P2_DATAO_REG_24__SCAN_IN), .S(n13160), .Z(
        P2_U3555) );
  MUX2_X1 U15334 ( .A(n13143), .B(P2_DATAO_REG_23__SCAN_IN), .S(n13160), .Z(
        P2_U3554) );
  MUX2_X1 U15335 ( .A(n13356), .B(P2_DATAO_REG_22__SCAN_IN), .S(n13160), .Z(
        P2_U3553) );
  MUX2_X1 U15336 ( .A(n13144), .B(P2_DATAO_REG_21__SCAN_IN), .S(n13160), .Z(
        P2_U3552) );
  MUX2_X1 U15337 ( .A(n13355), .B(P2_DATAO_REG_20__SCAN_IN), .S(n13160), .Z(
        P2_U3551) );
  MUX2_X1 U15338 ( .A(n13403), .B(P2_DATAO_REG_19__SCAN_IN), .S(n13160), .Z(
        P2_U3550) );
  MUX2_X1 U15339 ( .A(n13145), .B(P2_DATAO_REG_18__SCAN_IN), .S(n13160), .Z(
        P2_U3549) );
  MUX2_X1 U15340 ( .A(n13400), .B(P2_DATAO_REG_17__SCAN_IN), .S(n13160), .Z(
        P2_U3548) );
  MUX2_X1 U15341 ( .A(n13146), .B(P2_DATAO_REG_16__SCAN_IN), .S(n13160), .Z(
        P2_U3547) );
  MUX2_X1 U15342 ( .A(n13147), .B(P2_DATAO_REG_15__SCAN_IN), .S(n13160), .Z(
        P2_U3546) );
  MUX2_X1 U15343 ( .A(n13148), .B(P2_DATAO_REG_14__SCAN_IN), .S(n13160), .Z(
        P2_U3545) );
  MUX2_X1 U15344 ( .A(n13149), .B(P2_DATAO_REG_13__SCAN_IN), .S(n13160), .Z(
        P2_U3544) );
  MUX2_X1 U15345 ( .A(n13150), .B(P2_DATAO_REG_12__SCAN_IN), .S(n13160), .Z(
        P2_U3543) );
  MUX2_X1 U15346 ( .A(n13151), .B(P2_DATAO_REG_11__SCAN_IN), .S(n13160), .Z(
        P2_U3542) );
  MUX2_X1 U15347 ( .A(n13152), .B(P2_DATAO_REG_10__SCAN_IN), .S(n13160), .Z(
        P2_U3541) );
  MUX2_X1 U15348 ( .A(n13153), .B(P2_DATAO_REG_9__SCAN_IN), .S(n13160), .Z(
        P2_U3540) );
  MUX2_X1 U15349 ( .A(n13154), .B(P2_DATAO_REG_8__SCAN_IN), .S(n13160), .Z(
        P2_U3539) );
  MUX2_X1 U15350 ( .A(n13155), .B(P2_DATAO_REG_7__SCAN_IN), .S(n13160), .Z(
        P2_U3538) );
  MUX2_X1 U15351 ( .A(n13156), .B(P2_DATAO_REG_6__SCAN_IN), .S(n13160), .Z(
        P2_U3537) );
  MUX2_X1 U15352 ( .A(n13157), .B(P2_DATAO_REG_5__SCAN_IN), .S(n13160), .Z(
        P2_U3536) );
  MUX2_X1 U15353 ( .A(n13158), .B(P2_DATAO_REG_4__SCAN_IN), .S(n13160), .Z(
        P2_U3535) );
  MUX2_X1 U15354 ( .A(n13159), .B(P2_DATAO_REG_3__SCAN_IN), .S(n13160), .Z(
        P2_U3534) );
  MUX2_X1 U15355 ( .A(n8301), .B(P2_DATAO_REG_2__SCAN_IN), .S(n13160), .Z(
        P2_U3533) );
  MUX2_X1 U15356 ( .A(n7753), .B(P2_DATAO_REG_1__SCAN_IN), .S(n13160), .Z(
        P2_U3532) );
  MUX2_X1 U15357 ( .A(n8305), .B(P2_DATAO_REG_0__SCAN_IN), .S(n13160), .Z(
        P2_U3531) );
  OAI22_X1 U15358 ( .A1(n14834), .A2(n13162), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13161), .ZN(n13163) );
  AOI21_X1 U15359 ( .B1(n14789), .B2(P2_ADDR_REG_2__SCAN_IN), .A(n13163), .ZN(
        n13173) );
  OAI211_X1 U15360 ( .C1(n13166), .C2(n13165), .A(n14853), .B(n13164), .ZN(
        n13172) );
  INV_X1 U15361 ( .A(n13167), .ZN(n13181) );
  NAND3_X1 U15362 ( .A1(n14795), .A2(n13169), .A3(n13168), .ZN(n13170) );
  NAND3_X1 U15363 ( .A1(n14870), .A2(n13181), .A3(n13170), .ZN(n13171) );
  NAND3_X1 U15364 ( .A1(n13173), .A2(n13172), .A3(n13171), .ZN(P2_U3216) );
  INV_X1 U15365 ( .A(n13174), .ZN(n13175) );
  OAI211_X1 U15366 ( .C1(n13177), .C2(n13176), .A(n14853), .B(n13175), .ZN(
        n13188) );
  INV_X1 U15367 ( .A(n13178), .ZN(n13180) );
  MUX2_X1 U15368 ( .A(n9530), .B(P2_REG2_REG_3__SCAN_IN), .S(n13184), .Z(
        n13179) );
  NAND3_X1 U15369 ( .A1(n13181), .A2(n13180), .A3(n13179), .ZN(n13182) );
  NAND3_X1 U15370 ( .A1(n14870), .A2(n13183), .A3(n13182), .ZN(n13187) );
  AOI22_X1 U15371 ( .A1(n14868), .A2(n13184), .B1(P2_REG3_REG_3__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13186) );
  NAND2_X1 U15372 ( .A1(n14789), .A2(P2_ADDR_REG_3__SCAN_IN), .ZN(n13185) );
  NAND4_X1 U15373 ( .A1(n13188), .A2(n13187), .A3(n13186), .A4(n13185), .ZN(
        P2_U3217) );
  INV_X1 U15374 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n15370) );
  MUX2_X1 U15375 ( .A(n15370), .B(P2_REG1_REG_17__SCAN_IN), .S(n13211), .Z(
        n13191) );
  NAND2_X1 U15376 ( .A1(n13192), .A2(n13191), .ZN(n13206) );
  OAI211_X1 U15377 ( .C1(n13192), .C2(n13191), .A(n13206), .B(n14853), .ZN(
        n13205) );
  AND2_X1 U15378 ( .A1(P2_U3088), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n13194) );
  NOR2_X1 U15379 ( .A1(n14834), .A2(n13211), .ZN(n13193) );
  AOI211_X1 U15380 ( .C1(P2_ADDR_REG_17__SCAN_IN), .C2(n14789), .A(n13194), 
        .B(n13193), .ZN(n13204) );
  INV_X1 U15381 ( .A(n13195), .ZN(n13200) );
  AOI21_X1 U15382 ( .B1(n13211), .B2(P2_REG2_REG_17__SCAN_IN), .A(n13200), 
        .ZN(n13196) );
  OAI21_X1 U15383 ( .B1(P2_REG2_REG_17__SCAN_IN), .B2(n13211), .A(n13196), 
        .ZN(n13201) );
  INV_X1 U15384 ( .A(n13211), .ZN(n13197) );
  NAND2_X1 U15385 ( .A1(n13197), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n13199) );
  INV_X1 U15386 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n13212) );
  NAND2_X1 U15387 ( .A1(n13211), .A2(n13212), .ZN(n13198) );
  OAI211_X1 U15388 ( .C1(n13202), .C2(n13201), .A(n13210), .B(n14870), .ZN(
        n13203) );
  NAND3_X1 U15389 ( .A1(n13205), .A2(n13204), .A3(n13203), .ZN(P2_U3231) );
  OAI21_X1 U15390 ( .B1(n15370), .B2(n13211), .A(n13206), .ZN(n13207) );
  AND2_X1 U15391 ( .A1(n13207), .A2(n13214), .ZN(n13224) );
  OAI21_X1 U15392 ( .B1(n6606), .B2(P2_REG1_REG_18__SCAN_IN), .A(n14853), .ZN(
        n13220) );
  OAI21_X1 U15393 ( .B1(n14834), .B2(n6948), .A(n13209), .ZN(n13218) );
  OAI21_X1 U15394 ( .B1(n13212), .B2(n13211), .A(n13210), .ZN(n13213) );
  AOI21_X1 U15395 ( .B1(P2_REG2_REG_18__SCAN_IN), .B2(n13215), .A(n13222), 
        .ZN(n13216) );
  NOR2_X1 U15396 ( .A1(n13216), .A2(n14836), .ZN(n13217) );
  AOI211_X1 U15397 ( .C1(n14789), .C2(P2_ADDR_REG_18__SCAN_IN), .A(n13218), 
        .B(n13217), .ZN(n13219) );
  OAI21_X1 U15398 ( .B1(n13220), .B2(n13223), .A(n13219), .ZN(P2_U3232) );
  XNOR2_X1 U15399 ( .A(n13225), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n13227) );
  AOI22_X1 U15400 ( .A1(n13228), .A2(n14870), .B1(n14853), .B2(n13227), .ZN(
        n13230) );
  NAND2_X1 U15401 ( .A1(n13546), .A2(n13239), .ZN(n13238) );
  NAND2_X1 U15402 ( .A1(n13234), .A2(n13233), .ZN(n13452) );
  NOR2_X1 U15403 ( .A1(n13419), .A2(n13452), .ZN(n13241) );
  NOR2_X1 U15404 ( .A1(n13543), .A2(n13414), .ZN(n13236) );
  AOI211_X1 U15405 ( .C1(n13419), .C2(P2_REG2_REG_31__SCAN_IN), .A(n13241), 
        .B(n13236), .ZN(n13237) );
  OAI21_X1 U15406 ( .B1(n13450), .B2(n13432), .A(n13237), .ZN(P2_U3234) );
  OAI211_X1 U15407 ( .C1(n13546), .C2(n13239), .A(n13316), .B(n13238), .ZN(
        n13453) );
  NOR2_X1 U15408 ( .A1(n13546), .A2(n13414), .ZN(n13240) );
  AOI211_X1 U15409 ( .C1(n13419), .C2(P2_REG2_REG_30__SCAN_IN), .A(n13241), 
        .B(n13240), .ZN(n13242) );
  OAI21_X1 U15410 ( .B1(n13432), .B2(n13453), .A(n13242), .ZN(P2_U3235) );
  NAND2_X1 U15411 ( .A1(n13245), .A2(n13244), .ZN(n13463) );
  AOI21_X1 U15412 ( .B1(n13247), .B2(n13246), .A(n13534), .ZN(n13250) );
  OAI21_X1 U15413 ( .B1(n13251), .B2(n14877), .A(n13462), .ZN(n13252) );
  NAND2_X1 U15414 ( .A1(n13252), .A2(n13429), .ZN(n13260) );
  INV_X1 U15415 ( .A(n13272), .ZN(n13253) );
  AOI21_X1 U15416 ( .B1(n13464), .B2(n13253), .A(n13269), .ZN(n13254) );
  NAND2_X1 U15417 ( .A1(n13255), .A2(n13254), .ZN(n13461) );
  INV_X1 U15418 ( .A(n13461), .ZN(n13258) );
  INV_X1 U15419 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n13256) );
  OAI22_X1 U15420 ( .A1(n13550), .A2(n13414), .B1(n14884), .B2(n13256), .ZN(
        n13257) );
  AOI21_X1 U15421 ( .B1(n13258), .B2(n13444), .A(n13257), .ZN(n13259) );
  OAI211_X1 U15422 ( .C1(n13393), .C2(n13463), .A(n13260), .B(n13259), .ZN(
        P2_U3237) );
  XNOR2_X1 U15423 ( .A(n13261), .B(n13264), .ZN(n13263) );
  AOI21_X1 U15424 ( .B1(n13263), .B2(n13407), .A(n13262), .ZN(n13472) );
  NAND2_X1 U15425 ( .A1(n13265), .A2(n13264), .ZN(n13466) );
  NAND3_X1 U15426 ( .A1(n13467), .A2(n13466), .A3(n13442), .ZN(n13275) );
  OAI22_X1 U15427 ( .A1(n14884), .A2(n13267), .B1(n13266), .B2(n14877), .ZN(
        n13268) );
  AOI21_X1 U15428 ( .B1(n13469), .B2(n13440), .A(n13268), .ZN(n13274) );
  NAND2_X1 U15429 ( .A1(n13469), .A2(n13278), .ZN(n13270) );
  NAND2_X1 U15430 ( .A1(n13270), .A2(n13316), .ZN(n13271) );
  NOR2_X1 U15431 ( .A1(n13272), .A2(n13271), .ZN(n13468) );
  NAND2_X1 U15432 ( .A1(n13468), .A2(n13444), .ZN(n13273) );
  AND3_X1 U15433 ( .A1(n13275), .A2(n13274), .A3(n13273), .ZN(n13276) );
  OAI21_X1 U15434 ( .B1(n13419), .B2(n13472), .A(n13276), .ZN(P2_U3238) );
  XNOR2_X1 U15435 ( .A(n13277), .B(n13284), .ZN(n13477) );
  INV_X1 U15436 ( .A(n13278), .ZN(n13279) );
  AOI211_X1 U15437 ( .C1(n13474), .C2(n13300), .A(n13269), .B(n13279), .ZN(
        n13473) );
  INV_X1 U15438 ( .A(n13280), .ZN(n13281) );
  AOI22_X1 U15439 ( .A1(n13419), .A2(P2_REG2_REG_26__SCAN_IN), .B1(n13281), 
        .B2(n14487), .ZN(n13282) );
  OAI21_X1 U15440 ( .B1(n7401), .B2(n13414), .A(n13282), .ZN(n13288) );
  XOR2_X1 U15441 ( .A(n13284), .B(n13283), .Z(n13286) );
  AOI21_X1 U15442 ( .B1(n13286), .B2(n13407), .A(n13285), .ZN(n13476) );
  NOR2_X1 U15443 ( .A1(n13476), .A2(n13419), .ZN(n13287) );
  AOI211_X1 U15444 ( .C1(n13473), .C2(n13444), .A(n13288), .B(n13287), .ZN(
        n13289) );
  OAI21_X1 U15445 ( .B1(n13477), .B2(n13393), .A(n13289), .ZN(P2_U3239) );
  XNOR2_X1 U15446 ( .A(n13290), .B(n13292), .ZN(n13482) );
  OAI21_X1 U15447 ( .B1(n13293), .B2(n13292), .A(n13291), .ZN(n13296) );
  AOI222_X1 U15448 ( .A1(n13407), .A2(n13296), .B1(n13295), .B2(n13401), .C1(
        n13294), .C2(n13402), .ZN(n13479) );
  OAI22_X1 U15449 ( .A1(n13429), .A2(n13298), .B1(n13297), .B2(n14877), .ZN(
        n13299) );
  AOI21_X1 U15450 ( .B1(n13478), .B2(n13440), .A(n13299), .ZN(n13303) );
  AOI21_X1 U15451 ( .B1(n13317), .B2(n13478), .A(n13269), .ZN(n13301) );
  AND2_X1 U15452 ( .A1(n13301), .A2(n13300), .ZN(n13481) );
  NAND2_X1 U15453 ( .A1(n13481), .A2(n13444), .ZN(n13302) );
  OAI211_X1 U15454 ( .C1(n13479), .C2(n13419), .A(n13303), .B(n13302), .ZN(
        n13304) );
  AOI21_X1 U15455 ( .B1(n13442), .B2(n13482), .A(n13304), .ZN(n13305) );
  INV_X1 U15456 ( .A(n13305), .ZN(P2_U3240) );
  XNOR2_X1 U15457 ( .A(n13306), .B(n13310), .ZN(n13308) );
  AOI21_X1 U15458 ( .B1(n13308), .B2(n13407), .A(n13307), .ZN(n13488) );
  OAI21_X1 U15459 ( .B1(n6603), .B2(n13310), .A(n13309), .ZN(n13489) );
  INV_X1 U15460 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n13312) );
  OAI22_X1 U15461 ( .A1(n14884), .A2(n13312), .B1(n13311), .B2(n14877), .ZN(
        n13313) );
  AOI21_X1 U15462 ( .B1(n13486), .B2(n13440), .A(n13313), .ZN(n13319) );
  OR2_X1 U15463 ( .A1(n13325), .A2(n13314), .ZN(n13315) );
  AND3_X1 U15464 ( .A1(n13317), .A2(n13316), .A3(n13315), .ZN(n13485) );
  NAND2_X1 U15465 ( .A1(n13485), .A2(n13444), .ZN(n13318) );
  OAI211_X1 U15466 ( .C1(n13489), .C2(n13393), .A(n13319), .B(n13318), .ZN(
        n13320) );
  INV_X1 U15467 ( .A(n13320), .ZN(n13321) );
  OAI21_X1 U15468 ( .B1(n13419), .B2(n13488), .A(n13321), .ZN(P2_U3241) );
  XOR2_X1 U15469 ( .A(n13329), .B(n13322), .Z(n13490) );
  NAND2_X1 U15470 ( .A1(n13326), .A2(n13347), .ZN(n13323) );
  NAND2_X1 U15471 ( .A1(n13323), .A2(n13316), .ZN(n13324) );
  NOR2_X1 U15472 ( .A1(n13325), .A2(n13324), .ZN(n13492) );
  INV_X1 U15473 ( .A(n13326), .ZN(n13560) );
  INV_X1 U15474 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n13327) );
  OAI22_X1 U15475 ( .A1(n13560), .A2(n13414), .B1(n14884), .B2(n13327), .ZN(
        n13335) );
  INV_X1 U15476 ( .A(n13328), .ZN(n13332) );
  XNOR2_X1 U15477 ( .A(n13330), .B(n13329), .ZN(n13331) );
  AOI211_X1 U15478 ( .C1(n14487), .C2(n13332), .A(n13491), .B(n13493), .ZN(
        n13333) );
  NOR2_X1 U15479 ( .A1(n13333), .A2(n13419), .ZN(n13334) );
  AOI211_X1 U15480 ( .C1(n13492), .C2(n13444), .A(n13335), .B(n13334), .ZN(
        n13336) );
  OAI21_X1 U15481 ( .B1(n13490), .B2(n13393), .A(n13336), .ZN(P2_U3242) );
  XNOR2_X1 U15482 ( .A(n13342), .B(n13337), .ZN(n13339) );
  OAI21_X1 U15483 ( .B1(n13339), .B2(n13534), .A(n13338), .ZN(n13498) );
  OAI21_X1 U15484 ( .B1(n13342), .B2(n13341), .A(n13340), .ZN(n13497) );
  INV_X1 U15485 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n13344) );
  OAI22_X1 U15486 ( .A1(n13429), .A2(n13344), .B1(n13343), .B2(n14877), .ZN(
        n13345) );
  AOI21_X1 U15487 ( .B1(n13346), .B2(n13440), .A(n13345), .ZN(n13350) );
  AOI21_X1 U15488 ( .B1(n13346), .B2(n13358), .A(n13269), .ZN(n13348) );
  AND2_X1 U15489 ( .A1(n13348), .A2(n13347), .ZN(n13499) );
  NAND2_X1 U15490 ( .A1(n13499), .A2(n13444), .ZN(n13349) );
  OAI211_X1 U15491 ( .C1(n13497), .C2(n13393), .A(n13350), .B(n13349), .ZN(
        n13351) );
  AOI21_X1 U15492 ( .B1(n14884), .B2(n13498), .A(n13351), .ZN(n13352) );
  INV_X1 U15493 ( .A(n13352), .ZN(P2_U3243) );
  OAI21_X1 U15494 ( .B1(n13354), .B2(n13364), .A(n13353), .ZN(n13357) );
  AOI222_X1 U15495 ( .A1(n13407), .A2(n13357), .B1(n13356), .B2(n13402), .C1(
        n13355), .C2(n13401), .ZN(n13503) );
  AOI211_X1 U15496 ( .C1(n13359), .C2(n13374), .A(n13269), .B(n6906), .ZN(
        n13505) );
  NOR2_X1 U15497 ( .A1(n13567), .A2(n13414), .ZN(n13363) );
  OAI22_X1 U15498 ( .A1(n13429), .A2(n13361), .B1(n13360), .B2(n14877), .ZN(
        n13362) );
  AOI211_X1 U15499 ( .C1(n13505), .C2(n13444), .A(n13363), .B(n13362), .ZN(
        n13367) );
  XNOR2_X1 U15500 ( .A(n13365), .B(n13364), .ZN(n13506) );
  NAND2_X1 U15501 ( .A1(n13506), .A2(n13442), .ZN(n13366) );
  OAI211_X1 U15502 ( .C1(n13503), .C2(n13419), .A(n13367), .B(n13366), .ZN(
        P2_U3244) );
  XOR2_X1 U15503 ( .A(n13368), .B(n13370), .Z(n13513) );
  AOI21_X1 U15504 ( .B1(n13370), .B2(n13369), .A(n6608), .ZN(n13371) );
  OAI222_X1 U15505 ( .A1(n13538), .A2(n13373), .B1(n13536), .B2(n13372), .C1(
        n13534), .C2(n13371), .ZN(n13509) );
  INV_X1 U15506 ( .A(n13374), .ZN(n13375) );
  AOI211_X1 U15507 ( .C1(n13511), .C2(n13382), .A(n13269), .B(n13375), .ZN(
        n13510) );
  NAND2_X1 U15508 ( .A1(n13510), .A2(n13444), .ZN(n13378) );
  AOI22_X1 U15509 ( .A1(n13419), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n13376), 
        .B2(n14487), .ZN(n13377) );
  OAI211_X1 U15510 ( .C1(n7407), .C2(n13414), .A(n13378), .B(n13377), .ZN(
        n13379) );
  AOI21_X1 U15511 ( .B1(n13509), .B2(n14884), .A(n13379), .ZN(n13380) );
  OAI21_X1 U15512 ( .B1(n13513), .B2(n13393), .A(n13380), .ZN(P2_U3245) );
  XOR2_X1 U15513 ( .A(n13381), .B(n13387), .Z(n13518) );
  AOI211_X1 U15514 ( .C1(n13516), .C2(n13409), .A(n13269), .B(n7404), .ZN(
        n13515) );
  INV_X1 U15515 ( .A(n13516), .ZN(n13385) );
  AOI22_X1 U15516 ( .A1(n13419), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n13383), 
        .B2(n14487), .ZN(n13384) );
  OAI21_X1 U15517 ( .B1(n13385), .B2(n13414), .A(n13384), .ZN(n13386) );
  AOI21_X1 U15518 ( .B1(n13515), .B2(n13444), .A(n13386), .ZN(n13392) );
  XNOR2_X1 U15519 ( .A(n13388), .B(n13387), .ZN(n13390) );
  OAI21_X1 U15520 ( .B1(n13390), .B2(n13534), .A(n13389), .ZN(n13514) );
  NAND2_X1 U15521 ( .A1(n13514), .A2(n13429), .ZN(n13391) );
  OAI211_X1 U15522 ( .C1(n13518), .C2(n13393), .A(n13392), .B(n13391), .ZN(
        P2_U3246) );
  XNOR2_X1 U15523 ( .A(n13395), .B(n13394), .ZN(n13408) );
  INV_X1 U15524 ( .A(n13396), .ZN(n13397) );
  AOI21_X1 U15525 ( .B1(n13399), .B2(n13398), .A(n13397), .ZN(n13524) );
  AOI22_X1 U15526 ( .A1(n13403), .A2(n13402), .B1(n13401), .B2(n13400), .ZN(
        n13404) );
  OAI21_X1 U15527 ( .B1(n13524), .B2(n13405), .A(n13404), .ZN(n13406) );
  AOI21_X1 U15528 ( .B1(n13408), .B2(n13407), .A(n13406), .ZN(n13523) );
  INV_X1 U15529 ( .A(n13409), .ZN(n13410) );
  AOI211_X1 U15530 ( .C1(n13521), .C2(n13426), .A(n13269), .B(n13410), .ZN(
        n13520) );
  INV_X1 U15531 ( .A(n13411), .ZN(n13412) );
  AOI22_X1 U15532 ( .A1(n13419), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n13412), 
        .B2(n14487), .ZN(n13413) );
  OAI21_X1 U15533 ( .B1(n7405), .B2(n13414), .A(n13413), .ZN(n13417) );
  NOR2_X1 U15534 ( .A1(n13524), .A2(n13415), .ZN(n13416) );
  AOI211_X1 U15535 ( .C1(n13520), .C2(n13444), .A(n13417), .B(n13416), .ZN(
        n13418) );
  OAI21_X1 U15536 ( .B1(n13419), .B2(n13523), .A(n13418), .ZN(P2_U3247) );
  XOR2_X1 U15537 ( .A(n13423), .B(n13420), .Z(n13422) );
  OAI21_X1 U15538 ( .B1(n13422), .B2(n13534), .A(n13421), .ZN(n14501) );
  INV_X1 U15539 ( .A(n14501), .ZN(n13435) );
  XNOR2_X1 U15540 ( .A(n13424), .B(n13423), .ZN(n14503) );
  AOI21_X1 U15541 ( .B1(n13425), .B2(n14498), .A(n13269), .ZN(n13427) );
  NAND2_X1 U15542 ( .A1(n13427), .A2(n13426), .ZN(n14499) );
  OAI22_X1 U15543 ( .A1(n13429), .A2(n13212), .B1(n13428), .B2(n14877), .ZN(
        n13430) );
  AOI21_X1 U15544 ( .B1(n14498), .B2(n13440), .A(n13430), .ZN(n13431) );
  OAI21_X1 U15545 ( .B1(n14499), .B2(n13432), .A(n13431), .ZN(n13433) );
  AOI21_X1 U15546 ( .B1(n14503), .B2(n13442), .A(n13433), .ZN(n13434) );
  OAI21_X1 U15547 ( .B1(n13435), .B2(n13419), .A(n13434), .ZN(P2_U3248) );
  NAND2_X1 U15548 ( .A1(n13436), .A2(n13429), .ZN(n13449) );
  OAI22_X1 U15549 ( .A1(n13429), .A2(n13438), .B1(n13437), .B2(n14877), .ZN(
        n13439) );
  AOI21_X1 U15550 ( .B1(n13441), .B2(n13440), .A(n13439), .ZN(n13448) );
  NAND2_X1 U15551 ( .A1(n13443), .A2(n13442), .ZN(n13447) );
  NAND2_X1 U15552 ( .A1(n13445), .A2(n13444), .ZN(n13446) );
  NAND4_X1 U15553 ( .A1(n13449), .A2(n13448), .A3(n13447), .A4(n13446), .ZN(
        P2_U3252) );
  AND2_X1 U15554 ( .A1(n13453), .A2(n13452), .ZN(n13544) );
  MUX2_X1 U15555 ( .A(n13454), .B(n13544), .S(n14929), .Z(n13455) );
  OAI21_X1 U15556 ( .B1(n13546), .B2(n13540), .A(n13455), .ZN(P2_U3529) );
  AOI21_X1 U15557 ( .B1(n14899), .B2(n13457), .A(n13456), .ZN(n13458) );
  MUX2_X1 U15558 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n13547), .S(n14929), .Z(
        P2_U3528) );
  NAND3_X1 U15559 ( .A1(n13467), .A2(n13466), .A3(n14515), .ZN(n13471) );
  AOI21_X1 U15560 ( .B1(n14899), .B2(n13469), .A(n13468), .ZN(n13470) );
  NAND3_X1 U15561 ( .A1(n13472), .A2(n13471), .A3(n13470), .ZN(n13551) );
  MUX2_X1 U15562 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n13551), .S(n14929), .Z(
        P2_U3526) );
  AOI21_X1 U15563 ( .B1(n14899), .B2(n13474), .A(n13473), .ZN(n13475) );
  OAI211_X1 U15564 ( .C1(n13519), .C2(n13477), .A(n13476), .B(n13475), .ZN(
        n13552) );
  MUX2_X1 U15565 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n13552), .S(n14929), .Z(
        P2_U3525) );
  INV_X1 U15566 ( .A(n13478), .ZN(n13555) );
  INV_X1 U15567 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n13483) );
  INV_X1 U15568 ( .A(n13479), .ZN(n13480) );
  AOI211_X1 U15569 ( .C1(n14515), .C2(n13482), .A(n13481), .B(n13480), .ZN(
        n13553) );
  MUX2_X1 U15570 ( .A(n13483), .B(n13553), .S(n14929), .Z(n13484) );
  OAI21_X1 U15571 ( .B1(n13555), .B2(n13540), .A(n13484), .ZN(P2_U3524) );
  AOI21_X1 U15572 ( .B1(n14899), .B2(n13486), .A(n13485), .ZN(n13487) );
  OAI211_X1 U15573 ( .C1(n13489), .C2(n13519), .A(n13488), .B(n13487), .ZN(
        n13556) );
  MUX2_X1 U15574 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n13556), .S(n14929), .Z(
        P2_U3523) );
  NOR2_X1 U15575 ( .A1(n13490), .A2(n13519), .ZN(n13494) );
  NOR4_X1 U15576 ( .A1(n13494), .A2(n13493), .A3(n13492), .A4(n13491), .ZN(
        n13557) );
  MUX2_X1 U15577 ( .A(n13495), .B(n13557), .S(n14929), .Z(n13496) );
  OAI21_X1 U15578 ( .B1(n13560), .B2(n13540), .A(n13496), .ZN(P2_U3522) );
  INV_X1 U15579 ( .A(n13497), .ZN(n13500) );
  AOI211_X1 U15580 ( .C1(n13500), .C2(n14515), .A(n13499), .B(n13498), .ZN(
        n13561) );
  MUX2_X1 U15581 ( .A(n13501), .B(n13561), .S(n14929), .Z(n13502) );
  OAI21_X1 U15582 ( .B1(n6905), .B2(n13540), .A(n13502), .ZN(P2_U3521) );
  INV_X1 U15583 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n13507) );
  INV_X1 U15584 ( .A(n13503), .ZN(n13504) );
  AOI211_X1 U15585 ( .C1(n14515), .C2(n13506), .A(n13505), .B(n13504), .ZN(
        n13564) );
  MUX2_X1 U15586 ( .A(n13507), .B(n13564), .S(n14929), .Z(n13508) );
  OAI21_X1 U15587 ( .B1(n13567), .B2(n13540), .A(n13508), .ZN(P2_U3520) );
  AOI211_X1 U15588 ( .C1(n14899), .C2(n13511), .A(n13510), .B(n13509), .ZN(
        n13512) );
  OAI21_X1 U15589 ( .B1(n13519), .B2(n13513), .A(n13512), .ZN(n13568) );
  MUX2_X1 U15590 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n13568), .S(n14929), .Z(
        P2_U3519) );
  AOI211_X1 U15591 ( .C1(n14899), .C2(n13516), .A(n13515), .B(n13514), .ZN(
        n13517) );
  OAI21_X1 U15592 ( .B1(n13519), .B2(n13518), .A(n13517), .ZN(n13569) );
  MUX2_X1 U15593 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n13569), .S(n14929), .Z(
        P2_U3518) );
  AOI21_X1 U15594 ( .B1(n14899), .B2(n13521), .A(n13520), .ZN(n13522) );
  OAI211_X1 U15595 ( .C1(n13524), .C2(n14901), .A(n13523), .B(n13522), .ZN(
        n13570) );
  MUX2_X1 U15596 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n13570), .S(n14929), .Z(
        P2_U3517) );
  INV_X1 U15597 ( .A(n14489), .ZN(n13574) );
  XNOR2_X1 U15598 ( .A(n13525), .B(n13529), .ZN(n14496) );
  AOI211_X1 U15599 ( .C1(n14489), .C2(n13527), .A(n13269), .B(n13526), .ZN(
        n14484) );
  NAND3_X1 U15600 ( .A1(n13530), .A2(n13529), .A3(n13528), .ZN(n13531) );
  AND2_X1 U15601 ( .A1(n13532), .A2(n13531), .ZN(n13533) );
  OAI222_X1 U15602 ( .A1(n13538), .A2(n13537), .B1(n13536), .B2(n13535), .C1(
        n13534), .C2(n13533), .ZN(n14493) );
  AOI211_X1 U15603 ( .C1(n14496), .C2(n14515), .A(n14484), .B(n14493), .ZN(
        n13571) );
  MUX2_X1 U15604 ( .A(n7990), .B(n13571), .S(n14929), .Z(n13539) );
  OAI21_X1 U15605 ( .B1(n13574), .B2(n13540), .A(n13539), .ZN(P2_U3514) );
  INV_X1 U15606 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n13542) );
  MUX2_X1 U15607 ( .A(n15402), .B(n13544), .S(n14925), .Z(n13545) );
  OAI21_X1 U15608 ( .B1(n13546), .B2(n13573), .A(n13545), .ZN(P2_U3497) );
  MUX2_X1 U15609 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n13547), .S(n14925), .Z(
        P2_U3496) );
  OAI21_X1 U15610 ( .B1(n13550), .B2(n13573), .A(n13549), .ZN(P2_U3495) );
  MUX2_X1 U15611 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n13551), .S(n14925), .Z(
        P2_U3494) );
  MUX2_X1 U15612 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n13552), .S(n14925), .Z(
        P2_U3493) );
  MUX2_X1 U15613 ( .A(n15409), .B(n13553), .S(n14925), .Z(n13554) );
  OAI21_X1 U15614 ( .B1(n13555), .B2(n13573), .A(n13554), .ZN(P2_U3492) );
  MUX2_X1 U15615 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n13556), .S(n14925), .Z(
        P2_U3491) );
  INV_X1 U15616 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n13558) );
  MUX2_X1 U15617 ( .A(n13558), .B(n13557), .S(n14925), .Z(n13559) );
  OAI21_X1 U15618 ( .B1(n13560), .B2(n13573), .A(n13559), .ZN(P2_U3490) );
  INV_X1 U15619 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n13562) );
  MUX2_X1 U15620 ( .A(n13562), .B(n13561), .S(n14925), .Z(n13563) );
  OAI21_X1 U15621 ( .B1(n6905), .B2(n13573), .A(n13563), .ZN(P2_U3489) );
  INV_X1 U15622 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n13565) );
  MUX2_X1 U15623 ( .A(n13565), .B(n13564), .S(n14925), .Z(n13566) );
  OAI21_X1 U15624 ( .B1(n13567), .B2(n13573), .A(n13566), .ZN(P2_U3488) );
  MUX2_X1 U15625 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n13568), .S(n14925), .Z(
        P2_U3487) );
  MUX2_X1 U15626 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n13569), .S(n14925), .Z(
        P2_U3486) );
  MUX2_X1 U15627 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n13570), .S(n14925), .Z(
        P2_U3484) );
  INV_X1 U15628 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n15169) );
  MUX2_X1 U15629 ( .A(n15169), .B(n13571), .S(n14925), .Z(n13572) );
  OAI21_X1 U15630 ( .B1(n13574), .B2(n13573), .A(n13572), .ZN(P2_U3475) );
  INV_X1 U15631 ( .A(n13575), .ZN(n14246) );
  NAND3_X1 U15632 ( .A1(n13576), .A2(P2_IR_REG_31__SCAN_IN), .A3(
        P2_STATE_REG_SCAN_IN), .ZN(n13578) );
  OAI22_X1 U15633 ( .A1(n7468), .A2(n13578), .B1(n13577), .B2(n13588), .ZN(
        n13579) );
  INV_X1 U15634 ( .A(n13579), .ZN(n13580) );
  OAI21_X1 U15635 ( .B1(n14246), .B2(n13596), .A(n13580), .ZN(P2_U3296) );
  OAI222_X1 U15636 ( .A1(n13596), .A2(n13582), .B1(P2_U3088), .B2(n7740), .C1(
        n13581), .C2(n13594), .ZN(P2_U3298) );
  NAND2_X1 U15637 ( .A1(n13584), .A2(n13583), .ZN(n13586) );
  OAI211_X1 U15638 ( .C1(n13588), .C2(n13587), .A(n13586), .B(n13585), .ZN(
        P2_U3299) );
  AOI21_X1 U15639 ( .B1(P1_DATAO_REG_27__SCAN_IN), .B2(n13590), .A(n13589), 
        .ZN(n13591) );
  OAI21_X1 U15640 ( .B1(n13592), .B2(n13596), .A(n13591), .ZN(P2_U3300) );
  INV_X1 U15641 ( .A(n13593), .ZN(n14248) );
  OAI222_X1 U15642 ( .A1(P2_U3088), .A2(n13597), .B1(n13596), .B2(n14248), 
        .C1(n13595), .C2(n13594), .ZN(P2_U3301) );
  INV_X1 U15643 ( .A(n13599), .ZN(n13600) );
  MUX2_X1 U15644 ( .A(n13600), .B(n15330), .S(P2_STATE_REG_SCAN_IN), .Z(
        P2_U3327) );
  INV_X1 U15645 ( .A(n13601), .ZN(n13613) );
  NAND2_X1 U15646 ( .A1(n13891), .A2(n14742), .ZN(n14148) );
  OAI21_X1 U15647 ( .B1(n13604), .B2(n13603), .A(n13602), .ZN(n13605) );
  NAND2_X1 U15648 ( .A1(n13605), .A2(n14535), .ZN(n13612) );
  INV_X1 U15649 ( .A(n13606), .ZN(n13610) );
  OAI22_X1 U15650 ( .A1(n13715), .A2(n13608), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13607), .ZN(n13609) );
  AOI21_X1 U15651 ( .B1(n13610), .B2(n13717), .A(n13609), .ZN(n13611) );
  OAI211_X1 U15652 ( .C1(n13613), .C2(n14148), .A(n13612), .B(n13611), .ZN(
        P1_U3214) );
  OAI21_X1 U15653 ( .B1(n13615), .B2(n13614), .A(n13686), .ZN(n13616) );
  NAND2_X1 U15654 ( .A1(n13616), .A2(n14535), .ZN(n13622) );
  INV_X1 U15655 ( .A(n13978), .ZN(n13620) );
  AND2_X1 U15656 ( .A1(n13757), .A2(n13732), .ZN(n13617) );
  AOI21_X1 U15657 ( .B1(n13759), .B2(n13897), .A(n13617), .ZN(n14169) );
  INV_X1 U15658 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n13618) );
  OAI22_X1 U15659 ( .A1(n14169), .A2(n13715), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13618), .ZN(n13619) );
  AOI21_X1 U15660 ( .B1(n13620), .B2(n13717), .A(n13619), .ZN(n13621) );
  OAI211_X1 U15661 ( .C1(n14171), .C2(n13753), .A(n13622), .B(n13621), .ZN(
        P1_U3216) );
  INV_X1 U15662 ( .A(n14197), .ZN(n13631) );
  OAI211_X1 U15663 ( .C1(n13625), .C2(n13624), .A(n13623), .B(n14535), .ZN(
        n13630) );
  OAI22_X1 U15664 ( .A1(n13627), .A2(n14678), .B1(n13626), .B2(n13674), .ZN(
        n14196) );
  AND2_X1 U15665 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n13871) );
  NOR2_X1 U15666 ( .A1(n14542), .A2(n14041), .ZN(n13628) );
  AOI211_X1 U15667 ( .C1(n14537), .C2(n14196), .A(n13871), .B(n13628), .ZN(
        n13629) );
  OAI211_X1 U15668 ( .C1(n13631), .C2(n13753), .A(n13630), .B(n13629), .ZN(
        P1_U3219) );
  OAI21_X1 U15669 ( .B1(n13634), .B2(n13633), .A(n13632), .ZN(n13635) );
  NAND2_X1 U15670 ( .A1(n13635), .A2(n14535), .ZN(n13640) );
  INV_X1 U15671 ( .A(n13636), .ZN(n14012) );
  AOI22_X1 U15672 ( .A1(n13759), .A2(n13732), .B1(n13897), .B2(n13761), .ZN(
        n14004) );
  OAI22_X1 U15673 ( .A1(n14004), .A2(n13715), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13637), .ZN(n13638) );
  AOI21_X1 U15674 ( .B1(n14012), .B2(n13717), .A(n13638), .ZN(n13639) );
  OAI211_X1 U15675 ( .C1(n14183), .C2(n13753), .A(n13640), .B(n13639), .ZN(
        P1_U3223) );
  AND2_X1 U15676 ( .A1(n11649), .A2(n13641), .ZN(n13644) );
  OAI211_X1 U15677 ( .C1(n13644), .C2(n13643), .A(n14535), .B(n13642), .ZN(
        n13650) );
  NOR2_X1 U15678 ( .A1(n14542), .A2(n13645), .ZN(n13646) );
  AOI211_X1 U15679 ( .C1(n14537), .C2(n13648), .A(n13647), .B(n13646), .ZN(
        n13649) );
  OAI211_X1 U15680 ( .C1(n14393), .C2(n13753), .A(n13650), .B(n13649), .ZN(
        P1_U3224) );
  NAND2_X1 U15681 ( .A1(n13757), .A2(n13897), .ZN(n13652) );
  NAND2_X1 U15682 ( .A1(n13755), .A2(n13732), .ZN(n13651) );
  NAND2_X1 U15683 ( .A1(n13652), .A2(n13651), .ZN(n14158) );
  AOI22_X1 U15684 ( .A1(n14537), .A2(n14158), .B1(P1_REG3_REG_25__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13653) );
  OAI21_X1 U15685 ( .B1(n13946), .B2(n14542), .A(n13653), .ZN(n13659) );
  AOI21_X1 U15686 ( .B1(n13657), .B2(n13656), .A(n13727), .ZN(n13658) );
  INV_X1 U15687 ( .A(n13671), .ZN(n13662) );
  AOI21_X1 U15688 ( .B1(n6745), .B2(n13740), .A(n13660), .ZN(n13661) );
  OAI21_X1 U15689 ( .B1(n13662), .B2(n13661), .A(n14535), .ZN(n13668) );
  OR2_X1 U15690 ( .A1(n13663), .A2(n13674), .ZN(n13665) );
  NAND2_X1 U15691 ( .A1(n13764), .A2(n13732), .ZN(n13664) );
  NAND2_X1 U15692 ( .A1(n13665), .A2(n13664), .ZN(n14087) );
  AND2_X1 U15693 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n13798) );
  NOR2_X1 U15694 ( .A1(n14542), .A2(n14088), .ZN(n13666) );
  AOI211_X1 U15695 ( .C1(n14537), .C2(n14087), .A(n13798), .B(n13666), .ZN(
        n13667) );
  OAI211_X1 U15696 ( .C1(n14215), .C2(n13753), .A(n13668), .B(n13667), .ZN(
        P1_U3226) );
  INV_X1 U15697 ( .A(n14209), .ZN(n14074) );
  AND3_X1 U15698 ( .A1(n13671), .A2(n13670), .A3(n13669), .ZN(n13672) );
  OAI21_X1 U15699 ( .B1(n13673), .B2(n13672), .A(n14535), .ZN(n13679) );
  OR2_X1 U15700 ( .A1(n13746), .A2(n13674), .ZN(n13676) );
  NAND2_X1 U15701 ( .A1(n13763), .A2(n13732), .ZN(n13675) );
  NAND2_X1 U15702 ( .A1(n13676), .A2(n13675), .ZN(n14068) );
  AND2_X1 U15703 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n13818) );
  NOR2_X1 U15704 ( .A1(n14542), .A2(n14071), .ZN(n13677) );
  AOI211_X1 U15705 ( .C1(n14537), .C2(n14068), .A(n13818), .B(n13677), .ZN(
        n13678) );
  OAI211_X1 U15706 ( .C1(n14074), .C2(n13753), .A(n13679), .B(n13678), .ZN(
        P1_U3228) );
  NAND2_X1 U15707 ( .A1(n13758), .A2(n13897), .ZN(n13681) );
  NAND2_X1 U15708 ( .A1(n13756), .A2(n13732), .ZN(n13680) );
  NAND2_X1 U15709 ( .A1(n13681), .A2(n13680), .ZN(n13959) );
  AOI22_X1 U15710 ( .A1(n14537), .A2(n13959), .B1(P1_REG3_REG_24__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13682) );
  OAI21_X1 U15711 ( .B1(n13964), .B2(n14542), .A(n13682), .ZN(n13690) );
  INV_X1 U15712 ( .A(n13683), .ZN(n13688) );
  NAND3_X1 U15713 ( .A1(n13686), .A2(n13685), .A3(n13684), .ZN(n13687) );
  AOI21_X1 U15714 ( .B1(n13688), .B2(n13687), .A(n13727), .ZN(n13689) );
  AOI211_X1 U15715 ( .C1(n14533), .C2(n14165), .A(n13690), .B(n13689), .ZN(
        n13691) );
  INV_X1 U15716 ( .A(n13691), .ZN(P1_U3229) );
  XNOR2_X1 U15717 ( .A(n13693), .B(n13692), .ZN(n13698) );
  NOR2_X1 U15718 ( .A1(n14542), .A2(n14024), .ZN(n13696) );
  AND2_X1 U15719 ( .A1(n13762), .A2(n13897), .ZN(n13694) );
  AOI21_X1 U15720 ( .B1(n13760), .B2(n13732), .A(n13694), .ZN(n14022) );
  OAI22_X1 U15721 ( .A1(n14022), .A2(n13715), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n15196), .ZN(n13695) );
  AOI211_X1 U15722 ( .C1(n14029), .C2(n14533), .A(n13696), .B(n13695), .ZN(
        n13697) );
  OAI21_X1 U15723 ( .B1(n13698), .B2(n13727), .A(n13697), .ZN(P1_U3233) );
  XNOR2_X1 U15724 ( .A(n13700), .B(n13699), .ZN(n13708) );
  NAND2_X1 U15725 ( .A1(n14537), .A2(n13701), .ZN(n13702) );
  OAI211_X1 U15726 ( .C1(n14542), .C2(n13704), .A(n13703), .B(n13702), .ZN(
        n13705) );
  AOI21_X1 U15727 ( .B1(n13706), .B2(n14533), .A(n13705), .ZN(n13707) );
  OAI21_X1 U15728 ( .B1(n13708), .B2(n13727), .A(n13707), .ZN(P1_U3234) );
  OAI21_X1 U15729 ( .B1(n13711), .B2(n13710), .A(n13709), .ZN(n13712) );
  NAND2_X1 U15730 ( .A1(n13712), .A2(n14535), .ZN(n13719) );
  INV_X1 U15731 ( .A(n13713), .ZN(n13994) );
  AOI22_X1 U15732 ( .A1(n13760), .A2(n13897), .B1(n13732), .B2(n13758), .ZN(
        n13989) );
  INV_X1 U15733 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n13714) );
  OAI22_X1 U15734 ( .A1(n13989), .A2(n13715), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13714), .ZN(n13716) );
  AOI21_X1 U15735 ( .B1(n13994), .B2(n13717), .A(n13716), .ZN(n13718) );
  OAI211_X1 U15736 ( .C1(n13753), .C2(n13997), .A(n13719), .B(n13718), .ZN(
        P1_U3235) );
  AOI21_X1 U15737 ( .B1(n6677), .B2(n13721), .A(n13720), .ZN(n13728) );
  NAND2_X1 U15738 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n13840)
         );
  NAND2_X1 U15739 ( .A1(n13762), .A2(n13732), .ZN(n13723) );
  NAND2_X1 U15740 ( .A1(n13764), .A2(n13897), .ZN(n13722) );
  NAND2_X1 U15741 ( .A1(n13723), .A2(n13722), .ZN(n14203) );
  NAND2_X1 U15742 ( .A1(n14537), .A2(n14203), .ZN(n13724) );
  OAI211_X1 U15743 ( .C1(n14542), .C2(n14060), .A(n13840), .B(n13724), .ZN(
        n13725) );
  AOI21_X1 U15744 ( .B1(n14204), .B2(n14533), .A(n13725), .ZN(n13726) );
  OAI21_X1 U15745 ( .B1(n13728), .B2(n13727), .A(n13726), .ZN(P1_U3238) );
  OAI21_X1 U15746 ( .B1(n13731), .B2(n13730), .A(n13729), .ZN(n13738) );
  NAND2_X1 U15747 ( .A1(n14153), .A2(n14533), .ZN(n13736) );
  NAND2_X1 U15748 ( .A1(n13908), .A2(n13732), .ZN(n13734) );
  NAND2_X1 U15749 ( .A1(n13756), .A2(n13897), .ZN(n13733) );
  NAND2_X1 U15750 ( .A1(n13734), .A2(n13733), .ZN(n14152) );
  AOI22_X1 U15751 ( .A1(n14537), .A2(n14152), .B1(P1_REG3_REG_26__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13735) );
  OAI211_X1 U15752 ( .C1(n14542), .C2(n13934), .A(n13736), .B(n13735), .ZN(
        n13737) );
  AOI21_X1 U15753 ( .B1(n13738), .B2(n14535), .A(n13737), .ZN(n13739) );
  INV_X1 U15754 ( .A(n13739), .ZN(P1_U3240) );
  INV_X1 U15755 ( .A(n14115), .ZN(n14544) );
  INV_X1 U15756 ( .A(n13740), .ZN(n13744) );
  OAI21_X1 U15757 ( .B1(n13742), .B2(n13744), .A(n13741), .ZN(n13743) );
  OAI211_X1 U15758 ( .C1(n6745), .C2(n13744), .A(n13743), .B(n14535), .ZN(
        n13752) );
  OR2_X1 U15759 ( .A1(n13746), .A2(n14678), .ZN(n13748) );
  NAND2_X1 U15760 ( .A1(n13766), .A2(n13897), .ZN(n13747) );
  NAND2_X1 U15761 ( .A1(n13748), .A2(n13747), .ZN(n14100) );
  NAND2_X1 U15762 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n14622)
         );
  INV_X1 U15763 ( .A(n14622), .ZN(n13750) );
  NOR2_X1 U15764 ( .A1(n14542), .A2(n14111), .ZN(n13749) );
  AOI211_X1 U15765 ( .C1(n14537), .C2(n14100), .A(n13750), .B(n13749), .ZN(
        n13751) );
  OAI211_X1 U15766 ( .C1(n14544), .C2(n13753), .A(n13752), .B(n13751), .ZN(
        P1_U3241) );
  MUX2_X1 U15767 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n13899), .S(P1_U4016), .Z(
        P1_U3590) );
  MUX2_X1 U15768 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n13754), .S(n13777), .Z(
        P1_U3589) );
  MUX2_X1 U15769 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n13908), .S(n13777), .Z(
        P1_U3587) );
  MUX2_X1 U15770 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n13755), .S(n13777), .Z(
        P1_U3586) );
  MUX2_X1 U15771 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n13756), .S(n13777), .Z(
        P1_U3585) );
  MUX2_X1 U15772 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n13757), .S(n13777), .Z(
        P1_U3584) );
  MUX2_X1 U15773 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n13758), .S(n13777), .Z(
        P1_U3583) );
  MUX2_X1 U15774 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n13759), .S(n13777), .Z(
        P1_U3582) );
  MUX2_X1 U15775 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n13760), .S(n13777), .Z(
        P1_U3581) );
  MUX2_X1 U15776 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n13761), .S(n13777), .Z(
        P1_U3580) );
  MUX2_X1 U15777 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n13762), .S(P1_U4016), .Z(
        P1_U3579) );
  MUX2_X1 U15778 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n13763), .S(n13777), .Z(
        P1_U3578) );
  MUX2_X1 U15779 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n13764), .S(n13777), .Z(
        P1_U3577) );
  MUX2_X1 U15780 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n13765), .S(n13777), .Z(
        P1_U3576) );
  MUX2_X1 U15781 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n13766), .S(n13777), .Z(
        P1_U3574) );
  MUX2_X1 U15782 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n13767), .S(n13777), .Z(
        P1_U3573) );
  MUX2_X1 U15783 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n13768), .S(n13777), .Z(
        P1_U3572) );
  MUX2_X1 U15784 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n13769), .S(n13777), .Z(
        P1_U3571) );
  MUX2_X1 U15785 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n13770), .S(n13777), .Z(
        P1_U3570) );
  MUX2_X1 U15786 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n13771), .S(n13777), .Z(
        P1_U3569) );
  MUX2_X1 U15787 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n13772), .S(n13777), .Z(
        P1_U3568) );
  MUX2_X1 U15788 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n13773), .S(n13777), .Z(
        P1_U3567) );
  MUX2_X1 U15789 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n13774), .S(n13777), .Z(
        P1_U3566) );
  MUX2_X1 U15790 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n13775), .S(n13777), .Z(
        P1_U3564) );
  MUX2_X1 U15791 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n13776), .S(n13777), .Z(
        P1_U3563) );
  MUX2_X1 U15792 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n13778), .S(n13777), .Z(
        P1_U3562) );
  MUX2_X1 U15793 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n6770), .S(P1_U4016), .Z(
        P1_U3561) );
  MUX2_X1 U15794 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n13780), .S(P1_U4016), .Z(
        P1_U3560) );
  NAND2_X1 U15795 ( .A1(P1_REG2_REG_13__SCAN_IN), .A2(n13789), .ZN(n13782) );
  NAND2_X1 U15796 ( .A1(n13782), .A2(n13781), .ZN(n13785) );
  MUX2_X1 U15797 ( .A(P1_REG2_REG_14__SCAN_IN), .B(n13783), .S(n13806), .Z(
        n13784) );
  NAND2_X1 U15798 ( .A1(n13784), .A2(n13785), .ZN(n13799) );
  OAI211_X1 U15799 ( .C1(n13785), .C2(n13784), .A(n13866), .B(n13799), .ZN(
        n13796) );
  NAND2_X1 U15800 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n14539)
         );
  INV_X1 U15801 ( .A(n14539), .ZN(n13786) );
  AOI21_X1 U15802 ( .B1(n14604), .B2(P1_ADDR_REG_14__SCAN_IN), .A(n13786), 
        .ZN(n13795) );
  MUX2_X1 U15803 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n13787), .S(n13806), .Z(
        n13791) );
  NAND2_X1 U15804 ( .A1(n13791), .A2(n13790), .ZN(n13807) );
  OAI21_X1 U15805 ( .B1(n13791), .B2(n13790), .A(n13807), .ZN(n13792) );
  NAND2_X1 U15806 ( .A1(n14614), .A2(n13792), .ZN(n13794) );
  NAND2_X1 U15807 ( .A1(n14616), .A2(n13806), .ZN(n13793) );
  NAND4_X1 U15808 ( .A1(n13796), .A2(n13795), .A3(n13794), .A4(n13793), .ZN(
        P1_U3257) );
  INV_X1 U15809 ( .A(n13820), .ZN(n13828) );
  NOR2_X1 U15810 ( .A1(n13862), .A2(n13828), .ZN(n13797) );
  AOI211_X1 U15811 ( .C1(n14604), .C2(P1_ADDR_REG_16__SCAN_IN), .A(n13798), 
        .B(n13797), .ZN(n13816) );
  XNOR2_X1 U15812 ( .A(n13828), .B(P1_REG2_REG_16__SCAN_IN), .ZN(n13805) );
  NAND2_X1 U15813 ( .A1(n13806), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n13800) );
  NAND2_X1 U15814 ( .A1(n13800), .A2(n13799), .ZN(n13801) );
  INV_X1 U15815 ( .A(n13801), .ZN(n13803) );
  INV_X1 U15816 ( .A(n14615), .ZN(n13802) );
  XNOR2_X1 U15817 ( .A(n13801), .B(n14615), .ZN(n14609) );
  NOR2_X1 U15818 ( .A1(P1_REG2_REG_15__SCAN_IN), .A2(n14609), .ZN(n14608) );
  AOI21_X1 U15819 ( .B1(n13803), .B2(n13802), .A(n14608), .ZN(n13804) );
  NAND2_X1 U15820 ( .A1(n13805), .A2(n13804), .ZN(n13826) );
  OAI211_X1 U15821 ( .C1(n13805), .C2(n13804), .A(n13866), .B(n13826), .ZN(
        n13815) );
  OR2_X1 U15822 ( .A1(n13806), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n13808) );
  INV_X1 U15823 ( .A(n13809), .ZN(n13810) );
  XNOR2_X1 U15824 ( .A(n13809), .B(n14615), .ZN(n14612) );
  INV_X1 U15825 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n14611) );
  NAND2_X1 U15826 ( .A1(n14612), .A2(n14611), .ZN(n14610) );
  OAI21_X1 U15827 ( .B1(n13810), .B2(n14615), .A(n14610), .ZN(n13812) );
  XNOR2_X1 U15828 ( .A(n13820), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n13811) );
  AOI211_X1 U15829 ( .C1(n13812), .C2(n13811), .A(n13821), .B(n13847), .ZN(
        n13813) );
  INV_X1 U15830 ( .A(n13813), .ZN(n13814) );
  NAND3_X1 U15831 ( .A1(n13816), .A2(n13815), .A3(n13814), .ZN(P1_U3259) );
  NOR2_X1 U15832 ( .A1(n13862), .A2(n13838), .ZN(n13817) );
  AOI211_X1 U15833 ( .C1(n14604), .C2(P1_ADDR_REG_17__SCAN_IN), .A(n13818), 
        .B(n13817), .ZN(n13836) );
  INV_X1 U15834 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n13819) );
  XNOR2_X1 U15835 ( .A(n13844), .B(n13819), .ZN(n13825) );
  NAND2_X1 U15836 ( .A1(n13820), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n13823) );
  INV_X1 U15837 ( .A(n13821), .ZN(n13822) );
  OAI211_X1 U15838 ( .C1(n13825), .C2(n13824), .A(n14614), .B(n13846), .ZN(
        n13835) );
  OAI21_X1 U15839 ( .B1(n13828), .B2(n13827), .A(n13826), .ZN(n13833) );
  NAND2_X1 U15840 ( .A1(n13844), .A2(n13831), .ZN(n13829) );
  OAI21_X1 U15841 ( .B1(n13844), .B2(n13831), .A(n13829), .ZN(n13832) );
  NAND2_X1 U15842 ( .A1(n13838), .A2(n13831), .ZN(n13830) );
  OAI211_X1 U15843 ( .C1(n13838), .C2(n13831), .A(n13833), .B(n13830), .ZN(
        n13837) );
  OAI211_X1 U15844 ( .C1(n13833), .C2(n13832), .A(n13866), .B(n13837), .ZN(
        n13834) );
  NAND3_X1 U15845 ( .A1(n13836), .A2(n13835), .A3(n13834), .ZN(P1_U3260) );
  OAI21_X1 U15846 ( .B1(n13831), .B2(n13838), .A(n13837), .ZN(n13857) );
  XNOR2_X1 U15847 ( .A(n13857), .B(n13852), .ZN(n13839) );
  NAND2_X1 U15848 ( .A1(P1_REG2_REG_18__SCAN_IN), .A2(n13839), .ZN(n13860) );
  OAI211_X1 U15849 ( .C1(P1_REG2_REG_18__SCAN_IN), .C2(n13839), .A(n13866), 
        .B(n13860), .ZN(n13843) );
  INV_X1 U15850 ( .A(n13840), .ZN(n13841) );
  AOI21_X1 U15851 ( .B1(n14604), .B2(P1_ADDR_REG_18__SCAN_IN), .A(n13841), 
        .ZN(n13842) );
  OAI211_X1 U15852 ( .C1(n13862), .C2(n13852), .A(n13843), .B(n13842), .ZN(
        n13851) );
  NAND2_X1 U15853 ( .A1(n13844), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n13845) );
  AOI211_X1 U15854 ( .C1(n13849), .C2(n13848), .A(n13855), .B(n13847), .ZN(
        n13850) );
  OR2_X1 U15855 ( .A1(n13851), .A2(n13850), .ZN(P1_U3261) );
  INV_X1 U15856 ( .A(n14604), .ZN(n14624) );
  NOR2_X1 U15857 ( .A1(n13853), .A2(n13852), .ZN(n13854) );
  NOR2_X1 U15858 ( .A1(n13855), .A2(n13854), .ZN(n13856) );
  XNOR2_X1 U15859 ( .A(n13856), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n13867) );
  INV_X1 U15860 ( .A(n13867), .ZN(n13864) );
  NAND2_X1 U15861 ( .A1(n13858), .A2(n13857), .ZN(n13859) );
  NAND2_X1 U15862 ( .A1(n13860), .A2(n13859), .ZN(n13861) );
  XOR2_X1 U15863 ( .A(n13861), .B(P1_REG2_REG_19__SCAN_IN), .Z(n13865) );
  OAI21_X1 U15864 ( .B1(n13865), .B2(n14619), .A(n13862), .ZN(n13863) );
  AOI21_X1 U15865 ( .B1(n13864), .B2(n14614), .A(n13863), .ZN(n13870) );
  AOI22_X1 U15866 ( .A1(n13867), .A2(n14614), .B1(n13866), .B2(n13865), .ZN(
        n13869) );
  INV_X1 U15867 ( .A(n13871), .ZN(n13872) );
  INV_X1 U15868 ( .A(n13896), .ZN(n14133) );
  XNOR2_X1 U15869 ( .A(n13882), .B(n13880), .ZN(n13873) );
  NAND2_X1 U15870 ( .A1(n13873), .A2(n14109), .ZN(n14121) );
  NOR2_X1 U15871 ( .A1(n14113), .A2(n13874), .ZN(n13879) );
  NOR2_X1 U15872 ( .A1(n13875), .A2(n15224), .ZN(n13876) );
  NOR2_X1 U15873 ( .A1(n14678), .A2(n13876), .ZN(n13898) );
  INV_X1 U15874 ( .A(n13898), .ZN(n13878) );
  OR2_X1 U15875 ( .A1(n13878), .A2(n13877), .ZN(n14128) );
  NOR2_X1 U15876 ( .A1(n14674), .A2(n14128), .ZN(n13886) );
  AOI211_X1 U15877 ( .C1(n13880), .C2(n14662), .A(n13879), .B(n13886), .ZN(
        n13881) );
  OAI21_X1 U15878 ( .B1(n14121), .B2(n14117), .A(n13881), .ZN(P1_U3263) );
  INV_X1 U15879 ( .A(n13895), .ZN(n13884) );
  INV_X1 U15880 ( .A(n13882), .ZN(n13883) );
  OAI211_X1 U15881 ( .C1(n14130), .C2(n13884), .A(n13883), .B(n14109), .ZN(
        n14129) );
  AND2_X1 U15882 ( .A1(n14674), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n13885) );
  NOR2_X1 U15883 ( .A1(n13886), .A2(n13885), .ZN(n13889) );
  NAND2_X1 U15884 ( .A1(n13887), .A2(n14662), .ZN(n13888) );
  OAI211_X1 U15885 ( .C1(n14129), .C2(n14117), .A(n13889), .B(n13888), .ZN(
        P1_U3264) );
  NAND2_X1 U15886 ( .A1(n14140), .A2(n13913), .ZN(n13892) );
  INV_X1 U15887 ( .A(n13922), .ZN(n13893) );
  AOI21_X1 U15888 ( .B1(n13896), .B2(n13893), .A(n14663), .ZN(n13894) );
  NAND2_X1 U15889 ( .A1(n13896), .A2(n14662), .ZN(n13906) );
  NAND2_X1 U15890 ( .A1(n13913), .A2(n13897), .ZN(n14131) );
  INV_X1 U15891 ( .A(n14131), .ZN(n13903) );
  NAND2_X1 U15892 ( .A1(n13899), .A2(n13898), .ZN(n14132) );
  OAI22_X1 U15893 ( .A1(n13901), .A2(n14132), .B1(n13900), .B2(n14659), .ZN(
        n13902) );
  AOI21_X1 U15894 ( .B1(n14680), .B2(n13903), .A(n13902), .ZN(n13905) );
  NAND2_X1 U15895 ( .A1(n14674), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n13904) );
  NAND3_X1 U15896 ( .A1(n13906), .A2(n13905), .A3(n13904), .ZN(n13907) );
  AOI21_X1 U15897 ( .B1(n14135), .B2(n14669), .A(n13907), .ZN(n13917) );
  XNOR2_X1 U15898 ( .A(n13915), .B(n13914), .ZN(n14136) );
  NAND2_X1 U15899 ( .A1(n14136), .A2(n14675), .ZN(n13916) );
  OAI211_X1 U15900 ( .C1(n6519), .C2(n14095), .A(n13917), .B(n13916), .ZN(
        P1_U3356) );
  AOI211_X1 U15901 ( .C1(n14140), .C2(n6572), .A(n14663), .B(n13922), .ZN(
        n14138) );
  NAND2_X1 U15902 ( .A1(n14138), .A2(n14669), .ZN(n13927) );
  INV_X1 U15903 ( .A(n14139), .ZN(n13924) );
  OAI22_X1 U15904 ( .A1(n14674), .A2(n13924), .B1(n13923), .B2(n14659), .ZN(
        n13925) );
  AOI21_X1 U15905 ( .B1(P1_REG2_REG_28__SCAN_IN), .B2(n14674), .A(n13925), 
        .ZN(n13926) );
  OAI211_X1 U15906 ( .C1(n13911), .C2(n14089), .A(n13927), .B(n13926), .ZN(
        n13928) );
  AOI21_X1 U15907 ( .B1(n14141), .B2(n14676), .A(n13928), .ZN(n13929) );
  OAI21_X1 U15908 ( .B1(n14144), .B2(n14052), .A(n13929), .ZN(P1_U3265) );
  XNOR2_X1 U15909 ( .A(n13930), .B(n13932), .ZN(n14156) );
  XOR2_X1 U15910 ( .A(n13932), .B(n13931), .Z(n14150) );
  NAND2_X1 U15911 ( .A1(n14150), .A2(n14675), .ZN(n13941) );
  AOI211_X1 U15912 ( .C1(n14153), .C2(n13944), .A(n14663), .B(n13933), .ZN(
        n14151) );
  INV_X1 U15913 ( .A(n14152), .ZN(n13935) );
  OAI22_X1 U15914 ( .A1(n14674), .A2(n13935), .B1(n13934), .B2(n14659), .ZN(
        n13936) );
  AOI21_X1 U15915 ( .B1(P1_REG2_REG_26__SCAN_IN), .B2(n14674), .A(n13936), 
        .ZN(n13937) );
  OAI21_X1 U15916 ( .B1(n13938), .B2(n14089), .A(n13937), .ZN(n13939) );
  AOI21_X1 U15917 ( .B1(n14151), .B2(n14669), .A(n13939), .ZN(n13940) );
  OAI211_X1 U15918 ( .C1(n14156), .C2(n14095), .A(n13941), .B(n13940), .ZN(
        P1_U3267) );
  OAI21_X1 U15919 ( .B1(n13943), .B2(n13952), .A(n13942), .ZN(n14163) );
  INV_X1 U15920 ( .A(n13962), .ZN(n13945) );
  AOI211_X1 U15921 ( .C1(n14159), .C2(n13945), .A(n14663), .B(n7265), .ZN(
        n14157) );
  INV_X1 U15922 ( .A(n14158), .ZN(n13947) );
  OAI22_X1 U15923 ( .A1(n14674), .A2(n13947), .B1(n13946), .B2(n14659), .ZN(
        n13948) );
  AOI21_X1 U15924 ( .B1(P1_REG2_REG_25__SCAN_IN), .B2(n14674), .A(n13948), 
        .ZN(n13949) );
  OAI21_X1 U15925 ( .B1(n13950), .B2(n14089), .A(n13949), .ZN(n13951) );
  AOI21_X1 U15926 ( .B1(n14157), .B2(n14669), .A(n13951), .ZN(n13955) );
  XNOR2_X1 U15927 ( .A(n13953), .B(n13952), .ZN(n14160) );
  NAND2_X1 U15928 ( .A1(n14160), .A2(n14675), .ZN(n13954) );
  OAI211_X1 U15929 ( .C1(n14163), .C2(n14095), .A(n13955), .B(n13954), .ZN(
        P1_U3268) );
  INV_X1 U15930 ( .A(n13956), .ZN(n13958) );
  AOI21_X1 U15931 ( .B1(n13958), .B2(n13957), .A(n14737), .ZN(n13961) );
  AOI21_X1 U15932 ( .B1(n13961), .B2(n6765), .A(n13959), .ZN(n14167) );
  AOI211_X1 U15933 ( .C1(n14165), .C2(n6593), .A(n14663), .B(n13962), .ZN(
        n14164) );
  NOR2_X1 U15934 ( .A1(n13963), .A2(n14089), .ZN(n13967) );
  OAI22_X1 U15935 ( .A1(n14113), .A2(n13965), .B1(n13964), .B2(n14659), .ZN(
        n13966) );
  AOI211_X1 U15936 ( .C1(n14164), .C2(n14669), .A(n13967), .B(n13966), .ZN(
        n13973) );
  AOI21_X1 U15937 ( .B1(n13969), .B2(n13968), .A(n6620), .ZN(n14168) );
  INV_X1 U15938 ( .A(n14168), .ZN(n13971) );
  NAND2_X1 U15939 ( .A1(n13971), .A2(n13970), .ZN(n13972) );
  OAI211_X1 U15940 ( .C1(n14167), .C2(n14674), .A(n13973), .B(n13972), .ZN(
        P1_U3269) );
  XOR2_X1 U15941 ( .A(n13974), .B(n13976), .Z(n14175) );
  XOR2_X1 U15942 ( .A(n13975), .B(n13976), .Z(n14173) );
  OAI211_X1 U15943 ( .C1(n14171), .C2(n6516), .A(n14109), .B(n6593), .ZN(
        n14170) );
  NOR2_X1 U15944 ( .A1(n14113), .A2(n13977), .ZN(n13980) );
  OAI22_X1 U15945 ( .A1(n14169), .A2(n14674), .B1(n13978), .B2(n14659), .ZN(
        n13979) );
  AOI211_X1 U15946 ( .C1(n13981), .C2(n14662), .A(n13980), .B(n13979), .ZN(
        n13982) );
  OAI21_X1 U15947 ( .B1(n14170), .B2(n14117), .A(n13982), .ZN(n13983) );
  AOI21_X1 U15948 ( .B1(n14173), .B2(n14676), .A(n13983), .ZN(n13984) );
  OAI21_X1 U15949 ( .B1(n14175), .B2(n14052), .A(n13984), .ZN(P1_U3270) );
  XOR2_X1 U15950 ( .A(n13985), .B(n13988), .Z(n14179) );
  OAI21_X1 U15951 ( .B1(n13988), .B2(n13987), .A(n13986), .ZN(n13991) );
  INV_X1 U15952 ( .A(n13989), .ZN(n13990) );
  AOI21_X1 U15953 ( .B1(n13991), .B2(n14694), .A(n13990), .ZN(n14178) );
  INV_X1 U15954 ( .A(n14178), .ZN(n13999) );
  AOI21_X1 U15955 ( .B1(n12276), .B2(n14010), .A(n14663), .ZN(n13993) );
  AND2_X1 U15956 ( .A1(n13993), .A2(n13992), .ZN(n14176) );
  NAND2_X1 U15957 ( .A1(n14176), .A2(n14669), .ZN(n13996) );
  AOI22_X1 U15958 ( .A1(n14674), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n13994), 
        .B2(n14673), .ZN(n13995) );
  OAI211_X1 U15959 ( .C1(n14089), .C2(n13997), .A(n13996), .B(n13995), .ZN(
        n13998) );
  AOI21_X1 U15960 ( .B1(n13999), .B2(n14113), .A(n13998), .ZN(n14000) );
  OAI21_X1 U15961 ( .B1(n14179), .B2(n14095), .A(n14000), .ZN(P1_U3271) );
  OAI21_X1 U15962 ( .B1(n14001), .B2(n14006), .A(n14694), .ZN(n14002) );
  OR2_X1 U15963 ( .A1(n14003), .A2(n14002), .ZN(n14005) );
  NAND2_X1 U15964 ( .A1(n14005), .A2(n14004), .ZN(n14185) );
  INV_X1 U15965 ( .A(n14185), .ZN(n14018) );
  AND2_X1 U15966 ( .A1(n14007), .A2(n14006), .ZN(n14008) );
  OR2_X1 U15967 ( .A1(n14009), .A2(n14008), .ZN(n14180) );
  AOI21_X1 U15968 ( .B1(n14026), .B2(n14013), .A(n14663), .ZN(n14011) );
  NAND2_X1 U15969 ( .A1(n14011), .A2(n14010), .ZN(n14181) );
  AOI22_X1 U15970 ( .A1(n14674), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n14012), 
        .B2(n14673), .ZN(n14015) );
  NAND2_X1 U15971 ( .A1(n14013), .A2(n14662), .ZN(n14014) );
  OAI211_X1 U15972 ( .C1(n14181), .C2(n14117), .A(n14015), .B(n14014), .ZN(
        n14016) );
  AOI21_X1 U15973 ( .B1(n14180), .B2(n14676), .A(n14016), .ZN(n14017) );
  OAI21_X1 U15974 ( .B1(n14018), .B2(n14674), .A(n14017), .ZN(P1_U3272) );
  AND2_X1 U15975 ( .A1(n14035), .A2(n14019), .ZN(n14021) );
  OAI211_X1 U15976 ( .C1(n14021), .C2(n14030), .A(n14020), .B(n14694), .ZN(
        n14023) );
  NAND2_X1 U15977 ( .A1(n14023), .A2(n14022), .ZN(n14194) );
  INV_X1 U15978 ( .A(n14194), .ZN(n14034) );
  INV_X1 U15979 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n14025) );
  OAI22_X1 U15980 ( .A1(n14113), .A2(n14025), .B1(n14024), .B2(n14659), .ZN(
        n14028) );
  OAI211_X1 U15981 ( .C1(n14192), .C2(n14040), .A(n14109), .B(n14026), .ZN(
        n14190) );
  NOR2_X1 U15982 ( .A1(n14190), .A2(n14117), .ZN(n14027) );
  AOI211_X1 U15983 ( .C1(n14662), .C2(n14029), .A(n14028), .B(n14027), .ZN(
        n14033) );
  NAND2_X1 U15984 ( .A1(n14031), .A2(n14030), .ZN(n14188) );
  NAND3_X1 U15985 ( .A1(n14189), .A2(n14188), .A3(n14676), .ZN(n14032) );
  OAI211_X1 U15986 ( .C1(n14034), .C2(n14674), .A(n14033), .B(n14032), .ZN(
        P1_U3273) );
  INV_X1 U15987 ( .A(n14035), .ZN(n14036) );
  AOI21_X1 U15988 ( .B1(n14048), .B2(n14037), .A(n14036), .ZN(n14201) );
  NAND2_X1 U15989 ( .A1(n14197), .A2(n14058), .ZN(n14038) );
  NAND2_X1 U15990 ( .A1(n14038), .A2(n14109), .ZN(n14039) );
  NOR2_X1 U15991 ( .A1(n14040), .A2(n14039), .ZN(n14195) );
  INV_X1 U15992 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n14046) );
  NAND2_X1 U15993 ( .A1(n14197), .A2(n14662), .ZN(n14045) );
  INV_X1 U15994 ( .A(n14196), .ZN(n14042) );
  OAI22_X1 U15995 ( .A1(n14674), .A2(n14042), .B1(n14041), .B2(n14659), .ZN(
        n14043) );
  INV_X1 U15996 ( .A(n14043), .ZN(n14044) );
  OAI211_X1 U15997 ( .C1(n14113), .C2(n14046), .A(n14045), .B(n14044), .ZN(
        n14047) );
  AOI21_X1 U15998 ( .B1(n14195), .B2(n14669), .A(n14047), .ZN(n14051) );
  XNOR2_X1 U15999 ( .A(n14049), .B(n14048), .ZN(n14198) );
  NAND2_X1 U16000 ( .A1(n14198), .A2(n14676), .ZN(n14050) );
  OAI211_X1 U16001 ( .C1(n14201), .C2(n14052), .A(n14051), .B(n14050), .ZN(
        P1_U3274) );
  XNOR2_X1 U16002 ( .A(n14054), .B(n14053), .ZN(n14207) );
  OAI211_X1 U16003 ( .C1(n6684), .C2(n14056), .A(n14694), .B(n14055), .ZN(
        n14206) );
  INV_X1 U16004 ( .A(n14206), .ZN(n14057) );
  OAI21_X1 U16005 ( .B1(n14057), .B2(n14203), .A(n14113), .ZN(n14065) );
  INV_X1 U16006 ( .A(n14058), .ZN(n14059) );
  AOI211_X1 U16007 ( .C1(n14204), .C2(n14070), .A(n14663), .B(n14059), .ZN(
        n14202) );
  NOR2_X1 U16008 ( .A1(n7269), .A2(n14089), .ZN(n14063) );
  OAI22_X1 U16009 ( .A1(n14113), .A2(n14061), .B1(n14060), .B2(n14659), .ZN(
        n14062) );
  AOI211_X1 U16010 ( .C1(n14202), .C2(n14669), .A(n14063), .B(n14062), .ZN(
        n14064) );
  OAI211_X1 U16011 ( .C1(n14066), .C2(n14207), .A(n14065), .B(n14064), .ZN(
        P1_U3275) );
  XNOR2_X1 U16012 ( .A(n14067), .B(n14075), .ZN(n14069) );
  AOI21_X1 U16013 ( .B1(n14069), .B2(n14694), .A(n14068), .ZN(n14211) );
  AOI211_X1 U16014 ( .C1(n14209), .C2(n14086), .A(n14663), .B(n7270), .ZN(
        n14208) );
  INV_X1 U16015 ( .A(n14071), .ZN(n14072) );
  AOI22_X1 U16016 ( .A1(n14674), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n14072), 
        .B2(n14673), .ZN(n14073) );
  OAI21_X1 U16017 ( .B1(n14074), .B2(n14089), .A(n14073), .ZN(n14078) );
  XNOR2_X1 U16018 ( .A(n6750), .B(n14075), .ZN(n14212) );
  NOR2_X1 U16019 ( .A1(n14212), .A2(n14095), .ZN(n14077) );
  AOI211_X1 U16020 ( .C1(n14208), .C2(n14669), .A(n14078), .B(n14077), .ZN(
        n14079) );
  OAI21_X1 U16021 ( .B1(n14674), .B2(n14211), .A(n14079), .ZN(P1_U3276) );
  XNOR2_X1 U16022 ( .A(n14080), .B(n14085), .ZN(n14219) );
  NAND2_X1 U16023 ( .A1(n14097), .A2(n14081), .ZN(n14083) );
  OAI21_X1 U16024 ( .B1(n6680), .B2(n14085), .A(n14084), .ZN(n14217) );
  OAI211_X1 U16025 ( .C1(n14108), .C2(n14215), .A(n14086), .B(n14109), .ZN(
        n14214) );
  INV_X1 U16026 ( .A(n14087), .ZN(n14213) );
  OAI22_X1 U16027 ( .A1(n14674), .A2(n14213), .B1(n14088), .B2(n14659), .ZN(
        n14091) );
  NOR2_X1 U16028 ( .A1(n14215), .A2(n14089), .ZN(n14090) );
  AOI211_X1 U16029 ( .C1(n14674), .C2(P1_REG2_REG_16__SCAN_IN), .A(n14091), 
        .B(n14090), .ZN(n14092) );
  OAI21_X1 U16030 ( .B1(n14117), .B2(n14214), .A(n14092), .ZN(n14093) );
  AOI21_X1 U16031 ( .B1(n14217), .B2(n14675), .A(n14093), .ZN(n14094) );
  OAI21_X1 U16032 ( .B1(n14095), .B2(n14219), .A(n14094), .ZN(P1_U3277) );
  NAND2_X1 U16033 ( .A1(n14097), .A2(n14096), .ZN(n14099) );
  XNOR2_X1 U16034 ( .A(n14099), .B(n14098), .ZN(n14102) );
  INV_X1 U16035 ( .A(n14100), .ZN(n14101) );
  OAI21_X1 U16036 ( .B1(n14102), .B2(n14737), .A(n14101), .ZN(n14545) );
  INV_X1 U16037 ( .A(n14545), .ZN(n14120) );
  INV_X1 U16038 ( .A(n14103), .ZN(n14106) );
  OAI21_X1 U16039 ( .B1(n14106), .B2(n14105), .A(n14104), .ZN(n14547) );
  INV_X1 U16040 ( .A(n14108), .ZN(n14110) );
  OAI211_X1 U16041 ( .C1(n14544), .C2(n7264), .A(n14110), .B(n14109), .ZN(
        n14543) );
  OAI22_X1 U16042 ( .A1(n14113), .A2(n14112), .B1(n14111), .B2(n14659), .ZN(
        n14114) );
  AOI21_X1 U16043 ( .B1(n14115), .B2(n14662), .A(n14114), .ZN(n14116) );
  OAI21_X1 U16044 ( .B1(n14543), .B2(n14117), .A(n14116), .ZN(n14118) );
  AOI21_X1 U16045 ( .B1(n14547), .B2(n14676), .A(n14118), .ZN(n14119) );
  OAI21_X1 U16046 ( .B1(n14120), .B2(n14674), .A(n14119), .ZN(P1_U3278) );
  OAI211_X1 U16047 ( .C1(n14122), .C2(n14767), .A(n14121), .B(n14128), .ZN(
        n14224) );
  INV_X1 U16048 ( .A(n14123), .ZN(n14125) );
  MUX2_X1 U16049 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n14224), .S(n14788), .Z(
        P1_U3559) );
  OAI211_X1 U16050 ( .C1(n14130), .C2(n14767), .A(n14129), .B(n14128), .ZN(
        n14225) );
  MUX2_X1 U16051 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n14225), .S(n14788), .Z(
        P1_U3558) );
  OAI211_X1 U16052 ( .C1(n14133), .C2(n14767), .A(n14132), .B(n14131), .ZN(
        n14134) );
  MUX2_X1 U16053 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n14226), .S(n14788), .Z(
        P1_U3557) );
  AOI211_X1 U16054 ( .C1(n14140), .C2(n14742), .A(n14139), .B(n14138), .ZN(
        n14143) );
  NAND2_X1 U16055 ( .A1(n14141), .A2(n14771), .ZN(n14142) );
  INV_X1 U16056 ( .A(n14747), .ZN(n14763) );
  NAND2_X1 U16057 ( .A1(n14145), .A2(n14763), .ZN(n14147) );
  MUX2_X1 U16058 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n14228), .S(n14788), .Z(
        P1_U3555) );
  NAND2_X1 U16059 ( .A1(n14150), .A2(n14694), .ZN(n14155) );
  AOI211_X1 U16060 ( .C1(n14153), .C2(n14742), .A(n14152), .B(n14151), .ZN(
        n14154) );
  OAI211_X1 U16061 ( .C1(n14724), .C2(n14156), .A(n14155), .B(n14154), .ZN(
        n14229) );
  MUX2_X1 U16062 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n14229), .S(n14788), .Z(
        P1_U3554) );
  AOI211_X1 U16063 ( .C1(n14159), .C2(n14742), .A(n14158), .B(n14157), .ZN(
        n14162) );
  NAND2_X1 U16064 ( .A1(n14160), .A2(n14694), .ZN(n14161) );
  OAI211_X1 U16065 ( .C1(n14163), .C2(n14724), .A(n14162), .B(n14161), .ZN(
        n14230) );
  MUX2_X1 U16066 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n14230), .S(n14788), .Z(
        P1_U3553) );
  AOI21_X1 U16067 ( .B1(n14165), .B2(n14742), .A(n14164), .ZN(n14166) );
  OAI211_X1 U16068 ( .C1(n14724), .C2(n14168), .A(n14167), .B(n14166), .ZN(
        n14231) );
  MUX2_X1 U16069 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n14231), .S(n14788), .Z(
        P1_U3552) );
  OAI211_X1 U16070 ( .C1(n14171), .C2(n14767), .A(n14170), .B(n14169), .ZN(
        n14172) );
  AOI21_X1 U16071 ( .B1(n14173), .B2(n14771), .A(n14172), .ZN(n14174) );
  OAI21_X1 U16072 ( .B1(n14175), .B2(n14737), .A(n14174), .ZN(n14232) );
  MUX2_X1 U16073 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n14232), .S(n14788), .Z(
        P1_U3551) );
  AOI21_X1 U16074 ( .B1(n12276), .B2(n14742), .A(n14176), .ZN(n14177) );
  OAI211_X1 U16075 ( .C1(n14724), .C2(n14179), .A(n14178), .B(n14177), .ZN(
        n14233) );
  MUX2_X1 U16076 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n14233), .S(n14788), .Z(
        P1_U3550) );
  NAND2_X1 U16077 ( .A1(n14180), .A2(n14771), .ZN(n14182) );
  OAI211_X1 U16078 ( .C1(n14183), .C2(n14767), .A(n14182), .B(n14181), .ZN(
        n14184) );
  NOR2_X1 U16079 ( .A1(n14185), .A2(n14184), .ZN(n14235) );
  INV_X1 U16080 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n14186) );
  MUX2_X1 U16081 ( .A(n14235), .B(n14186), .S(n14786), .Z(n14187) );
  INV_X1 U16082 ( .A(n14187), .ZN(P1_U3549) );
  NAND3_X1 U16083 ( .A1(n14189), .A2(n14771), .A3(n14188), .ZN(n14191) );
  OAI211_X1 U16084 ( .C1(n14192), .C2(n14767), .A(n14191), .B(n14190), .ZN(
        n14193) );
  MUX2_X1 U16085 ( .A(n14237), .B(P1_REG1_REG_20__SCAN_IN), .S(n14786), .Z(
        P1_U3548) );
  AOI211_X1 U16086 ( .C1(n14197), .C2(n14742), .A(n14196), .B(n14195), .ZN(
        n14200) );
  NAND2_X1 U16087 ( .A1(n14198), .A2(n14771), .ZN(n14199) );
  OAI211_X1 U16088 ( .C1(n14201), .C2(n14737), .A(n14200), .B(n14199), .ZN(
        n14238) );
  MUX2_X1 U16089 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n14238), .S(n14788), .Z(
        P1_U3547) );
  AOI211_X1 U16090 ( .C1(n14204), .C2(n14742), .A(n14203), .B(n14202), .ZN(
        n14205) );
  OAI211_X1 U16091 ( .C1(n14724), .C2(n14207), .A(n14206), .B(n14205), .ZN(
        n14239) );
  MUX2_X1 U16092 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n14239), .S(n14788), .Z(
        P1_U3546) );
  AOI21_X1 U16093 ( .B1(n14209), .B2(n14742), .A(n14208), .ZN(n14210) );
  OAI211_X1 U16094 ( .C1(n14724), .C2(n14212), .A(n14211), .B(n14210), .ZN(
        n14240) );
  MUX2_X1 U16095 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n14240), .S(n14788), .Z(
        P1_U3545) );
  OAI211_X1 U16096 ( .C1(n14215), .C2(n14767), .A(n14214), .B(n14213), .ZN(
        n14216) );
  AOI21_X1 U16097 ( .B1(n14217), .B2(n14694), .A(n14216), .ZN(n14218) );
  OAI21_X1 U16098 ( .B1(n14724), .B2(n14219), .A(n14218), .ZN(n14241) );
  MUX2_X1 U16099 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n14241), .S(n14788), .Z(
        P1_U3544) );
  NOR2_X1 U16100 ( .A1(n14221), .A2(n14220), .ZN(n14222) );
  MUX2_X1 U16101 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n14224), .S(n14774), .Z(
        P1_U3527) );
  MUX2_X1 U16102 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n14225), .S(n14774), .Z(
        P1_U3526) );
  MUX2_X1 U16103 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n14226), .S(n14774), .Z(
        P1_U3525) );
  MUX2_X1 U16104 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n14229), .S(n14774), .Z(
        P1_U3522) );
  MUX2_X1 U16105 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n14230), .S(n14774), .Z(
        P1_U3521) );
  MUX2_X1 U16106 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n14231), .S(n14774), .Z(
        P1_U3520) );
  MUX2_X1 U16107 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n14232), .S(n14774), .Z(
        P1_U3519) );
  MUX2_X1 U16108 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n14233), .S(n14774), .Z(
        P1_U3518) );
  INV_X1 U16109 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n14234) );
  MUX2_X1 U16110 ( .A(n14235), .B(n14234), .S(n14772), .Z(n14236) );
  INV_X1 U16111 ( .A(n14236), .ZN(P1_U3517) );
  MUX2_X1 U16112 ( .A(n14237), .B(P1_REG0_REG_20__SCAN_IN), .S(n14772), .Z(
        P1_U3516) );
  MUX2_X1 U16113 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n14238), .S(n14774), .Z(
        P1_U3515) );
  MUX2_X1 U16114 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n14239), .S(n14774), .Z(
        P1_U3513) );
  MUX2_X1 U16115 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n14240), .S(n14774), .Z(
        P1_U3510) );
  MUX2_X1 U16116 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n14241), .S(n14774), .Z(
        P1_U3507) );
  NOR4_X1 U16117 ( .A1(n14242), .A2(P1_IR_REG_30__SCAN_IN), .A3(n9318), .A4(
        P1_U3086), .ZN(n14243) );
  AOI21_X1 U16118 ( .B1(n14244), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n14243), 
        .ZN(n14245) );
  OAI21_X1 U16119 ( .B1(n14246), .B2(n11860), .A(n14245), .ZN(P1_U3324) );
  OAI222_X1 U16120 ( .A1(P1_U3086), .A2(n14249), .B1(n11860), .B2(n14248), 
        .C1(n15197), .C2(n14247), .ZN(P1_U3329) );
  MUX2_X1 U16121 ( .A(n6796), .B(n14250), .S(P1_U3086), .Z(P1_U3333) );
  INV_X1 U16122 ( .A(n14252), .ZN(n14253) );
  MUX2_X1 U16123 ( .A(n14253), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  INV_X1 U16124 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n14598) );
  INV_X1 U16125 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n14625) );
  NOR2_X1 U16126 ( .A1(P3_ADDR_REG_15__SCAN_IN), .A2(n14625), .ZN(n14283) );
  INV_X1 U16127 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n14281) );
  XNOR2_X1 U16128 ( .A(P3_ADDR_REG_14__SCAN_IN), .B(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n14333) );
  INV_X1 U16129 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n14279) );
  INV_X1 U16130 ( .A(P3_ADDR_REG_12__SCAN_IN), .ZN(n14276) );
  XNOR2_X1 U16131 ( .A(P3_ADDR_REG_12__SCAN_IN), .B(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n14329) );
  INV_X1 U16132 ( .A(P3_ADDR_REG_11__SCAN_IN), .ZN(n14274) );
  INV_X1 U16133 ( .A(P3_ADDR_REG_10__SCAN_IN), .ZN(n15030) );
  XNOR2_X1 U16134 ( .A(n15030), .B(P1_ADDR_REG_10__SCAN_IN), .ZN(n14288) );
  INV_X1 U16135 ( .A(P3_ADDR_REG_9__SCAN_IN), .ZN(n14271) );
  INV_X1 U16136 ( .A(P3_ADDR_REG_8__SCAN_IN), .ZN(n14269) );
  INV_X1 U16137 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n14255) );
  NOR2_X1 U16138 ( .A1(n14257), .A2(n14258), .ZN(n14260) );
  NOR2_X1 U16139 ( .A1(n14261), .A2(n14974), .ZN(n14263) );
  INV_X1 U16140 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n15146) );
  NOR2_X1 U16141 ( .A1(P3_ADDR_REG_6__SCAN_IN), .A2(n15146), .ZN(n14308) );
  NOR2_X1 U16142 ( .A1(P3_ADDR_REG_7__SCAN_IN), .A2(n14264), .ZN(n14267) );
  INV_X1 U16143 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n14265) );
  XOR2_X1 U16144 ( .A(P3_ADDR_REG_8__SCAN_IN), .B(P1_ADDR_REG_8__SCAN_IN), .Z(
        n14289) );
  XNOR2_X1 U16145 ( .A(P3_ADDR_REG_9__SCAN_IN), .B(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n14320) );
  NAND2_X1 U16146 ( .A1(n14321), .A2(n14320), .ZN(n14270) );
  XNOR2_X1 U16147 ( .A(P3_ADDR_REG_11__SCAN_IN), .B(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n14326) );
  NAND2_X1 U16148 ( .A1(n14327), .A2(n14326), .ZN(n14273) );
  NAND2_X1 U16149 ( .A1(n14329), .A2(n14330), .ZN(n14275) );
  INV_X1 U16150 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n14277) );
  NAND2_X1 U16151 ( .A1(P1_ADDR_REG_13__SCAN_IN), .A2(n14277), .ZN(n14278) );
  NAND2_X1 U16152 ( .A1(n14333), .A2(n14332), .ZN(n14280) );
  INV_X1 U16153 ( .A(P3_ADDR_REG_15__SCAN_IN), .ZN(n14282) );
  OAI22_X1 U16154 ( .A1(n14283), .A2(n14336), .B1(P1_ADDR_REG_15__SCAN_IN), 
        .B2(n14282), .ZN(n14339) );
  XOR2_X1 U16155 ( .A(P1_ADDR_REG_16__SCAN_IN), .B(P3_ADDR_REG_16__SCAN_IN), 
        .Z(n14284) );
  XOR2_X1 U16156 ( .A(n14339), .B(n14284), .Z(n14597) );
  XOR2_X1 U16157 ( .A(P3_ADDR_REG_13__SCAN_IN), .B(P1_ADDR_REG_13__SCAN_IN), 
        .Z(n14285) );
  XOR2_X1 U16158 ( .A(n14286), .B(n14285), .Z(n14584) );
  INV_X1 U16159 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n14859) );
  INV_X1 U16160 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n14842) );
  XOR2_X1 U16161 ( .A(n14288), .B(n14287), .Z(n14389) );
  XOR2_X1 U16162 ( .A(n14290), .B(n14289), .Z(n14317) );
  NAND2_X1 U16163 ( .A1(P2_ADDR_REG_4__SCAN_IN), .A2(n14292), .ZN(n14303) );
  INV_X1 U16164 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n15434) );
  NAND2_X1 U16165 ( .A1(P2_ADDR_REG_1__SCAN_IN), .A2(n14295), .ZN(n14296) );
  AOI21_X1 U16166 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(n14938), .A(n14294), .ZN(
        n15428) );
  NOR2_X1 U16167 ( .A1(n15428), .A2(n9569), .ZN(n15437) );
  XNOR2_X1 U16168 ( .A(n14298), .B(n14297), .ZN(n14349) );
  NOR2_X1 U16169 ( .A1(n14350), .A2(n14349), .ZN(n14300) );
  INV_X1 U16170 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n14299) );
  NAND2_X1 U16171 ( .A1(n14350), .A2(n14349), .ZN(n14348) );
  XNOR2_X1 U16172 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(n14301), .ZN(n15433) );
  NAND2_X1 U16173 ( .A1(n15432), .A2(n15433), .ZN(n14302) );
  NOR2_X1 U16174 ( .A1(n15432), .A2(n15433), .ZN(n15431) );
  AOI21_X1 U16175 ( .B1(n15434), .B2(n14302), .A(n15431), .ZN(n15425) );
  XNOR2_X1 U16176 ( .A(n14306), .B(n14305), .ZN(n15427) );
  NAND2_X1 U16177 ( .A1(n14307), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n14311) );
  INV_X1 U16178 ( .A(n14308), .ZN(n15361) );
  OAI21_X1 U16179 ( .B1(n15223), .B2(P1_ADDR_REG_6__SCAN_IN), .A(n15361), .ZN(
        n14310) );
  XNOR2_X1 U16180 ( .A(n14310), .B(n14309), .ZN(n14375) );
  NAND2_X1 U16181 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n14312), .ZN(n14315) );
  XNOR2_X1 U16182 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n14313), .ZN(n15429) );
  NAND2_X1 U16183 ( .A1(n15430), .A2(n15429), .ZN(n14314) );
  NOR2_X1 U16184 ( .A1(n14317), .A2(n14316), .ZN(n14319) );
  XNOR2_X1 U16185 ( .A(n14321), .B(n14320), .ZN(n14323) );
  NAND2_X1 U16186 ( .A1(n14322), .A2(n14323), .ZN(n14324) );
  NAND2_X1 U16187 ( .A1(n14389), .A2(n14388), .ZN(n14325) );
  XNOR2_X1 U16188 ( .A(n14327), .B(n14326), .ZN(n14576) );
  NAND2_X1 U16189 ( .A1(n14577), .A2(n14576), .ZN(n14328) );
  NOR2_X1 U16190 ( .A1(n14577), .A2(n14576), .ZN(n14575) );
  XNOR2_X1 U16191 ( .A(n14330), .B(n14329), .ZN(n14580) );
  NAND2_X1 U16192 ( .A1(n14584), .A2(n14585), .ZN(n14331) );
  AOI21_X2 U16193 ( .B1(n11036), .B2(n14331), .A(n14583), .ZN(n14589) );
  XOR2_X1 U16194 ( .A(n14333), .B(n14332), .Z(n14588) );
  INV_X1 U16195 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n14334) );
  NAND2_X1 U16196 ( .A1(n14589), .A2(n14588), .ZN(n14587) );
  XNOR2_X1 U16197 ( .A(P1_ADDR_REG_15__SCAN_IN), .B(P3_ADDR_REG_15__SCAN_IN), 
        .ZN(n14337) );
  XOR2_X1 U16198 ( .A(n14337), .B(n14336), .Z(n14592) );
  INV_X1 U16199 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n15410) );
  NAND2_X1 U16200 ( .A1(n14593), .A2(n14592), .ZN(n14591) );
  INV_X1 U16201 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n14341) );
  NOR2_X1 U16202 ( .A1(P1_ADDR_REG_16__SCAN_IN), .A2(n14338), .ZN(n14340) );
  OAI22_X1 U16203 ( .A1(P3_ADDR_REG_16__SCAN_IN), .A2(n14341), .B1(n14340), 
        .B2(n14339), .ZN(n14342) );
  XOR2_X1 U16204 ( .A(P1_ADDR_REG_17__SCAN_IN), .B(n14342), .Z(n14343) );
  XNOR2_X1 U16205 ( .A(P3_ADDR_REG_17__SCAN_IN), .B(n14343), .ZN(n14401) );
  NOR2_X1 U16206 ( .A1(P1_ADDR_REG_17__SCAN_IN), .A2(n14342), .ZN(n14345) );
  AND2_X1 U16207 ( .A1(P3_ADDR_REG_17__SCAN_IN), .A2(n14343), .ZN(n14344) );
  NOR2_X1 U16208 ( .A1(n14345), .A2(n14344), .ZN(n14409) );
  XOR2_X1 U16209 ( .A(P3_ADDR_REG_18__SCAN_IN), .B(P1_ADDR_REG_18__SCAN_IN), 
        .Z(n14408) );
  XNOR2_X1 U16210 ( .A(n14409), .B(n14408), .ZN(n14404) );
  XNOR2_X1 U16211 ( .A(P2_ADDR_REG_18__SCAN_IN), .B(n14403), .ZN(SUB_1596_U62)
         );
  AOI21_X1 U16212 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n14346) );
  OAI21_X1 U16213 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(n14346), 
        .ZN(U28) );
  AOI21_X1 U16214 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(
        P3_RD_REG_SCAN_IN), .ZN(n14347) );
  OAI21_X1 U16215 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(n14347), 
        .ZN(U29) );
  OAI21_X1 U16216 ( .B1(n14350), .B2(n14349), .A(n14348), .ZN(n14351) );
  XNOR2_X1 U16217 ( .A(n14351), .B(P2_ADDR_REG_2__SCAN_IN), .ZN(SUB_1596_U61)
         );
  AOI22_X1 U16218 ( .A1(n14352), .A2(n14381), .B1(SI_6_), .B2(n14380), .ZN(
        n14353) );
  OAI21_X1 U16219 ( .B1(P3_U3151), .B2(n14354), .A(n14353), .ZN(P3_U3289) );
  INV_X1 U16220 ( .A(n14355), .ZN(n14356) );
  AOI22_X1 U16221 ( .A1(n14356), .A2(n14381), .B1(SI_4_), .B2(n14380), .ZN(
        n14357) );
  OAI21_X1 U16222 ( .B1(P3_U3151), .B2(n14358), .A(n14357), .ZN(P3_U3291) );
  INV_X1 U16223 ( .A(n14359), .ZN(n14360) );
  AOI22_X1 U16224 ( .A1(n14360), .A2(n14381), .B1(SI_2_), .B2(n14380), .ZN(
        n14361) );
  OAI21_X1 U16225 ( .B1(P3_U3151), .B2(n14362), .A(n14361), .ZN(P3_U3293) );
  NOR2_X1 U16226 ( .A1(n14368), .A2(n14363), .ZN(n14364) );
  AOI21_X1 U16227 ( .B1(n14365), .B2(n14381), .A(n14364), .ZN(n14366) );
  OAI21_X1 U16228 ( .B1(P3_U3151), .B2(n14367), .A(n14366), .ZN(P3_U3287) );
  OAI22_X1 U16229 ( .A1(n14371), .A2(n14370), .B1(n14369), .B2(n14368), .ZN(
        n14372) );
  INV_X1 U16230 ( .A(n14372), .ZN(n14373) );
  OAI21_X1 U16231 ( .B1(P3_U3151), .B2(n14374), .A(n14373), .ZN(P3_U3285) );
  XOR2_X1 U16232 ( .A(n14376), .B(n14375), .Z(SUB_1596_U57) );
  AOI22_X1 U16233 ( .A1(n14377), .A2(n14381), .B1(SI_14_), .B2(n14380), .ZN(
        n14378) );
  OAI21_X1 U16234 ( .B1(P3_U3151), .B2(n14379), .A(n14378), .ZN(P3_U3281) );
  AOI22_X1 U16235 ( .A1(n14382), .A2(n14381), .B1(SI_16_), .B2(n14380), .ZN(
        n14383) );
  OAI21_X1 U16236 ( .B1(P3_U3151), .B2(n14384), .A(n14383), .ZN(P3_U3279) );
  XNOR2_X1 U16237 ( .A(n6522), .B(P2_ADDR_REG_8__SCAN_IN), .ZN(SUB_1596_U55)
         );
  XNOR2_X1 U16238 ( .A(n14386), .B(n15353), .ZN(SUB_1596_U54) );
  AOI21_X1 U16239 ( .B1(n14389), .B2(n14388), .A(n14387), .ZN(n14390) );
  XNOR2_X1 U16240 ( .A(n14390), .B(n10173), .ZN(SUB_1596_U70) );
  INV_X1 U16241 ( .A(n14391), .ZN(n14396) );
  OAI21_X1 U16242 ( .B1(n14393), .B2(n14767), .A(n14392), .ZN(n14395) );
  AOI211_X1 U16243 ( .C1(n14763), .C2(n14396), .A(n14395), .B(n14394), .ZN(
        n14398) );
  INV_X1 U16244 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n14397) );
  AOI22_X1 U16245 ( .A1(n14774), .A2(n14398), .B1(n14397), .B2(n14772), .ZN(
        P1_U3495) );
  AOI22_X1 U16246 ( .A1(n14788), .A2(n14398), .B1(n15368), .B2(n14786), .ZN(
        P1_U3540) );
  OAI21_X1 U16247 ( .B1(n14401), .B2(n14400), .A(n14399), .ZN(n14402) );
  XNOR2_X1 U16248 ( .A(n14402), .B(P2_ADDR_REG_17__SCAN_IN), .ZN(SUB_1596_U63)
         );
  NOR2_X1 U16249 ( .A1(n14405), .A2(n14404), .ZN(n14406) );
  INV_X1 U16250 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n14411) );
  NOR2_X1 U16251 ( .A1(n14409), .A2(n14408), .ZN(n14410) );
  AOI21_X1 U16252 ( .B1(P3_ADDR_REG_18__SCAN_IN), .B2(n14411), .A(n14410), 
        .ZN(n14415) );
  XNOR2_X1 U16253 ( .A(n14412), .B(P2_ADDR_REG_19__SCAN_IN), .ZN(n14413) );
  XNOR2_X1 U16254 ( .A(n14413), .B(P1_ADDR_REG_19__SCAN_IN), .ZN(n14414) );
  XNOR2_X1 U16255 ( .A(n14415), .B(n14414), .ZN(n14416) );
  XNOR2_X1 U16256 ( .A(n14417), .B(n14416), .ZN(SUB_1596_U4) );
  NOR2_X1 U16257 ( .A1(n14419), .A2(n14418), .ZN(n14439) );
  AOI21_X1 U16258 ( .B1(n14439), .B2(n15049), .A(n14420), .ZN(n14425) );
  AOI22_X1 U16259 ( .A1(n14437), .A2(n14423), .B1(n15066), .B2(
        P3_REG2_REG_31__SCAN_IN), .ZN(n14421) );
  NAND2_X1 U16260 ( .A1(n14425), .A2(n14421), .ZN(P3_U3202) );
  AOI22_X1 U16261 ( .A1(n14423), .A2(n14440), .B1(P3_REG2_REG_30__SCAN_IN), 
        .B2(n15066), .ZN(n14424) );
  NAND2_X1 U16262 ( .A1(n14425), .A2(n14424), .ZN(P3_U3203) );
  XOR2_X1 U16263 ( .A(n14432), .B(n14426), .Z(n14429) );
  AOI222_X1 U16264 ( .A1(n15056), .A2(n14429), .B1(n14428), .B2(n15052), .C1(
        n14427), .C2(n15038), .ZN(n14448) );
  AOI22_X1 U16265 ( .A1(n15066), .A2(P3_REG2_REG_11__SCAN_IN), .B1(n14430), 
        .B2(n15058), .ZN(n14436) );
  OAI21_X1 U16266 ( .B1(n7165), .B2(n7164), .A(n14433), .ZN(n14451) );
  NOR2_X1 U16267 ( .A1(n14434), .A2(n15099), .ZN(n14450) );
  AOI22_X1 U16268 ( .A1(n14451), .A2(n15063), .B1(n14450), .B2(n15062), .ZN(
        n14435) );
  OAI211_X1 U16269 ( .C1(n15066), .C2(n14448), .A(n14436), .B(n14435), .ZN(
        P3_U3222) );
  AOI21_X1 U16270 ( .B1(n14437), .B2(n14441), .A(n14439), .ZN(n14452) );
  INV_X1 U16271 ( .A(P3_REG1_REG_31__SCAN_IN), .ZN(n14438) );
  AOI22_X1 U16272 ( .A1(n15131), .A2(n14452), .B1(n14438), .B2(n15129), .ZN(
        P3_U3490) );
  AOI21_X1 U16273 ( .B1(n14441), .B2(n14440), .A(n14439), .ZN(n14453) );
  INV_X1 U16274 ( .A(P3_REG1_REG_30__SCAN_IN), .ZN(n14442) );
  AOI22_X1 U16275 ( .A1(n15131), .A2(n14453), .B1(n14442), .B2(n15129), .ZN(
        P3_U3489) );
  NAND2_X1 U16276 ( .A1(n14443), .A2(n15094), .ZN(n14445) );
  INV_X1 U16277 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n14447) );
  AOI22_X1 U16278 ( .A1(n15131), .A2(n14454), .B1(n14447), .B2(n15129), .ZN(
        P3_U3471) );
  INV_X1 U16279 ( .A(n14448), .ZN(n14449) );
  AOI211_X1 U16280 ( .C1(n15094), .C2(n14451), .A(n14450), .B(n14449), .ZN(
        n14455) );
  AOI22_X1 U16281 ( .A1(n15131), .A2(n14455), .B1(n15377), .B2(n15129), .ZN(
        P3_U3470) );
  AOI22_X1 U16282 ( .A1(n15110), .A2(n14452), .B1(n11902), .B2(n15109), .ZN(
        P3_U3458) );
  AOI22_X1 U16283 ( .A1(n15110), .A2(n14453), .B1(n11841), .B2(n15109), .ZN(
        P3_U3457) );
  AOI22_X1 U16284 ( .A1(n15110), .A2(n14454), .B1(n8833), .B2(n15109), .ZN(
        P3_U3426) );
  AOI22_X1 U16285 ( .A1(n15110), .A2(n14455), .B1(n8606), .B2(n15109), .ZN(
        P3_U3423) );
  OAI21_X1 U16286 ( .B1(n6688), .B2(n14457), .A(n14456), .ZN(n14463) );
  NOR2_X1 U16287 ( .A1(n14511), .A2(n14458), .ZN(n14461) );
  OAI22_X1 U16288 ( .A1(n14471), .A2(n14469), .B1(n14470), .B2(n14459), .ZN(
        n14460) );
  AOI211_X1 U16289 ( .C1(n14463), .C2(n14462), .A(n14461), .B(n14460), .ZN(
        n14465) );
  OAI211_X1 U16290 ( .C1(n14467), .C2(n14466), .A(n14465), .B(n14464), .ZN(
        P2_U3187) );
  OAI22_X1 U16291 ( .A1(n14471), .A2(n14470), .B1(n14469), .B2(n14468), .ZN(
        n14478) );
  NAND2_X1 U16292 ( .A1(n14473), .A2(n14472), .ZN(n14475) );
  AOI21_X1 U16293 ( .B1(n14476), .B2(n14475), .A(n14474), .ZN(n14477) );
  AOI211_X1 U16294 ( .C1(n14480), .C2(n14479), .A(n14478), .B(n14477), .ZN(
        n14482) );
  OAI211_X1 U16295 ( .C1(n14467), .C2(n14483), .A(n14482), .B(n14481), .ZN(
        P2_U3198) );
  INV_X1 U16296 ( .A(n14484), .ZN(n14492) );
  INV_X1 U16297 ( .A(n14485), .ZN(n14486) );
  AOI22_X1 U16298 ( .A1(n14489), .A2(n14488), .B1(n14487), .B2(n14486), .ZN(
        n14490) );
  OAI21_X1 U16299 ( .B1(n14492), .B2(n14491), .A(n14490), .ZN(n14494) );
  AOI211_X1 U16300 ( .C1(n14496), .C2(n14495), .A(n14494), .B(n14493), .ZN(
        n14497) );
  AOI22_X1 U16301 ( .A1(n13419), .A2(n7991), .B1(n14497), .B2(n14884), .ZN(
        P2_U3250) );
  INV_X1 U16302 ( .A(n14498), .ZN(n14500) );
  INV_X1 U16303 ( .A(n14899), .ZN(n14919) );
  OAI21_X1 U16304 ( .B1(n14500), .B2(n14919), .A(n14499), .ZN(n14502) );
  AOI211_X1 U16305 ( .C1(n14515), .C2(n14503), .A(n14502), .B(n14501), .ZN(
        n14525) );
  AOI22_X1 U16306 ( .A1(n14929), .A2(n14525), .B1(n15370), .B2(n14930), .ZN(
        P2_U3516) );
  OAI21_X1 U16307 ( .B1(n14505), .B2(n14919), .A(n14504), .ZN(n14507) );
  AOI211_X1 U16308 ( .C1(n14508), .C2(n14515), .A(n14507), .B(n14506), .ZN(
        n14527) );
  AOI22_X1 U16309 ( .A1(n14929), .A2(n14527), .B1(n14509), .B2(n14930), .ZN(
        P2_U3515) );
  OAI21_X1 U16310 ( .B1(n14511), .B2(n14919), .A(n14510), .ZN(n14513) );
  AOI211_X1 U16311 ( .C1(n14515), .C2(n14514), .A(n14513), .B(n14512), .ZN(
        n14529) );
  AOI22_X1 U16312 ( .A1(n14929), .A2(n14529), .B1(n11162), .B2(n14930), .ZN(
        P2_U3513) );
  INV_X1 U16313 ( .A(n14516), .ZN(n14518) );
  OAI21_X1 U16314 ( .B1(n14518), .B2(n14919), .A(n14517), .ZN(n14519) );
  AOI21_X1 U16315 ( .B1(n14520), .B2(n14923), .A(n14519), .ZN(n14521) );
  INV_X1 U16316 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n14523) );
  AOI22_X1 U16317 ( .A1(n14929), .A2(n14530), .B1(n14523), .B2(n14930), .ZN(
        P2_U3511) );
  INV_X1 U16318 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n14524) );
  AOI22_X1 U16319 ( .A1(n14925), .A2(n14525), .B1(n14524), .B2(n14924), .ZN(
        P2_U3481) );
  INV_X1 U16320 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n14526) );
  AOI22_X1 U16321 ( .A1(n14925), .A2(n14527), .B1(n14526), .B2(n14924), .ZN(
        P2_U3478) );
  INV_X1 U16322 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n14528) );
  AOI22_X1 U16323 ( .A1(n14925), .A2(n14529), .B1(n14528), .B2(n14924), .ZN(
        P2_U3472) );
  AOI22_X1 U16324 ( .A1(n14925), .A2(n14530), .B1(n7944), .B2(n14924), .ZN(
        P2_U3466) );
  XNOR2_X1 U16325 ( .A(n14532), .B(n14531), .ZN(n14536) );
  AOI222_X1 U16326 ( .A1(n14538), .A2(n14537), .B1(n14536), .B2(n14535), .C1(
        n14534), .C2(n14533), .ZN(n14540) );
  OAI211_X1 U16327 ( .C1(n14542), .C2(n14541), .A(n14540), .B(n14539), .ZN(
        P1_U3215) );
  OAI21_X1 U16328 ( .B1(n14544), .B2(n14767), .A(n14543), .ZN(n14546) );
  AOI211_X1 U16329 ( .C1(n14771), .C2(n14547), .A(n14546), .B(n14545), .ZN(
        n14569) );
  AOI22_X1 U16330 ( .A1(n14788), .A2(n14569), .B1(n14611), .B2(n14786), .ZN(
        P1_U3543) );
  OAI211_X1 U16331 ( .C1(n14550), .C2(n14767), .A(n14549), .B(n14548), .ZN(
        n14554) );
  AND3_X1 U16332 ( .A1(n14552), .A2(n14771), .A3(n14551), .ZN(n14553) );
  AOI211_X1 U16333 ( .C1(n14555), .C2(n14694), .A(n14554), .B(n14553), .ZN(
        n14571) );
  AOI22_X1 U16334 ( .A1(n14788), .A2(n14571), .B1(n13787), .B2(n14786), .ZN(
        P1_U3542) );
  OAI21_X1 U16335 ( .B1(n14557), .B2(n14767), .A(n14556), .ZN(n14560) );
  INV_X1 U16336 ( .A(n14558), .ZN(n14559) );
  AOI211_X1 U16337 ( .C1(n14561), .C2(n14771), .A(n14560), .B(n14559), .ZN(
        n14572) );
  AOI22_X1 U16338 ( .A1(n14788), .A2(n14572), .B1(n10792), .B2(n14786), .ZN(
        P1_U3541) );
  INV_X1 U16339 ( .A(n14562), .ZN(n14563) );
  OAI21_X1 U16340 ( .B1(n14564), .B2(n14767), .A(n14563), .ZN(n14567) );
  INV_X1 U16341 ( .A(n14565), .ZN(n14566) );
  AOI211_X1 U16342 ( .C1(n14568), .C2(n14771), .A(n14567), .B(n14566), .ZN(
        n14574) );
  AOI22_X1 U16343 ( .A1(n14788), .A2(n14574), .B1(n11007), .B2(n14786), .ZN(
        P1_U3539) );
  AOI22_X1 U16344 ( .A1(n14774), .A2(n14569), .B1(n9746), .B2(n14772), .ZN(
        P1_U3504) );
  INV_X1 U16345 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n14570) );
  AOI22_X1 U16346 ( .A1(n14774), .A2(n14571), .B1(n14570), .B2(n14772), .ZN(
        P1_U3501) );
  AOI22_X1 U16347 ( .A1(n14774), .A2(n14572), .B1(n11201), .B2(n14772), .ZN(
        P1_U3498) );
  INV_X1 U16348 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n14573) );
  AOI22_X1 U16349 ( .A1(n14774), .A2(n14574), .B1(n14573), .B2(n14772), .ZN(
        P1_U3492) );
  AOI21_X1 U16350 ( .B1(n14577), .B2(n14576), .A(n14575), .ZN(n14578) );
  XNOR2_X1 U16351 ( .A(n14578), .B(n14842), .ZN(SUB_1596_U69) );
  AOI21_X1 U16352 ( .B1(n14581), .B2(n14580), .A(n14579), .ZN(n14582) );
  XNOR2_X1 U16353 ( .A(n14582), .B(n14859), .ZN(SUB_1596_U68) );
  AOI21_X1 U16354 ( .B1(n14585), .B2(n14584), .A(n14583), .ZN(n14586) );
  XNOR2_X1 U16355 ( .A(n14586), .B(n11036), .ZN(SUB_1596_U67) );
  OAI21_X1 U16356 ( .B1(n14589), .B2(n14588), .A(n14587), .ZN(n14590) );
  XNOR2_X1 U16357 ( .A(n14590), .B(P2_ADDR_REG_14__SCAN_IN), .ZN(SUB_1596_U66)
         );
  OAI21_X1 U16358 ( .B1(n14593), .B2(n14592), .A(n14591), .ZN(n14594) );
  XNOR2_X1 U16359 ( .A(n14594), .B(P2_ADDR_REG_15__SCAN_IN), .ZN(SUB_1596_U65)
         );
  AOI21_X1 U16360 ( .B1(n14597), .B2(n14596), .A(n14595), .ZN(n14599) );
  XNOR2_X1 U16361 ( .A(n14599), .B(n14598), .ZN(SUB_1596_U64) );
  OAI21_X1 U16362 ( .B1(n14601), .B2(P1_REG1_REG_0__SCAN_IN), .A(n14600), .ZN(
        n14603) );
  XNOR2_X1 U16363 ( .A(n14603), .B(n14602), .ZN(n14607) );
  AOI22_X1 U16364 ( .A1(n14604), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n14605) );
  OAI21_X1 U16365 ( .B1(n14607), .B2(n14606), .A(n14605), .ZN(P1_U3243) );
  AOI21_X1 U16366 ( .B1(n14609), .B2(P1_REG2_REG_15__SCAN_IN), .A(n14608), 
        .ZN(n14620) );
  OAI21_X1 U16367 ( .B1(n14612), .B2(n14611), .A(n14610), .ZN(n14613) );
  NAND2_X1 U16368 ( .A1(n14614), .A2(n14613), .ZN(n14618) );
  NAND2_X1 U16369 ( .A1(n14616), .A2(n14615), .ZN(n14617) );
  OAI211_X1 U16370 ( .C1(n14620), .C2(n14619), .A(n14618), .B(n14617), .ZN(
        n14621) );
  INV_X1 U16371 ( .A(n14621), .ZN(n14623) );
  OAI211_X1 U16372 ( .C1(n14625), .C2(n14624), .A(n14623), .B(n14622), .ZN(
        P1_U3258) );
  OAI21_X1 U16373 ( .B1(n14627), .B2(n14628), .A(n14626), .ZN(n14632) );
  XNOR2_X1 U16374 ( .A(n14629), .B(n14628), .ZN(n14746) );
  NOR2_X1 U16375 ( .A1(n14746), .A2(n14691), .ZN(n14630) );
  AOI211_X1 U16376 ( .C1(n14694), .C2(n14632), .A(n14631), .B(n14630), .ZN(
        n14745) );
  INV_X1 U16377 ( .A(n14633), .ZN(n14634) );
  AOI222_X1 U16378 ( .A1(n14743), .A2(n14662), .B1(P1_REG2_REG_7__SCAN_IN), 
        .B2(n14674), .C1(n14673), .C2(n14634), .ZN(n14639) );
  INV_X1 U16379 ( .A(n14746), .ZN(n14637) );
  AOI211_X1 U16380 ( .C1(n14743), .C2(n14636), .A(n14663), .B(n14635), .ZN(
        n14741) );
  AOI22_X1 U16381 ( .A1(n14637), .A2(n14670), .B1(n14669), .B2(n14741), .ZN(
        n14638) );
  OAI211_X1 U16382 ( .C1(n14674), .C2(n14745), .A(n14639), .B(n14638), .ZN(
        P1_U3286) );
  INV_X1 U16383 ( .A(n14691), .ZN(n14711) );
  XNOR2_X1 U16384 ( .A(n14640), .B(n14641), .ZN(n14731) );
  XNOR2_X1 U16385 ( .A(n14642), .B(n14641), .ZN(n14643) );
  NOR2_X1 U16386 ( .A1(n14643), .A2(n14737), .ZN(n14729) );
  AOI211_X1 U16387 ( .C1(n14711), .C2(n14731), .A(n14726), .B(n14729), .ZN(
        n14652) );
  INV_X1 U16388 ( .A(n14644), .ZN(n14645) );
  AOI222_X1 U16389 ( .A1(n14649), .A2(n14662), .B1(P1_REG2_REG_5__SCAN_IN), 
        .B2(n14674), .C1(n14673), .C2(n14645), .ZN(n14651) );
  INV_X1 U16390 ( .A(n14646), .ZN(n14648) );
  AOI211_X1 U16391 ( .C1(n14649), .C2(n14648), .A(n14663), .B(n6536), .ZN(
        n14727) );
  AOI22_X1 U16392 ( .A1(n14731), .A2(n14670), .B1(n14727), .B2(n14669), .ZN(
        n14650) );
  OAI211_X1 U16393 ( .C1(n14674), .C2(n14652), .A(n14651), .B(n14650), .ZN(
        P1_U3288) );
  XNOR2_X1 U16394 ( .A(n14653), .B(n14654), .ZN(n14718) );
  XNOR2_X1 U16395 ( .A(n14655), .B(n14654), .ZN(n14657) );
  OAI21_X1 U16396 ( .B1(n14657), .B2(n14737), .A(n14656), .ZN(n14658) );
  AOI21_X1 U16397 ( .B1(n14711), .B2(n14718), .A(n14658), .ZN(n14715) );
  OAI22_X1 U16398 ( .A1(n14680), .A2(n14660), .B1(P1_REG3_REG_3__SCAN_IN), 
        .B2(n14659), .ZN(n14661) );
  AOI21_X1 U16399 ( .B1(n14662), .B2(n14664), .A(n14661), .ZN(n14672) );
  AOI21_X1 U16400 ( .B1(n14665), .B2(n14664), .A(n14663), .ZN(n14667) );
  NAND2_X1 U16401 ( .A1(n14667), .A2(n14666), .ZN(n14713) );
  INV_X1 U16402 ( .A(n14713), .ZN(n14668) );
  AOI22_X1 U16403 ( .A1(n14718), .A2(n14670), .B1(n14669), .B2(n14668), .ZN(
        n14671) );
  OAI211_X1 U16404 ( .C1(n14674), .C2(n14715), .A(n14672), .B(n14671), .ZN(
        P1_U3290) );
  AOI22_X1 U16405 ( .A1(P1_REG2_REG_0__SCAN_IN), .A2(n14674), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(n14673), .ZN(n14683) );
  OAI21_X1 U16406 ( .B1(n14676), .B2(n14675), .A(n14688), .ZN(n14682) );
  OAI22_X1 U16407 ( .A1(n6719), .A2(n14678), .B1(n14677), .B2(n9434), .ZN(
        n14686) );
  NAND3_X1 U16408 ( .A1(n14680), .A2(n14679), .A3(n14686), .ZN(n14681) );
  NAND3_X1 U16409 ( .A1(n14683), .A2(n14682), .A3(n14681), .ZN(P1_U3293) );
  AND2_X1 U16410 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n14685), .ZN(P1_U3294) );
  AND2_X1 U16411 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n14685), .ZN(P1_U3295) );
  INV_X1 U16412 ( .A(n14685), .ZN(n14684) );
  INV_X1 U16413 ( .A(P1_D_REG_29__SCAN_IN), .ZN(n15238) );
  NOR2_X1 U16414 ( .A1(n14684), .A2(n15238), .ZN(P1_U3296) );
  AND2_X1 U16415 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n14685), .ZN(P1_U3297) );
  INV_X1 U16416 ( .A(P1_D_REG_27__SCAN_IN), .ZN(n15209) );
  NOR2_X1 U16417 ( .A1(n14684), .A2(n15209), .ZN(P1_U3298) );
  AND2_X1 U16418 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n14685), .ZN(P1_U3299) );
  AND2_X1 U16419 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n14685), .ZN(P1_U3300) );
  INV_X1 U16420 ( .A(P1_D_REG_24__SCAN_IN), .ZN(n15390) );
  NOR2_X1 U16421 ( .A1(n14684), .A2(n15390), .ZN(P1_U3301) );
  AND2_X1 U16422 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n14685), .ZN(P1_U3302) );
  AND2_X1 U16423 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n14685), .ZN(P1_U3303) );
  AND2_X1 U16424 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n14685), .ZN(P1_U3304) );
  AND2_X1 U16425 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n14685), .ZN(P1_U3305) );
  AND2_X1 U16426 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n14685), .ZN(P1_U3306) );
  AND2_X1 U16427 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n14685), .ZN(P1_U3307) );
  AND2_X1 U16428 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n14685), .ZN(P1_U3308) );
  AND2_X1 U16429 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n14685), .ZN(P1_U3309) );
  AND2_X1 U16430 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n14685), .ZN(P1_U3310) );
  AND2_X1 U16431 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n14685), .ZN(P1_U3311) );
  AND2_X1 U16432 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n14685), .ZN(P1_U3312) );
  AND2_X1 U16433 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n14685), .ZN(P1_U3313) );
  AND2_X1 U16434 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n14685), .ZN(P1_U3314) );
  AND2_X1 U16435 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n14685), .ZN(P1_U3315) );
  AND2_X1 U16436 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n14685), .ZN(P1_U3316) );
  INV_X1 U16437 ( .A(P1_D_REG_8__SCAN_IN), .ZN(n15280) );
  NOR2_X1 U16438 ( .A1(n14684), .A2(n15280), .ZN(P1_U3317) );
  INV_X1 U16439 ( .A(P1_D_REG_7__SCAN_IN), .ZN(n15213) );
  NOR2_X1 U16440 ( .A1(n14684), .A2(n15213), .ZN(P1_U3318) );
  AND2_X1 U16441 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n14685), .ZN(P1_U3319) );
  AND2_X1 U16442 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n14685), .ZN(P1_U3320) );
  AND2_X1 U16443 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n14685), .ZN(P1_U3321) );
  AND2_X1 U16444 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n14685), .ZN(P1_U3322) );
  AND2_X1 U16445 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n14685), .ZN(P1_U3323) );
  NAND2_X1 U16446 ( .A1(n14724), .A2(n14737), .ZN(n14687) );
  AOI21_X1 U16447 ( .B1(n14688), .B2(n14687), .A(n14686), .ZN(n14775) );
  INV_X1 U16448 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n14689) );
  AOI22_X1 U16449 ( .A1(n14774), .A2(n14775), .B1(n14689), .B2(n14772), .ZN(
        P1_U3459) );
  AOI21_X1 U16450 ( .B1(n14747), .B2(n14691), .A(n14690), .ZN(n14701) );
  INV_X1 U16451 ( .A(n14692), .ZN(n14695) );
  NAND3_X1 U16452 ( .A1(n14695), .A2(n14694), .A3(n14693), .ZN(n14697) );
  OAI211_X1 U16453 ( .C1(n14698), .C2(n14767), .A(n14697), .B(n14696), .ZN(
        n14700) );
  NOR3_X1 U16454 ( .A1(n14701), .A2(n14700), .A3(n14699), .ZN(n14776) );
  INV_X1 U16455 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n14702) );
  AOI22_X1 U16456 ( .A1(n14774), .A2(n14776), .B1(n14702), .B2(n14772), .ZN(
        P1_U3462) );
  INV_X1 U16457 ( .A(n14708), .ZN(n14710) );
  INV_X1 U16458 ( .A(n14703), .ZN(n14705) );
  AOI211_X1 U16459 ( .C1(n14706), .C2(n14742), .A(n14705), .B(n14704), .ZN(
        n14707) );
  OAI21_X1 U16460 ( .B1(n14708), .B2(n14747), .A(n14707), .ZN(n14709) );
  AOI21_X1 U16461 ( .B1(n14711), .B2(n14710), .A(n14709), .ZN(n14777) );
  INV_X1 U16462 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n14712) );
  AOI22_X1 U16463 ( .A1(n14774), .A2(n14777), .B1(n14712), .B2(n14772), .ZN(
        P1_U3465) );
  OAI21_X1 U16464 ( .B1(n14714), .B2(n14767), .A(n14713), .ZN(n14717) );
  INV_X1 U16465 ( .A(n14715), .ZN(n14716) );
  AOI211_X1 U16466 ( .C1(n14763), .C2(n14718), .A(n14717), .B(n14716), .ZN(
        n14779) );
  AOI22_X1 U16467 ( .A1(n14774), .A2(n14779), .B1(n9324), .B2(n14772), .ZN(
        P1_U3468) );
  AOI21_X1 U16468 ( .B1(n14720), .B2(n14742), .A(n14719), .ZN(n14722) );
  OAI211_X1 U16469 ( .C1(n14724), .C2(n14723), .A(n14722), .B(n14721), .ZN(
        n14725) );
  INV_X1 U16470 ( .A(n14725), .ZN(n14780) );
  AOI22_X1 U16471 ( .A1(n14774), .A2(n14780), .B1(n9452), .B2(n14772), .ZN(
        P1_U3471) );
  OR4_X1 U16472 ( .A1(n14729), .A2(n14728), .A3(n14727), .A4(n14726), .ZN(
        n14730) );
  AOI21_X1 U16473 ( .B1(n14731), .B2(n14771), .A(n14730), .ZN(n14781) );
  INV_X1 U16474 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n14732) );
  AOI22_X1 U16475 ( .A1(n14774), .A2(n14781), .B1(n14732), .B2(n14772), .ZN(
        P1_U3474) );
  NOR3_X1 U16476 ( .A1(n14735), .A2(n14734), .A3(n14733), .ZN(n14736) );
  OAI21_X1 U16477 ( .B1(n14738), .B2(n14737), .A(n14736), .ZN(n14739) );
  AOI21_X1 U16478 ( .B1(n14740), .B2(n14771), .A(n14739), .ZN(n14782) );
  AOI22_X1 U16479 ( .A1(n14774), .A2(n14782), .B1(n10393), .B2(n14772), .ZN(
        P1_U3477) );
  AOI21_X1 U16480 ( .B1(n14743), .B2(n14742), .A(n14741), .ZN(n14744) );
  OAI211_X1 U16481 ( .C1(n14747), .C2(n14746), .A(n14745), .B(n14744), .ZN(
        n14748) );
  INV_X1 U16482 ( .A(n14748), .ZN(n14783) );
  INV_X1 U16483 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n14749) );
  AOI22_X1 U16484 ( .A1(n14774), .A2(n14783), .B1(n14749), .B2(n14772), .ZN(
        P1_U3480) );
  AND2_X1 U16485 ( .A1(n14750), .A2(n14771), .ZN(n14755) );
  INV_X1 U16486 ( .A(n14751), .ZN(n14752) );
  NAND2_X1 U16487 ( .A1(n14753), .A2(n14752), .ZN(n14754) );
  NOR3_X1 U16488 ( .A1(n14756), .A2(n14755), .A3(n14754), .ZN(n14784) );
  INV_X1 U16489 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n14757) );
  AOI22_X1 U16490 ( .A1(n14774), .A2(n14784), .B1(n14757), .B2(n14772), .ZN(
        P1_U3483) );
  OAI21_X1 U16491 ( .B1(n14759), .B2(n14767), .A(n14758), .ZN(n14761) );
  AOI211_X1 U16492 ( .C1(n14763), .C2(n14762), .A(n14761), .B(n14760), .ZN(
        n14785) );
  INV_X1 U16493 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n14764) );
  AOI22_X1 U16494 ( .A1(n14774), .A2(n14785), .B1(n14764), .B2(n14772), .ZN(
        P1_U3486) );
  OAI211_X1 U16495 ( .C1(n14768), .C2(n14767), .A(n14766), .B(n14765), .ZN(
        n14769) );
  AOI21_X1 U16496 ( .B1(n14771), .B2(n14770), .A(n14769), .ZN(n14787) );
  INV_X1 U16497 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n14773) );
  AOI22_X1 U16498 ( .A1(n14774), .A2(n14787), .B1(n14773), .B2(n14772), .ZN(
        P1_U3489) );
  AOI22_X1 U16499 ( .A1(n14788), .A2(n14775), .B1(n9387), .B2(n14786), .ZN(
        P1_U3528) );
  AOI22_X1 U16500 ( .A1(n14788), .A2(n14776), .B1(n9596), .B2(n14786), .ZN(
        P1_U3529) );
  AOI22_X1 U16501 ( .A1(n14788), .A2(n14777), .B1(n9597), .B2(n14786), .ZN(
        P1_U3530) );
  INV_X1 U16502 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n14778) );
  AOI22_X1 U16503 ( .A1(n14788), .A2(n14779), .B1(n14778), .B2(n14786), .ZN(
        P1_U3531) );
  INV_X1 U16504 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n15133) );
  AOI22_X1 U16505 ( .A1(n14788), .A2(n14780), .B1(n15133), .B2(n14786), .ZN(
        P1_U3532) );
  AOI22_X1 U16506 ( .A1(n14788), .A2(n14781), .B1(n9754), .B2(n14786), .ZN(
        P1_U3533) );
  AOI22_X1 U16507 ( .A1(n14788), .A2(n14782), .B1(n9624), .B2(n14786), .ZN(
        P1_U3534) );
  AOI22_X1 U16508 ( .A1(n14788), .A2(n14783), .B1(n10409), .B2(n14786), .ZN(
        P1_U3535) );
  AOI22_X1 U16509 ( .A1(n14788), .A2(n14784), .B1(n10688), .B2(n14786), .ZN(
        P1_U3536) );
  AOI22_X1 U16510 ( .A1(n14788), .A2(n14785), .B1(n10707), .B2(n14786), .ZN(
        P1_U3537) );
  AOI22_X1 U16511 ( .A1(n14788), .A2(n14787), .B1(n10880), .B2(n14786), .ZN(
        P1_U3538) );
  NOR2_X1 U16512 ( .A1(n14789), .A2(P2_U3947), .ZN(P2_U3087) );
  AOI22_X1 U16513 ( .A1(n14789), .A2(P2_ADDR_REG_1__SCAN_IN), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(P2_U3088), .ZN(n14800) );
  XNOR2_X1 U16514 ( .A(n14790), .B(n15358), .ZN(n14792) );
  OAI22_X1 U16515 ( .A1(n14863), .A2(n14792), .B1(n14791), .B2(n14834), .ZN(
        n14793) );
  INV_X1 U16516 ( .A(n14793), .ZN(n14799) );
  NOR2_X1 U16517 ( .A1(n14794), .A2(n9565), .ZN(n14797) );
  OAI211_X1 U16518 ( .C1(n14797), .C2(n14796), .A(n14870), .B(n14795), .ZN(
        n14798) );
  NAND3_X1 U16519 ( .A1(n14800), .A2(n14799), .A3(n14798), .ZN(P2_U3215) );
  AOI211_X1 U16520 ( .C1(n14803), .C2(n14802), .A(n14863), .B(n14801), .ZN(
        n14804) );
  AOI211_X1 U16521 ( .C1(n14868), .C2(n14806), .A(n14805), .B(n14804), .ZN(
        n14812) );
  AOI211_X1 U16522 ( .C1(n14809), .C2(n14808), .A(n14836), .B(n14807), .ZN(
        n14810) );
  INV_X1 U16523 ( .A(n14810), .ZN(n14811) );
  OAI211_X1 U16524 ( .C1(n14874), .C2(n7037), .A(n14812), .B(n14811), .ZN(
        P2_U3221) );
  INV_X1 U16525 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n14826) );
  INV_X1 U16526 ( .A(n14813), .ZN(n14818) );
  AOI211_X1 U16527 ( .C1(n14816), .C2(n14815), .A(n14863), .B(n14814), .ZN(
        n14817) );
  AOI211_X1 U16528 ( .C1(n14868), .C2(n14819), .A(n14818), .B(n14817), .ZN(
        n14825) );
  AOI211_X1 U16529 ( .C1(n14822), .C2(n14821), .A(n14836), .B(n14820), .ZN(
        n14823) );
  INV_X1 U16530 ( .A(n14823), .ZN(n14824) );
  OAI211_X1 U16531 ( .C1(n14874), .C2(n14826), .A(n14825), .B(n14824), .ZN(
        P2_U3222) );
  AOI211_X1 U16532 ( .C1(n14829), .C2(n14828), .A(n14863), .B(n14827), .ZN(
        n14839) );
  INV_X1 U16533 ( .A(n14830), .ZN(n14833) );
  INV_X1 U16534 ( .A(n14831), .ZN(n14832) );
  AOI21_X1 U16535 ( .B1(n14833), .B2(n14832), .A(n14845), .ZN(n14837) );
  OAI22_X1 U16536 ( .A1(n14837), .A2(n14836), .B1(n14835), .B2(n14834), .ZN(
        n14838) );
  NOR2_X1 U16537 ( .A1(n14839), .A2(n14838), .ZN(n14841) );
  OAI211_X1 U16538 ( .C1(n14842), .C2(n14874), .A(n14841), .B(n14840), .ZN(
        P2_U3225) );
  OR3_X1 U16539 ( .A1(n14845), .A2(n14844), .A3(n14843), .ZN(n14846) );
  NAND2_X1 U16540 ( .A1(n14847), .A2(n14846), .ZN(n14856) );
  NAND2_X1 U16541 ( .A1(n14849), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n14848) );
  OAI21_X1 U16542 ( .B1(n14849), .B2(P2_REG1_REG_12__SCAN_IN), .A(n14848), 
        .ZN(n14851) );
  OAI21_X1 U16543 ( .B1(n14852), .B2(n14851), .A(n14850), .ZN(n14854) );
  AOI222_X1 U16544 ( .A1(n14856), .A2(n14870), .B1(n14855), .B2(n14868), .C1(
        n14854), .C2(n14853), .ZN(n14858) );
  OAI211_X1 U16545 ( .C1(n14859), .C2(n14874), .A(n14858), .B(n14857), .ZN(
        P2_U3226) );
  NOR2_X1 U16546 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n14860), .ZN(n14866) );
  INV_X1 U16547 ( .A(n14861), .ZN(n14862) );
  AOI211_X1 U16548 ( .C1(n7990), .C2(n14864), .A(n14863), .B(n14862), .ZN(
        n14865) );
  AOI211_X1 U16549 ( .C1(n14868), .C2(n14867), .A(n14866), .B(n14865), .ZN(
        n14873) );
  OAI211_X1 U16550 ( .C1(n14871), .C2(P2_REG2_REG_15__SCAN_IN), .A(n14870), 
        .B(n14869), .ZN(n14872) );
  OAI211_X1 U16551 ( .C1(n14874), .C2(n15410), .A(n14873), .B(n14872), .ZN(
        P2_U3229) );
  INV_X1 U16552 ( .A(n14875), .ZN(n14878) );
  OAI22_X1 U16553 ( .A1(n14878), .A2(n14876), .B1(n7761), .B2(n14877), .ZN(
        n14881) );
  INV_X1 U16554 ( .A(n14879), .ZN(n14880) );
  AOI211_X1 U16555 ( .C1(n14883), .C2(n14882), .A(n14881), .B(n14880), .ZN(
        n14885) );
  AOI22_X1 U16556 ( .A1(n13419), .A2(n9565), .B1(n14885), .B2(n14884), .ZN(
        P2_U3265) );
  AND2_X1 U16557 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n14887), .ZN(P2_U3266) );
  INV_X1 U16558 ( .A(n14887), .ZN(n14888) );
  INV_X1 U16559 ( .A(P2_D_REG_30__SCAN_IN), .ZN(n15245) );
  NOR2_X1 U16560 ( .A1(n14888), .A2(n15245), .ZN(P2_U3267) );
  INV_X1 U16561 ( .A(P2_D_REG_29__SCAN_IN), .ZN(n15294) );
  NOR2_X1 U16562 ( .A1(n14888), .A2(n15294), .ZN(P2_U3268) );
  AND2_X1 U16563 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n14887), .ZN(P2_U3269) );
  AND2_X1 U16564 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n14887), .ZN(P2_U3270) );
  INV_X1 U16565 ( .A(P2_D_REG_26__SCAN_IN), .ZN(n15395) );
  NOR2_X1 U16566 ( .A1(n14888), .A2(n15395), .ZN(P2_U3271) );
  AND2_X1 U16567 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n14887), .ZN(P2_U3272) );
  AND2_X1 U16568 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n14887), .ZN(P2_U3273) );
  AND2_X1 U16569 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n14887), .ZN(P2_U3274) );
  AND2_X1 U16570 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n14887), .ZN(P2_U3275) );
  AND2_X1 U16571 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n14887), .ZN(P2_U3276) );
  AND2_X1 U16572 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n14887), .ZN(P2_U3277) );
  INV_X1 U16573 ( .A(P2_D_REG_19__SCAN_IN), .ZN(n15375) );
  NOR2_X1 U16574 ( .A1(n14888), .A2(n15375), .ZN(P2_U3278) );
  AND2_X1 U16575 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n14887), .ZN(P2_U3279) );
  AND2_X1 U16576 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n14887), .ZN(P2_U3280) );
  AND2_X1 U16577 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n14887), .ZN(P2_U3281) );
  AND2_X1 U16578 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n14887), .ZN(P2_U3282) );
  INV_X1 U16579 ( .A(P2_D_REG_14__SCAN_IN), .ZN(n15267) );
  NOR2_X1 U16580 ( .A1(n14888), .A2(n15267), .ZN(P2_U3283) );
  AND2_X1 U16581 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n14887), .ZN(P2_U3284) );
  AND2_X1 U16582 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n14887), .ZN(P2_U3285) );
  AND2_X1 U16583 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n14887), .ZN(P2_U3286) );
  AND2_X1 U16584 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n14887), .ZN(P2_U3287) );
  AND2_X1 U16585 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n14887), .ZN(P2_U3288) );
  INV_X1 U16586 ( .A(P2_D_REG_8__SCAN_IN), .ZN(n15388) );
  NOR2_X1 U16587 ( .A1(n14888), .A2(n15388), .ZN(P2_U3289) );
  AND2_X1 U16588 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n14887), .ZN(P2_U3290) );
  INV_X1 U16589 ( .A(P2_D_REG_6__SCAN_IN), .ZN(n15242) );
  NOR2_X1 U16590 ( .A1(n14888), .A2(n15242), .ZN(P2_U3291) );
  AND2_X1 U16591 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n14887), .ZN(P2_U3292) );
  AND2_X1 U16592 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n14887), .ZN(P2_U3293) );
  AND2_X1 U16593 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n14887), .ZN(P2_U3294) );
  INV_X1 U16594 ( .A(P2_D_REG_2__SCAN_IN), .ZN(n15144) );
  NOR2_X1 U16595 ( .A1(n14888), .A2(n15144), .ZN(P2_U3295) );
  INV_X1 U16596 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n14889) );
  AOI22_X1 U16597 ( .A1(n14891), .A2(n14890), .B1(n14889), .B2(n14893), .ZN(
        P2_U3416) );
  INV_X1 U16598 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n14894) );
  AOI21_X1 U16599 ( .B1(n14894), .B2(n14893), .A(n14892), .ZN(P2_U3417) );
  AOI22_X1 U16600 ( .A1(n14925), .A2(n14895), .B1(n7760), .B2(n14924), .ZN(
        P2_U3430) );
  INV_X1 U16601 ( .A(n14896), .ZN(n14904) );
  AOI21_X1 U16602 ( .B1(n14899), .B2(n14898), .A(n14897), .ZN(n14900) );
  OAI21_X1 U16603 ( .B1(n14902), .B2(n14901), .A(n14900), .ZN(n14903) );
  AOI211_X1 U16604 ( .C1(n14906), .C2(n14905), .A(n14904), .B(n14903), .ZN(
        n14926) );
  AOI22_X1 U16605 ( .A1(n14925), .A2(n14926), .B1(n7809), .B2(n14924), .ZN(
        P2_U3442) );
  INV_X1 U16606 ( .A(n14907), .ZN(n14912) );
  OAI21_X1 U16607 ( .B1(n14909), .B2(n14919), .A(n14908), .ZN(n14911) );
  AOI211_X1 U16608 ( .C1(n14923), .C2(n14912), .A(n14911), .B(n14910), .ZN(
        n14927) );
  AOI22_X1 U16609 ( .A1(n14925), .A2(n14927), .B1(n7875), .B2(n14924), .ZN(
        P2_U3454) );
  OAI21_X1 U16610 ( .B1(n14914), .B2(n14919), .A(n14913), .ZN(n14916) );
  AOI211_X1 U16611 ( .C1(n14923), .C2(n14917), .A(n14916), .B(n14915), .ZN(
        n14928) );
  AOI22_X1 U16612 ( .A1(n14925), .A2(n14928), .B1(n7901), .B2(n14924), .ZN(
        P2_U3460) );
  OAI21_X1 U16613 ( .B1(n7402), .B2(n14919), .A(n14918), .ZN(n14921) );
  AOI211_X1 U16614 ( .C1(n14923), .C2(n14922), .A(n14921), .B(n14920), .ZN(
        n14931) );
  AOI22_X1 U16615 ( .A1(n14925), .A2(n14931), .B1(n7920), .B2(n14924), .ZN(
        P2_U3463) );
  AOI22_X1 U16616 ( .A1(n14929), .A2(n14926), .B1(n9546), .B2(n14930), .ZN(
        P2_U3503) );
  AOI22_X1 U16617 ( .A1(n14929), .A2(n14927), .B1(n9878), .B2(n14930), .ZN(
        P2_U3507) );
  AOI22_X1 U16618 ( .A1(n14929), .A2(n14928), .B1(n10163), .B2(n14930), .ZN(
        P2_U3509) );
  AOI22_X1 U16619 ( .A1(n14929), .A2(n14931), .B1(n11022), .B2(n14930), .ZN(
        P2_U3510) );
  NOR2_X1 U16620 ( .A1(P3_U3897), .A2(n15001), .ZN(P3_U3150) );
  AOI22_X1 U16621 ( .A1(n15013), .A2(P3_IR_REG_0__SCAN_IN), .B1(
        P3_REG3_REG_0__SCAN_IN), .B2(P3_U3151), .ZN(n14937) );
  NOR2_X1 U16622 ( .A1(n14932), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n14934) );
  NAND3_X1 U16623 ( .A1(n14948), .A2(n15023), .A3(n15018), .ZN(n14933) );
  OAI21_X1 U16624 ( .B1(n14935), .B2(n14934), .A(n14933), .ZN(n14936) );
  OAI211_X1 U16625 ( .C1(n14938), .C2(n15029), .A(n14937), .B(n14936), .ZN(
        P3_U3182) );
  AOI21_X1 U16626 ( .B1(n15115), .B2(n14940), .A(n14939), .ZN(n14945) );
  AOI21_X1 U16627 ( .B1(n14943), .B2(n14942), .A(n14941), .ZN(n14944) );
  OAI22_X1 U16628 ( .A1(n15018), .A2(n14945), .B1(n15023), .B2(n14944), .ZN(
        n14951) );
  XOR2_X1 U16629 ( .A(n14946), .B(n14947), .Z(n14949) );
  NOR2_X1 U16630 ( .A1(n14949), .A2(n14948), .ZN(n14950) );
  AOI211_X1 U16631 ( .C1(n15013), .C2(n14952), .A(n14951), .B(n14950), .ZN(
        n14955) );
  INV_X1 U16632 ( .A(n14953), .ZN(n14954) );
  OAI211_X1 U16633 ( .C1(n14956), .C2(n15029), .A(n14955), .B(n14954), .ZN(
        P3_U3185) );
  AOI21_X1 U16634 ( .B1(n15156), .B2(n14958), .A(n14957), .ZN(n14959) );
  OR2_X1 U16635 ( .A1(n14959), .A2(n15023), .ZN(n14970) );
  AOI21_X1 U16636 ( .B1(n15119), .B2(n14961), .A(n14960), .ZN(n14962) );
  OR2_X1 U16637 ( .A1(n14962), .A2(n15018), .ZN(n14969) );
  XNOR2_X1 U16638 ( .A(n14964), .B(n14963), .ZN(n14965) );
  NAND2_X1 U16639 ( .A1(n14965), .A2(n15015), .ZN(n14968) );
  NAND2_X1 U16640 ( .A1(n15013), .A2(n14966), .ZN(n14967) );
  AND4_X1 U16641 ( .A1(n14970), .A2(n14969), .A3(n14968), .A4(n14967), .ZN(
        n14973) );
  INV_X1 U16642 ( .A(n14971), .ZN(n14972) );
  OAI211_X1 U16643 ( .C1(n14974), .C2(n15029), .A(n14973), .B(n14972), .ZN(
        P3_U3187) );
  AOI21_X1 U16644 ( .B1(n14977), .B2(n14976), .A(n14975), .ZN(n14978) );
  OR2_X1 U16645 ( .A1(n14978), .A2(n15023), .ZN(n14990) );
  AOI21_X1 U16646 ( .B1(n14981), .B2(n14980), .A(n14979), .ZN(n14982) );
  OR2_X1 U16647 ( .A1(n14982), .A2(n15018), .ZN(n14989) );
  XNOR2_X1 U16648 ( .A(n14984), .B(n14983), .ZN(n14985) );
  NAND2_X1 U16649 ( .A1(n14985), .A2(n15015), .ZN(n14988) );
  NAND2_X1 U16650 ( .A1(n15013), .A2(n14986), .ZN(n14987) );
  AND4_X1 U16651 ( .A1(n14990), .A2(n14989), .A3(n14988), .A4(n14987), .ZN(
        n14992) );
  OAI211_X1 U16652 ( .C1(n15223), .C2(n15029), .A(n14992), .B(n14991), .ZN(
        P3_U3188) );
  AOI21_X1 U16653 ( .B1(n14994), .B2(n15316), .A(n14993), .ZN(n14998) );
  AOI21_X1 U16654 ( .B1(n14996), .B2(n15123), .A(n14995), .ZN(n14997) );
  OAI22_X1 U16655 ( .A1(n14998), .A2(n15023), .B1(n14997), .B2(n15018), .ZN(
        n14999) );
  AOI211_X1 U16656 ( .C1(P3_ADDR_REG_7__SCAN_IN), .C2(n15001), .A(n15000), .B(
        n14999), .ZN(n15007) );
  XNOR2_X1 U16657 ( .A(n15003), .B(n15002), .ZN(n15005) );
  AOI22_X1 U16658 ( .A1(n15005), .A2(n15015), .B1(n15004), .B2(n15013), .ZN(
        n15006) );
  NAND2_X1 U16659 ( .A1(n15007), .A2(n15006), .ZN(P3_U3189) );
  AOI21_X1 U16660 ( .B1(n15010), .B2(n15009), .A(n15008), .ZN(n15019) );
  XNOR2_X1 U16661 ( .A(n15012), .B(n15011), .ZN(n15016) );
  AOI22_X1 U16662 ( .A1(n15016), .A2(n15015), .B1(n15014), .B2(n15013), .ZN(
        n15017) );
  OAI21_X1 U16663 ( .B1(n15019), .B2(n15018), .A(n15017), .ZN(n15026) );
  AOI21_X1 U16664 ( .B1(n15022), .B2(n15021), .A(n15020), .ZN(n15024) );
  NOR2_X1 U16665 ( .A1(n15024), .A2(n15023), .ZN(n15025) );
  NOR2_X1 U16666 ( .A1(n15026), .A2(n15025), .ZN(n15028) );
  OAI211_X1 U16667 ( .C1(n15030), .C2(n15029), .A(n15028), .B(n15027), .ZN(
        P3_U3192) );
  INV_X1 U16668 ( .A(n15031), .ZN(n15045) );
  XNOR2_X1 U16669 ( .A(n15032), .B(n15035), .ZN(n15085) );
  AOI21_X1 U16670 ( .B1(n15035), .B2(n15034), .A(n15033), .ZN(n15044) );
  AOI22_X1 U16671 ( .A1(n15038), .A2(n15037), .B1(n15036), .B2(n15052), .ZN(
        n15042) );
  INV_X1 U16672 ( .A(n15039), .ZN(n15040) );
  NAND2_X1 U16673 ( .A1(n15085), .A2(n15040), .ZN(n15041) );
  OAI211_X1 U16674 ( .C1(n15044), .C2(n15043), .A(n15042), .B(n15041), .ZN(
        n15083) );
  AOI21_X1 U16675 ( .B1(n15045), .B2(n15085), .A(n15083), .ZN(n15050) );
  NOR2_X1 U16676 ( .A1(n15046), .A2(n15099), .ZN(n15084) );
  AOI22_X1 U16677 ( .A1(n15062), .A2(n15084), .B1(n15058), .B2(n15047), .ZN(
        n15048) );
  OAI221_X1 U16678 ( .B1(n15066), .B2(n15050), .C1(n15049), .C2(n15156), .A(
        n15048), .ZN(P3_U3228) );
  XNOR2_X1 U16679 ( .A(n15051), .B(n15059), .ZN(n15055) );
  AOI222_X1 U16680 ( .A1(n15056), .A2(n15055), .B1(n15054), .B2(n15038), .C1(
        n15053), .C2(n15052), .ZN(n15079) );
  AOI22_X1 U16681 ( .A1(n15066), .A2(P3_REG2_REG_4__SCAN_IN), .B1(n15058), 
        .B2(n15057), .ZN(n15065) );
  XNOR2_X1 U16682 ( .A(n15060), .B(n15059), .ZN(n15082) );
  NOR2_X1 U16683 ( .A1(n15061), .A2(n15099), .ZN(n15081) );
  AOI22_X1 U16684 ( .A1(n15063), .A2(n15082), .B1(n15081), .B2(n15062), .ZN(
        n15064) );
  OAI211_X1 U16685 ( .C1(n15066), .C2(n15079), .A(n15065), .B(n15064), .ZN(
        P3_U3229) );
  AOI211_X1 U16686 ( .C1(n15108), .C2(n15069), .A(n15068), .B(n15067), .ZN(
        n15112) );
  AOI22_X1 U16687 ( .A1(n15110), .A2(n15112), .B1(n8699), .B2(n15109), .ZN(
        P3_U3393) );
  INV_X1 U16688 ( .A(n15070), .ZN(n15074) );
  INV_X1 U16689 ( .A(n15071), .ZN(n15073) );
  AOI211_X1 U16690 ( .C1(n15074), .C2(n15108), .A(n15073), .B(n15072), .ZN(
        n15114) );
  AOI22_X1 U16691 ( .A1(n15110), .A2(n15114), .B1(n8723), .B2(n15109), .ZN(
        P3_U3396) );
  OAI22_X1 U16692 ( .A1(n15076), .A2(n15101), .B1(n15075), .B2(n15099), .ZN(
        n15077) );
  NOR2_X1 U16693 ( .A1(n15078), .A2(n15077), .ZN(n15116) );
  AOI22_X1 U16694 ( .A1(n15110), .A2(n15116), .B1(n8735), .B2(n15109), .ZN(
        P3_U3399) );
  INV_X1 U16695 ( .A(n15079), .ZN(n15080) );
  AOI211_X1 U16696 ( .C1(n15082), .C2(n15094), .A(n15081), .B(n15080), .ZN(
        n15118) );
  AOI22_X1 U16697 ( .A1(n15110), .A2(n15118), .B1(n8683), .B2(n15109), .ZN(
        P3_U3402) );
  AOI211_X1 U16698 ( .C1(n15085), .C2(n15108), .A(n15084), .B(n15083), .ZN(
        n15120) );
  AOI22_X1 U16699 ( .A1(n15110), .A2(n15120), .B1(n8752), .B2(n15109), .ZN(
        P3_U3405) );
  OAI22_X1 U16700 ( .A1(n15087), .A2(n15101), .B1(n15086), .B2(n15099), .ZN(
        n15088) );
  NOR2_X1 U16701 ( .A1(n15089), .A2(n15088), .ZN(n15122) );
  AOI22_X1 U16702 ( .A1(n15110), .A2(n15122), .B1(n8663), .B2(n15109), .ZN(
        P3_U3408) );
  OAI21_X1 U16703 ( .B1(n15091), .B2(n15101), .A(n15090), .ZN(n15092) );
  NOR2_X1 U16704 ( .A1(n15093), .A2(n15092), .ZN(n15124) );
  AOI22_X1 U16705 ( .A1(n15110), .A2(n15124), .B1(n8761), .B2(n15109), .ZN(
        P3_U3411) );
  NAND2_X1 U16706 ( .A1(n15095), .A2(n15094), .ZN(n15097) );
  AOI22_X1 U16707 ( .A1(n15110), .A2(n15126), .B1(n8782), .B2(n15109), .ZN(
        P3_U3414) );
  OAI22_X1 U16708 ( .A1(n15102), .A2(n15101), .B1(n15100), .B2(n15099), .ZN(
        n15103) );
  NOR2_X1 U16709 ( .A1(n15104), .A2(n15103), .ZN(n15128) );
  AOI22_X1 U16710 ( .A1(n15110), .A2(n15128), .B1(n8799), .B2(n15109), .ZN(
        P3_U3417) );
  AOI211_X1 U16711 ( .C1(n15108), .C2(n15107), .A(n15106), .B(n15105), .ZN(
        n15130) );
  AOI22_X1 U16712 ( .A1(n15110), .A2(n15130), .B1(n8613), .B2(n15109), .ZN(
        P3_U3420) );
  AOI22_X1 U16713 ( .A1(n15131), .A2(n15112), .B1(n15111), .B2(n15129), .ZN(
        P3_U3460) );
  AOI22_X1 U16714 ( .A1(n15131), .A2(n15114), .B1(n15113), .B2(n15129), .ZN(
        P3_U3461) );
  AOI22_X1 U16715 ( .A1(n15131), .A2(n15116), .B1(n15115), .B2(n15129), .ZN(
        P3_U3462) );
  AOI22_X1 U16716 ( .A1(n15131), .A2(n15118), .B1(n15117), .B2(n15129), .ZN(
        P3_U3463) );
  AOI22_X1 U16717 ( .A1(n15131), .A2(n15120), .B1(n15119), .B2(n15129), .ZN(
        P3_U3464) );
  AOI22_X1 U16718 ( .A1(n15131), .A2(n15122), .B1(n15121), .B2(n15129), .ZN(
        P3_U3465) );
  AOI22_X1 U16719 ( .A1(n15131), .A2(n15124), .B1(n15123), .B2(n15129), .ZN(
        P3_U3466) );
  AOI22_X1 U16720 ( .A1(n15131), .A2(n15126), .B1(n15125), .B2(n15129), .ZN(
        P3_U3467) );
  AOI22_X1 U16721 ( .A1(n15131), .A2(n15128), .B1(n15127), .B2(n15129), .ZN(
        P3_U3468) );
  AOI22_X1 U16722 ( .A1(n15131), .A2(n15130), .B1(n15269), .B2(n15129), .ZN(
        P3_U3469) );
  AOI22_X1 U16723 ( .A1(n15353), .A2(keyinput97), .B1(n15133), .B2(keyinput99), 
        .ZN(n15132) );
  OAI221_X1 U16724 ( .B1(n15353), .B2(keyinput97), .C1(n15133), .C2(keyinput99), .A(n15132), .ZN(n15142) );
  AOI22_X1 U16725 ( .A1(n15136), .A2(keyinput89), .B1(keyinput125), .B2(n15135), .ZN(n15134) );
  OAI221_X1 U16726 ( .B1(n15136), .B2(keyinput89), .C1(n15135), .C2(
        keyinput125), .A(n15134), .ZN(n15141) );
  AOI22_X1 U16727 ( .A1(n15378), .A2(keyinput105), .B1(n15379), .B2(keyinput47), .ZN(n15137) );
  OAI221_X1 U16728 ( .B1(n15378), .B2(keyinput105), .C1(n15379), .C2(
        keyinput47), .A(n15137), .ZN(n15140) );
  AOI22_X1 U16729 ( .A1(n13003), .A2(keyinput107), .B1(keyinput100), .B2(n8279), .ZN(n15138) );
  OAI221_X1 U16730 ( .B1(n13003), .B2(keyinput107), .C1(n8279), .C2(
        keyinput100), .A(n15138), .ZN(n15139) );
  NOR4_X1 U16731 ( .A1(n15142), .A2(n15141), .A3(n15140), .A4(n15139), .ZN(
        n15182) );
  AOI22_X1 U16732 ( .A1(n10688), .A2(keyinput46), .B1(keyinput55), .B2(n15144), 
        .ZN(n15143) );
  OAI221_X1 U16733 ( .B1(n10688), .B2(keyinput46), .C1(n15144), .C2(keyinput55), .A(n15143), .ZN(n15153) );
  AOI22_X1 U16734 ( .A1(n15146), .A2(keyinput19), .B1(n15377), .B2(keyinput2), 
        .ZN(n15145) );
  OAI221_X1 U16735 ( .B1(n15146), .B2(keyinput19), .C1(n15377), .C2(keyinput2), 
        .A(n15145), .ZN(n15152) );
  AOI22_X1 U16736 ( .A1(n13361), .A2(keyinput85), .B1(n8613), .B2(keyinput31), 
        .ZN(n15147) );
  OAI221_X1 U16737 ( .B1(n13361), .B2(keyinput85), .C1(n8613), .C2(keyinput31), 
        .A(n15147), .ZN(n15151) );
  XOR2_X1 U16738 ( .A(n8593), .B(keyinput76), .Z(n15149) );
  XNOR2_X1 U16739 ( .A(P2_IR_REG_12__SCAN_IN), .B(keyinput82), .ZN(n15148) );
  NAND2_X1 U16740 ( .A1(n15149), .A2(n15148), .ZN(n15150) );
  NOR4_X1 U16741 ( .A1(n15153), .A2(n15152), .A3(n15151), .A4(n15150), .ZN(
        n15181) );
  AOI22_X1 U16742 ( .A1(n15156), .A2(keyinput52), .B1(n15155), .B2(keyinput16), 
        .ZN(n15154) );
  OAI221_X1 U16743 ( .B1(n15156), .B2(keyinput52), .C1(n15155), .C2(keyinput16), .A(n15154), .ZN(n15165) );
  AOI22_X1 U16744 ( .A1(n15158), .A2(keyinput86), .B1(keyinput15), .B2(n10703), 
        .ZN(n15157) );
  OAI221_X1 U16745 ( .B1(n15158), .B2(keyinput86), .C1(n10703), .C2(keyinput15), .A(n15157), .ZN(n15164) );
  AOI22_X1 U16746 ( .A1(n15160), .A2(keyinput60), .B1(keyinput58), .B2(n13004), 
        .ZN(n15159) );
  OAI221_X1 U16747 ( .B1(n15160), .B2(keyinput60), .C1(n13004), .C2(keyinput58), .A(n15159), .ZN(n15163) );
  AOI22_X1 U16748 ( .A1(n15375), .A2(keyinput122), .B1(n15376), .B2(
        keyinput121), .ZN(n15161) );
  OAI221_X1 U16749 ( .B1(n15375), .B2(keyinput122), .C1(n15376), .C2(
        keyinput121), .A(n15161), .ZN(n15162) );
  NOR4_X1 U16750 ( .A1(n15165), .A2(n15164), .A3(n15163), .A4(n15162), .ZN(
        n15180) );
  AOI22_X1 U16751 ( .A1(P3_U3151), .A2(keyinput4), .B1(n15167), .B2(
        keyinput113), .ZN(n15166) );
  OAI221_X1 U16752 ( .B1(P3_U3151), .B2(keyinput4), .C1(n15167), .C2(
        keyinput113), .A(n15166), .ZN(n15178) );
  AOI22_X1 U16753 ( .A1(n15170), .A2(keyinput78), .B1(keyinput56), .B2(n15169), 
        .ZN(n15168) );
  OAI221_X1 U16754 ( .B1(n15170), .B2(keyinput78), .C1(n15169), .C2(keyinput56), .A(n15168), .ZN(n15177) );
  AOI22_X1 U16755 ( .A1(n15354), .A2(keyinput18), .B1(n15172), .B2(keyinput14), 
        .ZN(n15171) );
  OAI221_X1 U16756 ( .B1(n15354), .B2(keyinput18), .C1(n15172), .C2(keyinput14), .A(n15171), .ZN(n15176) );
  XOR2_X1 U16757 ( .A(n13587), .B(keyinput119), .Z(n15174) );
  XNOR2_X1 U16758 ( .A(n6756), .B(keyinput74), .ZN(n15173) );
  NAND2_X1 U16759 ( .A1(n15174), .A2(n15173), .ZN(n15175) );
  NOR4_X1 U16760 ( .A1(n15178), .A2(n15177), .A3(n15176), .A4(n15175), .ZN(
        n15179) );
  NAND4_X1 U16761 ( .A1(n15182), .A2(n15181), .A3(n15180), .A4(n15179), .ZN(
        n15344) );
  AOI22_X1 U16762 ( .A1(n15368), .A2(keyinput65), .B1(keyinput44), .B2(n11444), 
        .ZN(n15183) );
  OAI221_X1 U16763 ( .B1(n15368), .B2(keyinput65), .C1(n11444), .C2(keyinput44), .A(n15183), .ZN(n15192) );
  AOI22_X1 U16764 ( .A1(n15349), .A2(keyinput0), .B1(n10948), .B2(keyinput106), 
        .ZN(n15184) );
  OAI221_X1 U16765 ( .B1(n15349), .B2(keyinput0), .C1(n10948), .C2(keyinput106), .A(n15184), .ZN(n15191) );
  INV_X1 U16766 ( .A(keyinput77), .ZN(n15186) );
  AOI22_X1 U16767 ( .A1(n15370), .A2(keyinput102), .B1(P3_DATAO_REG_1__SCAN_IN), .B2(n15186), .ZN(n15185) );
  OAI221_X1 U16768 ( .B1(n15370), .B2(keyinput102), .C1(n15186), .C2(
        P3_DATAO_REG_1__SCAN_IN), .A(n15185), .ZN(n15190) );
  XNOR2_X1 U16769 ( .A(P2_IR_REG_23__SCAN_IN), .B(keyinput81), .ZN(n15188) );
  XNOR2_X1 U16770 ( .A(P1_REG3_REG_5__SCAN_IN), .B(keyinput61), .ZN(n15187) );
  NAND2_X1 U16771 ( .A1(n15188), .A2(n15187), .ZN(n15189) );
  NOR4_X1 U16772 ( .A1(n15192), .A2(n15191), .A3(n15190), .A4(n15189), .ZN(
        n15235) );
  AOI22_X1 U16773 ( .A1(n15194), .A2(keyinput73), .B1(n15355), .B2(keyinput41), 
        .ZN(n15193) );
  OAI221_X1 U16774 ( .B1(n15194), .B2(keyinput73), .C1(n15355), .C2(keyinput41), .A(n15193), .ZN(n15205) );
  AOI22_X1 U16775 ( .A1(n15197), .A2(keyinput95), .B1(keyinput27), .B2(n15196), 
        .ZN(n15195) );
  OAI221_X1 U16776 ( .B1(n15197), .B2(keyinput95), .C1(n15196), .C2(keyinput27), .A(n15195), .ZN(n15204) );
  INV_X1 U16777 ( .A(P3_REG3_REG_28__SCAN_IN), .ZN(n15199) );
  AOI22_X1 U16778 ( .A1(n15199), .A2(keyinput126), .B1(keyinput11), .B2(n15369), .ZN(n15198) );
  OAI221_X1 U16779 ( .B1(n15199), .B2(keyinput126), .C1(n15369), .C2(
        keyinput11), .A(n15198), .ZN(n15203) );
  XNOR2_X1 U16780 ( .A(P3_REG1_REG_21__SCAN_IN), .B(keyinput93), .ZN(n15201)
         );
  XNOR2_X1 U16781 ( .A(P2_IR_REG_19__SCAN_IN), .B(keyinput87), .ZN(n15200) );
  NAND2_X1 U16782 ( .A1(n15201), .A2(n15200), .ZN(n15202) );
  NOR4_X1 U16783 ( .A1(n15205), .A2(n15204), .A3(n15203), .A4(n15202), .ZN(
        n15234) );
  AOI22_X1 U16784 ( .A1(n15207), .A2(keyinput59), .B1(keyinput104), .B2(n14660), .ZN(n15206) );
  OAI221_X1 U16785 ( .B1(n15207), .B2(keyinput59), .C1(n14660), .C2(
        keyinput104), .A(n15206), .ZN(n15219) );
  AOI22_X1 U16786 ( .A1(n15210), .A2(keyinput79), .B1(n15209), .B2(keyinput114), .ZN(n15208) );
  OAI221_X1 U16787 ( .B1(n15210), .B2(keyinput79), .C1(n15209), .C2(
        keyinput114), .A(n15208), .ZN(n15218) );
  AOI22_X1 U16788 ( .A1(n15213), .A2(keyinput123), .B1(n15212), .B2(keyinput69), .ZN(n15211) );
  OAI221_X1 U16789 ( .B1(n15213), .B2(keyinput123), .C1(n15212), .C2(
        keyinput69), .A(n15211), .ZN(n15217) );
  XNOR2_X1 U16790 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(keyinput28), .ZN(n15215)
         );
  XNOR2_X1 U16791 ( .A(SI_3_), .B(keyinput23), .ZN(n15214) );
  NAND2_X1 U16792 ( .A1(n15215), .A2(n15214), .ZN(n15216) );
  NOR4_X1 U16793 ( .A1(n15219), .A2(n15218), .A3(n15217), .A4(n15216), .ZN(
        n15233) );
  AOI22_X1 U16794 ( .A1(n15221), .A2(keyinput22), .B1(keyinput127), .B2(n11162), .ZN(n15220) );
  OAI221_X1 U16795 ( .B1(n15221), .B2(keyinput22), .C1(n11162), .C2(
        keyinput127), .A(n15220), .ZN(n15231) );
  AOI22_X1 U16796 ( .A1(n15223), .A2(keyinput9), .B1(n15396), .B2(keyinput45), 
        .ZN(n15222) );
  OAI221_X1 U16797 ( .B1(n15223), .B2(keyinput9), .C1(n15396), .C2(keyinput45), 
        .A(n15222), .ZN(n15230) );
  XOR2_X1 U16798 ( .A(n15224), .B(keyinput13), .Z(n15228) );
  XNOR2_X1 U16799 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(keyinput110), .ZN(n15227)
         );
  XNOR2_X1 U16800 ( .A(P1_IR_REG_5__SCAN_IN), .B(keyinput3), .ZN(n15226) );
  XNOR2_X1 U16801 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(keyinput21), .ZN(n15225)
         );
  NAND4_X1 U16802 ( .A1(n15228), .A2(n15227), .A3(n15226), .A4(n15225), .ZN(
        n15229) );
  NOR3_X1 U16803 ( .A1(n15231), .A2(n15230), .A3(n15229), .ZN(n15232) );
  NAND4_X1 U16804 ( .A1(n15235), .A2(n15234), .A3(n15233), .A4(n15232), .ZN(
        n15343) );
  AOI22_X1 U16805 ( .A1(n15238), .A2(keyinput57), .B1(keyinput38), .B2(n15237), 
        .ZN(n15236) );
  OAI221_X1 U16806 ( .B1(n15238), .B2(keyinput57), .C1(n15237), .C2(keyinput38), .A(n15236), .ZN(n15249) );
  AOI22_X1 U16807 ( .A1(n15395), .A2(keyinput33), .B1(n15240), .B2(keyinput40), 
        .ZN(n15239) );
  OAI221_X1 U16808 ( .B1(n15395), .B2(keyinput33), .C1(n15240), .C2(keyinput40), .A(n15239), .ZN(n15248) );
  AOI22_X1 U16809 ( .A1(n15242), .A2(keyinput32), .B1(keyinput35), .B2(n15388), 
        .ZN(n15241) );
  OAI221_X1 U16810 ( .B1(n15242), .B2(keyinput32), .C1(n15388), .C2(keyinput35), .A(n15241), .ZN(n15247) );
  AOI22_X1 U16811 ( .A1(n15245), .A2(keyinput92), .B1(keyinput10), .B2(n15244), 
        .ZN(n15243) );
  OAI221_X1 U16812 ( .B1(n15245), .B2(keyinput92), .C1(n15244), .C2(keyinput10), .A(n15243), .ZN(n15246) );
  NOR4_X1 U16813 ( .A1(n15249), .A2(n15248), .A3(n15247), .A4(n15246), .ZN(
        n15289) );
  AOI22_X1 U16814 ( .A1(n15387), .A2(keyinput34), .B1(keyinput62), .B2(n9545), 
        .ZN(n15250) );
  OAI221_X1 U16815 ( .B1(n15387), .B2(keyinput34), .C1(n9545), .C2(keyinput62), 
        .A(n15250), .ZN(n15259) );
  AOI22_X1 U16816 ( .A1(n13977), .A2(keyinput26), .B1(keyinput101), .B2(n15385), .ZN(n15251) );
  OAI221_X1 U16817 ( .B1(n13977), .B2(keyinput26), .C1(n15385), .C2(
        keyinput101), .A(n15251), .ZN(n15258) );
  AOI22_X1 U16818 ( .A1(n15386), .A2(keyinput75), .B1(n15253), .B2(keyinput36), 
        .ZN(n15252) );
  OAI221_X1 U16819 ( .B1(n15386), .B2(keyinput75), .C1(n15253), .C2(keyinput36), .A(n15252), .ZN(n15257) );
  XOR2_X1 U16820 ( .A(n8654), .B(keyinput109), .Z(n15255) );
  XNOR2_X1 U16821 ( .A(SI_5_), .B(keyinput5), .ZN(n15254) );
  NAND2_X1 U16822 ( .A1(n15255), .A2(n15254), .ZN(n15256) );
  NOR4_X1 U16823 ( .A1(n15259), .A2(n15258), .A3(n15257), .A4(n15256), .ZN(
        n15288) );
  INV_X1 U16824 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n15389) );
  AOI22_X1 U16825 ( .A1(n15389), .A2(keyinput80), .B1(n15261), .B2(keyinput112), .ZN(n15260) );
  OAI221_X1 U16826 ( .B1(n15389), .B2(keyinput80), .C1(n15261), .C2(
        keyinput112), .A(n15260), .ZN(n15265) );
  XNOR2_X1 U16827 ( .A(n15262), .B(keyinput91), .ZN(n15264) );
  XNOR2_X1 U16828 ( .A(n15390), .B(keyinput120), .ZN(n15263) );
  OR3_X1 U16829 ( .A1(n15265), .A2(n15264), .A3(n15263), .ZN(n15273) );
  AOI22_X1 U16830 ( .A1(n15267), .A2(keyinput24), .B1(keyinput84), .B2(n10775), 
        .ZN(n15266) );
  OAI221_X1 U16831 ( .B1(n15267), .B2(keyinput24), .C1(n10775), .C2(keyinput84), .A(n15266), .ZN(n15272) );
  AOI22_X1 U16832 ( .A1(n15270), .A2(keyinput51), .B1(n15269), .B2(keyinput70), 
        .ZN(n15268) );
  OAI221_X1 U16833 ( .B1(n15270), .B2(keyinput51), .C1(n15269), .C2(keyinput70), .A(n15268), .ZN(n15271) );
  NOR3_X1 U16834 ( .A1(n15273), .A2(n15272), .A3(n15271), .ZN(n15287) );
  AOI22_X1 U16835 ( .A1(n10136), .A2(keyinput20), .B1(keyinput6), .B2(n10173), 
        .ZN(n15274) );
  OAI221_X1 U16836 ( .B1(n10136), .B2(keyinput20), .C1(n10173), .C2(keyinput6), 
        .A(n15274), .ZN(n15285) );
  AOI22_X1 U16837 ( .A1(n15409), .A2(keyinput117), .B1(n15276), .B2(keyinput39), .ZN(n15275) );
  OAI221_X1 U16838 ( .B1(n15409), .B2(keyinput117), .C1(n15276), .C2(
        keyinput39), .A(n15275), .ZN(n15284) );
  INV_X1 U16839 ( .A(P3_ADDR_REG_7__SCAN_IN), .ZN(n15278) );
  AOI22_X1 U16840 ( .A1(n7886), .A2(keyinput67), .B1(keyinput1), .B2(n15278), 
        .ZN(n15277) );
  OAI221_X1 U16841 ( .B1(n7886), .B2(keyinput67), .C1(n15278), .C2(keyinput1), 
        .A(n15277), .ZN(n15283) );
  AOI22_X1 U16842 ( .A1(n15281), .A2(keyinput83), .B1(keyinput94), .B2(n15280), 
        .ZN(n15279) );
  OAI221_X1 U16843 ( .B1(n15281), .B2(keyinput83), .C1(n15280), .C2(keyinput94), .A(n15279), .ZN(n15282) );
  NOR4_X1 U16844 ( .A1(n15285), .A2(n15284), .A3(n15283), .A4(n15282), .ZN(
        n15286) );
  NAND4_X1 U16845 ( .A1(n15289), .A2(n15288), .A3(n15287), .A4(n15286), .ZN(
        n15342) );
  AOI22_X1 U16846 ( .A1(n7851), .A2(keyinput7), .B1(keyinput116), .B2(n15291), 
        .ZN(n15290) );
  OAI221_X1 U16847 ( .B1(n7851), .B2(keyinput7), .C1(n15291), .C2(keyinput116), 
        .A(n15290), .ZN(n15302) );
  AOI22_X1 U16848 ( .A1(n15294), .A2(keyinput90), .B1(n15293), .B2(keyinput53), 
        .ZN(n15292) );
  OAI221_X1 U16849 ( .B1(n15294), .B2(keyinput90), .C1(n15293), .C2(keyinput53), .A(n15292), .ZN(n15301) );
  AOI22_X1 U16850 ( .A1(n15296), .A2(keyinput43), .B1(keyinput98), .B2(n15402), 
        .ZN(n15295) );
  OAI221_X1 U16851 ( .B1(n15296), .B2(keyinput43), .C1(n15402), .C2(keyinput98), .A(n15295), .ZN(n15300) );
  XOR2_X1 U16852 ( .A(n8205), .B(keyinput12), .Z(n15298) );
  XNOR2_X1 U16853 ( .A(P3_IR_REG_5__SCAN_IN), .B(keyinput54), .ZN(n15297) );
  NAND2_X1 U16854 ( .A1(n15298), .A2(n15297), .ZN(n15299) );
  NOR4_X1 U16855 ( .A1(n15302), .A2(n15301), .A3(n15300), .A4(n15299), .ZN(
        n15340) );
  AOI22_X1 U16856 ( .A1(n15304), .A2(keyinput63), .B1(n15403), .B2(keyinput115), .ZN(n15303) );
  OAI221_X1 U16857 ( .B1(n15304), .B2(keyinput63), .C1(n15403), .C2(
        keyinput115), .A(n15303), .ZN(n15313) );
  AOI22_X1 U16858 ( .A1(n13438), .A2(keyinput96), .B1(keyinput103), .B2(n15306), .ZN(n15305) );
  OAI221_X1 U16859 ( .B1(n13438), .B2(keyinput96), .C1(n15306), .C2(
        keyinput103), .A(n15305), .ZN(n15312) );
  AOI22_X1 U16860 ( .A1(n15308), .A2(keyinput42), .B1(keyinput72), .B2(n15350), 
        .ZN(n15307) );
  OAI221_X1 U16861 ( .B1(n15308), .B2(keyinput42), .C1(n15350), .C2(keyinput72), .A(n15307), .ZN(n15311) );
  AOI22_X1 U16862 ( .A1(n8799), .A2(keyinput71), .B1(n11772), .B2(keyinput50), 
        .ZN(n15309) );
  OAI221_X1 U16863 ( .B1(n8799), .B2(keyinput71), .C1(n11772), .C2(keyinput50), 
        .A(n15309), .ZN(n15310) );
  NOR4_X1 U16864 ( .A1(n15313), .A2(n15312), .A3(n15311), .A4(n15310), .ZN(
        n15339) );
  AOI22_X1 U16865 ( .A1(n15410), .A2(keyinput30), .B1(n11029), .B2(keyinput29), 
        .ZN(n15314) );
  OAI221_X1 U16866 ( .B1(n15410), .B2(keyinput30), .C1(n11029), .C2(keyinput29), .A(n15314), .ZN(n15323) );
  AOI22_X1 U16867 ( .A1(n8735), .A2(keyinput108), .B1(keyinput48), .B2(n9452), 
        .ZN(n15315) );
  OAI221_X1 U16868 ( .B1(n8735), .B2(keyinput108), .C1(n9452), .C2(keyinput48), 
        .A(n15315), .ZN(n15322) );
  XOR2_X1 U16869 ( .A(n15316), .B(keyinput64), .Z(n15320) );
  XOR2_X1 U16870 ( .A(n9420), .B(keyinput37), .Z(n15319) );
  XNOR2_X1 U16871 ( .A(P2_IR_REG_22__SCAN_IN), .B(keyinput88), .ZN(n15318) );
  XNOR2_X1 U16872 ( .A(P2_REG1_REG_0__SCAN_IN), .B(keyinput49), .ZN(n15317) );
  NAND4_X1 U16873 ( .A1(n15320), .A2(n15319), .A3(n15318), .A4(n15317), .ZN(
        n15321) );
  NOR3_X1 U16874 ( .A1(n15323), .A2(n15322), .A3(n15321), .ZN(n15338) );
  AOI22_X1 U16875 ( .A1(n15325), .A2(keyinput118), .B1(keyinput111), .B2(n7778), .ZN(n15324) );
  OAI221_X1 U16876 ( .B1(n15325), .B2(keyinput118), .C1(n7778), .C2(
        keyinput111), .A(n15324), .ZN(n15336) );
  AOI22_X1 U16877 ( .A1(n9624), .A2(keyinput25), .B1(keyinput68), .B2(n6951), 
        .ZN(n15326) );
  OAI221_X1 U16878 ( .B1(n9624), .B2(keyinput25), .C1(n6951), .C2(keyinput68), 
        .A(n15326), .ZN(n15335) );
  INV_X1 U16879 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n15328) );
  AOI22_X1 U16880 ( .A1(n15329), .A2(keyinput66), .B1(n15328), .B2(keyinput17), 
        .ZN(n15327) );
  OAI221_X1 U16881 ( .B1(n15329), .B2(keyinput66), .C1(n15328), .C2(keyinput17), .A(n15327), .ZN(n15334) );
  XNOR2_X1 U16882 ( .A(P3_REG1_REG_28__SCAN_IN), .B(keyinput124), .ZN(n15332)
         );
  XNOR2_X1 U16883 ( .A(n15330), .B(keyinput8), .ZN(n15331) );
  NAND2_X1 U16884 ( .A1(n15332), .A2(n15331), .ZN(n15333) );
  NOR4_X1 U16885 ( .A1(n15336), .A2(n15335), .A3(n15334), .A4(n15333), .ZN(
        n15337) );
  NAND4_X1 U16886 ( .A1(n15340), .A2(n15339), .A3(n15338), .A4(n15337), .ZN(
        n15341) );
  NOR4_X1 U16887 ( .A1(n15344), .A2(n15343), .A3(n15342), .A4(n15341), .ZN(
        n15348) );
  NAND2_X1 U16888 ( .A1(n15345), .A2(P3_U3897), .ZN(n15346) );
  OAI21_X1 U16889 ( .B1(P3_U3897), .B2(P3_DATAO_REG_25__SCAN_IN), .A(n15346), 
        .ZN(n15347) );
  XNOR2_X1 U16890 ( .A(n15348), .B(n15347), .ZN(n15424) );
  NOR4_X1 U16891 ( .A1(P3_IR_REG_5__SCAN_IN), .A2(P3_IR_REG_17__SCAN_IN), .A3(
        P3_REG3_REG_24__SCAN_IN), .A4(P3_ADDR_REG_7__SCAN_IN), .ZN(n15351) );
  NAND4_X1 U16892 ( .A1(n15352), .A2(n15351), .A3(n15350), .A4(n15349), .ZN(
        n15367) );
  NAND4_X1 U16893 ( .A1(P1_REG1_REG_4__SCAN_IN), .A2(P3_D_REG_14__SCAN_IN), 
        .A3(P2_REG0_REG_28__SCAN_IN), .A4(n15353), .ZN(n15366) );
  NAND4_X1 U16894 ( .A1(P3_IR_REG_30__SCAN_IN), .A2(n15355), .A3(n8654), .A4(
        n15354), .ZN(n15365) );
  NAND3_X1 U16895 ( .A1(n15357), .A2(P3_REG3_REG_28__SCAN_IN), .A3(n15356), 
        .ZN(n15360) );
  OR4_X1 U16896 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11772), .A3(n15358), .A4(
        n13587), .ZN(n15359) );
  NOR4_X1 U16897 ( .A1(n15361), .A2(n15360), .A3(P2_IR_REG_22__SCAN_IN), .A4(
        n15359), .ZN(n15362) );
  NAND2_X1 U16898 ( .A1(n15363), .A2(n15362), .ZN(n15364) );
  NOR4_X1 U16899 ( .A1(n15367), .A2(n15366), .A3(n15365), .A4(n15364), .ZN(
        n15422) );
  NAND4_X1 U16900 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P2_IR_REG_23__SCAN_IN), 
        .A3(n10948), .A4(n15368), .ZN(n15374) );
  NAND4_X1 U16901 ( .A1(P3_D_REG_21__SCAN_IN), .A2(P1_DATAO_REG_14__SCAN_IN), 
        .A3(n6756), .A4(P2_REG0_REG_15__SCAN_IN), .ZN(n15373) );
  NAND4_X1 U16902 ( .A1(P3_REG1_REG_21__SCAN_IN), .A2(P2_DATAO_REG_26__SCAN_IN), .A3(P1_REG3_REG_20__SCAN_IN), .A4(n15369), .ZN(n15372) );
  NAND4_X1 U16903 ( .A1(P2_REG3_REG_22__SCAN_IN), .A2(P3_DATAO_REG_1__SCAN_IN), 
        .A3(n15370), .A4(n11444), .ZN(n15371) );
  NOR4_X1 U16904 ( .A1(n15374), .A2(n15373), .A3(n15372), .A4(n15371), .ZN(
        n15421) );
  NAND4_X1 U16905 ( .A1(P3_REG0_REG_14__SCAN_IN), .A2(n15376), .A3(n13004), 
        .A4(n15375), .ZN(n15384) );
  NAND4_X1 U16906 ( .A1(P3_REG0_REG_10__SCAN_IN), .A2(P2_D_REG_2__SCAN_IN), 
        .A3(n15377), .A4(n10688), .ZN(n15383) );
  NAND4_X1 U16907 ( .A1(P2_REG2_REG_21__SCAN_IN), .A2(n15379), .A3(n15378), 
        .A4(n8279), .ZN(n15382) );
  NAND4_X1 U16908 ( .A1(n15380), .A2(SI_17_), .A3(P1_REG2_REG_9__SCAN_IN), 
        .A4(P3_REG2_REG_5__SCAN_IN), .ZN(n15381) );
  NOR4_X1 U16909 ( .A1(n15384), .A2(n15383), .A3(n15382), .A4(n15381), .ZN(
        n15420) );
  NOR4_X1 U16910 ( .A1(P2_REG1_REG_2__SCAN_IN), .A2(n15387), .A3(n15386), .A4(
        n15385), .ZN(n15394) );
  NOR4_X1 U16911 ( .A1(P1_REG0_REG_28__SCAN_IN), .A2(P1_REG2_REG_23__SCAN_IN), 
        .A3(P3_DATAO_REG_12__SCAN_IN), .A4(n15388), .ZN(n15393) );
  NOR4_X1 U16912 ( .A1(P3_REG1_REG_10__SCAN_IN), .A2(P1_REG0_REG_29__SCAN_IN), 
        .A3(P2_D_REG_14__SCAN_IN), .A4(n10775), .ZN(n15392) );
  NOR4_X1 U16913 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(SI_5_), .A3(n15390), 
        .A4(n15389), .ZN(n15391) );
  NAND4_X1 U16914 ( .A1(n15394), .A2(n15393), .A3(n15392), .A4(n15391), .ZN(
        n15418) );
  NOR4_X1 U16915 ( .A1(P2_DATAO_REG_11__SCAN_IN), .A2(P1_D_REG_29__SCAN_IN), 
        .A3(P3_DATAO_REG_6__SCAN_IN), .A4(n15395), .ZN(n15401) );
  NAND4_X1 U16916 ( .A1(SI_3_), .A2(P2_REG3_REG_10__SCAN_IN), .A3(
        P2_DATAO_REG_10__SCAN_IN), .A4(P2_DATAO_REG_25__SCAN_IN), .ZN(n15399)
         );
  NOR4_X1 U16917 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), 
        .A3(n15396), .A4(n11162), .ZN(n15397) );
  NAND2_X1 U16918 ( .A1(P1_REG2_REG_3__SCAN_IN), .A2(n15397), .ZN(n15398) );
  NOR4_X1 U16919 ( .A1(n15399), .A2(P1_B_REG_SCAN_IN), .A3(P1_D_REG_7__SCAN_IN), .A4(n15398), .ZN(n15400) );
  NAND3_X1 U16920 ( .A1(n15401), .A2(n15400), .A3(P1_D_REG_27__SCAN_IN), .ZN(
        n15417) );
  NAND4_X1 U16921 ( .A1(P1_REG3_REG_10__SCAN_IN), .A2(P3_DATAO_REG_4__SCAN_IN), 
        .A3(n15403), .A4(n15402), .ZN(n15408) );
  NAND4_X1 U16922 ( .A1(P3_REG2_REG_15__SCAN_IN), .A2(P2_B_REG_SCAN_IN), .A3(
        P2_D_REG_29__SCAN_IN), .A4(P2_REG2_REG_2__SCAN_IN), .ZN(n15407) );
  NAND4_X1 U16923 ( .A1(P3_REG2_REG_6__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), 
        .A3(P2_IR_REG_1__SCAN_IN), .A4(n15404), .ZN(n15406) );
  NAND4_X1 U16924 ( .A1(P1_REG3_REG_19__SCAN_IN), .A2(P1_REG0_REG_4__SCAN_IN), 
        .A3(P2_REG1_REG_26__SCAN_IN), .A4(n9624), .ZN(n15405) );
  OR4_X1 U16925 ( .A1(n15408), .A2(n15407), .A3(n15406), .A4(n15405), .ZN(
        n15416) );
  NOR4_X1 U16926 ( .A1(P1_D_REG_8__SCAN_IN), .A2(P2_REG3_REG_9__SCAN_IN), .A3(
        P2_REG3_REG_7__SCAN_IN), .A4(n8205), .ZN(n15414) );
  NOR4_X1 U16927 ( .A1(P3_REG0_REG_16__SCAN_IN), .A2(P1_REG2_REG_28__SCAN_IN), 
        .A3(n15409), .A4(n10173), .ZN(n15413) );
  NOR4_X1 U16928 ( .A1(P3_REG0_REG_3__SCAN_IN), .A2(P1_D_REG_0__SCAN_IN), .A3(
        n11029), .A4(n15410), .ZN(n15412) );
  NOR4_X1 U16929 ( .A1(P1_REG1_REG_24__SCAN_IN), .A2(P3_REG2_REG_7__SCAN_IN), 
        .A3(P2_REG2_REG_13__SCAN_IN), .A4(n8799), .ZN(n15411) );
  NAND4_X1 U16930 ( .A1(n15414), .A2(n15413), .A3(n15412), .A4(n15411), .ZN(
        n15415) );
  NOR4_X1 U16931 ( .A1(n15418), .A2(n15417), .A3(n15416), .A4(n15415), .ZN(
        n15419) );
  NAND4_X1 U16932 ( .A1(n15422), .A2(n15421), .A3(n15420), .A4(n15419), .ZN(
        n15423) );
  XNOR2_X1 U16933 ( .A(n15424), .B(n15423), .ZN(P3_U3516) );
  XOR2_X1 U16934 ( .A(n15425), .B(n15426), .Z(SUB_1596_U59) );
  XNOR2_X1 U16935 ( .A(n15427), .B(P2_ADDR_REG_5__SCAN_IN), .ZN(SUB_1596_U58)
         );
  AOI21_X1 U16936 ( .B1(n15428), .B2(n9569), .A(n15437), .ZN(SUB_1596_U53) );
  XOR2_X1 U16937 ( .A(n15430), .B(n15429), .Z(SUB_1596_U56) );
  AOI21_X1 U16938 ( .B1(n15433), .B2(n15432), .A(n15431), .ZN(n15435) );
  XNOR2_X1 U16939 ( .A(n15435), .B(n15434), .ZN(SUB_1596_U60) );
  XOR2_X1 U16940 ( .A(n15437), .B(n15436), .Z(SUB_1596_U5) );
  NAND2_X1 U7281 ( .A1(n7482), .A2(n7481), .ZN(n11973) );
  INV_X2 U7284 ( .A(n8439), .ZN(n8517) );
  INV_X1 U7313 ( .A(n8488), .ZN(n8157) );
  CLKBUF_X1 U7323 ( .A(n14076), .Z(n6750) );
  CLKBUF_X1 U7338 ( .A(n9187), .Z(n9185) );
  CLKBUF_X1 U7339 ( .A(P1_IR_REG_13__SCAN_IN), .Z(n6756) );
  CLKBUF_X1 U7347 ( .A(P1_IR_REG_8__SCAN_IN), .Z(n6751) );
  NAND2_X1 U7359 ( .A1(n14314), .A2(n14315), .ZN(n14316) );
  INV_X1 U7368 ( .A(n14362), .ZN(n9814) );
  XNOR2_X1 U7400 ( .A(n8655), .B(n8654), .ZN(n9721) );
  CLKBUF_X1 U7407 ( .A(n13960), .Z(n6765) );
  CLKBUF_X1 U7609 ( .A(n10724), .Z(n6523) );
  CLKBUF_X2 U8091 ( .A(n7746), .Z(n6538) );
endmodule

