

module b15_C_gen_AntiSAT_k_256_8 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, 
        READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, 
        CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, 
        REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, 
        FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput_f0, keyinput_f1, 
        keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, 
        keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, 
        keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, 
        keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, 
        keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, 
        keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, 
        keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, 
        keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, 
        keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, 
        keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, 
        keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, 
        keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, 
        keyinput_f62, keyinput_f63, keyinput_f64, keyinput_f65, keyinput_f66, 
        keyinput_f67, keyinput_f68, keyinput_f69, keyinput_f70, keyinput_f71, 
        keyinput_f72, keyinput_f73, keyinput_f74, keyinput_f75, keyinput_f76, 
        keyinput_f77, keyinput_f78, keyinput_f79, keyinput_f80, keyinput_f81, 
        keyinput_f82, keyinput_f83, keyinput_f84, keyinput_f85, keyinput_f86, 
        keyinput_f87, keyinput_f88, keyinput_f89, keyinput_f90, keyinput_f91, 
        keyinput_f92, keyinput_f93, keyinput_f94, keyinput_f95, keyinput_f96, 
        keyinput_f97, keyinput_f98, keyinput_f99, keyinput_f100, keyinput_f101, 
        keyinput_f102, keyinput_f103, keyinput_f104, keyinput_f105, 
        keyinput_f106, keyinput_f107, keyinput_f108, keyinput_f109, 
        keyinput_f110, keyinput_f111, keyinput_f112, keyinput_f113, 
        keyinput_f114, keyinput_f115, keyinput_f116, keyinput_f117, 
        keyinput_f118, keyinput_f119, keyinput_f120, keyinput_f121, 
        keyinput_f122, keyinput_f123, keyinput_f124, keyinput_f125, 
        keyinput_f126, keyinput_f127, keyinput_g0, keyinput_g1, keyinput_g2, 
        keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7, 
        keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12, 
        keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17, 
        keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22, 
        keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27, 
        keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32, 
        keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37, 
        keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42, 
        keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47, 
        keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52, 
        keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57, 
        keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62, 
        keyinput_g63, keyinput_g64, keyinput_g65, keyinput_g66, keyinput_g67, 
        keyinput_g68, keyinput_g69, keyinput_g70, keyinput_g71, keyinput_g72, 
        keyinput_g73, keyinput_g74, keyinput_g75, keyinput_g76, keyinput_g77, 
        keyinput_g78, keyinput_g79, keyinput_g80, keyinput_g81, keyinput_g82, 
        keyinput_g83, keyinput_g84, keyinput_g85, keyinput_g86, keyinput_g87, 
        keyinput_g88, keyinput_g89, keyinput_g90, keyinput_g91, keyinput_g92, 
        keyinput_g93, keyinput_g94, keyinput_g95, keyinput_g96, keyinput_g97, 
        keyinput_g98, keyinput_g99, keyinput_g100, keyinput_g101, 
        keyinput_g102, keyinput_g103, keyinput_g104, keyinput_g105, 
        keyinput_g106, keyinput_g107, keyinput_g108, keyinput_g109, 
        keyinput_g110, keyinput_g111, keyinput_g112, keyinput_g113, 
        keyinput_g114, keyinput_g115, keyinput_g116, keyinput_g117, 
        keyinput_g118, keyinput_g119, keyinput_g120, keyinput_g121, 
        keyinput_g122, keyinput_g123, keyinput_g124, keyinput_g125, 
        keyinput_g126, keyinput_g127, U3445, U3446, U3447, U3448, U3213, U3212, 
        U3211, U3210, U3209, U3208, U3207, U3206, U3205, U3204, U3203, U3202, 
        U3201, U3200, U3199, U3198, U3197, U3196, U3195, U3194, U3193, U3192, 
        U3191, U3190, U3189, U3188, U3187, U3186, U3185, U3184, U3183, U3182, 
        U3181, U3451, U3452, U3180, U3179, U3178, U3177, U3176, U3175, U3174, 
        U3173, U3172, U3171, U3170, U3169, U3168, U3167, U3166, U3165, U3164, 
        U3163, U3162, U3161, U3160, U3159, U3158, U3157, U3156, U3155, U3154, 
        U3153, U3152, U3151, U3453, U3150, U3149, U3148, U3147, U3146, U3145, 
        U3144, U3143, U3142, U3141, U3140, U3139, U3138, U3137, U3136, U3135, 
        U3134, U3133, U3132, U3131, U3130, U3129, U3128, U3127, U3126, U3125, 
        U3124, U3123, U3122, U3121, U3120, U3119, U3118, U3117, U3116, U3115, 
        U3114, U3113, U3112, U3111, U3110, U3109, U3108, U3107, U3106, U3105, 
        U3104, U3103, U3102, U3101, U3100, U3099, U3098, U3097, U3096, U3095, 
        U3094, U3093, U3092, U3091, U3090, U3089, U3088, U3087, U3086, U3085, 
        U3084, U3083, U3082, U3081, U3080, U3079, U3078, U3077, U3076, U3075, 
        U3074, U3073, U3072, U3071, U3070, U3069, U3068, U3067, U3066, U3065, 
        U3064, U3063, U3062, U3061, U3060, U3059, U3058, U3057, U3056, U3055, 
        U3054, U3053, U3052, U3051, U3050, U3049, U3048, U3047, U3046, U3045, 
        U3044, U3043, U3042, U3041, U3040, U3039, U3038, U3037, U3036, U3035, 
        U3034, U3033, U3032, U3031, U3030, U3029, U3028, U3027, U3026, U3025, 
        U3024, U3023, U3022, U3021, U3020, U3455, U3456, U3459, U3460, U3461, 
        U3019, U3462, U3463, U3464, U3465, U3018, U3017, U3016, U3015, U3014, 
        U3013, U3012, U3011, U3010, U3009, U3008, U3007, U3006, U3005, U3004, 
        U3003, U3002, U3001, U3000, U2999, U2998, U2997, U2996, U2995, U2994, 
        U2993, U2992, U2991, U2990, U2989, U2988, U2987, U2986, U2985, U2984, 
        U2983, U2982, U2981, U2980, U2979, U2978, U2977, U2976, U2975, U2974, 
        U2973, U2972, U2971, U2970, U2969, U2968, U2967, U2966, U2965, U2964, 
        U2963, U2962, U2961, U2960, U2959, U2958, U2957, U2956, U2955, U2954, 
        U2953, U2952, U2951, U2950, U2949, U2948, U2947, U2946, U2945, U2944, 
        U2943, U2942, U2941, U2940, U2939, U2938, U2937, U2936, U2935, U2934, 
        U2933, U2932, U2931, U2930, U2929, U2928, U2927, U2926, U2925, U2924, 
        U2923, U2922, U2921, U2920, U2919, U2918, U2917, U2916, U2915, U2914, 
        U2913, U2912, U2911, U2910, U2909, U2908, U2907, U2906, U2905, U2904, 
        U2903, U2902, U2901, U2900, U2899, U2898, U2897, U2896, U2895, U2894, 
        U2893, U2892, U2891, U2890, U2889, U2888, U2887, U2886, U2885, U2884, 
        U2883, U2882, U2881, U2880, U2879, U2878, U2877, U2876, U2875, U2874, 
        U2873, U2872, U2871, U2870, U2869, U2868, U2867, U2866, U2865, U2864, 
        U2863, U2862, U2861, U2860, U2859, U2858, U2857, U2856, U2855, U2854, 
        U2853, U2852, U2851, U2850, U2849, U2848, U2847, U2846, U2845, U2844, 
        U2843, U2842, U2841, U2840, U2839, U2838, U2837, U2836, U2835, U2834, 
        U2833, U2832, U2831, U2830, U2829, U2828, U2827, U2826, U2825, U2824, 
        U2823, U2822, U2821, U2820, U2819, U2818, U2817, U2816, U2815, U2814, 
        U2813, U2812, U2811, U2810, U2809, U2808, U2807, U2806, U2805, U2804, 
        U2803, U2802, U2801, U2800, U2799, U2798, U2797, U2796, U2795, U3468, 
        U2794, U3469, U3470, U2793, U3471, U2792, U3472, U2791, U3473, U2790, 
        U2789, U3474, U2788 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
         READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
         M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
         STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
         W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput_f0, keyinput_f1,
         keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6,
         keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11,
         keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16,
         keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21,
         keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26,
         keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31,
         keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36,
         keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41,
         keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46,
         keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51,
         keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56,
         keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61,
         keyinput_f62, keyinput_f63, keyinput_f64, keyinput_f65, keyinput_f66,
         keyinput_f67, keyinput_f68, keyinput_f69, keyinput_f70, keyinput_f71,
         keyinput_f72, keyinput_f73, keyinput_f74, keyinput_f75, keyinput_f76,
         keyinput_f77, keyinput_f78, keyinput_f79, keyinput_f80, keyinput_f81,
         keyinput_f82, keyinput_f83, keyinput_f84, keyinput_f85, keyinput_f86,
         keyinput_f87, keyinput_f88, keyinput_f89, keyinput_f90, keyinput_f91,
         keyinput_f92, keyinput_f93, keyinput_f94, keyinput_f95, keyinput_f96,
         keyinput_f97, keyinput_f98, keyinput_f99, keyinput_f100,
         keyinput_f101, keyinput_f102, keyinput_f103, keyinput_f104,
         keyinput_f105, keyinput_f106, keyinput_f107, keyinput_f108,
         keyinput_f109, keyinput_f110, keyinput_f111, keyinput_f112,
         keyinput_f113, keyinput_f114, keyinput_f115, keyinput_f116,
         keyinput_f117, keyinput_f118, keyinput_f119, keyinput_f120,
         keyinput_f121, keyinput_f122, keyinput_f123, keyinput_f124,
         keyinput_f125, keyinput_f126, keyinput_f127, keyinput_g0, keyinput_g1,
         keyinput_g2, keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6,
         keyinput_g7, keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11,
         keyinput_g12, keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16,
         keyinput_g17, keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21,
         keyinput_g22, keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26,
         keyinput_g27, keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31,
         keyinput_g32, keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36,
         keyinput_g37, keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41,
         keyinput_g42, keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46,
         keyinput_g47, keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51,
         keyinput_g52, keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56,
         keyinput_g57, keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61,
         keyinput_g62, keyinput_g63, keyinput_g64, keyinput_g65, keyinput_g66,
         keyinput_g67, keyinput_g68, keyinput_g69, keyinput_g70, keyinput_g71,
         keyinput_g72, keyinput_g73, keyinput_g74, keyinput_g75, keyinput_g76,
         keyinput_g77, keyinput_g78, keyinput_g79, keyinput_g80, keyinput_g81,
         keyinput_g82, keyinput_g83, keyinput_g84, keyinput_g85, keyinput_g86,
         keyinput_g87, keyinput_g88, keyinput_g89, keyinput_g90, keyinput_g91,
         keyinput_g92, keyinput_g93, keyinput_g94, keyinput_g95, keyinput_g96,
         keyinput_g97, keyinput_g98, keyinput_g99, keyinput_g100,
         keyinput_g101, keyinput_g102, keyinput_g103, keyinput_g104,
         keyinput_g105, keyinput_g106, keyinput_g107, keyinput_g108,
         keyinput_g109, keyinput_g110, keyinput_g111, keyinput_g112,
         keyinput_g113, keyinput_g114, keyinput_g115, keyinput_g116,
         keyinput_g117, keyinput_g118, keyinput_g119, keyinput_g120,
         keyinput_g121, keyinput_g122, keyinput_g123, keyinput_g124,
         keyinput_g125, keyinput_g126, keyinput_g127;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4027, n4028, n4029, n4030, n4031, n4032, n4033,
         n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043,
         n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053,
         n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063,
         n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073,
         n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083,
         n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093,
         n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103,
         n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113,
         n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123,
         n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133,
         n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143,
         n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153,
         n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163,
         n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173,
         n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183,
         n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193,
         n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203,
         n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213,
         n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223,
         n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233,
         n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243,
         n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253,
         n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263,
         n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273,
         n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283,
         n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293,
         n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303,
         n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313,
         n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323,
         n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333,
         n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343,
         n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353,
         n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363,
         n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373,
         n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383,
         n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393,
         n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403,
         n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413,
         n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423,
         n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433,
         n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443,
         n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453,
         n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463,
         n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473,
         n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483,
         n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493,
         n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503,
         n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513,
         n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523,
         n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533,
         n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543,
         n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553,
         n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563,
         n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573,
         n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583,
         n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593,
         n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603,
         n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613,
         n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623,
         n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633,
         n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643,
         n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653,
         n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663,
         n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673,
         n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683,
         n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693,
         n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703,
         n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713,
         n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723,
         n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733,
         n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743,
         n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753,
         n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763,
         n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773,
         n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783,
         n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793,
         n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803,
         n4804, n4805, n4806, n4807, n4808, n4810, n4811, n4812, n4813, n4814,
         n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824,
         n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834,
         n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844,
         n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854,
         n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864,
         n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874,
         n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884,
         n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894,
         n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904,
         n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914,
         n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924,
         n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934,
         n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944,
         n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954,
         n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964,
         n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974,
         n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984,
         n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994,
         n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004,
         n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014,
         n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024,
         n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034,
         n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044,
         n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054,
         n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064,
         n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074,
         n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084,
         n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094,
         n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104,
         n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114,
         n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124,
         n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134,
         n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144,
         n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154,
         n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164,
         n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174,
         n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184,
         n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194,
         n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204,
         n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214,
         n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224,
         n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234,
         n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244,
         n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254,
         n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264,
         n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274,
         n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284,
         n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294,
         n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304,
         n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314,
         n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324,
         n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334,
         n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344,
         n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354,
         n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364,
         n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374,
         n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384,
         n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394,
         n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404,
         n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414,
         n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424,
         n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434,
         n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444,
         n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454,
         n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464,
         n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474,
         n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484,
         n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494,
         n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504,
         n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514,
         n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524,
         n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534,
         n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544,
         n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554,
         n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564,
         n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574,
         n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584,
         n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594,
         n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604,
         n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614,
         n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624,
         n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634,
         n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644,
         n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654,
         n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664,
         n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674,
         n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684,
         n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694,
         n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704,
         n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714,
         n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724,
         n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734,
         n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744,
         n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754,
         n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764,
         n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774,
         n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784,
         n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794,
         n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804,
         n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814,
         n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824,
         n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834,
         n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844,
         n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854,
         n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864,
         n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874,
         n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884,
         n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894,
         n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904,
         n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914,
         n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924,
         n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934,
         n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944,
         n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954,
         n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964,
         n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974,
         n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984,
         n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994,
         n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004,
         n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014,
         n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024,
         n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034,
         n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044,
         n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054,
         n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064,
         n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074,
         n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084,
         n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094,
         n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104,
         n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114,
         n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124,
         n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134,
         n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144,
         n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154,
         n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164,
         n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174,
         n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184,
         n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194,
         n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204,
         n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214,
         n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224,
         n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234,
         n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244,
         n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254,
         n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264,
         n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274,
         n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284,
         n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294,
         n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304,
         n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314,
         n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324,
         n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334,
         n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344,
         n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354,
         n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364,
         n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374,
         n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384,
         n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394,
         n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404,
         n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414,
         n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424,
         n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434,
         n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444,
         n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454,
         n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464,
         n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474,
         n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484,
         n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494,
         n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504,
         n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514,
         n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524,
         n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534,
         n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544,
         n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554,
         n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564,
         n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574,
         n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584,
         n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594,
         n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604,
         n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614,
         n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624,
         n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634,
         n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644,
         n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654,
         n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664,
         n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674,
         n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684,
         n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694,
         n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704,
         n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714,
         n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724,
         n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734,
         n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744,
         n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754,
         n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764,
         n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774,
         n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784,
         n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794,
         n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804,
         n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814,
         n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824,
         n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834,
         n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844,
         n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854,
         n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864,
         n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874,
         n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884,
         n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894,
         n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904,
         n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914,
         n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924,
         n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934,
         n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944,
         n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954,
         n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964,
         n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974,
         n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984,
         n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994,
         n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004,
         n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014,
         n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024,
         n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034,
         n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044,
         n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054,
         n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064,
         n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074,
         n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084,
         n7085, n7086, n7087;

  BUF_X1 U3601 ( .A(n4092), .Z(n4093) );
  OAI21_X1 U3602 ( .B1(n4422), .B2(STATE2_REG_0__SCAN_IN), .A(n3431), .ZN(
        n3436) );
  CLKBUF_X2 U3603 ( .A(n3972), .Z(n4000) );
  CLKBUF_X2 U3604 ( .A(n3990), .Z(n3926) );
  CLKBUF_X2 U3605 ( .A(n3420), .Z(n3989) );
  CLKBUF_X2 U3606 ( .A(n3370), .Z(n3991) );
  CLKBUF_X2 U3607 ( .A(n3391), .Z(n3992) );
  CLKBUF_X2 U3608 ( .A(n3362), .Z(n3921) );
  NAND2_X2 U3610 ( .A1(n3256), .A2(n3255), .ZN(n4676) );
  AND2_X2 U3611 ( .A1(n3195), .A2(n4430), .ZN(n3972) );
  CLKBUF_X1 U3612 ( .A(n3827), .Z(n3153) );
  NOR2_X1 U3613 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATEBS16_REG_SCAN_IN), .ZN(
        n3827) );
  NAND2_X1 U3614 ( .A1(n3323), .A2(n3307), .ZN(n3308) );
  AND2_X2 U3615 ( .A1(n4538), .A2(n4431), .ZN(n3293) );
  OAI21_X1 U3616 ( .B1(n4650), .B2(n3655), .A(n3720), .ZN(n3475) );
  INV_X1 U3617 ( .A(n4668), .ZN(n4327) );
  XNOR2_X1 U3618 ( .A(n3380), .B(n3379), .ZN(n3440) );
  AOI211_X1 U3621 ( .C1(n4399), .C2(n4398), .A(n4400), .B(n4397), .ZN(n4404)
         );
  NAND2_X1 U3622 ( .A1(n4968), .A2(n3660), .ZN(n5358) );
  NAND2_X1 U3623 ( .A1(n5833), .A2(n5825), .ZN(n5827) );
  INV_X1 U3624 ( .A(n6247), .ZN(n6272) );
  AND2_X1 U3625 ( .A1(n3356), .A2(n3335), .ZN(n3154) );
  AND2_X1 U3626 ( .A1(n3440), .A2(n3441), .ZN(n3155) );
  AND2_X1 U3627 ( .A1(n4092), .A2(n4327), .ZN(n3156) );
  NAND2_X2 U3628 ( .A1(n3214), .A2(n3213), .ZN(n3318) );
  AND2_X2 U3629 ( .A1(n3333), .A2(n3330), .ZN(n3328) );
  BUF_X2 U3630 ( .A(n3235), .Z(n3323) );
  AND2_X4 U3631 ( .A1(n3197), .A2(n4538), .ZN(n3264) );
  AND2_X2 U3632 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n3189), .ZN(n3197)
         );
  AND2_X1 U3633 ( .A1(n3196), .A2(n3195), .ZN(n3157) );
  NAND4_X4 U3634 ( .A1(n3290), .A2(n3289), .A3(n3288), .A4(n3287), .ZN(n4094)
         );
  AND4_X2 U3635 ( .A1(n3282), .A2(n3281), .A3(n3280), .A4(n3279), .ZN(n3288)
         );
  AND2_X1 U3636 ( .A1(n4538), .A2(n4431), .ZN(n3158) );
  NOR2_X2 U3637 ( .A1(n4332), .A2(n3258), .ZN(n3340) );
  NAND2_X2 U3638 ( .A1(n3303), .A2(n3302), .ZN(n4668) );
  NAND2_X2 U3639 ( .A1(n3321), .A2(n4348), .ZN(n4030) );
  NAND2_X2 U3640 ( .A1(n3155), .A2(n3500), .ZN(n3533) );
  NAND2_X2 U3641 ( .A1(n5476), .A2(n5475), .ZN(n5497) );
  NAND2_X1 U3642 ( .A1(n5622), .A2(n3180), .ZN(n5874) );
  NAND2_X1 U3643 ( .A1(n4316), .A2(n6004), .ZN(n6001) );
  NAND2_X1 U3644 ( .A1(n4297), .A2(n4296), .ZN(n5476) );
  AND2_X1 U3645 ( .A1(n5336), .A2(n5363), .ZN(n5361) );
  NOR2_X1 U3646 ( .A1(n4969), .A2(n3659), .ZN(n3660) );
  AOI21_X1 U3647 ( .B1(n4275), .B2(n3704), .A(n3580), .ZN(n4969) );
  INV_X4 U3648 ( .A(n4664), .ZN(n3321) );
  OR2_X2 U3649 ( .A1(n3245), .A2(n3244), .ZN(n3324) );
  CLKBUF_X2 U3650 ( .A(n3259), .Z(n3399) );
  AOI21_X1 U3651 ( .B1(n5864), .B2(INSTADDRPOINTER_REG_29__SCAN_IN), .A(n5624), 
        .ZN(n5625) );
  AOI21_X1 U3652 ( .B1(n5732), .B2(n6357), .A(n5728), .ZN(n5729) );
  AOI211_X1 U3653 ( .C1(n6144), .C2(n5673), .A(n5655), .B(n5654), .ZN(n5656)
         );
  NOR2_X1 U3654 ( .A1(n5903), .A2(n5904), .ZN(n5902) );
  AOI21_X1 U3655 ( .B1(n5771), .B2(n5769), .A(n5770), .ZN(n5871) );
  OR2_X1 U3656 ( .A1(n5823), .A2(n5652), .ZN(n5653) );
  CLKBUF_X1 U3657 ( .A(n5651), .Z(n5823) );
  NAND2_X1 U3658 ( .A1(n3920), .A2(n3185), .ZN(n5820) );
  AND2_X1 U3659 ( .A1(n4407), .A2(n4406), .ZN(n4408) );
  INV_X1 U3660 ( .A(n5766), .ZN(n5636) );
  OR2_X1 U3661 ( .A1(n5779), .A2(n5778), .ZN(n5935) );
  OAI21_X1 U3662 ( .B1(n4398), .B2(n5776), .A(n3177), .ZN(n5779) );
  XNOR2_X1 U3663 ( .A(n4285), .B(n3574), .ZN(n4275) );
  NOR2_X1 U3664 ( .A1(n4881), .A2(n5237), .ZN(n6436) );
  CLKBUF_X1 U3665 ( .A(n4650), .Z(n6025) );
  AND2_X1 U3666 ( .A1(n4509), .A2(n4511), .ZN(n3474) );
  AND2_X1 U3667 ( .A1(n3439), .A2(n3438), .ZN(n3441) );
  AND2_X1 U3668 ( .A1(n3499), .A2(n3498), .ZN(n4998) );
  CLKBUF_X1 U3669 ( .A(n4547), .Z(n5237) );
  CLKBUF_X1 U3670 ( .A(n4517), .Z(n5414) );
  AOI21_X1 U3671 ( .B1(n3418), .B2(n3457), .A(n3417), .ZN(n3446) );
  NOR2_X1 U3672 ( .A1(n7014), .A2(n4926), .ZN(n6462) );
  NAND2_X1 U3673 ( .A1(n3453), .A2(n3456), .ZN(n3418) );
  CLKBUF_X1 U3675 ( .A(n4422), .Z(n6023) );
  NAND2_X1 U3676 ( .A1(n4644), .A2(n4645), .ZN(n4760) );
  NAND2_X1 U3677 ( .A1(n3484), .A2(n3483), .ZN(n6445) );
  AOI21_X1 U3678 ( .B1(n3479), .B2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(n3354), 
        .ZN(n3357) );
  NAND2_X1 U3679 ( .A1(n4321), .A2(n4986), .ZN(n5754) );
  CLKBUF_X1 U3680 ( .A(n4321), .Z(n4423) );
  CLKBUF_X1 U3681 ( .A(n3315), .Z(n4333) );
  BUF_X2 U3682 ( .A(n3343), .Z(n4413) );
  AND2_X1 U3683 ( .A1(n4612), .A2(n4672), .ZN(n3258) );
  AND2_X1 U3684 ( .A1(n3318), .A2(n3324), .ZN(n5491) );
  NAND2_X1 U3685 ( .A1(n3270), .A2(n4392), .ZN(n3315) );
  BUF_X2 U3686 ( .A(n4098), .Z(n5597) );
  NAND2_X1 U3687 ( .A1(n3160), .A2(n4023), .ZN(n4425) );
  OR2_X1 U3688 ( .A1(n3398), .A2(n3397), .ZN(n4279) );
  AND2_X1 U3689 ( .A1(n3324), .A2(n3305), .ZN(n3270) );
  BUF_X2 U3690 ( .A(n3323), .Z(n5492) );
  CLKBUF_X1 U3691 ( .A(n3321), .Z(n4417) );
  AND2_X2 U3692 ( .A1(n4664), .A2(n3323), .ZN(n4023) );
  INV_X1 U3693 ( .A(n3305), .ZN(n4672) );
  AND4_X2 U3694 ( .A1(n3234), .A2(n3233), .A3(n3232), .A4(n3231), .ZN(n3305)
         );
  OR2_X1 U3695 ( .A1(n3204), .A2(n3203), .ZN(n3235) );
  AND4_X1 U3696 ( .A1(n3208), .A2(n3207), .A3(n3206), .A4(n3205), .ZN(n3214)
         );
  AND4_X1 U3697 ( .A1(n3286), .A2(n3285), .A3(n3284), .A4(n3283), .ZN(n3287)
         );
  AND4_X1 U3698 ( .A1(n3278), .A2(n3277), .A3(n3276), .A4(n3275), .ZN(n3289)
         );
  AND4_X1 U3699 ( .A1(n3274), .A2(n3273), .A3(n3272), .A4(n3271), .ZN(n3290)
         );
  AND4_X1 U3700 ( .A1(n3268), .A2(n3267), .A3(n3266), .A4(n3265), .ZN(n3269)
         );
  AND4_X1 U3701 ( .A1(n3263), .A2(n3262), .A3(n3261), .A4(n3260), .ZN(n3179)
         );
  AND4_X1 U3702 ( .A1(n3212), .A2(n3211), .A3(n3210), .A4(n3209), .ZN(n3213)
         );
  AND4_X1 U3703 ( .A1(n3226), .A2(n3225), .A3(n3224), .A4(n3223), .ZN(n3232)
         );
  NAND2_X2 U3704 ( .A1(n6648), .A2(n7040), .ZN(n6655) );
  AND4_X1 U3705 ( .A1(n3218), .A2(n3217), .A3(n3216), .A4(n3215), .ZN(n3234)
         );
  AND4_X1 U3706 ( .A1(n3301), .A2(n3300), .A3(n3299), .A4(n3298), .ZN(n3302)
         );
  AND4_X1 U3707 ( .A1(n3250), .A2(n3249), .A3(n3248), .A4(n3247), .ZN(n3256)
         );
  NAND2_X2 U3708 ( .A1(STATE_REG_2__SCAN_IN), .A2(n6648), .ZN(n6654) );
  AND4_X1 U3709 ( .A1(n3297), .A2(n3296), .A3(n3295), .A4(n3294), .ZN(n3303)
         );
  AND4_X1 U3710 ( .A1(n3222), .A2(n3221), .A3(n3220), .A4(n3219), .ZN(n3233)
         );
  BUF_X2 U3711 ( .A(n3363), .Z(n3971) );
  BUF_X2 U3712 ( .A(n3264), .Z(n3836) );
  BUF_X2 U3713 ( .A(n3405), .Z(n3999) );
  BUF_X2 U3714 ( .A(n3404), .Z(n3997) );
  CLKBUF_X2 U3715 ( .A(n3487), .Z(n3386) );
  AND2_X2 U3716 ( .A1(n3196), .A2(n3195), .ZN(n3392) );
  BUF_X2 U3717 ( .A(n3364), .Z(n3988) );
  AND2_X2 U3718 ( .A1(n3196), .A2(n4538), .ZN(n3363) );
  AND2_X2 U3719 ( .A1(n4430), .A2(n4538), .ZN(n3370) );
  NOR2_X2 U3720 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3195) );
  AND2_X1 U3721 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4518) );
  NOR2_X1 U3722 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3190) );
  INV_X1 U3723 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3187) );
  NOR2_X2 U3725 ( .A1(n5208), .A2(n5209), .ZN(n4974) );
  AND2_X1 U3726 ( .A1(n4295), .A2(n3169), .ZN(n3159) );
  NOR2_X2 U3727 ( .A1(n5332), .A2(n5333), .ZN(n5312) );
  OR2_X2 U3728 ( .A1(n3462), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3453) );
  AND2_X1 U3729 ( .A1(n4676), .A2(n3305), .ZN(n3160) );
  NAND2_X1 U3730 ( .A1(n4023), .A2(n3305), .ZN(n3161) );
  BUF_X1 U3731 ( .A(n3292), .Z(n3162) );
  NAND2_X1 U3732 ( .A1(n4078), .A2(n4417), .ZN(n3163) );
  NAND2_X1 U3733 ( .A1(n4078), .A2(n4417), .ZN(n4344) );
  AND3_X2 U3734 ( .A1(n3320), .A2(n3319), .A3(n3342), .ZN(n4078) );
  AND2_X1 U3735 ( .A1(n4240), .A2(n4239), .ZN(n6354) );
  XNOR2_X1 U3736 ( .A(n3448), .B(n3447), .ZN(n4651) );
  XNOR2_X1 U3737 ( .A(n3446), .B(n3445), .ZN(n3448) );
  NAND2_X1 U3738 ( .A1(n3356), .A2(n3335), .ZN(n3164) );
  INV_X1 U3739 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3165) );
  NAND2_X1 U3740 ( .A1(n4308), .A2(n4307), .ZN(n3166) );
  NAND2_X1 U3741 ( .A1(n4308), .A2(n4307), .ZN(n5537) );
  BUF_X1 U3742 ( .A(n4215), .Z(n4650) );
  NOR2_X2 U3743 ( .A1(n4104), .A2(n4103), .ZN(n4639) );
  NOR2_X2 U3744 ( .A1(n4760), .A2(n4761), .ZN(n4803) );
  NAND2_X1 U3745 ( .A1(n3440), .A2(n3441), .ZN(n3167) );
  NAND2_X1 U3746 ( .A1(n6338), .A2(n3171), .ZN(n3168) );
  AND2_X1 U3747 ( .A1(n3168), .A2(n3169), .ZN(n5387) );
  OR2_X1 U3748 ( .A1(n3170), .A2(n5187), .ZN(n3169) );
  INV_X1 U3749 ( .A(n4293), .ZN(n3170) );
  AND2_X1 U3750 ( .A1(n4284), .A2(n4293), .ZN(n3171) );
  XNOR2_X1 U3751 ( .A(n3419), .B(n3164), .ZN(n4422) );
  AND2_X1 U3752 ( .A1(n3316), .A2(n3320), .ZN(n4321) );
  AND2_X1 U3753 ( .A1(n3198), .A2(n4431), .ZN(n3172) );
  AND2_X1 U3754 ( .A1(n3198), .A2(n4431), .ZN(n3259) );
  NAND2_X1 U3755 ( .A1(n3291), .A2(n3318), .ZN(n4392) );
  XNOR2_X1 U3756 ( .A(n3533), .B(n3534), .ZN(n4249) );
  NAND2_X1 U3757 ( .A1(n4220), .A2(n4219), .ZN(n6363) );
  AND2_X1 U3758 ( .A1(n4430), .A2(n4538), .ZN(n3173) );
  NAND2_X1 U3759 ( .A1(n4285), .A2(n4288), .ZN(n3174) );
  NOR2_X2 U3760 ( .A1(n5408), .A2(n5409), .ZN(n5407) );
  AND2_X4 U3761 ( .A1(n3196), .A2(n3198), .ZN(n3487) );
  AND2_X1 U3762 ( .A1(n5694), .A2(n5840), .ZN(n5788) );
  NAND2_X1 U3763 ( .A1(n3381), .A2(n3382), .ZN(n3419) );
  NAND2_X1 U3764 ( .A1(n3350), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3329) );
  AND2_X1 U3765 ( .A1(n3901), .A2(n3900), .ZN(n5787) );
  OR2_X1 U3766 ( .A1(n4294), .A2(n4306), .ZN(n4307) );
  INV_X1 U3767 ( .A(n3377), .ZN(n4241) );
  NAND2_X1 U3768 ( .A1(n4327), .A2(n4676), .ZN(n4352) );
  NAND2_X1 U3769 ( .A1(n4348), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3486) );
  NOR2_X2 U3770 ( .A1(n5820), .A2(n5822), .ZN(n5651) );
  INV_X1 U3771 ( .A(n4009), .ZN(n3983) );
  INV_X1 U3772 ( .A(n4019), .ZN(n3776) );
  AND2_X1 U3773 ( .A1(n5329), .A2(n5328), .ZN(n5355) );
  INV_X1 U3774 ( .A(n3153), .ZN(n4012) );
  INV_X1 U3775 ( .A(n3776), .ZN(n4014) );
  INV_X1 U3776 ( .A(n3655), .ZN(n3704) );
  NAND2_X1 U3777 ( .A1(n3154), .A2(n3419), .ZN(n3360) );
  AND3_X1 U3778 ( .A1(n4986), .A2(n4672), .A3(STATE2_REG_0__SCAN_IN), .ZN(
        n4062) );
  NAND2_X1 U3779 ( .A1(n3486), .A2(n3485), .ZN(n4074) );
  XNOR2_X1 U3780 ( .A(n4457), .B(n6445), .ZN(n4517) );
  OR3_X1 U3781 ( .A1(n5756), .A2(n6598), .A3(n5754), .ZN(n4419) );
  INV_X1 U3782 ( .A(n3720), .ZN(n4018) );
  NOR2_X1 U3783 ( .A1(n3962), .A2(n5650), .ZN(n3963) );
  CLKBUF_X1 U3784 ( .A(n5788), .Z(n5789) );
  CLKBUF_X1 U3785 ( .A(n5790), .Z(n5791) );
  INV_X1 U3786 ( .A(n5604), .ZN(n5850) );
  CLKBUF_X1 U3787 ( .A(n5603), .Z(n5604) );
  NOR2_X1 U3788 ( .A1(n3688), .A2(n5302), .ZN(n3692) );
  NAND2_X1 U3789 ( .A1(n3531), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3576)
         );
  NAND2_X1 U3790 ( .A1(n5705), .A2(n5621), .ZN(n5646) );
  AND2_X1 U3791 ( .A1(n5598), .A2(n4156), .ZN(n5609) );
  NOR2_X2 U3792 ( .A1(n6165), .A2(n5533), .ZN(n5598) );
  OR2_X1 U3793 ( .A1(n5553), .A2(n4302), .ZN(n4303) );
  AND2_X1 U3794 ( .A1(n5727), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4983) );
  OR2_X1 U3795 ( .A1(n5636), .A2(n6288), .ZN(n4407) );
  XNOR2_X1 U3796 ( .A(n5770), .B(n4390), .ZN(n5855) );
  INV_X1 U3797 ( .A(n4389), .ZN(n4390) );
  NAND2_X1 U3798 ( .A1(n5714), .A2(n5726), .ZN(n5715) );
  AOI21_X1 U3799 ( .B1(n5779), .B2(n4400), .A(n4397), .ZN(n4197) );
  CLKBUF_X1 U3800 ( .A(n3392), .Z(n3998) );
  CLKBUF_X1 U3801 ( .A(n3603), .Z(n3885) );
  INV_X1 U3802 ( .A(n3318), .ZN(n3307) );
  OR2_X1 U3803 ( .A1(n3564), .A2(n3563), .ZN(n4277) );
  OR2_X1 U3804 ( .A1(n3545), .A2(n3544), .ZN(n4266) );
  OR2_X1 U3805 ( .A1(n3519), .A2(n3518), .ZN(n4267) );
  INV_X1 U3806 ( .A(n4227), .ZN(n3434) );
  OR2_X1 U3807 ( .A1(n3376), .A2(n3375), .ZN(n3377) );
  INV_X2 U3808 ( .A(n4094), .ZN(n4348) );
  INV_X1 U3809 ( .A(n5790), .ZN(n3920) );
  NAND2_X1 U3810 ( .A1(n4636), .A2(n4635), .ZN(n3477) );
  OR2_X1 U3811 ( .A1(n4102), .A2(n4185), .ZN(n4142) );
  INV_X1 U3812 ( .A(n4182), .ZN(n4166) );
  INV_X1 U3813 ( .A(n4142), .ZN(n4134) );
  INV_X1 U3814 ( .A(n4194), .ZN(n4174) );
  NAND2_X1 U3815 ( .A1(n4102), .A2(n5597), .ZN(n4182) );
  NOR2_X1 U3816 ( .A1(n4352), .A2(n3323), .ZN(n3316) );
  NAND2_X1 U3817 ( .A1(n3337), .A2(n3336), .ZN(n3381) );
  AOI21_X1 U3818 ( .B1(n3348), .B2(n4664), .A(n3347), .ZN(n3349) );
  NAND2_X1 U3819 ( .A1(n3443), .A2(n3442), .ZN(n3444) );
  INV_X1 U3820 ( .A(n3440), .ZN(n3443) );
  NAND2_X1 U3821 ( .A1(n3360), .A2(n3359), .ZN(n3478) );
  OR2_X1 U3822 ( .A1(n4612), .A2(n3708), .ZN(n4429) );
  AND2_X1 U3823 ( .A1(n4428), .A2(n4357), .ZN(n4521) );
  AND2_X2 U3824 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4430) );
  INV_X1 U3825 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n5243) );
  AND2_X1 U3826 ( .A1(n3480), .A2(n4654), .ZN(n4925) );
  OAI21_X1 U3827 ( .B1(n6680), .B2(n4545), .A(n5738), .ZN(n4658) );
  INV_X1 U3828 ( .A(n4652), .ZN(n5089) );
  INV_X1 U3829 ( .A(n4413), .ZN(n6679) );
  NOR2_X2 U3830 ( .A1(n5774), .A2(n5775), .ZN(n4401) );
  OR2_X1 U3831 ( .A1(n4205), .A2(n5296), .ZN(n5467) );
  NOR2_X1 U3832 ( .A1(n3623), .A2(n6241), .ZN(n3661) );
  OR2_X1 U3833 ( .A1(n6675), .A2(n4086), .ZN(n5372) );
  OR2_X1 U3834 ( .A1(n6036), .A2(n4012), .ZN(n3943) );
  INV_X1 U3835 ( .A(n6335), .ZN(n4465) );
  NOR2_X1 U3836 ( .A1(n3324), .A2(n6590), .ZN(n4019) );
  NAND2_X1 U3837 ( .A1(n3939), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n3941)
         );
  OR2_X1 U3838 ( .A1(n3941), .A2(n3940), .ZN(n3962) );
  CLKBUF_X1 U3839 ( .A(n5820), .Z(n5821) );
  OR2_X1 U3840 ( .A1(n3896), .A2(n3895), .ZN(n3897) );
  NOR2_X1 U3841 ( .A1(n3857), .A2(n5898), .ZN(n3858) );
  OR2_X1 U3842 ( .A1(n5810), .A2(n4012), .ZN(n3860) );
  CLKBUF_X1 U3843 ( .A(n5694), .Z(n5695) );
  CLKBUF_X1 U3844 ( .A(n5696), .Z(n5697) );
  AND2_X1 U3845 ( .A1(PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n3810), .ZN(n3811)
         );
  NAND2_X1 U3846 ( .A1(n3811), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n3857)
         );
  NOR2_X1 U3847 ( .A1(n3762), .A2(n6212), .ZN(n3763) );
  CLKBUF_X1 U3848 ( .A(n5529), .Z(n5530) );
  CLKBUF_X1 U3849 ( .A(n5525), .Z(n5526) );
  AND2_X1 U3850 ( .A1(n3740), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3741)
         );
  CLKBUF_X1 U3851 ( .A(n5523), .Z(n5524) );
  CLKBUF_X1 U3852 ( .A(n5461), .Z(n5462) );
  CLKBUF_X1 U3853 ( .A(n5361), .Z(n5362) );
  NAND2_X1 U3854 ( .A1(n3692), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n3707)
         );
  NAND2_X1 U3855 ( .A1(n3677), .A2(n3676), .ZN(n5338) );
  AND3_X1 U3856 ( .A1(n3691), .A2(n3690), .A3(n3689), .ZN(n5339) );
  CLKBUF_X1 U3857 ( .A(n5336), .Z(n5337) );
  NAND2_X1 U3858 ( .A1(n3661), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3688)
         );
  CLKBUF_X1 U3859 ( .A(n5179), .Z(n5180) );
  NAND2_X1 U3860 ( .A1(n3627), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3623)
         );
  NAND2_X1 U3861 ( .A1(n3595), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3652)
         );
  INV_X1 U3862 ( .A(n3594), .ZN(n3595) );
  NOR2_X1 U3863 ( .A1(n4972), .A2(n4973), .ZN(n5329) );
  NOR2_X1 U3864 ( .A1(n3576), .A2(n3575), .ZN(n3577) );
  INV_X1 U3865 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3575) );
  CLKBUF_X1 U3866 ( .A(n4969), .Z(n4970) );
  OAI211_X1 U3867 ( .C1(n3550), .C2(n4012), .A(n3549), .B(n3548), .ZN(n4733)
         );
  NOR2_X1 U3868 ( .A1(n3526), .A2(n5290), .ZN(n3531) );
  INV_X1 U3869 ( .A(n3502), .ZN(n3503) );
  NAND2_X1 U3870 ( .A1(n3508), .A2(n3507), .ZN(n4701) );
  NAND2_X1 U3871 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3502) );
  CLKBUF_X1 U3872 ( .A(n4634), .Z(n4702) );
  NAND2_X1 U3873 ( .A1(n4491), .A2(n4490), .ZN(n4489) );
  AND2_X1 U3874 ( .A1(n6156), .A2(n5631), .ZN(n5940) );
  OAI21_X1 U3875 ( .B1(n6000), .B2(n5618), .A(n4294), .ZN(n5619) );
  AND2_X1 U3876 ( .A1(n4149), .A2(n4148), .ZN(n5533) );
  CLKBUF_X1 U3877 ( .A(n5913), .Z(n5914) );
  AND2_X1 U3878 ( .A1(n5554), .A2(n4304), .ZN(n5563) );
  NOR2_X2 U3879 ( .A1(n5182), .A2(n5183), .ZN(n5342) );
  AND2_X1 U3880 ( .A1(n5498), .A2(n4299), .ZN(n4300) );
  OR2_X1 U3881 ( .A1(n4294), .A2(n5573), .ZN(n4299) );
  NAND2_X1 U3882 ( .A1(n5312), .A2(n5313), .ZN(n5408) );
  OR2_X1 U3883 ( .A1(n4294), .A2(n4298), .ZN(n5498) );
  NAND2_X1 U3884 ( .A1(n4974), .A2(n4975), .ZN(n5332) );
  AND2_X1 U3885 ( .A1(n4360), .A2(n4481), .ZN(n5195) );
  NAND2_X1 U3886 ( .A1(n4803), .A2(n4804), .ZN(n5208) );
  AND2_X1 U3887 ( .A1(n4185), .A2(n5597), .ZN(n4483) );
  NOR2_X1 U3888 ( .A1(n4375), .A2(n5661), .ZN(n5577) );
  NAND2_X1 U3889 ( .A1(n4517), .A2(n6596), .ZN(n3499) );
  INV_X1 U3890 ( .A(n5238), .ZN(n6486) );
  INV_X1 U3891 ( .A(n4926), .ZN(n4820) );
  NAND2_X1 U3892 ( .A1(n4076), .A2(n4075), .ZN(n5756) );
  NOR2_X1 U3893 ( .A1(n6025), .A2(n3500), .ZN(n6028) );
  NOR2_X1 U3894 ( .A1(n6486), .A2(n4652), .ZN(n4860) );
  AND2_X1 U3895 ( .A1(n5240), .A2(n5414), .ZN(n6488) );
  NOR2_X1 U3896 ( .A1(n4734), .A2(n4652), .ZN(n4736) );
  NAND2_X1 U3897 ( .A1(n6596), .A2(n4658), .ZN(n4926) );
  OR2_X1 U3898 ( .A1(n4734), .A2(n5089), .ZN(n4660) );
  INV_X1 U3899 ( .A(n6496), .ZN(n6455) );
  OR3_X1 U3900 ( .A1(n6043), .A2(n7057), .A3(n7009), .ZN(n5763) );
  INV_X1 U3901 ( .A(n6276), .ZN(n6242) );
  AND2_X1 U3902 ( .A1(n6675), .A2(n4200), .ZN(n6277) );
  AND2_X1 U3903 ( .A1(n6231), .A2(n5372), .ZN(n6091) );
  INV_X1 U3904 ( .A(n6288), .ZN(n5846) );
  NAND2_X1 U3905 ( .A1(n6292), .A2(n5731), .ZN(n6288) );
  AND2_X1 U3906 ( .A1(n5860), .A2(n4613), .ZN(n6297) );
  INV_X1 U3907 ( .A(n5860), .ZN(n6299) );
  INV_X1 U3908 ( .A(n5861), .ZN(n6300) );
  NAND2_X1 U3909 ( .A1(n4611), .A2(n4610), .ZN(n5860) );
  XNOR2_X1 U3911 ( .A(n4090), .B(n4089), .ZN(n5727) );
  INV_X1 U3912 ( .A(n6039), .ZN(n6101) );
  OAI21_X1 U3913 ( .B1(n5829), .B2(n3185), .A(n5821), .ZN(n6047) );
  AOI21_X1 U3914 ( .B1(n5793), .B2(n5792), .A(n5829), .ZN(n6129) );
  INV_X1 U3915 ( .A(n5890), .ZN(n6106) );
  AND2_X1 U3916 ( .A1(n5406), .A2(n5405), .ZN(n6248) );
  INV_X1 U3917 ( .A(n6370), .ZN(n6144) );
  INV_X1 U3918 ( .A(n6148), .ZN(n6361) );
  NAND2_X1 U3919 ( .A1(n6148), .A2(n4513), .ZN(n6370) );
  INV_X1 U3920 ( .A(n6195), .ZN(n6366) );
  CLKBUF_X1 U3921 ( .A(n5646), .Z(n5881) );
  OR2_X1 U3922 ( .A1(n4375), .A2(n5752), .ZN(n5687) );
  INV_X1 U3923 ( .A(n6398), .ZN(n6418) );
  AND2_X1 U3924 ( .A1(n5199), .A2(n4573), .ZN(n6420) );
  INV_X1 U3925 ( .A(n6395), .ZN(n6412) );
  OR2_X1 U3926 ( .A1(n5199), .A2(n6414), .ZN(n5633) );
  INV_X1 U3927 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6558) );
  CLKBUF_X1 U3928 ( .A(n3462), .Z(n3463) );
  CLKBUF_X1 U3929 ( .A(n4651), .Z(n4652) );
  INV_X1 U3930 ( .A(n6021), .ZN(n6485) );
  CLKBUF_X1 U3931 ( .A(n4526), .Z(n4527) );
  INV_X1 U3932 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3188) );
  OR2_X1 U3933 ( .A1(n5756), .A2(n6666), .ZN(n5738) );
  NOR2_X1 U3934 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_3__SCAN_IN), .ZN(
        n6597) );
  INV_X1 U3935 ( .A(n6443), .ZN(n4794) );
  INV_X1 U3936 ( .A(n6436), .ZN(n5090) );
  NOR2_X1 U3937 ( .A1(n5137), .A2(n5138), .ZN(n5127) );
  AND2_X1 U3938 ( .A1(n6028), .A2(n5419), .ZN(n6479) );
  NAND2_X1 U3939 ( .A1(n4860), .A2(n5138), .ZN(n5248) );
  NAND2_X1 U3940 ( .A1(n5238), .A2(n4999), .ZN(n6527) );
  INV_X1 U3941 ( .A(n5257), .ZN(n6506) );
  INV_X1 U3942 ( .A(n6512), .ZN(n6463) );
  INV_X1 U3943 ( .A(n5249), .ZN(n6518) );
  INV_X1 U3944 ( .A(n6525), .ZN(n6469) );
  INV_X1 U3945 ( .A(n5275), .ZN(n6539) );
  AND2_X1 U3946 ( .A1(n4077), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6583) );
  INV_X1 U3947 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n6596) );
  INV_X1 U3948 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n6600) );
  INV_X1 U3949 ( .A(n6583), .ZN(n6598) );
  NAND2_X1 U3950 ( .A1(n5855), .A2(n4396), .ZN(n4409) );
  INV_X1 U3951 ( .A(n5718), .ZN(n5719) );
  OAI21_X1 U3952 ( .B1(n5746), .B2(n6395), .A(n5717), .ZN(n5718) );
  INV_X1 U3953 ( .A(n4294), .ZN(n6002) );
  INV_X2 U3954 ( .A(n4106), .ZN(n4102) );
  INV_X1 U3955 ( .A(n3436), .ZN(n3447) );
  NAND2_X1 U3956 ( .A1(n5342), .A2(n5343), .ZN(n5341) );
  AND2_X2 U3957 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4538) );
  OR2_X1 U3958 ( .A1(n4451), .A2(n4609), .ZN(n6561) );
  OR2_X1 U3959 ( .A1(n5704), .A2(n6398), .ZN(n3175) );
  OR4_X1 U3960 ( .A1(n5763), .A2(REIP_REG_31__SCAN_IN), .A3(n6975), .A4(n5762), 
        .ZN(n3176) );
  OR2_X1 U3961 ( .A1(n5774), .A2(n5773), .ZN(n3177) );
  NAND2_X1 U3962 ( .A1(n4294), .A2(n4306), .ZN(n3178) );
  AND2_X1 U3963 ( .A1(n4294), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n3180)
         );
  INV_X1 U3964 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n6241) );
  INV_X1 U3965 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n5382) );
  INV_X1 U3966 ( .A(n4578), .ZN(n4565) );
  AND2_X1 U3967 ( .A1(INSTADDRPOINTER_REG_30__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n3181) );
  NAND2_X1 U3968 ( .A1(n4100), .A2(n4099), .ZN(n3182) );
  AND2_X1 U3969 ( .A1(n4395), .A2(n6583), .ZN(n6292) );
  INV_X1 U3970 ( .A(n6292), .ZN(n4405) );
  INV_X1 U3971 ( .A(n5836), .ZN(n4396) );
  AND2_X1 U3972 ( .A1(n5922), .A2(n4311), .ZN(n3183) );
  OR2_X1 U3973 ( .A1(n5630), .A2(n5613), .ZN(n3184) );
  NAND2_X1 U3974 ( .A1(n3308), .A2(n4676), .ZN(n3342) );
  NAND2_X1 U3975 ( .A1(n4094), .A2(n4664), .ZN(n4106) );
  AND2_X1 U3976 ( .A1(n3919), .A2(n3918), .ZN(n3185) );
  AND2_X1 U3977 ( .A1(n4226), .A2(n4234), .ZN(n3186) );
  AND2_X1 U3978 ( .A1(n3342), .A2(n3321), .ZN(n3309) );
  OR2_X1 U3979 ( .A1(n3434), .A2(n3485), .ZN(n3431) );
  INV_X1 U3980 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4024) );
  AND2_X1 U3981 ( .A1(n4392), .A2(n3324), .ZN(n3246) );
  INV_X1 U3982 ( .A(n3569), .ZN(n3571) );
  AND3_X1 U3983 ( .A1(n3345), .A2(n4425), .A3(n3304), .ZN(n3313) );
  OR2_X1 U3984 ( .A1(n4040), .A2(n4039), .ZN(n4042) );
  AND2_X2 U3985 ( .A1(n4024), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3196)
         );
  OR2_X1 U3986 ( .A1(n3430), .A2(n3429), .ZN(n4227) );
  INV_X1 U3987 ( .A(n3441), .ZN(n3442) );
  AOI22_X1 U3988 ( .A1(n3264), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3293), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3208) );
  INV_X1 U3989 ( .A(n4676), .ZN(n4092) );
  INV_X1 U3990 ( .A(n6142), .ZN(n3744) );
  AND2_X1 U3991 ( .A1(n5563), .A2(n3178), .ZN(n4305) );
  NAND2_X1 U3992 ( .A1(n4294), .A2(n5486), .ZN(n4295) );
  INV_X1 U3993 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n4237) );
  OR2_X1 U3994 ( .A1(n3411), .A2(n3410), .ZN(n4228) );
  NOR2_X1 U3995 ( .A1(n3358), .A2(n3357), .ZN(n3359) );
  OR2_X1 U3996 ( .A1(n3497), .A2(n3496), .ZN(n4250) );
  AND4_X1 U3997 ( .A1(n3230), .A2(n3229), .A3(n3228), .A4(n3227), .ZN(n3231)
         );
  AND2_X1 U3998 ( .A1(n4061), .A2(n4060), .ZN(n4080) );
  INV_X1 U3999 ( .A(n5849), .ZN(n3830) );
  AND2_X1 U4000 ( .A1(n4102), .A2(n5776), .ZN(n4105) );
  AND2_X1 U4001 ( .A1(n5759), .A2(n3153), .ZN(n4015) );
  INV_X1 U4002 ( .A(n3809), .ZN(n3810) );
  NOR2_X1 U4003 ( .A1(n3652), .A2(n5382), .ZN(n3627) );
  NOR2_X1 U4004 ( .A1(n6162), .A2(n6163), .ZN(n4145) );
  NAND2_X1 U4005 ( .A1(n3305), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3485) );
  AND4_X1 U4007 ( .A1(n3254), .A2(n3253), .A3(n3252), .A4(n3251), .ZN(n3255)
         );
  NOR2_X1 U4008 ( .A1(n6646), .A2(n6219), .ZN(n6210) );
  NAND2_X1 U4009 ( .A1(n4105), .A2(n4990), .ZN(n4097) );
  NAND2_X1 U4010 ( .A1(n4664), .A2(n4676), .ZN(n4098) );
  NAND2_X1 U4011 ( .A1(n3963), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4087)
         );
  NOR2_X1 U4012 ( .A1(n4429), .A2(n6596), .ZN(n4009) );
  NOR2_X2 U4013 ( .A1(n5843), .A2(n4175), .ZN(n5831) );
  AND2_X1 U4014 ( .A1(n6161), .A2(n4385), .ZN(n5975) );
  AND2_X1 U4015 ( .A1(n3327), .A2(n3352), .ZN(n4924) );
  OAI21_X1 U4016 ( .B1(n3455), .B2(n3454), .A(n3456), .ZN(n3460) );
  AND2_X1 U4017 ( .A1(n6662), .A2(n4658), .ZN(n4686) );
  AND2_X1 U4018 ( .A1(n3321), .A2(n4986), .ZN(n3343) );
  NAND2_X1 U4019 ( .A1(n4209), .A2(REIP_REG_31__SCAN_IN), .ZN(n4210) );
  NAND2_X1 U4020 ( .A1(n3858), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n3896)
         );
  NOR2_X1 U4021 ( .A1(n3707), .A2(n5374), .ZN(n3740) );
  INV_X1 U4022 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n5302) );
  INV_X1 U4023 ( .A(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n5290) );
  NAND2_X1 U4024 ( .A1(n6675), .A2(n4204), .ZN(n6231) );
  AND2_X1 U4025 ( .A1(n4981), .A2(n4102), .ZN(n4103) );
  AND2_X1 U4027 ( .A1(n3794), .A2(n3793), .ZN(n5593) );
  AOI21_X1 U4028 ( .B1(n5716), .B2(INSTADDRPOINTER_REG_31__SCAN_IN), .A(n5715), 
        .ZN(n5717) );
  OR2_X1 U4029 ( .A1(n6149), .A2(n5959), .ZN(n5953) );
  OAI21_X1 U4030 ( .B1(n4315), .B2(n6004), .A(n4294), .ZN(n4317) );
  NAND2_X1 U4031 ( .A1(n5407), .A2(n5359), .ZN(n5182) );
  OR2_X1 U4032 ( .A1(n4375), .A2(n4374), .ZN(n6395) );
  INV_X1 U4033 ( .A(n4246), .ZN(n4853) );
  INV_X1 U4034 ( .A(n5127), .ZN(n5174) );
  INV_X1 U4035 ( .A(n6479), .ZN(n5456) );
  INV_X1 U4036 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n4854) );
  INV_X1 U4037 ( .A(n6548), .ZN(n5277) );
  AND2_X1 U4038 ( .A1(n4853), .A2(n6025), .ZN(n5238) );
  NAND2_X1 U4039 ( .A1(n3460), .A2(n3459), .ZN(n4547) );
  AND2_X1 U4040 ( .A1(n6600), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4077) );
  OR2_X1 U4041 ( .A1(n5753), .A2(n6598), .ZN(n4410) );
  NAND2_X1 U4042 ( .A1(n4419), .A2(n4410), .ZN(n6675) );
  NAND2_X1 U4043 ( .A1(n3176), .A2(n4210), .ZN(n4211) );
  NAND2_X1 U4044 ( .A1(n3741), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n3762)
         );
  AND2_X1 U4045 ( .A1(n5372), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6229) );
  INV_X1 U4046 ( .A(n6082), .ZN(n6258) );
  AND2_X1 U4047 ( .A1(n5372), .A2(n4983), .ZN(n6247) );
  AND2_X1 U4048 ( .A1(n6675), .A2(n4989), .ZN(n6276) );
  CLKBUF_X1 U4049 ( .A(n5312), .Z(n5331) );
  AND2_X1 U4050 ( .A1(n5860), .A2(n5491), .ZN(n6296) );
  NOR2_X1 U4051 ( .A1(n6333), .A2(n4465), .ZN(n6332) );
  INV_X1 U4052 ( .A(n4610), .ZN(n4579) );
  NOR2_X1 U4053 ( .A1(n3897), .A2(n5800), .ZN(n3939) );
  NAND2_X1 U4054 ( .A1(n3763), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n3809)
         );
  NAND2_X1 U4055 ( .A1(n3577), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3594)
         );
  NAND2_X1 U4056 ( .A1(n3503), .A2(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3526)
         );
  OR2_X1 U4057 ( .A1(n5577), .A2(n5575), .ZN(n5199) );
  INV_X1 U4058 ( .A(n5687), .ZN(n6414) );
  NAND2_X1 U4059 ( .A1(n4338), .A2(n6583), .ZN(n4375) );
  INV_X1 U4060 ( .A(n5414), .ZN(n6281) );
  INV_X1 U4061 ( .A(n4817), .ZN(n4848) );
  NOR2_X1 U4062 ( .A1(n4853), .A2(n4707), .ZN(n4713) );
  AND2_X1 U4063 ( .A1(n4713), .A2(n5138), .ZN(n4793) );
  INV_X1 U4064 ( .A(n5237), .ZN(n5138) );
  INV_X1 U4065 ( .A(n5420), .ZN(n5458) );
  INV_X1 U4066 ( .A(n6450), .ZN(n6478) );
  OR2_X1 U4067 ( .A1(n5005), .A2(n5004), .ZN(n5033) );
  AND2_X1 U4068 ( .A1(n4860), .A2(n5237), .ZN(n4997) );
  INV_X1 U4069 ( .A(n5248), .ZN(n5279) );
  AND2_X1 U4070 ( .A1(n5238), .A2(n5419), .ZN(n6548) );
  INV_X1 U4071 ( .A(n6527), .ZN(n6549) );
  INV_X1 U4072 ( .A(n5080), .ZN(n5063) );
  INV_X1 U4073 ( .A(n6493), .ZN(n6451) );
  INV_X1 U4074 ( .A(n5253), .ZN(n6533) );
  INV_X1 U4075 ( .A(n5267), .ZN(n6546) );
  NOR2_X1 U4076 ( .A1(n4212), .A2(n4211), .ZN(n4213) );
  INV_X1 U4077 ( .A(n6229), .ZN(n6273) );
  INV_X1 U4078 ( .A(n6371), .ZN(n6393) );
  NAND2_X1 U4079 ( .A1(n5372), .A2(n4091), .ZN(n6082) );
  INV_X1 U4080 ( .A(n6277), .ZN(n6218) );
  OR2_X1 U4081 ( .A1(n5824), .A2(n5823), .ZN(n6039) );
  INV_X1 U4082 ( .A(n4396), .ZN(n5854) );
  NAND2_X1 U4083 ( .A1(n5769), .A2(n5653), .ZN(n5680) );
  INV_X1 U4084 ( .A(n6297), .ZN(n6114) );
  OR3_X1 U4085 ( .A1(n5756), .A2(n4464), .A3(n4463), .ZN(n6335) );
  OR2_X1 U4086 ( .A1(n4419), .A2(n4418), .ZN(n4610) );
  NAND2_X1 U4087 ( .A1(n6195), .A2(n4494), .ZN(n6148) );
  OR2_X1 U4088 ( .A1(n6574), .A2(n6598), .ZN(n6195) );
  AND2_X1 U4089 ( .A1(n5630), .A2(n5629), .ZN(n6156) );
  AOI21_X1 U4090 ( .B1(n6420), .B2(n4382), .A(n5576), .ZN(n6186) );
  OR2_X1 U4091 ( .A1(n4375), .A2(n4347), .ZN(n6398) );
  INV_X1 U4092 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n5741) );
  AND2_X1 U4093 ( .A1(n4823), .A2(n4822), .ZN(n4852) );
  INV_X1 U4094 ( .A(n4768), .ZN(n4798) );
  OR2_X1 U4095 ( .A1(n4881), .A2(n5138), .ZN(n6443) );
  INV_X1 U4096 ( .A(n5097), .ZN(n5133) );
  INV_X1 U4097 ( .A(n5136), .ZN(n5177) );
  INV_X1 U4098 ( .A(n4997), .ZN(n5039) );
  NOR2_X1 U4099 ( .A1(n4929), .A2(n4928), .ZN(n4966) );
  NAND2_X1 U4100 ( .A1(n4736), .A2(n5237), .ZN(n4959) );
  NAND2_X1 U4101 ( .A1(n4409), .A2(n4408), .ZN(U2829) );
  NOR2_X2 U4102 ( .A1(n3187), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3198)
         );
  NOR2_X4 U4103 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4431) );
  AND2_X2 U4104 ( .A1(n3195), .A2(n4431), .ZN(n3364) );
  AOI22_X1 U4105 ( .A1(n3172), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3364), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3194) );
  NOR2_X2 U4106 ( .A1(n3188), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n5720)
         );
  AND2_X2 U4107 ( .A1(n5720), .A2(n3196), .ZN(n3362) );
  AOI22_X1 U4108 ( .A1(n3362), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3363), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3193) );
  INV_X1 U4109 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3189) );
  AND2_X2 U4110 ( .A1(n3197), .A2(n5720), .ZN(n3603) );
  AND2_X2 U4111 ( .A1(n3197), .A2(n3195), .ZN(n3404) );
  AOI22_X1 U4112 ( .A1(n3603), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3404), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3192) );
  AND2_X2 U4113 ( .A1(n4518), .A2(n3190), .ZN(n3990) );
  AOI22_X1 U4114 ( .A1(n3972), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n3990), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3191) );
  NAND4_X1 U4115 ( .A1(n3194), .A2(n3193), .A3(n3192), .A4(n3191), .ZN(n3204)
         );
  AOI22_X1 U4116 ( .A1(n3487), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3157), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3202) );
  AND2_X2 U4117 ( .A1(n5720), .A2(n4430), .ZN(n3292) );
  AOI22_X1 U4118 ( .A1(n3264), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3292), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3201) );
  AND2_X2 U4119 ( .A1(n3198), .A2(n4430), .ZN(n3420) );
  AOI22_X1 U4120 ( .A1(n3420), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3173), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3200) );
  AND2_X2 U4121 ( .A1(n5720), .A2(n4431), .ZN(n3405) );
  AOI22_X1 U4122 ( .A1(n3405), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3158), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3199) );
  NAND4_X1 U4123 ( .A1(n3202), .A2(n3201), .A3(n3200), .A4(n3199), .ZN(n3203)
         );
  AOI22_X1 U4124 ( .A1(n3362), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3972), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3207) );
  AOI22_X1 U4125 ( .A1(n3603), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3363), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3206) );
  AOI22_X1 U4126 ( .A1(n3420), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3370), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3205) );
  AOI22_X1 U4127 ( .A1(n3292), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3405), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3212) );
  AOI22_X1 U4128 ( .A1(n3487), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3392), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3211) );
  AOI22_X1 U4129 ( .A1(n3404), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3364), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3210) );
  AOI22_X1 U4130 ( .A1(n3259), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3990), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3209) );
  NAND2_X1 U4131 ( .A1(n3404), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3218) );
  NAND2_X1 U4132 ( .A1(n3487), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3217) );
  NAND2_X1 U4133 ( .A1(n3264), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3216)
         );
  NAND2_X1 U4134 ( .A1(n3292), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3215)
         );
  NAND2_X1 U4135 ( .A1(n3362), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3222) );
  NAND2_X1 U4136 ( .A1(n3363), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3221)
         );
  NAND2_X1 U4137 ( .A1(n3259), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3220) );
  NAND2_X1 U4138 ( .A1(n3972), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3219) );
  NAND2_X1 U4139 ( .A1(n3405), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3226) );
  NAND2_X1 U4140 ( .A1(n3392), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3225) );
  NAND2_X1 U4141 ( .A1(n3370), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3224)
         );
  NAND2_X1 U4142 ( .A1(n3293), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3223)
         );
  NAND2_X1 U4143 ( .A1(n3603), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3230)
         );
  NAND2_X1 U4144 ( .A1(n3420), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3229) );
  NAND2_X1 U4145 ( .A1(n3364), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3228) );
  NAND2_X1 U4146 ( .A1(n3990), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3227) );
  INV_X1 U4147 ( .A(n3235), .ZN(n3291) );
  BUF_X1 U4148 ( .A(n3292), .Z(n3391) );
  AOI22_X1 U4149 ( .A1(n3391), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3363), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3239) );
  AOI22_X1 U4150 ( .A1(n3404), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3364), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3238) );
  AOI22_X1 U4151 ( .A1(n3172), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3990), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3237) );
  AOI22_X1 U4152 ( .A1(n3157), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3370), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3236) );
  NAND4_X1 U4153 ( .A1(n3239), .A2(n3238), .A3(n3237), .A4(n3236), .ZN(n3245)
         );
  AOI22_X1 U4154 ( .A1(n3264), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3362), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3243) );
  AOI22_X1 U4155 ( .A1(n3405), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3420), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3242) );
  AOI22_X1 U4156 ( .A1(n3603), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3972), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3241) );
  AOI22_X1 U4157 ( .A1(n3487), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3293), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3240) );
  NAND4_X1 U4158 ( .A1(n3243), .A2(n3242), .A3(n3241), .A4(n3240), .ZN(n3244)
         );
  OAI21_X1 U4159 ( .B1(n3308), .B2(n4672), .A(n3246), .ZN(n4350) );
  INV_X1 U4160 ( .A(n4350), .ZN(n3257) );
  AOI22_X1 U4161 ( .A1(n3363), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3364), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3250) );
  AOI22_X1 U4162 ( .A1(n3264), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3293), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3249) );
  AOI22_X1 U4163 ( .A1(n3362), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3990), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3248) );
  AOI22_X1 U4164 ( .A1(n3259), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3370), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3247) );
  AOI22_X1 U4165 ( .A1(n3162), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3405), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3254) );
  AOI22_X1 U4166 ( .A1(n3487), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3392), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3253) );
  AOI22_X1 U4167 ( .A1(n3404), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3420), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3252) );
  AOI22_X1 U4168 ( .A1(n3603), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3972), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3251) );
  NAND2_X1 U4169 ( .A1(n3257), .A2(n4676), .ZN(n4332) );
  AOI22_X1 U4170 ( .A1(n3362), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3172), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3263) );
  AOI22_X1 U4171 ( .A1(n3487), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3392), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3262) );
  AOI22_X1 U4172 ( .A1(n3404), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n3363), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3261) );
  AOI22_X1 U4173 ( .A1(n3420), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3293), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3260) );
  AOI22_X1 U4174 ( .A1(n3264), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3405), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3268) );
  AOI22_X1 U4175 ( .A1(n3603), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3364), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3267) );
  AOI22_X1 U4176 ( .A1(n3972), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n3990), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3266) );
  AOI22_X1 U4177 ( .A1(n3292), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3370), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3265) );
  NAND2_X4 U4178 ( .A1(n3179), .A2(n3269), .ZN(n4664) );
  NAND2_X1 U4179 ( .A1(n3362), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3274) );
  NAND2_X1 U4180 ( .A1(n3603), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3273)
         );
  NAND2_X1 U4181 ( .A1(n3404), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3272) );
  NAND2_X1 U4182 ( .A1(n3363), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3271)
         );
  NAND2_X1 U4183 ( .A1(n3405), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3278) );
  NAND2_X1 U4184 ( .A1(n3487), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3277) );
  NAND2_X1 U4185 ( .A1(n3392), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3276) );
  NAND2_X1 U4186 ( .A1(n3293), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3275)
         );
  NAND2_X1 U4187 ( .A1(n3264), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3282)
         );
  NAND2_X1 U4188 ( .A1(n3162), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3281)
         );
  NAND2_X1 U4189 ( .A1(n3420), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3280) );
  NAND2_X1 U4190 ( .A1(n3370), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3279)
         );
  NAND2_X1 U4191 ( .A1(n3259), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3286) );
  NAND2_X1 U4192 ( .A1(n3364), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3285) );
  NAND2_X1 U4193 ( .A1(n3972), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3284) );
  NAND2_X1 U4194 ( .A1(n3990), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3283) );
  BUF_X4 U4195 ( .A(n4094), .Z(n4986) );
  NAND2_X1 U4196 ( .A1(n4333), .A2(n3343), .ZN(n3345) );
  NAND2_X1 U4197 ( .A1(STATE_REG_1__SCAN_IN), .A2(STATE_REG_2__SCAN_IN), .ZN(
        n6621) );
  OAI21_X1 U4198 ( .B1(STATE_REG_1__SCAN_IN), .B2(STATE_REG_2__SCAN_IN), .A(
        n6621), .ZN(n4201) );
  NAND2_X1 U4199 ( .A1(n3321), .A2(n4201), .ZN(n3317) );
  AOI22_X1 U4200 ( .A1(n3264), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3292), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3297) );
  AOI22_X1 U4201 ( .A1(n3487), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3392), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3296) );
  AOI22_X1 U4202 ( .A1(n3420), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3370), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3295) );
  AOI22_X1 U4203 ( .A1(n3405), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3293), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3294) );
  AOI22_X1 U4204 ( .A1(n3172), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3364), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3301) );
  AOI22_X1 U4205 ( .A1(n3972), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n3990), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3300) );
  AOI22_X1 U4206 ( .A1(n3362), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3363), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3299) );
  AOI22_X1 U4207 ( .A1(n3603), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3404), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3298) );
  AOI21_X1 U4208 ( .B1(n3317), .B2(n3291), .A(n4668), .ZN(n3304) );
  OR2_X1 U4209 ( .A1(n3318), .A2(n3305), .ZN(n3306) );
  INV_X1 U4210 ( .A(n3324), .ZN(n5731) );
  AOI21_X1 U4211 ( .B1(n4392), .B2(n3306), .A(n5731), .ZN(n3311) );
  OAI21_X1 U4212 ( .B1(n3315), .B2(n3461), .A(n4668), .ZN(n3310) );
  OAI211_X1 U4213 ( .C1(n4668), .C2(n3311), .A(n3310), .B(n3309), .ZN(n3312)
         );
  NAND2_X1 U4214 ( .A1(n3312), .A2(n4348), .ZN(n3338) );
  NAND3_X1 U4215 ( .A1(n3340), .A2(n3313), .A3(n3338), .ZN(n3314) );
  AND2_X2 U4216 ( .A1(n3314), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3350) );
  INV_X1 U4217 ( .A(n3315), .ZN(n3320) );
  INV_X1 U4218 ( .A(n3317), .ZN(n3325) );
  AND3_X1 U4219 ( .A1(n4348), .A2(n3318), .A3(n4668), .ZN(n3319) );
  INV_X1 U4220 ( .A(n4030), .ZN(n3322) );
  NAND2_X1 U4221 ( .A1(n3322), .A2(n3156), .ZN(n4606) );
  NOR2_X2 U4222 ( .A1(n4606), .A2(n5492), .ZN(n4424) );
  NAND2_X1 U4223 ( .A1(n4424), .A2(n5491), .ZN(n4342) );
  OAI211_X1 U4224 ( .C1(n5754), .C2(n3325), .A(n4344), .B(n4342), .ZN(n3326)
         );
  NAND2_X1 U4225 ( .A1(n3326), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3333) );
  NAND2_X1 U4226 ( .A1(n6597), .A2(n6596), .ZN(n4493) );
  INV_X1 U4227 ( .A(n4493), .ZN(n3482) );
  NAND2_X1 U4228 ( .A1(n4854), .A2(n6558), .ZN(n3327) );
  NAND2_X1 U4229 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n3352) );
  INV_X1 U4230 ( .A(n4077), .ZN(n3481) );
  AOI22_X1 U4231 ( .A1(n3482), .A2(n4924), .B1(n3481), .B2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3330) );
  NAND2_X2 U4232 ( .A1(n3329), .A2(n3328), .ZN(n3356) );
  INV_X1 U4233 ( .A(n3330), .ZN(n3331) );
  NOR2_X1 U4234 ( .A1(n3331), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3332)
         );
  NOR2_X1 U4235 ( .A1(n3333), .A2(n3332), .ZN(n3334) );
  INV_X1 U4236 ( .A(n3334), .ZN(n3335) );
  NAND2_X1 U4237 ( .A1(n3350), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3337) );
  MUX2_X1 U4238 ( .A(n4077), .B(n4493), .S(n6558), .Z(n3336) );
  INV_X1 U4239 ( .A(n3338), .ZN(n3339) );
  NAND2_X1 U4240 ( .A1(n3339), .A2(n3161), .ZN(n4356) );
  INV_X1 U4241 ( .A(n3340), .ZN(n3348) );
  NAND2_X1 U4242 ( .A1(n4668), .A2(n4986), .ZN(n4349) );
  NAND3_X1 U4243 ( .A1(n4349), .A2(n6597), .A3(STATE2_REG_0__SCAN_IN), .ZN(
        n3341) );
  AOI21_X1 U4244 ( .B1(n3156), .B2(n3461), .A(n3341), .ZN(n3346) );
  NAND2_X1 U4245 ( .A1(n3342), .A2(n4413), .ZN(n3344) );
  NAND4_X1 U4246 ( .A1(n3346), .A2(n3345), .A3(n4425), .A4(n3344), .ZN(n3347)
         );
  NAND2_X1 U4247 ( .A1(n4356), .A2(n3349), .ZN(n3382) );
  NAND2_X1 U4248 ( .A1(n3360), .A2(n3356), .ZN(n3355) );
  INV_X1 U4249 ( .A(n3352), .ZN(n3351) );
  NAND2_X1 U4250 ( .A1(n3351), .A2(n5243), .ZN(n4874) );
  NAND2_X1 U4251 ( .A1(n3352), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3353) );
  AND2_X1 U4252 ( .A1(n4874), .A2(n3353), .ZN(n4769) );
  OAI22_X1 U4253 ( .A1(n4769), .A2(n4493), .B1(n4077), .B2(n5243), .ZN(n3354)
         );
  NAND2_X1 U4254 ( .A1(n3355), .A2(n3357), .ZN(n3361) );
  INV_X1 U4255 ( .A(n3356), .ZN(n3358) );
  NAND2_X1 U4256 ( .A1(n3361), .A2(n3478), .ZN(n4526) );
  AOI22_X1 U4257 ( .A1(n3885), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3997), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3368) );
  AOI22_X1 U4258 ( .A1(n3921), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3971), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3367) );
  AOI22_X1 U4259 ( .A1(n3399), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3988), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3366) );
  AOI22_X1 U4260 ( .A1(n4000), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3926), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3365) );
  NAND4_X1 U4261 ( .A1(n3368), .A2(n3367), .A3(n3366), .A4(n3365), .ZN(n3376)
         );
  AOI22_X1 U4262 ( .A1(n3264), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n3992), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3374) );
  AOI22_X1 U4264 ( .A1(n3386), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3998), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3373) );
  AOI22_X1 U4265 ( .A1(n3989), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3991), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3372) );
  AOI22_X1 U4266 ( .A1(n3999), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3966), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3371) );
  NAND4_X1 U4267 ( .A1(n3374), .A2(n3373), .A3(n3372), .A4(n3371), .ZN(n3375)
         );
  OAI22_X2 U4268 ( .A1(n4526), .A2(STATE2_REG_0__SCAN_IN), .B1(n4241), .B2(
        n3485), .ZN(n3380) );
  INV_X1 U4269 ( .A(n3486), .ZN(n3378) );
  AOI22_X1 U4270 ( .A1(n3378), .A2(n3377), .B1(n4062), .B2(
        INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3379) );
  INV_X1 U4271 ( .A(n3381), .ZN(n3384) );
  INV_X1 U4272 ( .A(n3382), .ZN(n3383) );
  NAND2_X1 U4273 ( .A1(n3384), .A2(n3383), .ZN(n3385) );
  NAND2_X1 U4274 ( .A1(n3419), .A2(n3385), .ZN(n3462) );
  AOI22_X1 U4275 ( .A1(n3885), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3997), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3390) );
  AOI22_X1 U4276 ( .A1(n3264), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n3405), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3389) );
  AOI22_X1 U4277 ( .A1(n3921), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3988), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3388) );
  AOI22_X1 U4278 ( .A1(n3386), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3966), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3387) );
  NAND4_X1 U4279 ( .A1(n3390), .A2(n3389), .A3(n3388), .A4(n3387), .ZN(n3398)
         );
  AOI22_X1 U4280 ( .A1(n3992), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3369), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3396) );
  AOI22_X1 U4281 ( .A1(n3971), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3972), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3395) );
  AOI22_X1 U4282 ( .A1(n3399), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3990), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3394) );
  AOI22_X1 U4283 ( .A1(n3989), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3991), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3393) );
  NAND4_X1 U4284 ( .A1(n3396), .A2(n3395), .A3(n3394), .A4(n3393), .ZN(n3397)
         );
  NAND2_X1 U4285 ( .A1(n3305), .A2(n4279), .ZN(n4286) );
  INV_X1 U4286 ( .A(n4279), .ZN(n4289) );
  NAND2_X1 U4287 ( .A1(n4289), .A2(n3305), .ZN(n3412) );
  AOI22_X1 U4288 ( .A1(n3885), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3399), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3403) );
  AOI22_X1 U4289 ( .A1(n3386), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n3998), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3402) );
  AOI22_X1 U4290 ( .A1(n3264), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n3989), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3401) );
  AOI22_X1 U4291 ( .A1(n3921), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3988), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3400) );
  NAND4_X1 U4292 ( .A1(n3403), .A2(n3402), .A3(n3401), .A4(n3400), .ZN(n3411)
         );
  AOI22_X1 U4293 ( .A1(n3997), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n4000), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3409) );
  AOI22_X1 U4294 ( .A1(n3405), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3966), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3408) );
  AOI22_X1 U4295 ( .A1(n3971), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n3926), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3407) );
  AOI22_X1 U4296 ( .A1(n3992), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3991), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3406) );
  NAND4_X1 U4297 ( .A1(n3409), .A2(n3408), .A3(n3407), .A4(n3406), .ZN(n3410)
         );
  MUX2_X1 U4298 ( .A(n4286), .B(n3412), .S(n4228), .Z(n3413) );
  INV_X1 U4299 ( .A(n3413), .ZN(n3414) );
  NAND2_X1 U4300 ( .A1(n3414), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3456) );
  NAND2_X1 U4301 ( .A1(n4062), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3416) );
  AOI21_X1 U4302 ( .B1(n4348), .B2(n4228), .A(n6596), .ZN(n3415) );
  NAND3_X1 U4303 ( .A1(n3416), .A2(n3415), .A3(n4286), .ZN(n3457) );
  NOR2_X1 U4304 ( .A1(n4286), .A2(n6596), .ZN(n3417) );
  AOI22_X1 U4305 ( .A1(INSTQUEUE_REG_3__1__SCAN_IN), .A2(n3997), .B1(n3971), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3424) );
  AOI22_X1 U4306 ( .A1(INSTQUEUE_REG_15__1__SCAN_IN), .A2(n3836), .B1(n3992), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3423) );
  AOI22_X1 U4307 ( .A1(INSTQUEUE_REG_10__1__SCAN_IN), .A2(n3921), .B1(n3399), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3422) );
  AOI22_X1 U4308 ( .A1(n3989), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3991), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3421) );
  NAND4_X1 U4309 ( .A1(n3424), .A2(n3423), .A3(n3422), .A4(n3421), .ZN(n3430)
         );
  AOI22_X1 U4310 ( .A1(INSTQUEUE_REG_6__1__SCAN_IN), .A2(n3386), .B1(n3998), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3428) );
  AOI22_X1 U4311 ( .A1(n3885), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3988), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3427) );
  AOI22_X1 U4312 ( .A1(n3999), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3966), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3426) );
  AOI22_X1 U4313 ( .A1(n4000), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n3926), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3425) );
  NAND4_X1 U4314 ( .A1(n3428), .A2(n3427), .A3(n3426), .A4(n3425), .ZN(n3429)
         );
  NAND2_X1 U4315 ( .A1(n4062), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3433) );
  OR2_X1 U4316 ( .A1(n3485), .A2(n4279), .ZN(n3432) );
  OAI211_X1 U4317 ( .C1(n3486), .C2(n3434), .A(n3433), .B(n3432), .ZN(n3445)
         );
  NAND2_X1 U4318 ( .A1(n3436), .A2(n3445), .ZN(n3435) );
  NAND2_X1 U4319 ( .A1(n3446), .A2(n3435), .ZN(n3439) );
  INV_X1 U4320 ( .A(n3445), .ZN(n3437) );
  NAND2_X1 U4321 ( .A1(n3447), .A2(n3437), .ZN(n3438) );
  NAND2_X1 U4322 ( .A1(n3167), .A2(n3444), .ZN(n4215) );
  NAND2_X1 U4323 ( .A1(n3461), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3655) );
  INV_X2 U4324 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n6590) );
  NAND2_X1 U4325 ( .A1(n6590), .A2(STATEBS16_REG_SCAN_IN), .ZN(n3720) );
  NAND2_X1 U4326 ( .A1(n4651), .A2(n3704), .ZN(n3452) );
  AOI22_X1 U4327 ( .A1(n4019), .A2(EAX_REG_1__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n6590), .ZN(n3450) );
  AND2_X1 U4328 ( .A1(n5491), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3464) );
  NAND2_X1 U4329 ( .A1(n3464), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3449) );
  AND2_X1 U4330 ( .A1(n3450), .A2(n3449), .ZN(n3451) );
  NAND2_X1 U4331 ( .A1(n3452), .A2(n3451), .ZN(n4509) );
  INV_X1 U4332 ( .A(n3453), .ZN(n3455) );
  INV_X1 U4333 ( .A(n3457), .ZN(n3454) );
  INV_X1 U4334 ( .A(n3456), .ZN(n3458) );
  NAND2_X1 U4335 ( .A1(n3458), .A2(n3457), .ZN(n3459) );
  AOI21_X1 U4336 ( .B1(n4547), .B2(n3461), .A(n6590), .ZN(n4491) );
  OR2_X1 U4337 ( .A1(n3463), .A2(n3655), .ZN(n3469) );
  INV_X1 U4338 ( .A(n3464), .ZN(n3525) );
  INV_X1 U4339 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n5665) );
  NAND2_X1 U4340 ( .A1(PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n6590), .ZN(n3466)
         );
  NAND2_X1 U4341 ( .A1(n4019), .A2(EAX_REG_0__SCAN_IN), .ZN(n3465) );
  OAI211_X1 U4342 ( .C1(n3525), .C2(n5665), .A(n3466), .B(n3465), .ZN(n3467)
         );
  INV_X1 U4343 ( .A(n3467), .ZN(n3468) );
  NAND2_X1 U4344 ( .A1(n3469), .A2(n3468), .ZN(n4490) );
  INV_X1 U4345 ( .A(n4490), .ZN(n3470) );
  NAND2_X1 U4346 ( .A1(n3470), .A2(n3153), .ZN(n3471) );
  NAND2_X1 U4347 ( .A1(n4489), .A2(n3471), .ZN(n4511) );
  OR2_X2 U4348 ( .A1(n3475), .A2(n3474), .ZN(n4636) );
  OAI21_X1 U4349 ( .B1(PHYADDRPOINTER_REG_2__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_1__SCAN_IN), .A(n3502), .ZN(n6369) );
  AOI22_X1 U4350 ( .A1(n3153), .A2(n6369), .B1(n4018), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3473) );
  NAND2_X1 U4351 ( .A1(n4014), .A2(EAX_REG_2__SCAN_IN), .ZN(n3472) );
  OAI211_X1 U4352 ( .C1(n3525), .C2(n5741), .A(n3473), .B(n3472), .ZN(n4635)
         );
  NAND2_X1 U4353 ( .A1(n3475), .A2(n3474), .ZN(n3476) );
  NAND2_X1 U4354 ( .A1(n3477), .A2(n3476), .ZN(n4634) );
  NAND2_X1 U4355 ( .A1(n3479), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3484) );
  INV_X1 U4356 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6573) );
  NOR3_X1 U4357 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n5243), .A3(n4854), 
        .ZN(n6457) );
  NAND2_X1 U4358 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6457), .ZN(n6446) );
  NAND2_X1 U4359 ( .A1(n6573), .A2(n6446), .ZN(n3480) );
  NAND3_X1 U4360 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .ZN(n5042) );
  INV_X1 U4361 ( .A(n5042), .ZN(n4655) );
  NAND2_X1 U4362 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4655), .ZN(n4654) );
  AOI22_X1 U4363 ( .A1(n3482), .A2(n4925), .B1(n3481), .B2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3483) );
  AOI22_X1 U4364 ( .A1(n3992), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3999), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3491) );
  AOI22_X1 U4365 ( .A1(n3386), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3998), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3490) );
  AOI22_X1 U4366 ( .A1(n3831), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3926), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3489) );
  AOI22_X1 U4367 ( .A1(n3921), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3991), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3488) );
  NAND4_X1 U4368 ( .A1(n3491), .A2(n3490), .A3(n3489), .A4(n3488), .ZN(n3497)
         );
  AOI22_X1 U4369 ( .A1(n3971), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3399), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3495) );
  AOI22_X1 U4370 ( .A1(n3997), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n3989), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3494) );
  AOI22_X1 U4371 ( .A1(n3988), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n4000), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3493) );
  AOI22_X1 U4372 ( .A1(n3836), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n3966), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3492) );
  NAND4_X1 U4373 ( .A1(n3495), .A2(n3494), .A3(n3493), .A4(n3492), .ZN(n3496)
         );
  AOI22_X1 U4374 ( .A1(n4074), .A2(n4250), .B1(INSTQUEUE_REG_0__3__SCAN_IN), 
        .B2(n4062), .ZN(n3498) );
  INV_X1 U4375 ( .A(n4998), .ZN(n3500) );
  NAND2_X1 U4376 ( .A1(n3167), .A2(n4998), .ZN(n3501) );
  NAND2_X2 U4377 ( .A1(n3533), .A2(n3501), .ZN(n4246) );
  NAND2_X1 U4378 ( .A1(n4853), .A2(n3704), .ZN(n3508) );
  OAI21_X1 U4379 ( .B1(PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n3503), .A(n3526), 
        .ZN(n6360) );
  AOI22_X1 U4380 ( .A1(n3153), .A2(n6360), .B1(n4018), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3505) );
  NAND2_X1 U4381 ( .A1(n4014), .A2(EAX_REG_3__SCAN_IN), .ZN(n3504) );
  OAI211_X1 U4382 ( .C1(n3525), .C2(n3165), .A(n3505), .B(n3504), .ZN(n3506)
         );
  INV_X1 U4383 ( .A(n3506), .ZN(n3507) );
  AOI22_X1 U4384 ( .A1(n3831), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3997), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3512) );
  AOI22_X1 U4385 ( .A1(n3921), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3971), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3511) );
  AOI22_X1 U4386 ( .A1(n3399), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3988), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3510) );
  AOI22_X1 U4387 ( .A1(n4000), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n3926), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3509) );
  NAND4_X1 U4388 ( .A1(n3512), .A2(n3511), .A3(n3510), .A4(n3509), .ZN(n3519)
         );
  AOI22_X1 U4389 ( .A1(n3836), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n3992), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3517) );
  AOI22_X1 U4390 ( .A1(n3386), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3998), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3516) );
  INV_X1 U4391 ( .A(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3513) );
  AOI22_X1 U4392 ( .A1(n3989), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3991), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3515) );
  AOI22_X1 U4393 ( .A1(n3999), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3966), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3514) );
  NAND4_X1 U4394 ( .A1(n3517), .A2(n3516), .A3(n3515), .A4(n3514), .ZN(n3518)
         );
  NAND2_X1 U4395 ( .A1(n4074), .A2(n4267), .ZN(n3521) );
  NAND2_X1 U4396 ( .A1(n4062), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3520) );
  NAND2_X1 U4397 ( .A1(n3521), .A2(n3520), .ZN(n3534) );
  NAND2_X1 U4398 ( .A1(n4249), .A2(n3704), .ZN(n3530) );
  INV_X1 U4399 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n3524) );
  INV_X1 U4400 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n7056) );
  OAI21_X1 U4401 ( .B1(PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n7056), .A(n6590), 
        .ZN(n3523) );
  NAND2_X1 U4402 ( .A1(n4014), .A2(EAX_REG_4__SCAN_IN), .ZN(n3522) );
  OAI211_X1 U4403 ( .C1(n3525), .C2(n3524), .A(n3523), .B(n3522), .ZN(n3528)
         );
  AOI21_X1 U4404 ( .B1(n3526), .B2(n5290), .A(n3531), .ZN(n5285) );
  NAND2_X1 U4405 ( .A1(n5285), .A2(n3153), .ZN(n3527) );
  NAND2_X1 U4406 ( .A1(n3528), .A2(n3527), .ZN(n3529) );
  NAND2_X1 U4407 ( .A1(n3530), .A2(n3529), .ZN(n4642) );
  AND3_X2 U4408 ( .A1(n4634), .A2(n4701), .A3(n4642), .ZN(n4641) );
  OR2_X1 U4409 ( .A1(n3531), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3532) );
  NAND2_X1 U4410 ( .A1(n3576), .A2(n3532), .ZN(n6351) );
  INV_X1 U4411 ( .A(n6351), .ZN(n3550) );
  INV_X1 U4412 ( .A(n3533), .ZN(n3535) );
  NAND2_X1 U4413 ( .A1(n3535), .A2(n3534), .ZN(n3551) );
  AOI22_X1 U4414 ( .A1(n3921), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3971), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3539) );
  AOI22_X1 U4415 ( .A1(n3992), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3989), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3538) );
  AOI22_X1 U4416 ( .A1(n3988), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n4000), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3537) );
  AOI22_X1 U4417 ( .A1(n3999), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3966), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3536) );
  NAND4_X1 U4418 ( .A1(n3539), .A2(n3538), .A3(n3537), .A4(n3536), .ZN(n3545)
         );
  AOI22_X1 U4419 ( .A1(n3386), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3998), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3543) );
  AOI22_X1 U4420 ( .A1(n3997), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n3399), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3542) );
  AOI22_X1 U4421 ( .A1(n3831), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3926), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3541) );
  AOI22_X1 U4422 ( .A1(n3836), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n3991), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3540) );
  NAND4_X1 U4423 ( .A1(n3543), .A2(n3542), .A3(n3541), .A4(n3540), .ZN(n3544)
         );
  NAND2_X1 U4424 ( .A1(n4074), .A2(n4266), .ZN(n3547) );
  NAND2_X1 U4425 ( .A1(n4062), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3546) );
  NAND2_X1 U4426 ( .A1(n3547), .A2(n3546), .ZN(n3552) );
  XNOR2_X1 U4427 ( .A(n3551), .B(n3552), .ZN(n4257) );
  NAND2_X1 U4428 ( .A1(n4257), .A2(n3704), .ZN(n3549) );
  AOI22_X1 U4429 ( .A1(n4014), .A2(EAX_REG_5__SCAN_IN), .B1(n4018), .B2(
        PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3548) );
  AND2_X2 U4430 ( .A1(n4641), .A2(n4733), .ZN(n4813) );
  XNOR2_X1 U4431 ( .A(n3576), .B(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n4916) );
  INV_X1 U4432 ( .A(n3551), .ZN(n3553) );
  NAND2_X1 U4433 ( .A1(n3553), .A2(n3552), .ZN(n3569) );
  AOI22_X1 U4434 ( .A1(n3831), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3997), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3557) );
  AOI22_X1 U4435 ( .A1(n3921), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3971), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3556) );
  AOI22_X1 U4436 ( .A1(n3399), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3988), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3555) );
  AOI22_X1 U4437 ( .A1(n4000), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3926), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3554) );
  NAND4_X1 U4438 ( .A1(n3557), .A2(n3556), .A3(n3555), .A4(n3554), .ZN(n3564)
         );
  AOI22_X1 U4439 ( .A1(n3836), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n3992), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3562) );
  AOI22_X1 U4440 ( .A1(n3386), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3369), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3561) );
  INV_X1 U4441 ( .A(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3558) );
  AOI22_X1 U4442 ( .A1(n3989), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3991), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3560) );
  AOI22_X1 U4443 ( .A1(n3999), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3966), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3559) );
  NAND4_X1 U4444 ( .A1(n3562), .A2(n3561), .A3(n3560), .A4(n3559), .ZN(n3563)
         );
  NAND2_X1 U4445 ( .A1(n4074), .A2(n4277), .ZN(n3566) );
  NAND2_X1 U4446 ( .A1(n4062), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3565) );
  NAND2_X1 U4447 ( .A1(n3566), .A2(n3565), .ZN(n3570) );
  XNOR2_X1 U4448 ( .A(n3569), .B(n3570), .ZN(n4265) );
  NAND2_X1 U4449 ( .A1(n4265), .A2(n3704), .ZN(n3568) );
  AOI22_X1 U4450 ( .A1(n4014), .A2(EAX_REG_6__SCAN_IN), .B1(n4018), .B2(
        PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3567) );
  OAI211_X1 U4451 ( .C1(n4916), .C2(n4012), .A(n3568), .B(n3567), .ZN(n4814)
         );
  AND2_X2 U4452 ( .A1(n4813), .A2(n4814), .ZN(n4968) );
  NAND2_X1 U4453 ( .A1(n3571), .A2(n3570), .ZN(n4285) );
  NAND2_X1 U4454 ( .A1(n4074), .A2(n4279), .ZN(n3573) );
  NAND2_X1 U4455 ( .A1(n4062), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3572) );
  NAND2_X1 U4456 ( .A1(n3573), .A2(n3572), .ZN(n3574) );
  OAI21_X1 U4457 ( .B1(n3577), .B2(PHYADDRPOINTER_REG_7__SCAN_IN), .A(n3594), 
        .ZN(n6345) );
  NAND2_X1 U4458 ( .A1(n6345), .A2(n3153), .ZN(n3579) );
  AOI22_X1 U4459 ( .A1(n4014), .A2(EAX_REG_7__SCAN_IN), .B1(n4018), .B2(
        PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3578) );
  NAND2_X1 U4460 ( .A1(n3579), .A2(n3578), .ZN(n3580) );
  XNOR2_X1 U4461 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .B(n3594), .ZN(n5222) );
  AOI22_X1 U4462 ( .A1(n3997), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n3921), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3584) );
  AOI22_X1 U4463 ( .A1(n3836), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n3971), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3583) );
  AOI22_X1 U4464 ( .A1(n3386), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3992), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3582) );
  AOI22_X1 U4465 ( .A1(n3885), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3926), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3581) );
  NAND4_X1 U4466 ( .A1(n3584), .A2(n3583), .A3(n3582), .A4(n3581), .ZN(n3590)
         );
  AOI22_X1 U4467 ( .A1(n3369), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n4000), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3588) );
  AOI22_X1 U4468 ( .A1(n3399), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n3988), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3587) );
  AOI22_X1 U4469 ( .A1(n3999), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3966), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3586) );
  AOI22_X1 U4470 ( .A1(n3989), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3991), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3585) );
  NAND4_X1 U4471 ( .A1(n3588), .A2(n3587), .A3(n3586), .A4(n3585), .ZN(n3589)
         );
  OR2_X1 U4472 ( .A1(n3590), .A2(n3589), .ZN(n3591) );
  AOI22_X1 U4473 ( .A1(n3704), .A2(n3591), .B1(n4018), .B2(
        PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3593) );
  NAND2_X1 U4474 ( .A1(n4014), .A2(EAX_REG_8__SCAN_IN), .ZN(n3592) );
  OAI211_X1 U4475 ( .C1(n5222), .C2(n4012), .A(n3593), .B(n3592), .ZN(n4967)
         );
  XOR2_X1 U4476 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .B(n3661), .Z(n6234) );
  INV_X1 U4477 ( .A(n6234), .ZN(n5509) );
  INV_X1 U4478 ( .A(EAX_REG_12__SCAN_IN), .ZN(n3597) );
  INV_X1 U4479 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3596) );
  OAI22_X1 U4480 ( .A1(n3776), .A2(n3597), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n3596), .ZN(n3598) );
  NAND2_X1 U4481 ( .A1(n3598), .A2(n4012), .ZN(n3611) );
  AOI22_X1 U4482 ( .A1(n3386), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n3998), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3602) );
  AOI22_X1 U4483 ( .A1(n3921), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3988), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3601) );
  AOI22_X1 U4484 ( .A1(n4000), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3926), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3600) );
  AOI22_X1 U4485 ( .A1(n3966), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3991), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3599) );
  NAND4_X1 U4486 ( .A1(n3602), .A2(n3601), .A3(n3600), .A4(n3599), .ZN(n3609)
         );
  AOI22_X1 U4488 ( .A1(n3831), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3399), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3607) );
  AOI22_X1 U4489 ( .A1(n3997), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n3971), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3606) );
  AOI22_X1 U4490 ( .A1(n3836), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n3999), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3605) );
  AOI22_X1 U4491 ( .A1(n3992), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3989), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3604) );
  NAND4_X1 U4492 ( .A1(n3607), .A2(n3606), .A3(n3605), .A4(n3604), .ZN(n3608)
         );
  OAI21_X1 U4493 ( .B1(n3609), .B2(n3608), .A(n3704), .ZN(n3610) );
  NAND2_X1 U4494 ( .A1(n3611), .A2(n3610), .ZN(n3612) );
  AOI21_X1 U4495 ( .B1(n5509), .B2(n3153), .A(n3612), .ZN(n5356) );
  INV_X1 U4496 ( .A(n5356), .ZN(n3641) );
  AOI22_X1 U4497 ( .A1(n3992), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3971), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3616) );
  AOI22_X1 U4498 ( .A1(n3831), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3399), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3615) );
  AOI22_X1 U4499 ( .A1(n3921), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3988), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3614) );
  AOI22_X1 U4500 ( .A1(n3369), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n3966), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3613) );
  NAND4_X1 U4501 ( .A1(n3616), .A2(n3615), .A3(n3614), .A4(n3613), .ZN(n3622)
         );
  AOI22_X1 U4502 ( .A1(n3386), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3999), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3620) );
  AOI22_X1 U4503 ( .A1(n3989), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4000), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3619) );
  AOI22_X1 U4504 ( .A1(n3997), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3926), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3618) );
  AOI22_X1 U4505 ( .A1(n3836), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3991), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3617) );
  NAND4_X1 U4506 ( .A1(n3620), .A2(n3619), .A3(n3618), .A4(n3617), .ZN(n3621)
         );
  NOR2_X1 U4507 ( .A1(n3622), .A2(n3621), .ZN(n3626) );
  XNOR2_X1 U4508 ( .A(n3623), .B(n6241), .ZN(n6245) );
  NAND2_X1 U4509 ( .A1(n6245), .A2(n3153), .ZN(n3625) );
  AOI22_X1 U4510 ( .A1(n4014), .A2(EAX_REG_11__SCAN_IN), .B1(n4018), .B2(
        PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3624) );
  OAI211_X1 U4511 ( .C1(n3626), .C2(n3655), .A(n3625), .B(n3624), .ZN(n5403)
         );
  XOR2_X1 U4512 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .B(n3627), .Z(n5478) );
  AOI22_X1 U4513 ( .A1(n3921), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3971), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3631) );
  AOI22_X1 U4514 ( .A1(n3831), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3992), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3630) );
  AOI22_X1 U4515 ( .A1(n3836), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3998), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3629) );
  AOI22_X1 U4516 ( .A1(n3399), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3926), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3628) );
  NAND4_X1 U4517 ( .A1(n3631), .A2(n3630), .A3(n3629), .A4(n3628), .ZN(n3637)
         );
  AOI22_X1 U4518 ( .A1(n3997), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3989), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3635) );
  AOI22_X1 U4519 ( .A1(n3988), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n4000), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3634) );
  AOI22_X1 U4520 ( .A1(n3386), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3966), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3633) );
  AOI22_X1 U4521 ( .A1(n3999), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3991), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3632) );
  NAND4_X1 U4522 ( .A1(n3635), .A2(n3634), .A3(n3633), .A4(n3632), .ZN(n3636)
         );
  OR2_X1 U4523 ( .A1(n3637), .A2(n3636), .ZN(n3638) );
  AOI22_X1 U4524 ( .A1(n3704), .A2(n3638), .B1(n4018), .B2(
        PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3640) );
  NAND2_X1 U4525 ( .A1(n4014), .A2(EAX_REG_10__SCAN_IN), .ZN(n3639) );
  OAI211_X1 U4526 ( .C1(n5478), .C2(n4012), .A(n3640), .B(n3639), .ZN(n5307)
         );
  AND2_X1 U4527 ( .A1(n5403), .A2(n5307), .ZN(n5354) );
  AND2_X1 U4528 ( .A1(n3641), .A2(n5354), .ZN(n3657) );
  AOI22_X1 U4529 ( .A1(n3885), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3999), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3645) );
  AOI22_X1 U4530 ( .A1(INSTQUEUE_REG_0__1__SCAN_IN), .A2(n3836), .B1(n3998), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3644) );
  AOI22_X1 U4531 ( .A1(n3399), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3926), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3643) );
  AOI22_X1 U4532 ( .A1(n4000), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3991), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3642) );
  NAND4_X1 U4533 ( .A1(n3645), .A2(n3644), .A3(n3643), .A4(n3642), .ZN(n3651)
         );
  AOI22_X1 U4534 ( .A1(INSTQUEUE_REG_7__1__SCAN_IN), .A2(n3386), .B1(n3992), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3649) );
  AOI22_X1 U4535 ( .A1(INSTQUEUE_REG_15__1__SCAN_IN), .A2(n3971), .B1(n3989), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3648) );
  AOI22_X1 U4536 ( .A1(INSTQUEUE_REG_4__1__SCAN_IN), .A2(n3997), .B1(n3988), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3647) );
  AOI22_X1 U4537 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(n3921), .B1(n3966), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3646) );
  NAND4_X1 U4538 ( .A1(n3649), .A2(n3648), .A3(n3647), .A4(n3646), .ZN(n3650)
         );
  NOR2_X1 U4539 ( .A1(n3651), .A2(n3650), .ZN(n3656) );
  XNOR2_X1 U4540 ( .A(n3652), .B(n5382), .ZN(n5389) );
  NAND2_X1 U4541 ( .A1(n5389), .A2(n3153), .ZN(n3654) );
  AOI22_X1 U4542 ( .A1(n4014), .A2(EAX_REG_9__SCAN_IN), .B1(n4018), .B2(
        PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3653) );
  OAI211_X1 U4543 ( .C1(n3656), .C2(n3655), .A(n3654), .B(n3653), .ZN(n5328)
         );
  AND2_X1 U4544 ( .A1(n3657), .A2(n5328), .ZN(n3658) );
  NAND2_X1 U4545 ( .A1(n4967), .A2(n3658), .ZN(n3659) );
  XNOR2_X1 U4546 ( .A(n3688), .B(n5302), .ZN(n5558) );
  NAND2_X1 U4547 ( .A1(n5558), .A2(n3153), .ZN(n3664) );
  NOR2_X1 U4548 ( .A1(n3720), .A2(n5302), .ZN(n3662) );
  AOI21_X1 U4549 ( .B1(n4014), .B2(EAX_REG_13__SCAN_IN), .A(n3662), .ZN(n3663)
         );
  NAND2_X1 U4550 ( .A1(n3664), .A2(n3663), .ZN(n3676) );
  XNOR2_X2 U4551 ( .A(n5358), .B(n3676), .ZN(n5178) );
  AOI22_X1 U4552 ( .A1(n3831), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3997), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3668) );
  AOI22_X1 U4553 ( .A1(n3992), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3369), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3667) );
  AOI22_X1 U4554 ( .A1(n3386), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3989), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3666) );
  AOI22_X1 U4555 ( .A1(n4000), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3966), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3665) );
  NAND4_X1 U4556 ( .A1(n3668), .A2(n3667), .A3(n3666), .A4(n3665), .ZN(n3674)
         );
  AOI22_X1 U4557 ( .A1(n3836), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n3921), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3672) );
  AOI22_X1 U4558 ( .A1(n3999), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3988), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3671) );
  AOI22_X1 U4559 ( .A1(n3399), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3926), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3670) );
  AOI22_X1 U4560 ( .A1(n3971), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n3991), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3669) );
  NAND4_X1 U4561 ( .A1(n3672), .A2(n3671), .A3(n3670), .A4(n3669), .ZN(n3673)
         );
  OR2_X1 U4562 ( .A1(n3674), .A2(n3673), .ZN(n3675) );
  AND2_X1 U4563 ( .A1(n3704), .A2(n3675), .ZN(n5181) );
  NAND2_X1 U4564 ( .A1(n5178), .A2(n5181), .ZN(n5179) );
  INV_X1 U4565 ( .A(n5358), .ZN(n3677) );
  AOI22_X1 U4566 ( .A1(n3997), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3487), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3681) );
  AOI22_X1 U4567 ( .A1(n3831), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3989), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3680) );
  AOI22_X1 U4568 ( .A1(n3971), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n4000), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3679) );
  AOI22_X1 U4569 ( .A1(n3921), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3926), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3678) );
  NAND4_X1 U4570 ( .A1(n3681), .A2(n3680), .A3(n3679), .A4(n3678), .ZN(n3687)
         );
  AOI22_X1 U4571 ( .A1(n3836), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n3992), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3685) );
  AOI22_X1 U4572 ( .A1(n3999), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3998), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3684) );
  AOI22_X1 U4573 ( .A1(n3399), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3966), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3683) );
  AOI22_X1 U4574 ( .A1(n3988), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3991), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3682) );
  NAND4_X1 U4575 ( .A1(n3685), .A2(n3684), .A3(n3683), .A4(n3682), .ZN(n3686)
         );
  OAI21_X1 U4576 ( .B1(n3687), .B2(n3686), .A(n3704), .ZN(n3691) );
  XNOR2_X1 U4577 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .B(n3692), .ZN(n5567)
         );
  AOI22_X1 U4578 ( .A1(n3153), .A2(n5567), .B1(n4018), .B2(
        PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n3690) );
  NAND2_X1 U4579 ( .A1(n4014), .A2(EAX_REG_14__SCAN_IN), .ZN(n3689) );
  AOI21_X2 U4580 ( .B1(n5179), .B2(n5338), .A(n5339), .ZN(n5336) );
  XNOR2_X1 U4581 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .B(n3707), .ZN(n5547)
         );
  AOI22_X1 U4582 ( .A1(n3997), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3386), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3696) );
  AOI22_X1 U4583 ( .A1(n3921), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3999), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3695) );
  AOI22_X1 U4584 ( .A1(n3971), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n3988), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3694) );
  AOI22_X1 U4585 ( .A1(n4000), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3926), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3693) );
  NAND4_X1 U4586 ( .A1(n3696), .A2(n3695), .A3(n3694), .A4(n3693), .ZN(n3702)
         );
  AOI22_X1 U4587 ( .A1(n3836), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n3369), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3700) );
  AOI22_X1 U4588 ( .A1(n3399), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3989), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3699) );
  AOI22_X1 U4589 ( .A1(n3831), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3966), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3698) );
  AOI22_X1 U4590 ( .A1(n3992), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3991), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3697) );
  NAND4_X1 U4591 ( .A1(n3700), .A2(n3699), .A3(n3698), .A4(n3697), .ZN(n3701)
         );
  OR2_X1 U4592 ( .A1(n3702), .A2(n3701), .ZN(n3703) );
  AOI22_X1 U4593 ( .A1(n3704), .A2(n3703), .B1(n4018), .B2(
        PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3706) );
  NAND2_X1 U4594 ( .A1(n4014), .A2(EAX_REG_15__SCAN_IN), .ZN(n3705) );
  OAI211_X1 U4595 ( .C1(n5547), .C2(n4012), .A(n3706), .B(n3705), .ZN(n5363)
         );
  INV_X1 U4596 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n5374) );
  XNOR2_X1 U4597 ( .A(n3740), .B(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n5925)
         );
  NAND2_X1 U4598 ( .A1(n5925), .A2(n3153), .ZN(n3725) );
  NAND2_X1 U4599 ( .A1(n4672), .A2(n3324), .ZN(n3708) );
  AOI22_X1 U4600 ( .A1(n3831), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n3997), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3712) );
  AOI22_X1 U4601 ( .A1(n3836), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n3992), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3711) );
  AOI22_X1 U4602 ( .A1(n3487), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3369), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3710) );
  AOI22_X1 U4603 ( .A1(n3921), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3988), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3709) );
  NAND4_X1 U4604 ( .A1(n3712), .A2(n3711), .A3(n3710), .A4(n3709), .ZN(n3718)
         );
  AOI22_X1 U4605 ( .A1(n3971), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n4000), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3716) );
  AOI22_X1 U4606 ( .A1(n3999), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3966), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3715) );
  AOI22_X1 U4607 ( .A1(n3399), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3926), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3714) );
  AOI22_X1 U4608 ( .A1(n3989), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3991), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3713) );
  NAND4_X1 U4609 ( .A1(n3716), .A2(n3715), .A3(n3714), .A4(n3713), .ZN(n3717)
         );
  OR2_X1 U4610 ( .A1(n3718), .A2(n3717), .ZN(n3723) );
  INV_X1 U4611 ( .A(EAX_REG_16__SCAN_IN), .ZN(n3721) );
  INV_X1 U4612 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3719) );
  OAI22_X1 U4613 ( .A1(n3776), .A2(n3721), .B1(n3720), .B2(n3719), .ZN(n3722)
         );
  AOI21_X1 U4614 ( .B1(n4009), .B2(n3723), .A(n3722), .ZN(n3724) );
  NAND2_X1 U4615 ( .A1(n3725), .A2(n3724), .ZN(n5463) );
  NAND2_X1 U4616 ( .A1(n5361), .A2(n5463), .ZN(n5461) );
  INV_X1 U4617 ( .A(n5461), .ZN(n3745) );
  AOI22_X1 U4618 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(n3999), .B1(n3998), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3729) );
  AOI22_X1 U4619 ( .A1(n3836), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n3989), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3728) );
  AOI22_X1 U4620 ( .A1(n3831), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4000), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3727) );
  AOI22_X1 U4621 ( .A1(n3921), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3926), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3726) );
  NAND4_X1 U4622 ( .A1(n3729), .A2(n3728), .A3(n3727), .A4(n3726), .ZN(n3735)
         );
  AOI22_X1 U4623 ( .A1(n3997), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3971), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3733) );
  AOI22_X1 U4624 ( .A1(n3399), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3988), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3732) );
  AOI22_X1 U4625 ( .A1(INSTQUEUE_REG_8__1__SCAN_IN), .A2(n3487), .B1(n3966), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3731) );
  AOI22_X1 U4626 ( .A1(n3992), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3991), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3730) );
  NAND4_X1 U4627 ( .A1(n3733), .A2(n3732), .A3(n3731), .A4(n3730), .ZN(n3734)
         );
  NOR2_X1 U4628 ( .A1(n3735), .A2(n3734), .ZN(n3739) );
  NAND2_X1 U4629 ( .A1(n6590), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n3736)
         );
  NAND2_X1 U4630 ( .A1(n4012), .A2(n3736), .ZN(n3737) );
  AOI21_X1 U4631 ( .B1(n4014), .B2(EAX_REG_17__SCAN_IN), .A(n3737), .ZN(n3738)
         );
  OAI21_X1 U4632 ( .B1(n3983), .B2(n3739), .A(n3738), .ZN(n3743) );
  OAI21_X1 U4633 ( .B1(PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n3741), .A(n3762), 
        .ZN(n6227) );
  OR2_X1 U4634 ( .A1(n4012), .A2(n6227), .ZN(n3742) );
  NAND2_X1 U4635 ( .A1(n3743), .A2(n3742), .ZN(n6142) );
  NAND2_X1 U4636 ( .A1(n3745), .A2(n3744), .ZN(n5523) );
  AOI22_X1 U4637 ( .A1(n3836), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n3921), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3749) );
  AOI22_X1 U4638 ( .A1(n3386), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3971), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3748) );
  AOI22_X1 U4639 ( .A1(n3831), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3988), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3747) );
  AOI22_X1 U4640 ( .A1(n4000), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3926), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3746) );
  NAND4_X1 U4641 ( .A1(n3749), .A2(n3748), .A3(n3747), .A4(n3746), .ZN(n3755)
         );
  AOI22_X1 U4642 ( .A1(n3999), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3998), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3753) );
  AOI22_X1 U4643 ( .A1(n3399), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3989), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3752) );
  AOI22_X1 U4644 ( .A1(n3997), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3966), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3751) );
  AOI22_X1 U4645 ( .A1(n3992), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3991), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3750) );
  NAND4_X1 U4646 ( .A1(n3753), .A2(n3752), .A3(n3751), .A4(n3750), .ZN(n3754)
         );
  NOR2_X1 U4647 ( .A1(n3755), .A2(n3754), .ZN(n3759) );
  NAND2_X1 U4648 ( .A1(n6590), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n3756)
         );
  NAND2_X1 U4649 ( .A1(n4012), .A2(n3756), .ZN(n3757) );
  AOI21_X1 U4650 ( .B1(n4014), .B2(EAX_REG_18__SCAN_IN), .A(n3757), .ZN(n3758)
         );
  OAI21_X1 U4651 ( .B1(n3983), .B2(n3759), .A(n3758), .ZN(n3761) );
  XNOR2_X1 U4652 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .B(n3762), .ZN(n6214)
         );
  NAND2_X1 U4653 ( .A1(n3153), .A2(n6214), .ZN(n3760) );
  NAND2_X1 U4654 ( .A1(n3761), .A2(n3760), .ZN(n5527) );
  NOR2_X2 U4655 ( .A1(n5523), .A2(n5527), .ZN(n5525) );
  INV_X1 U4656 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n6212) );
  OR2_X1 U4657 ( .A1(n3763), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n3764)
         );
  NAND2_X1 U4658 ( .A1(n3764), .A2(n3809), .ZN(n6137) );
  INV_X1 U4659 ( .A(n6137), .ZN(n6096) );
  AOI22_X1 U4660 ( .A1(n3831), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3971), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3768) );
  AOI22_X1 U4661 ( .A1(n3836), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3992), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3767) );
  AOI22_X1 U4662 ( .A1(n3386), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3998), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3766) );
  AOI22_X1 U4663 ( .A1(n3997), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3991), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3765) );
  NAND4_X1 U4664 ( .A1(n3768), .A2(n3767), .A3(n3766), .A4(n3765), .ZN(n3774)
         );
  AOI22_X1 U4665 ( .A1(n3921), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3989), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3772) );
  AOI22_X1 U4666 ( .A1(n3399), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3988), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3771) );
  AOI22_X1 U4667 ( .A1(n3999), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3966), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3770) );
  AOI22_X1 U4668 ( .A1(n4000), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3926), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3769) );
  NAND4_X1 U4669 ( .A1(n3772), .A2(n3771), .A3(n3770), .A4(n3769), .ZN(n3773)
         );
  OR2_X1 U4670 ( .A1(n3774), .A2(n3773), .ZN(n3778) );
  NAND2_X1 U4671 ( .A1(n6590), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n3775)
         );
  OAI211_X1 U4672 ( .C1(n3776), .C2(n4622), .A(n4012), .B(n3775), .ZN(n3777)
         );
  AOI21_X1 U4673 ( .B1(n4009), .B2(n3778), .A(n3777), .ZN(n3779) );
  AOI21_X1 U4674 ( .B1(n6096), .B2(n3153), .A(n3779), .ZN(n5528) );
  AND2_X2 U4675 ( .A1(n5525), .A2(n5528), .ZN(n5529) );
  AOI22_X1 U4676 ( .A1(n3831), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3997), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3783) );
  AOI22_X1 U4677 ( .A1(n3921), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3971), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3782) );
  AOI22_X1 U4678 ( .A1(n3399), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n3988), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3781) );
  AOI22_X1 U4679 ( .A1(n4000), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3926), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3780) );
  NAND4_X1 U4680 ( .A1(n3783), .A2(n3782), .A3(n3781), .A4(n3780), .ZN(n3789)
         );
  AOI22_X1 U4681 ( .A1(n3836), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n3992), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3787) );
  AOI22_X1 U4682 ( .A1(n3487), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3369), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3786) );
  AOI22_X1 U4683 ( .A1(n3989), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3991), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3785) );
  AOI22_X1 U4684 ( .A1(n3999), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3966), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3784) );
  NAND4_X1 U4685 ( .A1(n3787), .A2(n3786), .A3(n3785), .A4(n3784), .ZN(n3788)
         );
  NOR2_X1 U4686 ( .A1(n3789), .A2(n3788), .ZN(n3792) );
  INV_X1 U4687 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n6089) );
  AOI21_X1 U4688 ( .B1(n6089), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3790) );
  AOI21_X1 U4689 ( .B1(n4014), .B2(EAX_REG_20__SCAN_IN), .A(n3790), .ZN(n3791)
         );
  OAI21_X1 U4690 ( .B1(n3983), .B2(n3792), .A(n3791), .ZN(n3794) );
  XNOR2_X1 U4691 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .B(n3809), .ZN(n6079)
         );
  NAND2_X1 U4692 ( .A1(n6079), .A2(n3153), .ZN(n3793) );
  NAND2_X1 U4693 ( .A1(n5529), .A2(n5593), .ZN(n5605) );
  AOI22_X1 U4694 ( .A1(n3836), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3992), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3798) );
  AOI22_X1 U4695 ( .A1(n3971), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n3399), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3797) );
  AOI22_X1 U4696 ( .A1(n3921), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3988), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3796) );
  AOI22_X1 U4697 ( .A1(n3998), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3966), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3795) );
  NAND4_X1 U4698 ( .A1(n3798), .A2(n3797), .A3(n3796), .A4(n3795), .ZN(n3804)
         );
  AOI22_X1 U4699 ( .A1(n3386), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3999), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3802) );
  AOI22_X1 U4700 ( .A1(n3997), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n4000), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3801) );
  AOI22_X1 U4701 ( .A1(n3831), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3926), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3800) );
  AOI22_X1 U4702 ( .A1(n3989), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3991), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3799) );
  NAND4_X1 U4703 ( .A1(n3802), .A2(n3801), .A3(n3800), .A4(n3799), .ZN(n3803)
         );
  NOR2_X1 U4704 ( .A1(n3804), .A2(n3803), .ZN(n3808) );
  NAND2_X1 U4705 ( .A1(n6590), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n3805)
         );
  NAND2_X1 U4706 ( .A1(n4012), .A2(n3805), .ZN(n3806) );
  AOI21_X1 U4707 ( .B1(n4014), .B2(EAX_REG_21__SCAN_IN), .A(n3806), .ZN(n3807)
         );
  OAI21_X1 U4708 ( .B1(n3983), .B2(n3808), .A(n3807), .ZN(n3813) );
  OAI21_X1 U4709 ( .B1(n3811), .B2(PHYADDRPOINTER_REG_21__SCAN_IN), .A(n3857), 
        .ZN(n6072) );
  OR2_X1 U4710 ( .A1(n6072), .A2(n4012), .ZN(n3812) );
  NAND2_X1 U4711 ( .A1(n3813), .A2(n3812), .ZN(n5606) );
  NOR2_X2 U4712 ( .A1(n5605), .A2(n5606), .ZN(n5603) );
  AOI22_X1 U4713 ( .A1(n3885), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3997), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3817) );
  AOI22_X1 U4714 ( .A1(n3921), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3971), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3816) );
  AOI22_X1 U4715 ( .A1(n3399), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3988), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3815) );
  AOI22_X1 U4716 ( .A1(n4000), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3926), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3814) );
  NAND4_X1 U4717 ( .A1(n3817), .A2(n3816), .A3(n3815), .A4(n3814), .ZN(n3823)
         );
  AOI22_X1 U4718 ( .A1(n3264), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3992), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3821) );
  AOI22_X1 U4719 ( .A1(n3487), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3369), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3820) );
  AOI22_X1 U4720 ( .A1(n3989), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3991), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3819) );
  AOI22_X1 U4721 ( .A1(n3999), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3966), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3818) );
  NAND4_X1 U4722 ( .A1(n3821), .A2(n3820), .A3(n3819), .A4(n3818), .ZN(n3822)
         );
  NOR2_X1 U4723 ( .A1(n3823), .A2(n3822), .ZN(n3826) );
  INV_X1 U4724 ( .A(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5898) );
  AOI21_X1 U4725 ( .B1(n5898), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3824) );
  AOI21_X1 U4726 ( .B1(n4014), .B2(EAX_REG_22__SCAN_IN), .A(n3824), .ZN(n3825)
         );
  OAI21_X1 U4727 ( .B1(n3983), .B2(n3826), .A(n3825), .ZN(n3829) );
  XNOR2_X1 U4728 ( .A(n3857), .B(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n6063)
         );
  NAND2_X1 U4729 ( .A1(n6063), .A2(n3153), .ZN(n3828) );
  NAND2_X1 U4730 ( .A1(n3829), .A2(n3828), .ZN(n5849) );
  NAND2_X1 U4731 ( .A1(n5603), .A2(n3830), .ZN(n5696) );
  AOI22_X1 U4732 ( .A1(n3831), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3997), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3835) );
  AOI22_X1 U4733 ( .A1(n3921), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3971), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3834) );
  AOI22_X1 U4734 ( .A1(n3399), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3988), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3833) );
  AOI22_X1 U4735 ( .A1(n4000), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3926), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3832) );
  NAND4_X1 U4736 ( .A1(n3835), .A2(n3834), .A3(n3833), .A4(n3832), .ZN(n3842)
         );
  AOI22_X1 U4737 ( .A1(n3836), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3992), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3840) );
  AOI22_X1 U4738 ( .A1(n3386), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3369), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3839) );
  AOI22_X1 U4739 ( .A1(n3989), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3991), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3838) );
  AOI22_X1 U4740 ( .A1(n3999), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3966), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3837) );
  NAND4_X1 U4741 ( .A1(n3840), .A2(n3839), .A3(n3838), .A4(n3837), .ZN(n3841)
         );
  NOR2_X1 U4742 ( .A1(n3842), .A2(n3841), .ZN(n3862) );
  AOI22_X1 U4743 ( .A1(n3487), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3369), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3846) );
  AOI22_X1 U4744 ( .A1(n3971), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n3988), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3845) );
  AOI22_X1 U4745 ( .A1(n3836), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n3966), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3844) );
  AOI22_X1 U4746 ( .A1(n3831), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n3926), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3843) );
  NAND4_X1 U4747 ( .A1(n3846), .A2(n3845), .A3(n3844), .A4(n3843), .ZN(n3852)
         );
  AOI22_X1 U4748 ( .A1(n3992), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n3999), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3850) );
  AOI22_X1 U4749 ( .A1(n3997), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n3399), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3849) );
  AOI22_X1 U4750 ( .A1(n3921), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4000), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3848) );
  AOI22_X1 U4751 ( .A1(n3989), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3991), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3847) );
  NAND4_X1 U4752 ( .A1(n3850), .A2(n3849), .A3(n3848), .A4(n3847), .ZN(n3851)
         );
  NOR2_X1 U4753 ( .A1(n3852), .A2(n3851), .ZN(n3863) );
  XNOR2_X1 U4754 ( .A(n3862), .B(n3863), .ZN(n3856) );
  NAND2_X1 U4755 ( .A1(n6590), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n3853)
         );
  NAND2_X1 U4756 ( .A1(n4012), .A2(n3853), .ZN(n3854) );
  AOI21_X1 U4757 ( .B1(n4014), .B2(EAX_REG_23__SCAN_IN), .A(n3854), .ZN(n3855)
         );
  OAI21_X1 U4758 ( .B1(n3983), .B2(n3856), .A(n3855), .ZN(n3861) );
  OR2_X1 U4759 ( .A1(n3858), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n3859)
         );
  NAND2_X1 U4760 ( .A1(n3896), .A2(n3859), .ZN(n5810) );
  NAND2_X1 U4761 ( .A1(n3861), .A2(n3860), .ZN(n5698) );
  NOR2_X2 U4762 ( .A1(n5696), .A2(n5698), .ZN(n5694) );
  OR2_X1 U4763 ( .A1(n3863), .A2(n3862), .ZN(n3880) );
  AOI22_X1 U4764 ( .A1(n3885), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3386), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3867) );
  AOI22_X1 U4765 ( .A1(n3999), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3369), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3866) );
  AOI22_X1 U4766 ( .A1(n3992), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n3989), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3865) );
  AOI22_X1 U4767 ( .A1(n3966), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n3991), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3864) );
  NAND4_X1 U4768 ( .A1(n3867), .A2(n3866), .A3(n3865), .A4(n3864), .ZN(n3873)
         );
  AOI22_X1 U4769 ( .A1(n3971), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n3399), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3871) );
  AOI22_X1 U4770 ( .A1(INSTQUEUE_REG_6__1__SCAN_IN), .A2(n3997), .B1(n3988), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3870) );
  AOI22_X1 U4771 ( .A1(n3921), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4000), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3869) );
  AOI22_X1 U4772 ( .A1(n3836), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n3926), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3868) );
  NAND4_X1 U4773 ( .A1(n3871), .A2(n3870), .A3(n3869), .A4(n3868), .ZN(n3872)
         );
  NOR2_X1 U4774 ( .A1(n3873), .A2(n3872), .ZN(n3879) );
  XNOR2_X1 U4775 ( .A(n3880), .B(n3879), .ZN(n3878) );
  XNOR2_X1 U4776 ( .A(n3896), .B(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n6054)
         );
  NAND2_X1 U4777 ( .A1(n4019), .A2(EAX_REG_24__SCAN_IN), .ZN(n3875) );
  NAND2_X1 U4778 ( .A1(n4018), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n3874)
         );
  OAI211_X1 U4779 ( .C1(n6054), .C2(n4012), .A(n3875), .B(n3874), .ZN(n3876)
         );
  INV_X1 U4780 ( .A(n3876), .ZN(n3877) );
  OAI21_X1 U4781 ( .B1(n3878), .B2(n3983), .A(n3877), .ZN(n5840) );
  OR2_X1 U4782 ( .A1(n3880), .A2(n3879), .ZN(n3902) );
  AOI22_X1 U4783 ( .A1(n3992), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n3999), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3884) );
  AOI22_X1 U4784 ( .A1(n3997), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3399), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3883) );
  AOI22_X1 U4785 ( .A1(n3971), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n3988), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3882) );
  AOI22_X1 U4786 ( .A1(n3921), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3926), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3881) );
  NAND4_X1 U4787 ( .A1(n3884), .A2(n3883), .A3(n3882), .A4(n3881), .ZN(n3891)
         );
  AOI22_X1 U4788 ( .A1(n3386), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3998), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3889) );
  AOI22_X1 U4789 ( .A1(n3885), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4000), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3888) );
  AOI22_X1 U4790 ( .A1(n3836), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3966), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3887) );
  AOI22_X1 U4791 ( .A1(n3989), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3991), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3886) );
  NAND4_X1 U4792 ( .A1(n3889), .A2(n3888), .A3(n3887), .A4(n3886), .ZN(n3890)
         );
  NOR2_X1 U4793 ( .A1(n3891), .A2(n3890), .ZN(n3903) );
  XNOR2_X1 U4794 ( .A(n3902), .B(n3903), .ZN(n3894) );
  INV_X1 U4795 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5800) );
  AOI21_X1 U4796 ( .B1(n5800), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3892) );
  AOI21_X1 U4797 ( .B1(n4014), .B2(EAX_REG_25__SCAN_IN), .A(n3892), .ZN(n3893)
         );
  OAI21_X1 U4798 ( .B1(n3894), .B2(n3983), .A(n3893), .ZN(n3901) );
  INV_X1 U4799 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n3895) );
  AND2_X1 U4800 ( .A1(n3897), .A2(n5800), .ZN(n3898) );
  OR2_X1 U4801 ( .A1(n3898), .A2(n3939), .ZN(n6132) );
  INV_X1 U4802 ( .A(n6132), .ZN(n3899) );
  NAND2_X1 U4803 ( .A1(n3899), .A2(n3153), .ZN(n3900) );
  NAND2_X1 U4804 ( .A1(n5788), .A2(n5787), .ZN(n5790) );
  NOR2_X1 U4805 ( .A1(n3903), .A2(n3902), .ZN(n3934) );
  AOI22_X1 U4806 ( .A1(n3831), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3997), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3907) );
  AOI22_X1 U4807 ( .A1(n3921), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3971), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3906) );
  AOI22_X1 U4808 ( .A1(n3399), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3988), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3905) );
  AOI22_X1 U4809 ( .A1(n4000), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3990), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3904) );
  NAND4_X1 U4810 ( .A1(n3907), .A2(n3906), .A3(n3905), .A4(n3904), .ZN(n3913)
         );
  AOI22_X1 U4811 ( .A1(n3836), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3992), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3911) );
  AOI22_X1 U4812 ( .A1(n3386), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3369), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3910) );
  AOI22_X1 U4813 ( .A1(n3989), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3991), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3909) );
  AOI22_X1 U4814 ( .A1(n3999), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3966), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3908) );
  NAND4_X1 U4815 ( .A1(n3911), .A2(n3910), .A3(n3909), .A4(n3908), .ZN(n3912)
         );
  OR2_X1 U4816 ( .A1(n3913), .A2(n3912), .ZN(n3933) );
  XNOR2_X1 U4817 ( .A(n3934), .B(n3933), .ZN(n3917) );
  NAND2_X1 U4818 ( .A1(n6590), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n3914)
         );
  NAND2_X1 U4819 ( .A1(n4012), .A2(n3914), .ZN(n3915) );
  AOI21_X1 U4820 ( .B1(n4014), .B2(EAX_REG_26__SCAN_IN), .A(n3915), .ZN(n3916)
         );
  OAI21_X1 U4821 ( .B1(n3917), .B2(n3983), .A(n3916), .ZN(n3919) );
  INV_X1 U4822 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n5882) );
  XNOR2_X1 U4823 ( .A(n3939), .B(n5882), .ZN(n6044) );
  NAND2_X1 U4824 ( .A1(n6044), .A2(n3153), .ZN(n3918) );
  AOI22_X1 U4825 ( .A1(n3997), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3992), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3925) );
  AOI22_X1 U4826 ( .A1(n3971), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n3399), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3924) );
  AOI22_X1 U4827 ( .A1(n3921), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n4000), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3923) );
  AOI22_X1 U4828 ( .A1(n3369), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3966), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3922) );
  NAND4_X1 U4829 ( .A1(n3925), .A2(n3924), .A3(n3923), .A4(n3922), .ZN(n3932)
         );
  AOI22_X1 U4830 ( .A1(n3487), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3999), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3930) );
  AOI22_X1 U4831 ( .A1(n3989), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3988), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3929) );
  AOI22_X1 U4832 ( .A1(n3831), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3926), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3928) );
  AOI22_X1 U4833 ( .A1(n3836), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n3991), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3927) );
  NAND4_X1 U4834 ( .A1(n3930), .A2(n3929), .A3(n3928), .A4(n3927), .ZN(n3931)
         );
  NOR2_X1 U4835 ( .A1(n3932), .A2(n3931), .ZN(n3956) );
  NAND2_X1 U4836 ( .A1(n3934), .A2(n3933), .ZN(n3955) );
  XNOR2_X1 U4837 ( .A(n3956), .B(n3955), .ZN(n3938) );
  NAND2_X1 U4838 ( .A1(n6590), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n3935)
         );
  NAND2_X1 U4839 ( .A1(n4012), .A2(n3935), .ZN(n3936) );
  AOI21_X1 U4840 ( .B1(n4014), .B2(EAX_REG_27__SCAN_IN), .A(n3936), .ZN(n3937)
         );
  OAI21_X1 U4841 ( .B1(n3938), .B2(n3983), .A(n3937), .ZN(n3944) );
  INV_X1 U4842 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n3940) );
  NAND2_X1 U4843 ( .A1(n3941), .A2(n3940), .ZN(n3942) );
  NAND2_X1 U4844 ( .A1(n3962), .A2(n3942), .ZN(n6036) );
  NAND2_X1 U4845 ( .A1(n3944), .A2(n3943), .ZN(n5822) );
  AOI22_X1 U4846 ( .A1(n3831), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3997), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3948) );
  AOI22_X1 U4847 ( .A1(n3921), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3971), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3947) );
  AOI22_X1 U4848 ( .A1(n3399), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3988), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3946) );
  AOI22_X1 U4849 ( .A1(n4000), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3990), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3945) );
  NAND4_X1 U4850 ( .A1(n3948), .A2(n3947), .A3(n3946), .A4(n3945), .ZN(n3954)
         );
  AOI22_X1 U4851 ( .A1(n3836), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3992), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3952) );
  AOI22_X1 U4852 ( .A1(n3487), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3998), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3951) );
  AOI22_X1 U4853 ( .A1(n3989), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3991), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3950) );
  AOI22_X1 U4854 ( .A1(n3999), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3966), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3949) );
  NAND4_X1 U4855 ( .A1(n3952), .A2(n3951), .A3(n3950), .A4(n3949), .ZN(n3953)
         );
  OR2_X1 U4856 ( .A1(n3954), .A2(n3953), .ZN(n3979) );
  NOR2_X1 U4857 ( .A1(n3956), .A2(n3955), .ZN(n3980) );
  XOR2_X1 U4858 ( .A(n3979), .B(n3980), .Z(n3957) );
  NAND2_X1 U4859 ( .A1(n3957), .A2(n4009), .ZN(n3961) );
  INV_X1 U4860 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5650) );
  NOR2_X1 U4861 ( .A1(n5650), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3958) );
  AOI211_X1 U4862 ( .C1(n4014), .C2(EAX_REG_28__SCAN_IN), .A(n3153), .B(n3958), 
        .ZN(n3960) );
  INV_X1 U4863 ( .A(n3962), .ZN(n3959) );
  XOR2_X1 U4864 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .B(n3959), .Z(n5673) );
  AOI22_X1 U4865 ( .A1(n3961), .A2(n3960), .B1(n3153), .B2(n5673), .ZN(n5652)
         );
  NAND2_X2 U4866 ( .A1(n5651), .A2(n5652), .ZN(n5769) );
  INV_X1 U4867 ( .A(n3963), .ZN(n3964) );
  INV_X1 U4868 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5772) );
  NAND2_X1 U4869 ( .A1(n3964), .A2(n5772), .ZN(n3965) );
  NAND2_X1 U4870 ( .A1(n4087), .A2(n3965), .ZN(n5869) );
  AOI22_X1 U4871 ( .A1(n3836), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3992), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3970) );
  AOI22_X1 U4872 ( .A1(n3386), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3966), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3969) );
  AOI22_X1 U4873 ( .A1(n3997), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3990), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3968) );
  AOI22_X1 U4874 ( .A1(n3831), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3991), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3967) );
  NAND4_X1 U4875 ( .A1(n3970), .A2(n3969), .A3(n3968), .A4(n3967), .ZN(n3978)
         );
  AOI22_X1 U4876 ( .A1(n3921), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3399), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3976) );
  AOI22_X1 U4877 ( .A1(n3999), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3998), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3975) );
  AOI22_X1 U4878 ( .A1(n3971), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3989), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3974) );
  AOI22_X1 U4879 ( .A1(n3988), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n4000), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3973) );
  NAND4_X1 U4880 ( .A1(n3976), .A2(n3975), .A3(n3974), .A4(n3973), .ZN(n3977)
         );
  NOR2_X1 U4881 ( .A1(n3978), .A2(n3977), .ZN(n3987) );
  NAND2_X1 U4882 ( .A1(n3980), .A2(n3979), .ZN(n3986) );
  XNOR2_X1 U4883 ( .A(n3987), .B(n3986), .ZN(n3984) );
  AOI21_X1 U4884 ( .B1(PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n6590), .A(n3153), 
        .ZN(n3982) );
  NAND2_X1 U4885 ( .A1(n4019), .A2(EAX_REG_29__SCAN_IN), .ZN(n3981) );
  OAI211_X1 U4886 ( .C1(n3984), .C2(n3983), .A(n3982), .B(n3981), .ZN(n3985)
         );
  OAI21_X1 U4887 ( .B1(n4012), .B2(n5869), .A(n3985), .ZN(n5771) );
  NOR2_X4 U4888 ( .A1(n5769), .A2(n5771), .ZN(n5770) );
  NOR2_X1 U4889 ( .A1(n3987), .A2(n3986), .ZN(n4008) );
  AOI22_X1 U4890 ( .A1(n3989), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3988), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3996) );
  AOI22_X1 U4891 ( .A1(n3386), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3966), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3995) );
  AOI22_X1 U4892 ( .A1(n3831), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3990), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3994) );
  AOI22_X1 U4893 ( .A1(n3992), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n3991), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3993) );
  NAND4_X1 U4894 ( .A1(n3996), .A2(n3995), .A3(n3994), .A4(n3993), .ZN(n4006)
         );
  AOI22_X1 U4895 ( .A1(n3264), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3997), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4004) );
  AOI22_X1 U4896 ( .A1(n3999), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3369), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4003) );
  AOI22_X1 U4897 ( .A1(n3971), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3399), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n4002) );
  AOI22_X1 U4898 ( .A1(n3921), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4000), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4001) );
  NAND4_X1 U4899 ( .A1(n4004), .A2(n4003), .A3(n4002), .A4(n4001), .ZN(n4005)
         );
  NOR2_X1 U4900 ( .A1(n4006), .A2(n4005), .ZN(n4007) );
  XNOR2_X1 U4901 ( .A(n4008), .B(n4007), .ZN(n4010) );
  NAND2_X1 U4902 ( .A1(n4010), .A2(n4009), .ZN(n4017) );
  NAND2_X1 U4903 ( .A1(n6590), .A2(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n4011)
         );
  NAND2_X1 U4904 ( .A1(n4012), .A2(n4011), .ZN(n4013) );
  AOI21_X1 U4905 ( .B1(n4014), .B2(EAX_REG_30__SCAN_IN), .A(n4013), .ZN(n4016)
         );
  XNOR2_X1 U4906 ( .A(n4087), .B(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5759)
         );
  AOI21_X1 U4907 ( .B1(n4017), .B2(n4016), .A(n4015), .ZN(n4389) );
  NAND2_X1 U4908 ( .A1(n5770), .A2(n4389), .ZN(n4022) );
  AOI22_X1 U4909 ( .A1(n4019), .A2(EAX_REG_31__SCAN_IN), .B1(n4018), .B2(
        PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4020) );
  INV_X1 U4910 ( .A(n4020), .ZN(n4021) );
  XNOR2_X2 U4911 ( .A(n4022), .B(n4021), .ZN(n5732) );
  INV_X1 U4912 ( .A(n5732), .ZN(n4214) );
  NAND2_X1 U4913 ( .A1(n4062), .A2(n4023), .ZN(n4063) );
  NAND2_X1 U4914 ( .A1(n4854), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4041) );
  NAND2_X1 U4915 ( .A1(n4024), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n4025) );
  NAND2_X1 U4916 ( .A1(n4041), .A2(n4025), .ZN(n4040) );
  NAND2_X1 U4917 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n6558), .ZN(n4039) );
  INV_X1 U4918 ( .A(n4039), .ZN(n4028) );
  XNOR2_X1 U4919 ( .A(n4040), .B(n4028), .ZN(n4081) );
  NAND2_X1 U4920 ( .A1(n4074), .A2(n4664), .ZN(n4027) );
  NAND2_X1 U4921 ( .A1(n4027), .A2(n5492), .ZN(n4036) );
  AOI21_X1 U4922 ( .B1(n5665), .B2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n4028), 
        .ZN(n4032) );
  NAND2_X1 U4923 ( .A1(n4074), .A2(n4032), .ZN(n4029) );
  NAND2_X1 U4924 ( .A1(n4029), .A2(n4063), .ZN(n4035) );
  NAND2_X1 U4925 ( .A1(n4417), .A2(n5492), .ZN(n4031) );
  NAND2_X1 U4926 ( .A1(n4030), .A2(n4031), .ZN(n4044) );
  NAND2_X1 U4927 ( .A1(n3305), .A2(n5492), .ZN(n4339) );
  AOI21_X1 U4928 ( .B1(n4339), .B2(n4032), .A(n4348), .ZN(n4033) );
  OR2_X1 U4929 ( .A1(n4044), .A2(n4033), .ZN(n4034) );
  OAI211_X1 U4930 ( .C1(n4036), .C2(n4081), .A(n4035), .B(n4034), .ZN(n4038)
         );
  NAND3_X1 U4931 ( .A1(n4036), .A2(STATE2_REG_0__SCAN_IN), .A3(n4081), .ZN(
        n4037) );
  OAI211_X1 U4932 ( .C1(n4063), .C2(n4081), .A(n4038), .B(n4037), .ZN(n4050)
         );
  NAND2_X1 U4933 ( .A1(n4042), .A2(n4041), .ZN(n4053) );
  NAND2_X1 U4934 ( .A1(n5243), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4054) );
  NAND2_X1 U4935 ( .A1(n5741), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4043) );
  NAND2_X1 U4936 ( .A1(n4054), .A2(n4043), .ZN(n4051) );
  XNOR2_X1 U4937 ( .A(n4053), .B(n4051), .ZN(n4079) );
  INV_X1 U4938 ( .A(n4062), .ZN(n4045) );
  NAND2_X1 U4939 ( .A1(n4074), .A2(n4079), .ZN(n4047) );
  INV_X1 U4940 ( .A(n4044), .ZN(n4046) );
  OAI211_X1 U4941 ( .C1(n4079), .C2(n4045), .A(n4047), .B(n4046), .ZN(n4049)
         );
  NOR2_X1 U4942 ( .A1(n4047), .A2(n4046), .ZN(n4048) );
  AOI21_X1 U4943 ( .B1(n4050), .B2(n4049), .A(n4048), .ZN(n4067) );
  INV_X1 U4944 ( .A(n4051), .ZN(n4052) );
  NAND2_X1 U4945 ( .A1(n4053), .A2(n4052), .ZN(n4055) );
  NAND2_X1 U4946 ( .A1(n4055), .A2(n4054), .ZN(n4059) );
  XNOR2_X1 U4947 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4057) );
  NOR2_X1 U4948 ( .A1(n3165), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4056)
         );
  AOI21_X1 U4949 ( .B1(n4059), .B2(n4057), .A(n4056), .ZN(n4070) );
  NAND3_X1 U4950 ( .A1(n4070), .A2(n3524), .A3(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n4061) );
  INV_X1 U4951 ( .A(n4057), .ZN(n4058) );
  XNOR2_X1 U4952 ( .A(n4059), .B(n4058), .ZN(n4060) );
  NOR2_X1 U4953 ( .A1(n4080), .A2(n4062), .ZN(n4066) );
  INV_X1 U4954 ( .A(n4063), .ZN(n4071) );
  INV_X1 U4955 ( .A(n4080), .ZN(n4064) );
  AOI22_X1 U4956 ( .A1(n4071), .A2(n4064), .B1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n6596), .ZN(n4065) );
  OAI21_X1 U4957 ( .B1(n4067), .B2(n4066), .A(n4065), .ZN(n4073) );
  INV_X1 U4958 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n6426) );
  NAND2_X1 U4959 ( .A1(n6426), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4069) );
  NOR2_X1 U4960 ( .A1(n6426), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4068)
         );
  AOI21_X1 U4961 ( .B1(n4070), .B2(n4069), .A(n4068), .ZN(n4083) );
  NAND2_X1 U4962 ( .A1(n4071), .A2(n4083), .ZN(n4072) );
  NAND2_X1 U4963 ( .A1(n4073), .A2(n4072), .ZN(n4076) );
  NAND2_X1 U4964 ( .A1(n4074), .A2(n4083), .ZN(n4075) );
  AND3_X1 U4965 ( .A1(n4081), .A2(n4080), .A3(n4079), .ZN(n4082) );
  OR2_X1 U4966 ( .A1(n4083), .A2(n4082), .ZN(n5747) );
  INV_X1 U4967 ( .A(n5747), .ZN(n4084) );
  NAND2_X1 U4968 ( .A1(n4078), .A2(n4084), .ZN(n5753) );
  INV_X1 U4969 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n6666) );
  NAND2_X1 U4970 ( .A1(n6600), .A2(n6590), .ZN(n6607) );
  NOR3_X1 U4971 ( .A1(n6596), .A2(n6666), .A3(n6607), .ZN(n6582) );
  NAND2_X1 U4972 ( .A1(n6596), .A2(n6590), .ZN(n6608) );
  INV_X1 U4973 ( .A(n6608), .ZN(n6601) );
  AND2_X1 U4974 ( .A1(n6597), .A2(n6601), .ZN(n6371) );
  NOR3_X1 U4975 ( .A1(STATEBS16_REG_SCAN_IN), .A2(n6608), .A3(n6600), .ZN(
        n6603) );
  OR2_X1 U4976 ( .A1(n6371), .A2(n6603), .ZN(n4085) );
  OR2_X1 U4977 ( .A1(n6582), .A2(n4085), .ZN(n4086) );
  INV_X1 U4978 ( .A(n4087), .ZN(n4088) );
  NAND2_X1 U4979 ( .A1(n4088), .A2(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n4090)
         );
  INV_X1 U4980 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4089) );
  NOR2_X1 U4981 ( .A1(n5727), .A2(n6600), .ZN(n4091) );
  NAND2_X4 U4982 ( .A1(n4093), .A2(n4986), .ZN(n4185) );
  INV_X1 U4983 ( .A(n4483), .ZN(n4196) );
  INV_X1 U4984 ( .A(n4102), .ZN(n4168) );
  OAI22_X1 U4985 ( .A1(n4196), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        EBX_REG_31__SCAN_IN), .B2(n4168), .ZN(n4198) );
  INV_X2 U4986 ( .A(n4098), .ZN(n5776) );
  INV_X1 U4987 ( .A(EBX_REG_1__SCAN_IN), .ZN(n4990) );
  INV_X1 U4988 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4574) );
  NAND2_X1 U4989 ( .A1(n4185), .A2(n4574), .ZN(n4095) );
  OAI211_X1 U4990 ( .C1(n4106), .C2(EBX_REG_1__SCAN_IN), .A(n4095), .B(n5597), 
        .ZN(n4096) );
  NAND2_X1 U4991 ( .A1(n4097), .A2(n4096), .ZN(n4101) );
  INV_X1 U4992 ( .A(n4101), .ZN(n4104) );
  NAND2_X1 U4993 ( .A1(n4185), .A2(EBX_REG_0__SCAN_IN), .ZN(n4100) );
  INV_X1 U4994 ( .A(EBX_REG_0__SCAN_IN), .ZN(n4633) );
  NAND2_X1 U4995 ( .A1(n5597), .A2(n4633), .ZN(n4099) );
  XNOR2_X1 U4996 ( .A(n4101), .B(n3182), .ZN(n4981) );
  INV_X1 U4997 ( .A(EBX_REG_2__SCAN_IN), .ZN(n5349) );
  NAND2_X1 U4998 ( .A1(n4194), .A2(n5349), .ZN(n4109) );
  OR2_X1 U4999 ( .A1(n4185), .A2(n5349), .ZN(n4108) );
  NAND2_X1 U5000 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n4168), .ZN(n4107)
         );
  NAND4_X1 U5001 ( .A1(n4142), .A2(n4109), .A3(n4108), .A4(n4107), .ZN(n4638)
         );
  NAND2_X1 U5002 ( .A1(n4639), .A2(n4638), .ZN(n4703) );
  NAND2_X1 U5003 ( .A1(n5776), .A2(EBX_REG_3__SCAN_IN), .ZN(n4111) );
  INV_X1 U5004 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n6408) );
  NAND2_X1 U5005 ( .A1(n4483), .A2(n6408), .ZN(n4110) );
  OAI211_X1 U5006 ( .C1(EBX_REG_3__SCAN_IN), .C2(n4182), .A(n4111), .B(n4110), 
        .ZN(n4704) );
  NOR2_X2 U5007 ( .A1(n4703), .A2(n4704), .ZN(n4644) );
  INV_X1 U5008 ( .A(EBX_REG_4__SCAN_IN), .ZN(n5283) );
  NAND2_X1 U5009 ( .A1(n4194), .A2(n5283), .ZN(n4114) );
  INV_X1 U5010 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n6403) );
  NAND2_X1 U5011 ( .A1(n4185), .A2(n6403), .ZN(n4112) );
  OAI211_X1 U5012 ( .C1(n4168), .C2(EBX_REG_4__SCAN_IN), .A(n4112), .B(n5597), 
        .ZN(n4113) );
  NAND2_X1 U5013 ( .A1(n4114), .A2(n4113), .ZN(n4645) );
  INV_X1 U5014 ( .A(EBX_REG_5__SCAN_IN), .ZN(n4763) );
  INV_X1 U5015 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n5688) );
  AOI22_X1 U5016 ( .A1(n4166), .A2(n4763), .B1(n4483), .B2(n5688), .ZN(n4115)
         );
  OAI21_X1 U5017 ( .B1(n5597), .B2(n4763), .A(n4115), .ZN(n4761) );
  INV_X1 U5018 ( .A(n4185), .ZN(n4171) );
  AOI21_X1 U5019 ( .B1(n4171), .B2(EBX_REG_6__SCAN_IN), .A(n4134), .ZN(n4117)
         );
  NAND2_X1 U5020 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n4168), .ZN(n4116)
         );
  OAI211_X1 U5021 ( .C1(EBX_REG_6__SCAN_IN), .C2(n4174), .A(n4117), .B(n4116), 
        .ZN(n4804) );
  INV_X1 U5022 ( .A(EBX_REG_7__SCAN_IN), .ZN(n5211) );
  INV_X1 U5023 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n6390) );
  AOI22_X1 U5024 ( .A1(n4166), .A2(n5211), .B1(n4483), .B2(n6390), .ZN(n4118)
         );
  OAI21_X1 U5025 ( .B1(n5597), .B2(n5211), .A(n4118), .ZN(n5209) );
  INV_X1 U5026 ( .A(EBX_REG_8__SCAN_IN), .ZN(n5220) );
  NAND2_X1 U5027 ( .A1(n4194), .A2(n5220), .ZN(n4121) );
  INV_X1 U5028 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n5200) );
  NAND2_X1 U5029 ( .A1(n4185), .A2(n5200), .ZN(n4119) );
  OAI211_X1 U5030 ( .C1(n4168), .C2(EBX_REG_8__SCAN_IN), .A(n4119), .B(n5597), 
        .ZN(n4120) );
  NAND2_X1 U5031 ( .A1(n4121), .A2(n4120), .ZN(n4975) );
  INV_X1 U5032 ( .A(EBX_REG_9__SCAN_IN), .ZN(n5334) );
  INV_X1 U5033 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n5486) );
  AOI22_X1 U5034 ( .A1(n4166), .A2(n5334), .B1(n4483), .B2(n5486), .ZN(n4122)
         );
  OAI21_X1 U5035 ( .B1(n5597), .B2(n5334), .A(n4122), .ZN(n5333) );
  INV_X1 U5036 ( .A(EBX_REG_10__SCAN_IN), .ZN(n4123) );
  NAND2_X1 U5037 ( .A1(n4194), .A2(n4123), .ZN(n4126) );
  OR2_X1 U5038 ( .A1(n4185), .A2(n4123), .ZN(n4125) );
  NAND2_X1 U5039 ( .A1(INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n4168), .ZN(n4124) );
  NAND4_X1 U5040 ( .A1(n4142), .A2(n4126), .A3(n4125), .A4(n4124), .ZN(n5313)
         );
  INV_X1 U5041 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n5573) );
  INV_X1 U5042 ( .A(EBX_REG_11__SCAN_IN), .ZN(n6243) );
  NAND2_X1 U5043 ( .A1(n4102), .A2(n6243), .ZN(n4127) );
  OAI211_X1 U5044 ( .C1(n5776), .C2(n5573), .A(n4185), .B(n4127), .ZN(n4128)
         );
  OAI21_X1 U5045 ( .B1(n4182), .B2(EBX_REG_11__SCAN_IN), .A(n4128), .ZN(n5409)
         );
  AOI21_X1 U5046 ( .B1(n4171), .B2(EBX_REG_12__SCAN_IN), .A(n4134), .ZN(n4130)
         );
  NAND2_X1 U5047 ( .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n4168), .ZN(n4129) );
  OAI211_X1 U5048 ( .C1(EBX_REG_12__SCAN_IN), .C2(n4174), .A(n4130), .B(n4129), 
        .ZN(n5359) );
  INV_X1 U5049 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5574) );
  INV_X1 U5050 ( .A(EBX_REG_13__SCAN_IN), .ZN(n4131) );
  NAND2_X1 U5051 ( .A1(n4102), .A2(n4131), .ZN(n4132) );
  OAI211_X1 U5052 ( .C1(n5776), .C2(n5574), .A(n4185), .B(n4132), .ZN(n4133)
         );
  OAI21_X1 U5053 ( .B1(n4182), .B2(EBX_REG_13__SCAN_IN), .A(n4133), .ZN(n5183)
         );
  AOI21_X1 U5054 ( .B1(n4171), .B2(EBX_REG_14__SCAN_IN), .A(n4134), .ZN(n4136)
         );
  NAND2_X1 U5055 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n4168), .ZN(n4135) );
  OAI211_X1 U5056 ( .C1(EBX_REG_14__SCAN_IN), .C2(n4174), .A(n4136), .B(n4135), 
        .ZN(n5343) );
  NAND2_X1 U5057 ( .A1(n5597), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n4137) );
  OAI211_X1 U5058 ( .C1(n4168), .C2(EBX_REG_15__SCAN_IN), .A(n4185), .B(n4137), 
        .ZN(n4138) );
  OAI21_X1 U5059 ( .B1(n4182), .B2(EBX_REG_15__SCAN_IN), .A(n4138), .ZN(n5365)
         );
  NOR2_X2 U5060 ( .A1(n5341), .A2(n5365), .ZN(n5464) );
  INV_X1 U5061 ( .A(EBX_REG_16__SCAN_IN), .ZN(n5496) );
  NAND2_X1 U5062 ( .A1(n4194), .A2(n5496), .ZN(n4141) );
  OR2_X1 U5063 ( .A1(n4185), .A2(n5496), .ZN(n4140) );
  NAND2_X1 U5064 ( .A1(INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n4168), .ZN(n4139) );
  NAND4_X1 U5065 ( .A1(n4142), .A2(n4141), .A3(n4140), .A4(n4139), .ZN(n5465)
         );
  NAND2_X1 U5066 ( .A1(n5464), .A2(n5465), .ZN(n6162) );
  NAND2_X1 U5067 ( .A1(n5597), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n4143) );
  OAI211_X1 U5068 ( .C1(n4168), .C2(EBX_REG_17__SCAN_IN), .A(n4185), .B(n4143), 
        .ZN(n4144) );
  OAI21_X1 U5069 ( .B1(n4182), .B2(EBX_REG_17__SCAN_IN), .A(n4144), .ZN(n6163)
         );
  INV_X1 U5070 ( .A(n4145), .ZN(n6165) );
  INV_X1 U5071 ( .A(EBX_REG_19__SCAN_IN), .ZN(n6100) );
  NAND2_X1 U5072 ( .A1(n4194), .A2(n6100), .ZN(n4149) );
  INV_X1 U5073 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n6004) );
  NAND2_X1 U5074 ( .A1(n4185), .A2(n6004), .ZN(n4147) );
  NAND2_X1 U5075 ( .A1(n4102), .A2(n6100), .ZN(n4146) );
  NAND3_X1 U5076 ( .A1(n4147), .A2(n5597), .A3(n4146), .ZN(n4148) );
  INV_X1 U5077 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5994) );
  NOR2_X1 U5078 ( .A1(n4168), .A2(EBX_REG_20__SCAN_IN), .ZN(n4150) );
  AOI21_X1 U5079 ( .B1(n4483), .B2(n5994), .A(n4150), .ZN(n5599) );
  OR2_X1 U5080 ( .A1(n4196), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n4152)
         );
  INV_X1 U5081 ( .A(EBX_REG_18__SCAN_IN), .ZN(n4151) );
  NAND2_X1 U5082 ( .A1(n4102), .A2(n4151), .ZN(n5517) );
  NAND2_X1 U5083 ( .A1(n4152), .A2(n5517), .ZN(n5594) );
  NAND2_X1 U5084 ( .A1(n5776), .A2(EBX_REG_20__SCAN_IN), .ZN(n4154) );
  NAND2_X1 U5085 ( .A1(n5594), .A2(n5597), .ZN(n4153) );
  OAI211_X1 U5086 ( .C1(n5599), .C2(n5594), .A(n4154), .B(n4153), .ZN(n4155)
         );
  INV_X1 U5087 ( .A(n4155), .ZN(n4156) );
  OR2_X1 U5088 ( .A1(n4196), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n4158)
         );
  NAND2_X1 U5089 ( .A1(n5776), .A2(EBX_REG_21__SCAN_IN), .ZN(n4157) );
  OAI211_X1 U5090 ( .C1(n4182), .C2(EBX_REG_21__SCAN_IN), .A(n4158), .B(n4157), 
        .ZN(n4159) );
  INV_X1 U5091 ( .A(n4159), .ZN(n5608) );
  NAND2_X1 U5092 ( .A1(n5609), .A2(n5608), .ZN(n4376) );
  INV_X1 U5093 ( .A(EBX_REG_23__SCAN_IN), .ZN(n5811) );
  NAND2_X1 U5094 ( .A1(n4166), .A2(n5811), .ZN(n4162) );
  NAND2_X1 U5095 ( .A1(n5597), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4160) );
  OAI211_X1 U5096 ( .C1(n4168), .C2(EBX_REG_23__SCAN_IN), .A(n4185), .B(n4160), 
        .ZN(n4161) );
  AND2_X1 U5097 ( .A1(n4162), .A2(n4161), .ZN(n4378) );
  NAND2_X1 U5098 ( .A1(n4168), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n4164) );
  NAND2_X1 U5099 ( .A1(n4171), .A2(EBX_REG_22__SCAN_IN), .ZN(n4163) );
  OAI211_X1 U5100 ( .C1(n4174), .C2(EBX_REG_22__SCAN_IN), .A(n4164), .B(n4163), 
        .ZN(n4377) );
  NAND2_X1 U5101 ( .A1(n4378), .A2(n4377), .ZN(n4165) );
  OR2_X2 U5102 ( .A1(n4376), .A2(n4165), .ZN(n5843) );
  INV_X1 U5103 ( .A(EBX_REG_25__SCAN_IN), .ZN(n5801) );
  NAND2_X1 U5104 ( .A1(n4166), .A2(n5801), .ZN(n4170) );
  NAND2_X1 U5105 ( .A1(n4098), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n4167) );
  OAI211_X1 U5106 ( .C1(n4168), .C2(EBX_REG_25__SCAN_IN), .A(n4185), .B(n4167), 
        .ZN(n4169) );
  AND2_X1 U5107 ( .A1(n4170), .A2(n4169), .ZN(n5794) );
  NAND2_X1 U5108 ( .A1(n4168), .A2(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n4173) );
  NAND2_X1 U5109 ( .A1(n4171), .A2(EBX_REG_24__SCAN_IN), .ZN(n4172) );
  OAI211_X1 U5110 ( .C1(n4174), .C2(EBX_REG_24__SCAN_IN), .A(n4173), .B(n4172), 
        .ZN(n5842) );
  NAND2_X1 U5111 ( .A1(n5794), .A2(n5842), .ZN(n4175) );
  INV_X1 U5112 ( .A(EBX_REG_26__SCAN_IN), .ZN(n6053) );
  NAND2_X1 U5113 ( .A1(n4194), .A2(n6053), .ZN(n4179) );
  INV_X1 U5114 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5879) );
  NAND2_X1 U5115 ( .A1(n4185), .A2(n5879), .ZN(n4177) );
  NAND2_X1 U5116 ( .A1(n4102), .A2(n6053), .ZN(n4176) );
  NAND3_X1 U5117 ( .A1(n4177), .A2(n4098), .A3(n4176), .ZN(n4178) );
  NAND2_X1 U5118 ( .A1(n4179), .A2(n4178), .ZN(n5830) );
  AND2_X2 U5119 ( .A1(n5831), .A2(n5830), .ZN(n5833) );
  OR2_X1 U5120 ( .A1(n4196), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n4181)
         );
  NAND2_X1 U5121 ( .A1(n5776), .A2(EBX_REG_27__SCAN_IN), .ZN(n4180) );
  OAI211_X1 U5122 ( .C1(n4182), .C2(EBX_REG_27__SCAN_IN), .A(n4181), .B(n4180), 
        .ZN(n4183) );
  INV_X1 U5123 ( .A(n4183), .ZN(n5825) );
  INV_X1 U5124 ( .A(EBX_REG_28__SCAN_IN), .ZN(n4186) );
  NAND2_X1 U5125 ( .A1(n4194), .A2(n4186), .ZN(n4190) );
  INV_X1 U5126 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n4184) );
  NAND2_X1 U5127 ( .A1(n4185), .A2(n4184), .ZN(n4188) );
  NAND2_X1 U5128 ( .A1(n4102), .A2(n4186), .ZN(n4187) );
  NAND3_X1 U5129 ( .A1(n4188), .A2(n4098), .A3(n4187), .ZN(n4189) );
  AND2_X1 U5130 ( .A1(n4190), .A2(n4189), .ZN(n5668) );
  NOR2_X2 U5131 ( .A1(n5827), .A2(n5668), .ZN(n4191) );
  INV_X1 U5132 ( .A(n4191), .ZN(n5774) );
  OR2_X1 U5133 ( .A1(n4196), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4193)
         );
  INV_X1 U5134 ( .A(EBX_REG_29__SCAN_IN), .ZN(n5818) );
  NAND2_X1 U5135 ( .A1(n4102), .A2(n5818), .ZN(n4192) );
  NAND2_X1 U5136 ( .A1(n4193), .A2(n4192), .ZN(n5775) );
  INV_X1 U5137 ( .A(n4401), .ZN(n4398) );
  NAND2_X1 U5138 ( .A1(n4194), .A2(n5818), .ZN(n5773) );
  AND2_X1 U5139 ( .A1(n4168), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4195)
         );
  AOI21_X1 U5140 ( .B1(n4196), .B2(EBX_REG_30__SCAN_IN), .A(n4195), .ZN(n4400)
         );
  NOR2_X1 U5141 ( .A1(n4401), .A2(n5776), .ZN(n4397) );
  XOR2_X1 U5142 ( .A(n4198), .B(n4197), .Z(n5746) );
  NOR2_X1 U5143 ( .A1(READY_N), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4984) );
  INV_X1 U5144 ( .A(EBX_REG_31__SCAN_IN), .ZN(n5745) );
  OR2_X1 U5145 ( .A1(n4984), .A2(n5745), .ZN(n4199) );
  NOR2_X1 U5146 ( .A1(n4168), .A2(n4199), .ZN(n4200) );
  OR2_X1 U5147 ( .A1(n4201), .A2(STATE_REG_0__SCAN_IN), .ZN(n6615) );
  INV_X1 U5148 ( .A(n6615), .ZN(n4462) );
  NAND2_X1 U5149 ( .A1(n4462), .A2(n4984), .ZN(n6588) );
  NAND2_X1 U5150 ( .A1(n4413), .A2(n6588), .ZN(n4988) );
  NOR2_X1 U5151 ( .A1(n4988), .A2(n5745), .ZN(n4202) );
  AOI22_X1 U5152 ( .A1(PHYADDRPOINTER_REG_31__SCAN_IN), .A2(n6229), .B1(n6675), 
        .B2(n4202), .ZN(n4203) );
  OAI21_X1 U5153 ( .B1(n5746), .B2(n6218), .A(n4203), .ZN(n4212) );
  INV_X1 U5154 ( .A(REIP_REG_20__SCAN_IN), .ZN(n6773) );
  INV_X1 U5155 ( .A(REIP_REG_17__SCAN_IN), .ZN(n6646) );
  NAND2_X1 U5156 ( .A1(n4417), .A2(n6615), .ZN(n4322) );
  AND3_X1 U5157 ( .A1(n4322), .A2(n4984), .A3(n4986), .ZN(n4204) );
  INV_X1 U5158 ( .A(REIP_REG_14__SCAN_IN), .ZN(n6644) );
  INV_X1 U5159 ( .A(REIP_REG_12__SCAN_IN), .ZN(n6640) );
  INV_X1 U5160 ( .A(REIP_REG_5__SCAN_IN), .ZN(n6631) );
  INV_X1 U5161 ( .A(REIP_REG_4__SCAN_IN), .ZN(n6630) );
  NAND3_X1 U5162 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_3__SCAN_IN), .A3(
        REIP_REG_2__SCAN_IN), .ZN(n5289) );
  OR2_X1 U5163 ( .A1(n6630), .A2(n5289), .ZN(n5213) );
  NOR2_X1 U5164 ( .A1(n6631), .A2(n5213), .ZN(n5214) );
  INV_X1 U5165 ( .A(REIP_REG_10__SCAN_IN), .ZN(n6638) );
  INV_X1 U5166 ( .A(REIP_REG_9__SCAN_IN), .ZN(n6637) );
  NAND3_X1 U5167 ( .A1(REIP_REG_8__SCAN_IN), .A2(REIP_REG_7__SCAN_IN), .A3(
        REIP_REG_6__SCAN_IN), .ZN(n5216) );
  NOR3_X1 U5168 ( .A1(n6638), .A2(n6637), .A3(n5216), .ZN(n6240) );
  NAND3_X1 U5169 ( .A1(REIP_REG_11__SCAN_IN), .A2(n5214), .A3(n6240), .ZN(
        n6230) );
  NOR2_X1 U5170 ( .A1(n6640), .A2(n6230), .ZN(n5297) );
  NAND2_X1 U5171 ( .A1(REIP_REG_13__SCAN_IN), .A2(n5297), .ZN(n5397) );
  NOR2_X1 U5172 ( .A1(n6644), .A2(n5397), .ZN(n5369) );
  NAND2_X1 U5173 ( .A1(REIP_REG_15__SCAN_IN), .A2(n5369), .ZN(n4205) );
  NOR2_X1 U5174 ( .A1(n6231), .A2(n4205), .ZN(n5468) );
  NAND2_X1 U5175 ( .A1(REIP_REG_16__SCAN_IN), .A2(n5468), .ZN(n6219) );
  NAND3_X1 U5176 ( .A1(REIP_REG_18__SCAN_IN), .A2(REIP_REG_19__SCAN_IN), .A3(
        n6210), .ZN(n6080) );
  NOR2_X1 U5177 ( .A1(n6773), .A2(n6080), .ZN(n6074) );
  NAND3_X1 U5178 ( .A1(REIP_REG_22__SCAN_IN), .A2(REIP_REG_21__SCAN_IN), .A3(
        n6074), .ZN(n5809) );
  INV_X1 U5179 ( .A(REIP_REG_23__SCAN_IN), .ZN(n7027) );
  NOR2_X1 U5180 ( .A1(n5809), .A2(n7027), .ZN(n5798) );
  AND3_X1 U5181 ( .A1(REIP_REG_24__SCAN_IN), .A2(REIP_REG_26__SCAN_IN), .A3(
        REIP_REG_25__SCAN_IN), .ZN(n4206) );
  NAND2_X1 U5182 ( .A1(n5798), .A2(n4206), .ZN(n6043) );
  INV_X1 U5183 ( .A(REIP_REG_28__SCAN_IN), .ZN(n7057) );
  INV_X1 U5184 ( .A(REIP_REG_27__SCAN_IN), .ZN(n7009) );
  INV_X1 U5185 ( .A(REIP_REG_30__SCAN_IN), .ZN(n6975) );
  INV_X1 U5186 ( .A(REIP_REG_29__SCAN_IN), .ZN(n5762) );
  INV_X1 U5187 ( .A(n5763), .ZN(n5784) );
  INV_X1 U5188 ( .A(REIP_REG_16__SCAN_IN), .ZN(n7038) );
  INV_X1 U5189 ( .A(n5372), .ZN(n5296) );
  NOR3_X1 U5190 ( .A1(n6646), .A2(n7038), .A3(n5467), .ZN(n6090) );
  NAND4_X1 U5191 ( .A1(REIP_REG_20__SCAN_IN), .A2(n6090), .A3(
        REIP_REG_18__SCAN_IN), .A4(REIP_REG_19__SCAN_IN), .ZN(n6061) );
  NAND2_X1 U5192 ( .A1(REIP_REG_22__SCAN_IN), .A2(REIP_REG_21__SCAN_IN), .ZN(
        n6066) );
  NOR3_X1 U5193 ( .A1(n7027), .A2(n6061), .A3(n6066), .ZN(n5797) );
  AOI21_X1 U5194 ( .B1(n5797), .B2(n4206), .A(n6091), .ZN(n6050) );
  AND2_X1 U5195 ( .A1(REIP_REG_28__SCAN_IN), .A2(REIP_REG_27__SCAN_IN), .ZN(
        n4207) );
  NOR2_X1 U5196 ( .A1(n6231), .A2(n4207), .ZN(n4208) );
  OR2_X1 U5197 ( .A1(n6050), .A2(n4208), .ZN(n5678) );
  AOI21_X1 U5198 ( .B1(n5784), .B2(n5762), .A(n5678), .ZN(n5782) );
  OAI21_X1 U5199 ( .B1(REIP_REG_30__SCAN_IN), .B2(n6231), .A(n5782), .ZN(n4209) );
  OAI21_X1 U5200 ( .B1(n4214), .B2(n6082), .A(n4213), .ZN(U2796) );
  INV_X1 U5201 ( .A(n4215), .ZN(n4216) );
  NAND2_X1 U5202 ( .A1(n4216), .A2(n4023), .ZN(n4220) );
  NAND2_X1 U5203 ( .A1(n4227), .A2(n4228), .ZN(n4242) );
  XNOR2_X1 U5204 ( .A(n4242), .B(n4241), .ZN(n4218) );
  NAND2_X1 U5205 ( .A1(n4348), .A2(n4676), .ZN(n4221) );
  INV_X1 U5206 ( .A(n4221), .ZN(n4217) );
  AOI21_X1 U5207 ( .B1(n4218), .B2(n4413), .A(n4217), .ZN(n4219) );
  NAND2_X1 U5208 ( .A1(n6363), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n4236)
         );
  INV_X1 U5209 ( .A(n4023), .ZN(n4245) );
  OAI21_X1 U5210 ( .B1(n6679), .B2(n4228), .A(n4221), .ZN(n4222) );
  INV_X1 U5211 ( .A(n4222), .ZN(n4223) );
  OAI21_X2 U5212 ( .B1(n4547), .B2(n4245), .A(n4223), .ZN(n4480) );
  NAND2_X1 U5213 ( .A1(n4480), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4224)
         );
  NAND2_X1 U5214 ( .A1(n4224), .A2(n4574), .ZN(n4226) );
  AND2_X1 U5215 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4225) );
  NAND2_X1 U5216 ( .A1(n4480), .A2(n4225), .ZN(n4234) );
  NAND2_X1 U5217 ( .A1(n4023), .A2(n4651), .ZN(n4233) );
  OAI21_X1 U5218 ( .B1(n4228), .B2(n4227), .A(n4242), .ZN(n4230) );
  INV_X1 U5219 ( .A(n4352), .ZN(n4229) );
  OAI211_X1 U5220 ( .C1(n4230), .C2(n6679), .A(n4229), .B(n5492), .ZN(n4231)
         );
  INV_X1 U5221 ( .A(n4231), .ZN(n4232) );
  NAND2_X1 U5222 ( .A1(n4233), .A2(n4232), .ZN(n4512) );
  INV_X1 U5223 ( .A(n4234), .ZN(n4235) );
  AOI21_X1 U5224 ( .B1(n4512), .B2(n3186), .A(n4235), .ZN(n6362) );
  NAND2_X1 U5225 ( .A1(n4236), .A2(n6362), .ZN(n4240) );
  INV_X1 U5226 ( .A(n6363), .ZN(n4238) );
  NAND2_X1 U5227 ( .A1(n4238), .A2(n4237), .ZN(n4239) );
  NAND2_X1 U5228 ( .A1(n4242), .A2(n4241), .ZN(n4251) );
  XNOR2_X1 U5229 ( .A(n4251), .B(n4250), .ZN(n4243) );
  OR2_X1 U5230 ( .A1(n4243), .A2(n6679), .ZN(n4244) );
  OAI21_X2 U5231 ( .B1(n4246), .B2(n4245), .A(n4244), .ZN(n4247) );
  XNOR2_X1 U5232 ( .A(n4247), .B(n6408), .ZN(n6352) );
  NAND2_X1 U5233 ( .A1(n6354), .A2(n6352), .ZN(n6353) );
  NAND2_X1 U5234 ( .A1(n4247), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4248)
         );
  NAND2_X1 U5235 ( .A1(n6353), .A2(n4248), .ZN(n4695) );
  NAND2_X1 U5236 ( .A1(n4249), .A2(n4023), .ZN(n4254) );
  NAND2_X1 U5237 ( .A1(n4251), .A2(n4250), .ZN(n4269) );
  XNOR2_X1 U5238 ( .A(n4269), .B(n4267), .ZN(n4252) );
  NAND2_X1 U5239 ( .A1(n4252), .A2(n4413), .ZN(n4253) );
  NAND2_X1 U5240 ( .A1(n4254), .A2(n4253), .ZN(n4255) );
  XNOR2_X1 U5241 ( .A(n4255), .B(n6403), .ZN(n4694) );
  NAND2_X1 U5242 ( .A1(n4695), .A2(n4694), .ZN(n4693) );
  NAND2_X1 U5243 ( .A1(n4255), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4256)
         );
  NAND2_X1 U5244 ( .A1(n4693), .A2(n4256), .ZN(n5681) );
  NAND2_X1 U5245 ( .A1(n4257), .A2(n4023), .ZN(n4262) );
  INV_X1 U5246 ( .A(n4267), .ZN(n4258) );
  OR2_X1 U5247 ( .A1(n4269), .A2(n4258), .ZN(n4259) );
  XNOR2_X1 U5248 ( .A(n4259), .B(n4266), .ZN(n4260) );
  NAND2_X1 U5249 ( .A1(n4260), .A2(n4413), .ZN(n4261) );
  NAND2_X1 U5250 ( .A1(n4262), .A2(n4261), .ZN(n4263) );
  XNOR2_X1 U5251 ( .A(n4263), .B(n5688), .ZN(n5684) );
  NAND2_X1 U5252 ( .A1(n5681), .A2(n5684), .ZN(n5682) );
  NAND2_X1 U5253 ( .A1(n4263), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4264)
         );
  NAND2_X1 U5254 ( .A1(n5682), .A2(n4264), .ZN(n4799) );
  NAND2_X1 U5255 ( .A1(n4265), .A2(n4023), .ZN(n4272) );
  NAND2_X1 U5256 ( .A1(n4267), .A2(n4266), .ZN(n4268) );
  OR2_X1 U5257 ( .A1(n4269), .A2(n4268), .ZN(n4276) );
  XNOR2_X1 U5258 ( .A(n4276), .B(n4277), .ZN(n4270) );
  NAND2_X1 U5259 ( .A1(n4270), .A2(n4413), .ZN(n4271) );
  NAND2_X1 U5260 ( .A1(n4272), .A2(n4271), .ZN(n4273) );
  INV_X1 U5261 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n4808) );
  XNOR2_X1 U5262 ( .A(n4273), .B(n4808), .ZN(n4802) );
  NAND2_X1 U5263 ( .A1(n4799), .A2(n4802), .ZN(n4800) );
  NAND2_X1 U5264 ( .A1(n4273), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n4274)
         );
  NAND2_X1 U5265 ( .A1(n4800), .A2(n4274), .ZN(n6337) );
  NAND2_X1 U5266 ( .A1(n4275), .A2(n4023), .ZN(n4282) );
  INV_X1 U5267 ( .A(n4276), .ZN(n4278) );
  NAND2_X1 U5268 ( .A1(n4278), .A2(n4277), .ZN(n4290) );
  XNOR2_X1 U5269 ( .A(n4290), .B(n4279), .ZN(n4280) );
  NAND2_X1 U5270 ( .A1(n4280), .A2(n4413), .ZN(n4281) );
  NAND2_X1 U5271 ( .A1(n4282), .A2(n4281), .ZN(n4283) );
  XNOR2_X1 U5272 ( .A(n4283), .B(n6390), .ZN(n6340) );
  NAND2_X1 U5273 ( .A1(n6337), .A2(n6340), .ZN(n6338) );
  NAND2_X1 U5274 ( .A1(n4283), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n4284)
         );
  NAND2_X1 U5275 ( .A1(n6338), .A2(n4284), .ZN(n5185) );
  NAND2_X1 U5276 ( .A1(n4023), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4287) );
  NOR2_X1 U5277 ( .A1(n4287), .A2(n4286), .ZN(n4288) );
  NAND2_X4 U5278 ( .A1(n4285), .A2(n4288), .ZN(n4294) );
  OR3_X1 U5279 ( .A1(n4290), .A2(n4289), .A3(n6679), .ZN(n4291) );
  NAND2_X1 U5280 ( .A1(n3174), .A2(n4291), .ZN(n4292) );
  XNOR2_X1 U5281 ( .A(n4292), .B(n5200), .ZN(n5187) );
  NAND2_X1 U5282 ( .A1(n5185), .A2(n5187), .ZN(n5186) );
  NAND2_X1 U5283 ( .A1(n4292), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n4293)
         );
  NAND2_X1 U5284 ( .A1(n3159), .A2(n3168), .ZN(n4297) );
  OR2_X1 U5285 ( .A1(n4294), .A2(n5486), .ZN(n4296) );
  INV_X1 U5286 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n4298) );
  NAND2_X1 U5287 ( .A1(n4294), .A2(n4298), .ZN(n5475) );
  AND2_X1 U5288 ( .A1(n4294), .A2(n5573), .ZN(n4301) );
  OAI21_X2 U5289 ( .B1(n5497), .B2(n4301), .A(n4300), .ZN(n5505) );
  INV_X1 U5290 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n5572) );
  NOR2_X1 U5291 ( .A1(n4294), .A2(n5572), .ZN(n5553) );
  XNOR2_X1 U5292 ( .A(n4294), .B(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5556)
         );
  INV_X1 U5293 ( .A(n5556), .ZN(n4302) );
  OR2_X2 U5294 ( .A1(n5505), .A2(n4303), .ZN(n5564) );
  NAND2_X1 U5295 ( .A1(n4294), .A2(n5572), .ZN(n5554) );
  NAND2_X1 U5296 ( .A1(n4294), .A2(n5574), .ZN(n4304) );
  INV_X1 U5297 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n4306) );
  NAND2_X1 U5298 ( .A1(n5564), .A2(n4305), .ZN(n4308) );
  INV_X1 U5299 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5539) );
  NOR2_X1 U5300 ( .A1(n4294), .A2(n5539), .ZN(n4310) );
  NAND2_X1 U5301 ( .A1(n4294), .A2(n5539), .ZN(n4309) );
  OAI21_X1 U5302 ( .B1(n5537), .B2(n4310), .A(n4309), .ZN(n5913) );
  INV_X1 U5303 ( .A(n5913), .ZN(n4312) );
  INV_X1 U5304 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5923) );
  NAND2_X1 U5305 ( .A1(n4294), .A2(n5923), .ZN(n5922) );
  NAND2_X1 U5306 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n4366) );
  NAND2_X1 U5307 ( .A1(n4294), .A2(n4366), .ZN(n4311) );
  NAND2_X1 U5308 ( .A1(n4312), .A2(n3183), .ZN(n4315) );
  NAND2_X1 U5309 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5617) );
  INV_X1 U5310 ( .A(n5617), .ZN(n5976) );
  AND2_X1 U5311 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n4367) );
  NAND3_X1 U5312 ( .A1(n4294), .A2(n5976), .A3(n4367), .ZN(n4318) );
  INV_X1 U5313 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n6160) );
  INV_X1 U5314 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n6019) );
  NAND3_X1 U5315 ( .A1(n6160), .A2(n5923), .A3(n6019), .ZN(n4313) );
  NAND2_X1 U5316 ( .A1(n6002), .A2(n4313), .ZN(n4314) );
  NAND2_X1 U5317 ( .A1(n4315), .A2(n4314), .ZN(n5616) );
  INV_X1 U5318 ( .A(n5616), .ZN(n4316) );
  NAND2_X1 U5319 ( .A1(n6001), .A2(n4317), .ZN(n5909) );
  XNOR2_X1 U5320 ( .A(n4294), .B(n5994), .ZN(n5908) );
  OAI22_X1 U5321 ( .A1(n5909), .A2(n5908), .B1(n4294), .B2(n5994), .ZN(n5903)
         );
  XNOR2_X1 U5322 ( .A(n6002), .B(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5904)
         );
  NOR2_X1 U5323 ( .A1(n4294), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5895)
         );
  NAND2_X1 U5324 ( .A1(n5902), .A2(n5895), .ZN(n5888) );
  OAI21_X1 U5325 ( .B1(n4315), .B2(n4318), .A(n5888), .ZN(n4319) );
  XNOR2_X1 U5326 ( .A(n4319), .B(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5704)
         );
  NAND2_X1 U5327 ( .A1(n4664), .A2(n6615), .ZN(n4320) );
  NOR2_X1 U5328 ( .A1(READY_N), .A2(n5747), .ZN(n4447) );
  NAND2_X1 U5329 ( .A1(n4320), .A2(n4447), .ZN(n4329) );
  INV_X1 U5330 ( .A(READY_N), .ZN(n7028) );
  AND2_X1 U5331 ( .A1(n4322), .A2(n7028), .ZN(n4325) );
  INV_X1 U5332 ( .A(n5491), .ZN(n4323) );
  NAND2_X1 U5333 ( .A1(n4323), .A2(n4986), .ZN(n4324) );
  AOI21_X1 U5334 ( .B1(n4423), .B2(n4325), .A(n4324), .ZN(n4326) );
  OR2_X1 U5335 ( .A1(n5756), .A2(n4326), .ZN(n4328) );
  MUX2_X1 U5336 ( .A(n4329), .B(n4328), .S(n4327), .Z(n4337) );
  NOR2_X1 U5337 ( .A1(n4429), .A2(n4417), .ZN(n4357) );
  NAND2_X1 U5338 ( .A1(n4429), .A2(n4348), .ZN(n4330) );
  NAND2_X1 U5339 ( .A1(n4330), .A2(n4327), .ZN(n4331) );
  NOR2_X1 U5340 ( .A1(n4332), .A2(n4331), .ZN(n4341) );
  NAND2_X1 U5341 ( .A1(n4333), .A2(n4986), .ZN(n4335) );
  INV_X1 U5342 ( .A(n4612), .ZN(n4334) );
  MUX2_X1 U5343 ( .A(n4335), .B(n6679), .S(n4334), .Z(n4353) );
  AOI21_X1 U5344 ( .B1(n4341), .B2(n4353), .A(n4078), .ZN(n4442) );
  AOI21_X1 U5345 ( .B1(n5756), .B2(n4357), .A(n4442), .ZN(n4336) );
  NAND2_X1 U5346 ( .A1(n4337), .A2(n4336), .ZN(n4338) );
  INV_X1 U5347 ( .A(n4030), .ZN(n4978) );
  NAND2_X1 U5348 ( .A1(n4341), .A2(n4978), .ZN(n4519) );
  INV_X1 U5349 ( .A(n4339), .ZN(n4340) );
  NAND2_X1 U5350 ( .A1(n4341), .A2(n4340), .ZN(n4488) );
  NAND2_X1 U5351 ( .A1(n4519), .A2(n4488), .ZN(n5748) );
  CLKBUF_X1 U5352 ( .A(n4342), .Z(n4343) );
  NAND2_X1 U5353 ( .A1(n4423), .A2(n4102), .ZN(n4345) );
  OAI211_X1 U5354 ( .C1(n4343), .C2(n3305), .A(n4345), .B(n3163), .ZN(n4346)
         );
  NOR2_X1 U5355 ( .A1(n5748), .A2(n4346), .ZN(n4347) );
  NAND2_X1 U5356 ( .A1(n4348), .A2(n4664), .ZN(n4412) );
  OR2_X1 U5357 ( .A1(n4412), .A2(n4668), .ZN(n4443) );
  NAND4_X1 U5358 ( .A1(n4483), .A2(n4443), .A3(n5491), .A4(n4349), .ZN(n4351)
         );
  AOI22_X1 U5359 ( .A1(n4352), .A2(n4351), .B1(n4350), .B2(n5776), .ZN(n4354)
         );
  AND2_X1 U5360 ( .A1(n4354), .A2(n4353), .ZN(n4355) );
  AND2_X1 U5361 ( .A1(n4356), .A2(n4355), .ZN(n4428) );
  INV_X1 U5362 ( .A(n4521), .ZN(n5752) );
  NOR2_X1 U5363 ( .A1(n6390), .A2(n5200), .ZN(n5485) );
  NAND3_X1 U5364 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .A3(n5485), .ZN(n4362) );
  AOI21_X1 U5365 ( .B1(INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .A(INSTADDRPOINTER_REG_2__SCAN_IN), 
        .ZN(n6416) );
  INV_X1 U5366 ( .A(n6416), .ZN(n4805) );
  NOR2_X1 U5367 ( .A1(n6408), .A2(n6403), .ZN(n6392) );
  NAND2_X1 U5368 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n6392), .ZN(n4807)
         );
  NOR2_X1 U5369 ( .A1(n4808), .A2(n4807), .ZN(n4361) );
  NAND2_X1 U5370 ( .A1(n4805), .A2(n4361), .ZN(n5194) );
  OR2_X1 U5371 ( .A1(n4362), .A2(n5194), .ZN(n4381) );
  OR2_X1 U5372 ( .A1(n4425), .A2(n4986), .ZN(n4358) );
  AND2_X1 U5373 ( .A1(n4428), .A2(n4358), .ZN(n4359) );
  NOR2_X1 U5374 ( .A1(n4375), .A2(n4359), .ZN(n5575) );
  INV_X1 U5375 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n5736) );
  NAND2_X1 U5376 ( .A1(n5575), .A2(n5736), .ZN(n4360) );
  AND2_X1 U5377 ( .A1(n4375), .A2(n6393), .ZN(n4569) );
  INV_X1 U5378 ( .A(n4569), .ZN(n4481) );
  NAND2_X1 U5379 ( .A1(n4078), .A2(n4664), .ZN(n5661) );
  NOR2_X1 U5380 ( .A1(n4237), .A2(n4574), .ZN(n6415) );
  NAND2_X1 U5381 ( .A1(n6415), .A2(n4361), .ZN(n5198) );
  NOR2_X1 U5382 ( .A1(n5198), .A2(n4362), .ZN(n4382) );
  INV_X1 U5383 ( .A(n4382), .ZN(n4363) );
  NAND2_X1 U5384 ( .A1(n5199), .A2(n4363), .ZN(n4364) );
  NAND2_X1 U5385 ( .A1(n5195), .A2(n4364), .ZN(n4369) );
  AOI21_X1 U5386 ( .B1(n6414), .B2(n4381), .A(n4369), .ZN(n5579) );
  NAND3_X1 U5387 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_12__SCAN_IN), .A3(INSTADDRPOINTER_REG_13__SCAN_IN), 
        .ZN(n5586) );
  NOR2_X1 U5388 ( .A1(n4306), .A2(n5586), .ZN(n6169) );
  NAND3_X1 U5389 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .A3(n6169), .ZN(n4383) );
  NOR2_X1 U5390 ( .A1(n6160), .A2(n4383), .ZN(n6012) );
  INV_X1 U5391 ( .A(n6012), .ZN(n5991) );
  NAND2_X1 U5392 ( .A1(n5633), .A2(n5991), .ZN(n4365) );
  NAND2_X1 U5393 ( .A1(n5579), .A2(n4365), .ZN(n6159) );
  INV_X1 U5394 ( .A(n4366), .ZN(n4368) );
  NAND2_X1 U5395 ( .A1(n4368), .A2(n4367), .ZN(n4384) );
  OR2_X1 U5396 ( .A1(n6159), .A2(n4384), .ZN(n4371) );
  OR2_X1 U5397 ( .A1(INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n5577), .ZN(n4573)
         );
  NOR2_X1 U5398 ( .A1(n6420), .A2(n6414), .ZN(n5626) );
  INV_X1 U5399 ( .A(n4369), .ZN(n4370) );
  NAND2_X1 U5400 ( .A1(n5626), .A2(n4370), .ZN(n5992) );
  NAND2_X1 U5401 ( .A1(n4371), .A2(n5992), .ZN(n5973) );
  NAND2_X1 U5402 ( .A1(n5633), .A2(n5617), .ZN(n4372) );
  AND2_X1 U5403 ( .A1(n5973), .A2(n4372), .ZN(n5630) );
  INV_X1 U5404 ( .A(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5613) );
  NAND2_X1 U5405 ( .A1(n4423), .A2(n4413), .ZN(n6587) );
  OAI21_X1 U5406 ( .B1(n4343), .B2(n4672), .A(n6587), .ZN(n4373) );
  INV_X1 U5407 ( .A(n4373), .ZN(n4374) );
  INV_X1 U5408 ( .A(n4377), .ZN(n5852) );
  INV_X1 U5409 ( .A(n4378), .ZN(n4379) );
  OAI21_X1 U5410 ( .B1(n4376), .B2(n5852), .A(n4379), .ZN(n4380) );
  NAND2_X1 U5411 ( .A1(n4380), .A2(n5843), .ZN(n5808) );
  NOR2_X1 U5412 ( .A1(n5687), .A2(n4381), .ZN(n5576) );
  NOR2_X1 U5413 ( .A1(n6186), .A2(n4383), .ZN(n6161) );
  INV_X1 U5414 ( .A(n4384), .ZN(n4385) );
  NAND3_X1 U5415 ( .A1(n5975), .A2(n5976), .A3(n5613), .ZN(n4386) );
  NAND2_X1 U5416 ( .A1(n6371), .A2(REIP_REG_23__SCAN_IN), .ZN(n5701) );
  OAI211_X1 U5417 ( .C1(n6395), .C2(n5808), .A(n4386), .B(n5701), .ZN(n4387)
         );
  INV_X1 U5418 ( .A(n4387), .ZN(n4388) );
  NAND3_X1 U5419 ( .A1(n3175), .A2(n3184), .A3(n4388), .ZN(U2995) );
  NAND2_X1 U5420 ( .A1(n5756), .A2(n4521), .ZN(n4446) );
  NAND2_X1 U5421 ( .A1(n5731), .A2(n3305), .ZN(n4391) );
  OR2_X1 U5422 ( .A1(n4392), .A2(n4391), .ZN(n4607) );
  INV_X1 U5423 ( .A(n4607), .ZN(n4393) );
  NAND3_X1 U5424 ( .A1(n4393), .A2(n3156), .A3(n4102), .ZN(n4394) );
  NAND2_X1 U5425 ( .A1(n4446), .A2(n4394), .ZN(n4395) );
  NAND2_X1 U5426 ( .A1(n6292), .A2(n3324), .ZN(n5836) );
  INV_X1 U5427 ( .A(n5774), .ZN(n4399) );
  INV_X1 U5428 ( .A(n4400), .ZN(n4402) );
  AOI211_X1 U5429 ( .C1(n5776), .C2(n5774), .A(n4402), .B(n4401), .ZN(n4403)
         );
  NOR2_X1 U5430 ( .A1(n4404), .A2(n4403), .ZN(n5766) );
  INV_X1 U5431 ( .A(EBX_REG_30__SCAN_IN), .ZN(n5761) );
  NAND2_X1 U5432 ( .A1(n4405), .A2(EBX_REG_30__SCAN_IN), .ZN(n4406) );
  NOR2_X2 U5433 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATE2_REG_3__SCAN_IN), .ZN(
        n6484) );
  INV_X1 U5434 ( .A(n6484), .ZN(n6498) );
  NOR2_X1 U5435 ( .A1(n6498), .A2(STATE2_REG_1__SCAN_IN), .ZN(n6187) );
  INV_X1 U5436 ( .A(n4419), .ZN(n4416) );
  AOI211_X1 U5437 ( .C1(MEMORYFETCH_REG_SCAN_IN), .C2(n4410), .A(n6187), .B(
        n4416), .ZN(n4411) );
  INV_X1 U5438 ( .A(n4411), .ZN(U2788) );
  INV_X1 U5439 ( .A(n6675), .ZN(n4415) );
  INV_X1 U5440 ( .A(n4412), .ZN(n4980) );
  OR2_X1 U5441 ( .A1(n4413), .A2(n4980), .ZN(n5757) );
  OAI21_X1 U5442 ( .B1(n6187), .B2(READREQUEST_REG_SCAN_IN), .A(n4415), .ZN(
        n4414) );
  OAI21_X1 U5443 ( .B1(n4415), .B2(n5757), .A(n4414), .ZN(U3474) );
  OR2_X1 U5444 ( .A1(n4419), .A2(n4664), .ZN(n4502) );
  INV_X1 U5445 ( .A(EAX_REG_15__SCAN_IN), .ZN(n4421) );
  INV_X1 U5446 ( .A(LWORD_REG_15__SCAN_IN), .ZN(n4420) );
  OAI21_X1 U5447 ( .B1(n4417), .B2(n7028), .A(n4416), .ZN(n4507) );
  INV_X1 U5448 ( .A(n4507), .ZN(n4578) );
  NAND2_X1 U5449 ( .A1(n4664), .A2(n7028), .ZN(n4418) );
  INV_X1 U5450 ( .A(DATAI_15_), .ZN(n6795) );
  OAI222_X1 U5451 ( .A1(n4502), .A2(n4421), .B1(n4420), .B2(n4578), .C1(n4610), 
        .C2(n6795), .ZN(U2954) );
  INV_X1 U5452 ( .A(n6023), .ZN(n4982) );
  INV_X1 U5453 ( .A(n4423), .ZN(n4438) );
  INV_X1 U5454 ( .A(n4424), .ZN(n4426) );
  AND4_X1 U5455 ( .A1(n3163), .A2(n4438), .A3(n4426), .A4(n4425), .ZN(n4427)
         );
  NAND2_X1 U5456 ( .A1(n4428), .A2(n4427), .ZN(n5658) );
  NAND2_X1 U5457 ( .A1(n4982), .A2(n5658), .ZN(n4433) );
  INV_X1 U5458 ( .A(n4429), .ZN(n5657) );
  CLKBUF_X1 U5459 ( .A(n4430), .Z(n4435) );
  INV_X1 U5460 ( .A(n4435), .ZN(n5737) );
  INV_X1 U5461 ( .A(n4431), .ZN(n4436) );
  NAND3_X1 U5462 ( .A1(n5657), .A2(n5737), .A3(n4436), .ZN(n4432) );
  OAI211_X1 U5463 ( .C1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .C2(n5661), .A(n4433), .B(n4432), .ZN(n6562) );
  NOR2_X1 U5464 ( .A1(n6600), .A2(n5736), .ZN(n4437) );
  INV_X1 U5465 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n4434) );
  AOI22_X1 U5466 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n4434), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n4574), .ZN(n5735) );
  NOR2_X1 U5467 ( .A1(n5738), .A2(n4435), .ZN(n5722) );
  AOI222_X1 U5468 ( .A1(n6562), .A2(n6597), .B1(n4437), .B2(n5735), .C1(n4436), 
        .C2(n5722), .ZN(n4456) );
  NAND2_X1 U5469 ( .A1(n5661), .A2(n4438), .ZN(n4440) );
  AOI21_X1 U5470 ( .B1(n4168), .B2(n6615), .A(READY_N), .ZN(n4439) );
  NAND2_X1 U5471 ( .A1(n4440), .A2(n4439), .ZN(n4441) );
  OR2_X1 U5472 ( .A1(n5756), .A2(n4441), .ZN(n4445) );
  INV_X1 U5473 ( .A(n4442), .ZN(n4444) );
  NAND4_X1 U5474 ( .A1(n4446), .A2(n4445), .A3(n4444), .A4(n4443), .ZN(n4451)
         );
  OR2_X1 U5475 ( .A1(n5756), .A2(n4519), .ZN(n4450) );
  INV_X1 U5476 ( .A(n4447), .ZN(n4448) );
  OR2_X1 U5477 ( .A1(n3163), .A2(n4448), .ZN(n4449) );
  NAND2_X1 U5478 ( .A1(n4450), .A2(n4449), .ZN(n4609) );
  NAND2_X1 U5479 ( .A1(n6561), .A2(n6583), .ZN(n4454) );
  NOR2_X1 U5480 ( .A1(n6600), .A2(n6590), .ZN(n4545) );
  NAND2_X1 U5481 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n4545), .ZN(n6663) );
  INV_X1 U5482 ( .A(n6663), .ZN(n4452) );
  NAND2_X1 U5483 ( .A1(FLUSH_REG_SCAN_IN), .A2(n4452), .ZN(n4453) );
  NAND2_X1 U5484 ( .A1(n4454), .A2(n4453), .ZN(n4460) );
  NOR2_X1 U5485 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n6666), .ZN(n6662) );
  NOR2_X1 U5486 ( .A1(n4460), .A2(n6662), .ZN(n5743) );
  NAND2_X1 U5487 ( .A1(n5743), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4455) );
  OAI21_X1 U5488 ( .B1(n4456), .B2(n5743), .A(n4455), .ZN(U3460) );
  INV_X1 U5489 ( .A(n6445), .ZN(n5091) );
  NOR2_X1 U5490 ( .A1(n4457), .A2(n5091), .ZN(n4458) );
  XNOR2_X1 U5491 ( .A(n4458), .B(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n5288)
         );
  OR2_X1 U5492 ( .A1(n3163), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4459) );
  OR2_X1 U5493 ( .A1(n5288), .A2(n4459), .ZN(n4537) );
  NAND2_X1 U5494 ( .A1(n4460), .A2(n6666), .ZN(n4461) );
  INV_X1 U5495 ( .A(n5743), .ZN(n5664) );
  OAI22_X1 U5496 ( .A1(n4537), .A2(n4461), .B1(n5664), .B2(n3524), .ZN(U3455)
         );
  INV_X1 U5497 ( .A(EAX_REG_25__SCAN_IN), .ZN(n4467) );
  AND2_X1 U5498 ( .A1(n5661), .A2(n6587), .ZN(n4464) );
  NAND2_X1 U5499 ( .A1(n4462), .A2(n6583), .ZN(n4463) );
  NAND2_X1 U5500 ( .A1(n4465), .A2(n4986), .ZN(n4631) );
  NAND2_X1 U5501 ( .A1(n4545), .A2(n6596), .ZN(n6584) );
  INV_X2 U5502 ( .A(n6584), .ZN(n6333) );
  AOI22_X1 U5503 ( .A1(n6333), .A2(UWORD_REG_9__SCAN_IN), .B1(n6332), .B2(
        DATAO_REG_25__SCAN_IN), .ZN(n4466) );
  OAI21_X1 U5504 ( .B1(n4467), .B2(n4631), .A(n4466), .ZN(U2898) );
  INV_X1 U5505 ( .A(EAX_REG_26__SCAN_IN), .ZN(n4469) );
  AOI22_X1 U5506 ( .A1(n6333), .A2(UWORD_REG_10__SCAN_IN), .B1(n6332), .B2(
        DATAO_REG_26__SCAN_IN), .ZN(n4468) );
  OAI21_X1 U5507 ( .B1(n4469), .B2(n4631), .A(n4468), .ZN(U2897) );
  INV_X1 U5508 ( .A(EAX_REG_24__SCAN_IN), .ZN(n4471) );
  AOI22_X1 U5509 ( .A1(n6333), .A2(UWORD_REG_8__SCAN_IN), .B1(n6332), .B2(
        DATAO_REG_24__SCAN_IN), .ZN(n4470) );
  OAI21_X1 U5510 ( .B1(n4471), .B2(n4631), .A(n4470), .ZN(U2899) );
  INV_X1 U5511 ( .A(EAX_REG_28__SCAN_IN), .ZN(n4473) );
  AOI22_X1 U5512 ( .A1(n6333), .A2(UWORD_REG_12__SCAN_IN), .B1(n6332), .B2(
        DATAO_REG_28__SCAN_IN), .ZN(n4472) );
  OAI21_X1 U5513 ( .B1(n4473), .B2(n4631), .A(n4472), .ZN(U2895) );
  INV_X1 U5514 ( .A(EAX_REG_29__SCAN_IN), .ZN(n4475) );
  AOI22_X1 U5515 ( .A1(n6333), .A2(UWORD_REG_13__SCAN_IN), .B1(n6332), .B2(
        DATAO_REG_29__SCAN_IN), .ZN(n4474) );
  OAI21_X1 U5516 ( .B1(n4475), .B2(n4631), .A(n4474), .ZN(U2894) );
  INV_X1 U5517 ( .A(EAX_REG_27__SCAN_IN), .ZN(n4477) );
  AOI22_X1 U5518 ( .A1(n6333), .A2(UWORD_REG_11__SCAN_IN), .B1(n6332), .B2(
        DATAO_REG_27__SCAN_IN), .ZN(n4476) );
  OAI21_X1 U5519 ( .B1(n4477), .B2(n4631), .A(n4476), .ZN(U2896) );
  INV_X1 U5520 ( .A(EAX_REG_30__SCAN_IN), .ZN(n4479) );
  AOI22_X1 U5521 ( .A1(n6333), .A2(UWORD_REG_14__SCAN_IN), .B1(n6332), .B2(
        DATAO_REG_30__SCAN_IN), .ZN(n4478) );
  OAI21_X1 U5522 ( .B1(n4479), .B2(n4631), .A(n4478), .ZN(U2893) );
  XNOR2_X1 U5523 ( .A(n4480), .B(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4501)
         );
  INV_X1 U5524 ( .A(n5577), .ZN(n4482) );
  NAND2_X1 U5525 ( .A1(n4482), .A2(n4481), .ZN(n4486) );
  NAND2_X1 U5526 ( .A1(n4483), .A2(n5736), .ZN(n4484) );
  NAND2_X1 U5527 ( .A1(n3182), .A2(n4484), .ZN(n5229) );
  INV_X1 U5528 ( .A(REIP_REG_0__SCAN_IN), .ZN(n6672) );
  OAI22_X1 U5529 ( .A1(n6395), .A2(n5229), .B1(n6672), .B2(n6393), .ZN(n4485)
         );
  NOR2_X1 U5530 ( .A1(n6414), .A2(n5575), .ZN(n5580) );
  NOR2_X1 U5531 ( .A1(n5580), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4568)
         );
  AOI211_X1 U5532 ( .C1(INSTADDRPOINTER_REG_0__SCAN_IN), .C2(n4486), .A(n4485), 
        .B(n4568), .ZN(n4487) );
  OAI21_X1 U5533 ( .B1(n4501), .B2(n6398), .A(n4487), .ZN(U3018) );
  OR2_X1 U5534 ( .A1(n5756), .A2(n4488), .ZN(n6574) );
  OAI21_X1 U5535 ( .B1(n4491), .B2(n4490), .A(n4489), .ZN(n5236) );
  INV_X1 U5536 ( .A(n5236), .ZN(n4499) );
  NAND3_X1 U5537 ( .A1(n6596), .A2(STATEBS16_REG_SCAN_IN), .A3(
        STATE2_REG_1__SCAN_IN), .ZN(n6610) );
  INV_X1 U5538 ( .A(n6610), .ZN(n4492) );
  NAND2_X1 U5539 ( .A1(n4492), .A2(n6484), .ZN(n5930) );
  INV_X2 U5540 ( .A(n5930), .ZN(n6357) );
  NAND2_X1 U5541 ( .A1(n6498), .A2(n4493), .ZN(n6676) );
  NAND2_X1 U5542 ( .A1(n6676), .A2(n6596), .ZN(n4494) );
  NAND2_X1 U5543 ( .A1(n6596), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4496) );
  NAND2_X1 U5544 ( .A1(n7056), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4495) );
  NAND2_X1 U5545 ( .A1(n4496), .A2(n4495), .ZN(n4513) );
  OAI21_X1 U5546 ( .B1(n6361), .B2(n4513), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n4497) );
  OAI21_X1 U5547 ( .B1(n6672), .B2(n6393), .A(n4497), .ZN(n4498) );
  AOI21_X1 U5548 ( .B1(n4499), .B2(n6357), .A(n4498), .ZN(n4500) );
  OAI21_X1 U5549 ( .B1(n4501), .B2(n6195), .A(n4500), .ZN(U2986) );
  INV_X2 U5550 ( .A(n4502), .ZN(n4603) );
  AOI22_X1 U5551 ( .A1(LWORD_REG_4__SCAN_IN), .A2(n4507), .B1(n4603), .B2(
        EAX_REG_4__SCAN_IN), .ZN(n4503) );
  NAND2_X1 U5552 ( .A1(n4579), .A2(DATAI_4_), .ZN(n4587) );
  NAND2_X1 U5553 ( .A1(n4503), .A2(n4587), .ZN(U2943) );
  AOI22_X1 U5554 ( .A1(LWORD_REG_11__SCAN_IN), .A2(n4507), .B1(n4603), .B2(
        EAX_REG_11__SCAN_IN), .ZN(n4504) );
  NAND2_X1 U5555 ( .A1(n4579), .A2(DATAI_11_), .ZN(n4561) );
  NAND2_X1 U5556 ( .A1(n4504), .A2(n4561), .ZN(U2950) );
  AOI22_X1 U5557 ( .A1(LWORD_REG_6__SCAN_IN), .A2(n4507), .B1(n4603), .B2(
        EAX_REG_6__SCAN_IN), .ZN(n4505) );
  NAND2_X1 U5558 ( .A1(n4579), .A2(DATAI_6_), .ZN(n4591) );
  NAND2_X1 U5559 ( .A1(n4505), .A2(n4591), .ZN(U2945) );
  AOI22_X1 U5560 ( .A1(LWORD_REG_5__SCAN_IN), .A2(n4507), .B1(n4603), .B2(
        EAX_REG_5__SCAN_IN), .ZN(n4506) );
  NAND2_X1 U5561 ( .A1(n4579), .A2(DATAI_5_), .ZN(n4589) );
  NAND2_X1 U5562 ( .A1(n4506), .A2(n4589), .ZN(U2944) );
  AOI22_X1 U5563 ( .A1(LWORD_REG_3__SCAN_IN), .A2(n4507), .B1(n4603), .B2(
        EAX_REG_3__SCAN_IN), .ZN(n4508) );
  NAND2_X1 U5564 ( .A1(n4579), .A2(DATAI_3_), .ZN(n4604) );
  NAND2_X1 U5565 ( .A1(n4508), .A2(n4604), .ZN(U2942) );
  INV_X1 U5566 ( .A(n3474), .ZN(n4510) );
  OAI21_X1 U5567 ( .B1(n4511), .B2(n4509), .A(n4510), .ZN(n4996) );
  XOR2_X1 U5568 ( .A(n3186), .B(n4512), .Z(n4567) );
  NAND2_X1 U5569 ( .A1(n4567), .A2(n6366), .ZN(n4516) );
  INV_X1 U5570 ( .A(REIP_REG_1__SCAN_IN), .ZN(n6667) );
  NOR2_X1 U5571 ( .A1(n6393), .A2(n6667), .ZN(n4572) );
  NOR2_X1 U5572 ( .A1(n6370), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n4514)
         );
  AOI211_X1 U5573 ( .C1(n6361), .C2(PHYADDRPOINTER_REG_1__SCAN_IN), .A(n4572), 
        .B(n4514), .ZN(n4515) );
  OAI211_X1 U5574 ( .C1(n5930), .C2(n4996), .A(n4516), .B(n4515), .ZN(U2985)
         );
  XNOR2_X1 U5575 ( .A(n4518), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4524)
         );
  INV_X1 U5576 ( .A(n4519), .ZN(n4520) );
  OR2_X1 U5577 ( .A1(n4521), .A2(n4520), .ZN(n4532) );
  NAND2_X1 U5578 ( .A1(n5737), .A2(n5741), .ZN(n4528) );
  XNOR2_X1 U5579 ( .A(n4528), .B(n3165), .ZN(n4522) );
  NAND2_X1 U5580 ( .A1(n4532), .A2(n4522), .ZN(n4523) );
  OAI21_X1 U5581 ( .B1(n4524), .B2(n5661), .A(n4523), .ZN(n4525) );
  AOI21_X1 U5582 ( .B1(n5414), .B2(n5658), .A(n4525), .ZN(n5721) );
  INV_X1 U5583 ( .A(n5658), .ZN(n4534) );
  OAI21_X1 U5584 ( .B1(n5741), .B2(n5737), .A(n4528), .ZN(n4531) );
  XNOR2_X1 U5585 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4529) );
  NOR2_X1 U5586 ( .A1(n5661), .A2(n4529), .ZN(n4530) );
  AOI21_X1 U5587 ( .B1(n4532), .B2(n4531), .A(n4530), .ZN(n4533) );
  OAI21_X1 U5588 ( .B1(n4527), .B2(n4534), .A(n4533), .ZN(n6568) );
  NAND3_X1 U5589 ( .A1(n6568), .A2(n6600), .A3(n6561), .ZN(n4541) );
  INV_X1 U5590 ( .A(FLUSH_REG_SCAN_IN), .ZN(n7080) );
  NAND2_X1 U5591 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n7080), .ZN(n4535) );
  OAI21_X1 U5592 ( .B1(n6561), .B2(STATE2_REG_1__SCAN_IN), .A(n4535), .ZN(
        n4539) );
  NAND2_X1 U5593 ( .A1(n4539), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4536) );
  AND2_X1 U5594 ( .A1(n4537), .A2(n4536), .ZN(n4542) );
  NAND2_X1 U5595 ( .A1(n4539), .A2(n4538), .ZN(n4540) );
  OAI211_X1 U5596 ( .C1(n5721), .C2(n4541), .A(n4542), .B(n4540), .ZN(n6577)
         );
  NAND2_X1 U5597 ( .A1(n4542), .A2(n4431), .ZN(n4543) );
  NAND2_X1 U5598 ( .A1(n6577), .A2(n4543), .ZN(n4546) );
  AOI21_X1 U5599 ( .B1(n4546), .B2(n7080), .A(n6663), .ZN(n4544) );
  INV_X1 U5600 ( .A(n6607), .ZN(n6680) );
  OR2_X1 U5601 ( .A1(n4544), .A2(n4820), .ZN(n6425) );
  NAND2_X1 U5602 ( .A1(n4546), .A2(n4545), .ZN(n6595) );
  INV_X1 U5603 ( .A(n6595), .ZN(n4549) );
  NOR2_X1 U5604 ( .A1(STATE2_REG_3__SCAN_IN), .A2(n6600), .ZN(n6032) );
  OAI22_X1 U5605 ( .A1(n5237), .A2(n6498), .B1(n3463), .B2(n6032), .ZN(n4548)
         );
  OAI21_X1 U5606 ( .B1(n4549), .B2(n4548), .A(n6425), .ZN(n4550) );
  OAI21_X1 U5607 ( .B1(n6425), .B2(n6558), .A(n4550), .ZN(U3465) );
  AOI22_X1 U5608 ( .A1(LWORD_REG_2__SCAN_IN), .A2(n4565), .B1(n4603), .B2(
        EAX_REG_2__SCAN_IN), .ZN(n4551) );
  NAND2_X1 U5609 ( .A1(n4579), .A2(DATAI_2_), .ZN(n4583) );
  NAND2_X1 U5610 ( .A1(n4551), .A2(n4583), .ZN(U2941) );
  AOI22_X1 U5611 ( .A1(LWORD_REG_1__SCAN_IN), .A2(n4565), .B1(n4603), .B2(
        EAX_REG_1__SCAN_IN), .ZN(n4552) );
  NAND2_X1 U5612 ( .A1(n4579), .A2(DATAI_1_), .ZN(n4585) );
  NAND2_X1 U5613 ( .A1(n4552), .A2(n4585), .ZN(U2940) );
  AOI22_X1 U5614 ( .A1(UWORD_REG_13__SCAN_IN), .A2(n4565), .B1(n4603), .B2(
        EAX_REG_29__SCAN_IN), .ZN(n4553) );
  NAND2_X1 U5615 ( .A1(n4579), .A2(DATAI_13_), .ZN(n4563) );
  NAND2_X1 U5616 ( .A1(n4553), .A2(n4563), .ZN(U2937) );
  AOI22_X1 U5617 ( .A1(UWORD_REG_14__SCAN_IN), .A2(n4565), .B1(n4603), .B2(
        EAX_REG_30__SCAN_IN), .ZN(n4554) );
  INV_X1 U5618 ( .A(DATAI_14_), .ZN(n5345) );
  OR2_X1 U5619 ( .A1(n4610), .A2(n5345), .ZN(n4581) );
  NAND2_X1 U5620 ( .A1(n4554), .A2(n4581), .ZN(U2938) );
  AOI22_X1 U5621 ( .A1(UWORD_REG_9__SCAN_IN), .A2(n4565), .B1(n4603), .B2(
        EAX_REG_25__SCAN_IN), .ZN(n4555) );
  NAND2_X1 U5622 ( .A1(n4579), .A2(DATAI_9_), .ZN(n4558) );
  NAND2_X1 U5623 ( .A1(n4555), .A2(n4558), .ZN(U2933) );
  AOI22_X1 U5624 ( .A1(LWORD_REG_7__SCAN_IN), .A2(n4565), .B1(n4603), .B2(
        EAX_REG_7__SCAN_IN), .ZN(n4556) );
  NAND2_X1 U5625 ( .A1(n4579), .A2(DATAI_7_), .ZN(n4593) );
  NAND2_X1 U5626 ( .A1(n4556), .A2(n4593), .ZN(U2946) );
  AOI22_X1 U5627 ( .A1(UWORD_REG_10__SCAN_IN), .A2(n4565), .B1(n4603), .B2(
        EAX_REG_26__SCAN_IN), .ZN(n4557) );
  INV_X1 U5628 ( .A(DATAI_10_), .ZN(n5330) );
  OR2_X1 U5629 ( .A1(n4610), .A2(n5330), .ZN(n4599) );
  NAND2_X1 U5630 ( .A1(n4557), .A2(n4599), .ZN(U2934) );
  AOI22_X1 U5631 ( .A1(LWORD_REG_9__SCAN_IN), .A2(n4565), .B1(n4603), .B2(
        EAX_REG_9__SCAN_IN), .ZN(n4559) );
  NAND2_X1 U5632 ( .A1(n4559), .A2(n4558), .ZN(U2948) );
  AOI22_X1 U5633 ( .A1(UWORD_REG_12__SCAN_IN), .A2(n4565), .B1(n4603), .B2(
        EAX_REG_28__SCAN_IN), .ZN(n4560) );
  NAND2_X1 U5634 ( .A1(n4579), .A2(DATAI_12_), .ZN(n4597) );
  NAND2_X1 U5635 ( .A1(n4560), .A2(n4597), .ZN(U2936) );
  AOI22_X1 U5636 ( .A1(UWORD_REG_11__SCAN_IN), .A2(n4565), .B1(n4603), .B2(
        EAX_REG_27__SCAN_IN), .ZN(n4562) );
  NAND2_X1 U5637 ( .A1(n4562), .A2(n4561), .ZN(U2935) );
  AOI22_X1 U5638 ( .A1(LWORD_REG_13__SCAN_IN), .A2(n4565), .B1(n4603), .B2(
        EAX_REG_13__SCAN_IN), .ZN(n4564) );
  NAND2_X1 U5639 ( .A1(n4564), .A2(n4563), .ZN(U2952) );
  AOI22_X1 U5640 ( .A1(LWORD_REG_0__SCAN_IN), .A2(n4565), .B1(n4603), .B2(
        EAX_REG_0__SCAN_IN), .ZN(n4566) );
  NAND2_X1 U5641 ( .A1(n4579), .A2(DATAI_0_), .ZN(n4601) );
  NAND2_X1 U5642 ( .A1(n4566), .A2(n4601), .ZN(U2939) );
  INV_X1 U5643 ( .A(n4567), .ZN(n4577) );
  XNOR2_X1 U5644 ( .A(n4981), .B(n4102), .ZN(n4615) );
  OAI21_X1 U5645 ( .B1(n4569), .B2(n4568), .A(INSTADDRPOINTER_REG_1__SCAN_IN), 
        .ZN(n4570) );
  INV_X1 U5646 ( .A(n4570), .ZN(n4571) );
  AOI211_X1 U5647 ( .C1(n6412), .C2(n4615), .A(n4572), .B(n4571), .ZN(n4576)
         );
  NAND3_X1 U5648 ( .A1(n5633), .A2(n4574), .A3(n4573), .ZN(n4575) );
  OAI211_X1 U5649 ( .C1(n4577), .C2(n6398), .A(n4576), .B(n4575), .ZN(U3017)
         );
  AOI22_X1 U5650 ( .A1(UWORD_REG_8__SCAN_IN), .A2(n4565), .B1(n4603), .B2(
        EAX_REG_24__SCAN_IN), .ZN(n4580) );
  NAND2_X1 U5651 ( .A1(n4579), .A2(DATAI_8_), .ZN(n4595) );
  NAND2_X1 U5652 ( .A1(n4580), .A2(n4595), .ZN(U2932) );
  AOI22_X1 U5653 ( .A1(LWORD_REG_14__SCAN_IN), .A2(n4565), .B1(n4603), .B2(
        EAX_REG_14__SCAN_IN), .ZN(n4582) );
  NAND2_X1 U5654 ( .A1(n4582), .A2(n4581), .ZN(U2953) );
  AOI22_X1 U5655 ( .A1(UWORD_REG_2__SCAN_IN), .A2(n4507), .B1(n4603), .B2(
        EAX_REG_18__SCAN_IN), .ZN(n4584) );
  NAND2_X1 U5656 ( .A1(n4584), .A2(n4583), .ZN(U2926) );
  AOI22_X1 U5657 ( .A1(UWORD_REG_1__SCAN_IN), .A2(n4507), .B1(n4603), .B2(
        EAX_REG_17__SCAN_IN), .ZN(n4586) );
  NAND2_X1 U5658 ( .A1(n4586), .A2(n4585), .ZN(U2925) );
  AOI22_X1 U5659 ( .A1(UWORD_REG_4__SCAN_IN), .A2(n4507), .B1(n4603), .B2(
        EAX_REG_20__SCAN_IN), .ZN(n4588) );
  NAND2_X1 U5660 ( .A1(n4588), .A2(n4587), .ZN(U2928) );
  AOI22_X1 U5661 ( .A1(UWORD_REG_5__SCAN_IN), .A2(n4507), .B1(n4603), .B2(
        EAX_REG_21__SCAN_IN), .ZN(n4590) );
  NAND2_X1 U5662 ( .A1(n4590), .A2(n4589), .ZN(U2929) );
  AOI22_X1 U5663 ( .A1(UWORD_REG_6__SCAN_IN), .A2(n4507), .B1(n4603), .B2(
        EAX_REG_22__SCAN_IN), .ZN(n4592) );
  NAND2_X1 U5664 ( .A1(n4592), .A2(n4591), .ZN(U2930) );
  AOI22_X1 U5665 ( .A1(UWORD_REG_7__SCAN_IN), .A2(n4565), .B1(n4603), .B2(
        EAX_REG_23__SCAN_IN), .ZN(n4594) );
  NAND2_X1 U5666 ( .A1(n4594), .A2(n4593), .ZN(U2931) );
  AOI22_X1 U5667 ( .A1(LWORD_REG_8__SCAN_IN), .A2(n4565), .B1(n4603), .B2(
        EAX_REG_8__SCAN_IN), .ZN(n4596) );
  NAND2_X1 U5668 ( .A1(n4596), .A2(n4595), .ZN(U2947) );
  AOI22_X1 U5669 ( .A1(LWORD_REG_12__SCAN_IN), .A2(n4565), .B1(n4603), .B2(
        EAX_REG_12__SCAN_IN), .ZN(n4598) );
  NAND2_X1 U5670 ( .A1(n4598), .A2(n4597), .ZN(U2951) );
  AOI22_X1 U5671 ( .A1(LWORD_REG_10__SCAN_IN), .A2(n4565), .B1(n4603), .B2(
        EAX_REG_10__SCAN_IN), .ZN(n4600) );
  NAND2_X1 U5672 ( .A1(n4600), .A2(n4599), .ZN(U2949) );
  AOI22_X1 U5673 ( .A1(UWORD_REG_0__SCAN_IN), .A2(n4565), .B1(n4603), .B2(
        EAX_REG_16__SCAN_IN), .ZN(n4602) );
  NAND2_X1 U5674 ( .A1(n4602), .A2(n4601), .ZN(U2924) );
  AOI22_X1 U5675 ( .A1(UWORD_REG_3__SCAN_IN), .A2(n4565), .B1(n4603), .B2(
        EAX_REG_19__SCAN_IN), .ZN(n4605) );
  NAND2_X1 U5676 ( .A1(n4605), .A2(n4604), .ZN(U2927) );
  NOR2_X1 U5677 ( .A1(n4606), .A2(n4607), .ZN(n4608) );
  OAI21_X1 U5678 ( .B1(n4609), .B2(n4608), .A(n6583), .ZN(n4611) );
  NAND2_X1 U5679 ( .A1(n4612), .A2(n3324), .ZN(n4613) );
  INV_X1 U5680 ( .A(n4613), .ZN(n4614) );
  NAND2_X1 U5681 ( .A1(n5860), .A2(n4614), .ZN(n5411) );
  INV_X1 U5682 ( .A(DATAI_0_), .ZN(n6945) );
  INV_X1 U5683 ( .A(EAX_REG_0__SCAN_IN), .ZN(n6336) );
  OAI222_X1 U5684 ( .A1(n5236), .A2(n6114), .B1(n5411), .B2(n6945), .C1(n5860), 
        .C2(n6336), .ZN(U2891) );
  INV_X1 U5685 ( .A(DATAI_1_), .ZN(n6995) );
  INV_X1 U5686 ( .A(EAX_REG_1__SCAN_IN), .ZN(n6331) );
  OAI222_X1 U5687 ( .A1(n4996), .A2(n6114), .B1(n5411), .B2(n6995), .C1(n5860), 
        .C2(n6331), .ZN(U2890) );
  AOI22_X1 U5688 ( .A1(n5846), .A2(n4615), .B1(n4405), .B2(EBX_REG_1__SCAN_IN), 
        .ZN(n4616) );
  OAI21_X1 U5689 ( .B1(n4996), .B2(n5836), .A(n4616), .ZN(U2858) );
  INV_X1 U5690 ( .A(EAX_REG_23__SCAN_IN), .ZN(n4618) );
  AOI22_X1 U5691 ( .A1(n6333), .A2(UWORD_REG_7__SCAN_IN), .B1(n6323), .B2(
        DATAO_REG_23__SCAN_IN), .ZN(n4617) );
  OAI21_X1 U5692 ( .B1(n4618), .B2(n4631), .A(n4617), .ZN(U2900) );
  INV_X1 U5693 ( .A(EAX_REG_18__SCAN_IN), .ZN(n4620) );
  AOI22_X1 U5694 ( .A1(n6333), .A2(UWORD_REG_2__SCAN_IN), .B1(n6323), .B2(
        DATAO_REG_18__SCAN_IN), .ZN(n4619) );
  OAI21_X1 U5695 ( .B1(n4620), .B2(n4631), .A(n4619), .ZN(U2905) );
  INV_X1 U5696 ( .A(EAX_REG_19__SCAN_IN), .ZN(n4622) );
  AOI22_X1 U5697 ( .A1(n6333), .A2(UWORD_REG_3__SCAN_IN), .B1(n6323), .B2(
        DATAO_REG_19__SCAN_IN), .ZN(n4621) );
  OAI21_X1 U5698 ( .B1(n4622), .B2(n4631), .A(n4621), .ZN(U2904) );
  INV_X1 U5699 ( .A(EAX_REG_17__SCAN_IN), .ZN(n4624) );
  AOI22_X1 U5700 ( .A1(n6333), .A2(UWORD_REG_1__SCAN_IN), .B1(n6323), .B2(
        DATAO_REG_17__SCAN_IN), .ZN(n4623) );
  OAI21_X1 U5701 ( .B1(n4624), .B2(n4631), .A(n4623), .ZN(U2906) );
  INV_X1 U5702 ( .A(EAX_REG_20__SCAN_IN), .ZN(n4626) );
  AOI22_X1 U5703 ( .A1(n6333), .A2(UWORD_REG_4__SCAN_IN), .B1(n6323), .B2(
        DATAO_REG_20__SCAN_IN), .ZN(n4625) );
  OAI21_X1 U5704 ( .B1(n4626), .B2(n4631), .A(n4625), .ZN(U2903) );
  INV_X1 U5705 ( .A(EAX_REG_22__SCAN_IN), .ZN(n4628) );
  AOI22_X1 U5706 ( .A1(n6333), .A2(UWORD_REG_6__SCAN_IN), .B1(n6323), .B2(
        DATAO_REG_22__SCAN_IN), .ZN(n4627) );
  OAI21_X1 U5707 ( .B1(n4628), .B2(n4631), .A(n4627), .ZN(U2901) );
  AOI22_X1 U5708 ( .A1(n6333), .A2(UWORD_REG_0__SCAN_IN), .B1(n6323), .B2(
        DATAO_REG_16__SCAN_IN), .ZN(n4629) );
  OAI21_X1 U5709 ( .B1(n3721), .B2(n4631), .A(n4629), .ZN(U2907) );
  INV_X1 U5710 ( .A(EAX_REG_21__SCAN_IN), .ZN(n4632) );
  AOI22_X1 U5711 ( .A1(n6333), .A2(UWORD_REG_5__SCAN_IN), .B1(n6323), .B2(
        DATAO_REG_21__SCAN_IN), .ZN(n4630) );
  OAI21_X1 U5712 ( .B1(n4632), .B2(n4631), .A(n4630), .ZN(U2902) );
  OAI222_X1 U5713 ( .A1(n5229), .A2(n6288), .B1(n6292), .B2(n4633), .C1(n5236), 
        .C2(n5854), .ZN(U2859) );
  NOR2_X1 U5714 ( .A1(n4636), .A2(n4635), .ZN(n4637) );
  NOR2_X1 U5715 ( .A1(n4702), .A2(n4637), .ZN(n6365) );
  INV_X1 U5716 ( .A(n6365), .ZN(n4640) );
  INV_X1 U5717 ( .A(DATAI_2_), .ZN(n7014) );
  INV_X1 U5718 ( .A(EAX_REG_2__SCAN_IN), .ZN(n6329) );
  OAI222_X1 U5719 ( .A1(n4640), .A2(n6114), .B1(n5411), .B2(n7014), .C1(n5860), 
        .C2(n6329), .ZN(U2889) );
  XNOR2_X1 U5720 ( .A(n4639), .B(n4638), .ZN(n6410) );
  OAI222_X1 U5721 ( .A1(n5836), .A2(n4640), .B1(n5349), .B2(n6292), .C1(n6288), 
        .C2(n6410), .ZN(U2857) );
  AOI21_X1 U5722 ( .B1(n4702), .B2(n4701), .A(n4642), .ZN(n4643) );
  NOR2_X1 U5723 ( .A1(n4641), .A2(n4643), .ZN(n5293) );
  INV_X1 U5724 ( .A(n5293), .ZN(n4649) );
  OR2_X1 U5725 ( .A1(n4645), .A2(n4644), .ZN(n4646) );
  NAND2_X1 U5726 ( .A1(n4646), .A2(n4760), .ZN(n6394) );
  INV_X1 U5727 ( .A(n6394), .ZN(n4647) );
  AOI22_X1 U5728 ( .A1(n5846), .A2(n4647), .B1(n4405), .B2(EBX_REG_4__SCAN_IN), 
        .ZN(n4648) );
  OAI21_X1 U5729 ( .B1(n4649), .B2(n5836), .A(n4648), .ZN(U2855) );
  INV_X1 U5730 ( .A(DATAI_4_), .ZN(n7005) );
  INV_X1 U5731 ( .A(EAX_REG_4__SCAN_IN), .ZN(n6325) );
  OAI222_X1 U5732 ( .A1(n4649), .A2(n6114), .B1(n5411), .B2(n7005), .C1(n5860), 
        .C2(n6325), .ZN(U2887) );
  OR2_X1 U5733 ( .A1(n6025), .A2(n4998), .ZN(n4734) );
  INV_X1 U5734 ( .A(n4660), .ZN(n4653) );
  NAND2_X1 U5735 ( .A1(n6484), .A2(n7056), .ZN(n6033) );
  OAI21_X1 U5736 ( .B1(n4653), .B2(n5930), .A(n6033), .ZN(n4657) );
  INV_X1 U5737 ( .A(n3463), .ZN(n6487) );
  AND2_X1 U5738 ( .A1(n5414), .A2(n6487), .ZN(n4855) );
  NOR2_X1 U5739 ( .A1(n4527), .A2(n6023), .ZN(n6448) );
  INV_X1 U5740 ( .A(n4654), .ZN(n4687) );
  AOI21_X1 U5741 ( .B1(n4855), .B2(n6448), .A(n4687), .ZN(n4659) );
  OAI21_X1 U5742 ( .B1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n6666), .A(n4820), 
        .ZN(n6496) );
  OAI21_X1 U5743 ( .B1(n6484), .B2(n4655), .A(n6455), .ZN(n4656) );
  AOI21_X1 U5744 ( .B1(n4657), .B2(n4659), .A(n4656), .ZN(n4692) );
  INV_X1 U5745 ( .A(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4663) );
  NOR2_X2 U5746 ( .A1(n4660), .A2(n5237), .ZN(n4846) );
  NAND2_X1 U5747 ( .A1(n6357), .A2(DATAI_16_), .ZN(n6494) );
  INV_X1 U5748 ( .A(n6494), .ZN(n6452) );
  NAND2_X1 U5749 ( .A1(n4686), .A2(n4986), .ZN(n6493) );
  AOI22_X1 U5750 ( .A1(n4846), .A2(n6452), .B1(n4687), .B2(n6451), .ZN(n4662)
         );
  NOR2_X1 U5751 ( .A1(n6945), .A2(n4926), .ZN(n5115) );
  OAI22_X1 U5752 ( .A1(n4659), .A2(n6498), .B1(n5042), .B2(n6590), .ZN(n4688)
         );
  NOR2_X2 U5753 ( .A1(n4660), .A2(n5138), .ZN(n5082) );
  AND2_X1 U5754 ( .A1(n6357), .A2(DATAI_24_), .ZN(n6502) );
  AOI22_X1 U5755 ( .A1(n5115), .A2(n4688), .B1(n5082), .B2(n6502), .ZN(n4661)
         );
  OAI211_X1 U5756 ( .C1(n4692), .C2(n4663), .A(n4662), .B(n4661), .ZN(U3140)
         );
  INV_X1 U5757 ( .A(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4667) );
  NAND2_X1 U5758 ( .A1(n6357), .A2(DATAI_17_), .ZN(n5435) );
  INV_X1 U5759 ( .A(n5435), .ZN(n6508) );
  NAND2_X1 U5760 ( .A1(n4686), .A2(n4664), .ZN(n5257) );
  AOI22_X1 U5761 ( .A1(n4846), .A2(n6508), .B1(n4687), .B2(n6506), .ZN(n4666)
         );
  NOR2_X1 U5762 ( .A1(n6995), .A2(n4926), .ZN(n5101) );
  AND2_X1 U5763 ( .A1(n6357), .A2(DATAI_25_), .ZN(n6507) );
  AOI22_X1 U5764 ( .A1(n5101), .A2(n4688), .B1(n5082), .B2(n6507), .ZN(n4665)
         );
  OAI211_X1 U5765 ( .C1(n4692), .C2(n4667), .A(n4666), .B(n4665), .ZN(U3141)
         );
  INV_X1 U5766 ( .A(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4671) );
  NAND2_X1 U5767 ( .A1(n6357), .A2(DATAI_18_), .ZN(n6513) );
  INV_X1 U5768 ( .A(n6513), .ZN(n6464) );
  NAND2_X1 U5769 ( .A1(n4686), .A2(n4668), .ZN(n6512) );
  AOI22_X1 U5770 ( .A1(n4846), .A2(n6464), .B1(n4687), .B2(n6463), .ZN(n4670)
         );
  AND2_X1 U5771 ( .A1(n6357), .A2(DATAI_26_), .ZN(n6515) );
  AOI22_X1 U5772 ( .A1(n6462), .A2(n4688), .B1(n5082), .B2(n6515), .ZN(n4669)
         );
  OAI211_X1 U5773 ( .C1(n4692), .C2(n4671), .A(n4670), .B(n4669), .ZN(U3142)
         );
  INV_X1 U5774 ( .A(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4675) );
  NAND2_X1 U5775 ( .A1(n6357), .A2(DATAI_20_), .ZN(n6526) );
  INV_X1 U5776 ( .A(n6526), .ZN(n6470) );
  NAND2_X1 U5777 ( .A1(n4686), .A2(n4672), .ZN(n6525) );
  AOI22_X1 U5778 ( .A1(n4846), .A2(n6470), .B1(n4687), .B2(n6469), .ZN(n4674)
         );
  NOR2_X1 U5779 ( .A1(n7005), .A2(n4926), .ZN(n5119) );
  AND2_X1 U5780 ( .A1(n6357), .A2(DATAI_28_), .ZN(n6529) );
  AOI22_X1 U5781 ( .A1(n5119), .A2(n4688), .B1(n5082), .B2(n6529), .ZN(n4673)
         );
  OAI211_X1 U5782 ( .C1(n4692), .C2(n4675), .A(n4674), .B(n4673), .ZN(U3144)
         );
  INV_X1 U5783 ( .A(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4679) );
  NAND2_X1 U5784 ( .A1(n6357), .A2(DATAI_19_), .ZN(n5427) );
  INV_X1 U5785 ( .A(n5427), .ZN(n6520) );
  NAND2_X1 U5786 ( .A1(n4686), .A2(n4676), .ZN(n5249) );
  AOI22_X1 U5787 ( .A1(n4846), .A2(n6520), .B1(n4687), .B2(n6518), .ZN(n4678)
         );
  INV_X1 U5788 ( .A(DATAI_3_), .ZN(n6986) );
  NOR2_X1 U5789 ( .A1(n6986), .A2(n4926), .ZN(n6431) );
  AND2_X1 U5790 ( .A1(n6357), .A2(DATAI_27_), .ZN(n6519) );
  AOI22_X1 U5791 ( .A1(n6431), .A2(n4688), .B1(n5082), .B2(n6519), .ZN(n4677)
         );
  OAI211_X1 U5792 ( .C1(n4692), .C2(n4679), .A(n4678), .B(n4677), .ZN(U3143)
         );
  INV_X1 U5793 ( .A(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4682) );
  NAND2_X1 U5794 ( .A1(n6357), .A2(DATAI_23_), .ZN(n5443) );
  INV_X1 U5795 ( .A(n5443), .ZN(n6550) );
  NAND2_X1 U5796 ( .A1(n4686), .A2(n3324), .ZN(n5267) );
  AOI22_X1 U5797 ( .A1(n4846), .A2(n6550), .B1(n4687), .B2(n6546), .ZN(n4681)
         );
  INV_X1 U5798 ( .A(DATAI_7_), .ZN(n5040) );
  NOR2_X1 U5799 ( .A1(n5040), .A2(n4926), .ZN(n5129) );
  AND2_X1 U5800 ( .A1(n6357), .A2(DATAI_31_), .ZN(n6547) );
  AOI22_X1 U5801 ( .A1(n5129), .A2(n4688), .B1(n5082), .B2(n6547), .ZN(n4680)
         );
  OAI211_X1 U5802 ( .C1(n4692), .C2(n4682), .A(n4681), .B(n4680), .ZN(U3147)
         );
  INV_X1 U5803 ( .A(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4685) );
  NAND2_X1 U5804 ( .A1(n6357), .A2(DATAI_22_), .ZN(n5439) );
  INV_X1 U5805 ( .A(n5439), .ZN(n6541) );
  NAND2_X1 U5806 ( .A1(n4686), .A2(n3318), .ZN(n5275) );
  AOI22_X1 U5807 ( .A1(n4846), .A2(n6541), .B1(n4687), .B2(n6539), .ZN(n4684)
         );
  INV_X1 U5808 ( .A(DATAI_6_), .ZN(n4815) );
  NOR2_X1 U5809 ( .A1(n4815), .A2(n4926), .ZN(n5108) );
  AND2_X1 U5810 ( .A1(n6357), .A2(DATAI_30_), .ZN(n6540) );
  AOI22_X1 U5811 ( .A1(n5108), .A2(n4688), .B1(n5082), .B2(n6540), .ZN(n4683)
         );
  OAI211_X1 U5812 ( .C1(n4692), .C2(n4685), .A(n4684), .B(n4683), .ZN(U3146)
         );
  INV_X1 U5813 ( .A(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4691) );
  NAND2_X1 U5814 ( .A1(n6357), .A2(DATAI_21_), .ZN(n5431) );
  INV_X1 U5815 ( .A(n5431), .ZN(n6535) );
  NAND2_X1 U5816 ( .A1(n4686), .A2(n5492), .ZN(n5253) );
  AOI22_X1 U5817 ( .A1(n4846), .A2(n6535), .B1(n4687), .B2(n6533), .ZN(n4690)
         );
  INV_X1 U5818 ( .A(DATAI_5_), .ZN(n6881) );
  NOR2_X1 U5819 ( .A1(n6881), .A2(n4926), .ZN(n6438) );
  NAND2_X1 U5820 ( .A1(n6357), .A2(DATAI_29_), .ZN(n6442) );
  INV_X1 U5821 ( .A(n6442), .ZN(n6534) );
  AOI22_X1 U5822 ( .A1(n6438), .A2(n4688), .B1(n5082), .B2(n6534), .ZN(n4689)
         );
  OAI211_X1 U5823 ( .C1(n4692), .C2(n4691), .A(n4690), .B(n4689), .ZN(U3145)
         );
  OR2_X1 U5824 ( .A1(n4695), .A2(n4694), .ZN(n4696) );
  NAND2_X1 U5825 ( .A1(n4693), .A2(n4696), .ZN(n6399) );
  INV_X1 U5826 ( .A(n5285), .ZN(n4698) );
  INV_X1 U5827 ( .A(n6393), .ZN(n6411) );
  AOI22_X1 U5828 ( .A1(n6361), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .B1(n6411), 
        .B2(REIP_REG_4__SCAN_IN), .ZN(n4697) );
  OAI21_X1 U5829 ( .B1(n4698), .B2(n6370), .A(n4697), .ZN(n4699) );
  AOI21_X1 U5830 ( .B1(n5293), .B2(n6357), .A(n4699), .ZN(n4700) );
  OAI21_X1 U5831 ( .B1(n6399), .B2(n6195), .A(n4700), .ZN(U2982) );
  XOR2_X1 U5832 ( .A(n4702), .B(n4701), .Z(n6356) );
  INV_X1 U5833 ( .A(n6356), .ZN(n4706) );
  AOI21_X1 U5834 ( .B1(n4704), .B2(n4703), .A(n4644), .ZN(n6405) );
  AOI22_X1 U5835 ( .A1(n5846), .A2(n6405), .B1(EBX_REG_3__SCAN_IN), .B2(n4405), 
        .ZN(n4705) );
  OAI21_X1 U5836 ( .B1(n4706), .B2(n5836), .A(n4705), .ZN(U2856) );
  INV_X1 U5837 ( .A(EAX_REG_3__SCAN_IN), .ZN(n6327) );
  OAI222_X1 U5838 ( .A1(n4706), .A2(n6114), .B1(n5411), .B2(n6986), .C1(n5860), 
        .C2(n6327), .ZN(U2888) );
  INV_X1 U5839 ( .A(n6519), .ZN(n6434) );
  NAND2_X1 U5840 ( .A1(n6025), .A2(n5089), .ZN(n4707) );
  NAND2_X1 U5841 ( .A1(n4713), .A2(n5237), .ZN(n4817) );
  AND2_X1 U5842 ( .A1(n6023), .A2(n4527), .ZN(n5000) );
  NAND2_X1 U5843 ( .A1(n6281), .A2(n5000), .ZN(n4825) );
  INV_X1 U5844 ( .A(n4825), .ZN(n4708) );
  NAND3_X1 U5845 ( .A1(n6573), .A2(n5243), .A3(n4854), .ZN(n4819) );
  NOR2_X1 U5846 ( .A1(n6558), .A2(n4819), .ZN(n4730) );
  AOI21_X1 U5847 ( .B1(n4708), .B2(n6487), .A(n4730), .ZN(n4712) );
  AOI21_X1 U5848 ( .B1(n4713), .B2(STATEBS16_REG_SCAN_IN), .A(n6498), .ZN(
        n4710) );
  AOI22_X1 U5849 ( .A1(n4712), .A2(n4710), .B1(n6498), .B2(n4819), .ZN(n4709)
         );
  NAND2_X1 U5850 ( .A1(n6455), .A2(n4709), .ZN(n4729) );
  INV_X1 U5851 ( .A(n4710), .ZN(n4711) );
  OAI22_X1 U5852 ( .A1(n4712), .A2(n4711), .B1(n6590), .B2(n4819), .ZN(n4728)
         );
  AOI22_X1 U5853 ( .A1(INSTQUEUE_REG_1__3__SCAN_IN), .A2(n4729), .B1(n6431), 
        .B2(n4728), .ZN(n4715) );
  AOI22_X1 U5854 ( .A1(n4793), .A2(n6520), .B1(n6518), .B2(n4730), .ZN(n4714)
         );
  OAI211_X1 U5855 ( .C1(n6434), .C2(n4817), .A(n4715), .B(n4714), .ZN(U3031)
         );
  INV_X1 U5856 ( .A(n6515), .ZN(n6430) );
  AOI22_X1 U5857 ( .A1(INSTQUEUE_REG_1__2__SCAN_IN), .A2(n4729), .B1(n6462), 
        .B2(n4728), .ZN(n4717) );
  AOI22_X1 U5858 ( .A1(n4793), .A2(n6464), .B1(n6463), .B2(n4730), .ZN(n4716)
         );
  OAI211_X1 U5859 ( .C1(n6430), .C2(n4817), .A(n4717), .B(n4716), .ZN(U3030)
         );
  INV_X1 U5860 ( .A(n6507), .ZN(n5156) );
  AOI22_X1 U5861 ( .A1(INSTQUEUE_REG_1__1__SCAN_IN), .A2(n4729), .B1(n5101), 
        .B2(n4728), .ZN(n4719) );
  AOI22_X1 U5862 ( .A1(n4793), .A2(n6508), .B1(n6506), .B2(n4730), .ZN(n4718)
         );
  OAI211_X1 U5863 ( .C1(n5156), .C2(n4817), .A(n4719), .B(n4718), .ZN(U3029)
         );
  INV_X1 U5864 ( .A(n6502), .ZN(n5146) );
  AOI22_X1 U5865 ( .A1(INSTQUEUE_REG_1__0__SCAN_IN), .A2(n4729), .B1(n5115), 
        .B2(n4728), .ZN(n4721) );
  AOI22_X1 U5866 ( .A1(n4793), .A2(n6452), .B1(n6451), .B2(n4730), .ZN(n4720)
         );
  OAI211_X1 U5867 ( .C1(n5146), .C2(n4817), .A(n4721), .B(n4720), .ZN(U3028)
         );
  AOI22_X1 U5868 ( .A1(INSTQUEUE_REG_1__5__SCAN_IN), .A2(n4729), .B1(n6438), 
        .B2(n4728), .ZN(n4723) );
  AOI22_X1 U5869 ( .A1(n4793), .A2(n6535), .B1(n6533), .B2(n4730), .ZN(n4722)
         );
  OAI211_X1 U5870 ( .C1(n6442), .C2(n4817), .A(n4723), .B(n4722), .ZN(U3033)
         );
  INV_X1 U5871 ( .A(n6529), .ZN(n5164) );
  AOI22_X1 U5872 ( .A1(INSTQUEUE_REG_1__4__SCAN_IN), .A2(n4729), .B1(n5119), 
        .B2(n4728), .ZN(n4725) );
  AOI22_X1 U5873 ( .A1(n4793), .A2(n6470), .B1(n6469), .B2(n4730), .ZN(n4724)
         );
  OAI211_X1 U5874 ( .C1(n5164), .C2(n4817), .A(n4725), .B(n4724), .ZN(U3032)
         );
  INV_X1 U5875 ( .A(n6547), .ZN(n5160) );
  AOI22_X1 U5876 ( .A1(INSTQUEUE_REG_1__7__SCAN_IN), .A2(n4729), .B1(n5129), 
        .B2(n4728), .ZN(n4727) );
  AOI22_X1 U5877 ( .A1(n4793), .A2(n6550), .B1(n6546), .B2(n4730), .ZN(n4726)
         );
  OAI211_X1 U5878 ( .C1(n5160), .C2(n4817), .A(n4727), .B(n4726), .ZN(U3035)
         );
  INV_X1 U5879 ( .A(n6540), .ZN(n5168) );
  AOI22_X1 U5880 ( .A1(INSTQUEUE_REG_1__6__SCAN_IN), .A2(n4729), .B1(n5108), 
        .B2(n4728), .ZN(n4732) );
  AOI22_X1 U5881 ( .A1(n4793), .A2(n6541), .B1(n6539), .B2(n4730), .ZN(n4731)
         );
  OAI211_X1 U5882 ( .C1(n5168), .C2(n4817), .A(n4732), .B(n4731), .ZN(U3034)
         );
  XOR2_X1 U5883 ( .A(n4641), .B(n4733), .Z(n6347) );
  INV_X1 U5884 ( .A(n6347), .ZN(n4762) );
  INV_X1 U5885 ( .A(EAX_REG_5__SCAN_IN), .ZN(n6322) );
  OAI222_X1 U5886 ( .A1(n6114), .A2(n4762), .B1(n5411), .B2(n6881), .C1(n5860), 
        .C2(n6322), .ZN(U2886) );
  NAND2_X1 U5887 ( .A1(n4736), .A2(n5138), .ZN(n5080) );
  NOR2_X1 U5888 ( .A1(n4527), .A2(n4982), .ZN(n5092) );
  NAND2_X1 U5889 ( .A1(n4854), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n5088) );
  NOR2_X1 U5890 ( .A1(n6573), .A2(n5088), .ZN(n4923) );
  AND2_X1 U5891 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4923), .ZN(n4757)
         );
  AOI21_X1 U5892 ( .B1(n4855), .B2(n5092), .A(n4757), .ZN(n4737) );
  NAND2_X1 U5893 ( .A1(STATE2_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4735) );
  OAI22_X1 U5894 ( .A1(n4737), .A2(n6498), .B1(n4735), .B2(n5088), .ZN(n4755)
         );
  AOI22_X1 U5895 ( .A1(n5063), .A2(n6508), .B1(n5101), .B2(n4755), .ZN(n4742)
         );
  NAND2_X1 U5896 ( .A1(n4736), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4871) );
  NAND2_X1 U5897 ( .A1(n4737), .A2(n4871), .ZN(n4740) );
  INV_X1 U5898 ( .A(n4923), .ZN(n4738) );
  NAND2_X1 U5899 ( .A1(n6498), .A2(n4738), .ZN(n4739) );
  OAI211_X1 U5900 ( .C1(n6498), .C2(n4740), .A(n6455), .B(n4739), .ZN(n4756)
         );
  AOI22_X1 U5901 ( .A1(n6506), .A2(n4757), .B1(INSTQUEUE_REG_13__1__SCAN_IN), 
        .B2(n4756), .ZN(n4741) );
  OAI211_X1 U5902 ( .C1(n5156), .C2(n4959), .A(n4742), .B(n4741), .ZN(U3125)
         );
  AOI22_X1 U5903 ( .A1(n5063), .A2(n6520), .B1(n6431), .B2(n4755), .ZN(n4744)
         );
  AOI22_X1 U5904 ( .A1(n6518), .A2(n4757), .B1(INSTQUEUE_REG_13__3__SCAN_IN), 
        .B2(n4756), .ZN(n4743) );
  OAI211_X1 U5905 ( .C1(n6434), .C2(n4959), .A(n4744), .B(n4743), .ZN(U3127)
         );
  AOI22_X1 U5906 ( .A1(n5063), .A2(n6550), .B1(n5129), .B2(n4755), .ZN(n4746)
         );
  AOI22_X1 U5907 ( .A1(n6546), .A2(n4757), .B1(INSTQUEUE_REG_13__7__SCAN_IN), 
        .B2(n4756), .ZN(n4745) );
  OAI211_X1 U5908 ( .C1(n5160), .C2(n4959), .A(n4746), .B(n4745), .ZN(U3131)
         );
  AOI22_X1 U5909 ( .A1(n5063), .A2(n6535), .B1(n6438), .B2(n4755), .ZN(n4748)
         );
  AOI22_X1 U5910 ( .A1(n6533), .A2(n4757), .B1(INSTQUEUE_REG_13__5__SCAN_IN), 
        .B2(n4756), .ZN(n4747) );
  OAI211_X1 U5911 ( .C1(n6442), .C2(n4959), .A(n4748), .B(n4747), .ZN(U3129)
         );
  AOI22_X1 U5912 ( .A1(n5063), .A2(n6452), .B1(n5115), .B2(n4755), .ZN(n4750)
         );
  AOI22_X1 U5913 ( .A1(n6451), .A2(n4757), .B1(INSTQUEUE_REG_13__0__SCAN_IN), 
        .B2(n4756), .ZN(n4749) );
  OAI211_X1 U5914 ( .C1(n5146), .C2(n4959), .A(n4750), .B(n4749), .ZN(U3124)
         );
  AOI22_X1 U5915 ( .A1(n5063), .A2(n6470), .B1(n5119), .B2(n4755), .ZN(n4752)
         );
  AOI22_X1 U5916 ( .A1(n6469), .A2(n4757), .B1(INSTQUEUE_REG_13__4__SCAN_IN), 
        .B2(n4756), .ZN(n4751) );
  OAI211_X1 U5917 ( .C1(n5164), .C2(n4959), .A(n4752), .B(n4751), .ZN(U3128)
         );
  AOI22_X1 U5918 ( .A1(n5063), .A2(n6464), .B1(n6462), .B2(n4755), .ZN(n4754)
         );
  AOI22_X1 U5919 ( .A1(n6463), .A2(n4757), .B1(INSTQUEUE_REG_13__2__SCAN_IN), 
        .B2(n4756), .ZN(n4753) );
  OAI211_X1 U5920 ( .C1(n6430), .C2(n4959), .A(n4754), .B(n4753), .ZN(U3126)
         );
  AOI22_X1 U5921 ( .A1(n5063), .A2(n6541), .B1(n5108), .B2(n4755), .ZN(n4759)
         );
  AOI22_X1 U5922 ( .A1(n6539), .A2(n4757), .B1(INSTQUEUE_REG_13__6__SCAN_IN), 
        .B2(n4756), .ZN(n4758) );
  OAI211_X1 U5923 ( .C1(n5168), .C2(n4959), .A(n4759), .B(n4758), .ZN(U3130)
         );
  AOI21_X1 U5924 ( .B1(n4761), .B2(n4760), .A(n4803), .ZN(n6262) );
  INV_X1 U5925 ( .A(n6262), .ZN(n4764) );
  OAI222_X1 U5926 ( .A1(n4764), .A2(n6288), .B1(n4763), .B2(n6292), .C1(n5854), 
        .C2(n4762), .ZN(U2854) );
  NAND3_X1 U5927 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n6573), .A3(n5243), .ZN(n4877) );
  NOR2_X1 U5928 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4877), .ZN(n4791)
         );
  AND2_X1 U5929 ( .A1(n6025), .A2(n4652), .ZN(n4765) );
  NAND2_X1 U5930 ( .A1(n4246), .A2(n4765), .ZN(n4881) );
  OAI21_X1 U5931 ( .B1(n4794), .B2(n4793), .A(n6033), .ZN(n4766) );
  AND2_X1 U5932 ( .A1(n4527), .A2(n4982), .ZN(n5240) );
  NAND2_X1 U5933 ( .A1(n6281), .A2(n5240), .ZN(n4873) );
  NAND2_X1 U5934 ( .A1(n4766), .A2(n4873), .ZN(n4767) );
  NOR2_X1 U5935 ( .A1(n4769), .A2(n6590), .ZN(n5417) );
  OAI21_X1 U5936 ( .B1(n4924), .B2(n6590), .A(n4820), .ZN(n5043) );
  NOR2_X1 U5937 ( .A1(n5417), .A2(n5043), .ZN(n5247) );
  OAI221_X1 U5938 ( .B1(n4791), .B2(n6666), .C1(n4791), .C2(n4767), .A(n5247), 
        .ZN(n4768) );
  INV_X1 U5939 ( .A(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4772) );
  AND2_X1 U5940 ( .A1(n4769), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5242) );
  INV_X1 U5941 ( .A(n5242), .ZN(n4927) );
  NAND2_X1 U5942 ( .A1(n4924), .A2(n6573), .ZN(n5413) );
  OAI22_X1 U5943 ( .A1(n4873), .A2(n6498), .B1(n4927), .B2(n5413), .ZN(n4792)
         );
  AOI22_X1 U5944 ( .A1(n6462), .A2(n4792), .B1(n6463), .B2(n4791), .ZN(n4771)
         );
  AOI22_X1 U5945 ( .A1(n4794), .A2(n6464), .B1(n4793), .B2(n6515), .ZN(n4770)
         );
  OAI211_X1 U5946 ( .C1(n4798), .C2(n4772), .A(n4771), .B(n4770), .ZN(U3038)
         );
  INV_X1 U5947 ( .A(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4775) );
  AOI22_X1 U5948 ( .A1(n5108), .A2(n4792), .B1(n6539), .B2(n4791), .ZN(n4774)
         );
  AOI22_X1 U5949 ( .A1(n4794), .A2(n6541), .B1(n4793), .B2(n6540), .ZN(n4773)
         );
  OAI211_X1 U5950 ( .C1(n4798), .C2(n4775), .A(n4774), .B(n4773), .ZN(U3042)
         );
  INV_X1 U5951 ( .A(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4778) );
  AOI22_X1 U5952 ( .A1(n6438), .A2(n4792), .B1(n6533), .B2(n4791), .ZN(n4777)
         );
  AOI22_X1 U5953 ( .A1(n4794), .A2(n6535), .B1(n4793), .B2(n6534), .ZN(n4776)
         );
  OAI211_X1 U5954 ( .C1(n4798), .C2(n4778), .A(n4777), .B(n4776), .ZN(U3041)
         );
  INV_X1 U5955 ( .A(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4781) );
  AOI22_X1 U5956 ( .A1(n5119), .A2(n4792), .B1(n6469), .B2(n4791), .ZN(n4780)
         );
  AOI22_X1 U5957 ( .A1(n4794), .A2(n6470), .B1(n4793), .B2(n6529), .ZN(n4779)
         );
  OAI211_X1 U5958 ( .C1(n4798), .C2(n4781), .A(n4780), .B(n4779), .ZN(U3040)
         );
  INV_X1 U5959 ( .A(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4784) );
  AOI22_X1 U5960 ( .A1(n6431), .A2(n4792), .B1(n6518), .B2(n4791), .ZN(n4783)
         );
  AOI22_X1 U5961 ( .A1(n4794), .A2(n6520), .B1(n4793), .B2(n6519), .ZN(n4782)
         );
  OAI211_X1 U5962 ( .C1(n4798), .C2(n4784), .A(n4783), .B(n4782), .ZN(U3039)
         );
  INV_X1 U5963 ( .A(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4787) );
  AOI22_X1 U5964 ( .A1(n5115), .A2(n4792), .B1(n6451), .B2(n4791), .ZN(n4786)
         );
  AOI22_X1 U5965 ( .A1(n4794), .A2(n6452), .B1(n4793), .B2(n6502), .ZN(n4785)
         );
  OAI211_X1 U5966 ( .C1(n4798), .C2(n4787), .A(n4786), .B(n4785), .ZN(U3036)
         );
  INV_X1 U5967 ( .A(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4790) );
  AOI22_X1 U5968 ( .A1(n5101), .A2(n4792), .B1(n6506), .B2(n4791), .ZN(n4789)
         );
  AOI22_X1 U5969 ( .A1(n4794), .A2(n6508), .B1(n4793), .B2(n6507), .ZN(n4788)
         );
  OAI211_X1 U5970 ( .C1(n4798), .C2(n4790), .A(n4789), .B(n4788), .ZN(U3037)
         );
  INV_X1 U5971 ( .A(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4797) );
  AOI22_X1 U5972 ( .A1(n5129), .A2(n4792), .B1(n6546), .B2(n4791), .ZN(n4796)
         );
  AOI22_X1 U5973 ( .A1(n4794), .A2(n6550), .B1(n4793), .B2(n6547), .ZN(n4795)
         );
  OAI211_X1 U5974 ( .C1(n4798), .C2(n4797), .A(n4796), .B(n4795), .ZN(U3043)
         );
  CLKBUF_X1 U5975 ( .A(n4800), .Z(n4801) );
  OAI21_X1 U5976 ( .B1(n4799), .B2(n4802), .A(n4801), .ZN(n4921) );
  OAI21_X1 U5977 ( .B1(n4804), .B2(n4803), .A(n5208), .ZN(n5322) );
  INV_X1 U5978 ( .A(n5322), .ZN(n4811) );
  AND2_X1 U5979 ( .A1(n6411), .A2(REIP_REG_6__SCAN_IN), .ZN(n4918) );
  NAND2_X1 U5981 ( .A1(n6392), .A2(n4805), .ZN(n5686) );
  INV_X1 U5982 ( .A(n5199), .ZN(n4806) );
  OAI21_X1 U5983 ( .B1(n4806), .B2(n6415), .A(n5195), .ZN(n6417) );
  AOI221_X1 U5984 ( .B1(n5688), .B2(n5633), .C1(n5686), .C2(n5633), .A(n6417), 
        .ZN(n5685) );
  AOI21_X1 U5985 ( .B1(n6415), .B2(n6420), .A(n6414), .ZN(n5193) );
  OR2_X1 U5986 ( .A1(n6416), .A2(n5193), .ZN(n6409) );
  OAI33_X1 U5987 ( .A1(1'b0), .A2(n5685), .A3(n4808), .B1(
        INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n4807), .B3(n6409), .ZN(n4810) );
  AOI211_X1 U5988 ( .C1(n6412), .C2(n4811), .A(n4918), .B(n4810), .ZN(n4812)
         );
  OAI21_X1 U5989 ( .B1(n6398), .B2(n4921), .A(n4812), .ZN(U3012) );
  OAI21_X1 U5990 ( .B1(n4813), .B2(n4814), .A(n4971), .ZN(n5326) );
  INV_X1 U5991 ( .A(EAX_REG_6__SCAN_IN), .ZN(n6320) );
  OAI222_X1 U5992 ( .A1(n5326), .A2(n6114), .B1(n5411), .B2(n4815), .C1(n5860), 
        .C2(n6320), .ZN(U2885) );
  INV_X1 U5993 ( .A(EBX_REG_6__SCAN_IN), .ZN(n4816) );
  OAI222_X1 U5994 ( .A1(n5326), .A2(n5836), .B1(n6292), .B2(n4816), .C1(n5322), 
        .C2(n6288), .ZN(U2853) );
  NOR3_X1 U5995 ( .A1(n4848), .A2(n4846), .A3(n6498), .ZN(n4818) );
  INV_X1 U5996 ( .A(n6033), .ZN(n5134) );
  OAI21_X1 U5997 ( .B1(n4818), .B2(n5134), .A(n4825), .ZN(n4823) );
  NOR2_X1 U5998 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4819), .ZN(n4845)
         );
  INV_X1 U5999 ( .A(n4845), .ZN(n4821) );
  NOR2_X1 U6000 ( .A1(n4924), .A2(n4925), .ZN(n4824) );
  OAI21_X1 U6001 ( .B1(n4824), .B2(n6590), .A(n4820), .ZN(n5094) );
  AOI211_X1 U6002 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n4821), .A(n5417), .B(
        n5094), .ZN(n4822) );
  INV_X1 U6003 ( .A(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4828) );
  AOI22_X1 U6004 ( .A1(n4846), .A2(n6534), .B1(n6533), .B2(n4845), .ZN(n4827)
         );
  INV_X1 U6005 ( .A(n4824), .ZN(n5098) );
  OAI22_X1 U6006 ( .A1(n4825), .A2(n6498), .B1(n4927), .B2(n5098), .ZN(n4847)
         );
  AOI22_X1 U6007 ( .A1(n4848), .A2(n6535), .B1(n6438), .B2(n4847), .ZN(n4826)
         );
  OAI211_X1 U6008 ( .C1(n4852), .C2(n4828), .A(n4827), .B(n4826), .ZN(U3025)
         );
  INV_X1 U6009 ( .A(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4831) );
  AOI22_X1 U6010 ( .A1(n4846), .A2(n6547), .B1(n6546), .B2(n4845), .ZN(n4830)
         );
  AOI22_X1 U6011 ( .A1(n4848), .A2(n6550), .B1(n5129), .B2(n4847), .ZN(n4829)
         );
  OAI211_X1 U6012 ( .C1(n4852), .C2(n4831), .A(n4830), .B(n4829), .ZN(U3027)
         );
  AOI22_X1 U6013 ( .A1(n4846), .A2(n6529), .B1(n6469), .B2(n4845), .ZN(n4833)
         );
  AOI22_X1 U6014 ( .A1(n4848), .A2(n6470), .B1(n5119), .B2(n4847), .ZN(n4832)
         );
  OAI211_X1 U6015 ( .C1(n4852), .C2(n3513), .A(n4833), .B(n4832), .ZN(U3024)
         );
  INV_X1 U6016 ( .A(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4836) );
  AOI22_X1 U6017 ( .A1(n4846), .A2(n6502), .B1(n6451), .B2(n4845), .ZN(n4835)
         );
  AOI22_X1 U6018 ( .A1(n4848), .A2(n6452), .B1(n5115), .B2(n4847), .ZN(n4834)
         );
  OAI211_X1 U6019 ( .C1(n4852), .C2(n4836), .A(n4835), .B(n4834), .ZN(U3020)
         );
  AOI22_X1 U6020 ( .A1(n4846), .A2(n6540), .B1(n6539), .B2(n4845), .ZN(n4838)
         );
  AOI22_X1 U6021 ( .A1(n4848), .A2(n6541), .B1(n5108), .B2(n4847), .ZN(n4837)
         );
  OAI211_X1 U6022 ( .C1(n4852), .C2(n3558), .A(n4838), .B(n4837), .ZN(U3026)
         );
  INV_X1 U6023 ( .A(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4841) );
  AOI22_X1 U6024 ( .A1(n4846), .A2(n6519), .B1(n6518), .B2(n4845), .ZN(n4840)
         );
  AOI22_X1 U6025 ( .A1(n4848), .A2(n6520), .B1(n6431), .B2(n4847), .ZN(n4839)
         );
  OAI211_X1 U6026 ( .C1(n4852), .C2(n4841), .A(n4840), .B(n4839), .ZN(U3023)
         );
  INV_X1 U6027 ( .A(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4844) );
  AOI22_X1 U6028 ( .A1(n4846), .A2(n6515), .B1(n6463), .B2(n4845), .ZN(n4843)
         );
  AOI22_X1 U6029 ( .A1(n4848), .A2(n6464), .B1(n6462), .B2(n4847), .ZN(n4842)
         );
  OAI211_X1 U6030 ( .C1(n4852), .C2(n4844), .A(n4843), .B(n4842), .ZN(U3022)
         );
  INV_X1 U6031 ( .A(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4851) );
  AOI22_X1 U6032 ( .A1(n4846), .A2(n6507), .B1(n6506), .B2(n4845), .ZN(n4850)
         );
  AOI22_X1 U6033 ( .A1(n4848), .A2(n6508), .B1(n5101), .B2(n4847), .ZN(n4849)
         );
  OAI211_X1 U6034 ( .C1(n4852), .C2(n4851), .A(n4850), .B(n4849), .ZN(U3021)
         );
  AOI21_X1 U6035 ( .B1(n4860), .B2(STATEBS16_REG_SCAN_IN), .A(n6498), .ZN(
        n4857) );
  NAND3_X1 U6036 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n5243), .A3(n4854), .ZN(n5002) );
  NOR2_X1 U6037 ( .A1(n6558), .A2(n5002), .ZN(n4861) );
  AOI21_X1 U6038 ( .B1(n4855), .B2(n5000), .A(n4861), .ZN(n4859) );
  AOI22_X1 U6039 ( .A1(n4857), .A2(n4859), .B1(n6498), .B2(n5002), .ZN(n4856)
         );
  NAND2_X1 U6040 ( .A1(n6455), .A2(n4856), .ZN(n4911) );
  INV_X1 U6041 ( .A(n4857), .ZN(n4858) );
  OAI22_X1 U6042 ( .A1(n4859), .A2(n4858), .B1(n6590), .B2(n5002), .ZN(n4910)
         );
  AOI22_X1 U6043 ( .A1(INSTQUEUE_REG_9__2__SCAN_IN), .A2(n4911), .B1(n6462), 
        .B2(n4910), .ZN(n4864) );
  INV_X1 U6044 ( .A(n4861), .ZN(n4912) );
  OAI22_X1 U6045 ( .A1(n5248), .A2(n6513), .B1(n6512), .B2(n4912), .ZN(n4862)
         );
  AOI21_X1 U6046 ( .B1(n6515), .B2(n4997), .A(n4862), .ZN(n4863) );
  NAND2_X1 U6047 ( .A1(n4864), .A2(n4863), .ZN(U3094) );
  AOI22_X1 U6048 ( .A1(INSTQUEUE_REG_9__3__SCAN_IN), .A2(n4911), .B1(n6431), 
        .B2(n4910), .ZN(n4867) );
  OAI22_X1 U6049 ( .A1(n5248), .A2(n5427), .B1(n5249), .B2(n4912), .ZN(n4865)
         );
  AOI21_X1 U6050 ( .B1(n6519), .B2(n4997), .A(n4865), .ZN(n4866) );
  NAND2_X1 U6051 ( .A1(n4867), .A2(n4866), .ZN(U3095) );
  AOI22_X1 U6052 ( .A1(INSTQUEUE_REG_9__5__SCAN_IN), .A2(n4911), .B1(n6438), 
        .B2(n4910), .ZN(n4870) );
  OAI22_X1 U6053 ( .A1(n5248), .A2(n5431), .B1(n5253), .B2(n4912), .ZN(n4868)
         );
  AOI21_X1 U6054 ( .B1(n6534), .B2(n4997), .A(n4868), .ZN(n4869) );
  NAND2_X1 U6055 ( .A1(n4870), .A2(n4869), .ZN(U3097) );
  NAND2_X1 U6056 ( .A1(n4871), .A2(n6486), .ZN(n6030) );
  AND2_X1 U6057 ( .A1(n4652), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6021) );
  NAND2_X1 U6058 ( .A1(n6021), .A2(n6025), .ZN(n4872) );
  OAI21_X1 U6059 ( .B1(n6030), .B2(n4872), .A(n6484), .ZN(n4880) );
  OR2_X1 U6060 ( .A1(n4873), .A2(n3463), .ZN(n4875) );
  INV_X1 U6061 ( .A(n4874), .ZN(n6489) );
  NAND2_X1 U6062 ( .A1(n6489), .A2(n6573), .ZN(n6427) );
  NAND2_X1 U6063 ( .A1(n4875), .A2(n6427), .ZN(n4879) );
  INV_X1 U6064 ( .A(n4879), .ZN(n4876) );
  OAI22_X1 U6065 ( .A1(n4880), .A2(n4876), .B1(n4877), .B2(n6590), .ZN(n6437)
         );
  INV_X1 U6066 ( .A(n6437), .ZN(n4897) );
  INV_X1 U6067 ( .A(n5129), .ZN(n6554) );
  AOI21_X1 U6068 ( .B1(n6498), .B2(n4877), .A(n6496), .ZN(n4878) );
  OAI21_X1 U6069 ( .B1(n4880), .B2(n4879), .A(n4878), .ZN(n6439) );
  NOR2_X1 U6070 ( .A1(n6443), .A2(n5160), .ZN(n4883) );
  OAI22_X1 U6071 ( .A1(n5090), .A2(n5443), .B1(n5267), .B2(n6427), .ZN(n4882)
         );
  AOI211_X1 U6072 ( .C1(n6439), .C2(INSTQUEUE_REG_3__7__SCAN_IN), .A(n4883), 
        .B(n4882), .ZN(n4884) );
  OAI21_X1 U6073 ( .B1(n4897), .B2(n6554), .A(n4884), .ZN(U3051) );
  INV_X1 U6074 ( .A(n5119), .ZN(n6532) );
  NOR2_X1 U6075 ( .A1(n6443), .A2(n5164), .ZN(n4886) );
  OAI22_X1 U6076 ( .A1(n5090), .A2(n6526), .B1(n6525), .B2(n6427), .ZN(n4885)
         );
  AOI211_X1 U6077 ( .C1(n6439), .C2(INSTQUEUE_REG_3__4__SCAN_IN), .A(n4886), 
        .B(n4885), .ZN(n4887) );
  OAI21_X1 U6078 ( .B1(n4897), .B2(n6532), .A(n4887), .ZN(U3048) );
  INV_X1 U6079 ( .A(n5115), .ZN(n6505) );
  NOR2_X1 U6080 ( .A1(n6443), .A2(n5146), .ZN(n4889) );
  OAI22_X1 U6081 ( .A1(n5090), .A2(n6494), .B1(n6493), .B2(n6427), .ZN(n4888)
         );
  AOI211_X1 U6082 ( .C1(n6439), .C2(INSTQUEUE_REG_3__0__SCAN_IN), .A(n4889), 
        .B(n4888), .ZN(n4890) );
  OAI21_X1 U6083 ( .B1(n4897), .B2(n6505), .A(n4890), .ZN(U3044) );
  INV_X1 U6084 ( .A(n5108), .ZN(n6544) );
  NOR2_X1 U6085 ( .A1(n6443), .A2(n5168), .ZN(n4892) );
  OAI22_X1 U6086 ( .A1(n5090), .A2(n5439), .B1(n5275), .B2(n6427), .ZN(n4891)
         );
  AOI211_X1 U6087 ( .C1(n6439), .C2(INSTQUEUE_REG_3__6__SCAN_IN), .A(n4892), 
        .B(n4891), .ZN(n4893) );
  OAI21_X1 U6088 ( .B1(n4897), .B2(n6544), .A(n4893), .ZN(U3050) );
  INV_X1 U6089 ( .A(n5101), .ZN(n6511) );
  NOR2_X1 U6090 ( .A1(n6443), .A2(n5156), .ZN(n4895) );
  OAI22_X1 U6091 ( .A1(n5090), .A2(n5435), .B1(n5257), .B2(n6427), .ZN(n4894)
         );
  AOI211_X1 U6092 ( .C1(n6439), .C2(INSTQUEUE_REG_3__1__SCAN_IN), .A(n4895), 
        .B(n4894), .ZN(n4896) );
  OAI21_X1 U6093 ( .B1(n4897), .B2(n6511), .A(n4896), .ZN(U3045) );
  AOI22_X1 U6094 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n4911), .B1(n5115), 
        .B2(n4910), .ZN(n4900) );
  OAI22_X1 U6095 ( .A1(n5248), .A2(n6494), .B1(n6493), .B2(n4912), .ZN(n4898)
         );
  AOI21_X1 U6096 ( .B1(n6502), .B2(n4997), .A(n4898), .ZN(n4899) );
  NAND2_X1 U6097 ( .A1(n4900), .A2(n4899), .ZN(U3092) );
  AOI22_X1 U6098 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(n4911), .B1(n5101), 
        .B2(n4910), .ZN(n4903) );
  OAI22_X1 U6099 ( .A1(n5248), .A2(n5435), .B1(n5257), .B2(n4912), .ZN(n4901)
         );
  AOI21_X1 U6100 ( .B1(n6507), .B2(n4997), .A(n4901), .ZN(n4902) );
  NAND2_X1 U6101 ( .A1(n4903), .A2(n4902), .ZN(U3093) );
  AOI22_X1 U6102 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n4911), .B1(n5119), 
        .B2(n4910), .ZN(n4906) );
  OAI22_X1 U6103 ( .A1(n5248), .A2(n6526), .B1(n6525), .B2(n4912), .ZN(n4904)
         );
  AOI21_X1 U6104 ( .B1(n6529), .B2(n4997), .A(n4904), .ZN(n4905) );
  NAND2_X1 U6105 ( .A1(n4906), .A2(n4905), .ZN(U3096) );
  AOI22_X1 U6106 ( .A1(INSTQUEUE_REG_9__6__SCAN_IN), .A2(n4911), .B1(n5108), 
        .B2(n4910), .ZN(n4909) );
  OAI22_X1 U6107 ( .A1(n5248), .A2(n5439), .B1(n5275), .B2(n4912), .ZN(n4907)
         );
  AOI21_X1 U6108 ( .B1(n6540), .B2(n4997), .A(n4907), .ZN(n4908) );
  NAND2_X1 U6109 ( .A1(n4909), .A2(n4908), .ZN(U3098) );
  AOI22_X1 U6110 ( .A1(INSTQUEUE_REG_9__7__SCAN_IN), .A2(n4911), .B1(n5129), 
        .B2(n4910), .ZN(n4915) );
  OAI22_X1 U6111 ( .A1(n5248), .A2(n5443), .B1(n5267), .B2(n4912), .ZN(n4913)
         );
  AOI21_X1 U6112 ( .B1(n6547), .B2(n4997), .A(n4913), .ZN(n4914) );
  NAND2_X1 U6113 ( .A1(n4915), .A2(n4914), .ZN(U3099) );
  INV_X1 U6114 ( .A(n4916), .ZN(n5320) );
  NOR2_X1 U6115 ( .A1(n6370), .A2(n5320), .ZN(n4917) );
  AOI211_X1 U6116 ( .C1(n6361), .C2(PHYADDRPOINTER_REG_6__SCAN_IN), .A(n4918), 
        .B(n4917), .ZN(n4920) );
  OR2_X1 U6117 ( .A1(n5326), .A2(n5930), .ZN(n4919) );
  OAI211_X1 U6118 ( .C1(n4921), .C2(n6195), .A(n4920), .B(n4919), .ZN(U2980)
         );
  AND2_X1 U6119 ( .A1(n4652), .A2(n5138), .ZN(n4999) );
  AOI21_X1 U6120 ( .B1(n6527), .B2(n4959), .A(n7056), .ZN(n4922) );
  AOI211_X1 U6121 ( .C1(n5092), .C2(n6445), .A(n6498), .B(n4922), .ZN(n4929)
         );
  AND2_X1 U6122 ( .A1(n6558), .A2(n4923), .ZN(n4960) );
  INV_X1 U6123 ( .A(n4924), .ZN(n5048) );
  NAND2_X1 U6124 ( .A1(n5048), .A2(n4925), .ZN(n5007) );
  AOI21_X1 U6125 ( .B1(n5007), .B2(STATE2_REG_2__SCAN_IN), .A(n4926), .ZN(
        n5003) );
  OAI211_X1 U6126 ( .C1(n6666), .C2(n4960), .A(n4927), .B(n5003), .ZN(n4928)
         );
  INV_X1 U6127 ( .A(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n4933) );
  NAND2_X1 U6128 ( .A1(n5092), .A2(n6484), .ZN(n5100) );
  INV_X1 U6129 ( .A(n5417), .ZN(n5099) );
  OAI22_X1 U6130 ( .A1(n5100), .A2(n6281), .B1(n5007), .B2(n5099), .ZN(n4962)
         );
  NOR2_X1 U6131 ( .A1(n6527), .A2(n6434), .ZN(n4931) );
  INV_X1 U6132 ( .A(n4960), .ZN(n4954) );
  OAI22_X1 U6133 ( .A1(n4959), .A2(n5427), .B1(n5249), .B2(n4954), .ZN(n4930)
         );
  AOI211_X1 U6134 ( .C1(n6431), .C2(n4962), .A(n4931), .B(n4930), .ZN(n4932)
         );
  OAI21_X1 U6135 ( .B1(n4966), .B2(n4933), .A(n4932), .ZN(U3119) );
  INV_X1 U6136 ( .A(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n4937) );
  NOR2_X1 U6137 ( .A1(n6527), .A2(n6430), .ZN(n4935) );
  OAI22_X1 U6138 ( .A1(n4959), .A2(n6513), .B1(n6512), .B2(n4954), .ZN(n4934)
         );
  AOI211_X1 U6139 ( .C1(n6462), .C2(n4962), .A(n4935), .B(n4934), .ZN(n4936)
         );
  OAI21_X1 U6140 ( .B1(n4966), .B2(n4937), .A(n4936), .ZN(U3118) );
  INV_X1 U6141 ( .A(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n4941) );
  NOR2_X1 U6142 ( .A1(n6527), .A2(n5156), .ZN(n4939) );
  OAI22_X1 U6143 ( .A1(n4959), .A2(n5435), .B1(n5257), .B2(n4954), .ZN(n4938)
         );
  AOI211_X1 U6144 ( .C1(n5101), .C2(n4962), .A(n4939), .B(n4938), .ZN(n4940)
         );
  OAI21_X1 U6145 ( .B1(n4966), .B2(n4941), .A(n4940), .ZN(U3117) );
  INV_X1 U6146 ( .A(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n4945) );
  NOR2_X1 U6147 ( .A1(n6527), .A2(n6442), .ZN(n4943) );
  OAI22_X1 U6148 ( .A1(n4959), .A2(n5431), .B1(n5253), .B2(n4954), .ZN(n4942)
         );
  AOI211_X1 U6149 ( .C1(n6438), .C2(n4962), .A(n4943), .B(n4942), .ZN(n4944)
         );
  OAI21_X1 U6150 ( .B1(n4966), .B2(n4945), .A(n4944), .ZN(U3121) );
  INV_X1 U6151 ( .A(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n4949) );
  NOR2_X1 U6152 ( .A1(n6527), .A2(n5164), .ZN(n4947) );
  OAI22_X1 U6153 ( .A1(n4959), .A2(n6526), .B1(n6525), .B2(n4954), .ZN(n4946)
         );
  AOI211_X1 U6154 ( .C1(n5119), .C2(n4962), .A(n4947), .B(n4946), .ZN(n4948)
         );
  OAI21_X1 U6155 ( .B1(n4966), .B2(n4949), .A(n4948), .ZN(U3120) );
  INV_X1 U6156 ( .A(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n4953) );
  NOR2_X1 U6157 ( .A1(n6527), .A2(n5168), .ZN(n4951) );
  OAI22_X1 U6158 ( .A1(n4959), .A2(n5439), .B1(n5275), .B2(n4954), .ZN(n4950)
         );
  AOI211_X1 U6159 ( .C1(n5108), .C2(n4962), .A(n4951), .B(n4950), .ZN(n4952)
         );
  OAI21_X1 U6160 ( .B1(n4966), .B2(n4953), .A(n4952), .ZN(U3122) );
  INV_X1 U6161 ( .A(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n4958) );
  NOR2_X1 U6162 ( .A1(n6527), .A2(n5160), .ZN(n4956) );
  OAI22_X1 U6163 ( .A1(n4959), .A2(n5443), .B1(n5267), .B2(n4954), .ZN(n4955)
         );
  AOI211_X1 U6164 ( .C1(n5129), .C2(n4962), .A(n4956), .B(n4955), .ZN(n4957)
         );
  OAI21_X1 U6165 ( .B1(n4966), .B2(n4958), .A(n4957), .ZN(U3123) );
  INV_X1 U6166 ( .A(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n4965) );
  INV_X1 U6167 ( .A(n4959), .ZN(n4961) );
  AOI22_X1 U6168 ( .A1(n4961), .A2(n6452), .B1(n6451), .B2(n4960), .ZN(n4964)
         );
  AOI22_X1 U6169 ( .A1(n6502), .A2(n6549), .B1(n5115), .B2(n4962), .ZN(n4963)
         );
  OAI211_X1 U6170 ( .C1(n4966), .C2(n4965), .A(n4964), .B(n4963), .ZN(U3116)
         );
  INV_X1 U6171 ( .A(n4967), .ZN(n4973) );
  INV_X1 U6172 ( .A(n4968), .ZN(n4971) );
  OR2_X1 U6173 ( .A1(n4971), .A2(n4970), .ZN(n4972) );
  AOI21_X1 U6174 ( .B1(n4973), .B2(n4972), .A(n5329), .ZN(n5190) );
  INV_X1 U6175 ( .A(n5190), .ZN(n5228) );
  CLKBUF_X1 U6176 ( .A(n4974), .Z(n5207) );
  OR2_X1 U6177 ( .A1(n4975), .A2(n5207), .ZN(n4976) );
  NAND2_X1 U6178 ( .A1(n4976), .A2(n5332), .ZN(n5219) );
  INV_X1 U6179 ( .A(n5219), .ZN(n5204) );
  AOI22_X1 U6180 ( .A1(n5846), .A2(n5204), .B1(n4405), .B2(EBX_REG_8__SCAN_IN), 
        .ZN(n4977) );
  OAI21_X1 U6181 ( .B1(n5228), .B2(n5836), .A(n4977), .ZN(U2851) );
  NAND2_X1 U6182 ( .A1(n6675), .A2(n4978), .ZN(n4979) );
  NAND2_X1 U6183 ( .A1(n4979), .A2(n6082), .ZN(n6283) );
  INV_X1 U6184 ( .A(n6283), .ZN(n5235) );
  NAND2_X1 U6185 ( .A1(n6675), .A2(n4980), .ZN(n6280) );
  INV_X1 U6186 ( .A(n6280), .ZN(n5232) );
  AOI22_X1 U6187 ( .A1(n4982), .A2(n5232), .B1(n6277), .B2(n4981), .ZN(n4995)
         );
  INV_X1 U6188 ( .A(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n4993) );
  OAI22_X1 U6189 ( .A1(n6273), .A2(n4993), .B1(n6667), .B2(n5372), .ZN(n4992)
         );
  INV_X1 U6190 ( .A(n4984), .ZN(n4985) );
  NAND3_X1 U6191 ( .A1(n4986), .A2(n5745), .A3(n4985), .ZN(n4987) );
  NAND2_X1 U6192 ( .A1(n4988), .A2(n4987), .ZN(n4989) );
  OAI22_X1 U6193 ( .A1(n6242), .A2(n4990), .B1(n6231), .B2(REIP_REG_1__SCAN_IN), .ZN(n4991) );
  AOI211_X1 U6194 ( .C1(n6247), .C2(n4993), .A(n4992), .B(n4991), .ZN(n4994)
         );
  OAI211_X1 U6195 ( .C1(n4996), .C2(n5235), .A(n4995), .B(n4994), .ZN(U2826)
         );
  NAND2_X1 U6196 ( .A1(n6028), .A2(n4999), .ZN(n6450) );
  NAND3_X1 U6197 ( .A1(n5039), .A2(n6484), .A3(n6450), .ZN(n5001) );
  AND2_X1 U6198 ( .A1(n5000), .A2(n5414), .ZN(n5006) );
  AOI21_X1 U6199 ( .B1(n5001), .B2(n6033), .A(n5006), .ZN(n5005) );
  NOR2_X1 U6200 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5002), .ZN(n5011)
         );
  OAI211_X1 U6201 ( .C1(n6666), .C2(n5011), .A(n5099), .B(n5003), .ZN(n5004)
         );
  NAND2_X1 U6202 ( .A1(n5033), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n5014) );
  NAND2_X1 U6203 ( .A1(n5006), .A2(n6484), .ZN(n5010) );
  INV_X1 U6204 ( .A(n5007), .ZN(n5008) );
  NAND2_X1 U6205 ( .A1(n5008), .A2(n5242), .ZN(n5009) );
  NAND2_X1 U6206 ( .A1(n5010), .A2(n5009), .ZN(n5036) );
  INV_X1 U6207 ( .A(n5011), .ZN(n5034) );
  OAI22_X1 U6208 ( .A1(n6450), .A2(n5156), .B1(n5257), .B2(n5034), .ZN(n5012)
         );
  AOI21_X1 U6209 ( .B1(n5101), .B2(n5036), .A(n5012), .ZN(n5013) );
  OAI211_X1 U6210 ( .C1(n5039), .C2(n5435), .A(n5014), .B(n5013), .ZN(U3085)
         );
  NAND2_X1 U6211 ( .A1(n5033), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n5017) );
  OAI22_X1 U6212 ( .A1(n6450), .A2(n6430), .B1(n6512), .B2(n5034), .ZN(n5015)
         );
  AOI21_X1 U6213 ( .B1(n6462), .B2(n5036), .A(n5015), .ZN(n5016) );
  OAI211_X1 U6214 ( .C1(n5039), .C2(n6513), .A(n5017), .B(n5016), .ZN(U3086)
         );
  NAND2_X1 U6215 ( .A1(n5033), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n5020) );
  OAI22_X1 U6216 ( .A1(n6450), .A2(n6434), .B1(n5249), .B2(n5034), .ZN(n5018)
         );
  AOI21_X1 U6217 ( .B1(n6431), .B2(n5036), .A(n5018), .ZN(n5019) );
  OAI211_X1 U6218 ( .C1(n5039), .C2(n5427), .A(n5020), .B(n5019), .ZN(U3087)
         );
  NAND2_X1 U6219 ( .A1(n5033), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n5023) );
  OAI22_X1 U6220 ( .A1(n6450), .A2(n5146), .B1(n6493), .B2(n5034), .ZN(n5021)
         );
  AOI21_X1 U6221 ( .B1(n5115), .B2(n5036), .A(n5021), .ZN(n5022) );
  OAI211_X1 U6222 ( .C1(n5039), .C2(n6494), .A(n5023), .B(n5022), .ZN(U3084)
         );
  NAND2_X1 U6223 ( .A1(n5033), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n5026) );
  OAI22_X1 U6224 ( .A1(n6450), .A2(n6442), .B1(n5253), .B2(n5034), .ZN(n5024)
         );
  AOI21_X1 U6225 ( .B1(n6438), .B2(n5036), .A(n5024), .ZN(n5025) );
  OAI211_X1 U6226 ( .C1(n5039), .C2(n5431), .A(n5026), .B(n5025), .ZN(U3089)
         );
  NAND2_X1 U6227 ( .A1(n5033), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n5029) );
  OAI22_X1 U6228 ( .A1(n6450), .A2(n5160), .B1(n5267), .B2(n5034), .ZN(n5027)
         );
  AOI21_X1 U6229 ( .B1(n5129), .B2(n5036), .A(n5027), .ZN(n5028) );
  OAI211_X1 U6230 ( .C1(n5039), .C2(n5443), .A(n5029), .B(n5028), .ZN(U3091)
         );
  NAND2_X1 U6231 ( .A1(n5033), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n5032) );
  OAI22_X1 U6232 ( .A1(n6450), .A2(n5164), .B1(n6525), .B2(n5034), .ZN(n5030)
         );
  AOI21_X1 U6233 ( .B1(n5119), .B2(n5036), .A(n5030), .ZN(n5031) );
  OAI211_X1 U6234 ( .C1(n5039), .C2(n6526), .A(n5032), .B(n5031), .ZN(U3088)
         );
  NAND2_X1 U6235 ( .A1(n5033), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n5038) );
  OAI22_X1 U6236 ( .A1(n6450), .A2(n5168), .B1(n5275), .B2(n5034), .ZN(n5035)
         );
  AOI21_X1 U6237 ( .B1(n5108), .B2(n5036), .A(n5035), .ZN(n5037) );
  OAI211_X1 U6238 ( .C1(n5039), .C2(n5439), .A(n5038), .B(n5037), .ZN(U3090)
         );
  XOR2_X1 U6239 ( .A(n4970), .B(n4971), .Z(n6342) );
  INV_X1 U6240 ( .A(n6342), .ZN(n5210) );
  INV_X1 U6241 ( .A(EAX_REG_7__SCAN_IN), .ZN(n6318) );
  OAI222_X1 U6242 ( .A1(n6114), .A2(n5210), .B1(n5411), .B2(n5040), .C1(n5860), 
        .C2(n6318), .ZN(U2884) );
  INV_X1 U6243 ( .A(DATAI_8_), .ZN(n6811) );
  INV_X1 U6244 ( .A(EAX_REG_8__SCAN_IN), .ZN(n6316) );
  OAI222_X1 U6245 ( .A1(n5228), .A2(n6114), .B1(n5411), .B2(n6811), .C1(n5860), 
        .C2(n6316), .ZN(U2883) );
  NAND2_X1 U6246 ( .A1(n6448), .A2(n5414), .ZN(n5050) );
  NAND2_X1 U6247 ( .A1(n5080), .A2(n6484), .ZN(n5041) );
  OAI21_X1 U6248 ( .B1(n5041), .B2(n5082), .A(n6033), .ZN(n5046) );
  NOR2_X1 U6249 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5042), .ZN(n5062)
         );
  OAI21_X1 U6250 ( .B1(n5062), .B2(n6666), .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), 
        .ZN(n5045) );
  NOR2_X1 U6251 ( .A1(n5242), .A2(n5043), .ZN(n5424) );
  INV_X1 U6252 ( .A(n5424), .ZN(n5044) );
  AOI211_X2 U6253 ( .C1(n5050), .C2(n5046), .A(n5045), .B(n5044), .ZN(n5087)
         );
  INV_X1 U6254 ( .A(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n5053) );
  INV_X1 U6255 ( .A(n5062), .ZN(n5079) );
  OAI22_X1 U6256 ( .A1(n5080), .A2(n5164), .B1(n6525), .B2(n5079), .ZN(n5047)
         );
  INV_X1 U6257 ( .A(n5047), .ZN(n5052) );
  NOR2_X1 U6258 ( .A1(n5048), .A2(n6573), .ZN(n5241) );
  INV_X1 U6259 ( .A(n5241), .ZN(n5049) );
  OAI22_X1 U6260 ( .A1(n5050), .A2(n6498), .B1(n5049), .B2(n5099), .ZN(n5083)
         );
  AOI22_X1 U6261 ( .A1(n5119), .A2(n5083), .B1(n5082), .B2(n6470), .ZN(n5051)
         );
  OAI211_X1 U6262 ( .C1(n5087), .C2(n5053), .A(n5052), .B(n5051), .ZN(U3136)
         );
  INV_X1 U6263 ( .A(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n5057) );
  OAI22_X1 U6264 ( .A1(n5080), .A2(n6430), .B1(n6512), .B2(n5079), .ZN(n5054)
         );
  INV_X1 U6265 ( .A(n5054), .ZN(n5056) );
  AOI22_X1 U6266 ( .A1(n6462), .A2(n5083), .B1(n5082), .B2(n6464), .ZN(n5055)
         );
  OAI211_X1 U6267 ( .C1(n5087), .C2(n5057), .A(n5056), .B(n5055), .ZN(U3134)
         );
  INV_X1 U6268 ( .A(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n5061) );
  OAI22_X1 U6269 ( .A1(n5080), .A2(n5156), .B1(n5257), .B2(n5079), .ZN(n5058)
         );
  INV_X1 U6270 ( .A(n5058), .ZN(n5060) );
  AOI22_X1 U6271 ( .A1(n5101), .A2(n5083), .B1(n5082), .B2(n6508), .ZN(n5059)
         );
  OAI211_X1 U6272 ( .C1(n5087), .C2(n5061), .A(n5060), .B(n5059), .ZN(U3133)
         );
  INV_X1 U6273 ( .A(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n5066) );
  AOI22_X1 U6274 ( .A1(n5063), .A2(n6502), .B1(n6451), .B2(n5062), .ZN(n5065)
         );
  AOI22_X1 U6275 ( .A1(n5115), .A2(n5083), .B1(n5082), .B2(n6452), .ZN(n5064)
         );
  OAI211_X1 U6276 ( .C1(n5087), .C2(n5066), .A(n5065), .B(n5064), .ZN(U3132)
         );
  INV_X1 U6277 ( .A(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n5070) );
  OAI22_X1 U6278 ( .A1(n5080), .A2(n5168), .B1(n5275), .B2(n5079), .ZN(n5067)
         );
  INV_X1 U6279 ( .A(n5067), .ZN(n5069) );
  AOI22_X1 U6280 ( .A1(n5108), .A2(n5083), .B1(n5082), .B2(n6541), .ZN(n5068)
         );
  OAI211_X1 U6281 ( .C1(n5087), .C2(n5070), .A(n5069), .B(n5068), .ZN(U3138)
         );
  INV_X1 U6282 ( .A(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n5074) );
  OAI22_X1 U6283 ( .A1(n5080), .A2(n6434), .B1(n5249), .B2(n5079), .ZN(n5071)
         );
  INV_X1 U6284 ( .A(n5071), .ZN(n5073) );
  AOI22_X1 U6285 ( .A1(n6431), .A2(n5083), .B1(n5082), .B2(n6520), .ZN(n5072)
         );
  OAI211_X1 U6286 ( .C1(n5087), .C2(n5074), .A(n5073), .B(n5072), .ZN(U3135)
         );
  INV_X1 U6287 ( .A(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n5078) );
  OAI22_X1 U6288 ( .A1(n5080), .A2(n5160), .B1(n5267), .B2(n5079), .ZN(n5075)
         );
  INV_X1 U6289 ( .A(n5075), .ZN(n5077) );
  AOI22_X1 U6290 ( .A1(n5129), .A2(n5083), .B1(n5082), .B2(n6550), .ZN(n5076)
         );
  OAI211_X1 U6291 ( .C1(n5087), .C2(n5078), .A(n5077), .B(n5076), .ZN(U3139)
         );
  INV_X1 U6292 ( .A(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n5086) );
  OAI22_X1 U6293 ( .A1(n5080), .A2(n6442), .B1(n5253), .B2(n5079), .ZN(n5081)
         );
  INV_X1 U6294 ( .A(n5081), .ZN(n5085) );
  AOI22_X1 U6295 ( .A1(n6438), .A2(n5083), .B1(n5082), .B2(n6535), .ZN(n5084)
         );
  OAI211_X1 U6296 ( .C1(n5087), .C2(n5086), .A(n5085), .B(n5084), .ZN(U3137)
         );
  OR2_X1 U6297 ( .A1(n5088), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n5141)
         );
  NOR2_X1 U6298 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5141), .ZN(n5126)
         );
  NAND2_X1 U6299 ( .A1(n6028), .A2(n5089), .ZN(n5137) );
  AOI21_X1 U6300 ( .B1(n5090), .B2(n5174), .A(n7056), .ZN(n5093) );
  AND2_X1 U6301 ( .A1(n5092), .A2(n5091), .ZN(n5135) );
  NOR2_X1 U6302 ( .A1(n5093), .A2(n5135), .ZN(n5095) );
  AOI211_X1 U6303 ( .C1(n6484), .C2(n5095), .A(n5242), .B(n5094), .ZN(n5096)
         );
  OAI21_X1 U6304 ( .B1(n5126), .B2(n6666), .A(n5096), .ZN(n5097) );
  INV_X1 U6305 ( .A(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n5104) );
  AOI22_X1 U6306 ( .A1(n5127), .A2(n6508), .B1(n6506), .B2(n5126), .ZN(n5103)
         );
  OAI22_X1 U6307 ( .A1(n5100), .A2(n5414), .B1(n5099), .B2(n5098), .ZN(n5128)
         );
  AOI22_X1 U6308 ( .A1(n6436), .A2(n6507), .B1(n5101), .B2(n5128), .ZN(n5102)
         );
  OAI211_X1 U6309 ( .C1(n5133), .C2(n5104), .A(n5103), .B(n5102), .ZN(U3053)
         );
  INV_X1 U6310 ( .A(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n5107) );
  AOI22_X1 U6311 ( .A1(n5127), .A2(n6520), .B1(n6518), .B2(n5126), .ZN(n5106)
         );
  AOI22_X1 U6312 ( .A1(n6436), .A2(n6519), .B1(n6431), .B2(n5128), .ZN(n5105)
         );
  OAI211_X1 U6313 ( .C1(n5133), .C2(n5107), .A(n5106), .B(n5105), .ZN(U3055)
         );
  INV_X1 U6314 ( .A(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n5111) );
  AOI22_X1 U6315 ( .A1(n5127), .A2(n6541), .B1(n6539), .B2(n5126), .ZN(n5110)
         );
  AOI22_X1 U6316 ( .A1(n6436), .A2(n6540), .B1(n5108), .B2(n5128), .ZN(n5109)
         );
  OAI211_X1 U6317 ( .C1(n5133), .C2(n5111), .A(n5110), .B(n5109), .ZN(U3058)
         );
  INV_X1 U6318 ( .A(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n5114) );
  AOI22_X1 U6319 ( .A1(n5127), .A2(n6464), .B1(n6463), .B2(n5126), .ZN(n5113)
         );
  AOI22_X1 U6320 ( .A1(n6436), .A2(n6515), .B1(n6462), .B2(n5128), .ZN(n5112)
         );
  OAI211_X1 U6321 ( .C1(n5133), .C2(n5114), .A(n5113), .B(n5112), .ZN(U3054)
         );
  INV_X1 U6322 ( .A(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n5118) );
  AOI22_X1 U6323 ( .A1(n5127), .A2(n6452), .B1(n6451), .B2(n5126), .ZN(n5117)
         );
  AOI22_X1 U6324 ( .A1(n6436), .A2(n6502), .B1(n5115), .B2(n5128), .ZN(n5116)
         );
  OAI211_X1 U6325 ( .C1(n5133), .C2(n5118), .A(n5117), .B(n5116), .ZN(U3052)
         );
  INV_X1 U6326 ( .A(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n5122) );
  AOI22_X1 U6327 ( .A1(n5127), .A2(n6470), .B1(n6469), .B2(n5126), .ZN(n5121)
         );
  AOI22_X1 U6328 ( .A1(n6436), .A2(n6529), .B1(n5119), .B2(n5128), .ZN(n5120)
         );
  OAI211_X1 U6329 ( .C1(n5133), .C2(n5122), .A(n5121), .B(n5120), .ZN(U3056)
         );
  INV_X1 U6330 ( .A(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n5125) );
  AOI22_X1 U6331 ( .A1(n5127), .A2(n6535), .B1(n6533), .B2(n5126), .ZN(n5124)
         );
  AOI22_X1 U6332 ( .A1(n6436), .A2(n6534), .B1(n6438), .B2(n5128), .ZN(n5123)
         );
  OAI211_X1 U6333 ( .C1(n5133), .C2(n5125), .A(n5124), .B(n5123), .ZN(U3057)
         );
  INV_X1 U6334 ( .A(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n5132) );
  AOI22_X1 U6335 ( .A1(n5127), .A2(n6550), .B1(n6546), .B2(n5126), .ZN(n5131)
         );
  AOI22_X1 U6336 ( .A1(n6436), .A2(n6547), .B1(n5129), .B2(n5128), .ZN(n5130)
         );
  OAI211_X1 U6337 ( .C1(n5133), .C2(n5132), .A(n5131), .B(n5130), .ZN(U3059)
         );
  AOI21_X1 U6338 ( .B1(n5137), .B2(n6484), .A(n5134), .ZN(n5140) );
  NOR2_X1 U6339 ( .A1(n6558), .A2(n5141), .ZN(n5172) );
  AOI21_X1 U6340 ( .B1(n5135), .B2(n6487), .A(n5172), .ZN(n5143) );
  OAI22_X1 U6341 ( .A1(n5140), .A2(n5143), .B1(n5141), .B2(n6590), .ZN(n5136)
         );
  INV_X1 U6342 ( .A(n5137), .ZN(n5139) );
  NAND2_X1 U6343 ( .A1(n5139), .A2(n5138), .ZN(n5420) );
  INV_X1 U6344 ( .A(n5140), .ZN(n5142) );
  AOI22_X1 U6345 ( .A1(n5143), .A2(n5142), .B1(n5141), .B2(n6498), .ZN(n5144)
         );
  NAND2_X1 U6346 ( .A1(n6455), .A2(n5144), .ZN(n5171) );
  AOI22_X1 U6347 ( .A1(n6451), .A2(n5172), .B1(INSTQUEUE_REG_5__0__SCAN_IN), 
        .B2(n5171), .ZN(n5145) );
  OAI21_X1 U6348 ( .B1(n5174), .B2(n5146), .A(n5145), .ZN(n5147) );
  AOI21_X1 U6349 ( .B1(n6452), .B2(n5458), .A(n5147), .ZN(n5148) );
  OAI21_X1 U6350 ( .B1(n5177), .B2(n6505), .A(n5148), .ZN(U3060) );
  INV_X1 U6351 ( .A(n6431), .ZN(n6523) );
  AOI22_X1 U6352 ( .A1(n6518), .A2(n5172), .B1(INSTQUEUE_REG_5__3__SCAN_IN), 
        .B2(n5171), .ZN(n5149) );
  OAI21_X1 U6353 ( .B1(n5174), .B2(n6434), .A(n5149), .ZN(n5150) );
  AOI21_X1 U6354 ( .B1(n6520), .B2(n5458), .A(n5150), .ZN(n5151) );
  OAI21_X1 U6355 ( .B1(n5177), .B2(n6523), .A(n5151), .ZN(U3063) );
  INV_X1 U6356 ( .A(n6462), .ZN(n5452) );
  AOI22_X1 U6357 ( .A1(n6463), .A2(n5172), .B1(INSTQUEUE_REG_5__2__SCAN_IN), 
        .B2(n5171), .ZN(n5152) );
  OAI21_X1 U6358 ( .B1(n5174), .B2(n6430), .A(n5152), .ZN(n5153) );
  AOI21_X1 U6359 ( .B1(n6464), .B2(n5458), .A(n5153), .ZN(n5154) );
  OAI21_X1 U6360 ( .B1(n5177), .B2(n5452), .A(n5154), .ZN(U3062) );
  AOI22_X1 U6361 ( .A1(n6506), .A2(n5172), .B1(INSTQUEUE_REG_5__1__SCAN_IN), 
        .B2(n5171), .ZN(n5155) );
  OAI21_X1 U6362 ( .B1(n5174), .B2(n5156), .A(n5155), .ZN(n5157) );
  AOI21_X1 U6363 ( .B1(n6508), .B2(n5458), .A(n5157), .ZN(n5158) );
  OAI21_X1 U6364 ( .B1(n5177), .B2(n6511), .A(n5158), .ZN(U3061) );
  AOI22_X1 U6365 ( .A1(n6546), .A2(n5172), .B1(INSTQUEUE_REG_5__7__SCAN_IN), 
        .B2(n5171), .ZN(n5159) );
  OAI21_X1 U6366 ( .B1(n5174), .B2(n5160), .A(n5159), .ZN(n5161) );
  AOI21_X1 U6367 ( .B1(n6550), .B2(n5458), .A(n5161), .ZN(n5162) );
  OAI21_X1 U6368 ( .B1(n5177), .B2(n6554), .A(n5162), .ZN(U3067) );
  AOI22_X1 U6369 ( .A1(n6469), .A2(n5172), .B1(INSTQUEUE_REG_5__4__SCAN_IN), 
        .B2(n5171), .ZN(n5163) );
  OAI21_X1 U6370 ( .B1(n5174), .B2(n5164), .A(n5163), .ZN(n5165) );
  AOI21_X1 U6371 ( .B1(n6470), .B2(n5458), .A(n5165), .ZN(n5166) );
  OAI21_X1 U6372 ( .B1(n5177), .B2(n6532), .A(n5166), .ZN(U3064) );
  AOI22_X1 U6373 ( .A1(n6539), .A2(n5172), .B1(INSTQUEUE_REG_5__6__SCAN_IN), 
        .B2(n5171), .ZN(n5167) );
  OAI21_X1 U6374 ( .B1(n5174), .B2(n5168), .A(n5167), .ZN(n5169) );
  AOI21_X1 U6375 ( .B1(n6541), .B2(n5458), .A(n5169), .ZN(n5170) );
  OAI21_X1 U6376 ( .B1(n5177), .B2(n6544), .A(n5170), .ZN(U3066) );
  INV_X1 U6377 ( .A(n6438), .ZN(n6538) );
  AOI22_X1 U6378 ( .A1(n6533), .A2(n5172), .B1(INSTQUEUE_REG_5__5__SCAN_IN), 
        .B2(n5171), .ZN(n5173) );
  OAI21_X1 U6379 ( .B1(n5174), .B2(n6442), .A(n5173), .ZN(n5175) );
  AOI21_X1 U6380 ( .B1(n6535), .B2(n5458), .A(n5175), .ZN(n5176) );
  OAI21_X1 U6381 ( .B1(n5177), .B2(n6538), .A(n5176), .ZN(U3065) );
  OAI21_X1 U6382 ( .B1(n5178), .B2(n5181), .A(n5180), .ZN(n5562) );
  AOI21_X1 U6383 ( .B1(n5183), .B2(n5182), .A(n5342), .ZN(n6180) );
  AOI22_X1 U6384 ( .A1(n5846), .A2(n6180), .B1(n4405), .B2(EBX_REG_13__SCAN_IN), .ZN(n5184) );
  OAI21_X1 U6385 ( .B1(n5562), .B2(n5854), .A(n5184), .ZN(U2846) );
  OAI21_X1 U6386 ( .B1(n5185), .B2(n5187), .A(n5186), .ZN(n5206) );
  INV_X1 U6387 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n5224) );
  NAND2_X1 U6388 ( .A1(n6144), .A2(n5222), .ZN(n5188) );
  NAND2_X1 U6389 ( .A1(n6371), .A2(REIP_REG_8__SCAN_IN), .ZN(n5192) );
  OAI211_X1 U6390 ( .C1(n6148), .C2(n5224), .A(n5188), .B(n5192), .ZN(n5189)
         );
  AOI21_X1 U6391 ( .B1(n5190), .B2(n6357), .A(n5189), .ZN(n5191) );
  OAI21_X1 U6392 ( .B1(n5206), .B2(n6195), .A(n5191), .ZN(U2978) );
  INV_X1 U6393 ( .A(n5192), .ZN(n5203) );
  NOR2_X1 U6394 ( .A1(n5193), .A2(n5194), .ZN(n6386) );
  OAI21_X1 U6395 ( .B1(INSTADDRPOINTER_REG_7__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_8__SCAN_IN), .A(n6386), .ZN(n5201) );
  INV_X1 U6396 ( .A(n5194), .ZN(n5196) );
  OAI21_X1 U6397 ( .B1(n5196), .B2(n5687), .A(n5195), .ZN(n5197) );
  AOI21_X1 U6398 ( .B1(n5199), .B2(n5198), .A(n5197), .ZN(n6391) );
  OAI22_X1 U6399 ( .A1(n5485), .A2(n5201), .B1(n6391), .B2(n5200), .ZN(n5202)
         );
  AOI211_X1 U6400 ( .C1(n6412), .C2(n5204), .A(n5203), .B(n5202), .ZN(n5205)
         );
  OAI21_X1 U6401 ( .B1(n5206), .B2(n6398), .A(n5205), .ZN(U3010) );
  AOI21_X1 U6402 ( .B1(n5209), .B2(n5208), .A(n5207), .ZN(n6385) );
  INV_X1 U6403 ( .A(n6385), .ZN(n5212) );
  OAI222_X1 U6404 ( .A1(n5212), .A2(n6288), .B1(n5211), .B2(n6292), .C1(n5854), 
        .C2(n5210), .ZN(U2852) );
  INV_X1 U6405 ( .A(REIP_REG_8__SCAN_IN), .ZN(n6636) );
  NOR2_X1 U6406 ( .A1(n6231), .A2(n5213), .ZN(n6267) );
  AND2_X1 U6407 ( .A1(n6267), .A2(REIP_REG_5__SCAN_IN), .ZN(n6239) );
  NAND3_X1 U6408 ( .A1(REIP_REG_7__SCAN_IN), .A2(REIP_REG_6__SCAN_IN), .A3(
        n6239), .ZN(n5309) );
  NAND2_X1 U6409 ( .A1(n6636), .A2(n5309), .ZN(n5226) );
  OR2_X1 U6410 ( .A1(n6231), .A2(n5214), .ZN(n5215) );
  NAND2_X1 U6411 ( .A1(n5215), .A2(n5372), .ZN(n6266) );
  INV_X1 U6412 ( .A(n6266), .ZN(n5218) );
  INV_X1 U6413 ( .A(n6231), .ZN(n5371) );
  NAND2_X1 U6414 ( .A1(n5371), .A2(n5216), .ZN(n5217) );
  NAND2_X1 U6415 ( .A1(n5218), .A2(n5217), .ZN(n5379) );
  OAI22_X1 U6416 ( .A1(n5220), .A2(n6242), .B1(n6218), .B2(n5219), .ZN(n5221)
         );
  AOI211_X1 U6417 ( .C1(n6247), .C2(n5222), .A(n5221), .B(n6411), .ZN(n5223)
         );
  OAI21_X1 U6418 ( .B1(n5224), .B2(n6273), .A(n5223), .ZN(n5225) );
  AOI21_X1 U6419 ( .B1(n5226), .B2(n5379), .A(n5225), .ZN(n5227) );
  OAI21_X1 U6420 ( .B1(n5228), .B2(n6082), .A(n5227), .ZN(U2819) );
  NAND2_X1 U6421 ( .A1(n6273), .A2(n6272), .ZN(n5231) );
  OAI22_X1 U6422 ( .A1(n6091), .A2(n6672), .B1(n6218), .B2(n5229), .ZN(n5230)
         );
  AOI21_X1 U6423 ( .B1(n5231), .B2(PHYADDRPOINTER_REG_0__SCAN_IN), .A(n5230), 
        .ZN(n5234) );
  AOI22_X1 U6424 ( .A1(n6487), .A2(n5232), .B1(n6276), .B2(EBX_REG_0__SCAN_IN), 
        .ZN(n5233) );
  OAI211_X1 U6425 ( .C1(n5236), .C2(n5235), .A(n5234), .B(n5233), .ZN(U2827)
         );
  INV_X1 U6426 ( .A(DATAI_13_), .ZN(n6848) );
  INV_X1 U6427 ( .A(EAX_REG_13__SCAN_IN), .ZN(n6307) );
  OAI222_X1 U6428 ( .A1(n5562), .A2(n6114), .B1(n5411), .B2(n6848), .C1(n6307), 
        .C2(n5860), .ZN(U2878) );
  AND2_X1 U6429 ( .A1(n4652), .A2(n5237), .ZN(n5419) );
  NAND3_X1 U6430 ( .A1(n5277), .A2(n5248), .A3(n6484), .ZN(n5239) );
  NAND2_X1 U6431 ( .A1(n5239), .A2(n6033), .ZN(n5245) );
  AOI22_X1 U6432 ( .A1(n5245), .A2(n6488), .B1(n5242), .B2(n5241), .ZN(n5282)
         );
  INV_X1 U6433 ( .A(n6488), .ZN(n5244) );
  NAND3_X1 U6434 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n5243), .ZN(n6497) );
  OR2_X1 U6435 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6497), .ZN(n5276)
         );
  AOI22_X1 U6436 ( .A1(n5245), .A2(n5244), .B1(STATE2_REG_3__SCAN_IN), .B2(
        n5276), .ZN(n5246) );
  OAI211_X1 U6437 ( .C1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C2(n6590), .A(n5247), .B(n5246), .ZN(n5274) );
  NAND2_X1 U6438 ( .A1(n5274), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n5252)
         );
  OAI22_X1 U6439 ( .A1(n5277), .A2(n5427), .B1(n5276), .B2(n5249), .ZN(n5250)
         );
  AOI21_X1 U6440 ( .B1(n5279), .B2(n6519), .A(n5250), .ZN(n5251) );
  OAI211_X1 U6441 ( .C1(n5282), .C2(n6523), .A(n5252), .B(n5251), .ZN(U3103)
         );
  NAND2_X1 U6442 ( .A1(n5274), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n5256)
         );
  OAI22_X1 U6443 ( .A1(n5277), .A2(n5431), .B1(n5276), .B2(n5253), .ZN(n5254)
         );
  AOI21_X1 U6444 ( .B1(n5279), .B2(n6534), .A(n5254), .ZN(n5255) );
  OAI211_X1 U6445 ( .C1(n5282), .C2(n6538), .A(n5256), .B(n5255), .ZN(U3105)
         );
  NAND2_X1 U6446 ( .A1(n5274), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n5260)
         );
  OAI22_X1 U6447 ( .A1(n5277), .A2(n5435), .B1(n5276), .B2(n5257), .ZN(n5258)
         );
  AOI21_X1 U6448 ( .B1(n5279), .B2(n6507), .A(n5258), .ZN(n5259) );
  OAI211_X1 U6449 ( .C1(n5282), .C2(n6511), .A(n5260), .B(n5259), .ZN(U3101)
         );
  NAND2_X1 U6450 ( .A1(n5274), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n5263)
         );
  OAI22_X1 U6451 ( .A1(n5277), .A2(n6513), .B1(n5276), .B2(n6512), .ZN(n5261)
         );
  AOI21_X1 U6452 ( .B1(n5279), .B2(n6515), .A(n5261), .ZN(n5262) );
  OAI211_X1 U6453 ( .C1(n5282), .C2(n5452), .A(n5263), .B(n5262), .ZN(U3102)
         );
  NAND2_X1 U6454 ( .A1(n5274), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n5266)
         );
  OAI22_X1 U6455 ( .A1(n5277), .A2(n6526), .B1(n5276), .B2(n6525), .ZN(n5264)
         );
  AOI21_X1 U6456 ( .B1(n5279), .B2(n6529), .A(n5264), .ZN(n5265) );
  OAI211_X1 U6457 ( .C1(n5282), .C2(n6532), .A(n5266), .B(n5265), .ZN(U3104)
         );
  NAND2_X1 U6458 ( .A1(n5274), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n5270)
         );
  OAI22_X1 U6459 ( .A1(n5277), .A2(n5443), .B1(n5276), .B2(n5267), .ZN(n5268)
         );
  AOI21_X1 U6460 ( .B1(n5279), .B2(n6547), .A(n5268), .ZN(n5269) );
  OAI211_X1 U6461 ( .C1(n5282), .C2(n6554), .A(n5270), .B(n5269), .ZN(U3107)
         );
  NAND2_X1 U6462 ( .A1(n5274), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n5273)
         );
  OAI22_X1 U6463 ( .A1(n5277), .A2(n6494), .B1(n6493), .B2(n5276), .ZN(n5271)
         );
  AOI21_X1 U6464 ( .B1(n5279), .B2(n6502), .A(n5271), .ZN(n5272) );
  OAI211_X1 U6465 ( .C1(n5282), .C2(n6505), .A(n5273), .B(n5272), .ZN(U3100)
         );
  NAND2_X1 U6466 ( .A1(n5274), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n5281)
         );
  OAI22_X1 U6467 ( .A1(n5277), .A2(n5439), .B1(n5276), .B2(n5275), .ZN(n5278)
         );
  AOI21_X1 U6468 ( .B1(n5279), .B2(n6540), .A(n5278), .ZN(n5280) );
  OAI211_X1 U6469 ( .C1(n5282), .C2(n6544), .A(n5281), .B(n5280), .ZN(U3106)
         );
  OR3_X1 U6470 ( .A1(n6231), .A2(REIP_REG_4__SCAN_IN), .A3(n5289), .ZN(n5287)
         );
  OAI22_X1 U6471 ( .A1(n5283), .A2(n6242), .B1(n6218), .B2(n6394), .ZN(n5284)
         );
  AOI211_X1 U6472 ( .C1(n6247), .C2(n5285), .A(n5284), .B(n6411), .ZN(n5286)
         );
  OAI211_X1 U6473 ( .C1(n5288), .C2(n6280), .A(n5287), .B(n5286), .ZN(n5292)
         );
  INV_X1 U6474 ( .A(n6091), .ZN(n5295) );
  OAI21_X1 U6475 ( .B1(n5296), .B2(n5289), .A(n5295), .ZN(n6286) );
  OAI22_X1 U6476 ( .A1(n6286), .A2(n6630), .B1(n5290), .B2(n6273), .ZN(n5291)
         );
  AOI211_X1 U6477 ( .C1(n5293), .C2(n6283), .A(n5292), .B(n5291), .ZN(n5294)
         );
  INV_X1 U6478 ( .A(n5294), .ZN(U2823) );
  OAI21_X1 U6479 ( .B1(n5296), .B2(n6230), .A(n5295), .ZN(n6251) );
  INV_X1 U6480 ( .A(n6251), .ZN(n5305) );
  INV_X1 U6481 ( .A(REIP_REG_13__SCAN_IN), .ZN(n6642) );
  AOI22_X1 U6482 ( .A1(n6640), .A2(REIP_REG_13__SCAN_IN), .B1(n6642), .B2(
        n5297), .ZN(n5300) );
  INV_X1 U6483 ( .A(n5558), .ZN(n5298) );
  NAND2_X1 U6484 ( .A1(n6247), .A2(n5298), .ZN(n5299) );
  OAI21_X1 U6485 ( .B1(n6231), .B2(n5300), .A(n5299), .ZN(n5304) );
  AOI22_X1 U6486 ( .A1(EBX_REG_13__SCAN_IN), .A2(n6276), .B1(n6277), .B2(n6180), .ZN(n5301) );
  OAI211_X1 U6487 ( .C1(n6273), .C2(n5302), .A(n5301), .B(n6393), .ZN(n5303)
         );
  AOI211_X1 U6488 ( .C1(REIP_REG_13__SCAN_IN), .C2(n5305), .A(n5304), .B(n5303), .ZN(n5306) );
  OAI21_X1 U6489 ( .B1(n5562), .B2(n6082), .A(n5306), .ZN(U2814) );
  INV_X1 U6490 ( .A(n5307), .ZN(n5308) );
  INV_X1 U6491 ( .A(n5355), .ZN(n5327) );
  AND2_X1 U6492 ( .A1(n5355), .A2(n5307), .ZN(n5404) );
  AOI21_X1 U6493 ( .B1(n5308), .B2(n5327), .A(n5404), .ZN(n5482) );
  INV_X1 U6494 ( .A(n5482), .ZN(n5394) );
  NOR2_X1 U6495 ( .A1(n6636), .A2(n5309), .ZN(n5385) );
  XNOR2_X1 U6496 ( .A(REIP_REG_10__SCAN_IN), .B(n6637), .ZN(n5317) );
  INV_X1 U6497 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n5311) );
  NAND2_X1 U6498 ( .A1(n5379), .A2(REIP_REG_10__SCAN_IN), .ZN(n5310) );
  OAI211_X1 U6499 ( .C1(n6273), .C2(n5311), .A(n5310), .B(n6393), .ZN(n5316)
         );
  OAI21_X1 U6500 ( .B1(n5313), .B2(n5331), .A(n5408), .ZN(n5484) );
  AOI22_X1 U6501 ( .A1(EBX_REG_10__SCAN_IN), .A2(n6276), .B1(n5478), .B2(n6247), .ZN(n5314) );
  OAI21_X1 U6502 ( .B1(n6218), .B2(n5484), .A(n5314), .ZN(n5315) );
  AOI211_X1 U6503 ( .C1(n5385), .C2(n5317), .A(n5316), .B(n5315), .ZN(n5318)
         );
  OAI21_X1 U6504 ( .B1(n5394), .B2(n6082), .A(n5318), .ZN(U2817) );
  INV_X1 U6505 ( .A(n6239), .ZN(n6253) );
  NOR2_X1 U6506 ( .A1(REIP_REG_6__SCAN_IN), .A2(n6253), .ZN(n6259) );
  INV_X1 U6507 ( .A(n6259), .ZN(n5319) );
  OAI21_X1 U6508 ( .B1(n6272), .B2(n5320), .A(n5319), .ZN(n5324) );
  AOI22_X1 U6509 ( .A1(EBX_REG_6__SCAN_IN), .A2(n6276), .B1(
        PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n6229), .ZN(n5321) );
  OAI211_X1 U6510 ( .C1(n6218), .C2(n5322), .A(n5321), .B(n6393), .ZN(n5323)
         );
  AOI211_X1 U6511 ( .C1(REIP_REG_6__SCAN_IN), .C2(n6266), .A(n5324), .B(n5323), 
        .ZN(n5325) );
  OAI21_X1 U6512 ( .B1(n6082), .B2(n5326), .A(n5325), .ZN(U2821) );
  OAI21_X1 U6513 ( .B1(n5329), .B2(n5328), .A(n5327), .ZN(n5393) );
  INV_X1 U6514 ( .A(DATAI_9_), .ZN(n6846) );
  INV_X1 U6515 ( .A(EAX_REG_9__SCAN_IN), .ZN(n6314) );
  OAI222_X1 U6516 ( .A1(n5393), .A2(n6114), .B1(n5411), .B2(n6846), .C1(n5860), 
        .C2(n6314), .ZN(U2882) );
  INV_X1 U6517 ( .A(EAX_REG_10__SCAN_IN), .ZN(n6312) );
  OAI222_X1 U6518 ( .A1(n5394), .A2(n6114), .B1(n5411), .B2(n5330), .C1(n5860), 
        .C2(n6312), .ZN(U2881) );
  AOI21_X1 U6519 ( .B1(n5333), .B2(n5332), .A(n5331), .ZN(n6379) );
  INV_X1 U6520 ( .A(n6379), .ZN(n5335) );
  OAI222_X1 U6521 ( .A1(n5335), .A2(n6288), .B1(n5334), .B2(n6292), .C1(n5393), 
        .C2(n5854), .ZN(U2850) );
  AND3_X1 U6522 ( .A1(n5180), .A2(n5339), .A3(n5338), .ZN(n5340) );
  OR2_X1 U6523 ( .A1(n5337), .A2(n5340), .ZN(n5571) );
  INV_X1 U6524 ( .A(EBX_REG_14__SCAN_IN), .ZN(n5344) );
  OAI21_X1 U6525 ( .B1(n5343), .B2(n5342), .A(n5341), .ZN(n5585) );
  OAI222_X1 U6526 ( .A1(n5571), .A2(n5854), .B1(n6292), .B2(n5344), .C1(n5585), 
        .C2(n6288), .ZN(U2845) );
  INV_X1 U6527 ( .A(EAX_REG_14__SCAN_IN), .ZN(n6305) );
  OAI222_X1 U6528 ( .A1(n5571), .A2(n6114), .B1(n5411), .B2(n5345), .C1(n5860), 
        .C2(n6305), .ZN(U2877) );
  NAND2_X1 U6529 ( .A1(n6365), .A2(n6283), .ZN(n5353) );
  OAI21_X1 U6530 ( .B1(n6231), .B2(REIP_REG_1__SCAN_IN), .A(n5372), .ZN(n6270)
         );
  INV_X1 U6531 ( .A(REIP_REG_2__SCAN_IN), .ZN(n5346) );
  NAND3_X1 U6532 ( .A1(n5371), .A2(REIP_REG_1__SCAN_IN), .A3(n5346), .ZN(n5348) );
  NAND2_X1 U6533 ( .A1(n6229), .A2(PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n5347)
         );
  OAI211_X1 U6534 ( .C1(n6272), .C2(n6369), .A(n5348), .B(n5347), .ZN(n5351)
         );
  OAI22_X1 U6535 ( .A1(n6242), .A2(n5349), .B1(n4527), .B2(n6280), .ZN(n5350)
         );
  AOI211_X1 U6536 ( .C1(REIP_REG_2__SCAN_IN), .C2(n6270), .A(n5351), .B(n5350), 
        .ZN(n5352) );
  OAI211_X1 U6537 ( .C1(n6410), .C2(n6218), .A(n5353), .B(n5352), .ZN(U2825)
         );
  NAND2_X1 U6538 ( .A1(n5355), .A2(n5354), .ZN(n5405) );
  NAND2_X1 U6539 ( .A1(n5405), .A2(n5356), .ZN(n5357) );
  AND2_X1 U6540 ( .A1(n5358), .A2(n5357), .ZN(n6235) );
  INV_X1 U6541 ( .A(n6235), .ZN(n5402) );
  XOR2_X1 U6542 ( .A(n5407), .B(n5359), .Z(n6228) );
  AOI22_X1 U6543 ( .A1(n5846), .A2(n6228), .B1(EBX_REG_12__SCAN_IN), .B2(n4405), .ZN(n5360) );
  OAI21_X1 U6544 ( .B1(n5402), .B2(n5836), .A(n5360), .ZN(U2847) );
  NOR2_X1 U6545 ( .A1(n5337), .A2(n5363), .ZN(n5364) );
  OR2_X1 U6546 ( .A1(n5362), .A2(n5364), .ZN(n5548) );
  AOI21_X1 U6547 ( .B1(n5365), .B2(n5341), .A(n5464), .ZN(n5541) );
  INV_X1 U6548 ( .A(n5547), .ZN(n5368) );
  INV_X1 U6549 ( .A(REIP_REG_15__SCAN_IN), .ZN(n5366) );
  NAND2_X1 U6550 ( .A1(n5369), .A2(n5366), .ZN(n5367) );
  OAI22_X1 U6551 ( .A1(n6272), .A2(n5368), .B1(n6231), .B2(n5367), .ZN(n5376)
         );
  INV_X1 U6552 ( .A(n5369), .ZN(n5370) );
  NAND2_X1 U6553 ( .A1(n5371), .A2(n5370), .ZN(n5396) );
  NAND2_X1 U6554 ( .A1(n5396), .A2(n5372), .ZN(n5400) );
  AOI22_X1 U6555 ( .A1(EBX_REG_15__SCAN_IN), .A2(n6276), .B1(
        REIP_REG_15__SCAN_IN), .B2(n5400), .ZN(n5373) );
  OAI211_X1 U6556 ( .C1(n6273), .C2(n5374), .A(n5373), .B(n6393), .ZN(n5375)
         );
  AOI211_X1 U6557 ( .C1(n5541), .C2(n6277), .A(n5376), .B(n5375), .ZN(n5377)
         );
  OAI21_X1 U6558 ( .B1(n5548), .B2(n6082), .A(n5377), .ZN(U2812) );
  AOI22_X1 U6559 ( .A1(n5846), .A2(n5541), .B1(EBX_REG_15__SCAN_IN), .B2(n4405), .ZN(n5378) );
  OAI21_X1 U6560 ( .B1(n5548), .B2(n5836), .A(n5378), .ZN(U2844) );
  INV_X1 U6561 ( .A(n5379), .ZN(n5380) );
  OAI22_X1 U6562 ( .A1(n5380), .A2(n6637), .B1(n5389), .B2(n6272), .ZN(n5384)
         );
  AOI22_X1 U6563 ( .A1(EBX_REG_9__SCAN_IN), .A2(n6276), .B1(n6277), .B2(n6379), 
        .ZN(n5381) );
  OAI211_X1 U6564 ( .C1(n6273), .C2(n5382), .A(n5381), .B(n6393), .ZN(n5383)
         );
  AOI211_X1 U6565 ( .C1(n5385), .C2(n6637), .A(n5384), .B(n5383), .ZN(n5386)
         );
  OAI21_X1 U6566 ( .B1(n5393), .B2(n6082), .A(n5386), .ZN(U2818) );
  XNOR2_X1 U6567 ( .A(n4294), .B(n5486), .ZN(n5388) );
  XNOR2_X1 U6568 ( .A(n5387), .B(n5388), .ZN(n6381) );
  NAND2_X1 U6569 ( .A1(n6381), .A2(n6366), .ZN(n5392) );
  AND2_X1 U6570 ( .A1(n6411), .A2(REIP_REG_9__SCAN_IN), .ZN(n6378) );
  NOR2_X1 U6571 ( .A1(n6370), .A2(n5389), .ZN(n5390) );
  AOI211_X1 U6572 ( .C1(n6361), .C2(PHYADDRPOINTER_REG_9__SCAN_IN), .A(n6378), 
        .B(n5390), .ZN(n5391) );
  OAI211_X1 U6573 ( .C1(n5930), .C2(n5393), .A(n5392), .B(n5391), .ZN(U2977)
         );
  OAI222_X1 U6574 ( .A1(n5484), .A2(n6288), .B1(n6292), .B2(n4123), .C1(n5394), 
        .C2(n5854), .ZN(U2849) );
  OAI22_X1 U6575 ( .A1(n6218), .A2(n5585), .B1(n5567), .B2(n6272), .ZN(n5399)
         );
  AOI22_X1 U6576 ( .A1(EBX_REG_14__SCAN_IN), .A2(n6276), .B1(
        PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n6229), .ZN(n5395) );
  OAI211_X1 U6577 ( .C1(n5397), .C2(n5396), .A(n5395), .B(n6393), .ZN(n5398)
         );
  AOI211_X1 U6578 ( .C1(REIP_REG_14__SCAN_IN), .C2(n5400), .A(n5399), .B(n5398), .ZN(n5401) );
  OAI21_X1 U6579 ( .B1(n5571), .B2(n6082), .A(n5401), .ZN(U2813) );
  INV_X1 U6580 ( .A(DATAI_12_), .ZN(n7015) );
  OAI222_X1 U6581 ( .A1(n5402), .A2(n6114), .B1(n5411), .B2(n7015), .C1(n5860), 
        .C2(n3597), .ZN(U2879) );
  OR2_X1 U6582 ( .A1(n5404), .A2(n5403), .ZN(n5406) );
  INV_X1 U6583 ( .A(n6248), .ZN(n5412) );
  AOI21_X1 U6584 ( .B1(n5409), .B2(n5408), .A(n5407), .ZN(n6372) );
  AOI22_X1 U6585 ( .A1(n5846), .A2(n6372), .B1(n4405), .B2(EBX_REG_11__SCAN_IN), .ZN(n5410) );
  OAI21_X1 U6586 ( .B1(n5412), .B2(n5854), .A(n5410), .ZN(U2848) );
  OAI222_X1 U6587 ( .A1(n5548), .A2(n6114), .B1(n5411), .B2(n6795), .C1(n5860), 
        .C2(n4421), .ZN(U2876) );
  INV_X1 U6588 ( .A(DATAI_11_), .ZN(n6769) );
  INV_X1 U6589 ( .A(EAX_REG_11__SCAN_IN), .ZN(n6310) );
  OAI222_X1 U6590 ( .A1(n5412), .A2(n6114), .B1(n5411), .B2(n6769), .C1(n5860), 
        .C2(n6310), .ZN(U2880) );
  INV_X1 U6591 ( .A(n5413), .ZN(n5418) );
  INV_X1 U6592 ( .A(n6448), .ZN(n5415) );
  NOR3_X1 U6593 ( .A1(n5415), .A2(n5414), .A3(n6498), .ZN(n5416) );
  AOI21_X1 U6594 ( .B1(n5418), .B2(n5417), .A(n5416), .ZN(n5460) );
  NAND2_X1 U6595 ( .A1(n6558), .A2(n6457), .ZN(n5423) );
  INV_X1 U6596 ( .A(n5423), .ZN(n5454) );
  NAND3_X1 U6597 ( .A1(n6484), .A2(n5420), .A3(n5456), .ZN(n5421) );
  AOI21_X1 U6598 ( .B1(n5421), .B2(n6033), .A(n6448), .ZN(n5422) );
  AOI21_X1 U6599 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n5423), .A(n5422), .ZN(
        n5425) );
  NAND3_X1 U6600 ( .A1(n6573), .A2(n5425), .A3(n5424), .ZN(n5453) );
  AOI22_X1 U6601 ( .A1(n6518), .A2(n5454), .B1(INSTQUEUE_REG_6__3__SCAN_IN), 
        .B2(n5453), .ZN(n5426) );
  OAI21_X1 U6602 ( .B1(n5456), .B2(n5427), .A(n5426), .ZN(n5428) );
  AOI21_X1 U6603 ( .B1(n6519), .B2(n5458), .A(n5428), .ZN(n5429) );
  OAI21_X1 U6604 ( .B1(n5460), .B2(n6523), .A(n5429), .ZN(U3071) );
  AOI22_X1 U6605 ( .A1(n6533), .A2(n5454), .B1(INSTQUEUE_REG_6__5__SCAN_IN), 
        .B2(n5453), .ZN(n5430) );
  OAI21_X1 U6606 ( .B1(n5456), .B2(n5431), .A(n5430), .ZN(n5432) );
  AOI21_X1 U6607 ( .B1(n6534), .B2(n5458), .A(n5432), .ZN(n5433) );
  OAI21_X1 U6608 ( .B1(n5460), .B2(n6538), .A(n5433), .ZN(U3073) );
  AOI22_X1 U6609 ( .A1(n6506), .A2(n5454), .B1(INSTQUEUE_REG_6__1__SCAN_IN), 
        .B2(n5453), .ZN(n5434) );
  OAI21_X1 U6610 ( .B1(n5456), .B2(n5435), .A(n5434), .ZN(n5436) );
  AOI21_X1 U6611 ( .B1(n6507), .B2(n5458), .A(n5436), .ZN(n5437) );
  OAI21_X1 U6612 ( .B1(n5460), .B2(n6511), .A(n5437), .ZN(U3069) );
  AOI22_X1 U6613 ( .A1(n6539), .A2(n5454), .B1(INSTQUEUE_REG_6__6__SCAN_IN), 
        .B2(n5453), .ZN(n5438) );
  OAI21_X1 U6614 ( .B1(n5456), .B2(n5439), .A(n5438), .ZN(n5440) );
  AOI21_X1 U6615 ( .B1(n6540), .B2(n5458), .A(n5440), .ZN(n5441) );
  OAI21_X1 U6616 ( .B1(n5460), .B2(n6544), .A(n5441), .ZN(U3074) );
  AOI22_X1 U6617 ( .A1(n6546), .A2(n5454), .B1(INSTQUEUE_REG_6__7__SCAN_IN), 
        .B2(n5453), .ZN(n5442) );
  OAI21_X1 U6618 ( .B1(n5456), .B2(n5443), .A(n5442), .ZN(n5444) );
  AOI21_X1 U6619 ( .B1(n6547), .B2(n5458), .A(n5444), .ZN(n5445) );
  OAI21_X1 U6620 ( .B1(n5460), .B2(n6554), .A(n5445), .ZN(U3075) );
  AOI22_X1 U6621 ( .A1(n6451), .A2(n5454), .B1(INSTQUEUE_REG_6__0__SCAN_IN), 
        .B2(n5453), .ZN(n5446) );
  OAI21_X1 U6622 ( .B1(n5456), .B2(n6494), .A(n5446), .ZN(n5447) );
  AOI21_X1 U6623 ( .B1(n6502), .B2(n5458), .A(n5447), .ZN(n5448) );
  OAI21_X1 U6624 ( .B1(n5460), .B2(n6505), .A(n5448), .ZN(U3068) );
  AOI22_X1 U6625 ( .A1(n6463), .A2(n5454), .B1(INSTQUEUE_REG_6__2__SCAN_IN), 
        .B2(n5453), .ZN(n5449) );
  OAI21_X1 U6626 ( .B1(n5456), .B2(n6513), .A(n5449), .ZN(n5450) );
  AOI21_X1 U6627 ( .B1(n6515), .B2(n5458), .A(n5450), .ZN(n5451) );
  OAI21_X1 U6628 ( .B1(n5460), .B2(n5452), .A(n5451), .ZN(U3070) );
  AOI22_X1 U6629 ( .A1(n6469), .A2(n5454), .B1(INSTQUEUE_REG_6__4__SCAN_IN), 
        .B2(n5453), .ZN(n5455) );
  OAI21_X1 U6630 ( .B1(n5456), .B2(n6526), .A(n5455), .ZN(n5457) );
  AOI21_X1 U6631 ( .B1(n6529), .B2(n5458), .A(n5457), .ZN(n5459) );
  OAI21_X1 U6632 ( .B1(n5460), .B2(n6532), .A(n5459), .ZN(U3072) );
  OAI21_X1 U6633 ( .B1(n5362), .B2(n5463), .A(n5462), .ZN(n5929) );
  INV_X1 U6634 ( .A(n5925), .ZN(n5473) );
  XNOR2_X1 U6635 ( .A(n5465), .B(n5464), .ZN(n6170) );
  AOI21_X1 U6636 ( .B1(n6229), .B2(PHYADDRPOINTER_REG_16__SCAN_IN), .A(n6411), 
        .ZN(n5466) );
  OAI21_X1 U6637 ( .B1(n6218), .B2(n6170), .A(n5466), .ZN(n5472) );
  NAND2_X1 U6638 ( .A1(n5467), .A2(REIP_REG_16__SCAN_IN), .ZN(n5470) );
  AOI22_X1 U6639 ( .A1(EBX_REG_16__SCAN_IN), .A2(n6276), .B1(n5468), .B2(n7038), .ZN(n5469) );
  OAI21_X1 U6640 ( .B1(n6091), .B2(n5470), .A(n5469), .ZN(n5471) );
  AOI211_X1 U6641 ( .C1(n6247), .C2(n5473), .A(n5472), .B(n5471), .ZN(n5474)
         );
  OAI21_X1 U6642 ( .B1(n5929), .B2(n6082), .A(n5474), .ZN(U2811) );
  NAND2_X1 U6643 ( .A1(n5498), .A2(n5475), .ZN(n5477) );
  XOR2_X1 U6644 ( .A(n5477), .B(n5476), .Z(n5490) );
  INV_X1 U6645 ( .A(n5478), .ZN(n5480) );
  AOI22_X1 U6646 ( .A1(n6361), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .B1(n6411), 
        .B2(REIP_REG_10__SCAN_IN), .ZN(n5479) );
  OAI21_X1 U6647 ( .B1(n5480), .B2(n6370), .A(n5479), .ZN(n5481) );
  AOI21_X1 U6648 ( .B1(n5482), .B2(n6357), .A(n5481), .ZN(n5483) );
  OAI21_X1 U6649 ( .B1(n5490), .B2(n6195), .A(n5483), .ZN(U2976) );
  INV_X1 U6650 ( .A(n5633), .ZN(n5713) );
  OAI21_X1 U6651 ( .B1(n5713), .B2(n5485), .A(n6391), .ZN(n6380) );
  OAI22_X1 U6652 ( .A1(n6395), .A2(n5484), .B1(n6638), .B2(n6393), .ZN(n5488)
         );
  NAND2_X1 U6653 ( .A1(n5485), .A2(n6386), .ZN(n6384) );
  AOI221_X1 U6654 ( .B1(INSTADDRPOINTER_REG_9__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .C1(n5486), .C2(n4298), .A(n6384), 
        .ZN(n5487) );
  AOI211_X1 U6655 ( .C1(INSTADDRPOINTER_REG_10__SCAN_IN), .C2(n6380), .A(n5488), .B(n5487), .ZN(n5489) );
  OAI21_X1 U6656 ( .B1(n5490), .B2(n6398), .A(n5489), .ZN(U3008) );
  AOI22_X1 U6657 ( .A1(n6296), .A2(DATAI_16_), .B1(n6299), .B2(
        EAX_REG_16__SCAN_IN), .ZN(n5495) );
  NOR2_X1 U6658 ( .A1(n5731), .A2(n5492), .ZN(n5493) );
  NAND2_X1 U6659 ( .A1(n5860), .A2(n5493), .ZN(n5861) );
  NAND2_X1 U6660 ( .A1(n6300), .A2(DATAI_0_), .ZN(n5494) );
  OAI211_X1 U6661 ( .C1(n5929), .C2(n6114), .A(n5495), .B(n5494), .ZN(U2875)
         );
  OAI222_X1 U6662 ( .A1(n5836), .A2(n5929), .B1(n5496), .B2(n6292), .C1(n6288), 
        .C2(n6170), .ZN(U2843) );
  NAND2_X1 U6663 ( .A1(n5497), .A2(n5498), .ZN(n5500) );
  XNOR2_X1 U6664 ( .A(n4294), .B(n5573), .ZN(n5499) );
  XNOR2_X1 U6665 ( .A(n5500), .B(n5499), .ZN(n6373) );
  INV_X1 U6666 ( .A(n6373), .ZN(n5504) );
  AOI22_X1 U6667 ( .A1(n6361), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .B1(n6411), 
        .B2(REIP_REG_11__SCAN_IN), .ZN(n5501) );
  OAI21_X1 U6668 ( .B1(n6245), .B2(n6370), .A(n5501), .ZN(n5502) );
  AOI21_X1 U6669 ( .B1(n6248), .B2(n6357), .A(n5502), .ZN(n5503) );
  OAI21_X1 U6670 ( .B1(n5504), .B2(n6195), .A(n5503), .ZN(U2975) );
  INV_X1 U6671 ( .A(n5554), .ZN(n5506) );
  NOR2_X1 U6672 ( .A1(n5553), .A2(n5506), .ZN(n5507) );
  XNOR2_X1 U6673 ( .A(n5505), .B(n5507), .ZN(n5516) );
  AOI22_X1 U6674 ( .A1(n6361), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .B1(n6411), 
        .B2(REIP_REG_12__SCAN_IN), .ZN(n5508) );
  OAI21_X1 U6675 ( .B1(n5509), .B2(n6370), .A(n5508), .ZN(n5510) );
  AOI21_X1 U6676 ( .B1(n6235), .B2(n6357), .A(n5510), .ZN(n5511) );
  OAI21_X1 U6677 ( .B1(n5516), .B2(n6195), .A(n5511), .ZN(U2974) );
  NOR3_X1 U6678 ( .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n6186), .A3(n5573), 
        .ZN(n5513) );
  NOR2_X1 U6679 ( .A1(n6393), .A2(n6640), .ZN(n5512) );
  AOI211_X1 U6680 ( .C1(n6412), .C2(n6228), .A(n5513), .B(n5512), .ZN(n5515)
         );
  NAND2_X1 U6681 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n5579), .ZN(n6374) );
  NAND3_X1 U6682 ( .A1(n5992), .A2(INSTADDRPOINTER_REG_12__SCAN_IN), .A3(n6374), .ZN(n5514) );
  OAI211_X1 U6683 ( .C1(n5516), .C2(n6398), .A(n5515), .B(n5514), .ZN(U3006)
         );
  INV_X1 U6684 ( .A(n5517), .ZN(n5518) );
  NAND2_X1 U6685 ( .A1(n5518), .A2(n5776), .ZN(n5519) );
  OAI21_X1 U6686 ( .B1(n5594), .B2(n5776), .A(n5519), .ZN(n5520) );
  INV_X1 U6687 ( .A(n6165), .ZN(n5521) );
  NAND2_X1 U6688 ( .A1(n5520), .A2(n5521), .ZN(n5534) );
  OR2_X1 U6689 ( .A1(n5521), .A2(n5520), .ZN(n5522) );
  NAND2_X1 U6690 ( .A1(n5534), .A2(n5522), .ZN(n6217) );
  AOI21_X1 U6691 ( .B1(n5527), .B2(n5524), .A(n5526), .ZN(n6293) );
  INV_X1 U6692 ( .A(n6293), .ZN(n5921) );
  OAI222_X1 U6693 ( .A1(n6217), .A2(n6288), .B1(n6292), .B2(n4151), .C1(n5921), 
        .C2(n5854), .ZN(U2841) );
  INV_X1 U6694 ( .A(n5528), .ZN(n5532) );
  INV_X1 U6695 ( .A(n5526), .ZN(n5531) );
  AOI21_X1 U6696 ( .B1(n5532), .B2(n5531), .A(n5530), .ZN(n6133) );
  INV_X1 U6697 ( .A(n6133), .ZN(n5536) );
  XNOR2_X1 U6698 ( .A(n5534), .B(n5533), .ZN(n6008) );
  INV_X1 U6699 ( .A(n6008), .ZN(n6097) );
  AOI22_X1 U6700 ( .A1(n5846), .A2(n6097), .B1(EBX_REG_19__SCAN_IN), .B2(n4405), .ZN(n5535) );
  OAI21_X1 U6701 ( .B1(n5536), .B2(n5854), .A(n5535), .ZN(U2840) );
  XNOR2_X1 U6702 ( .A(n4294), .B(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5538)
         );
  XNOR2_X1 U6703 ( .A(n3166), .B(n5538), .ZN(n5552) );
  OAI21_X1 U6704 ( .B1(n5713), .B2(n6169), .A(n5579), .ZN(n6173) );
  INV_X1 U6705 ( .A(n6186), .ZN(n6375) );
  AND2_X1 U6706 ( .A1(n6375), .A2(n6169), .ZN(n5540) );
  AOI22_X1 U6707 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n6173), .B1(n5540), .B2(n5539), .ZN(n5543) );
  AND2_X1 U6708 ( .A1(n6411), .A2(REIP_REG_15__SCAN_IN), .ZN(n5544) );
  AOI21_X1 U6709 ( .B1(n6412), .B2(n5541), .A(n5544), .ZN(n5542) );
  OAI211_X1 U6710 ( .C1(n5552), .C2(n6398), .A(n5543), .B(n5542), .ZN(U3003)
         );
  INV_X1 U6711 ( .A(n5544), .ZN(n5545) );
  OAI21_X1 U6712 ( .B1(n6148), .B2(n5374), .A(n5545), .ZN(n5546) );
  AOI21_X1 U6713 ( .B1(n6144), .B2(n5547), .A(n5546), .ZN(n5551) );
  INV_X1 U6714 ( .A(n5548), .ZN(n5549) );
  NAND2_X1 U6715 ( .A1(n5549), .A2(n6357), .ZN(n5550) );
  OAI211_X1 U6716 ( .C1(n5552), .C2(n6195), .A(n5551), .B(n5550), .ZN(U2971)
         );
  OR2_X1 U6717 ( .A1(n5505), .A2(n5553), .ZN(n5555) );
  NAND2_X1 U6718 ( .A1(n5555), .A2(n5554), .ZN(n5557) );
  XNOR2_X1 U6719 ( .A(n5557), .B(n5556), .ZN(n6182) );
  NAND2_X1 U6720 ( .A1(n6182), .A2(n6366), .ZN(n5561) );
  AND2_X1 U6721 ( .A1(n6411), .A2(REIP_REG_13__SCAN_IN), .ZN(n6179) );
  NOR2_X1 U6722 ( .A1(n6370), .A2(n5558), .ZN(n5559) );
  AOI211_X1 U6723 ( .C1(n6361), .C2(PHYADDRPOINTER_REG_13__SCAN_IN), .A(n6179), 
        .B(n5559), .ZN(n5560) );
  OAI211_X1 U6724 ( .C1(n5930), .C2(n5562), .A(n5561), .B(n5560), .ZN(U2973)
         );
  NAND2_X1 U6725 ( .A1(n5564), .A2(n5563), .ZN(n5566) );
  XNOR2_X1 U6726 ( .A(n4294), .B(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5565)
         );
  XNOR2_X1 U6727 ( .A(n5566), .B(n5565), .ZN(n5584) );
  NAND2_X1 U6728 ( .A1(n5584), .A2(n6366), .ZN(n5570) );
  AND2_X1 U6729 ( .A1(n6411), .A2(REIP_REG_14__SCAN_IN), .ZN(n5588) );
  NOR2_X1 U6730 ( .A1(n6370), .A2(n5567), .ZN(n5568) );
  AOI211_X1 U6731 ( .C1(n6361), .C2(PHYADDRPOINTER_REG_14__SCAN_IN), .A(n5588), 
        .B(n5568), .ZN(n5569) );
  OAI211_X1 U6732 ( .C1(n5930), .C2(n5571), .A(n5570), .B(n5569), .ZN(U2972)
         );
  NOR2_X1 U6733 ( .A1(n5573), .A2(n5572), .ZN(n5581) );
  NAND2_X1 U6734 ( .A1(n5574), .A2(n5581), .ZN(n6185) );
  INV_X1 U6735 ( .A(n6185), .ZN(n5583) );
  OR2_X1 U6736 ( .A1(n5576), .A2(n5575), .ZN(n5582) );
  NAND2_X1 U6737 ( .A1(n5577), .A2(n5586), .ZN(n5578) );
  OAI211_X1 U6738 ( .C1(n5581), .C2(n5580), .A(n5579), .B(n5578), .ZN(n6181)
         );
  AOI21_X1 U6739 ( .B1(n5583), .B2(n5582), .A(n6181), .ZN(n5592) );
  NAND2_X1 U6740 ( .A1(n5584), .A2(n6418), .ZN(n5591) );
  INV_X1 U6741 ( .A(n5585), .ZN(n5589) );
  NOR3_X1 U6742 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n6186), .A3(n5586), 
        .ZN(n5587) );
  AOI211_X1 U6743 ( .C1(n6412), .C2(n5589), .A(n5588), .B(n5587), .ZN(n5590)
         );
  OAI211_X1 U6744 ( .C1(n4306), .C2(n5592), .A(n5591), .B(n5590), .ZN(U3004)
         );
  XOR2_X1 U6745 ( .A(n5593), .B(n5530), .Z(n6122) );
  INV_X1 U6746 ( .A(n6122), .ZN(n6083) );
  INV_X1 U6747 ( .A(EBX_REG_20__SCAN_IN), .ZN(n5602) );
  INV_X1 U6748 ( .A(n5594), .ZN(n5595) );
  NAND2_X1 U6749 ( .A1(n5598), .A2(n5595), .ZN(n5596) );
  OAI21_X1 U6750 ( .B1(n5598), .B2(n5597), .A(n5596), .ZN(n5601) );
  INV_X1 U6751 ( .A(n5599), .ZN(n5600) );
  XNOR2_X1 U6752 ( .A(n5601), .B(n5600), .ZN(n5997) );
  INV_X1 U6753 ( .A(n5997), .ZN(n6081) );
  OAI222_X1 U6754 ( .A1(n6083), .A2(n5854), .B1(n6292), .B2(n5602), .C1(n6288), 
        .C2(n6081), .ZN(U2839) );
  NAND2_X1 U6755 ( .A1(n5605), .A2(n5606), .ZN(n5607) );
  AND2_X1 U6756 ( .A1(n5850), .A2(n5607), .ZN(n6119) );
  INV_X1 U6757 ( .A(n6119), .ZN(n5612) );
  INV_X1 U6758 ( .A(EBX_REG_21__SCAN_IN), .ZN(n5611) );
  OR2_X1 U6759 ( .A1(n5609), .A2(n5608), .ZN(n5610) );
  NAND2_X1 U6760 ( .A1(n4376), .A2(n5610), .ZN(n6075) );
  OAI222_X1 U6761 ( .A1(n5612), .A2(n5836), .B1(n5611), .B2(n6292), .C1(n6288), 
        .C2(n6075), .ZN(U2838) );
  INV_X1 U6762 ( .A(n6001), .ZN(n5615) );
  NOR2_X1 U6763 ( .A1(INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5977) );
  INV_X1 U6764 ( .A(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5968) );
  AND4_X1 U6765 ( .A1(n5977), .A2(n5968), .A3(n5994), .A4(n5613), .ZN(n5614)
         );
  NAND2_X1 U6766 ( .A1(n5615), .A2(n5614), .ZN(n5620) );
  NAND2_X1 U6767 ( .A1(n5616), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n6000) );
  NAND2_X1 U6768 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5627) );
  NOR2_X1 U6769 ( .A1(n5617), .A2(n5627), .ZN(n5634) );
  NAND2_X1 U6770 ( .A1(n5634), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5618) );
  NAND2_X1 U6771 ( .A1(n5620), .A2(n5619), .ZN(n5647) );
  XNOR2_X1 U6772 ( .A(n4294), .B(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n6128)
         );
  NAND2_X1 U6773 ( .A1(n5647), .A2(n6128), .ZN(n5705) );
  INV_X1 U6774 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n6155) );
  NAND2_X1 U6775 ( .A1(n4294), .A2(n6155), .ZN(n5621) );
  INV_X1 U6776 ( .A(n5646), .ZN(n5622) );
  NAND2_X1 U6777 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5943) );
  NOR2_X2 U6778 ( .A1(n5874), .A2(n5943), .ZN(n5864) );
  NOR2_X1 U6779 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5945) );
  NAND2_X1 U6780 ( .A1(n5945), .A2(n5879), .ZN(n5623) );
  NOR2_X1 U6781 ( .A1(n4294), .A2(n5623), .ZN(n5707) );
  NAND2_X1 U6782 ( .A1(n5646), .A2(n5707), .ZN(n5865) );
  NOR2_X1 U6783 ( .A1(n5865), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5624)
         );
  INV_X1 U6784 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5706) );
  XNOR2_X1 U6785 ( .A(n5625), .B(n5706), .ZN(n5645) );
  INV_X1 U6786 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5931) );
  INV_X1 U6787 ( .A(n5626), .ZN(n5628) );
  NAND2_X1 U6788 ( .A1(n5628), .A2(n5627), .ZN(n5629) );
  NAND2_X1 U6789 ( .A1(INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5959) );
  NAND2_X1 U6790 ( .A1(n5633), .A2(n5959), .ZN(n5631) );
  NAND2_X1 U6791 ( .A1(n5633), .A2(n5943), .ZN(n5632) );
  NAND2_X1 U6792 ( .A1(n5940), .A2(n5632), .ZN(n5937) );
  AOI21_X1 U6793 ( .B1(n5931), .B2(n5633), .A(n5937), .ZN(n5712) );
  INV_X1 U6794 ( .A(n5712), .ZN(n5638) );
  NAND2_X1 U6795 ( .A1(n5975), .A2(n5634), .ZN(n6149) );
  NOR2_X1 U6796 ( .A1(n5953), .A2(n5943), .ZN(n5932) );
  NAND3_X1 U6797 ( .A1(n5932), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .A3(n5706), .ZN(n5635) );
  NAND2_X1 U6798 ( .A1(n6371), .A2(REIP_REG_30__SCAN_IN), .ZN(n5640) );
  OAI211_X1 U6799 ( .C1(n6395), .C2(n5636), .A(n5635), .B(n5640), .ZN(n5637)
         );
  AOI21_X1 U6800 ( .B1(n5638), .B2(INSTADDRPOINTER_REG_30__SCAN_IN), .A(n5637), 
        .ZN(n5639) );
  OAI21_X1 U6801 ( .B1(n5645), .B2(n6398), .A(n5639), .ZN(U2988) );
  INV_X1 U6802 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5642) );
  NAND2_X1 U6803 ( .A1(n6144), .A2(n5759), .ZN(n5641) );
  OAI211_X1 U6804 ( .C1(n5642), .C2(n6148), .A(n5641), .B(n5640), .ZN(n5643)
         );
  AOI21_X1 U6805 ( .B1(n5855), .B2(n6357), .A(n5643), .ZN(n5644) );
  OAI21_X1 U6806 ( .B1(n5645), .B2(n6195), .A(n5644), .ZN(U2956) );
  NAND3_X1 U6807 ( .A1(n5622), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .A3(n4294), .ZN(n5648) );
  NOR2_X1 U6808 ( .A1(INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5960) );
  NAND3_X1 U6809 ( .A1(n5647), .A2(n6002), .A3(n5960), .ZN(n5873) );
  AOI22_X1 U6810 ( .A1(n5648), .A2(n5873), .B1(INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n5879), .ZN(n5649) );
  XNOR2_X1 U6811 ( .A(n5649), .B(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5949)
         );
  NAND2_X1 U6812 ( .A1(n6411), .A2(REIP_REG_28__SCAN_IN), .ZN(n5941) );
  OAI21_X1 U6813 ( .B1(n6148), .B2(n5650), .A(n5941), .ZN(n5655) );
  NOR2_X1 U6814 ( .A1(n5680), .A2(n5930), .ZN(n5654) );
  OAI21_X1 U6815 ( .B1(n6195), .B2(n5949), .A(n5656), .ZN(U2958) );
  AOI22_X1 U6816 ( .A1(n6487), .A2(n5658), .B1(n5657), .B2(n5665), .ZN(n6557)
         );
  INV_X1 U6817 ( .A(n6597), .ZN(n5660) );
  INV_X1 U6818 ( .A(n5738), .ZN(n6589) );
  AOI22_X1 U6819 ( .A1(n6589), .A2(n5665), .B1(STATE2_REG_1__SCAN_IN), .B2(
        n5736), .ZN(n5659) );
  OAI21_X1 U6820 ( .B1(n6557), .B2(n5660), .A(n5659), .ZN(n5662) );
  NOR2_X1 U6821 ( .A1(n5661), .A2(n5665), .ZN(n6559) );
  AOI22_X1 U6822 ( .A1(n5664), .A2(n5662), .B1(n6597), .B2(n6559), .ZN(n5663)
         );
  OAI21_X1 U6823 ( .B1(n5665), .B2(n5664), .A(n5663), .ZN(U3461) );
  AOI22_X1 U6824 ( .A1(n6296), .A2(DATAI_28_), .B1(n6299), .B2(
        EAX_REG_28__SCAN_IN), .ZN(n5667) );
  NAND2_X1 U6825 ( .A1(n6300), .A2(DATAI_12_), .ZN(n5666) );
  OAI211_X1 U6826 ( .C1(n5680), .C2(n6114), .A(n5667), .B(n5666), .ZN(U2863)
         );
  INV_X1 U6827 ( .A(n5827), .ZN(n5670) );
  INV_X1 U6828 ( .A(n5668), .ZN(n5669) );
  OAI21_X1 U6829 ( .B1(n5670), .B2(n5669), .A(n5774), .ZN(n5942) );
  INV_X1 U6830 ( .A(n5942), .ZN(n5671) );
  AOI22_X1 U6831 ( .A1(n5671), .A2(n5846), .B1(EBX_REG_28__SCAN_IN), .B2(n4405), .ZN(n5672) );
  OAI21_X1 U6832 ( .B1(n5680), .B2(n5854), .A(n5672), .ZN(U2831) );
  AOI22_X1 U6833 ( .A1(PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n6229), .B1(n6247), 
        .B2(n5673), .ZN(n5675) );
  NAND2_X1 U6834 ( .A1(n6276), .A2(EBX_REG_28__SCAN_IN), .ZN(n5674) );
  OAI211_X1 U6835 ( .C1(n6218), .C2(n5942), .A(n5675), .B(n5674), .ZN(n5677)
         );
  NOR3_X1 U6836 ( .A1(n6043), .A2(REIP_REG_28__SCAN_IN), .A3(n7009), .ZN(n5676) );
  AOI211_X1 U6837 ( .C1(REIP_REG_28__SCAN_IN), .C2(n5678), .A(n5677), .B(n5676), .ZN(n5679) );
  OAI21_X1 U6838 ( .B1(n5680), .B2(n6082), .A(n5679), .ZN(U2799) );
  CLKBUF_X1 U6839 ( .A(n5682), .Z(n5683) );
  OAI21_X1 U6840 ( .B1(n5681), .B2(n5684), .A(n5683), .ZN(n6346) );
  AOI221_X1 U6841 ( .B1(n5687), .B2(n5688), .C1(n5686), .C2(n5688), .A(n5685), 
        .ZN(n5692) );
  NAND4_X1 U6842 ( .A1(n6415), .A2(n6392), .A3(n6420), .A4(n5688), .ZN(n5690)
         );
  NAND2_X1 U6843 ( .A1(n6412), .A2(n6262), .ZN(n5689) );
  OAI211_X1 U6844 ( .C1(n6631), .C2(n6393), .A(n5690), .B(n5689), .ZN(n5691)
         );
  NOR2_X1 U6845 ( .A1(n5692), .A2(n5691), .ZN(n5693) );
  OAI21_X1 U6846 ( .B1(n6398), .B2(n6346), .A(n5693), .ZN(U3013) );
  AND2_X1 U6847 ( .A1(n5697), .A2(n5698), .ZN(n5699) );
  NOR2_X1 U6848 ( .A1(n5695), .A2(n5699), .ZN(n6109) );
  NAND2_X1 U6849 ( .A1(n6361), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5700)
         );
  OAI211_X1 U6850 ( .C1(n6370), .C2(n5810), .A(n5701), .B(n5700), .ZN(n5702)
         );
  AOI21_X1 U6851 ( .B1(n6109), .B2(n6357), .A(n5702), .ZN(n5703) );
  OAI21_X1 U6852 ( .B1(n5704), .B2(n6195), .A(n5703), .ZN(U2963) );
  NAND2_X1 U6853 ( .A1(n5864), .A2(n3181), .ZN(n5710) );
  INV_X1 U6855 ( .A(n6127), .ZN(n5708) );
  NAND4_X1 U6856 ( .A1(n5708), .A2(n5707), .A3(n5706), .A4(n5931), .ZN(n5709)
         );
  NAND2_X1 U6857 ( .A1(n5710), .A2(n5709), .ZN(n5711) );
  XNOR2_X1 U6858 ( .A(n5711), .B(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n5730)
         );
  OAI21_X1 U6859 ( .B1(INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n5713), .A(n5712), 
        .ZN(n5716) );
  NAND4_X1 U6860 ( .A1(n5932), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_30__SCAN_IN), .A4(n4434), .ZN(n5714) );
  NAND2_X1 U6861 ( .A1(n6411), .A2(REIP_REG_31__SCAN_IN), .ZN(n5726) );
  OAI21_X1 U6862 ( .B1(n5730), .B2(n6398), .A(n5719), .ZN(U2987) );
  INV_X1 U6863 ( .A(n5720), .ZN(n5724) );
  INV_X1 U6864 ( .A(n5721), .ZN(n6556) );
  AOI22_X1 U6865 ( .A1(n6556), .A2(n6597), .B1(n3989), .B2(n6589), .ZN(n5723)
         );
  NOR2_X1 U6866 ( .A1(n5743), .A2(n5722), .ZN(n5742) );
  OAI222_X1 U6867 ( .A1(n5738), .A2(n5724), .B1(n5743), .B2(n5723), .C1(n3165), 
        .C2(n5742), .ZN(U3456) );
  NAND2_X1 U6868 ( .A1(n6361), .A2(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n5725)
         );
  OAI211_X1 U6869 ( .C1(n6370), .C2(n5727), .A(n5726), .B(n5725), .ZN(n5728)
         );
  OAI21_X1 U6870 ( .B1(n5730), .B2(n6195), .A(n5729), .ZN(U2955) );
  NAND3_X1 U6871 ( .A1(n5732), .A2(n5731), .A3(n5860), .ZN(n5734) );
  AOI22_X1 U6872 ( .A1(n6296), .A2(DATAI_31_), .B1(EAX_REG_31__SCAN_IN), .B2(
        n6299), .ZN(n5733) );
  NAND2_X1 U6873 ( .A1(n5734), .A2(n5733), .ZN(U2860) );
  NOR3_X1 U6874 ( .A1(n6600), .A2(n5736), .A3(n5735), .ZN(n5740) );
  NOR3_X1 U6875 ( .A1(n5738), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n5737), 
        .ZN(n5739) );
  AOI211_X1 U6876 ( .C1(n6568), .C2(n6597), .A(n5740), .B(n5739), .ZN(n5744)
         );
  OAI22_X1 U6877 ( .A1(n5744), .A2(n5743), .B1(n5742), .B2(n5741), .ZN(U3459)
         );
  OAI22_X1 U6878 ( .A1(n5746), .A2(n6288), .B1(n6292), .B2(n5745), .ZN(U2828)
         );
  NAND2_X1 U6879 ( .A1(n4078), .A2(n5747), .ZN(n5751) );
  INV_X1 U6880 ( .A(n5754), .ZN(n5749) );
  OAI21_X1 U6881 ( .B1(n5749), .B2(n5748), .A(n5756), .ZN(n5750) );
  OAI211_X1 U6882 ( .C1(n5752), .C2(n5756), .A(n5751), .B(n5750), .ZN(n6575)
         );
  AND2_X1 U6883 ( .A1(n5754), .A2(n5753), .ZN(n5755) );
  AOI21_X1 U6884 ( .B1(n5756), .B2(n4030), .A(n5755), .ZN(n6188) );
  NAND2_X1 U6885 ( .A1(n5757), .A2(n6615), .ZN(n5758) );
  NAND2_X1 U6886 ( .A1(n5758), .A2(n7028), .ZN(n6677) );
  AND2_X1 U6887 ( .A1(n6188), .A2(n6677), .ZN(n6578) );
  NOR2_X1 U6888 ( .A1(n6578), .A2(n6598), .ZN(n6196) );
  MUX2_X1 U6889 ( .A(MORE_REG_SCAN_IN), .B(n6575), .S(n6196), .Z(U3471) );
  NAND2_X1 U6890 ( .A1(n5855), .A2(n6258), .ZN(n5768) );
  AOI22_X1 U6891 ( .A1(PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n6229), .B1(n6247), 
        .B2(n5759), .ZN(n5760) );
  OAI21_X1 U6892 ( .B1(n6242), .B2(n5761), .A(n5760), .ZN(n5765) );
  NOR3_X1 U6893 ( .A1(n5763), .A2(REIP_REG_30__SCAN_IN), .A3(n5762), .ZN(n5764) );
  AOI211_X1 U6894 ( .C1(n6277), .C2(n5766), .A(n5765), .B(n5764), .ZN(n5767)
         );
  OAI211_X1 U6895 ( .C1(n5782), .C2(n6975), .A(n5768), .B(n5767), .ZN(U2797)
         );
  INV_X1 U6896 ( .A(n5871), .ZN(n5819) );
  OAI22_X1 U6897 ( .A1(n5772), .A2(n6273), .B1(n6272), .B2(n5869), .ZN(n5781)
         );
  OAI211_X1 U6898 ( .C1(n5776), .C2(n5775), .A(n5774), .B(n5773), .ZN(n5777)
         );
  INV_X1 U6899 ( .A(n5777), .ZN(n5778) );
  NOR2_X1 U6900 ( .A1(n5935), .A2(n6218), .ZN(n5780) );
  AOI211_X1 U6901 ( .C1(n6276), .C2(EBX_REG_29__SCAN_IN), .A(n5781), .B(n5780), 
        .ZN(n5786) );
  INV_X1 U6902 ( .A(n5782), .ZN(n5783) );
  OAI21_X1 U6903 ( .B1(REIP_REG_29__SCAN_IN), .B2(n5784), .A(n5783), .ZN(n5785) );
  OAI211_X1 U6904 ( .C1(n5819), .C2(n6082), .A(n5786), .B(n5785), .ZN(U2798)
         );
  INV_X1 U6905 ( .A(n5787), .ZN(n5793) );
  INV_X1 U6906 ( .A(n5789), .ZN(n5792) );
  INV_X1 U6907 ( .A(n5791), .ZN(n5829) );
  NAND2_X1 U6908 ( .A1(REIP_REG_24__SCAN_IN), .A2(n5798), .ZN(n6045) );
  OAI22_X1 U6909 ( .A1(REIP_REG_25__SCAN_IN), .A2(n6045), .B1(n6132), .B2(
        n6272), .ZN(n5806) );
  INV_X1 U6910 ( .A(n5843), .ZN(n5795) );
  AOI21_X1 U6911 ( .B1(n5795), .B2(n5842), .A(n5794), .ZN(n5796) );
  OR2_X1 U6912 ( .A1(n5796), .A2(n5831), .ZN(n5837) );
  NOR2_X1 U6913 ( .A1(n6091), .A2(n5797), .ZN(n6055) );
  INV_X1 U6914 ( .A(REIP_REG_24__SCAN_IN), .ZN(n6962) );
  NAND2_X1 U6915 ( .A1(n6962), .A2(n5798), .ZN(n6057) );
  INV_X1 U6916 ( .A(n6057), .ZN(n5799) );
  OAI21_X1 U6917 ( .B1(n6055), .B2(n5799), .A(REIP_REG_25__SCAN_IN), .ZN(n5804) );
  OAI22_X1 U6918 ( .A1(n5801), .A2(n6242), .B1(n5800), .B2(n6273), .ZN(n5802)
         );
  INV_X1 U6919 ( .A(n5802), .ZN(n5803) );
  OAI211_X1 U6920 ( .C1(n6218), .C2(n5837), .A(n5804), .B(n5803), .ZN(n5805)
         );
  AOI211_X1 U6921 ( .C1(n6129), .C2(n6258), .A(n5806), .B(n5805), .ZN(n5807)
         );
  INV_X1 U6922 ( .A(n5807), .ZN(U2802) );
  INV_X1 U6923 ( .A(n6109), .ZN(n5848) );
  INV_X1 U6924 ( .A(n5808), .ZN(n5845) );
  NAND2_X1 U6925 ( .A1(n6229), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5815)
         );
  NAND2_X1 U6926 ( .A1(n7027), .A2(n5809), .ZN(n5813) );
  OAI22_X1 U6927 ( .A1(n5811), .A2(n6242), .B1(n5810), .B2(n6272), .ZN(n5812)
         );
  AOI21_X1 U6928 ( .B1(n5813), .B2(n6055), .A(n5812), .ZN(n5814) );
  NAND2_X1 U6929 ( .A1(n5815), .A2(n5814), .ZN(n5816) );
  AOI21_X1 U6930 ( .B1(n5845), .B2(n6277), .A(n5816), .ZN(n5817) );
  OAI21_X1 U6931 ( .B1(n5848), .B2(n6082), .A(n5817), .ZN(U2804) );
  OAI222_X1 U6932 ( .A1(n5854), .A2(n5819), .B1(n5818), .B2(n6292), .C1(n5935), 
        .C2(n6288), .ZN(U2830) );
  AND2_X1 U6933 ( .A1(n5821), .A2(n5822), .ZN(n5824) );
  INV_X1 U6934 ( .A(EBX_REG_27__SCAN_IN), .ZN(n5828) );
  OR2_X1 U6935 ( .A1(n5833), .A2(n5825), .ZN(n5826) );
  NAND2_X1 U6936 ( .A1(n5827), .A2(n5826), .ZN(n6038) );
  OAI222_X1 U6937 ( .A1(n5836), .A2(n6039), .B1(n5828), .B2(n6292), .C1(n6038), 
        .C2(n6288), .ZN(U2832) );
  NOR2_X1 U6938 ( .A1(n5831), .A2(n5830), .ZN(n5832) );
  OR2_X1 U6939 ( .A1(n5833), .A2(n5832), .ZN(n6046) );
  INV_X1 U6940 ( .A(n6046), .ZN(n5834) );
  AOI22_X1 U6941 ( .A1(n5846), .A2(n5834), .B1(EBX_REG_26__SCAN_IN), .B2(n4405), .ZN(n5835) );
  OAI21_X1 U6942 ( .B1(n6047), .B2(n5836), .A(n5835), .ZN(U2833) );
  INV_X1 U6943 ( .A(n6129), .ZN(n5839) );
  INV_X1 U6944 ( .A(n5837), .ZN(n6151) );
  AOI22_X1 U6945 ( .A1(n5846), .A2(n6151), .B1(EBX_REG_25__SCAN_IN), .B2(n4405), .ZN(n5838) );
  OAI21_X1 U6946 ( .B1(n5839), .B2(n5854), .A(n5838), .ZN(U2834) );
  NOR2_X1 U6947 ( .A1(n5695), .A2(n5840), .ZN(n5841) );
  OR2_X1 U6948 ( .A1(n5789), .A2(n5841), .ZN(n5890) );
  XNOR2_X1 U6949 ( .A(n5843), .B(n5842), .ZN(n6056) );
  AOI22_X1 U6950 ( .A1(n5846), .A2(n6056), .B1(EBX_REG_24__SCAN_IN), .B2(n4405), .ZN(n5844) );
  OAI21_X1 U6951 ( .B1(n5890), .B2(n5854), .A(n5844), .ZN(U2835) );
  AOI22_X1 U6952 ( .A1(n5846), .A2(n5845), .B1(EBX_REG_23__SCAN_IN), .B2(n4405), .ZN(n5847) );
  OAI21_X1 U6953 ( .B1(n5848), .B2(n5854), .A(n5847), .ZN(U2836) );
  NAND2_X1 U6954 ( .A1(n5850), .A2(n5849), .ZN(n5851) );
  NAND2_X1 U6955 ( .A1(n5697), .A2(n5851), .ZN(n6115) );
  XNOR2_X1 U6956 ( .A(n4376), .B(n5852), .ZN(n6064) );
  INV_X1 U6957 ( .A(EBX_REG_22__SCAN_IN), .ZN(n5853) );
  OAI222_X1 U6958 ( .A1(n5854), .A2(n6115), .B1(n6288), .B2(n6064), .C1(n5853), 
        .C2(n6292), .ZN(U2837) );
  NAND2_X1 U6959 ( .A1(n5855), .A2(n6297), .ZN(n5857) );
  AOI22_X1 U6960 ( .A1(n6296), .A2(DATAI_30_), .B1(n6299), .B2(
        EAX_REG_30__SCAN_IN), .ZN(n5856) );
  OAI211_X1 U6961 ( .C1(n5861), .C2(n5345), .A(n5857), .B(n5856), .ZN(U2861)
         );
  NAND2_X1 U6962 ( .A1(n5871), .A2(n6297), .ZN(n5859) );
  AOI22_X1 U6963 ( .A1(n6296), .A2(DATAI_29_), .B1(n6299), .B2(
        EAX_REG_29__SCAN_IN), .ZN(n5858) );
  OAI211_X1 U6964 ( .C1(n5861), .C2(n6848), .A(n5859), .B(n5858), .ZN(U2862)
         );
  OAI22_X1 U6965 ( .A1(n5861), .A2(n5330), .B1(n4469), .B2(n5860), .ZN(n5862)
         );
  AOI21_X1 U6966 ( .B1(n6296), .B2(DATAI_26_), .A(n5862), .ZN(n5863) );
  OAI21_X1 U6967 ( .B1(n6047), .B2(n6114), .A(n5863), .ZN(U2865) );
  INV_X1 U6968 ( .A(n5864), .ZN(n5866) );
  NAND2_X1 U6969 ( .A1(n5866), .A2(n5865), .ZN(n5867) );
  XNOR2_X1 U6970 ( .A(n5867), .B(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5939)
         );
  NAND2_X1 U6971 ( .A1(n6371), .A2(REIP_REG_29__SCAN_IN), .ZN(n5933) );
  NAND2_X1 U6972 ( .A1(n6361), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5868)
         );
  OAI211_X1 U6973 ( .C1(n6370), .C2(n5869), .A(n5933), .B(n5868), .ZN(n5870)
         );
  AOI21_X1 U6974 ( .B1(n5871), .B2(n6357), .A(n5870), .ZN(n5872) );
  OAI21_X1 U6975 ( .B1(n5939), .B2(n6195), .A(n5872), .ZN(U2957) );
  NAND2_X1 U6976 ( .A1(n5874), .A2(n5873), .ZN(n5875) );
  XNOR2_X1 U6977 ( .A(n5875), .B(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5957)
         );
  NOR2_X1 U6978 ( .A1(n6393), .A2(n7009), .ZN(n5950) );
  AOI21_X1 U6979 ( .B1(n6361), .B2(PHYADDRPOINTER_REG_27__SCAN_IN), .A(n5950), 
        .ZN(n5876) );
  OAI21_X1 U6980 ( .B1(n6036), .B2(n6370), .A(n5876), .ZN(n5877) );
  AOI21_X1 U6981 ( .B1(n6101), .B2(n6357), .A(n5877), .ZN(n5878) );
  OAI21_X1 U6982 ( .B1(n5957), .B2(n6195), .A(n5878), .ZN(U2959) );
  XNOR2_X1 U6983 ( .A(n4294), .B(n5879), .ZN(n5880) );
  XNOR2_X1 U6984 ( .A(n5881), .B(n5880), .ZN(n5966) );
  NAND2_X1 U6985 ( .A1(n6411), .A2(REIP_REG_26__SCAN_IN), .ZN(n5958) );
  OAI21_X1 U6986 ( .B1(n6148), .B2(n5882), .A(n5958), .ZN(n5884) );
  NOR2_X1 U6987 ( .A1(n6047), .A2(n5930), .ZN(n5883) );
  AOI211_X1 U6988 ( .C1(n6144), .C2(n6044), .A(n5884), .B(n5883), .ZN(n5885)
         );
  OAI21_X1 U6989 ( .B1(n6195), .B2(n5966), .A(n5885), .ZN(U2960) );
  INV_X1 U6990 ( .A(n5902), .ZN(n5886) );
  OAI21_X1 U6991 ( .B1(n6002), .B2(INSTADDRPOINTER_REG_21__SCAN_IN), .A(n5886), 
        .ZN(n5897) );
  NAND3_X1 U6992 ( .A1(n4294), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5887) );
  OAI22_X1 U6993 ( .A1(n5888), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .B1(n5897), .B2(n5887), .ZN(n5889) );
  XNOR2_X1 U6994 ( .A(n5889), .B(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5972)
         );
  INV_X1 U6995 ( .A(n6054), .ZN(n5892) );
  AND2_X1 U6996 ( .A1(n6411), .A2(REIP_REG_24__SCAN_IN), .ZN(n5970) );
  AOI21_X1 U6997 ( .B1(n6361), .B2(PHYADDRPOINTER_REG_24__SCAN_IN), .A(n5970), 
        .ZN(n5891) );
  OAI21_X1 U6998 ( .B1(n5892), .B2(n6370), .A(n5891), .ZN(n5893) );
  AOI21_X1 U6999 ( .B1(n6106), .B2(n6357), .A(n5893), .ZN(n5894) );
  OAI21_X1 U7000 ( .B1(n5972), .B2(n6195), .A(n5894), .ZN(U2962) );
  AOI21_X1 U7001 ( .B1(INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n4294), .A(n5895), 
        .ZN(n5896) );
  XNOR2_X1 U7002 ( .A(n5897), .B(n5896), .ZN(n5981) );
  NAND2_X1 U7003 ( .A1(n6411), .A2(REIP_REG_22__SCAN_IN), .ZN(n5974) );
  OAI21_X1 U7004 ( .B1(n6148), .B2(n5898), .A(n5974), .ZN(n5900) );
  NOR2_X1 U7005 ( .A1(n6115), .A2(n5930), .ZN(n5899) );
  AOI211_X1 U7006 ( .C1(n6144), .C2(n6063), .A(n5900), .B(n5899), .ZN(n5901)
         );
  OAI21_X1 U7007 ( .B1(n5981), .B2(n6195), .A(n5901), .ZN(U2964) );
  AOI21_X1 U7008 ( .B1(n5904), .B2(n5903), .A(n5902), .ZN(n5988) );
  NAND2_X1 U7009 ( .A1(n6411), .A2(REIP_REG_21__SCAN_IN), .ZN(n5982) );
  NAND2_X1 U7010 ( .A1(n6361), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n5905)
         );
  OAI211_X1 U7011 ( .C1(n6370), .C2(n6072), .A(n5982), .B(n5905), .ZN(n5906)
         );
  AOI21_X1 U7012 ( .B1(n6119), .B2(n6357), .A(n5906), .ZN(n5907) );
  OAI21_X1 U7013 ( .B1(n5988), .B2(n6195), .A(n5907), .ZN(U2965) );
  XNOR2_X1 U7014 ( .A(n5909), .B(n5908), .ZN(n5999) );
  NAND2_X1 U7015 ( .A1(n6144), .A2(n6079), .ZN(n5910) );
  NAND2_X1 U7016 ( .A1(n6411), .A2(REIP_REG_20__SCAN_IN), .ZN(n5989) );
  OAI211_X1 U7017 ( .C1(n6148), .C2(n6089), .A(n5910), .B(n5989), .ZN(n5911)
         );
  AOI21_X1 U7018 ( .B1(n6122), .B2(n6357), .A(n5911), .ZN(n5912) );
  OAI21_X1 U7019 ( .B1(n5999), .B2(n6195), .A(n5912), .ZN(U2966) );
  NAND2_X1 U7020 ( .A1(n6371), .A2(REIP_REG_18__SCAN_IN), .ZN(n6015) );
  NOR2_X1 U7021 ( .A1(n4294), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5915)
         );
  NAND2_X1 U7022 ( .A1(n5914), .A2(n5915), .ZN(n6140) );
  NAND3_X1 U7023 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n4294), .A3(n5922), .ZN(n5916) );
  OAI22_X1 U7024 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n6140), .B1(n5916), .B2(n5914), .ZN(n5917) );
  XNOR2_X1 U7025 ( .A(n6019), .B(n5917), .ZN(n6017) );
  NAND2_X1 U7026 ( .A1(n6366), .A2(n6017), .ZN(n5918) );
  OAI211_X1 U7027 ( .C1(n6148), .C2(n6212), .A(n6015), .B(n5918), .ZN(n5919)
         );
  AOI21_X1 U7028 ( .B1(n6144), .B2(n6214), .A(n5919), .ZN(n5920) );
  OAI21_X1 U7029 ( .B1(n5921), .B2(n5930), .A(n5920), .ZN(U2968) );
  OAI21_X1 U7030 ( .B1(n4294), .B2(n5923), .A(n5922), .ZN(n5924) );
  XOR2_X1 U7031 ( .A(n5924), .B(n5914), .Z(n6174) );
  NAND2_X1 U7032 ( .A1(n6174), .A2(n6366), .ZN(n5928) );
  AND2_X1 U7033 ( .A1(n6411), .A2(REIP_REG_16__SCAN_IN), .ZN(n6171) );
  NOR2_X1 U7034 ( .A1(n6370), .A2(n5925), .ZN(n5926) );
  AOI211_X1 U7035 ( .C1(n6361), .C2(PHYADDRPOINTER_REG_16__SCAN_IN), .A(n6171), 
        .B(n5926), .ZN(n5927) );
  OAI211_X1 U7036 ( .C1(n5930), .C2(n5929), .A(n5928), .B(n5927), .ZN(U2970)
         );
  NAND2_X1 U7037 ( .A1(n5932), .A2(n5931), .ZN(n5934) );
  OAI211_X1 U7038 ( .C1(n6395), .C2(n5935), .A(n5934), .B(n5933), .ZN(n5936)
         );
  AOI21_X1 U7039 ( .B1(INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n5937), .A(n5936), 
        .ZN(n5938) );
  OAI21_X1 U7040 ( .B1(n5939), .B2(n6398), .A(n5938), .ZN(U2989) );
  INV_X1 U7041 ( .A(n5940), .ZN(n5955) );
  OAI21_X1 U7042 ( .B1(n5942), .B2(n6395), .A(n5941), .ZN(n5947) );
  INV_X1 U7043 ( .A(n5943), .ZN(n5944) );
  NOR3_X1 U7044 ( .A1(n5953), .A2(n5945), .A3(n5944), .ZN(n5946) );
  AOI211_X1 U7045 ( .C1(INSTADDRPOINTER_REG_28__SCAN_IN), .C2(n5955), .A(n5947), .B(n5946), .ZN(n5948) );
  OAI21_X1 U7046 ( .B1(n5949), .B2(n6398), .A(n5948), .ZN(U2990) );
  INV_X1 U7047 ( .A(n6038), .ZN(n5951) );
  AOI21_X1 U7048 ( .B1(n6412), .B2(n5951), .A(n5950), .ZN(n5952) );
  OAI21_X1 U7049 ( .B1(n5953), .B2(INSTADDRPOINTER_REG_27__SCAN_IN), .A(n5952), 
        .ZN(n5954) );
  AOI21_X1 U7050 ( .B1(n5955), .B2(INSTADDRPOINTER_REG_27__SCAN_IN), .A(n5954), 
        .ZN(n5956) );
  OAI21_X1 U7051 ( .B1(n5957), .B2(n6398), .A(n5956), .ZN(U2991) );
  INV_X1 U7052 ( .A(n6156), .ZN(n5964) );
  OAI21_X1 U7053 ( .B1(n6395), .B2(n6046), .A(n5958), .ZN(n5963) );
  INV_X1 U7054 ( .A(n5959), .ZN(n5961) );
  NOR3_X1 U7055 ( .A1(n6149), .A2(n5961), .A3(n5960), .ZN(n5962) );
  AOI211_X1 U7056 ( .C1(INSTADDRPOINTER_REG_26__SCAN_IN), .C2(n5964), .A(n5963), .B(n5962), .ZN(n5965) );
  OAI21_X1 U7057 ( .B1(n5966), .B2(n6398), .A(n5965), .ZN(U2992) );
  NAND3_X1 U7058 ( .A1(n5975), .A2(n5976), .A3(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5967) );
  AOI21_X1 U7059 ( .B1(n5968), .B2(n5967), .A(n6156), .ZN(n5969) );
  AOI211_X1 U7060 ( .C1(n6412), .C2(n6056), .A(n5970), .B(n5969), .ZN(n5971)
         );
  OAI21_X1 U7061 ( .B1(n5972), .B2(n6398), .A(n5971), .ZN(U2994) );
  INV_X1 U7062 ( .A(n5973), .ZN(n5986) );
  OAI21_X1 U7063 ( .B1(n6395), .B2(n6064), .A(n5974), .ZN(n5979) );
  INV_X1 U7064 ( .A(n5975), .ZN(n5983) );
  NOR3_X1 U7065 ( .A1(n5983), .A2(n5977), .A3(n5976), .ZN(n5978) );
  AOI211_X1 U7066 ( .C1(n5986), .C2(INSTADDRPOINTER_REG_22__SCAN_IN), .A(n5979), .B(n5978), .ZN(n5980) );
  OAI21_X1 U7067 ( .B1(n5981), .B2(n6398), .A(n5980), .ZN(U2996) );
  OAI21_X1 U7068 ( .B1(n6395), .B2(n6075), .A(n5982), .ZN(n5985) );
  NOR2_X1 U7069 ( .A1(n5983), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5984)
         );
  AOI211_X1 U7070 ( .C1(n5986), .C2(INSTADDRPOINTER_REG_21__SCAN_IN), .A(n5985), .B(n5984), .ZN(n5987) );
  OAI21_X1 U7071 ( .B1(n5988), .B2(n6398), .A(n5987), .ZN(U2997) );
  NAND4_X1 U7072 ( .A1(n5994), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_19__SCAN_IN), .A4(n6375), .ZN(n5990) );
  OAI21_X1 U7073 ( .B1(n5991), .B2(n5990), .A(n5989), .ZN(n5996) );
  OR2_X1 U7074 ( .A1(n6159), .A2(n6019), .ZN(n5993) );
  NAND2_X1 U7075 ( .A1(n5993), .A2(n5992), .ZN(n6005) );
  NAND4_X1 U7076 ( .A1(n6012), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .A3(n6004), .A4(n6375), .ZN(n6006) );
  AOI21_X1 U7077 ( .B1(n6005), .B2(n6006), .A(n5994), .ZN(n5995) );
  AOI211_X1 U7078 ( .C1(n6412), .C2(n5997), .A(n5996), .B(n5995), .ZN(n5998)
         );
  OAI21_X1 U7079 ( .B1(n5999), .B2(n6398), .A(n5998), .ZN(U2998) );
  NAND2_X1 U7080 ( .A1(n6001), .A2(n6000), .ZN(n6003) );
  XNOR2_X1 U7081 ( .A(n6003), .B(n6002), .ZN(n6134) );
  NOR2_X1 U7082 ( .A1(n6005), .A2(n6004), .ZN(n6010) );
  NAND2_X1 U7083 ( .A1(n6371), .A2(REIP_REG_19__SCAN_IN), .ZN(n6007) );
  OAI211_X1 U7084 ( .C1(n6395), .C2(n6008), .A(n6007), .B(n6006), .ZN(n6009)
         );
  AOI211_X1 U7085 ( .C1(n6134), .C2(n6418), .A(n6010), .B(n6009), .ZN(n6011)
         );
  INV_X1 U7086 ( .A(n6011), .ZN(U2999) );
  INV_X1 U7087 ( .A(n6159), .ZN(n6020) );
  AND2_X1 U7088 ( .A1(n6375), .A2(n6012), .ZN(n6013) );
  NAND2_X1 U7089 ( .A1(n6019), .A2(n6013), .ZN(n6014) );
  OAI211_X1 U7090 ( .C1(n6395), .C2(n6217), .A(n6015), .B(n6014), .ZN(n6016)
         );
  AOI21_X1 U7091 ( .B1(n6418), .B2(n6017), .A(n6016), .ZN(n6018) );
  OAI21_X1 U7092 ( .B1(n6020), .B2(n6019), .A(n6018), .ZN(U3000) );
  OAI211_X1 U7093 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n4652), .A(n6485), .B(
        n6484), .ZN(n6022) );
  OAI21_X1 U7094 ( .B1(n6032), .B2(n6023), .A(n6022), .ZN(n6024) );
  MUX2_X1 U7095 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n6024), .S(n6425), 
        .Z(U3464) );
  XNOR2_X1 U7096 ( .A(n6485), .B(n6025), .ZN(n6026) );
  OAI22_X1 U7097 ( .A1(n6026), .A2(n6498), .B1(n4527), .B2(n6032), .ZN(n6027)
         );
  MUX2_X1 U7098 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n6027), .S(n6425), 
        .Z(U3463) );
  INV_X1 U7099 ( .A(n6028), .ZN(n6029) );
  NOR2_X1 U7100 ( .A1(n6029), .A2(n6485), .ZN(n6444) );
  NOR2_X1 U7101 ( .A1(n6030), .A2(n6444), .ZN(n6031) );
  OAI222_X1 U7102 ( .A1(n4246), .A2(n6033), .B1(n6281), .B2(n6032), .C1(n6498), 
        .C2(n6031), .ZN(n6034) );
  MUX2_X1 U7103 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B(n6034), .S(n6425), 
        .Z(U3462) );
  AND2_X1 U7104 ( .A1(n6323), .A2(DATAO_REG_31__SCAN_IN), .ZN(U2892) );
  AOI22_X1 U7105 ( .A1(EBX_REG_27__SCAN_IN), .A2(n6276), .B1(
        PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n6229), .ZN(n6035) );
  OAI21_X1 U7106 ( .B1(n6036), .B2(n6272), .A(n6035), .ZN(n6037) );
  AOI21_X1 U7107 ( .B1(REIP_REG_27__SCAN_IN), .B2(n6050), .A(n6037), .ZN(n6042) );
  OAI22_X1 U7108 ( .A1(n6039), .A2(n6082), .B1(n6038), .B2(n6218), .ZN(n6040)
         );
  INV_X1 U7109 ( .A(n6040), .ZN(n6041) );
  OAI211_X1 U7110 ( .C1(REIP_REG_27__SCAN_IN), .C2(n6043), .A(n6042), .B(n6041), .ZN(U2800) );
  AOI22_X1 U7111 ( .A1(PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n6229), .B1(n6044), 
        .B2(n6247), .ZN(n6052) );
  INV_X1 U7112 ( .A(REIP_REG_25__SCAN_IN), .ZN(n6652) );
  INV_X1 U7113 ( .A(REIP_REG_26__SCAN_IN), .ZN(n6957) );
  OAI21_X1 U7114 ( .B1(n6652), .B2(n6045), .A(n6957), .ZN(n6049) );
  OAI22_X1 U7115 ( .A1(n6047), .A2(n6082), .B1(n6046), .B2(n6218), .ZN(n6048)
         );
  AOI21_X1 U7116 ( .B1(n6050), .B2(n6049), .A(n6048), .ZN(n6051) );
  OAI211_X1 U7117 ( .C1(n6053), .C2(n6242), .A(n6052), .B(n6051), .ZN(U2801)
         );
  AOI22_X1 U7118 ( .A1(EBX_REG_24__SCAN_IN), .A2(n6276), .B1(
        PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n6229), .ZN(n6060) );
  AOI22_X1 U7119 ( .A1(REIP_REG_24__SCAN_IN), .A2(n6055), .B1(n6054), .B2(
        n6247), .ZN(n6059) );
  AOI22_X1 U7120 ( .A1(n6106), .A2(n6258), .B1(n6277), .B2(n6056), .ZN(n6058)
         );
  NAND4_X1 U7121 ( .A1(n6060), .A2(n6059), .A3(n6058), .A4(n6057), .ZN(U2803)
         );
  AOI22_X1 U7122 ( .A1(EBX_REG_22__SCAN_IN), .A2(n6276), .B1(
        PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n6229), .ZN(n6070) );
  INV_X1 U7123 ( .A(n6061), .ZN(n6062) );
  NOR2_X1 U7124 ( .A1(n6091), .A2(n6062), .ZN(n6086) );
  AOI22_X1 U7125 ( .A1(n6063), .A2(n6247), .B1(REIP_REG_22__SCAN_IN), .B2(
        n6086), .ZN(n6069) );
  OAI22_X1 U7126 ( .A1(n6115), .A2(n6082), .B1(n6064), .B2(n6218), .ZN(n6065)
         );
  INV_X1 U7127 ( .A(n6065), .ZN(n6068) );
  OAI211_X1 U7128 ( .C1(REIP_REG_22__SCAN_IN), .C2(REIP_REG_21__SCAN_IN), .A(
        n6074), .B(n6066), .ZN(n6067) );
  NAND4_X1 U7129 ( .A1(n6070), .A2(n6069), .A3(n6068), .A4(n6067), .ZN(U2805)
         );
  INV_X1 U7130 ( .A(REIP_REG_21__SCAN_IN), .ZN(n6649) );
  AOI22_X1 U7131 ( .A1(EBX_REG_21__SCAN_IN), .A2(n6276), .B1(
        PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n6229), .ZN(n6071) );
  OAI21_X1 U7132 ( .B1(n6072), .B2(n6272), .A(n6071), .ZN(n6073) );
  AOI221_X1 U7133 ( .B1(n6086), .B2(REIP_REG_21__SCAN_IN), .C1(n6074), .C2(
        n6649), .A(n6073), .ZN(n6078) );
  INV_X1 U7134 ( .A(n6075), .ZN(n6076) );
  AOI22_X1 U7135 ( .A1(n6119), .A2(n6258), .B1(n6277), .B2(n6076), .ZN(n6077)
         );
  NAND2_X1 U7136 ( .A1(n6078), .A2(n6077), .ZN(U2806) );
  AOI22_X1 U7137 ( .A1(EBX_REG_20__SCAN_IN), .A2(n6276), .B1(n6079), .B2(n6247), .ZN(n6088) );
  NAND2_X1 U7138 ( .A1(n6080), .A2(n6773), .ZN(n6085) );
  OAI22_X1 U7139 ( .A1(n6083), .A2(n6082), .B1(n6081), .B2(n6218), .ZN(n6084)
         );
  AOI21_X1 U7140 ( .B1(n6086), .B2(n6085), .A(n6084), .ZN(n6087) );
  OAI211_X1 U7141 ( .C1(n6089), .C2(n6273), .A(n6088), .B(n6087), .ZN(U2807)
         );
  NOR2_X1 U7142 ( .A1(n6091), .A2(n6090), .ZN(n6223) );
  INV_X1 U7143 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n6094) );
  NAND2_X1 U7144 ( .A1(REIP_REG_18__SCAN_IN), .A2(REIP_REG_19__SCAN_IN), .ZN(
        n6092) );
  OAI211_X1 U7145 ( .C1(REIP_REG_18__SCAN_IN), .C2(REIP_REG_19__SCAN_IN), .A(
        n6210), .B(n6092), .ZN(n6093) );
  OAI211_X1 U7146 ( .C1(n6273), .C2(n6094), .A(n6093), .B(n6393), .ZN(n6095)
         );
  AOI21_X1 U7147 ( .B1(REIP_REG_19__SCAN_IN), .B2(n6223), .A(n6095), .ZN(n6099) );
  AOI222_X1 U7148 ( .A1(n6097), .A2(n6277), .B1(n6258), .B2(n6133), .C1(n6096), 
        .C2(n6247), .ZN(n6098) );
  OAI211_X1 U7149 ( .C1(n6100), .C2(n6242), .A(n6099), .B(n6098), .ZN(U2808)
         );
  AOI22_X1 U7150 ( .A1(n6101), .A2(n6297), .B1(n6296), .B2(DATAI_27_), .ZN(
        n6103) );
  AOI22_X1 U7151 ( .A1(n6300), .A2(DATAI_11_), .B1(EAX_REG_27__SCAN_IN), .B2(
        n6299), .ZN(n6102) );
  NAND2_X1 U7152 ( .A1(n6103), .A2(n6102), .ZN(U2864) );
  AOI22_X1 U7153 ( .A1(n6129), .A2(n6297), .B1(n6296), .B2(DATAI_25_), .ZN(
        n6105) );
  AOI22_X1 U7154 ( .A1(n6300), .A2(DATAI_9_), .B1(EAX_REG_25__SCAN_IN), .B2(
        n6299), .ZN(n6104) );
  NAND2_X1 U7155 ( .A1(n6105), .A2(n6104), .ZN(U2866) );
  AOI22_X1 U7156 ( .A1(n6106), .A2(n6297), .B1(n6296), .B2(DATAI_24_), .ZN(
        n6108) );
  AOI22_X1 U7157 ( .A1(n6300), .A2(DATAI_8_), .B1(EAX_REG_24__SCAN_IN), .B2(
        n6299), .ZN(n6107) );
  NAND2_X1 U7158 ( .A1(n6108), .A2(n6107), .ZN(U2867) );
  AOI22_X1 U7159 ( .A1(n6109), .A2(n6297), .B1(n6296), .B2(DATAI_23_), .ZN(
        n6111) );
  AOI22_X1 U7160 ( .A1(n6300), .A2(DATAI_7_), .B1(EAX_REG_23__SCAN_IN), .B2(
        n6299), .ZN(n6110) );
  NAND2_X1 U7161 ( .A1(n6111), .A2(n6110), .ZN(U2868) );
  INV_X1 U7162 ( .A(n6296), .ZN(n6113) );
  INV_X1 U7163 ( .A(DATAI_22_), .ZN(n6112) );
  OAI22_X1 U7164 ( .A1(n6115), .A2(n6114), .B1(n6113), .B2(n6112), .ZN(n6116)
         );
  INV_X1 U7165 ( .A(n6116), .ZN(n6118) );
  AOI22_X1 U7166 ( .A1(n6300), .A2(DATAI_6_), .B1(EAX_REG_22__SCAN_IN), .B2(
        n6299), .ZN(n6117) );
  NAND2_X1 U7167 ( .A1(n6118), .A2(n6117), .ZN(U2869) );
  AOI22_X1 U7168 ( .A1(n6119), .A2(n6297), .B1(n6296), .B2(DATAI_21_), .ZN(
        n6121) );
  AOI22_X1 U7169 ( .A1(n6300), .A2(DATAI_5_), .B1(EAX_REG_21__SCAN_IN), .B2(
        n6299), .ZN(n6120) );
  NAND2_X1 U7170 ( .A1(n6121), .A2(n6120), .ZN(U2870) );
  AOI22_X1 U7171 ( .A1(n6122), .A2(n6297), .B1(n6296), .B2(DATAI_20_), .ZN(
        n6124) );
  AOI22_X1 U7172 ( .A1(n6300), .A2(DATAI_4_), .B1(EAX_REG_20__SCAN_IN), .B2(
        n6299), .ZN(n6123) );
  NAND2_X1 U7173 ( .A1(n6124), .A2(n6123), .ZN(U2871) );
  AOI22_X1 U7174 ( .A1(n6133), .A2(n6297), .B1(n6296), .B2(DATAI_19_), .ZN(
        n6126) );
  AOI22_X1 U7175 ( .A1(n6300), .A2(DATAI_3_), .B1(EAX_REG_19__SCAN_IN), .B2(
        n6299), .ZN(n6125) );
  NAND2_X1 U7176 ( .A1(n6126), .A2(n6125), .ZN(U2872) );
  AOI22_X1 U7177 ( .A1(n6411), .A2(REIP_REG_25__SCAN_IN), .B1(n6361), .B2(
        PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n6131) );
  OAI21_X1 U7178 ( .B1(n5647), .B2(n6128), .A(n6127), .ZN(n6152) );
  AOI22_X1 U7179 ( .A1(n6129), .A2(n6357), .B1(n6366), .B2(n6152), .ZN(n6130)
         );
  OAI211_X1 U7180 ( .C1(n6370), .C2(n6132), .A(n6131), .B(n6130), .ZN(U2961)
         );
  AOI22_X1 U7181 ( .A1(n6371), .A2(REIP_REG_19__SCAN_IN), .B1(n6361), .B2(
        PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n6136) );
  AOI22_X1 U7182 ( .A1(n6134), .A2(n6366), .B1(n6357), .B2(n6133), .ZN(n6135)
         );
  OAI211_X1 U7183 ( .C1(n6370), .C2(n6137), .A(n6136), .B(n6135), .ZN(U2967)
         );
  INV_X1 U7184 ( .A(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n6220) );
  NAND2_X1 U7185 ( .A1(n4294), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n6138) );
  OR2_X1 U7186 ( .A1(n5914), .A2(n6138), .ZN(n6139) );
  NAND2_X1 U7187 ( .A1(n6140), .A2(n6139), .ZN(n6141) );
  XNOR2_X1 U7188 ( .A(n6141), .B(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n6168)
         );
  INV_X1 U7189 ( .A(n6168), .ZN(n6146) );
  INV_X1 U7190 ( .A(n6227), .ZN(n6145) );
  NAND2_X1 U7191 ( .A1(n5462), .A2(n6142), .ZN(n6143) );
  AND2_X1 U7192 ( .A1(n5524), .A2(n6143), .ZN(n6298) );
  AOI222_X1 U7193 ( .A1(n6146), .A2(n6366), .B1(n6145), .B2(n6144), .C1(n6357), 
        .C2(n6298), .ZN(n6147) );
  NAND2_X1 U7194 ( .A1(n6371), .A2(REIP_REG_17__SCAN_IN), .ZN(n6157) );
  OAI211_X1 U7195 ( .C1(n6220), .C2(n6148), .A(n6147), .B(n6157), .ZN(U2969)
         );
  INV_X1 U7196 ( .A(n6149), .ZN(n6150) );
  AOI22_X1 U7197 ( .A1(REIP_REG_25__SCAN_IN), .A2(n6371), .B1(n6150), .B2(
        n6155), .ZN(n6154) );
  AOI22_X1 U7198 ( .A1(n6152), .A2(n6418), .B1(n6412), .B2(n6151), .ZN(n6153)
         );
  OAI211_X1 U7199 ( .C1(n6156), .C2(n6155), .A(n6154), .B(n6153), .ZN(U2993)
         );
  INV_X1 U7200 ( .A(n6157), .ZN(n6158) );
  AOI221_X1 U7201 ( .B1(n6161), .B2(n6160), .C1(n6159), .C2(
        INSTADDRPOINTER_REG_17__SCAN_IN), .A(n6158), .ZN(n6167) );
  NAND2_X1 U7202 ( .A1(n6163), .A2(n6162), .ZN(n6164) );
  NAND2_X1 U7203 ( .A1(n6165), .A2(n6164), .ZN(n6287) );
  INV_X1 U7204 ( .A(n6287), .ZN(n6224) );
  NAND2_X1 U7205 ( .A1(n6412), .A2(n6224), .ZN(n6166) );
  OAI211_X1 U7206 ( .C1(n6168), .C2(n6398), .A(n6167), .B(n6166), .ZN(U3001)
         );
  AND2_X1 U7207 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n6178) );
  OAI211_X1 U7208 ( .C1(INSTADDRPOINTER_REG_15__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .A(n6169), .B(n6375), .ZN(n6177) );
  INV_X1 U7209 ( .A(n6170), .ZN(n6172) );
  AOI21_X1 U7210 ( .B1(n6412), .B2(n6172), .A(n6171), .ZN(n6176) );
  AOI22_X1 U7211 ( .A1(n6174), .A2(n6418), .B1(INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n6173), .ZN(n6175) );
  OAI211_X1 U7212 ( .C1(n6178), .C2(n6177), .A(n6176), .B(n6175), .ZN(U3002)
         );
  AOI21_X1 U7213 ( .B1(n6412), .B2(n6180), .A(n6179), .ZN(n6184) );
  AOI22_X1 U7214 ( .A1(n6182), .A2(n6418), .B1(INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n6181), .ZN(n6183) );
  OAI211_X1 U7215 ( .C1(n6186), .C2(n6185), .A(n6184), .B(n6183), .ZN(U3005)
         );
  INV_X1 U7216 ( .A(STATE_REG_2__SCAN_IN), .ZN(n7040) );
  INV_X1 U7217 ( .A(STATE_REG_0__SCAN_IN), .ZN(n6854) );
  AOI21_X1 U7218 ( .B1(STATE_REG_1__SCAN_IN), .B2(n7040), .A(n6854), .ZN(n6193) );
  INV_X1 U7219 ( .A(ADS_N_REG_SCAN_IN), .ZN(n7060) );
  INV_X1 U7220 ( .A(STATE_REG_1__SCAN_IN), .ZN(n6736) );
  NOR2_X1 U7221 ( .A1(STATE_REG_0__SCAN_IN), .A2(n6736), .ZN(n6653) );
  INV_X1 U7222 ( .A(n6653), .ZN(n7084) );
  INV_X1 U7223 ( .A(n7084), .ZN(n6648) );
  AOI21_X1 U7224 ( .B1(n6193), .B2(n7060), .A(n6648), .ZN(U2789) );
  INV_X1 U7225 ( .A(n6187), .ZN(n6191) );
  INV_X1 U7226 ( .A(n6188), .ZN(n6189) );
  OAI21_X1 U7227 ( .B1(n6189), .B2(n6598), .A(CODEFETCH_REG_SCAN_IN), .ZN(
        n6190) );
  OAI21_X1 U7228 ( .B1(n6191), .B2(n6596), .A(n6190), .ZN(U2790) );
  INV_X1 U7229 ( .A(D_C_N_REG_SCAN_IN), .ZN(n6948) );
  NOR2_X1 U7230 ( .A1(STATE_REG_0__SCAN_IN), .A2(STATE_REG_2__SCAN_IN), .ZN(
        n6194) );
  NOR2_X1 U7231 ( .A1(n6648), .A2(n6194), .ZN(n6192) );
  AOI22_X1 U7232 ( .A1(CODEFETCH_REG_SCAN_IN), .A2(n6648), .B1(n6948), .B2(
        n6192), .ZN(U2791) );
  NOR2_X2 U7233 ( .A1(n6648), .A2(n6193), .ZN(n6661) );
  OAI21_X1 U7234 ( .B1(BS16_N), .B2(n6194), .A(n6661), .ZN(n6659) );
  OAI21_X1 U7235 ( .B1(n6661), .B2(n7056), .A(n6659), .ZN(U2792) );
  OAI21_X1 U7236 ( .B1(n6196), .B2(n7080), .A(n6195), .ZN(U2793) );
  NOR4_X1 U7237 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(DATAWIDTH_REG_4__SCAN_IN), 
        .A3(DATAWIDTH_REG_19__SCAN_IN), .A4(DATAWIDTH_REG_11__SCAN_IN), .ZN(
        n6200) );
  NOR4_X1 U7238 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(
        DATAWIDTH_REG_15__SCAN_IN), .A3(DATAWIDTH_REG_23__SCAN_IN), .A4(
        DATAWIDTH_REG_21__SCAN_IN), .ZN(n6199) );
  NOR4_X1 U7239 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(
        DATAWIDTH_REG_29__SCAN_IN), .A3(DATAWIDTH_REG_30__SCAN_IN), .A4(
        DATAWIDTH_REG_31__SCAN_IN), .ZN(n6198) );
  NOR4_X1 U7240 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(
        DATAWIDTH_REG_25__SCAN_IN), .A3(DATAWIDTH_REG_26__SCAN_IN), .A4(
        DATAWIDTH_REG_27__SCAN_IN), .ZN(n6197) );
  NAND4_X1 U7241 ( .A1(n6200), .A2(n6199), .A3(n6198), .A4(n6197), .ZN(n6206)
         );
  NOR4_X1 U7242 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(DATAWIDTH_REG_7__SCAN_IN), 
        .A3(DATAWIDTH_REG_22__SCAN_IN), .A4(DATAWIDTH_REG_12__SCAN_IN), .ZN(
        n6204) );
  AOI211_X1 U7243 ( .C1(DATAWIDTH_REG_0__SCAN_IN), .C2(
        DATAWIDTH_REG_1__SCAN_IN), .A(DATAWIDTH_REG_14__SCAN_IN), .B(
        DATAWIDTH_REG_5__SCAN_IN), .ZN(n6203) );
  NOR4_X1 U7244 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(DATAWIDTH_REG_20__SCAN_IN), .A3(DATAWIDTH_REG_8__SCAN_IN), .A4(DATAWIDTH_REG_17__SCAN_IN), .ZN(n6202) );
  NOR4_X1 U7245 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(DATAWIDTH_REG_10__SCAN_IN), .A3(DATAWIDTH_REG_16__SCAN_IN), .A4(DATAWIDTH_REG_13__SCAN_IN), .ZN(n6201)
         );
  NAND4_X1 U7246 ( .A1(n6204), .A2(n6203), .A3(n6202), .A4(n6201), .ZN(n6205)
         );
  NOR2_X1 U7247 ( .A1(n6206), .A2(n6205), .ZN(n6670) );
  INV_X1 U7248 ( .A(BYTEENABLE_REG_1__SCAN_IN), .ZN(n6656) );
  NOR3_X1 U7249 ( .A1(REIP_REG_0__SCAN_IN), .A2(DATAWIDTH_REG_0__SCAN_IN), 
        .A3(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6208) );
  OAI21_X1 U7250 ( .B1(REIP_REG_1__SCAN_IN), .B2(n6208), .A(n6670), .ZN(n6207)
         );
  OAI21_X1 U7251 ( .B1(n6670), .B2(n6656), .A(n6207), .ZN(U2794) );
  INV_X1 U7252 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6660) );
  AOI21_X1 U7253 ( .B1(n6667), .B2(n6660), .A(n6208), .ZN(n6209) );
  INV_X1 U7254 ( .A(BYTEENABLE_REG_3__SCAN_IN), .ZN(n6978) );
  INV_X1 U7255 ( .A(n6670), .ZN(n6673) );
  AOI22_X1 U7256 ( .A1(n6670), .A2(n6209), .B1(n6978), .B2(n6673), .ZN(U2795)
         );
  INV_X1 U7257 ( .A(REIP_REG_18__SCAN_IN), .ZN(n6762) );
  AOI22_X1 U7258 ( .A1(REIP_REG_18__SCAN_IN), .A2(n6223), .B1(n6210), .B2(
        n6762), .ZN(n6211) );
  OAI211_X1 U7259 ( .C1(n6273), .C2(n6212), .A(n6211), .B(n6393), .ZN(n6213)
         );
  AOI21_X1 U7260 ( .B1(EBX_REG_18__SCAN_IN), .B2(n6276), .A(n6213), .ZN(n6216)
         );
  AOI22_X1 U7261 ( .A1(n6293), .A2(n6258), .B1(n6247), .B2(n6214), .ZN(n6215)
         );
  OAI211_X1 U7262 ( .C1(n6218), .C2(n6217), .A(n6216), .B(n6215), .ZN(U2809)
         );
  NAND2_X1 U7263 ( .A1(n6646), .A2(n6219), .ZN(n6222) );
  INV_X1 U7264 ( .A(EBX_REG_17__SCAN_IN), .ZN(n6291) );
  OAI22_X1 U7265 ( .A1(n6291), .A2(n6242), .B1(n6220), .B2(n6273), .ZN(n6221)
         );
  AOI211_X1 U7266 ( .C1(n6223), .C2(n6222), .A(n6411), .B(n6221), .ZN(n6226)
         );
  AOI22_X1 U7267 ( .A1(n6298), .A2(n6258), .B1(n6277), .B2(n6224), .ZN(n6225)
         );
  OAI211_X1 U7268 ( .C1(n6227), .C2(n6272), .A(n6226), .B(n6225), .ZN(U2810)
         );
  AOI22_X1 U7269 ( .A1(PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n6229), .B1(n6277), 
        .B2(n6228), .ZN(n6238) );
  NOR3_X1 U7270 ( .A1(n6231), .A2(REIP_REG_12__SCAN_IN), .A3(n6230), .ZN(n6233) );
  NOR2_X1 U7271 ( .A1(n6640), .A2(n6251), .ZN(n6232) );
  AOI211_X1 U7272 ( .C1(n6276), .C2(EBX_REG_12__SCAN_IN), .A(n6233), .B(n6232), 
        .ZN(n6237) );
  AOI22_X1 U7273 ( .A1(n6235), .A2(n6258), .B1(n6234), .B2(n6247), .ZN(n6236)
         );
  NAND4_X1 U7274 ( .A1(n6238), .A2(n6237), .A3(n6236), .A4(n6393), .ZN(U2815)
         );
  AOI21_X1 U7275 ( .B1(n6240), .B2(n6239), .A(REIP_REG_11__SCAN_IN), .ZN(n6252) );
  OAI22_X1 U7276 ( .A1(n6243), .A2(n6242), .B1(n6241), .B2(n6273), .ZN(n6244)
         );
  AOI211_X1 U7277 ( .C1(n6277), .C2(n6372), .A(n6411), .B(n6244), .ZN(n6250)
         );
  INV_X1 U7278 ( .A(n6245), .ZN(n6246) );
  AOI22_X1 U7279 ( .A1(n6248), .A2(n6258), .B1(n6247), .B2(n6246), .ZN(n6249)
         );
  OAI211_X1 U7280 ( .C1(n6252), .C2(n6251), .A(n6250), .B(n6249), .ZN(U2816)
         );
  INV_X1 U7281 ( .A(REIP_REG_6__SCAN_IN), .ZN(n6633) );
  NOR3_X1 U7282 ( .A1(n6253), .A2(REIP_REG_7__SCAN_IN), .A3(n6633), .ZN(n6257)
         );
  INV_X1 U7283 ( .A(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n6255) );
  AOI22_X1 U7284 ( .A1(EBX_REG_7__SCAN_IN), .A2(n6276), .B1(n6277), .B2(n6385), 
        .ZN(n6254) );
  OAI211_X1 U7285 ( .C1(n6273), .C2(n6255), .A(n6393), .B(n6254), .ZN(n6256)
         );
  AOI211_X1 U7286 ( .C1(n6342), .C2(n6258), .A(n6257), .B(n6256), .ZN(n6261)
         );
  OAI21_X1 U7287 ( .B1(n6259), .B2(n6266), .A(REIP_REG_7__SCAN_IN), .ZN(n6260)
         );
  OAI211_X1 U7288 ( .C1(n6272), .C2(n6345), .A(n6261), .B(n6260), .ZN(U2820)
         );
  INV_X1 U7289 ( .A(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n6264) );
  AOI22_X1 U7290 ( .A1(EBX_REG_5__SCAN_IN), .A2(n6276), .B1(n6277), .B2(n6262), 
        .ZN(n6263) );
  OAI211_X1 U7291 ( .C1(n6273), .C2(n6264), .A(n6393), .B(n6263), .ZN(n6265)
         );
  AOI21_X1 U7292 ( .B1(n6347), .B2(n6283), .A(n6265), .ZN(n6269) );
  OAI21_X1 U7293 ( .B1(REIP_REG_5__SCAN_IN), .B2(n6267), .A(n6266), .ZN(n6268)
         );
  OAI211_X1 U7294 ( .C1(n6272), .C2(n6351), .A(n6269), .B(n6268), .ZN(U2822)
         );
  INV_X1 U7295 ( .A(REIP_REG_3__SCAN_IN), .ZN(n6629) );
  INV_X1 U7296 ( .A(n6270), .ZN(n6271) );
  NAND2_X1 U7297 ( .A1(n6271), .A2(REIP_REG_2__SCAN_IN), .ZN(n6285) );
  INV_X1 U7298 ( .A(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n6274) );
  OAI22_X1 U7299 ( .A1(n6274), .A2(n6273), .B1(n6272), .B2(n6360), .ZN(n6275)
         );
  AOI21_X1 U7300 ( .B1(n6276), .B2(EBX_REG_3__SCAN_IN), .A(n6275), .ZN(n6279)
         );
  NAND2_X1 U7301 ( .A1(n6277), .A2(n6405), .ZN(n6278) );
  OAI211_X1 U7302 ( .C1(n6281), .C2(n6280), .A(n6279), .B(n6278), .ZN(n6282)
         );
  AOI21_X1 U7303 ( .B1(n6356), .B2(n6283), .A(n6282), .ZN(n6284) );
  OAI221_X1 U7304 ( .B1(n6286), .B2(n6629), .C1(n6286), .C2(n6285), .A(n6284), 
        .ZN(U2824) );
  NOR2_X1 U7305 ( .A1(n6288), .A2(n6287), .ZN(n6289) );
  AOI21_X1 U7306 ( .B1(n6298), .B2(n4396), .A(n6289), .ZN(n6290) );
  OAI21_X1 U7307 ( .B1(n6292), .B2(n6291), .A(n6290), .ZN(U2842) );
  AOI22_X1 U7308 ( .A1(n6293), .A2(n6297), .B1(n6296), .B2(DATAI_18_), .ZN(
        n6295) );
  AOI22_X1 U7309 ( .A1(n6300), .A2(DATAI_2_), .B1(EAX_REG_18__SCAN_IN), .B2(
        n6299), .ZN(n6294) );
  NAND2_X1 U7310 ( .A1(n6295), .A2(n6294), .ZN(U2873) );
  AOI22_X1 U7311 ( .A1(n6298), .A2(n6297), .B1(n6296), .B2(DATAI_17_), .ZN(
        n6302) );
  AOI22_X1 U7312 ( .A1(n6300), .A2(DATAI_1_), .B1(EAX_REG_17__SCAN_IN), .B2(
        n6299), .ZN(n6301) );
  NAND2_X1 U7313 ( .A1(n6302), .A2(n6301), .ZN(U2874) );
  AOI22_X1 U7314 ( .A1(n6333), .A2(LWORD_REG_15__SCAN_IN), .B1(n6323), .B2(
        DATAO_REG_15__SCAN_IN), .ZN(n6303) );
  OAI21_X1 U7315 ( .B1(n4421), .B2(n6335), .A(n6303), .ZN(U2908) );
  AOI22_X1 U7316 ( .A1(n6333), .A2(LWORD_REG_14__SCAN_IN), .B1(n6323), .B2(
        DATAO_REG_14__SCAN_IN), .ZN(n6304) );
  OAI21_X1 U7317 ( .B1(n6305), .B2(n6335), .A(n6304), .ZN(U2909) );
  AOI22_X1 U7318 ( .A1(n6333), .A2(LWORD_REG_13__SCAN_IN), .B1(n6323), .B2(
        DATAO_REG_13__SCAN_IN), .ZN(n6306) );
  OAI21_X1 U7319 ( .B1(n6307), .B2(n6335), .A(n6306), .ZN(U2910) );
  AOI22_X1 U7320 ( .A1(n6333), .A2(LWORD_REG_12__SCAN_IN), .B1(n6323), .B2(
        DATAO_REG_12__SCAN_IN), .ZN(n6308) );
  OAI21_X1 U7321 ( .B1(n3597), .B2(n6335), .A(n6308), .ZN(U2911) );
  AOI22_X1 U7322 ( .A1(n6333), .A2(LWORD_REG_11__SCAN_IN), .B1(n6323), .B2(
        DATAO_REG_11__SCAN_IN), .ZN(n6309) );
  OAI21_X1 U7323 ( .B1(n6310), .B2(n6335), .A(n6309), .ZN(U2912) );
  AOI22_X1 U7324 ( .A1(n6333), .A2(LWORD_REG_10__SCAN_IN), .B1(n6323), .B2(
        DATAO_REG_10__SCAN_IN), .ZN(n6311) );
  OAI21_X1 U7325 ( .B1(n6312), .B2(n6335), .A(n6311), .ZN(U2913) );
  AOI22_X1 U7326 ( .A1(n6333), .A2(LWORD_REG_9__SCAN_IN), .B1(n6323), .B2(
        DATAO_REG_9__SCAN_IN), .ZN(n6313) );
  OAI21_X1 U7327 ( .B1(n6314), .B2(n6335), .A(n6313), .ZN(U2914) );
  AOI22_X1 U7328 ( .A1(n6333), .A2(LWORD_REG_8__SCAN_IN), .B1(n6323), .B2(
        DATAO_REG_8__SCAN_IN), .ZN(n6315) );
  OAI21_X1 U7329 ( .B1(n6316), .B2(n6335), .A(n6315), .ZN(U2915) );
  AOI22_X1 U7330 ( .A1(n6333), .A2(LWORD_REG_7__SCAN_IN), .B1(n6323), .B2(
        DATAO_REG_7__SCAN_IN), .ZN(n6317) );
  OAI21_X1 U7331 ( .B1(n6318), .B2(n6335), .A(n6317), .ZN(U2916) );
  AOI22_X1 U7332 ( .A1(n6333), .A2(LWORD_REG_6__SCAN_IN), .B1(n6323), .B2(
        DATAO_REG_6__SCAN_IN), .ZN(n6319) );
  OAI21_X1 U7333 ( .B1(n6320), .B2(n6335), .A(n6319), .ZN(U2917) );
  AOI22_X1 U7334 ( .A1(n6333), .A2(LWORD_REG_5__SCAN_IN), .B1(n6323), .B2(
        DATAO_REG_5__SCAN_IN), .ZN(n6321) );
  OAI21_X1 U7335 ( .B1(n6322), .B2(n6335), .A(n6321), .ZN(U2918) );
  AOI22_X1 U7336 ( .A1(n6333), .A2(LWORD_REG_4__SCAN_IN), .B1(n6323), .B2(
        DATAO_REG_4__SCAN_IN), .ZN(n6324) );
  OAI21_X1 U7337 ( .B1(n6325), .B2(n6335), .A(n6324), .ZN(U2919) );
  AOI22_X1 U7338 ( .A1(n6333), .A2(LWORD_REG_3__SCAN_IN), .B1(n6332), .B2(
        DATAO_REG_3__SCAN_IN), .ZN(n6326) );
  OAI21_X1 U7339 ( .B1(n6327), .B2(n6335), .A(n6326), .ZN(U2920) );
  AOI22_X1 U7340 ( .A1(n6333), .A2(LWORD_REG_2__SCAN_IN), .B1(n6332), .B2(
        DATAO_REG_2__SCAN_IN), .ZN(n6328) );
  OAI21_X1 U7341 ( .B1(n6329), .B2(n6335), .A(n6328), .ZN(U2921) );
  AOI22_X1 U7342 ( .A1(n6333), .A2(LWORD_REG_1__SCAN_IN), .B1(n6332), .B2(
        DATAO_REG_1__SCAN_IN), .ZN(n6330) );
  OAI21_X1 U7343 ( .B1(n6331), .B2(n6335), .A(n6330), .ZN(U2922) );
  AOI22_X1 U7344 ( .A1(n6333), .A2(LWORD_REG_0__SCAN_IN), .B1(n6332), .B2(
        DATAO_REG_0__SCAN_IN), .ZN(n6334) );
  OAI21_X1 U7345 ( .B1(n6336), .B2(n6335), .A(n6334), .ZN(U2923) );
  AOI22_X1 U7346 ( .A1(n6371), .A2(REIP_REG_7__SCAN_IN), .B1(n6361), .B2(
        PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n6344) );
  CLKBUF_X1 U7347 ( .A(n6338), .Z(n6339) );
  OAI21_X1 U7348 ( .B1(n6337), .B2(n6340), .A(n6339), .ZN(n6341) );
  INV_X1 U7349 ( .A(n6341), .ZN(n6387) );
  AOI22_X1 U7350 ( .A1(n6387), .A2(n6366), .B1(n6357), .B2(n6342), .ZN(n6343)
         );
  OAI211_X1 U7351 ( .C1(n6370), .C2(n6345), .A(n6344), .B(n6343), .ZN(U2979)
         );
  AOI22_X1 U7352 ( .A1(n6371), .A2(REIP_REG_5__SCAN_IN), .B1(n6361), .B2(
        PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n6350) );
  INV_X1 U7353 ( .A(n6346), .ZN(n6348) );
  AOI22_X1 U7354 ( .A1(n6348), .A2(n6366), .B1(n6357), .B2(n6347), .ZN(n6349)
         );
  OAI211_X1 U7355 ( .C1(n6370), .C2(n6351), .A(n6350), .B(n6349), .ZN(U2981)
         );
  AOI22_X1 U7356 ( .A1(n6371), .A2(REIP_REG_3__SCAN_IN), .B1(n6361), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n6359) );
  OAI21_X1 U7357 ( .B1(n6352), .B2(n6354), .A(n6353), .ZN(n6355) );
  INV_X1 U7358 ( .A(n6355), .ZN(n6404) );
  AOI22_X1 U7359 ( .A1(n6357), .A2(n6356), .B1(n6404), .B2(n6366), .ZN(n6358)
         );
  OAI211_X1 U7360 ( .C1(n6370), .C2(n6360), .A(n6359), .B(n6358), .ZN(U2983)
         );
  AOI22_X1 U7361 ( .A1(n6411), .A2(REIP_REG_2__SCAN_IN), .B1(n6361), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n6368) );
  XOR2_X1 U7362 ( .A(n6363), .B(INSTADDRPOINTER_REG_2__SCAN_IN), .Z(n6364) );
  XNOR2_X1 U7363 ( .A(n6362), .B(n6364), .ZN(n6419) );
  AOI22_X1 U7364 ( .A1(n6419), .A2(n6366), .B1(n6365), .B2(n6357), .ZN(n6367)
         );
  OAI211_X1 U7365 ( .C1(n6370), .C2(n6369), .A(n6368), .B(n6367), .ZN(U2984)
         );
  INV_X1 U7366 ( .A(REIP_REG_11__SCAN_IN), .ZN(n6639) );
  AOI22_X1 U7367 ( .A1(n6373), .A2(n6418), .B1(n6412), .B2(n6372), .ZN(n6377)
         );
  OAI21_X1 U7368 ( .B1(INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n6375), .A(n6374), 
        .ZN(n6376) );
  OAI211_X1 U7369 ( .C1(n6639), .C2(n6393), .A(n6377), .B(n6376), .ZN(U3007)
         );
  AOI21_X1 U7370 ( .B1(n6412), .B2(n6379), .A(n6378), .ZN(n6383) );
  AOI22_X1 U7371 ( .A1(n6381), .A2(n6418), .B1(INSTADDRPOINTER_REG_9__SCAN_IN), 
        .B2(n6380), .ZN(n6382) );
  OAI211_X1 U7372 ( .C1(INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n6384), .A(n6383), 
        .B(n6382), .ZN(U3009) );
  AOI22_X1 U7373 ( .A1(n6412), .A2(n6385), .B1(n6411), .B2(REIP_REG_7__SCAN_IN), .ZN(n6389) );
  AOI22_X1 U7374 ( .A1(n6387), .A2(n6418), .B1(n6386), .B2(n6390), .ZN(n6388)
         );
  OAI211_X1 U7375 ( .C1(n6391), .C2(n6390), .A(n6389), .B(n6388), .ZN(U3011)
         );
  AOI21_X1 U7376 ( .B1(n6414), .B2(n6416), .A(n6417), .ZN(n6407) );
  AOI211_X1 U7377 ( .C1(n6408), .C2(n6403), .A(n6392), .B(n6409), .ZN(n6401)
         );
  OAI22_X1 U7378 ( .A1(n6395), .A2(n6394), .B1(n6630), .B2(n6393), .ZN(n6396)
         );
  INV_X1 U7379 ( .A(n6396), .ZN(n6397) );
  OAI21_X1 U7380 ( .B1(n6399), .B2(n6398), .A(n6397), .ZN(n6400) );
  NOR2_X1 U7381 ( .A1(n6401), .A2(n6400), .ZN(n6402) );
  OAI21_X1 U7382 ( .B1(n6407), .B2(n6403), .A(n6402), .ZN(U3014) );
  AOI222_X1 U7383 ( .A1(REIP_REG_3__SCAN_IN), .A2(n6371), .B1(n6412), .B2(
        n6405), .C1(n6418), .C2(n6404), .ZN(n6406) );
  OAI221_X1 U7384 ( .B1(INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n6409), .C1(n6408), .C2(n6407), .A(n6406), .ZN(U3015) );
  INV_X1 U7385 ( .A(n6410), .ZN(n6413) );
  AOI22_X1 U7386 ( .A1(n6413), .A2(n6412), .B1(n6411), .B2(REIP_REG_2__SCAN_IN), .ZN(n6424) );
  OAI221_X1 U7387 ( .B1(n6416), .B2(n6415), .C1(n6416), .C2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .A(n6414), .ZN(n6423) );
  AOI22_X1 U7388 ( .A1(n6419), .A2(n6418), .B1(INSTADDRPOINTER_REG_2__SCAN_IN), 
        .B2(n6417), .ZN(n6422) );
  NAND3_X1 U7389 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n6420), .A3(n4237), 
        .ZN(n6421) );
  NAND4_X1 U7390 ( .A1(n6424), .A2(n6423), .A3(n6422), .A4(n6421), .ZN(U3016)
         );
  NOR2_X1 U7391 ( .A1(n6426), .A2(n6425), .ZN(U3019) );
  INV_X1 U7392 ( .A(n6427), .ZN(n6435) );
  AOI22_X1 U7393 ( .A1(n6436), .A2(n6464), .B1(n6463), .B2(n6435), .ZN(n6429)
         );
  AOI22_X1 U7394 ( .A1(INSTQUEUE_REG_3__2__SCAN_IN), .A2(n6439), .B1(n6462), 
        .B2(n6437), .ZN(n6428) );
  OAI211_X1 U7395 ( .C1(n6443), .C2(n6430), .A(n6429), .B(n6428), .ZN(U3046)
         );
  AOI22_X1 U7396 ( .A1(n6436), .A2(n6520), .B1(n6518), .B2(n6435), .ZN(n6433)
         );
  AOI22_X1 U7397 ( .A1(INSTQUEUE_REG_3__3__SCAN_IN), .A2(n6439), .B1(n6431), 
        .B2(n6437), .ZN(n6432) );
  OAI211_X1 U7398 ( .C1(n6443), .C2(n6434), .A(n6433), .B(n6432), .ZN(U3047)
         );
  AOI22_X1 U7399 ( .A1(n6436), .A2(n6535), .B1(n6533), .B2(n6435), .ZN(n6441)
         );
  AOI22_X1 U7400 ( .A1(INSTQUEUE_REG_3__5__SCAN_IN), .A2(n6439), .B1(n6438), 
        .B2(n6437), .ZN(n6440) );
  OAI211_X1 U7401 ( .C1(n6443), .C2(n6442), .A(n6441), .B(n6440), .ZN(U3049)
         );
  NOR2_X1 U7402 ( .A1(n6444), .A2(n6498), .ZN(n6454) );
  NOR2_X1 U7403 ( .A1(n3463), .A2(n6445), .ZN(n6447) );
  INV_X1 U7404 ( .A(n6446), .ZN(n6477) );
  AOI21_X1 U7405 ( .B1(n6448), .B2(n6447), .A(n6477), .ZN(n6453) );
  INV_X1 U7406 ( .A(n6453), .ZN(n6449) );
  AOI22_X1 U7407 ( .A1(n6454), .A2(n6449), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n6457), .ZN(n6483) );
  AOI22_X1 U7408 ( .A1(n6478), .A2(n6452), .B1(n6451), .B2(n6477), .ZN(n6459)
         );
  NAND2_X1 U7409 ( .A1(n6454), .A2(n6453), .ZN(n6456) );
  OAI211_X1 U7410 ( .C1(n6457), .C2(n6484), .A(n6456), .B(n6455), .ZN(n6480)
         );
  AOI22_X1 U7411 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n6480), .B1(n6502), 
        .B2(n6479), .ZN(n6458) );
  OAI211_X1 U7412 ( .C1(n6483), .C2(n6505), .A(n6459), .B(n6458), .ZN(U3076)
         );
  AOI22_X1 U7413 ( .A1(n6507), .A2(n6479), .B1(n6506), .B2(n6477), .ZN(n6461)
         );
  AOI22_X1 U7414 ( .A1(n6480), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n6508), 
        .B2(n6478), .ZN(n6460) );
  OAI211_X1 U7415 ( .C1(n6483), .C2(n6511), .A(n6461), .B(n6460), .ZN(U3077)
         );
  AOI22_X1 U7416 ( .A1(n6515), .A2(n6479), .B1(n6463), .B2(n6477), .ZN(n6466)
         );
  AOI22_X1 U7417 ( .A1(n6480), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n6464), 
        .B2(n6478), .ZN(n6465) );
  OAI211_X1 U7418 ( .C1(n6483), .C2(n5452), .A(n6466), .B(n6465), .ZN(U3078)
         );
  AOI22_X1 U7419 ( .A1(n6478), .A2(n6520), .B1(n6518), .B2(n6477), .ZN(n6468)
         );
  AOI22_X1 U7420 ( .A1(INSTQUEUE_REG_7__3__SCAN_IN), .A2(n6480), .B1(n6519), 
        .B2(n6479), .ZN(n6467) );
  OAI211_X1 U7421 ( .C1(n6483), .C2(n6523), .A(n6468), .B(n6467), .ZN(U3079)
         );
  AOI22_X1 U7422 ( .A1(n6529), .A2(n6479), .B1(n6469), .B2(n6477), .ZN(n6472)
         );
  AOI22_X1 U7423 ( .A1(n6480), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n6470), 
        .B2(n6478), .ZN(n6471) );
  OAI211_X1 U7424 ( .C1(n6483), .C2(n6532), .A(n6472), .B(n6471), .ZN(U3080)
         );
  AOI22_X1 U7425 ( .A1(n6534), .A2(n6479), .B1(n6533), .B2(n6477), .ZN(n6474)
         );
  AOI22_X1 U7426 ( .A1(n6480), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n6535), 
        .B2(n6478), .ZN(n6473) );
  OAI211_X1 U7427 ( .C1(n6483), .C2(n6538), .A(n6474), .B(n6473), .ZN(U3081)
         );
  AOI22_X1 U7428 ( .A1(n6478), .A2(n6541), .B1(n6539), .B2(n6477), .ZN(n6476)
         );
  AOI22_X1 U7429 ( .A1(INSTQUEUE_REG_7__6__SCAN_IN), .A2(n6480), .B1(n6540), 
        .B2(n6479), .ZN(n6475) );
  OAI211_X1 U7430 ( .C1(n6483), .C2(n6544), .A(n6476), .B(n6475), .ZN(U3082)
         );
  AOI22_X1 U7431 ( .A1(n6478), .A2(n6550), .B1(n6546), .B2(n6477), .ZN(n6482)
         );
  AOI22_X1 U7432 ( .A1(INSTQUEUE_REG_7__7__SCAN_IN), .A2(n6480), .B1(n6547), 
        .B2(n6479), .ZN(n6481) );
  OAI211_X1 U7433 ( .C1(n6483), .C2(n6554), .A(n6482), .B(n6481), .ZN(U3083)
         );
  OAI21_X1 U7434 ( .B1(n6486), .B2(n6485), .A(n6484), .ZN(n6501) );
  INV_X1 U7435 ( .A(n6501), .ZN(n6492) );
  NAND2_X1 U7436 ( .A1(n6488), .A2(n6487), .ZN(n6490) );
  NAND2_X1 U7437 ( .A1(n6489), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6524) );
  NAND2_X1 U7438 ( .A1(n6490), .A2(n6524), .ZN(n6500) );
  INV_X1 U7439 ( .A(n6497), .ZN(n6491) );
  AOI22_X1 U7440 ( .A1(n6492), .A2(n6500), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n6491), .ZN(n6555) );
  OAI22_X1 U7441 ( .A1(n6527), .A2(n6494), .B1(n6493), .B2(n6524), .ZN(n6495)
         );
  INV_X1 U7442 ( .A(n6495), .ZN(n6504) );
  AOI21_X1 U7443 ( .B1(n6498), .B2(n6497), .A(n6496), .ZN(n6499) );
  OAI21_X1 U7444 ( .B1(n6501), .B2(n6500), .A(n6499), .ZN(n6551) );
  AOI22_X1 U7445 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n6551), .B1(n6502), 
        .B2(n6548), .ZN(n6503) );
  OAI211_X1 U7446 ( .C1(n6555), .C2(n6505), .A(n6504), .B(n6503), .ZN(U3108)
         );
  INV_X1 U7447 ( .A(n6524), .ZN(n6545) );
  AOI22_X1 U7448 ( .A1(n6548), .A2(n6507), .B1(n6506), .B2(n6545), .ZN(n6510)
         );
  AOI22_X1 U7449 ( .A1(n6551), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n6508), 
        .B2(n6549), .ZN(n6509) );
  OAI211_X1 U7450 ( .C1(n6555), .C2(n6511), .A(n6510), .B(n6509), .ZN(U3109)
         );
  OAI22_X1 U7451 ( .A1(n6527), .A2(n6513), .B1(n6512), .B2(n6524), .ZN(n6514)
         );
  INV_X1 U7452 ( .A(n6514), .ZN(n6517) );
  AOI22_X1 U7453 ( .A1(INSTQUEUE_REG_11__2__SCAN_IN), .A2(n6551), .B1(n6515), 
        .B2(n6548), .ZN(n6516) );
  OAI211_X1 U7454 ( .C1(n6555), .C2(n5452), .A(n6517), .B(n6516), .ZN(U3110)
         );
  AOI22_X1 U7455 ( .A1(n6548), .A2(n6519), .B1(n6518), .B2(n6545), .ZN(n6522)
         );
  AOI22_X1 U7456 ( .A1(n6551), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n6520), 
        .B2(n6549), .ZN(n6521) );
  OAI211_X1 U7457 ( .C1(n6555), .C2(n6523), .A(n6522), .B(n6521), .ZN(U3111)
         );
  OAI22_X1 U7458 ( .A1(n6527), .A2(n6526), .B1(n6525), .B2(n6524), .ZN(n6528)
         );
  INV_X1 U7459 ( .A(n6528), .ZN(n6531) );
  AOI22_X1 U7460 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n6551), .B1(n6529), 
        .B2(n6548), .ZN(n6530) );
  OAI211_X1 U7461 ( .C1(n6555), .C2(n6532), .A(n6531), .B(n6530), .ZN(U3112)
         );
  AOI22_X1 U7462 ( .A1(n6548), .A2(n6534), .B1(n6533), .B2(n6545), .ZN(n6537)
         );
  AOI22_X1 U7463 ( .A1(n6551), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n6535), 
        .B2(n6549), .ZN(n6536) );
  OAI211_X1 U7464 ( .C1(n6555), .C2(n6538), .A(n6537), .B(n6536), .ZN(U3113)
         );
  AOI22_X1 U7465 ( .A1(n6548), .A2(n6540), .B1(n6539), .B2(n6545), .ZN(n6543)
         );
  AOI22_X1 U7466 ( .A1(n6551), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n6541), 
        .B2(n6549), .ZN(n6542) );
  OAI211_X1 U7467 ( .C1(n6555), .C2(n6544), .A(n6543), .B(n6542), .ZN(U3114)
         );
  AOI22_X1 U7468 ( .A1(n6548), .A2(n6547), .B1(n6546), .B2(n6545), .ZN(n6553)
         );
  AOI22_X1 U7469 ( .A1(n6551), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n6550), 
        .B2(n6549), .ZN(n6552) );
  OAI211_X1 U7470 ( .C1(n6555), .C2(n6554), .A(n6553), .B(n6552), .ZN(U3115)
         );
  AND2_X1 U7471 ( .A1(n6561), .A2(n6556), .ZN(n6572) );
  INV_X1 U7472 ( .A(n6557), .ZN(n6560) );
  NOR3_X1 U7473 ( .A1(n6560), .A2(n6559), .A3(n6558), .ZN(n6564) );
  NAND2_X1 U7474 ( .A1(n6564), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6566) );
  INV_X1 U7475 ( .A(n6561), .ZN(n6567) );
  INV_X1 U7476 ( .A(n6562), .ZN(n6563) );
  OAI22_X1 U7477 ( .A1(n6564), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B1(n6567), .B2(n6563), .ZN(n6565) );
  NAND2_X1 U7478 ( .A1(n6566), .A2(n6565), .ZN(n6570) );
  NAND2_X1 U7479 ( .A1(n6561), .A2(n6568), .ZN(n6569) );
  AOI222_X1 U7480 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n6570), .B1(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n6569), .C1(n6570), .C2(n6569), 
        .ZN(n6571) );
  AOI222_X1 U7481 ( .A1(n6573), .A2(n6572), .B1(n6573), .B2(n6571), .C1(n6572), 
        .C2(n6571), .ZN(n6581) );
  INV_X1 U7482 ( .A(n6574), .ZN(n6576) );
  NOR3_X1 U7483 ( .A1(n6577), .A2(n6576), .A3(n6575), .ZN(n6580) );
  OAI21_X1 U7484 ( .B1(FLUSH_REG_SCAN_IN), .B2(MORE_REG_SCAN_IN), .A(n6578), 
        .ZN(n6579) );
  OAI211_X1 U7485 ( .C1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .C2(n6581), .A(n6580), .B(n6579), .ZN(n6585) );
  AOI21_X1 U7486 ( .B1(n6583), .B2(n6585), .A(n6582), .ZN(n6594) );
  OAI22_X1 U7487 ( .A1(n6585), .A2(n6598), .B1(n6584), .B2(n7028), .ZN(n6586)
         );
  OAI21_X1 U7488 ( .B1(n6588), .B2(n6587), .A(n6586), .ZN(n6665) );
  AOI21_X1 U7489 ( .B1(n6680), .B2(n6589), .A(STATE2_REG_0__SCAN_IN), .ZN(
        n6592) );
  NAND2_X1 U7490 ( .A1(READY_N), .A2(n6590), .ZN(n6606) );
  AOI21_X1 U7491 ( .B1(n6606), .B2(n6665), .A(n6596), .ZN(n6591) );
  AOI21_X1 U7492 ( .B1(n6665), .B2(n6592), .A(n6591), .ZN(n6593) );
  OAI211_X1 U7493 ( .C1(n6596), .C2(n6595), .A(n6594), .B(n6593), .ZN(U3148)
         );
  NAND2_X1 U7494 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n6597), .ZN(n6599) );
  OAI21_X1 U7495 ( .B1(READY_N), .B2(n6599), .A(n6598), .ZN(n6604) );
  AOI211_X1 U7496 ( .C1(n6665), .C2(n6606), .A(n6601), .B(n6600), .ZN(n6602)
         );
  AOI211_X1 U7497 ( .C1(n6665), .C2(n6604), .A(n6603), .B(n6602), .ZN(n6605)
         );
  INV_X1 U7498 ( .A(n6605), .ZN(U3149) );
  NAND4_X1 U7499 ( .A1(n6608), .A2(n6607), .A3(n6606), .A4(n6663), .ZN(n6609)
         );
  NAND2_X1 U7500 ( .A1(n6610), .A2(n6609), .ZN(U3150) );
  INV_X1 U7501 ( .A(n6661), .ZN(n6658) );
  AND2_X1 U7502 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(n6658), .ZN(U3151) );
  AND2_X1 U7503 ( .A1(DATAWIDTH_REG_30__SCAN_IN), .A2(n6658), .ZN(U3152) );
  AND2_X1 U7504 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(n6658), .ZN(U3153) );
  AND2_X1 U7505 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(n6658), .ZN(U3154) );
  AND2_X1 U7506 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(n6658), .ZN(U3155) );
  AND2_X1 U7507 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(n6658), .ZN(U3156) );
  AND2_X1 U7508 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(n6658), .ZN(U3157) );
  AND2_X1 U7509 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(n6658), .ZN(U3158) );
  INV_X1 U7510 ( .A(DATAWIDTH_REG_23__SCAN_IN), .ZN(n6782) );
  NOR2_X1 U7511 ( .A1(n6661), .A2(n6782), .ZN(U3159) );
  INV_X1 U7512 ( .A(DATAWIDTH_REG_22__SCAN_IN), .ZN(n6772) );
  NOR2_X1 U7513 ( .A1(n6661), .A2(n6772), .ZN(U3160) );
  INV_X1 U7514 ( .A(DATAWIDTH_REG_21__SCAN_IN), .ZN(n7008) );
  NOR2_X1 U7515 ( .A1(n6661), .A2(n7008), .ZN(U3161) );
  AND2_X1 U7516 ( .A1(n6658), .A2(DATAWIDTH_REG_20__SCAN_IN), .ZN(U3162) );
  INV_X1 U7517 ( .A(DATAWIDTH_REG_19__SCAN_IN), .ZN(n7051) );
  NOR2_X1 U7518 ( .A1(n6661), .A2(n7051), .ZN(U3163) );
  INV_X1 U7519 ( .A(DATAWIDTH_REG_18__SCAN_IN), .ZN(n6991) );
  NOR2_X1 U7520 ( .A1(n6661), .A2(n6991), .ZN(U3164) );
  INV_X1 U7521 ( .A(DATAWIDTH_REG_17__SCAN_IN), .ZN(n6849) );
  NOR2_X1 U7522 ( .A1(n6661), .A2(n6849), .ZN(U3165) );
  AND2_X1 U7523 ( .A1(n6658), .A2(DATAWIDTH_REG_16__SCAN_IN), .ZN(U3166) );
  AND2_X1 U7524 ( .A1(n6658), .A2(DATAWIDTH_REG_15__SCAN_IN), .ZN(U3167) );
  INV_X1 U7525 ( .A(DATAWIDTH_REG_14__SCAN_IN), .ZN(n6814) );
  NOR2_X1 U7526 ( .A1(n6661), .A2(n6814), .ZN(U3168) );
  INV_X1 U7527 ( .A(DATAWIDTH_REG_13__SCAN_IN), .ZN(n6851) );
  NOR2_X1 U7528 ( .A1(n6661), .A2(n6851), .ZN(U3169) );
  INV_X1 U7529 ( .A(DATAWIDTH_REG_12__SCAN_IN), .ZN(n6760) );
  NOR2_X1 U7530 ( .A1(n6661), .A2(n6760), .ZN(U3170) );
  INV_X1 U7531 ( .A(DATAWIDTH_REG_11__SCAN_IN), .ZN(n7022) );
  NOR2_X1 U7532 ( .A1(n6661), .A2(n7022), .ZN(U3171) );
  AND2_X1 U7533 ( .A1(n6658), .A2(DATAWIDTH_REG_10__SCAN_IN), .ZN(U3172) );
  AND2_X1 U7534 ( .A1(n6658), .A2(DATAWIDTH_REG_9__SCAN_IN), .ZN(U3173) );
  INV_X1 U7535 ( .A(DATAWIDTH_REG_8__SCAN_IN), .ZN(n6954) );
  NOR2_X1 U7536 ( .A1(n6661), .A2(n6954), .ZN(U3174) );
  AND2_X1 U7537 ( .A1(n6658), .A2(DATAWIDTH_REG_7__SCAN_IN), .ZN(U3175) );
  INV_X1 U7538 ( .A(DATAWIDTH_REG_6__SCAN_IN), .ZN(n7011) );
  NOR2_X1 U7539 ( .A1(n6661), .A2(n7011), .ZN(U3176) );
  INV_X1 U7540 ( .A(DATAWIDTH_REG_5__SCAN_IN), .ZN(n6798) );
  NOR2_X1 U7541 ( .A1(n6661), .A2(n6798), .ZN(U3177) );
  INV_X1 U7542 ( .A(DATAWIDTH_REG_4__SCAN_IN), .ZN(n7053) );
  NOR2_X1 U7543 ( .A1(n6661), .A2(n7053), .ZN(U3178) );
  AND2_X1 U7544 ( .A1(n6658), .A2(DATAWIDTH_REG_3__SCAN_IN), .ZN(U3179) );
  AND2_X1 U7545 ( .A1(n6658), .A2(DATAWIDTH_REG_2__SCAN_IN), .ZN(U3180) );
  INV_X1 U7546 ( .A(n6621), .ZN(n6613) );
  NAND2_X1 U7547 ( .A1(STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n6619) );
  INV_X1 U7548 ( .A(n6619), .ZN(n6617) );
  AOI21_X1 U7549 ( .B1(STATE_REG_1__SCAN_IN), .B2(READY_N), .A(n6617), .ZN(
        n6612) );
  INV_X1 U7550 ( .A(HOLD), .ZN(n6785) );
  NOR2_X1 U7551 ( .A1(n6736), .A2(n6785), .ZN(n6614) );
  INV_X1 U7552 ( .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6808) );
  OAI21_X1 U7553 ( .B1(n6614), .B2(n6808), .A(n7084), .ZN(n6611) );
  OAI211_X1 U7554 ( .C1(NA_N), .C2(n7040), .A(n6854), .B(n6621), .ZN(n6622) );
  OAI211_X1 U7555 ( .C1(n6613), .C2(n6612), .A(n6611), .B(n6622), .ZN(U3181)
         );
  AOI21_X1 U7556 ( .B1(REQUESTPENDING_REG_SCAN_IN), .B2(STATE_REG_0__SCAN_IN), 
        .A(n6614), .ZN(n6616) );
  NAND2_X1 U7557 ( .A1(READY_N), .A2(STATE_REG_1__SCAN_IN), .ZN(n6620) );
  OAI211_X1 U7558 ( .C1(n6617), .C2(n6616), .A(n6615), .B(n6620), .ZN(U3182)
         );
  NOR2_X1 U7559 ( .A1(NA_N), .A2(n7028), .ZN(n6624) );
  OAI211_X1 U7560 ( .C1(n6624), .C2(n6736), .A(HOLD), .B(n6808), .ZN(n6618) );
  OAI211_X1 U7561 ( .C1(n6621), .C2(n6620), .A(n6619), .B(n6618), .ZN(n6623)
         );
  OAI21_X1 U7562 ( .B1(n6854), .B2(n6623), .A(n6622), .ZN(n6626) );
  NAND4_X1 U7563 ( .A1(STATE_REG_0__SCAN_IN), .A2(STATE_REG_1__SCAN_IN), .A3(
        REQUESTPENDING_REG_SCAN_IN), .A4(n6624), .ZN(n6625) );
  NAND2_X1 U7564 ( .A1(n6626), .A2(n6625), .ZN(U3183) );
  INV_X1 U7565 ( .A(ADDRESS_REG_0__SCAN_IN), .ZN(n6627) );
  INV_X1 U7566 ( .A(n7084), .ZN(n7085) );
  OAI222_X1 U7567 ( .A1(n6655), .A2(n5346), .B1(n6627), .B2(n7085), .C1(n6667), 
        .C2(n6654), .ZN(U3184) );
  INV_X1 U7568 ( .A(ADDRESS_REG_1__SCAN_IN), .ZN(n6628) );
  OAI222_X1 U7569 ( .A1(n6654), .A2(n5346), .B1(n6628), .B2(n7085), .C1(n6629), 
        .C2(n6655), .ZN(U3185) );
  INV_X1 U7570 ( .A(ADDRESS_REG_2__SCAN_IN), .ZN(n6823) );
  OAI222_X1 U7571 ( .A1(n6654), .A2(n6629), .B1(n6823), .B2(n7085), .C1(n6630), 
        .C2(n6655), .ZN(U3186) );
  INV_X1 U7572 ( .A(ADDRESS_REG_3__SCAN_IN), .ZN(n6833) );
  OAI222_X1 U7573 ( .A1(n6654), .A2(n6630), .B1(n6833), .B2(n7085), .C1(n6631), 
        .C2(n6655), .ZN(U3187) );
  INV_X1 U7574 ( .A(ADDRESS_REG_4__SCAN_IN), .ZN(n6835) );
  OAI222_X1 U7575 ( .A1(n6655), .A2(n6633), .B1(n6835), .B2(n7085), .C1(n6631), 
        .C2(n6654), .ZN(U3188) );
  INV_X1 U7576 ( .A(ADDRESS_REG_5__SCAN_IN), .ZN(n6632) );
  INV_X1 U7577 ( .A(REIP_REG_7__SCAN_IN), .ZN(n6635) );
  OAI222_X1 U7578 ( .A1(n6654), .A2(n6633), .B1(n6632), .B2(n7085), .C1(n6635), 
        .C2(n6655), .ZN(U3189) );
  INV_X1 U7579 ( .A(ADDRESS_REG_6__SCAN_IN), .ZN(n6634) );
  OAI222_X1 U7580 ( .A1(n6654), .A2(n6635), .B1(n6634), .B2(n7085), .C1(n6636), 
        .C2(n6655), .ZN(U3190) );
  INV_X1 U7581 ( .A(ADDRESS_REG_7__SCAN_IN), .ZN(n7041) );
  OAI222_X1 U7582 ( .A1(n6654), .A2(n6636), .B1(n7041), .B2(n7085), .C1(n6637), 
        .C2(n6655), .ZN(U3191) );
  INV_X1 U7583 ( .A(ADDRESS_REG_8__SCAN_IN), .ZN(n6976) );
  OAI222_X1 U7584 ( .A1(n6654), .A2(n6637), .B1(n6976), .B2(n7085), .C1(n6638), 
        .C2(n6655), .ZN(U3192) );
  INV_X1 U7585 ( .A(ADDRESS_REG_9__SCAN_IN), .ZN(n6763) );
  OAI222_X1 U7586 ( .A1(n6654), .A2(n6638), .B1(n6763), .B2(n6653), .C1(n6639), 
        .C2(n6655), .ZN(U3193) );
  INV_X1 U7587 ( .A(ADDRESS_REG_10__SCAN_IN), .ZN(n7050) );
  OAI222_X1 U7588 ( .A1(n6654), .A2(n6639), .B1(n7050), .B2(n7085), .C1(n6640), 
        .C2(n6655), .ZN(U3194) );
  INV_X1 U7589 ( .A(ADDRESS_REG_11__SCAN_IN), .ZN(n7059) );
  OAI222_X1 U7590 ( .A1(n6654), .A2(n6640), .B1(n7059), .B2(n6653), .C1(n6642), 
        .C2(n6655), .ZN(U3195) );
  INV_X1 U7591 ( .A(ADDRESS_REG_12__SCAN_IN), .ZN(n6641) );
  OAI222_X1 U7592 ( .A1(n6654), .A2(n6642), .B1(n6641), .B2(n6648), .C1(n6644), 
        .C2(n6655), .ZN(U3196) );
  INV_X1 U7593 ( .A(ADDRESS_REG_13__SCAN_IN), .ZN(n6643) );
  OAI222_X1 U7594 ( .A1(n6654), .A2(n6644), .B1(n6643), .B2(n7085), .C1(n5366), 
        .C2(n6655), .ZN(U3197) );
  INV_X1 U7595 ( .A(ADDRESS_REG_14__SCAN_IN), .ZN(n6645) );
  OAI222_X1 U7596 ( .A1(n6654), .A2(n5366), .B1(n6645), .B2(n6653), .C1(n7038), 
        .C2(n6655), .ZN(U3198) );
  INV_X1 U7597 ( .A(ADDRESS_REG_15__SCAN_IN), .ZN(n7021) );
  OAI222_X1 U7598 ( .A1(n6654), .A2(n7038), .B1(n7021), .B2(n6653), .C1(n6646), 
        .C2(n6655), .ZN(U3199) );
  INV_X1 U7599 ( .A(ADDRESS_REG_16__SCAN_IN), .ZN(n6959) );
  OAI222_X1 U7600 ( .A1(n6655), .A2(n6762), .B1(n6959), .B2(n6653), .C1(n6646), 
        .C2(n6654), .ZN(U3200) );
  INV_X1 U7601 ( .A(REIP_REG_19__SCAN_IN), .ZN(n7031) );
  INV_X1 U7602 ( .A(ADDRESS_REG_17__SCAN_IN), .ZN(n6947) );
  OAI222_X1 U7603 ( .A1(n6655), .A2(n7031), .B1(n6947), .B2(n6653), .C1(n6762), 
        .C2(n6654), .ZN(U3201) );
  INV_X1 U7604 ( .A(ADDRESS_REG_18__SCAN_IN), .ZN(n6647) );
  OAI222_X1 U7605 ( .A1(n6654), .A2(n7031), .B1(n6647), .B2(n6653), .C1(n6773), 
        .C2(n6655), .ZN(U3202) );
  INV_X1 U7606 ( .A(ADDRESS_REG_19__SCAN_IN), .ZN(n6960) );
  OAI222_X1 U7607 ( .A1(n6654), .A2(n6773), .B1(n6960), .B2(n6648), .C1(n6649), 
        .C2(n6655), .ZN(U3203) );
  INV_X1 U7608 ( .A(ADDRESS_REG_20__SCAN_IN), .ZN(n6939) );
  INV_X1 U7609 ( .A(REIP_REG_22__SCAN_IN), .ZN(n6825) );
  OAI222_X1 U7610 ( .A1(n6654), .A2(n6649), .B1(n6939), .B2(n6653), .C1(n6825), 
        .C2(n6655), .ZN(U3204) );
  INV_X1 U7611 ( .A(ADDRESS_REG_21__SCAN_IN), .ZN(n6650) );
  OAI222_X1 U7612 ( .A1(n6654), .A2(n6825), .B1(n6650), .B2(n7085), .C1(n7027), 
        .C2(n6655), .ZN(U3205) );
  INV_X1 U7613 ( .A(ADDRESS_REG_22__SCAN_IN), .ZN(n6970) );
  OAI222_X1 U7614 ( .A1(n6654), .A2(n7027), .B1(n6970), .B2(n6653), .C1(n6962), 
        .C2(n6655), .ZN(U3206) );
  INV_X1 U7615 ( .A(ADDRESS_REG_23__SCAN_IN), .ZN(n6989) );
  OAI222_X1 U7616 ( .A1(n6655), .A2(n6652), .B1(n6989), .B2(n7085), .C1(n6962), 
        .C2(n6654), .ZN(U3207) );
  INV_X1 U7617 ( .A(ADDRESS_REG_24__SCAN_IN), .ZN(n6651) );
  OAI222_X1 U7618 ( .A1(n6654), .A2(n6652), .B1(n6651), .B2(n7085), .C1(n6957), 
        .C2(n6655), .ZN(U3208) );
  INV_X1 U7619 ( .A(ADDRESS_REG_25__SCAN_IN), .ZN(n6988) );
  OAI222_X1 U7620 ( .A1(n6654), .A2(n6957), .B1(n6988), .B2(n7085), .C1(n7009), 
        .C2(n6655), .ZN(U3209) );
  INV_X1 U7621 ( .A(ADDRESS_REG_26__SCAN_IN), .ZN(n6985) );
  OAI222_X1 U7622 ( .A1(n6654), .A2(n7009), .B1(n6985), .B2(n7085), .C1(n7057), 
        .C2(n6655), .ZN(U3210) );
  INV_X1 U7623 ( .A(ADDRESS_REG_27__SCAN_IN), .ZN(n6809) );
  OAI222_X1 U7624 ( .A1(n6654), .A2(n7057), .B1(n6809), .B2(n7085), .C1(n5762), 
        .C2(n6655), .ZN(U3211) );
  INV_X1 U7625 ( .A(ADDRESS_REG_28__SCAN_IN), .ZN(n7044) );
  OAI222_X1 U7626 ( .A1(n6654), .A2(n5762), .B1(n7044), .B2(n6653), .C1(n6975), 
        .C2(n6655), .ZN(U3212) );
  INV_X1 U7627 ( .A(REIP_REG_31__SCAN_IN), .ZN(n6973) );
  INV_X1 U7628 ( .A(ADDRESS_REG_29__SCAN_IN), .ZN(n6853) );
  OAI222_X1 U7629 ( .A1(n6655), .A2(n6973), .B1(n6853), .B2(n7085), .C1(n6975), 
        .C2(n6654), .ZN(U3213) );
  INV_X1 U7630 ( .A(BYTEENABLE_REG_2__SCAN_IN), .ZN(n6839) );
  INV_X1 U7631 ( .A(BE_N_REG_2__SCAN_IN), .ZN(n6784) );
  AOI22_X1 U7632 ( .A1(n7085), .A2(n6839), .B1(n6784), .B2(n7084), .ZN(U3446)
         );
  INV_X1 U7633 ( .A(BE_N_REG_1__SCAN_IN), .ZN(n6813) );
  AOI22_X1 U7634 ( .A1(n7085), .A2(n6656), .B1(n6813), .B2(n7084), .ZN(U3447)
         );
  INV_X1 U7635 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n6674) );
  INV_X1 U7636 ( .A(BE_N_REG_0__SCAN_IN), .ZN(n6838) );
  AOI22_X1 U7637 ( .A1(n7085), .A2(n6674), .B1(n6838), .B2(n7084), .ZN(U3448)
         );
  INV_X1 U7638 ( .A(DATAWIDTH_REG_0__SCAN_IN), .ZN(n7025) );
  INV_X1 U7639 ( .A(n6659), .ZN(n6657) );
  AOI21_X1 U7640 ( .B1(n7025), .B2(n6658), .A(n6657), .ZN(U3451) );
  OAI21_X1 U7641 ( .B1(n6661), .B2(n6660), .A(n6659), .ZN(U3452) );
  INV_X1 U7642 ( .A(n6662), .ZN(n6664) );
  OAI211_X1 U7643 ( .C1(n6666), .C2(n6665), .A(n6664), .B(n6663), .ZN(U3453)
         );
  AOI21_X1 U7644 ( .B1(REIP_REG_0__SCAN_IN), .B2(DATAWIDTH_REG_0__SCAN_IN), 
        .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6668) );
  AOI22_X1 U7645 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_0__SCAN_IN), .B1(
        n6668), .B2(n6667), .ZN(n6669) );
  AOI22_X1 U7646 ( .A1(n6670), .A2(n6669), .B1(n6839), .B2(n6673), .ZN(U3468)
         );
  NOR2_X1 U7647 ( .A1(n6673), .A2(REIP_REG_1__SCAN_IN), .ZN(n6671) );
  AOI22_X1 U7648 ( .A1(n6674), .A2(n6673), .B1(n6672), .B2(n6671), .ZN(U3469)
         );
  INV_X1 U7649 ( .A(W_R_N_REG_SCAN_IN), .ZN(n6793) );
  AOI22_X1 U7650 ( .A1(n7085), .A2(READREQUEST_REG_SCAN_IN), .B1(n6793), .B2(
        n7084), .ZN(U3470) );
  AOI211_X1 U7651 ( .C1(n6333), .C2(n7028), .A(n6676), .B(n6675), .ZN(n6684)
         );
  INV_X1 U7652 ( .A(n6677), .ZN(n6678) );
  OAI211_X1 U7653 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n6679), .A(n6678), .B(
        STATE2_REG_2__SCAN_IN), .ZN(n6681) );
  AOI21_X1 U7654 ( .B1(n6681), .B2(STATE2_REG_0__SCAN_IN), .A(n6680), .ZN(
        n6683) );
  NAND2_X1 U7655 ( .A1(n6684), .A2(REQUESTPENDING_REG_SCAN_IN), .ZN(n6682) );
  OAI21_X1 U7656 ( .B1(n6684), .B2(n6683), .A(n6682), .ZN(U3472) );
  INV_X1 U7657 ( .A(MEMORYFETCH_REG_SCAN_IN), .ZN(n6845) );
  INV_X1 U7658 ( .A(M_IO_N_REG_SCAN_IN), .ZN(n6685) );
  AOI22_X1 U7659 ( .A1(n7085), .A2(n6845), .B1(n6685), .B2(n7084), .ZN(U3473)
         );
  OAI22_X1 U7660 ( .A1(REIP_REG_16__SCAN_IN), .A2(keyinput_g66), .B1(
        keyinput_g12), .B2(DATAI_19_), .ZN(n6686) );
  AOI221_X1 U7661 ( .B1(REIP_REG_16__SCAN_IN), .B2(keyinput_g66), .C1(
        DATAI_19_), .C2(keyinput_g12), .A(n6686), .ZN(n6693) );
  OAI22_X1 U7662 ( .A1(DATAI_18_), .A2(keyinput_g13), .B1(
        ADDRESS_REG_25__SCAN_IN), .B2(keyinput_g75), .ZN(n6687) );
  AOI221_X1 U7663 ( .B1(DATAI_18_), .B2(keyinput_g13), .C1(keyinput_g75), .C2(
        ADDRESS_REG_25__SCAN_IN), .A(n6687), .ZN(n6692) );
  OAI22_X1 U7664 ( .A1(BYTEENABLE_REG_1__SCAN_IN), .A2(keyinput_g48), .B1(
        DATAWIDTH_REG_6__SCAN_IN), .B2(keyinput_g110), .ZN(n6688) );
  AOI221_X1 U7665 ( .B1(BYTEENABLE_REG_1__SCAN_IN), .B2(keyinput_g48), .C1(
        keyinput_g110), .C2(DATAWIDTH_REG_6__SCAN_IN), .A(n6688), .ZN(n6691)
         );
  OAI22_X1 U7666 ( .A1(DATAI_7_), .A2(keyinput_g24), .B1(DATAI_1_), .B2(
        keyinput_g30), .ZN(n6689) );
  AOI221_X1 U7667 ( .B1(DATAI_7_), .B2(keyinput_g24), .C1(keyinput_g30), .C2(
        DATAI_1_), .A(n6689), .ZN(n6690) );
  NAND4_X1 U7668 ( .A1(n6693), .A2(n6692), .A3(n6691), .A4(n6690), .ZN(n6721)
         );
  OAI22_X1 U7669 ( .A1(M_IO_N_REG_SCAN_IN), .A2(keyinput_g40), .B1(
        keyinput_g87), .B2(ADDRESS_REG_13__SCAN_IN), .ZN(n6694) );
  AOI221_X1 U7670 ( .B1(M_IO_N_REG_SCAN_IN), .B2(keyinput_g40), .C1(
        ADDRESS_REG_13__SCAN_IN), .C2(keyinput_g87), .A(n6694), .ZN(n6701) );
  OAI22_X1 U7671 ( .A1(DATAWIDTH_REG_15__SCAN_IN), .A2(keyinput_g119), .B1(
        ADDRESS_REG_11__SCAN_IN), .B2(keyinput_g89), .ZN(n6695) );
  AOI221_X1 U7672 ( .B1(DATAWIDTH_REG_15__SCAN_IN), .B2(keyinput_g119), .C1(
        keyinput_g89), .C2(ADDRESS_REG_11__SCAN_IN), .A(n6695), .ZN(n6700) );
  OAI22_X1 U7673 ( .A1(REIP_REG_28__SCAN_IN), .A2(keyinput_g54), .B1(DATAI_17_), .B2(keyinput_g14), .ZN(n6696) );
  AOI221_X1 U7674 ( .B1(REIP_REG_28__SCAN_IN), .B2(keyinput_g54), .C1(
        keyinput_g14), .C2(DATAI_17_), .A(n6696), .ZN(n6699) );
  OAI22_X1 U7675 ( .A1(REIP_REG_31__SCAN_IN), .A2(keyinput_g51), .B1(
        keyinput_g94), .B2(ADDRESS_REG_6__SCAN_IN), .ZN(n6697) );
  AOI221_X1 U7676 ( .B1(REIP_REG_31__SCAN_IN), .B2(keyinput_g51), .C1(
        ADDRESS_REG_6__SCAN_IN), .C2(keyinput_g94), .A(n6697), .ZN(n6698) );
  NAND4_X1 U7677 ( .A1(n6701), .A2(n6700), .A3(n6699), .A4(n6698), .ZN(n6720)
         );
  OAI22_X1 U7678 ( .A1(DATAI_28_), .A2(keyinput_g3), .B1(keyinput_g85), .B2(
        ADDRESS_REG_15__SCAN_IN), .ZN(n6702) );
  AOI221_X1 U7679 ( .B1(DATAI_28_), .B2(keyinput_g3), .C1(
        ADDRESS_REG_15__SCAN_IN), .C2(keyinput_g85), .A(n6702), .ZN(n6709) );
  OAI22_X1 U7680 ( .A1(ADDRESS_REG_18__SCAN_IN), .A2(keyinput_g82), .B1(
        ADDRESS_REG_16__SCAN_IN), .B2(keyinput_g84), .ZN(n6703) );
  AOI221_X1 U7681 ( .B1(ADDRESS_REG_18__SCAN_IN), .B2(keyinput_g82), .C1(
        keyinput_g84), .C2(ADDRESS_REG_16__SCAN_IN), .A(n6703), .ZN(n6708) );
  OAI22_X1 U7682 ( .A1(READY_N), .A2(keyinput_g35), .B1(keyinput_g105), .B2(
        DATAWIDTH_REG_1__SCAN_IN), .ZN(n6704) );
  AOI221_X1 U7683 ( .B1(READY_N), .B2(keyinput_g35), .C1(
        DATAWIDTH_REG_1__SCAN_IN), .C2(keyinput_g105), .A(n6704), .ZN(n6707)
         );
  OAI22_X1 U7684 ( .A1(DATAWIDTH_REG_7__SCAN_IN), .A2(keyinput_g111), .B1(
        ADDRESS_REG_1__SCAN_IN), .B2(keyinput_g99), .ZN(n6705) );
  AOI221_X1 U7685 ( .B1(DATAWIDTH_REG_7__SCAN_IN), .B2(keyinput_g111), .C1(
        keyinput_g99), .C2(ADDRESS_REG_1__SCAN_IN), .A(n6705), .ZN(n6706) );
  NAND4_X1 U7686 ( .A1(n6709), .A2(n6708), .A3(n6707), .A4(n6706), .ZN(n6719)
         );
  OAI22_X1 U7687 ( .A1(REIP_REG_21__SCAN_IN), .A2(keyinput_g61), .B1(
        keyinput_g120), .B2(DATAWIDTH_REG_16__SCAN_IN), .ZN(n6710) );
  AOI221_X1 U7688 ( .B1(REIP_REG_21__SCAN_IN), .B2(keyinput_g61), .C1(
        DATAWIDTH_REG_16__SCAN_IN), .C2(keyinput_g120), .A(n6710), .ZN(n6717)
         );
  OAI22_X1 U7689 ( .A1(DATAI_23_), .A2(keyinput_g8), .B1(keyinput_g26), .B2(
        DATAI_5_), .ZN(n6711) );
  AOI221_X1 U7690 ( .B1(DATAI_23_), .B2(keyinput_g8), .C1(DATAI_5_), .C2(
        keyinput_g26), .A(n6711), .ZN(n6716) );
  OAI22_X1 U7691 ( .A1(REIP_REG_17__SCAN_IN), .A2(keyinput_g65), .B1(DATAI_3_), 
        .B2(keyinput_g28), .ZN(n6712) );
  AOI221_X1 U7692 ( .B1(REIP_REG_17__SCAN_IN), .B2(keyinput_g65), .C1(
        keyinput_g28), .C2(DATAI_3_), .A(n6712), .ZN(n6715) );
  OAI22_X1 U7693 ( .A1(n7022), .A2(keyinput_g115), .B1(keyinput_g56), .B2(
        REIP_REG_26__SCAN_IN), .ZN(n6713) );
  AOI221_X1 U7694 ( .B1(n7022), .B2(keyinput_g115), .C1(REIP_REG_26__SCAN_IN), 
        .C2(keyinput_g56), .A(n6713), .ZN(n6714) );
  NAND4_X1 U7695 ( .A1(n6717), .A2(n6716), .A3(n6715), .A4(n6714), .ZN(n6718)
         );
  NOR4_X1 U7696 ( .A1(n6721), .A2(n6720), .A3(n6719), .A4(n6718), .ZN(n7083)
         );
  OAI22_X1 U7697 ( .A1(ADDRESS_REG_21__SCAN_IN), .A2(keyinput_g79), .B1(
        ADDRESS_REG_5__SCAN_IN), .B2(keyinput_g95), .ZN(n6722) );
  AOI221_X1 U7698 ( .B1(ADDRESS_REG_21__SCAN_IN), .B2(keyinput_g79), .C1(
        keyinput_g95), .C2(ADDRESS_REG_5__SCAN_IN), .A(n6722), .ZN(n6729) );
  OAI22_X1 U7699 ( .A1(DATAI_14_), .A2(keyinput_g17), .B1(
        DATAWIDTH_REG_3__SCAN_IN), .B2(keyinput_g107), .ZN(n6723) );
  AOI221_X1 U7700 ( .B1(DATAI_14_), .B2(keyinput_g17), .C1(keyinput_g107), 
        .C2(DATAWIDTH_REG_3__SCAN_IN), .A(n6723), .ZN(n6728) );
  OAI22_X1 U7701 ( .A1(ADDRESS_REG_12__SCAN_IN), .A2(keyinput_g88), .B1(
        ADDRESS_REG_14__SCAN_IN), .B2(keyinput_g86), .ZN(n6724) );
  AOI221_X1 U7702 ( .B1(ADDRESS_REG_12__SCAN_IN), .B2(keyinput_g88), .C1(
        keyinput_g86), .C2(ADDRESS_REG_14__SCAN_IN), .A(n6724), .ZN(n6727) );
  OAI22_X1 U7703 ( .A1(DATAI_30_), .A2(keyinput_g1), .B1(keyinput_g44), .B2(
        MORE_REG_SCAN_IN), .ZN(n6725) );
  AOI221_X1 U7704 ( .B1(DATAI_30_), .B2(keyinput_g1), .C1(MORE_REG_SCAN_IN), 
        .C2(keyinput_g44), .A(n6725), .ZN(n6726) );
  NAND4_X1 U7705 ( .A1(n6729), .A2(n6728), .A3(n6727), .A4(n6726), .ZN(n6866)
         );
  OAI22_X1 U7706 ( .A1(ADDRESS_REG_7__SCAN_IN), .A2(keyinput_g93), .B1(
        keyinput_g90), .B2(ADDRESS_REG_10__SCAN_IN), .ZN(n6730) );
  AOI221_X1 U7707 ( .B1(ADDRESS_REG_7__SCAN_IN), .B2(keyinput_g93), .C1(
        ADDRESS_REG_10__SCAN_IN), .C2(keyinput_g90), .A(n6730), .ZN(n6756) );
  OAI22_X1 U7708 ( .A1(DATAI_20_), .A2(keyinput_g11), .B1(keyinput_g33), .B2(
        NA_N), .ZN(n6731) );
  AOI221_X1 U7709 ( .B1(DATAI_20_), .B2(keyinput_g11), .C1(NA_N), .C2(
        keyinput_g33), .A(n6731), .ZN(n6734) );
  OAI22_X1 U7710 ( .A1(REIP_REG_25__SCAN_IN), .A2(keyinput_g57), .B1(DATAI_6_), 
        .B2(keyinput_g25), .ZN(n6732) );
  AOI221_X1 U7711 ( .B1(REIP_REG_25__SCAN_IN), .B2(keyinput_g57), .C1(
        keyinput_g25), .C2(DATAI_6_), .A(n6732), .ZN(n6733) );
  OAI211_X1 U7712 ( .C1(n6736), .C2(keyinput_g102), .A(n6734), .B(n6733), .ZN(
        n6735) );
  AOI21_X1 U7713 ( .B1(n6736), .B2(keyinput_g102), .A(n6735), .ZN(n6755) );
  AOI22_X1 U7714 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(keyinput_g114), .B1(
        DATAI_24_), .B2(keyinput_g7), .ZN(n6737) );
  OAI221_X1 U7715 ( .B1(DATAWIDTH_REG_10__SCAN_IN), .B2(keyinput_g114), .C1(
        DATAI_24_), .C2(keyinput_g7), .A(n6737), .ZN(n6744) );
  AOI22_X1 U7716 ( .A1(ADDRESS_REG_17__SCAN_IN), .A2(keyinput_g83), .B1(
        ADDRESS_REG_24__SCAN_IN), .B2(keyinput_g76), .ZN(n6738) );
  OAI221_X1 U7717 ( .B1(ADDRESS_REG_17__SCAN_IN), .B2(keyinput_g83), .C1(
        ADDRESS_REG_24__SCAN_IN), .C2(keyinput_g76), .A(n6738), .ZN(n6743) );
  AOI22_X1 U7718 ( .A1(ADDRESS_REG_22__SCAN_IN), .A2(keyinput_g78), .B1(
        DATAWIDTH_REG_20__SCAN_IN), .B2(keyinput_g124), .ZN(n6739) );
  OAI221_X1 U7719 ( .B1(ADDRESS_REG_22__SCAN_IN), .B2(keyinput_g78), .C1(
        DATAWIDTH_REG_20__SCAN_IN), .C2(keyinput_g124), .A(n6739), .ZN(n6742)
         );
  AOI22_X1 U7720 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(keyinput_g112), .B1(
        DATAI_10_), .B2(keyinput_g21), .ZN(n6740) );
  OAI221_X1 U7721 ( .B1(DATAWIDTH_REG_8__SCAN_IN), .B2(keyinput_g112), .C1(
        DATAI_10_), .C2(keyinput_g21), .A(n6740), .ZN(n6741) );
  NOR4_X1 U7722 ( .A1(n6744), .A2(n6743), .A3(n6742), .A4(n6741), .ZN(n6754)
         );
  AOI22_X1 U7723 ( .A1(BYTEENABLE_REG_0__SCAN_IN), .A2(keyinput_g47), .B1(
        REIP_REG_30__SCAN_IN), .B2(keyinput_g52), .ZN(n6745) );
  OAI221_X1 U7724 ( .B1(BYTEENABLE_REG_0__SCAN_IN), .B2(keyinput_g47), .C1(
        REIP_REG_30__SCAN_IN), .C2(keyinput_g52), .A(n6745), .ZN(n6752) );
  AOI22_X1 U7725 ( .A1(DATAWIDTH_REG_0__SCAN_IN), .A2(keyinput_g104), .B1(
        DATAWIDTH_REG_9__SCAN_IN), .B2(keyinput_g113), .ZN(n6746) );
  OAI221_X1 U7726 ( .B1(DATAWIDTH_REG_0__SCAN_IN), .B2(keyinput_g104), .C1(
        DATAWIDTH_REG_9__SCAN_IN), .C2(keyinput_g113), .A(n6746), .ZN(n6751)
         );
  AOI22_X1 U7727 ( .A1(ADDRESS_REG_0__SCAN_IN), .A2(keyinput_g100), .B1(
        REIP_REG_24__SCAN_IN), .B2(keyinput_g58), .ZN(n6747) );
  OAI221_X1 U7728 ( .B1(ADDRESS_REG_0__SCAN_IN), .B2(keyinput_g100), .C1(
        REIP_REG_24__SCAN_IN), .C2(keyinput_g58), .A(n6747), .ZN(n6750) );
  AOI22_X1 U7729 ( .A1(BYTEENABLE_REG_3__SCAN_IN), .A2(keyinput_g50), .B1(
        DATAWIDTH_REG_2__SCAN_IN), .B2(keyinput_g106), .ZN(n6748) );
  OAI221_X1 U7730 ( .B1(BYTEENABLE_REG_3__SCAN_IN), .B2(keyinput_g50), .C1(
        DATAWIDTH_REG_2__SCAN_IN), .C2(keyinput_g106), .A(n6748), .ZN(n6749)
         );
  NOR4_X1 U7731 ( .A1(n6752), .A2(n6751), .A3(n6750), .A4(n6749), .ZN(n6753)
         );
  NAND4_X1 U7732 ( .A1(n6756), .A2(n6755), .A3(n6754), .A4(n6753), .ZN(n6865)
         );
  AOI22_X1 U7733 ( .A1(n6976), .A2(keyinput_g92), .B1(keyinput_g122), .B2(
        n6991), .ZN(n6757) );
  OAI221_X1 U7734 ( .B1(n6976), .B2(keyinput_g92), .C1(n6991), .C2(
        keyinput_g122), .A(n6757), .ZN(n6767) );
  INV_X1 U7735 ( .A(DATAI_31_), .ZN(n6956) );
  AOI22_X1 U7736 ( .A1(n6956), .A2(keyinput_g0), .B1(keyinput_g74), .B2(n6985), 
        .ZN(n6758) );
  OAI221_X1 U7737 ( .B1(n6956), .B2(keyinput_g0), .C1(n6985), .C2(keyinput_g74), .A(n6758), .ZN(n6766) );
  INV_X1 U7738 ( .A(DATAI_25_), .ZN(n6942) );
  AOI22_X1 U7739 ( .A1(n6760), .A2(keyinput_g116), .B1(n6942), .B2(keyinput_g6), .ZN(n6759) );
  OAI221_X1 U7740 ( .B1(n6760), .B2(keyinput_g116), .C1(n6942), .C2(
        keyinput_g6), .A(n6759), .ZN(n6765) );
  AOI22_X1 U7741 ( .A1(n6763), .A2(keyinput_g91), .B1(n6762), .B2(keyinput_g64), .ZN(n6761) );
  OAI221_X1 U7742 ( .B1(n6763), .B2(keyinput_g91), .C1(n6762), .C2(
        keyinput_g64), .A(n6761), .ZN(n6764) );
  NOR4_X1 U7743 ( .A1(n6767), .A2(n6766), .A3(n6765), .A4(n6764), .ZN(n6806)
         );
  INV_X1 U7744 ( .A(DATAI_29_), .ZN(n7054) );
  AOI22_X1 U7745 ( .A1(n7054), .A2(keyinput_g2), .B1(keyinput_g20), .B2(n6769), 
        .ZN(n6768) );
  OAI221_X1 U7746 ( .B1(n7054), .B2(keyinput_g2), .C1(n6769), .C2(keyinput_g20), .A(n6768), .ZN(n6778) );
  AOI22_X1 U7747 ( .A1(n7005), .A2(keyinput_g27), .B1(n7015), .B2(keyinput_g19), .ZN(n6770) );
  OAI221_X1 U7748 ( .B1(n7005), .B2(keyinput_g27), .C1(n7015), .C2(
        keyinput_g19), .A(n6770), .ZN(n6777) );
  AOI22_X1 U7749 ( .A1(n6773), .A2(keyinput_g62), .B1(keyinput_g126), .B2(
        n6772), .ZN(n6771) );
  OAI221_X1 U7750 ( .B1(n6773), .B2(keyinput_g62), .C1(n6772), .C2(
        keyinput_g126), .A(n6771), .ZN(n6776) );
  INV_X1 U7751 ( .A(CODEFETCH_REG_SCAN_IN), .ZN(n7043) );
  AOI22_X1 U7752 ( .A1(n7008), .A2(keyinput_g125), .B1(n7043), .B2(
        keyinput_g39), .ZN(n6774) );
  OAI221_X1 U7753 ( .B1(n7008), .B2(keyinput_g125), .C1(n7043), .C2(
        keyinput_g39), .A(n6774), .ZN(n6775) );
  NOR4_X1 U7754 ( .A1(n6778), .A2(n6777), .A3(n6776), .A4(n6775), .ZN(n6805)
         );
  INV_X1 U7755 ( .A(DATAI_16_), .ZN(n6780) );
  AOI22_X1 U7756 ( .A1(n6780), .A2(keyinput_g15), .B1(n6112), .B2(keyinput_g9), 
        .ZN(n6779) );
  OAI221_X1 U7757 ( .B1(n6780), .B2(keyinput_g15), .C1(n6112), .C2(keyinput_g9), .A(n6779), .ZN(n6790) );
  AOI22_X1 U7758 ( .A1(n6782), .A2(keyinput_g127), .B1(n7014), .B2(
        keyinput_g29), .ZN(n6781) );
  OAI221_X1 U7759 ( .B1(n6782), .B2(keyinput_g127), .C1(n7014), .C2(
        keyinput_g29), .A(n6781), .ZN(n6789) );
  AOI22_X1 U7760 ( .A1(n6785), .A2(keyinput_g36), .B1(n6784), .B2(keyinput_g68), .ZN(n6783) );
  OAI221_X1 U7761 ( .B1(n6785), .B2(keyinput_g36), .C1(n6784), .C2(
        keyinput_g68), .A(n6783), .ZN(n6788) );
  INV_X1 U7762 ( .A(DATAI_26_), .ZN(n6979) );
  AOI22_X1 U7763 ( .A1(n7060), .A2(keyinput_g38), .B1(n6979), .B2(keyinput_g5), 
        .ZN(n6786) );
  OAI221_X1 U7764 ( .B1(n7060), .B2(keyinput_g38), .C1(n6979), .C2(keyinput_g5), .A(n6786), .ZN(n6787) );
  NOR4_X1 U7765 ( .A1(n6790), .A2(n6789), .A3(n6788), .A4(n6787), .ZN(n6804)
         );
  INV_X1 U7766 ( .A(BS16_N), .ZN(n6792) );
  AOI22_X1 U7767 ( .A1(n6793), .A2(keyinput_g46), .B1(keyinput_g34), .B2(n6792), .ZN(n6791) );
  OAI221_X1 U7768 ( .B1(n6793), .B2(keyinput_g46), .C1(n6792), .C2(
        keyinput_g34), .A(n6791), .ZN(n6802) );
  AOI22_X1 U7769 ( .A1(n7009), .A2(keyinput_g55), .B1(keyinput_g16), .B2(n6795), .ZN(n6794) );
  OAI221_X1 U7770 ( .B1(n7009), .B2(keyinput_g55), .C1(n6795), .C2(
        keyinput_g16), .A(n6794), .ZN(n6801) );
  INV_X1 U7771 ( .A(DATAI_21_), .ZN(n7006) );
  AOI22_X1 U7772 ( .A1(n7006), .A2(keyinput_g10), .B1(keyinput_g41), .B2(n6948), .ZN(n6796) );
  OAI221_X1 U7773 ( .B1(n7006), .B2(keyinput_g10), .C1(n6948), .C2(
        keyinput_g41), .A(n6796), .ZN(n6800) );
  AOI22_X1 U7774 ( .A1(n6798), .A2(keyinput_g109), .B1(keyinput_g77), .B2(
        n6989), .ZN(n6797) );
  OAI221_X1 U7775 ( .B1(n6798), .B2(keyinput_g109), .C1(n6989), .C2(
        keyinput_g77), .A(n6797), .ZN(n6799) );
  NOR4_X1 U7776 ( .A1(n6802), .A2(n6801), .A3(n6800), .A4(n6799), .ZN(n6803)
         );
  NAND4_X1 U7777 ( .A1(n6806), .A2(n6805), .A3(n6804), .A4(n6803), .ZN(n6864)
         );
  AOI22_X1 U7778 ( .A1(n6809), .A2(keyinput_g73), .B1(n6808), .B2(keyinput_g42), .ZN(n6807) );
  OAI221_X1 U7779 ( .B1(n6809), .B2(keyinput_g73), .C1(n6808), .C2(
        keyinput_g42), .A(n6807), .ZN(n6820) );
  AOI22_X1 U7780 ( .A1(n5762), .A2(keyinput_g53), .B1(keyinput_g23), .B2(n6811), .ZN(n6810) );
  OAI221_X1 U7781 ( .B1(n5762), .B2(keyinput_g53), .C1(n6811), .C2(
        keyinput_g23), .A(n6810), .ZN(n6819) );
  AOI22_X1 U7782 ( .A1(n6814), .A2(keyinput_g118), .B1(n6813), .B2(
        keyinput_g69), .ZN(n6812) );
  OAI221_X1 U7783 ( .B1(n6814), .B2(keyinput_g118), .C1(n6813), .C2(
        keyinput_g69), .A(n6812), .ZN(n6818) );
  INV_X1 U7784 ( .A(DATAI_27_), .ZN(n6963) );
  INV_X1 U7785 ( .A(BE_N_REG_3__SCAN_IN), .ZN(n6816) );
  AOI22_X1 U7786 ( .A1(n6963), .A2(keyinput_g4), .B1(keyinput_g67), .B2(n6816), 
        .ZN(n6815) );
  OAI221_X1 U7787 ( .B1(n6963), .B2(keyinput_g4), .C1(n6816), .C2(keyinput_g67), .A(n6815), .ZN(n6817) );
  NOR4_X1 U7788 ( .A1(n6820), .A2(n6819), .A3(n6818), .A4(n6817), .ZN(n6862)
         );
  AOI22_X1 U7789 ( .A1(n7044), .A2(keyinput_g72), .B1(n7027), .B2(keyinput_g59), .ZN(n6821) );
  OAI221_X1 U7790 ( .B1(n7044), .B2(keyinput_g72), .C1(n7027), .C2(
        keyinput_g59), .A(n6821), .ZN(n6831) );
  AOI22_X1 U7791 ( .A1(n6823), .A2(keyinput_g98), .B1(n7031), .B2(keyinput_g63), .ZN(n6822) );
  OAI221_X1 U7792 ( .B1(n6823), .B2(keyinput_g98), .C1(n7031), .C2(
        keyinput_g63), .A(n6822), .ZN(n6830) );
  AOI22_X1 U7793 ( .A1(n6825), .A2(keyinput_g60), .B1(keyinput_g108), .B2(
        n7053), .ZN(n6824) );
  OAI221_X1 U7794 ( .B1(n6825), .B2(keyinput_g60), .C1(n7053), .C2(
        keyinput_g108), .A(n6824), .ZN(n6829) );
  INV_X1 U7795 ( .A(READREQUEST_REG_SCAN_IN), .ZN(n6827) );
  AOI22_X1 U7796 ( .A1(n7051), .A2(keyinput_g123), .B1(n6827), .B2(
        keyinput_g37), .ZN(n6826) );
  OAI221_X1 U7797 ( .B1(n7051), .B2(keyinput_g123), .C1(n6827), .C2(
        keyinput_g37), .A(n6826), .ZN(n6828) );
  NOR4_X1 U7798 ( .A1(n6831), .A2(n6830), .A3(n6829), .A4(n6828), .ZN(n6861)
         );
  AOI22_X1 U7799 ( .A1(n6833), .A2(keyinput_g97), .B1(n7056), .B2(keyinput_g43), .ZN(n6832) );
  OAI221_X1 U7800 ( .B1(n6833), .B2(keyinput_g97), .C1(n7056), .C2(
        keyinput_g43), .A(n6832), .ZN(n6843) );
  AOI22_X1 U7801 ( .A1(n6939), .A2(keyinput_g80), .B1(n6835), .B2(keyinput_g96), .ZN(n6834) );
  OAI221_X1 U7802 ( .B1(n6939), .B2(keyinput_g80), .C1(n6835), .C2(
        keyinput_g96), .A(n6834), .ZN(n6842) );
  AOI22_X1 U7803 ( .A1(n7040), .A2(keyinput_g101), .B1(keyinput_g31), .B2(
        n6945), .ZN(n6836) );
  OAI221_X1 U7804 ( .B1(n7040), .B2(keyinput_g101), .C1(n6945), .C2(
        keyinput_g31), .A(n6836), .ZN(n6841) );
  AOI22_X1 U7805 ( .A1(n6839), .A2(keyinput_g49), .B1(keyinput_g70), .B2(n6838), .ZN(n6837) );
  OAI221_X1 U7806 ( .B1(n6839), .B2(keyinput_g49), .C1(n6838), .C2(
        keyinput_g70), .A(n6837), .ZN(n6840) );
  NOR4_X1 U7807 ( .A1(n6843), .A2(n6842), .A3(n6841), .A4(n6840), .ZN(n6860)
         );
  AOI22_X1 U7808 ( .A1(n6846), .A2(keyinput_g22), .B1(keyinput_g32), .B2(n6845), .ZN(n6844) );
  OAI221_X1 U7809 ( .B1(n6846), .B2(keyinput_g22), .C1(n6845), .C2(
        keyinput_g32), .A(n6844), .ZN(n6858) );
  AOI22_X1 U7810 ( .A1(n6849), .A2(keyinput_g121), .B1(n6848), .B2(
        keyinput_g18), .ZN(n6847) );
  OAI221_X1 U7811 ( .B1(n6849), .B2(keyinput_g121), .C1(n6848), .C2(
        keyinput_g18), .A(n6847), .ZN(n6857) );
  AOI22_X1 U7812 ( .A1(n6851), .A2(keyinput_g117), .B1(keyinput_g81), .B2(
        n6960), .ZN(n6850) );
  OAI221_X1 U7813 ( .B1(n6851), .B2(keyinput_g117), .C1(n6960), .C2(
        keyinput_g81), .A(n6850), .ZN(n6856) );
  AOI22_X1 U7814 ( .A1(n6854), .A2(keyinput_g103), .B1(keyinput_g71), .B2(
        n6853), .ZN(n6852) );
  OAI221_X1 U7815 ( .B1(n6854), .B2(keyinput_g103), .C1(n6853), .C2(
        keyinput_g71), .A(n6852), .ZN(n6855) );
  NOR4_X1 U7816 ( .A1(n6858), .A2(n6857), .A3(n6856), .A4(n6855), .ZN(n6859)
         );
  NAND4_X1 U7817 ( .A1(n6862), .A2(n6861), .A3(n6860), .A4(n6859), .ZN(n6863)
         );
  NOR4_X1 U7818 ( .A1(n6866), .A2(n6865), .A3(n6864), .A4(n6863), .ZN(n7082)
         );
  AOI22_X1 U7819 ( .A1(keyinput_f118), .A2(DATAWIDTH_REG_14__SCAN_IN), .B1(
        REIP_REG_18__SCAN_IN), .B2(keyinput_f64), .ZN(n6867) );
  OAI221_X1 U7820 ( .B1(keyinput_f118), .B2(DATAWIDTH_REG_14__SCAN_IN), .C1(
        REIP_REG_18__SCAN_IN), .C2(keyinput_f64), .A(n6867), .ZN(n6874) );
  AOI22_X1 U7821 ( .A1(DATAI_6_), .A2(keyinput_f25), .B1(DATAI_14_), .B2(
        keyinput_f17), .ZN(n6868) );
  OAI221_X1 U7822 ( .B1(DATAI_6_), .B2(keyinput_f25), .C1(DATAI_14_), .C2(
        keyinput_f17), .A(n6868), .ZN(n6873) );
  AOI22_X1 U7823 ( .A1(keyinput_f82), .A2(ADDRESS_REG_18__SCAN_IN), .B1(
        REQUESTPENDING_REG_SCAN_IN), .B2(keyinput_f42), .ZN(n6869) );
  OAI221_X1 U7824 ( .B1(keyinput_f82), .B2(ADDRESS_REG_18__SCAN_IN), .C1(
        REQUESTPENDING_REG_SCAN_IN), .C2(keyinput_f42), .A(n6869), .ZN(n6872)
         );
  AOI22_X1 U7825 ( .A1(keyinput_f109), .A2(DATAWIDTH_REG_5__SCAN_IN), .B1(
        DATAI_30_), .B2(keyinput_f1), .ZN(n6870) );
  OAI221_X1 U7826 ( .B1(keyinput_f109), .B2(DATAWIDTH_REG_5__SCAN_IN), .C1(
        DATAI_30_), .C2(keyinput_f1), .A(n6870), .ZN(n6871) );
  NOR4_X1 U7827 ( .A1(n6874), .A2(n6873), .A3(n6872), .A4(n6871), .ZN(n7075)
         );
  AOI22_X1 U7828 ( .A1(keyinput_f69), .A2(BE_N_REG_1__SCAN_IN), .B1(
        keyinput_f49), .B2(BYTEENABLE_REG_2__SCAN_IN), .ZN(n6875) );
  OAI221_X1 U7829 ( .B1(keyinput_f69), .B2(BE_N_REG_1__SCAN_IN), .C1(
        keyinput_f49), .C2(BYTEENABLE_REG_2__SCAN_IN), .A(n6875), .ZN(n6901)
         );
  OAI22_X1 U7830 ( .A1(REIP_REG_21__SCAN_IN), .A2(keyinput_f61), .B1(
        keyinput_f73), .B2(ADDRESS_REG_27__SCAN_IN), .ZN(n6876) );
  AOI221_X1 U7831 ( .B1(REIP_REG_21__SCAN_IN), .B2(keyinput_f61), .C1(
        ADDRESS_REG_27__SCAN_IN), .C2(keyinput_f73), .A(n6876), .ZN(n6880) );
  AOI22_X1 U7832 ( .A1(MEMORYFETCH_REG_SCAN_IN), .A2(keyinput_f32), .B1(
        DATAI_11_), .B2(keyinput_f20), .ZN(n6877) );
  OAI221_X1 U7833 ( .B1(MEMORYFETCH_REG_SCAN_IN), .B2(keyinput_f32), .C1(
        DATAI_11_), .C2(keyinput_f20), .A(n6877), .ZN(n6878) );
  AOI21_X1 U7834 ( .B1(keyinput_f26), .B2(n6881), .A(n6878), .ZN(n6879) );
  OAI211_X1 U7835 ( .C1(keyinput_f26), .C2(n6881), .A(n6880), .B(n6879), .ZN(
        n6900) );
  OAI22_X1 U7836 ( .A1(keyinput_f91), .A2(ADDRESS_REG_9__SCAN_IN), .B1(
        keyinput_f98), .B2(ADDRESS_REG_2__SCAN_IN), .ZN(n6882) );
  AOI221_X1 U7837 ( .B1(keyinput_f91), .B2(ADDRESS_REG_9__SCAN_IN), .C1(
        ADDRESS_REG_2__SCAN_IN), .C2(keyinput_f98), .A(n6882), .ZN(n6889) );
  OAI22_X1 U7838 ( .A1(keyinput_f71), .A2(ADDRESS_REG_29__SCAN_IN), .B1(
        keyinput_f94), .B2(ADDRESS_REG_6__SCAN_IN), .ZN(n6883) );
  AOI221_X1 U7839 ( .B1(keyinput_f71), .B2(ADDRESS_REG_29__SCAN_IN), .C1(
        ADDRESS_REG_6__SCAN_IN), .C2(keyinput_f94), .A(n6883), .ZN(n6888) );
  OAI22_X1 U7840 ( .A1(keyinput_f106), .A2(DATAWIDTH_REG_2__SCAN_IN), .B1(
        keyinput_f67), .B2(BE_N_REG_3__SCAN_IN), .ZN(n6884) );
  AOI221_X1 U7841 ( .B1(keyinput_f106), .B2(DATAWIDTH_REG_2__SCAN_IN), .C1(
        BE_N_REG_3__SCAN_IN), .C2(keyinput_f67), .A(n6884), .ZN(n6887) );
  OAI22_X1 U7842 ( .A1(REIP_REG_20__SCAN_IN), .A2(keyinput_f62), .B1(
        keyinput_f11), .B2(DATAI_20_), .ZN(n6885) );
  AOI221_X1 U7843 ( .B1(REIP_REG_20__SCAN_IN), .B2(keyinput_f62), .C1(
        DATAI_20_), .C2(keyinput_f11), .A(n6885), .ZN(n6886) );
  NAND4_X1 U7844 ( .A1(n6889), .A2(n6888), .A3(n6887), .A4(n6886), .ZN(n6899)
         );
  OAI22_X1 U7845 ( .A1(STATE_REG_0__SCAN_IN), .A2(keyinput_f103), .B1(
        STATE_REG_1__SCAN_IN), .B2(keyinput_f102), .ZN(n6890) );
  AOI221_X1 U7846 ( .B1(STATE_REG_0__SCAN_IN), .B2(keyinput_f103), .C1(
        keyinput_f102), .C2(STATE_REG_1__SCAN_IN), .A(n6890), .ZN(n6897) );
  OAI22_X1 U7847 ( .A1(DATAI_16_), .A2(keyinput_f15), .B1(keyinput_f111), .B2(
        DATAWIDTH_REG_7__SCAN_IN), .ZN(n6891) );
  AOI221_X1 U7848 ( .B1(DATAI_16_), .B2(keyinput_f15), .C1(
        DATAWIDTH_REG_7__SCAN_IN), .C2(keyinput_f111), .A(n6891), .ZN(n6896)
         );
  OAI22_X1 U7849 ( .A1(keyinput_f68), .A2(BE_N_REG_2__SCAN_IN), .B1(
        keyinput_f99), .B2(ADDRESS_REG_1__SCAN_IN), .ZN(n6892) );
  AOI221_X1 U7850 ( .B1(keyinput_f68), .B2(BE_N_REG_2__SCAN_IN), .C1(
        ADDRESS_REG_1__SCAN_IN), .C2(keyinput_f99), .A(n6892), .ZN(n6895) );
  OAI22_X1 U7851 ( .A1(keyinput_f48), .A2(BYTEENABLE_REG_1__SCAN_IN), .B1(
        keyinput_f76), .B2(ADDRESS_REG_24__SCAN_IN), .ZN(n6893) );
  AOI221_X1 U7852 ( .B1(keyinput_f48), .B2(BYTEENABLE_REG_1__SCAN_IN), .C1(
        ADDRESS_REG_24__SCAN_IN), .C2(keyinput_f76), .A(n6893), .ZN(n6894) );
  NAND4_X1 U7853 ( .A1(n6897), .A2(n6896), .A3(n6895), .A4(n6894), .ZN(n6898)
         );
  NOR4_X1 U7854 ( .A1(n6901), .A2(n6900), .A3(n6899), .A4(n6898), .ZN(n7074)
         );
  OAI22_X1 U7855 ( .A1(REIP_REG_17__SCAN_IN), .A2(keyinput_f65), .B1(
        BE_N_REG_0__SCAN_IN), .B2(keyinput_f70), .ZN(n6902) );
  AOI221_X1 U7856 ( .B1(REIP_REG_17__SCAN_IN), .B2(keyinput_f65), .C1(
        keyinput_f70), .C2(BE_N_REG_0__SCAN_IN), .A(n6902), .ZN(n6909) );
  OAI22_X1 U7857 ( .A1(REIP_REG_22__SCAN_IN), .A2(keyinput_f60), .B1(
        keyinput_f37), .B2(READREQUEST_REG_SCAN_IN), .ZN(n6903) );
  AOI221_X1 U7858 ( .B1(REIP_REG_22__SCAN_IN), .B2(keyinput_f60), .C1(
        READREQUEST_REG_SCAN_IN), .C2(keyinput_f37), .A(n6903), .ZN(n6908) );
  OAI22_X1 U7859 ( .A1(DATAI_22_), .A2(keyinput_f9), .B1(
        DATAWIDTH_REG_22__SCAN_IN), .B2(keyinput_f126), .ZN(n6904) );
  AOI221_X1 U7860 ( .B1(DATAI_22_), .B2(keyinput_f9), .C1(keyinput_f126), .C2(
        DATAWIDTH_REG_22__SCAN_IN), .A(n6904), .ZN(n6907) );
  OAI22_X1 U7861 ( .A1(keyinput_f79), .A2(ADDRESS_REG_21__SCAN_IN), .B1(
        keyinput_f40), .B2(M_IO_N_REG_SCAN_IN), .ZN(n6905) );
  AOI221_X1 U7862 ( .B1(keyinput_f79), .B2(ADDRESS_REG_21__SCAN_IN), .C1(
        M_IO_N_REG_SCAN_IN), .C2(keyinput_f40), .A(n6905), .ZN(n6906) );
  NAND4_X1 U7863 ( .A1(n6909), .A2(n6908), .A3(n6907), .A4(n6906), .ZN(n6937)
         );
  OAI22_X1 U7864 ( .A1(keyinput_f116), .A2(DATAWIDTH_REG_12__SCAN_IN), .B1(
        keyinput_f87), .B2(ADDRESS_REG_13__SCAN_IN), .ZN(n6910) );
  AOI221_X1 U7865 ( .B1(keyinput_f116), .B2(DATAWIDTH_REG_12__SCAN_IN), .C1(
        ADDRESS_REG_13__SCAN_IN), .C2(keyinput_f87), .A(n6910), .ZN(n6917) );
  OAI22_X1 U7866 ( .A1(DATAI_10_), .A2(keyinput_f21), .B1(keyinput_f24), .B2(
        DATAI_7_), .ZN(n6911) );
  AOI221_X1 U7867 ( .B1(DATAI_10_), .B2(keyinput_f21), .C1(DATAI_7_), .C2(
        keyinput_f24), .A(n6911), .ZN(n6916) );
  OAI22_X1 U7868 ( .A1(REIP_REG_25__SCAN_IN), .A2(keyinput_f57), .B1(
        keyinput_f96), .B2(ADDRESS_REG_4__SCAN_IN), .ZN(n6912) );
  AOI221_X1 U7869 ( .B1(REIP_REG_25__SCAN_IN), .B2(keyinput_f57), .C1(
        ADDRESS_REG_4__SCAN_IN), .C2(keyinput_f96), .A(n6912), .ZN(n6915) );
  OAI22_X1 U7870 ( .A1(keyinput_f113), .A2(DATAWIDTH_REG_9__SCAN_IN), .B1(
        keyinput_f97), .B2(ADDRESS_REG_3__SCAN_IN), .ZN(n6913) );
  AOI221_X1 U7871 ( .B1(keyinput_f113), .B2(DATAWIDTH_REG_9__SCAN_IN), .C1(
        ADDRESS_REG_3__SCAN_IN), .C2(keyinput_f97), .A(n6913), .ZN(n6914) );
  NAND4_X1 U7872 ( .A1(n6917), .A2(n6916), .A3(n6915), .A4(n6914), .ZN(n6936)
         );
  OAI22_X1 U7873 ( .A1(DATAI_8_), .A2(keyinput_f23), .B1(
        DATAWIDTH_REG_10__SCAN_IN), .B2(keyinput_f114), .ZN(n6918) );
  AOI221_X1 U7874 ( .B1(DATAI_8_), .B2(keyinput_f23), .C1(keyinput_f114), .C2(
        DATAWIDTH_REG_10__SCAN_IN), .A(n6918), .ZN(n6925) );
  OAI22_X1 U7875 ( .A1(DATAI_18_), .A2(keyinput_f13), .B1(keyinput_f46), .B2(
        W_R_N_REG_SCAN_IN), .ZN(n6919) );
  AOI221_X1 U7876 ( .B1(DATAI_18_), .B2(keyinput_f13), .C1(W_R_N_REG_SCAN_IN), 
        .C2(keyinput_f46), .A(n6919), .ZN(n6924) );
  OAI22_X1 U7877 ( .A1(keyinput_f120), .A2(DATAWIDTH_REG_16__SCAN_IN), .B1(
        keyinput_f95), .B2(ADDRESS_REG_5__SCAN_IN), .ZN(n6920) );
  AOI221_X1 U7878 ( .B1(keyinput_f120), .B2(DATAWIDTH_REG_16__SCAN_IN), .C1(
        ADDRESS_REG_5__SCAN_IN), .C2(keyinput_f95), .A(n6920), .ZN(n6923) );
  OAI22_X1 U7879 ( .A1(DATAI_13_), .A2(keyinput_f18), .B1(keyinput_f47), .B2(
        BYTEENABLE_REG_0__SCAN_IN), .ZN(n6921) );
  AOI221_X1 U7880 ( .B1(DATAI_13_), .B2(keyinput_f18), .C1(
        BYTEENABLE_REG_0__SCAN_IN), .C2(keyinput_f47), .A(n6921), .ZN(n6922)
         );
  NAND4_X1 U7881 ( .A1(n6925), .A2(n6924), .A3(n6923), .A4(n6922), .ZN(n6935)
         );
  OAI22_X1 U7882 ( .A1(keyinput_f117), .A2(DATAWIDTH_REG_13__SCAN_IN), .B1(
        keyinput_f107), .B2(DATAWIDTH_REG_3__SCAN_IN), .ZN(n6926) );
  AOI221_X1 U7883 ( .B1(keyinput_f117), .B2(DATAWIDTH_REG_13__SCAN_IN), .C1(
        DATAWIDTH_REG_3__SCAN_IN), .C2(keyinput_f107), .A(n6926), .ZN(n6933)
         );
  OAI22_X1 U7884 ( .A1(DATAI_15_), .A2(keyinput_f16), .B1(
        ADDRESS_REG_12__SCAN_IN), .B2(keyinput_f88), .ZN(n6927) );
  AOI221_X1 U7885 ( .B1(DATAI_15_), .B2(keyinput_f16), .C1(keyinput_f88), .C2(
        ADDRESS_REG_12__SCAN_IN), .A(n6927), .ZN(n6932) );
  OAI22_X1 U7886 ( .A1(DATAI_9_), .A2(keyinput_f22), .B1(
        ADDRESS_REG_14__SCAN_IN), .B2(keyinput_f86), .ZN(n6928) );
  AOI221_X1 U7887 ( .B1(DATAI_9_), .B2(keyinput_f22), .C1(keyinput_f86), .C2(
        ADDRESS_REG_14__SCAN_IN), .A(n6928), .ZN(n6931) );
  OAI22_X1 U7888 ( .A1(DATAI_19_), .A2(keyinput_f12), .B1(keyinput_f14), .B2(
        DATAI_17_), .ZN(n6929) );
  AOI221_X1 U7889 ( .B1(DATAI_19_), .B2(keyinput_f12), .C1(DATAI_17_), .C2(
        keyinput_f14), .A(n6929), .ZN(n6930) );
  NAND4_X1 U7890 ( .A1(n6933), .A2(n6932), .A3(n6931), .A4(n6930), .ZN(n6934)
         );
  NOR4_X1 U7891 ( .A1(n6937), .A2(n6936), .A3(n6935), .A4(n6934), .ZN(n7073)
         );
  AOI22_X1 U7892 ( .A1(HOLD), .A2(keyinput_f36), .B1(n6939), .B2(keyinput_f80), 
        .ZN(n6938) );
  OAI221_X1 U7893 ( .B1(HOLD), .B2(keyinput_f36), .C1(n6939), .C2(keyinput_f80), .A(n6938), .ZN(n6952) );
  INV_X1 U7894 ( .A(keyinput_f124), .ZN(n6941) );
  AOI22_X1 U7895 ( .A1(n6942), .A2(keyinput_f6), .B1(DATAWIDTH_REG_20__SCAN_IN), .B2(n6941), .ZN(n6940) );
  OAI221_X1 U7896 ( .B1(n6942), .B2(keyinput_f6), .C1(n6941), .C2(
        DATAWIDTH_REG_20__SCAN_IN), .A(n6940), .ZN(n6951) );
  INV_X1 U7897 ( .A(DATAI_23_), .ZN(n6944) );
  AOI22_X1 U7898 ( .A1(n6945), .A2(keyinput_f31), .B1(n6944), .B2(keyinput_f8), 
        .ZN(n6943) );
  OAI221_X1 U7899 ( .B1(n6945), .B2(keyinput_f31), .C1(n6944), .C2(keyinput_f8), .A(n6943), .ZN(n6950) );
  AOI22_X1 U7900 ( .A1(n6948), .A2(keyinput_f41), .B1(keyinput_f83), .B2(n6947), .ZN(n6946) );
  OAI221_X1 U7901 ( .B1(n6948), .B2(keyinput_f41), .C1(n6947), .C2(
        keyinput_f83), .A(n6946), .ZN(n6949) );
  NOR4_X1 U7902 ( .A1(n6952), .A2(n6951), .A3(n6950), .A4(n6949), .ZN(n7003)
         );
  AOI22_X1 U7903 ( .A1(n5762), .A2(keyinput_f53), .B1(keyinput_f112), .B2(
        n6954), .ZN(n6953) );
  OAI221_X1 U7904 ( .B1(n5762), .B2(keyinput_f53), .C1(n6954), .C2(
        keyinput_f112), .A(n6953), .ZN(n6967) );
  AOI22_X1 U7905 ( .A1(n6957), .A2(keyinput_f56), .B1(keyinput_f0), .B2(n6956), 
        .ZN(n6955) );
  OAI221_X1 U7906 ( .B1(n6957), .B2(keyinput_f56), .C1(n6956), .C2(keyinput_f0), .A(n6955), .ZN(n6966) );
  AOI22_X1 U7907 ( .A1(n6960), .A2(keyinput_f81), .B1(keyinput_f84), .B2(n6959), .ZN(n6958) );
  OAI221_X1 U7908 ( .B1(n6960), .B2(keyinput_f81), .C1(n6959), .C2(
        keyinput_f84), .A(n6958), .ZN(n6965) );
  AOI22_X1 U7909 ( .A1(n6963), .A2(keyinput_f4), .B1(n6962), .B2(keyinput_f58), 
        .ZN(n6961) );
  OAI221_X1 U7910 ( .B1(n6963), .B2(keyinput_f4), .C1(n6962), .C2(keyinput_f58), .A(n6961), .ZN(n6964) );
  NOR4_X1 U7911 ( .A1(n6967), .A2(n6966), .A3(n6965), .A4(n6964), .ZN(n7002)
         );
  INV_X1 U7912 ( .A(DATAI_24_), .ZN(n6969) );
  AOI22_X1 U7913 ( .A1(n6970), .A2(keyinput_f78), .B1(n6969), .B2(keyinput_f7), 
        .ZN(n6968) );
  OAI221_X1 U7914 ( .B1(n6970), .B2(keyinput_f78), .C1(n6969), .C2(keyinput_f7), .A(n6968), .ZN(n6983) );
  INV_X1 U7915 ( .A(keyinput_f121), .ZN(n6972) );
  AOI22_X1 U7916 ( .A1(n6973), .A2(keyinput_f51), .B1(
        DATAWIDTH_REG_17__SCAN_IN), .B2(n6972), .ZN(n6971) );
  OAI221_X1 U7917 ( .B1(n6973), .B2(keyinput_f51), .C1(n6972), .C2(
        DATAWIDTH_REG_17__SCAN_IN), .A(n6971), .ZN(n6982) );
  AOI22_X1 U7918 ( .A1(n6976), .A2(keyinput_f92), .B1(n6975), .B2(keyinput_f52), .ZN(n6974) );
  OAI221_X1 U7919 ( .B1(n6976), .B2(keyinput_f92), .C1(n6975), .C2(
        keyinput_f52), .A(n6974), .ZN(n6981) );
  AOI22_X1 U7920 ( .A1(n6979), .A2(keyinput_f5), .B1(keyinput_f50), .B2(n6978), 
        .ZN(n6977) );
  OAI221_X1 U7921 ( .B1(n6979), .B2(keyinput_f5), .C1(n6978), .C2(keyinput_f50), .A(n6977), .ZN(n6980) );
  NOR4_X1 U7922 ( .A1(n6983), .A2(n6982), .A3(n6981), .A4(n6980), .ZN(n7001)
         );
  AOI22_X1 U7923 ( .A1(n6986), .A2(keyinput_f28), .B1(keyinput_f74), .B2(n6985), .ZN(n6984) );
  OAI221_X1 U7924 ( .B1(n6986), .B2(keyinput_f28), .C1(n6985), .C2(
        keyinput_f74), .A(n6984), .ZN(n6999) );
  AOI22_X1 U7925 ( .A1(n6989), .A2(keyinput_f77), .B1(keyinput_f75), .B2(n6988), .ZN(n6987) );
  OAI221_X1 U7926 ( .B1(n6989), .B2(keyinput_f77), .C1(n6988), .C2(
        keyinput_f75), .A(n6987), .ZN(n6998) );
  INV_X1 U7927 ( .A(DATAI_28_), .ZN(n6992) );
  AOI22_X1 U7928 ( .A1(n6992), .A2(keyinput_f3), .B1(keyinput_f122), .B2(n6991), .ZN(n6990) );
  OAI221_X1 U7929 ( .B1(n6992), .B2(keyinput_f3), .C1(n6991), .C2(
        keyinput_f122), .A(n6990), .ZN(n6997) );
  INV_X1 U7930 ( .A(keyinput_f119), .ZN(n6994) );
  AOI22_X1 U7931 ( .A1(n6995), .A2(keyinput_f30), .B1(
        DATAWIDTH_REG_15__SCAN_IN), .B2(n6994), .ZN(n6993) );
  OAI221_X1 U7932 ( .B1(n6995), .B2(keyinput_f30), .C1(n6994), .C2(
        DATAWIDTH_REG_15__SCAN_IN), .A(n6993), .ZN(n6996) );
  NOR4_X1 U7933 ( .A1(n6999), .A2(n6998), .A3(n6997), .A4(n6996), .ZN(n7000)
         );
  NAND4_X1 U7934 ( .A1(n7003), .A2(n7002), .A3(n7001), .A4(n7000), .ZN(n7071)
         );
  OAI22_X1 U7935 ( .A1(n7006), .A2(keyinput_f10), .B1(n7005), .B2(keyinput_f27), .ZN(n7004) );
  AOI221_X1 U7936 ( .B1(n7006), .B2(keyinput_f10), .C1(keyinput_f27), .C2(
        n7005), .A(n7004), .ZN(n7019) );
  OAI22_X1 U7937 ( .A1(n7009), .A2(keyinput_f55), .B1(n7008), .B2(
        keyinput_f125), .ZN(n7007) );
  AOI221_X1 U7938 ( .B1(n7009), .B2(keyinput_f55), .C1(keyinput_f125), .C2(
        n7008), .A(n7007), .ZN(n7018) );
  INV_X1 U7939 ( .A(MORE_REG_SCAN_IN), .ZN(n7012) );
  OAI22_X1 U7940 ( .A1(n7012), .A2(keyinput_f44), .B1(n7011), .B2(
        keyinput_f110), .ZN(n7010) );
  AOI221_X1 U7941 ( .B1(n7012), .B2(keyinput_f44), .C1(keyinput_f110), .C2(
        n7011), .A(n7010), .ZN(n7017) );
  OAI22_X1 U7942 ( .A1(n7015), .A2(keyinput_f19), .B1(n7014), .B2(keyinput_f29), .ZN(n7013) );
  AOI221_X1 U7943 ( .B1(n7015), .B2(keyinput_f19), .C1(keyinput_f29), .C2(
        n7014), .A(n7013), .ZN(n7016) );
  NAND4_X1 U7944 ( .A1(n7019), .A2(n7018), .A3(n7017), .A4(n7016), .ZN(n7070)
         );
  OAI22_X1 U7945 ( .A1(keyinput_f115), .A2(n7022), .B1(n7021), .B2(
        keyinput_f85), .ZN(n7020) );
  AOI221_X1 U7946 ( .B1(n7022), .B2(keyinput_f115), .C1(n7021), .C2(
        keyinput_f85), .A(n7020), .ZN(n7035) );
  INV_X1 U7947 ( .A(keyinput_f105), .ZN(n7024) );
  OAI22_X1 U7948 ( .A1(keyinput_f104), .A2(n7025), .B1(n7024), .B2(
        DATAWIDTH_REG_1__SCAN_IN), .ZN(n7023) );
  AOI221_X1 U7949 ( .B1(n7025), .B2(keyinput_f104), .C1(n7024), .C2(
        DATAWIDTH_REG_1__SCAN_IN), .A(n7023), .ZN(n7034) );
  OAI22_X1 U7950 ( .A1(n7028), .A2(keyinput_f35), .B1(n7027), .B2(keyinput_f59), .ZN(n7026) );
  AOI221_X1 U7951 ( .B1(n7028), .B2(keyinput_f35), .C1(keyinput_f59), .C2(
        n7027), .A(n7026), .ZN(n7033) );
  INV_X1 U7952 ( .A(keyinput_f34), .ZN(n7030) );
  OAI22_X1 U7953 ( .A1(n7031), .A2(keyinput_f63), .B1(n7030), .B2(BS16_N), 
        .ZN(n7029) );
  AOI221_X1 U7954 ( .B1(n7031), .B2(keyinput_f63), .C1(BS16_N), .C2(n7030), 
        .A(n7029), .ZN(n7032) );
  NAND4_X1 U7955 ( .A1(n7035), .A2(n7034), .A3(n7033), .A4(n7032), .ZN(n7069)
         );
  INV_X1 U7956 ( .A(keyinput_f33), .ZN(n7037) );
  OAI22_X1 U7957 ( .A1(n7038), .A2(keyinput_f66), .B1(n7037), .B2(NA_N), .ZN(
        n7036) );
  AOI221_X1 U7958 ( .B1(n7038), .B2(keyinput_f66), .C1(NA_N), .C2(n7037), .A(
        n7036), .ZN(n7067) );
  XOR2_X1 U7959 ( .A(ADDRESS_REG_0__SCAN_IN), .B(keyinput_f100), .Z(n7048) );
  XOR2_X1 U7960 ( .A(keyinput_f127), .B(DATAWIDTH_REG_23__SCAN_IN), .Z(n7047)
         );
  AOI22_X1 U7961 ( .A1(n7041), .A2(keyinput_f93), .B1(n7040), .B2(
        keyinput_f101), .ZN(n7039) );
  OAI221_X1 U7962 ( .B1(n7041), .B2(keyinput_f93), .C1(n7040), .C2(
        keyinput_f101), .A(n7039), .ZN(n7046) );
  AOI22_X1 U7963 ( .A1(n7044), .A2(keyinput_f72), .B1(n7043), .B2(keyinput_f39), .ZN(n7042) );
  OAI221_X1 U7964 ( .B1(n7044), .B2(keyinput_f72), .C1(n7043), .C2(
        keyinput_f39), .A(n7042), .ZN(n7045) );
  NOR4_X1 U7965 ( .A1(n7048), .A2(n7047), .A3(n7046), .A4(n7045), .ZN(n7066)
         );
  OAI22_X1 U7966 ( .A1(keyinput_f123), .A2(n7051), .B1(n7050), .B2(
        keyinput_f90), .ZN(n7049) );
  AOI221_X1 U7967 ( .B1(n7051), .B2(keyinput_f123), .C1(n7050), .C2(
        keyinput_f90), .A(n7049), .ZN(n7065) );
  AOI22_X1 U7968 ( .A1(n7054), .A2(keyinput_f2), .B1(keyinput_f108), .B2(n7053), .ZN(n7052) );
  OAI221_X1 U7969 ( .B1(n7054), .B2(keyinput_f2), .C1(n7053), .C2(
        keyinput_f108), .A(n7052), .ZN(n7063) );
  AOI22_X1 U7970 ( .A1(n7057), .A2(keyinput_f54), .B1(n7056), .B2(keyinput_f43), .ZN(n7055) );
  OAI221_X1 U7971 ( .B1(n7057), .B2(keyinput_f54), .C1(n7056), .C2(
        keyinput_f43), .A(n7055), .ZN(n7062) );
  AOI22_X1 U7972 ( .A1(n7060), .A2(keyinput_f38), .B1(keyinput_f89), .B2(n7059), .ZN(n7058) );
  OAI221_X1 U7973 ( .B1(n7060), .B2(keyinput_f38), .C1(n7059), .C2(
        keyinput_f89), .A(n7058), .ZN(n7061) );
  NOR3_X1 U7974 ( .A1(n7063), .A2(n7062), .A3(n7061), .ZN(n7064) );
  NAND4_X1 U7975 ( .A1(n7067), .A2(n7066), .A3(n7065), .A4(n7064), .ZN(n7068)
         );
  NOR4_X1 U7976 ( .A1(n7071), .A2(n7070), .A3(n7069), .A4(n7068), .ZN(n7072)
         );
  NAND4_X1 U7977 ( .A1(n7075), .A2(n7074), .A3(n7073), .A4(n7072), .ZN(n7077)
         );
  AOI21_X1 U7978 ( .B1(keyinput_f45), .B2(n7077), .A(keyinput_g45), .ZN(n7079)
         );
  INV_X1 U7979 ( .A(keyinput_f45), .ZN(n7076) );
  AOI21_X1 U7980 ( .B1(n7077), .B2(n7076), .A(n7080), .ZN(n7078) );
  AOI22_X1 U7981 ( .A1(n7080), .A2(n7079), .B1(keyinput_g45), .B2(n7078), .ZN(
        n7081) );
  AOI21_X1 U7982 ( .B1(n7083), .B2(n7082), .A(n7081), .ZN(n7087) );
  AOI22_X1 U7983 ( .A1(n7085), .A2(BYTEENABLE_REG_3__SCAN_IN), .B1(
        BE_N_REG_3__SCAN_IN), .B2(n7084), .ZN(n7086) );
  XNOR2_X1 U7984 ( .A(n7087), .B(n7086), .ZN(U3445) );
  CLKBUF_X2 U3609 ( .A(n3293), .Z(n3966) );
  BUF_X1 U3674 ( .A(n3478), .Z(n4457) );
  CLKBUF_X1 U3619 ( .A(n3392), .Z(n3369) );
  CLKBUF_X1 U3620 ( .A(n3350), .Z(n3479) );
  CLKBUF_X1 U3724 ( .A(n4105), .Z(n4194) );
  CLKBUF_X1 U3910 ( .A(n3308), .Z(n4612) );
  CLKBUF_X1 U4006 ( .A(n3307), .Z(n3461) );
  CLKBUF_X1 U4026 ( .A(n5705), .Z(n6127) );
  CLKBUF_X1 U4263 ( .A(n6332), .Z(n6323) );
  CLKBUF_X1 U4487 ( .A(n3603), .Z(n3831) );
endmodule

