

module b20_C_AntiSAT_k_256_8 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, 
        keyinput128, keyinput129, keyinput130, keyinput131, keyinput132, 
        keyinput133, keyinput134, keyinput135, keyinput136, keyinput137, 
        keyinput138, keyinput139, keyinput140, keyinput141, keyinput142, 
        keyinput143, keyinput144, keyinput145, keyinput146, keyinput147, 
        keyinput148, keyinput149, keyinput150, keyinput151, keyinput152, 
        keyinput153, keyinput154, keyinput155, keyinput156, keyinput157, 
        keyinput158, keyinput159, keyinput160, keyinput161, keyinput162, 
        keyinput163, keyinput164, keyinput165, keyinput166, keyinput167, 
        keyinput168, keyinput169, keyinput170, keyinput171, keyinput172, 
        keyinput173, keyinput174, keyinput175, keyinput176, keyinput177, 
        keyinput178, keyinput179, keyinput180, keyinput181, keyinput182, 
        keyinput183, keyinput184, keyinput185, keyinput186, keyinput187, 
        keyinput188, keyinput189, keyinput190, keyinput191, keyinput192, 
        keyinput193, keyinput194, keyinput195, keyinput196, keyinput197, 
        keyinput198, keyinput199, keyinput200, keyinput201, keyinput202, 
        keyinput203, keyinput204, keyinput205, keyinput206, keyinput207, 
        keyinput208, keyinput209, keyinput210, keyinput211, keyinput212, 
        keyinput213, keyinput214, keyinput215, keyinput216, keyinput217, 
        keyinput218, keyinput219, keyinput220, keyinput221, keyinput222, 
        keyinput223, keyinput224, keyinput225, keyinput226, keyinput227, 
        keyinput228, keyinput229, keyinput230, keyinput231, keyinput232, 
        keyinput233, keyinput234, keyinput235, keyinput236, keyinput237, 
        keyinput238, keyinput239, keyinput240, keyinput241, keyinput242, 
        keyinput243, keyinput244, keyinput245, keyinput246, keyinput247, 
        keyinput248, keyinput249, keyinput250, keyinput251, keyinput252, 
        keyinput253, keyinput254, keyinput255, ADD_1068_U4, ADD_1068_U55, 
        ADD_1068_U56, ADD_1068_U57, ADD_1068_U58, ADD_1068_U59, ADD_1068_U60, 
        ADD_1068_U61, ADD_1068_U62, ADD_1068_U63, ADD_1068_U47, ADD_1068_U48, 
        ADD_1068_U49, ADD_1068_U50, ADD_1068_U51, ADD_1068_U52, ADD_1068_U53, 
        ADD_1068_U54, ADD_1068_U5, ADD_1068_U46, U126, U123, P1_U3355, 
        P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, 
        P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, 
        P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, 
        P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, 
        P1_U3326, P1_U3325, P1_U3324, P1_U3439, P1_U3440, P1_U3323, P1_U3322, 
        P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, 
        P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, 
        P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, 
        P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, 
        P1_U3453, P1_U3456, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, 
        P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, 
        P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3509, P1_U3510, 
        P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, P1_U3517, 
        P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, P1_U3524, 
        P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, P1_U3531, 
        P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, P1_U3538, 
        P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, P1_U3545, 
        P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, P1_U3552, 
        P1_U3553, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, P1_U3288, 
        P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, 
        P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, 
        P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, 
        P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, P1_U3261, 
        P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, 
        P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, 
        P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3554, P1_U3555, P1_U3556, 
        P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, P1_U3563, 
        P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, P1_U3570, 
        P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, P1_U3577, 
        P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, P1_U3584, 
        P1_U3585, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, P1_U3237, 
        P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, 
        P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, 
        P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, 
        P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U3973, P2_U3295, 
        P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, 
        P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, 
        P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, 
        P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, 
        P2_U3266, P2_U3265, P2_U3264, P2_U3376, P2_U3377, P2_U3263, P2_U3262, 
        P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, 
        P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, 
        P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3390, P2_U3393, P2_U3396, P2_U3399, P2_U3402, P2_U3405, P2_U3408, 
        P2_U3411, P2_U3414, P2_U3417, P2_U3420, P2_U3423, P2_U3426, P2_U3429, 
        P2_U3432, P2_U3435, P2_U3438, P2_U3441, P2_U3444, P2_U3446, P2_U3447, 
        P2_U3448, P2_U3449, P2_U3450, P2_U3451, P2_U3452, P2_U3453, P2_U3454, 
        P2_U3455, P2_U3456, P2_U3457, P2_U3458, P2_U3459, P2_U3460, P2_U3461, 
        P2_U3462, P2_U3463, P2_U3464, P2_U3465, P2_U3466, P2_U3467, P2_U3468, 
        P2_U3469, P2_U3470, P2_U3471, P2_U3472, P2_U3473, P2_U3474, P2_U3475, 
        P2_U3476, P2_U3477, P2_U3478, P2_U3479, P2_U3480, P2_U3481, P2_U3482, 
        P2_U3483, P2_U3484, P2_U3485, P2_U3486, P2_U3487, P2_U3488, P2_U3489, 
        P2_U3490, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, 
        P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, 
        P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, 
        P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, P2_U3207, 
        P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, 
        P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, 
        P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, 
        P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3491, P2_U3492, P2_U3493, 
        P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, 
        P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, 
        P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, 
        P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, 
        P2_U3522, P2_U3296, P2_U3181, P2_U3180, P2_U3179, P2_U3178, P2_U3177, 
        P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, P2_U3171, P2_U3170, 
        P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, P2_U3164, P2_U3163, 
        P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, P2_U3157, P2_U3156, 
        P2_U3155, P2_U3154, P2_U3153, P2_U3151, P2_U3150, P2_U3893 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127, keyinput128, keyinput129,
         keyinput130, keyinput131, keyinput132, keyinput133, keyinput134,
         keyinput135, keyinput136, keyinput137, keyinput138, keyinput139,
         keyinput140, keyinput141, keyinput142, keyinput143, keyinput144,
         keyinput145, keyinput146, keyinput147, keyinput148, keyinput149,
         keyinput150, keyinput151, keyinput152, keyinput153, keyinput154,
         keyinput155, keyinput156, keyinput157, keyinput158, keyinput159,
         keyinput160, keyinput161, keyinput162, keyinput163, keyinput164,
         keyinput165, keyinput166, keyinput167, keyinput168, keyinput169,
         keyinput170, keyinput171, keyinput172, keyinput173, keyinput174,
         keyinput175, keyinput176, keyinput177, keyinput178, keyinput179,
         keyinput180, keyinput181, keyinput182, keyinput183, keyinput184,
         keyinput185, keyinput186, keyinput187, keyinput188, keyinput189,
         keyinput190, keyinput191, keyinput192, keyinput193, keyinput194,
         keyinput195, keyinput196, keyinput197, keyinput198, keyinput199,
         keyinput200, keyinput201, keyinput202, keyinput203, keyinput204,
         keyinput205, keyinput206, keyinput207, keyinput208, keyinput209,
         keyinput210, keyinput211, keyinput212, keyinput213, keyinput214,
         keyinput215, keyinput216, keyinput217, keyinput218, keyinput219,
         keyinput220, keyinput221, keyinput222, keyinput223, keyinput224,
         keyinput225, keyinput226, keyinput227, keyinput228, keyinput229,
         keyinput230, keyinput231, keyinput232, keyinput233, keyinput234,
         keyinput235, keyinput236, keyinput237, keyinput238, keyinput239,
         keyinput240, keyinput241, keyinput242, keyinput243, keyinput244,
         keyinput245, keyinput246, keyinput247, keyinput248, keyinput249,
         keyinput250, keyinput251, keyinput252, keyinput253, keyinput254,
         keyinput255;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515,
         n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525,
         n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535,
         n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545,
         n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555,
         n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565,
         n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575,
         n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585,
         n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595,
         n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605,
         n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615,
         n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625,
         n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635,
         n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645,
         n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655,
         n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665,
         n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675,
         n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685,
         n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695,
         n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705,
         n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715,
         n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725,
         n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735,
         n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745,
         n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755,
         n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765,
         n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775,
         n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785,
         n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795,
         n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805,
         n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815,
         n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825,
         n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835,
         n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845,
         n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855,
         n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865,
         n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875,
         n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885,
         n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895,
         n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905,
         n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915,
         n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925,
         n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935,
         n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945,
         n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955,
         n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965,
         n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975,
         n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985,
         n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995,
         n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005,
         n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015,
         n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025,
         n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035,
         n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045,
         n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055,
         n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065,
         n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075,
         n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085,
         n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095,
         n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105,
         n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115,
         n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125,
         n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135,
         n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145,
         n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155,
         n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165,
         n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175,
         n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185,
         n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195,
         n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205,
         n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215,
         n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225,
         n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235,
         n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245,
         n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255,
         n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265,
         n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275,
         n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285,
         n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295,
         n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305,
         n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315,
         n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325,
         n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335,
         n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345,
         n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355,
         n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365,
         n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375,
         n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385,
         n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395,
         n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405,
         n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415,
         n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425,
         n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435,
         n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445,
         n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455,
         n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465,
         n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475,
         n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485,
         n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495,
         n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505,
         n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515,
         n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525,
         n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535,
         n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545,
         n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555,
         n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565,
         n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575,
         n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585,
         n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595,
         n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605,
         n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615,
         n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625,
         n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635,
         n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645,
         n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655,
         n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665,
         n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675,
         n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685,
         n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695,
         n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705,
         n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715,
         n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725,
         n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735,
         n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745,
         n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755,
         n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765,
         n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775,
         n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785,
         n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795,
         n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805,
         n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815,
         n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825,
         n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835,
         n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845,
         n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855,
         n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865,
         n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875,
         n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885,
         n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895,
         n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905,
         n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915,
         n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925,
         n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935,
         n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945,
         n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955,
         n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965,
         n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975,
         n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985,
         n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995,
         n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005,
         n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015,
         n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025,
         n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035,
         n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045,
         n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055,
         n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065,
         n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075,
         n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085,
         n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095,
         n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105,
         n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115,
         n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125,
         n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135,
         n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145,
         n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155,
         n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165,
         n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175,
         n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185,
         n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195,
         n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205,
         n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215,
         n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225,
         n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235,
         n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245,
         n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255,
         n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265,
         n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275,
         n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285,
         n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295,
         n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305,
         n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315,
         n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325,
         n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335,
         n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345,
         n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355,
         n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365,
         n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375,
         n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385,
         n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395,
         n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405,
         n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415,
         n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425,
         n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435,
         n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445,
         n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455,
         n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465,
         n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475,
         n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485,
         n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495,
         n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505,
         n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515,
         n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525,
         n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535,
         n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545,
         n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555,
         n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565,
         n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575,
         n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585,
         n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595,
         n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605,
         n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615,
         n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625,
         n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635,
         n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645,
         n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655,
         n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665,
         n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675,
         n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685,
         n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695,
         n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705,
         n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715,
         n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725,
         n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735,
         n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745,
         n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755,
         n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765,
         n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775,
         n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785,
         n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795,
         n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805,
         n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815,
         n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825,
         n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835,
         n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845,
         n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855,
         n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865,
         n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875,
         n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885,
         n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895,
         n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905,
         n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915,
         n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925,
         n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935,
         n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945,
         n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955,
         n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965,
         n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975,
         n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985,
         n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995,
         n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005,
         n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015,
         n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025,
         n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035,
         n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045,
         n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055,
         n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065,
         n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075,
         n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085,
         n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095,
         n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105,
         n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115,
         n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125,
         n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135,
         n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145,
         n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155,
         n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165,
         n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175,
         n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185,
         n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195,
         n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205,
         n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215,
         n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225,
         n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235,
         n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245,
         n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255,
         n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265,
         n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275,
         n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285,
         n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295,
         n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305,
         n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315,
         n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325,
         n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335,
         n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345,
         n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355,
         n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365,
         n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375,
         n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385,
         n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395,
         n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405,
         n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415,
         n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425,
         n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435,
         n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445,
         n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455,
         n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465,
         n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475,
         n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485,
         n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495,
         n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505,
         n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515,
         n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525,
         n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535,
         n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545,
         n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555,
         n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565,
         n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575,
         n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585,
         n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595,
         n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605,
         n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615,
         n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625,
         n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635,
         n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645,
         n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655,
         n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665,
         n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675,
         n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685,
         n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695,
         n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705,
         n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715,
         n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725,
         n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735,
         n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745,
         n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755,
         n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765,
         n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775,
         n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785,
         n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795,
         n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805,
         n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815,
         n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825,
         n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835,
         n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845,
         n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855,
         n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865,
         n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875,
         n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885,
         n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895,
         n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905,
         n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915,
         n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925,
         n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935,
         n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945,
         n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955,
         n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965,
         n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975,
         n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985,
         n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995,
         n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005,
         n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015,
         n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025,
         n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035,
         n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045,
         n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055,
         n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065,
         n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075,
         n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085,
         n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095,
         n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105,
         n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115,
         n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125,
         n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135,
         n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145,
         n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155,
         n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165,
         n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175,
         n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185,
         n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195,
         n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205,
         n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215,
         n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225,
         n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235,
         n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245,
         n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255,
         n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265,
         n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275,
         n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285,
         n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295,
         n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305,
         n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315,
         n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325,
         n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335,
         n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345,
         n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355,
         n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365,
         n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375,
         n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385,
         n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395,
         n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405,
         n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415,
         n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425,
         n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435,
         n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445,
         n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455,
         n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465,
         n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475,
         n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485,
         n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495,
         n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505,
         n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515,
         n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525,
         n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535,
         n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545,
         n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555,
         n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565,
         n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575,
         n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585,
         n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595,
         n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605,
         n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615,
         n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625,
         n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635,
         n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645,
         n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655,
         n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665,
         n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675,
         n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685,
         n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695,
         n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705,
         n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715,
         n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725,
         n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735,
         n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745,
         n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755,
         n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765,
         n8766, n8767, n8768, n8769, n8770, n8771, n8773, n8774, n8775, n8776,
         n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786,
         n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796,
         n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806,
         n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816,
         n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826,
         n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836,
         n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846,
         n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856,
         n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866,
         n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876,
         n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886,
         n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896,
         n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906,
         n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916,
         n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926,
         n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936,
         n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946,
         n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956,
         n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966,
         n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976,
         n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986,
         n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996,
         n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006,
         n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016,
         n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026,
         n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036,
         n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046,
         n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056,
         n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066,
         n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076,
         n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086,
         n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096,
         n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106,
         n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116,
         n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126,
         n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136,
         n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146,
         n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156,
         n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166,
         n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176,
         n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186,
         n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196,
         n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206,
         n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216,
         n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226,
         n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236,
         n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246,
         n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256,
         n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266,
         n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276,
         n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286,
         n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296,
         n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306,
         n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316,
         n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326,
         n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336,
         n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346,
         n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356,
         n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366,
         n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376,
         n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386,
         n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396,
         n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406,
         n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416,
         n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426,
         n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436,
         n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446,
         n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456,
         n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466,
         n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476,
         n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486,
         n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496,
         n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506,
         n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516,
         n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526,
         n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536,
         n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546,
         n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556,
         n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566,
         n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576,
         n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586,
         n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596,
         n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606,
         n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616,
         n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626,
         n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636,
         n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646,
         n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656,
         n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666,
         n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676,
         n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686,
         n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696,
         n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706,
         n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716,
         n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726,
         n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736,
         n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746,
         n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756,
         n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766,
         n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776,
         n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786,
         n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796,
         n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806,
         n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816,
         n9817, n9818, n9819, n9820, n9821, n9822, n9824, n9825, n9826, n9827,
         n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837,
         n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847,
         n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857,
         n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867,
         n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877,
         n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887,
         n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897,
         n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907,
         n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917,
         n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927,
         n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938,
         n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948,
         n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958,
         n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968,
         n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978,
         n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988,
         n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998,
         n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
         n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
         n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
         n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
         n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
         n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
         n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247,
         n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255,
         n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263,
         n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271,
         n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279,
         n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287,
         n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295,
         n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303,
         n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311,
         n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319,
         n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327,
         n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335,
         n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343,
         n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351,
         n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359,
         n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367,
         n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375,
         n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383,
         n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391,
         n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399,
         n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407,
         n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415,
         n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423,
         n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431,
         n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439,
         n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447,
         n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455,
         n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463,
         n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471,
         n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479,
         n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487,
         n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495,
         n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503,
         n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511,
         n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519,
         n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527,
         n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535,
         n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543,
         n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551,
         n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559,
         n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567,
         n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575,
         n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583,
         n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591,
         n10592, n10593, n10594, n10595, n10596, n10597, n10598;

  INV_X4 U5012 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  NAND2_X1 U5013 ( .A1(n6891), .A2(n6892), .ZN(n8189) );
  AND2_X1 U5014 ( .A1(n5317), .A2(n5316), .ZN(n9898) );
  NAND4_X1 U5015 ( .A1(n5248), .A2(n5247), .A3(n5246), .A4(n5245), .ZN(n9263)
         );
  NAND2_X1 U5016 ( .A1(n5346), .A2(n5345), .ZN(n5353) );
  BUF_X1 U5017 ( .A(n6052), .Z(n4514) );
  INV_X2 U5018 ( .A(n6709), .ZN(n5718) );
  CLKBUF_X3 U5019 ( .A(n6255), .Z(n4517) );
  AND2_X1 U5020 ( .A1(n8773), .A2(n8161), .ZN(n6216) );
  NAND2_X1 U5021 ( .A1(n8773), .A2(n6190), .ZN(n6255) );
  BUF_X4 U5022 ( .A(n7328), .Z(n4507) );
  NAND2_X1 U5023 ( .A1(n6581), .A2(n6582), .ZN(n6587) );
  AND2_X1 U5024 ( .A1(n4821), .A2(n5836), .ZN(n4820) );
  XNOR2_X1 U5025 ( .A(n6156), .B(n6155), .ZN(n6581) );
  INV_X1 U5026 ( .A(n9096), .ZN(n8983) );
  AOI21_X1 U5027 ( .B1(n9345), .B2(n9908), .A(n5796), .ZN(n6640) );
  OR2_X1 U5028 ( .A1(n8592), .A2(n5099), .ZN(n5096) );
  INV_X1 U5029 ( .A(n8087), .ZN(n8090) );
  NAND2_X1 U5030 ( .A1(n5096), .A2(n5094), .ZN(n8567) );
  INV_X1 U5031 ( .A(n8075), .ZN(n6460) );
  AND2_X1 U5032 ( .A1(n9150), .A2(n9223), .ZN(n5835) );
  INV_X1 U5033 ( .A(n8962), .ZN(n5559) );
  INV_X1 U5034 ( .A(n8189), .ZN(n8196) );
  INV_X1 U5035 ( .A(n4517), .ZN(n6532) );
  OR2_X1 U5036 ( .A1(n7776), .A2(n4808), .ZN(n4806) );
  OAI21_X1 U5037 ( .B1(n7879), .B2(n6409), .A(n6408), .ZN(n7895) );
  OR2_X1 U5038 ( .A1(n7900), .A2(n8015), .ZN(n6571) );
  INV_X1 U5039 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n6246) );
  BUF_X1 U5040 ( .A(n6234), .Z(n6308) );
  INV_X1 U5042 ( .A(n9107), .ZN(n7059) );
  NAND2_X1 U5043 ( .A1(n9170), .A2(n9010), .ZN(n9115) );
  AND2_X1 U5044 ( .A1(n5297), .A2(n5296), .ZN(n7353) );
  INV_X1 U5045 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n6161) );
  OR2_X1 U5046 ( .A1(n4618), .A2(n6890), .ZN(n4617) );
  AND4_X1 U5047 ( .A1(n6244), .A2(n6243), .A3(n6242), .A4(n6241), .ZN(n7953)
         );
  NAND2_X1 U5048 ( .A1(n8590), .A2(n8034), .ZN(n8575) );
  NAND2_X1 U5049 ( .A1(n5026), .A2(n6337), .ZN(n10139) );
  XNOR2_X1 U5050 ( .A(n6185), .B(n8764), .ZN(n6191) );
  NAND2_X1 U5051 ( .A1(n8917), .A2(n8921), .ZN(n8836) );
  NOR2_X1 U5052 ( .A1(P2_ADDR_REG_19__SCAN_IN), .A2(P1_ADDR_REG_19__SCAN_IN), 
        .ZN(n7269) );
  NAND2_X2 U5053 ( .A1(n6233), .A2(n5135), .ZN(n8318) );
  BUF_X1 U5054 ( .A(n6191), .Z(n8773) );
  XNOR2_X1 U5055 ( .A(n6262), .B(n6261), .ZN(n7780) );
  NAND2_X1 U5056 ( .A1(n6189), .A2(n8161), .ZN(n7328) );
  INV_X2 U5057 ( .A(n9561), .ZN(n9857) );
  NAND2_X2 U5058 ( .A1(n8567), .A2(n6477), .ZN(n8552) );
  NAND2_X2 U5059 ( .A1(n6953), .A2(n6954), .ZN(n7025) );
  AND2_X2 U5060 ( .A1(n5843), .A2(n7026), .ZN(n6953) );
  NAND2_X2 U5061 ( .A1(n5353), .A2(n5352), .ZN(n5370) );
  NAND3_X2 U5062 ( .A1(n5912), .A2(n4854), .A3(n5911), .ZN(n7598) );
  INV_X1 U5063 ( .A(n4517), .ZN(n4506) );
  NOR2_X2 U5064 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n4834) );
  NAND2_X2 U5065 ( .A1(n7650), .A2(n5920), .ZN(n5927) );
  OAI21_X2 U5066 ( .B1(n9156), .B2(n9108), .A(n9155), .ZN(n7152) );
  NAND2_X2 U5067 ( .A1(n8973), .A2(n9152), .ZN(n9156) );
  NAND2_X2 U5068 ( .A1(n5879), .A2(n5881), .ZN(n7140) );
  NOR2_X2 U5069 ( .A1(n8398), .A2(n4628), .ZN(n8417) );
  INV_X1 U5070 ( .A(n7936), .ZN(n5431) );
  INV_X4 U5071 ( .A(n7936), .ZN(n5011) );
  XNOR2_X2 U5072 ( .A(n5961), .B(n5962), .ZN(n8790) );
  NAND2_X2 U5073 ( .A1(n4835), .A2(n4836), .ZN(n5961) );
  OAI21_X2 U5074 ( .B1(n8604), .B2(n6572), .A(n8032), .ZN(n8588) );
  NAND2_X2 U5075 ( .A1(n5557), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5558) );
  AND3_X1 U5076 ( .A1(n8943), .A2(n4518), .A3(n4610), .ZN(n6131) );
  NAND2_X1 U5077 ( .A1(n4850), .A2(n4851), .ZN(n8943) );
  NAND2_X1 U5078 ( .A1(n4738), .A2(n4536), .ZN(n9350) );
  AOI21_X1 U5079 ( .B1(n6118), .B2(n9549), .A(n6117), .ZN(n9365) );
  AOI21_X1 U5080 ( .B1(n8482), .B2(n8623), .A(n8481), .ZN(n8638) );
  NAND2_X1 U5081 ( .A1(n9398), .A2(n9145), .ZN(n9383) );
  OAI22_X1 U5082 ( .A1(n8508), .A2(n8514), .B1(n8521), .B2(n8714), .ZN(n8500)
         );
  CLKBUF_X1 U5083 ( .A(n8855), .Z(n4511) );
  AND2_X1 U5084 ( .A1(n5116), .A2(n4527), .ZN(n5115) );
  NAND2_X1 U5085 ( .A1(n8963), .A2(n8962), .ZN(n9665) );
  NAND2_X1 U5086 ( .A1(n8790), .A2(n8792), .ZN(n8791) );
  NAND2_X1 U5087 ( .A1(n8093), .A2(n8084), .ZN(n8105) );
  OAI21_X1 U5088 ( .B1(n8575), .B2(n6573), .A(n8036), .ZN(n8565) );
  XNOR2_X1 U5089 ( .A(n7931), .B(SI_29_), .ZN(n8159) );
  XNOR2_X1 U5090 ( .A(n7929), .B(n7928), .ZN(n7931) );
  AOI21_X1 U5091 ( .B1(n7895), .B2(n7896), .A(n7898), .ZN(n8617) );
  NAND2_X1 U5092 ( .A1(n6509), .A2(n6508), .ZN(n8714) );
  NAND2_X1 U5093 ( .A1(n5475), .A2(n5474), .ZN(n9025) );
  NAND2_X1 U5094 ( .A1(n5471), .A2(n5470), .ZN(n5490) );
  CLKBUF_X1 U5095 ( .A(n8926), .Z(n4622) );
  NAND2_X1 U5096 ( .A1(n5360), .A2(n5359), .ZN(n7660) );
  NAND2_X1 U5097 ( .A1(n4830), .A2(n5899), .ZN(n4829) );
  NAND2_X1 U5098 ( .A1(n5414), .A2(n5413), .ZN(n8842) );
  NAND2_X1 U5099 ( .A1(n6355), .A2(n6354), .ZN(n10146) );
  NAND2_X1 U5100 ( .A1(n5378), .A2(n5377), .ZN(n7538) );
  NAND2_X1 U5101 ( .A1(n5354), .A2(n5370), .ZN(n6696) );
  AND2_X1 U5102 ( .A1(n5898), .A2(n5897), .ZN(n7336) );
  NAND2_X2 U5103 ( .A1(n7104), .A2(n9869), .ZN(n9561) );
  INV_X1 U5104 ( .A(n7409), .ZN(n7219) );
  INV_X1 U5105 ( .A(n7125), .ZN(n7307) );
  NAND2_X1 U5106 ( .A1(n9564), .A2(n9659), .ZN(n9908) );
  AND2_X1 U5107 ( .A1(n6293), .A2(n6292), .ZN(n10120) );
  AND3_X1 U5108 ( .A1(n5283), .A2(n5282), .A3(n5281), .ZN(n7409) );
  CLKBUF_X3 U5109 ( .A(n5850), .Z(n6066) );
  CLKBUF_X1 U5110 ( .A(n5908), .Z(n6072) );
  INV_X1 U5111 ( .A(n5908), .ZN(n4508) );
  AND4_X1 U5112 ( .A1(n6221), .A2(n6220), .A3(n6219), .A4(n6218), .ZN(n6689)
         );
  NAND2_X1 U5113 ( .A1(n6169), .A2(n10410), .ZN(n6392) );
  AND3_X1 U5114 ( .A1(n5237), .A2(n5236), .A3(n5235), .ZN(n9893) );
  CLKBUF_X1 U5115 ( .A(n5833), .Z(n4621) );
  BUF_X2 U5116 ( .A(n6216), .Z(n6491) );
  INV_X1 U5117 ( .A(n6216), .ZN(n6543) );
  NAND2_X1 U5118 ( .A1(n5259), .A2(n5258), .ZN(n5271) );
  INV_X1 U5119 ( .A(n9888), .ZN(n7112) );
  NAND4_X1 U5120 ( .A1(n5194), .A2(n5193), .A3(n5192), .A4(n5191), .ZN(n7074)
         );
  NAND2_X1 U5121 ( .A1(n5835), .A2(n5833), .ZN(n7631) );
  INV_X1 U5122 ( .A(n6380), .ZN(n6169) );
  NAND2_X1 U5123 ( .A1(n5835), .A2(n6657), .ZN(n5844) );
  CLKBUF_X1 U5124 ( .A(n5687), .Z(n5595) );
  OR2_X1 U5125 ( .A1(n5687), .A2(n6961), .ZN(n5171) );
  AND3_X1 U5126 ( .A1(n5220), .A2(n5219), .A3(n5218), .ZN(n9888) );
  INV_X1 U5127 ( .A(n6225), .ZN(n4509) );
  INV_X2 U5128 ( .A(n5206), .ZN(n5295) );
  NOR2_X1 U5129 ( .A1(n9734), .A2(n9739), .ZN(n5810) );
  NAND2_X1 U5130 ( .A1(n8962), .A2(n5011), .ZN(n5206) );
  NAND2_X1 U5131 ( .A1(n8767), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6185) );
  INV_X1 U5132 ( .A(n9726), .ZN(n5169) );
  NAND2_X1 U5133 ( .A1(n9720), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5166) );
  NAND2_X1 U5134 ( .A1(n5532), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5556) );
  INV_X1 U5135 ( .A(n5806), .ZN(n9734) );
  INV_X1 U5136 ( .A(n6779), .ZN(n4799) );
  XNOR2_X1 U5137 ( .A(n5177), .B(n5176), .ZN(n5757) );
  XNOR2_X1 U5138 ( .A(n5179), .B(n5178), .ZN(n8163) );
  OR2_X1 U5139 ( .A1(n5164), .A2(n5276), .ZN(n5162) );
  NAND2_X1 U5140 ( .A1(n4753), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5179) );
  NAND2_X2 U5141 ( .A1(n6235), .A2(n4815), .ZN(n6760) );
  OAI21_X1 U5142 ( .B1(n7936), .B2(n6667), .A(n5002), .ZN(n5209) );
  NAND2_X1 U5143 ( .A1(n6215), .A2(n6214), .ZN(n9935) );
  AND2_X1 U5144 ( .A1(n4552), .A2(n5178), .ZN(n4794) );
  AND2_X2 U5145 ( .A1(n5215), .A2(n5148), .ZN(n5275) );
  NOR2_X1 U5146 ( .A1(n5153), .A2(n5152), .ZN(n5154) );
  AND3_X1 U5147 ( .A1(n6142), .A2(n6141), .A3(n6351), .ZN(n6143) );
  AND2_X1 U5148 ( .A1(n5155), .A2(n4915), .ZN(n4914) );
  AND2_X1 U5149 ( .A1(n6212), .A2(n4818), .ZN(n6234) );
  BUF_X1 U5150 ( .A(n6212), .Z(n6213) );
  NAND2_X1 U5151 ( .A1(n7268), .A2(n4951), .ZN(n5182) );
  AND2_X1 U5152 ( .A1(P2_ADDR_REG_19__SCAN_IN), .A2(P1_ADDR_REG_19__SCAN_IN), 
        .ZN(n7268) );
  INV_X1 U5153 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n5372) );
  INV_X1 U5154 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n5279) );
  INV_X4 U5155 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X1 U5156 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5149) );
  NOR2_X1 U5157 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n5150) );
  INV_X1 U5158 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n6447) );
  INV_X1 U5159 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n6351) );
  INV_X1 U5160 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n6248) );
  NOR2_X1 U5161 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_5__SCAN_IN), .ZN(
        n5048) );
  NOR2_X1 U5162 ( .A1(P2_IR_REG_4__SCAN_IN), .A2(P2_IR_REG_6__SCAN_IN), .ZN(
        n5047) );
  NOR2_X1 U5163 ( .A1(P2_IR_REG_14__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), .ZN(
        n6145) );
  INV_X1 U5164 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n6617) );
  INV_X1 U5165 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n6550) );
  INV_X1 U5166 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n6597) );
  NAND2_X1 U5167 ( .A1(n7048), .A2(n5872), .ZN(n4510) );
  AND2_X1 U5168 ( .A1(n8918), .A2(n8919), .ZN(n4512) );
  NAND2_X2 U5169 ( .A1(n8808), .A2(n8809), .ZN(n7048) );
  NAND2_X1 U5170 ( .A1(n8791), .A2(n5964), .ZN(n8855) );
  AND2_X1 U5171 ( .A1(n5858), .A2(n5860), .ZN(n7027) );
  OR2_X1 U5172 ( .A1(n5857), .A2(n5856), .ZN(n5858) );
  NAND2_X2 U5173 ( .A1(n7946), .A2(n7949), .ZN(n6561) );
  INV_X1 U5174 ( .A(n5844), .ZN(n4513) );
  INV_X1 U5175 ( .A(n5844), .ZN(n6071) );
  AND2_X2 U5176 ( .A1(n4853), .A2(n4852), .ZN(n8941) );
  NAND2_X1 U5177 ( .A1(n7030), .A2(n5860), .ZN(n8808) );
  NOR2_X2 U5178 ( .A1(n6150), .A2(n6149), .ZN(n6151) );
  AND2_X2 U5179 ( .A1(n4834), .A2(n4833), .ZN(n5215) );
  OAI21_X2 U5180 ( .B1(n7121), .B2(n6285), .A(n6284), .ZN(n7290) );
  NAND2_X2 U5181 ( .A1(n4516), .A2(n5850), .ZN(n5861) );
  INV_X2 U5182 ( .A(n5908), .ZN(n6068) );
  BUF_X4 U5183 ( .A(n6052), .Z(n4515) );
  INV_X1 U5184 ( .A(n5844), .ZN(n6052) );
  NAND3_X1 U5185 ( .A1(n6657), .A2(n5834), .A3(n7631), .ZN(n4516) );
  NAND2_X2 U5186 ( .A1(n5992), .A2(n8866), .ZN(n8816) );
  OR2_X2 U5187 ( .A1(n8880), .A2(n6048), .ZN(n4853) );
  AOI21_X2 U5188 ( .B1(n8799), .B2(n8878), .A(n8877), .ZN(n8880) );
  OAI21_X2 U5189 ( .B1(n8909), .B2(n8904), .A(n8800), .ZN(n8799) );
  NAND2_X1 U5190 ( .A1(n5038), .A2(n5035), .ZN(n4722) );
  NOR2_X1 U5191 ( .A1(n5037), .A2(n5036), .ZN(n5035) );
  AND2_X1 U5192 ( .A1(n8576), .A2(n4550), .ZN(n5100) );
  INV_X1 U5193 ( .A(n5391), .ZN(n4998) );
  XNOR2_X1 U5194 ( .A(n8547), .B(n8533), .ZN(n8548) );
  NAND2_X1 U5195 ( .A1(n5110), .A2(n5109), .ZN(n6507) );
  OR2_X1 U5196 ( .A1(n4527), .A2(n5114), .ZN(n5109) );
  OAI21_X1 U5197 ( .B1(n5038), .B2(n4578), .A(n5031), .ZN(n5030) );
  NAND2_X1 U5198 ( .A1(n5034), .A2(n5033), .ZN(n5032) );
  AOI21_X1 U5199 ( .B1(n4707), .B2(n8042), .A(n4706), .ZN(n4705) );
  NOR2_X1 U5200 ( .A1(n8657), .A2(n8533), .ZN(n4706) );
  INV_X1 U5201 ( .A(n8049), .ZN(n4707) );
  OAI21_X1 U5202 ( .B1(n4732), .B2(n4583), .A(n4731), .ZN(n8080) );
  NOR2_X1 U5203 ( .A1(n8105), .A2(n8069), .ZN(n4731) );
  OR2_X1 U5204 ( .A1(n6349), .A2(n5093), .ZN(n5092) );
  INV_X1 U5205 ( .A(n6335), .ZN(n5093) );
  INV_X1 U5206 ( .A(n8828), .ZN(n4842) );
  INV_X1 U5207 ( .A(n4979), .ZN(n4978) );
  AND2_X1 U5208 ( .A1(n4985), .A2(n4983), .ZN(n4982) );
  INV_X1 U5209 ( .A(n5528), .ZN(n4983) );
  NAND2_X1 U5210 ( .A1(n5326), .A2(n5325), .ZN(n5345) );
  NAND2_X1 U5211 ( .A1(n8270), .A2(n8180), .ZN(n8184) );
  NOR2_X1 U5212 ( .A1(n5067), .A2(n5068), .ZN(n5066) );
  INV_X1 U5213 ( .A(n6892), .ZN(n5051) );
  OAI21_X1 U5214 ( .B1(n6674), .B2(P2_D_REG_0__SCAN_IN), .A(n6692), .ZN(n6886)
         );
  INV_X1 U5215 ( .A(n6191), .ZN(n6189) );
  NAND2_X1 U5216 ( .A1(n6762), .A2(n6761), .ZN(n6763) );
  NAND2_X1 U5217 ( .A1(n4798), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n4797) );
  NAND2_X1 U5218 ( .A1(n9966), .A2(n7766), .ZN(n4814) );
  NAND2_X1 U5219 ( .A1(n9976), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n7766) );
  NAND2_X1 U5220 ( .A1(n4589), .A2(n5131), .ZN(n5126) );
  AND2_X1 U5221 ( .A1(n8702), .A2(n8502), .ZN(n5132) );
  INV_X1 U5222 ( .A(n5133), .ZN(n5129) );
  OR2_X1 U5223 ( .A1(n8175), .A2(n8306), .ZN(n8048) );
  OR2_X1 U5224 ( .A1(n8714), .A2(n8298), .ZN(n8060) );
  NAND2_X1 U5225 ( .A1(n8714), .A2(n8298), .ZN(n8059) );
  NAND2_X1 U5226 ( .A1(n6593), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6618) );
  NOR2_X1 U5227 ( .A1(n4547), .A2(n4525), .ZN(n4848) );
  NOR2_X1 U5228 ( .A1(n9373), .A2(n6119), .ZN(n5792) );
  OR2_X1 U5229 ( .A1(n6119), .A2(n7024), .ZN(n9080) );
  OR2_X1 U5230 ( .A1(n9375), .A2(n8947), .ZN(n9081) );
  OR2_X1 U5231 ( .A1(n9392), .A2(n6056), .ZN(n9078) );
  NAND2_X1 U5232 ( .A1(n9392), .A2(n6056), .ZN(n9195) );
  OR2_X1 U5233 ( .A1(n9404), .A2(n8945), .ZN(n9145) );
  OR2_X1 U5234 ( .A1(n8842), .A2(n7700), .ZN(n9014) );
  NAND2_X1 U5235 ( .A1(n8072), .A2(n8071), .ZN(n8074) );
  NAND2_X1 U5236 ( .A1(n4913), .A2(n4849), .ZN(n5743) );
  AND2_X1 U5237 ( .A1(n4914), .A2(n5513), .ZN(n4849) );
  AOI21_X1 U5238 ( .B1(n4996), .B2(n4528), .A(n4585), .ZN(n4995) );
  NAND2_X1 U5239 ( .A1(n5408), .A2(n5398), .ZN(n5409) );
  AND2_X1 U5240 ( .A1(n5369), .A2(n5351), .ZN(n5352) );
  INV_X1 U5241 ( .A(n5309), .ZN(n5310) );
  NAND2_X1 U5242 ( .A1(n5060), .A2(n5059), .ZN(n5058) );
  OR2_X1 U5243 ( .A1(n8197), .A2(n5061), .ZN(n5060) );
  NAND2_X1 U5244 ( .A1(n8197), .A2(n5062), .ZN(n5059) );
  AND2_X1 U5245 ( .A1(n5062), .A2(n8203), .ZN(n5061) );
  INV_X1 U5246 ( .A(n7622), .ZN(n5077) );
  INV_X1 U5247 ( .A(n7717), .ZN(n5078) );
  INV_X1 U5248 ( .A(n8184), .ZN(n8182) );
  OR2_X1 U5249 ( .A1(n8250), .A2(n4680), .ZN(n4676) );
  AND2_X1 U5250 ( .A1(n4681), .A2(n4685), .ZN(n4679) );
  NAND2_X1 U5251 ( .A1(n4952), .A2(n4954), .ZN(n4618) );
  AOI21_X1 U5252 ( .B1(n4955), .B2(n8090), .A(n8104), .ZN(n4954) );
  OAI21_X1 U5253 ( .B1(n4953), .B2(n5013), .A(n5012), .ZN(n4952) );
  NAND2_X1 U5254 ( .A1(n8088), .A2(n8136), .ZN(n5012) );
  AND2_X1 U5255 ( .A1(n8691), .A2(n8082), .ZN(n8146) );
  INV_X1 U5256 ( .A(n6229), .ZN(n6540) );
  INV_X1 U5257 ( .A(n6152), .ZN(n6376) );
  OR2_X1 U5258 ( .A1(n6376), .A2(P2_IR_REG_11__SCAN_IN), .ZN(n6388) );
  XNOR2_X1 U5259 ( .A(n8635), .B(n8494), .ZN(n8484) );
  NAND2_X1 U5260 ( .A1(n6183), .A2(n6182), .ZN(n6530) );
  INV_X1 U5261 ( .A(n6521), .ZN(n6183) );
  OR2_X1 U5262 ( .A1(n8736), .A2(n8580), .ZN(n6477) );
  AND2_X1 U5263 ( .A1(n7965), .A2(n7286), .ZN(n7975) );
  NAND2_X1 U5264 ( .A1(n6587), .A2(n7936), .ZN(n6263) );
  AOI21_X1 U5265 ( .B1(n5118), .B2(n4519), .A(n4581), .ZN(n5117) );
  NAND2_X1 U5266 ( .A1(n8552), .A2(n5118), .ZN(n5116) );
  AOI21_X1 U5267 ( .B1(n5100), .B2(n5098), .A(n5141), .ZN(n5097) );
  INV_X1 U5268 ( .A(n6457), .ZN(n5098) );
  NOR2_X1 U5269 ( .A1(n8008), .A2(n5105), .ZN(n5104) );
  INV_X1 U5270 ( .A(n6386), .ZN(n5105) );
  AND2_X1 U5271 ( .A1(n9665), .A2(n9335), .ZN(n9209) );
  AND4_X1 U5272 ( .A1(n5407), .A2(n5406), .A3(n5405), .A4(n5404), .ZN(n7606)
         );
  NAND2_X1 U5273 ( .A1(n5792), .A2(n6635), .ZN(n9339) );
  NOR2_X1 U5274 ( .A1(n5584), .A2(n4792), .ZN(n4791) );
  INV_X1 U5275 ( .A(n5572), .ZN(n4792) );
  AND2_X1 U5276 ( .A1(n4744), .A2(n4742), .ZN(n4619) );
  INV_X1 U5277 ( .A(n7872), .ZN(n9578) );
  NAND2_X1 U5278 ( .A1(n5574), .A2(n5573), .ZN(n5587) );
  NAND2_X1 U5279 ( .A1(n7269), .A2(n5180), .ZN(n5181) );
  INV_X1 U5280 ( .A(P1_RD_REG_SCAN_IN), .ZN(n5180) );
  INV_X1 U5281 ( .A(n6587), .ZN(n6655) );
  OAI21_X1 U5282 ( .B1(n5694), .B2(n4779), .A(n4777), .ZN(n5738) );
  AOI21_X1 U5283 ( .B1(n4778), .B2(n4780), .A(n4600), .ZN(n4777) );
  INV_X1 U5284 ( .A(n4780), .ZN(n4779) );
  NAND2_X1 U5285 ( .A1(n4908), .A2(n8985), .ZN(n8991) );
  AND2_X1 U5286 ( .A1(n4904), .A2(n4903), .ZN(n8989) );
  AOI21_X1 U5287 ( .B1(n4567), .B2(n5146), .A(n4909), .ZN(n4903) );
  NOR2_X1 U5288 ( .A1(n5022), .A2(n5023), .ZN(n5018) );
  AND2_X1 U5289 ( .A1(n5019), .A2(n5016), .ZN(n5015) );
  NAND2_X1 U5290 ( .A1(n8011), .A2(n5020), .ZN(n5019) );
  AND2_X1 U5291 ( .A1(n8014), .A2(n8128), .ZN(n5016) );
  NOR2_X1 U5292 ( .A1(n5023), .A2(n5021), .ZN(n5020) );
  NAND2_X1 U5293 ( .A1(n4723), .A2(n5039), .ZN(n5038) );
  NAND2_X1 U5294 ( .A1(n8030), .A2(n8090), .ZN(n5039) );
  INV_X1 U5295 ( .A(n8043), .ZN(n4709) );
  AOI21_X1 U5296 ( .B1(n4710), .B2(n8090), .A(n4886), .ZN(n4703) );
  NAND2_X1 U5297 ( .A1(n8052), .A2(n8047), .ZN(n4710) );
  AOI21_X1 U5298 ( .B1(n9039), .B2(n4910), .A(n9533), .ZN(n9045) );
  INV_X1 U5299 ( .A(n9062), .ZN(n4928) );
  NAND2_X1 U5300 ( .A1(n5029), .A2(n8055), .ZN(n5028) );
  NAND2_X1 U5301 ( .A1(n8061), .A2(n8501), .ZN(n4733) );
  INV_X1 U5302 ( .A(n7189), .ZN(n4830) );
  NOR2_X1 U5303 ( .A1(n9428), .A2(n9448), .ZN(n4930) );
  AND2_X1 U5304 ( .A1(n8719), .A2(n8242), .ZN(n8056) );
  NAND2_X1 U5305 ( .A1(n4948), .A2(n9096), .ZN(n4947) );
  NOR2_X1 U5306 ( .A1(n9665), .A2(n9101), .ZN(n4950) );
  AND2_X1 U5307 ( .A1(n4971), .A2(n4599), .ZN(n4967) );
  NOR2_X1 U5308 ( .A1(n7177), .A2(n4660), .ZN(n7082) );
  INV_X1 U5309 ( .A(n7174), .ZN(n4660) );
  NOR2_X1 U5310 ( .A1(n7016), .A2(n5044), .ZN(n5043) );
  INV_X1 U5311 ( .A(n7012), .ZN(n5044) );
  OR2_X1 U5312 ( .A1(n8686), .A2(n7675), .ZN(n7995) );
  AND2_X1 U5313 ( .A1(n5144), .A2(n7425), .ZN(n7427) );
  NAND2_X1 U5314 ( .A1(n7424), .A2(n7423), .ZN(n7425) );
  NOR2_X1 U5315 ( .A1(n6886), .A2(n6888), .ZN(n6887) );
  AND2_X1 U5316 ( .A1(n6890), .A2(n6889), .ZN(n6891) );
  NOR2_X1 U5317 ( .A1(n4687), .A2(n8192), .ZN(n4686) );
  AND2_X1 U5318 ( .A1(n8137), .A2(n8093), .ZN(n5014) );
  OR2_X1 U5319 ( .A1(n8695), .A2(n8083), .ZN(n8137) );
  OR2_X1 U5320 ( .A1(n7762), .A2(n9951), .ZN(n7763) );
  NAND2_X1 U5321 ( .A1(n4805), .A2(n4804), .ZN(n4803) );
  NAND2_X1 U5322 ( .A1(n7778), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n4804) );
  NAND2_X1 U5323 ( .A1(n4959), .A2(n4957), .ZN(n8093) );
  NOR2_X1 U5324 ( .A1(n6548), .A2(n4958), .ZN(n4957) );
  INV_X1 U5325 ( .A(n6539), .ZN(n4958) );
  NOR2_X1 U5326 ( .A1(n7982), .A2(n4866), .ZN(n4865) );
  INV_X1 U5327 ( .A(n7983), .ZN(n4866) );
  NAND2_X1 U5328 ( .A1(n4860), .A2(n7986), .ZN(n4863) );
  OR2_X1 U5329 ( .A1(n6334), .A2(n5092), .ZN(n5090) );
  INV_X1 U5330 ( .A(n5092), .ZN(n4631) );
  NAND2_X1 U5331 ( .A1(n10139), .A2(n6346), .ZN(n7987) );
  OR2_X1 U5332 ( .A1(n8708), .A2(n8293), .ZN(n8062) );
  AND2_X1 U5333 ( .A1(n8708), .A2(n8293), .ZN(n8064) );
  NOR2_X1 U5334 ( .A1(n8056), .A2(n4886), .ZN(n4885) );
  NAND2_X1 U5335 ( .A1(n4588), .A2(n5120), .ZN(n5114) );
  OR2_X1 U5336 ( .A1(n8719), .A2(n8242), .ZN(n8107) );
  NOR2_X1 U5337 ( .A1(n8110), .A2(n4519), .ZN(n5119) );
  OR2_X1 U5338 ( .A1(n8736), .A2(n8554), .ZN(n8039) );
  OR2_X1 U5339 ( .A1(n8666), .A2(n8597), .ZN(n8035) );
  OR2_X1 U5340 ( .A1(n8671), .A2(n8225), .ZN(n8034) );
  OR2_X1 U5341 ( .A1(n8750), .A2(n8595), .ZN(n8025) );
  OR2_X1 U5342 ( .A1(n8757), .A2(n7916), .ZN(n8024) );
  INV_X1 U5343 ( .A(n6374), .ZN(n5107) );
  NOR2_X1 U5344 ( .A1(n4531), .A2(P2_IR_REG_22__SCAN_IN), .ZN(n5103) );
  INV_X1 U5345 ( .A(n5835), .ZN(n4821) );
  AOI21_X1 U5346 ( .B1(n4522), .B2(n4839), .A(n4569), .ZN(n4836) );
  NAND3_X1 U5347 ( .A1(n6657), .A2(n5834), .A3(n7631), .ZN(n5908) );
  NOR2_X1 U5348 ( .A1(n4943), .A2(n4577), .ZN(n4940) );
  NOR2_X1 U5349 ( .A1(n4919), .A2(n4918), .ZN(n4917) );
  INV_X1 U5350 ( .A(n9069), .ZN(n4918) );
  NOR2_X1 U5351 ( .A1(n9367), .A2(n4784), .ZN(n4783) );
  INV_X1 U5352 ( .A(n5693), .ZN(n4784) );
  NOR2_X1 U5353 ( .A1(n9404), .A2(n9420), .ZN(n4656) );
  INV_X1 U5354 ( .A(n4762), .ZN(n4761) );
  OAI21_X1 U5355 ( .B1(n9103), .B2(n4763), .A(n5465), .ZN(n4762) );
  INV_X1 U5356 ( .A(n5446), .ZN(n4763) );
  NOR2_X1 U5357 ( .A1(n7601), .A2(n4643), .ZN(n4642) );
  INV_X1 U5358 ( .A(n9898), .ZN(n4643) );
  AND2_X1 U5359 ( .A1(n9113), .A2(n8990), .ZN(n4750) );
  NAND2_X1 U5360 ( .A1(n8965), .A2(n8966), .ZN(n8973) );
  OR2_X1 U5361 ( .A1(n5852), .A2(n9888), .ZN(n8966) );
  NAND2_X1 U5362 ( .A1(n5852), .A2(n9888), .ZN(n9152) );
  OR2_X1 U5363 ( .A1(n7024), .A2(n8944), .ZN(n4737) );
  INV_X1 U5364 ( .A(n9065), .ZN(n4734) );
  AND2_X1 U5365 ( .A1(n9131), .A2(n9427), .ZN(n4735) );
  OR2_X1 U5366 ( .A1(n5147), .A2(n8901), .ZN(n9579) );
  INV_X1 U5367 ( .A(n4757), .ZN(n4756) );
  OAI21_X1 U5368 ( .B1(n9115), .B2(n4758), .A(n7633), .ZN(n4757) );
  INV_X1 U5369 ( .A(n5387), .ZN(n4758) );
  AOI21_X1 U5370 ( .B1(n4991), .B2(n4993), .A(n4989), .ZN(n4988) );
  INV_X1 U5371 ( .A(n5677), .ZN(n4989) );
  NAND2_X1 U5372 ( .A1(n5645), .A2(n5644), .ZN(n5656) );
  NOR2_X1 U5373 ( .A1(n5585), .A2(n5586), .ZN(n4971) );
  AOI22_X1 U5374 ( .A1(n5586), .A2(n4970), .B1(n4972), .B2(n5585), .ZN(n4969)
         );
  INV_X1 U5375 ( .A(n5573), .ZN(n4970) );
  NAND2_X1 U5376 ( .A1(n5573), .A2(SI_20_), .ZN(n4972) );
  INV_X1 U5377 ( .A(n4975), .ZN(n4974) );
  OAI21_X1 U5378 ( .B1(n4978), .B2(n4976), .A(n5546), .ZN(n4975) );
  NAND2_X1 U5379 ( .A1(n5452), .A2(n5451), .ZN(n5468) );
  NAND2_X1 U5380 ( .A1(n5345), .A2(n5328), .ZN(n5329) );
  AOI21_X1 U5381 ( .B1(n5321), .B2(n4964), .A(n4576), .ZN(n4963) );
  INV_X1 U5382 ( .A(n5313), .ZN(n4964) );
  NAND2_X1 U5383 ( .A1(n4962), .A2(n4960), .ZN(n5346) );
  AND2_X1 U5384 ( .A1(n4963), .A2(n4961), .ZN(n4960) );
  INV_X1 U5385 ( .A(n5329), .ZN(n4961) );
  NAND2_X1 U5386 ( .A1(n4714), .A2(n4713), .ZN(n5311) );
  AOI21_X1 U5387 ( .B1(n4716), .B2(n4718), .A(n4575), .ZN(n4713) );
  NAND2_X1 U5388 ( .A1(n5271), .A2(n4716), .ZN(n4714) );
  XNOR2_X1 U5389 ( .A(n5312), .B(SI_6_), .ZN(n5309) );
  XNOR2_X1 U5390 ( .A(n5294), .B(SI_5_), .ZN(n5291) );
  INV_X1 U5391 ( .A(n7003), .ZN(n5046) );
  INV_X1 U5392 ( .A(n7004), .ZN(n5045) );
  INV_X1 U5393 ( .A(n5043), .ZN(n5041) );
  INV_X1 U5394 ( .A(n8312), .ZN(n6346) );
  INV_X1 U5395 ( .A(n8502), .ZN(n8200) );
  XNOR2_X1 U5396 ( .A(n6964), .B(n6224), .ZN(n6893) );
  AOI21_X1 U5397 ( .B1(n4542), .B2(n4697), .A(n4695), .ZN(n4694) );
  INV_X1 U5398 ( .A(n8188), .ZN(n8239) );
  AOI21_X1 U5399 ( .B1(n7911), .B2(n8608), .A(n4664), .ZN(n4662) );
  NAND2_X1 U5400 ( .A1(n4666), .A2(n4665), .ZN(n4664) );
  NAND2_X1 U5401 ( .A1(n7910), .A2(n8608), .ZN(n4665) );
  NAND2_X1 U5402 ( .A1(n8182), .A2(n8181), .ZN(n8248) );
  NAND2_X1 U5403 ( .A1(n6176), .A2(n6175), .ZN(n6470) );
  NOR2_X1 U5404 ( .A1(n4671), .A2(n7426), .ZN(n4668) );
  AND2_X1 U5405 ( .A1(n7458), .A2(n5070), .ZN(n5069) );
  NAND2_X1 U5406 ( .A1(n7571), .A2(n8309), .ZN(n5070) );
  NOR2_X1 U5407 ( .A1(n7571), .A2(n8309), .ZN(n5068) );
  AND2_X1 U5408 ( .A1(n5066), .A2(n7436), .ZN(n4670) );
  XNOR2_X1 U5409 ( .A(n10120), .B(n8189), .ZN(n7084) );
  INV_X1 U5410 ( .A(n4686), .ZN(n4683) );
  AOI21_X1 U5411 ( .B1(n4686), .B2(n4682), .A(n4688), .ZN(n4681) );
  INV_X1 U5412 ( .A(n8238), .ZN(n4682) );
  NOR2_X1 U5413 ( .A1(n4691), .A2(n4689), .ZN(n4688) );
  NAND2_X1 U5414 ( .A1(n7623), .A2(n5075), .ZN(n5074) );
  NAND2_X1 U5415 ( .A1(n4800), .A2(n4799), .ZN(n4798) );
  NAND2_X1 U5416 ( .A1(n6763), .A2(n6779), .ZN(n4801) );
  INV_X1 U5417 ( .A(n4814), .ZN(n5139) );
  OR2_X1 U5418 ( .A1(n10011), .A2(n10010), .ZN(n4805) );
  XNOR2_X1 U5419 ( .A(n4803), .B(n4802), .ZN(n10025) );
  XNOR2_X1 U5420 ( .A(n8324), .B(n8321), .ZN(n7797) );
  OR2_X1 U5421 ( .A1(n8323), .A2(n7825), .ZN(n4808) );
  OR2_X1 U5422 ( .A1(n4537), .A2(n8323), .ZN(n4807) );
  NAND2_X1 U5423 ( .A1(n6181), .A2(n6180), .ZN(n6519) );
  NAND2_X1 U5424 ( .A1(n6172), .A2(n10299), .ZN(n6426) );
  INV_X1 U5425 ( .A(n6414), .ZN(n6172) );
  AOI21_X1 U5426 ( .B1(n4865), .B2(n4863), .A(n4862), .ZN(n4861) );
  INV_X1 U5427 ( .A(n4865), .ZN(n4864) );
  INV_X1 U5428 ( .A(n4863), .ZN(n4868) );
  NAND2_X1 U5429 ( .A1(n5026), .A2(n5024), .ZN(n7983) );
  NOR2_X1 U5430 ( .A1(n6346), .A2(n5025), .ZN(n5024) );
  INV_X1 U5431 ( .A(n6337), .ZN(n5025) );
  NAND2_X1 U5432 ( .A1(n6696), .A2(n6203), .ZN(n5026) );
  NAND2_X1 U5433 ( .A1(n4870), .A2(n4869), .ZN(n7395) );
  AOI21_X1 U5434 ( .B1(n4871), .B2(n4874), .A(n6320), .ZN(n4869) );
  INV_X1 U5435 ( .A(n7975), .ZN(n4874) );
  NAND2_X1 U5436 ( .A1(n7120), .A2(n7970), .ZN(n7287) );
  INV_X1 U5437 ( .A(n8111), .ZN(n6981) );
  NAND2_X1 U5438 ( .A1(n6587), .A2(n4560), .ZN(n4898) );
  NAND2_X1 U5439 ( .A1(n4582), .A2(n6587), .ZN(n4897) );
  NAND2_X1 U5440 ( .A1(n8159), .A2(n6203), .ZN(n4959) );
  NAND2_X1 U5441 ( .A1(n5134), .A2(n5133), .ZN(n8493) );
  OR2_X1 U5442 ( .A1(n8500), .A2(n6527), .ZN(n5134) );
  INV_X1 U5443 ( .A(n4876), .ZN(n4875) );
  OAI21_X1 U5444 ( .B1(n4877), .B2(n6576), .A(n8059), .ZN(n4876) );
  AOI21_X1 U5445 ( .B1(n4883), .B2(n4885), .A(n4882), .ZN(n4881) );
  INV_X1 U5446 ( .A(n8107), .ZN(n4882) );
  INV_X1 U5447 ( .A(n4888), .ZN(n4883) );
  INV_X1 U5448 ( .A(n4885), .ZN(n4884) );
  AND2_X1 U5449 ( .A1(n8060), .A2(n8059), .ZN(n8514) );
  NAND2_X1 U5450 ( .A1(n8725), .A2(n8541), .ZN(n5120) );
  NOR2_X1 U5451 ( .A1(n4889), .A2(n8109), .ZN(n4888) );
  INV_X1 U5452 ( .A(n8047), .ZN(n4889) );
  NAND2_X1 U5453 ( .A1(n6479), .A2(n6478), .ZN(n8175) );
  NOR2_X1 U5454 ( .A1(n5102), .A2(n5095), .ZN(n5094) );
  INV_X1 U5455 ( .A(n5097), .ZN(n5095) );
  NAND2_X1 U5456 ( .A1(n6413), .A2(n6412), .ZN(n8682) );
  NAND2_X1 U5457 ( .A1(n5106), .A2(n6386), .ZN(n7736) );
  INV_X1 U5458 ( .A(n8598), .ZN(n8620) );
  INV_X1 U5459 ( .A(n8596), .ZN(n8618) );
  AND4_X1 U5460 ( .A1(n6397), .A2(n6396), .A3(n6395), .A4(n6394), .ZN(n7734)
         );
  NAND2_X2 U5461 ( .A1(n6559), .A2(n6644), .ZN(n8623) );
  NAND2_X1 U5462 ( .A1(n6606), .A2(n6607), .ZN(n6674) );
  NAND2_X1 U5463 ( .A1(n6594), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6598) );
  OR2_X1 U5464 ( .A1(n6279), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n6286) );
  NAND2_X1 U5465 ( .A1(n6246), .A2(n4818), .ZN(n4817) );
  NAND2_X1 U5466 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n4819) );
  AOI22_X1 U5467 ( .A1(n4508), .A2(n5840), .B1(n6071), .B2(n6958), .ZN(n5841)
         );
  AOI21_X1 U5468 ( .B1(n4848), .B2(n4845), .A(n4584), .ZN(n4844) );
  INV_X1 U5469 ( .A(n6008), .ZN(n4845) );
  INV_X1 U5470 ( .A(n4848), .ZN(n4846) );
  NAND2_X1 U5471 ( .A1(n7140), .A2(n7142), .ZN(n4832) );
  NAND2_X1 U5472 ( .A1(n4510), .A2(n5884), .ZN(n7141) );
  AOI21_X1 U5473 ( .B1(n4852), .B2(n6048), .A(n6061), .ZN(n4851) );
  OR2_X1 U5474 ( .A1(n8939), .A2(n8940), .ZN(n6061) );
  OR4_X1 U5475 ( .A1(n9209), .A2(n9137), .A3(n9218), .A4(n9136), .ZN(n9225) );
  CLKBUF_X1 U5476 ( .A(n5264), .Z(n5731) );
  INV_X1 U5477 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n5155) );
  INV_X1 U5478 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n4915) );
  INV_X1 U5479 ( .A(n5792), .ZN(n6120) );
  AND2_X1 U5480 ( .A1(n9080), .A2(n9073), .ZN(n9135) );
  NOR2_X1 U5481 ( .A1(n9135), .A2(n4781), .ZN(n4780) );
  INV_X1 U5482 ( .A(n5708), .ZN(n4781) );
  OAI21_X1 U5483 ( .B1(n9397), .B2(n5674), .A(n5673), .ZN(n9382) );
  AND2_X1 U5484 ( .A1(n9142), .A2(n9188), .ZN(n9412) );
  AOI21_X1 U5485 ( .B1(n4771), .B2(n4770), .A(n4545), .ZN(n4769) );
  INV_X1 U5486 ( .A(n5636), .ZN(n4771) );
  AND2_X1 U5487 ( .A1(n5615), .A2(n5614), .ZN(n4770) );
  NOR2_X1 U5488 ( .A1(n5636), .A2(n4773), .ZN(n4772) );
  INV_X1 U5489 ( .A(n5614), .ZN(n4773) );
  INV_X1 U5490 ( .A(n9131), .ZN(n9428) );
  OAI21_X1 U5491 ( .B1(n5571), .B2(n4788), .A(n4785), .ZN(n5600) );
  INV_X1 U5492 ( .A(n4791), .ZN(n4788) );
  NAND2_X1 U5493 ( .A1(n5571), .A2(n5142), .ZN(n4793) );
  OAI21_X1 U5494 ( .B1(n9510), .B2(n5543), .A(n5542), .ZN(n9498) );
  NOR2_X1 U5495 ( .A1(n9554), .A2(n9537), .ZN(n9536) );
  AOI21_X1 U5496 ( .B1(n4747), .B2(n4746), .A(n4745), .ZN(n4744) );
  INV_X1 U5497 ( .A(n9006), .ZN(n4746) );
  INV_X1 U5498 ( .A(n9014), .ZN(n4745) );
  NAND2_X1 U5499 ( .A1(n7489), .A2(n9115), .ZN(n7488) );
  NOR2_X1 U5500 ( .A1(n4644), .A2(n7538), .ZN(n7639) );
  OR2_X1 U5501 ( .A1(n9262), .A2(n7409), .ZN(n8990) );
  OAI22_X1 U5502 ( .A1(n7213), .A2(n9111), .B1(n7219), .B2(n9262), .ZN(n7238)
         );
  INV_X1 U5503 ( .A(n7212), .ZN(n9111) );
  NAND2_X1 U5504 ( .A1(n5713), .A2(n5712), .ZN(n6119) );
  INV_X1 U5505 ( .A(n5234), .ZN(n5560) );
  XNOR2_X1 U5506 ( .A(n7939), .B(n7938), .ZN(n8961) );
  NAND2_X1 U5507 ( .A1(n8074), .A2(n7935), .ZN(n7939) );
  NAND2_X1 U5508 ( .A1(n8074), .A2(n8073), .ZN(n9091) );
  OR2_X1 U5509 ( .A1(n8072), .A2(n8071), .ZN(n8073) );
  NAND2_X1 U5510 ( .A1(n5696), .A2(n5695), .ZN(n5698) );
  INV_X1 U5511 ( .A(n5709), .ZN(n5008) );
  XNOR2_X1 U5512 ( .A(n5676), .B(n5675), .ZN(n8784) );
  NAND2_X1 U5513 ( .A1(n5656), .A2(n5655), .ZN(n5676) );
  NAND2_X1 U5514 ( .A1(n5626), .A2(n5625), .ZN(n5638) );
  OAI21_X1 U5515 ( .B1(n5490), .B2(n4981), .A(n4979), .ZN(n5548) );
  NAND2_X1 U5516 ( .A1(n4984), .A2(n4985), .ZN(n5529) );
  NAND2_X1 U5517 ( .A1(n5490), .A2(n4986), .ZN(n4984) );
  OAI21_X1 U5518 ( .B1(n5490), .B2(n5489), .A(n5488), .ZN(n5506) );
  OAI21_X1 U5519 ( .B1(n5370), .B2(n4520), .A(n4996), .ZN(n5430) );
  XNOR2_X1 U5520 ( .A(n5410), .B(n5409), .ZN(n6718) );
  NAND2_X1 U5521 ( .A1(n4999), .A2(n5391), .ZN(n5410) );
  NAND2_X1 U5522 ( .A1(n5370), .A2(n5000), .ZN(n4999) );
  NAND2_X1 U5523 ( .A1(n7088), .A2(n7087), .ZN(n7424) );
  NOR2_X1 U5524 ( .A1(n4530), .A2(n8267), .ZN(n5055) );
  NAND2_X1 U5525 ( .A1(n5058), .A2(n5063), .ZN(n5057) );
  NAND2_X1 U5526 ( .A1(n8197), .A2(n5064), .ZN(n5063) );
  NAND2_X1 U5527 ( .A1(n6529), .A2(n6528), .ZN(n8635) );
  NAND2_X1 U5528 ( .A1(n5081), .A2(n5079), .ZN(n8250) );
  NAND2_X1 U5529 ( .A1(n5083), .A2(n5080), .ZN(n5079) );
  NOR2_X1 U5530 ( .A1(n8247), .A2(n8183), .ZN(n5082) );
  NAND2_X1 U5531 ( .A1(n4618), .A2(n8092), .ZN(n4616) );
  NAND2_X1 U5532 ( .A1(n6537), .A2(n6536), .ZN(n8494) );
  INV_X1 U5533 ( .A(n8242), .ZN(n8534) );
  NAND2_X1 U5534 ( .A1(n6496), .A2(n6495), .ZN(n8533) );
  NAND4_X1 U5535 ( .A1(n6300), .A2(n6299), .A3(n6298), .A4(n6297), .ZN(n8315)
         );
  NAND2_X1 U5536 ( .A1(n4539), .A2(n5085), .ZN(n5084) );
  OAI21_X1 U5537 ( .B1(n4811), .B2(n8420), .A(n8443), .ZN(n4810) );
  NAND2_X1 U5538 ( .A1(n6488), .A2(n6487), .ZN(n8547) );
  AND2_X1 U5539 ( .A1(n10103), .A2(n7285), .ZN(n8562) );
  INV_X1 U5540 ( .A(n8560), .ZN(n8627) );
  NAND2_X1 U5541 ( .A1(n6160), .A2(n6159), .ZN(n8702) );
  AOI21_X1 U5542 ( .B1(n4636), .B2(n8623), .A(n4633), .ZN(n8700) );
  NAND2_X1 U5543 ( .A1(n4635), .A2(n4634), .ZN(n4633) );
  XNOR2_X1 U5544 ( .A(n8493), .B(n8492), .ZN(n4636) );
  NAND2_X1 U5545 ( .A1(n8509), .A2(n8618), .ZN(n4634) );
  NAND2_X1 U5546 ( .A1(n6391), .A2(n6390), .ZN(n8005) );
  XNOR2_X1 U5547 ( .A(n6459), .B(n6550), .ZN(n8463) );
  NAND2_X1 U5548 ( .A1(n5577), .A2(n5576), .ZN(n9485) );
  AND2_X1 U5549 ( .A1(n6094), .A2(n6085), .ZN(n8942) );
  AND2_X1 U5550 ( .A1(n6094), .A2(n9233), .ZN(n9764) );
  NAND2_X1 U5551 ( .A1(n4935), .A2(n4934), .ZN(n4933) );
  NAND2_X1 U5552 ( .A1(n4938), .A2(n4932), .ZN(n4931) );
  INV_X1 U5553 ( .A(n4625), .ZN(n4624) );
  OAI21_X1 U5554 ( .B1(n9220), .B2(n9230), .A(n9098), .ZN(n4625) );
  NOR2_X1 U5555 ( .A1(n4949), .A2(n8983), .ZN(n4626) );
  NOR2_X1 U5556 ( .A1(n9332), .A2(n9578), .ZN(n9586) );
  NAND2_X1 U5557 ( .A1(n5730), .A2(n5729), .ZN(n9349) );
  INV_X1 U5558 ( .A(n9351), .ZN(n5794) );
  INV_X1 U5559 ( .A(n9350), .ZN(n5795) );
  OR2_X1 U5560 ( .A1(n7953), .A2(n10109), .ZN(n7962) );
  NAND2_X1 U5561 ( .A1(n4613), .A2(n4612), .ZN(n7973) );
  NAND2_X1 U5562 ( .A1(n4615), .A2(n4614), .ZN(n4613) );
  INV_X1 U5563 ( .A(n7959), .ZN(n4615) );
  NAND2_X1 U5564 ( .A1(n7961), .A2(n7960), .ZN(n4614) );
  NAND2_X1 U5565 ( .A1(n4726), .A2(n4724), .ZN(n7981) );
  NAND2_X1 U5566 ( .A1(n7983), .A2(n4549), .ZN(n4724) );
  NOR2_X1 U5567 ( .A1(n7994), .A2(n8090), .ZN(n5027) );
  AOI21_X1 U5568 ( .B1(n8971), .B2(n8970), .A(n8969), .ZN(n8982) );
  NOR2_X1 U5569 ( .A1(n4906), .A2(n8983), .ZN(n4905) );
  INV_X1 U5570 ( .A(n5146), .ZN(n4906) );
  INV_X1 U5571 ( .A(n9162), .ZN(n4907) );
  INV_X1 U5572 ( .A(n8007), .ZN(n5021) );
  INV_X1 U5573 ( .A(n8006), .ZN(n5023) );
  OR2_X1 U5574 ( .A1(n9003), .A2(n9002), .ZN(n9009) );
  INV_X1 U5575 ( .A(n8032), .ZN(n5036) );
  INV_X1 U5576 ( .A(n8033), .ZN(n5037) );
  AOI21_X1 U5577 ( .B1(n8023), .B2(n8022), .A(n8606), .ZN(n8028) );
  NOR2_X1 U5578 ( .A1(n8037), .A2(n8087), .ZN(n5033) );
  NOR2_X1 U5579 ( .A1(n8031), .A2(n8090), .ZN(n5031) );
  OR3_X1 U5580 ( .A1(n9024), .A2(n9023), .A3(n9175), .ZN(n9029) );
  AND2_X1 U5581 ( .A1(n4711), .A2(n8090), .ZN(n4704) );
  AND2_X1 U5582 ( .A1(n8548), .A2(n8045), .ZN(n4711) );
  AND2_X1 U5583 ( .A1(n4708), .A2(n8087), .ZN(n4701) );
  OAI21_X1 U5584 ( .B1(n4705), .B2(n8090), .A(n4703), .ZN(n4702) );
  NOR2_X1 U5585 ( .A1(n8049), .A2(n4709), .ZN(n4708) );
  NAND2_X1 U5586 ( .A1(n4930), .A2(n4925), .ZN(n4924) );
  INV_X1 U5587 ( .A(n4927), .ZN(n4925) );
  AOI21_X1 U5588 ( .B1(n9057), .B2(n9058), .A(n4928), .ZN(n4927) );
  AOI21_X1 U5589 ( .B1(n5006), .B2(n5008), .A(n5005), .ZN(n5004) );
  INV_X1 U5590 ( .A(n5723), .ZN(n5005) );
  INV_X1 U5591 ( .A(n6577), .ZN(n4895) );
  NOR2_X1 U5592 ( .A1(n4895), .A2(n4892), .ZN(n4891) );
  INV_X1 U5593 ( .A(n8067), .ZN(n4892) );
  AND2_X1 U5594 ( .A1(n4829), .A2(n5884), .ZN(n4826) );
  NAND2_X1 U5595 ( .A1(n4587), .A2(n4829), .ZN(n4822) );
  INV_X1 U5596 ( .A(n5899), .ZN(n4831) );
  OR2_X1 U5597 ( .A1(n8835), .A2(n4839), .ZN(n4838) );
  INV_X1 U5598 ( .A(n5949), .ZN(n4839) );
  MUX2_X1 U5599 ( .A(n9052), .B(n9051), .S(n9096), .Z(n9059) );
  NOR2_X1 U5600 ( .A1(n4926), .A2(n4922), .ZN(n4921) );
  INV_X1 U5601 ( .A(n4930), .ZN(n4926) );
  NAND2_X1 U5602 ( .A1(n9412), .A2(n9057), .ZN(n4922) );
  NOR2_X1 U5603 ( .A1(n4923), .A2(n4920), .ZN(n4919) );
  INV_X1 U5604 ( .A(n9412), .ZN(n4920) );
  AND2_X1 U5605 ( .A1(n4929), .A2(n4924), .ZN(n4923) );
  INV_X1 U5606 ( .A(n9068), .ZN(n4929) );
  OR2_X1 U5607 ( .A1(n9349), .A2(n6939), .ZN(n9202) );
  INV_X1 U5608 ( .A(n4992), .ZN(n4991) );
  OAI21_X1 U5609 ( .B1(n5644), .B2(n4993), .A(n5675), .ZN(n4992) );
  INV_X1 U5610 ( .A(n5655), .ZN(n4993) );
  NAND2_X1 U5611 ( .A1(n4981), .A2(n5544), .ZN(n4976) );
  NOR2_X1 U5612 ( .A1(n4978), .A2(n5547), .ZN(n4977) );
  INV_X1 U5613 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n5324) );
  INV_X1 U5614 ( .A(n4717), .ZN(n4716) );
  OAI21_X1 U5615 ( .B1(n5270), .B2(n4718), .A(n5292), .ZN(n4717) );
  INV_X1 U5616 ( .A(n5291), .ZN(n5292) );
  INV_X1 U5617 ( .A(n5274), .ZN(n4718) );
  INV_X1 U5618 ( .A(n8195), .ZN(n5062) );
  INV_X1 U5619 ( .A(n8258), .ZN(n4695) );
  INV_X1 U5620 ( .A(n7914), .ZN(n4666) );
  NAND2_X1 U5621 ( .A1(n4681), .A2(n4683), .ZN(n4680) );
  INV_X1 U5622 ( .A(n8089), .ZN(n5013) );
  NAND2_X1 U5623 ( .A1(n10001), .A2(n7790), .ZN(n7791) );
  NAND2_X1 U5624 ( .A1(n10034), .A2(n7793), .ZN(n7794) );
  OAI21_X1 U5625 ( .B1(n8350), .B2(n10395), .A(n8349), .ZN(n8376) );
  NAND2_X1 U5626 ( .A1(n8401), .A2(n4620), .ZN(n8429) );
  NAND2_X1 U5627 ( .A1(n8399), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n4620) );
  NAND2_X1 U5628 ( .A1(n8592), .A2(n6457), .ZN(n5101) );
  INV_X1 U5629 ( .A(n8314), .ZN(n7161) );
  NAND2_X1 U5630 ( .A1(n8313), .A2(n4725), .ZN(n7979) );
  INV_X1 U5631 ( .A(n10134), .ZN(n4725) );
  AOI21_X1 U5632 ( .B1(n7975), .B2(n4873), .A(n4872), .ZN(n4871) );
  INV_X1 U5633 ( .A(n7970), .ZN(n4873) );
  NAND2_X1 U5634 ( .A1(n5127), .A2(n6538), .ZN(n5124) );
  AOI21_X1 U5635 ( .B1(n5123), .B2(n6538), .A(n5130), .ZN(n5122) );
  AND2_X1 U5636 ( .A1(n8635), .A2(n8494), .ZN(n5130) );
  INV_X1 U5637 ( .A(n5126), .ZN(n5123) );
  NAND2_X1 U5638 ( .A1(n8708), .A2(n8509), .ZN(n5133) );
  NAND2_X1 U5639 ( .A1(n4881), .A2(n4884), .ZN(n4877) );
  NOR2_X1 U5640 ( .A1(n4880), .A2(n6576), .ZN(n4879) );
  INV_X1 U5641 ( .A(n4881), .ZN(n4880) );
  NOR2_X1 U5642 ( .A1(n5114), .A2(n5112), .ZN(n5111) );
  INV_X1 U5643 ( .A(n5118), .ZN(n5112) );
  NAND2_X1 U5644 ( .A1(n6398), .A2(n6148), .ZN(n5088) );
  AOI21_X1 U5645 ( .B1(n4523), .B2(n4846), .A(n4557), .ZN(n4840) );
  NOR2_X1 U5646 ( .A1(n4946), .A2(n4937), .ZN(n4936) );
  INV_X1 U5647 ( .A(n9089), .ZN(n4937) );
  AND2_X1 U5648 ( .A1(n9674), .A2(n4656), .ZN(n4655) );
  AND2_X1 U5649 ( .A1(n4786), .A2(n4789), .ZN(n4785) );
  NAND2_X1 U5650 ( .A1(n4791), .A2(n4787), .ZN(n4786) );
  AND2_X1 U5651 ( .A1(n4543), .A2(n5583), .ZN(n4789) );
  INV_X1 U5652 ( .A(n5142), .ZN(n4787) );
  NOR2_X1 U5653 ( .A1(n9470), .A2(n4648), .ZN(n4647) );
  INV_X1 U5654 ( .A(n4649), .ZN(n4648) );
  NOR2_X1 U5655 ( .A1(n9485), .A2(n9502), .ZN(n4649) );
  OR2_X1 U5656 ( .A1(n9264), .A2(n9893), .ZN(n9155) );
  NAND2_X1 U5657 ( .A1(n6958), .A2(n4752), .ZN(n5765) );
  NAND2_X1 U5658 ( .A1(n9153), .A2(n5765), .ZN(n9107) );
  NAND2_X1 U5659 ( .A1(n9236), .A2(n9230), .ZN(n5836) );
  NAND2_X1 U5660 ( .A1(n9433), .A2(n4653), .ZN(n9373) );
  AND2_X1 U5661 ( .A1(n4655), .A2(n4654), .ZN(n4653) );
  NAND2_X1 U5662 ( .A1(n9433), .A2(n9682), .ZN(n9417) );
  AND2_X1 U5663 ( .A1(n9686), .A2(n9450), .ZN(n9433) );
  NAND2_X1 U5664 ( .A1(n4639), .A2(n4638), .ZN(n4637) );
  AND2_X1 U5665 ( .A1(n9099), .A2(n4621), .ZN(n9096) );
  NOR2_X1 U5666 ( .A1(n7105), .A2(n7112), .ZN(n7278) );
  OAI21_X1 U5667 ( .B1(n7931), .B2(SI_29_), .A(n7930), .ZN(n8072) );
  NAND2_X1 U5668 ( .A1(n5638), .A2(n5637), .ZN(n5645) );
  AOI21_X1 U5669 ( .B1(n4969), .B2(n4967), .A(n4601), .ZN(n4966) );
  NAND2_X1 U5670 ( .A1(n4969), .A2(n4599), .ZN(n4968) );
  AOI21_X1 U5671 ( .B1(n4982), .B2(n4987), .A(n4980), .ZN(n4979) );
  INV_X1 U5672 ( .A(n5527), .ZN(n4980) );
  INV_X1 U5673 ( .A(n4982), .ZN(n4981) );
  AOI21_X1 U5674 ( .B1(n4986), .B2(n5489), .A(n4574), .ZN(n4985) );
  AND2_X1 U5675 ( .A1(n5485), .A2(SI_15_), .ZN(n5489) );
  INV_X1 U5676 ( .A(n4997), .ZN(n4996) );
  OAI21_X1 U5677 ( .B1(n5000), .B2(n4520), .A(n5408), .ZN(n4997) );
  NAND2_X1 U5678 ( .A1(n5390), .A2(SI_10_), .ZN(n5391) );
  NOR2_X1 U5679 ( .A1(n5392), .A2(n5001), .ZN(n5000) );
  INV_X1 U5680 ( .A(n5369), .ZN(n5001) );
  INV_X1 U5681 ( .A(n5388), .ZN(n5392) );
  NOR2_X2 U5682 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n5373) );
  XNOR2_X1 U5683 ( .A(n5389), .B(SI_10_), .ZN(n5388) );
  NAND2_X1 U5684 ( .A1(n7936), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n5002) );
  INV_X1 U5685 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4951) );
  AOI21_X1 U5686 ( .B1(n8238), .B2(n8239), .A(n4555), .ZN(n4691) );
  NAND2_X1 U5687 ( .A1(n5053), .A2(n5052), .ZN(n6894) );
  NAND2_X1 U5688 ( .A1(n6891), .A2(n4553), .ZN(n5053) );
  NOR2_X1 U5689 ( .A1(n8247), .A2(n8541), .ZN(n5080) );
  NAND2_X1 U5690 ( .A1(n4586), .A2(n8248), .ZN(n8212) );
  NAND2_X1 U5691 ( .A1(n5046), .A2(n5045), .ZN(n7013) );
  XNOR2_X1 U5692 ( .A(n10139), .B(n8196), .ZN(n7418) );
  NAND2_X1 U5693 ( .A1(n7428), .A2(n8311), .ZN(n7438) );
  OAI211_X1 U5694 ( .C1(n6891), .C2(n4509), .A(n5050), .B(n5049), .ZN(n6964)
         );
  NAND2_X1 U5695 ( .A1(n6225), .A2(n5051), .ZN(n5050) );
  OR3_X1 U5696 ( .A1(n6896), .A2(n10147), .A3(n8090), .ZN(n6895) );
  INV_X1 U5697 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n6142) );
  AND2_X1 U5698 ( .A1(n7331), .A2(n7330), .ZN(n8082) );
  OR2_X1 U5699 ( .A1(n9925), .A2(n7225), .ZN(n9927) );
  INV_X1 U5700 ( .A(n4797), .ZN(n4796) );
  NAND2_X1 U5701 ( .A1(n4797), .A2(n4801), .ZN(n6787) );
  NAND2_X1 U5702 ( .A1(n7782), .A2(n7781), .ZN(n7783) );
  NAND2_X1 U5703 ( .A1(n7765), .A2(n9961), .ZN(n9966) );
  NAND2_X1 U5704 ( .A1(n10002), .A2(n10003), .ZN(n10001) );
  INV_X1 U5705 ( .A(n4803), .ZN(n7769) );
  NAND2_X1 U5706 ( .A1(n10035), .A2(n10036), .ZN(n10034) );
  NOR2_X1 U5707 ( .A1(n10060), .A2(n4629), .ZN(n10087) );
  AND2_X1 U5708 ( .A1(n7774), .A2(n10050), .ZN(n4629) );
  NOR2_X1 U5709 ( .A1(n10087), .A2(n10086), .ZN(n10085) );
  NAND2_X1 U5710 ( .A1(n7797), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n8326) );
  AND3_X1 U5711 ( .A1(n4806), .A2(n4807), .A3(n4608), .ZN(n8370) );
  NOR2_X1 U5712 ( .A1(n8402), .A2(n8624), .ZN(n4628) );
  XNOR2_X1 U5713 ( .A(n8429), .B(n8424), .ZN(n8403) );
  INV_X1 U5714 ( .A(n5088), .ZN(n5085) );
  OR2_X1 U5715 ( .A1(n8418), .A2(n8419), .ZN(n4813) );
  NAND2_X1 U5716 ( .A1(n6179), .A2(n6178), .ZN(n6510) );
  INV_X1 U5717 ( .A(n6501), .ZN(n6179) );
  AND2_X1 U5718 ( .A1(n5101), .A2(n4550), .ZN(n8577) );
  AND2_X1 U5719 ( .A1(n5101), .A2(n5100), .ZN(n8578) );
  AND3_X1 U5720 ( .A1(n6444), .A2(n6443), .A3(n6442), .ZN(n8595) );
  AND3_X1 U5721 ( .A1(n6467), .A2(n6466), .A3(n6465), .ZN(n8597) );
  NAND2_X1 U5722 ( .A1(n6174), .A2(n6173), .ZN(n6453) );
  INV_X1 U5723 ( .A(n6438), .ZN(n6174) );
  NAND2_X1 U5724 ( .A1(n6171), .A2(n6170), .ZN(n6402) );
  INV_X1 U5725 ( .A(n6392), .ZN(n6171) );
  NAND2_X1 U5726 ( .A1(n4861), .A2(n4864), .ZN(n4858) );
  AND2_X1 U5727 ( .A1(n5090), .A2(n6348), .ZN(n5091) );
  NAND2_X1 U5728 ( .A1(n6168), .A2(n6167), .ZN(n6357) );
  INV_X1 U5729 ( .A(n6339), .ZN(n6168) );
  NAND2_X1 U5730 ( .A1(n7397), .A2(n6335), .ZN(n7449) );
  OR2_X1 U5731 ( .A1(n6327), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n6339) );
  OR2_X1 U5732 ( .A1(n10128), .A2(n7161), .ZN(n7394) );
  NAND2_X1 U5733 ( .A1(n7316), .A2(n6334), .ZN(n7397) );
  NAND2_X1 U5734 ( .A1(n6166), .A2(n6165), .ZN(n6327) );
  INV_X1 U5735 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n6165) );
  INV_X1 U5736 ( .A(n6313), .ZN(n6166) );
  OR2_X1 U5737 ( .A1(n6295), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n6313) );
  AND4_X1 U5738 ( .A1(n6260), .A2(n6259), .A3(n6258), .A4(n6257), .ZN(n7123)
         );
  NAND2_X1 U5739 ( .A1(n6162), .A2(n6161), .ZN(n6272) );
  INV_X1 U5740 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n6162) );
  NAND2_X1 U5741 ( .A1(n6164), .A2(n6163), .ZN(n6295) );
  INV_X1 U5742 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n6163) );
  INV_X1 U5743 ( .A(n6272), .ZN(n6164) );
  NAND2_X1 U5744 ( .A1(n6580), .A2(n7201), .ZN(n7520) );
  AND2_X1 U5745 ( .A1(n7513), .A2(n8444), .ZN(n7942) );
  AND3_X1 U5746 ( .A1(n6877), .A2(n6630), .A3(n6641), .ZN(n7197) );
  AND2_X1 U5747 ( .A1(n8087), .A2(n6608), .ZN(n7198) );
  AND2_X1 U5748 ( .A1(n8470), .A2(n8469), .ZN(n8692) );
  NAND2_X1 U5749 ( .A1(n8494), .A2(n8620), .ZN(n4635) );
  AND2_X1 U5750 ( .A1(n8058), .A2(n8062), .ZN(n8501) );
  INV_X1 U5751 ( .A(n5100), .ZN(n5099) );
  AND4_X1 U5752 ( .A1(n6373), .A2(n6372), .A3(n6371), .A4(n6370), .ZN(n7675)
         );
  INV_X1 U5753 ( .A(n10147), .ZN(n10119) );
  NAND2_X1 U5754 ( .A1(n6157), .A2(n6155), .ZN(n5089) );
  NAND2_X1 U5755 ( .A1(n4674), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6156) );
  NOR2_X1 U5756 ( .A1(P2_IR_REG_27__SCAN_IN), .A2(P2_IR_REG_26__SCAN_IN), .ZN(
        n4673) );
  INV_X1 U5757 ( .A(n6582), .ZN(n8450) );
  NAND2_X1 U5758 ( .A1(n6557), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6553) );
  NOR2_X1 U5759 ( .A1(n6388), .A2(n5086), .ZN(n6551) );
  NAND2_X1 U5760 ( .A1(n4539), .A2(n5087), .ZN(n5086) );
  NOR2_X1 U5761 ( .A1(n5088), .A2(P2_IR_REG_18__SCAN_IN), .ZN(n5087) );
  NOR2_X1 U5762 ( .A1(n6388), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n6399) );
  AND2_X1 U5763 ( .A1(n6309), .A2(n6322), .ZN(n7787) );
  NOR2_X1 U5764 ( .A1(n5302), .A2(n5301), .ZN(n5337) );
  INV_X1 U5765 ( .A(n8845), .ZN(n4852) );
  AOI21_X1 U5766 ( .B1(n9263), .B2(n6068), .A(n5868), .ZN(n5873) );
  XNOR2_X1 U5767 ( .A(n5864), .B(n6066), .ZN(n5869) );
  AND2_X1 U5768 ( .A1(n5337), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n5361) );
  OR2_X1 U5769 ( .A1(n5578), .A2(n8890), .ZN(n5593) );
  AND2_X1 U5770 ( .A1(n4596), .A2(n4939), .ZN(n4938) );
  NAND2_X1 U5771 ( .A1(n4540), .A2(n4940), .ZN(n4939) );
  NAND2_X1 U5772 ( .A1(n4945), .A2(n4948), .ZN(n4941) );
  NAND2_X1 U5773 ( .A1(n4936), .A2(n9136), .ZN(n4932) );
  AOI211_X1 U5774 ( .C1(n9077), .C2(n9145), .A(n9076), .B(n9075), .ZN(n9079)
         );
  NAND2_X1 U5775 ( .A1(n4540), .A2(n4942), .ZN(n4934) );
  INV_X1 U5776 ( .A(n4943), .ZN(n4942) );
  INV_X1 U5777 ( .A(n4936), .ZN(n4935) );
  INV_X1 U5778 ( .A(n8944), .ZN(n9232) );
  AND2_X1 U5779 ( .A1(n5692), .A2(n5691), .ZN(n6056) );
  AND4_X1 U5780 ( .A1(n5445), .A2(n5444), .A3(n5443), .A4(n5442), .ZN(n7605)
         );
  AND4_X1 U5781 ( .A1(n5425), .A2(n5424), .A3(n5423), .A4(n5422), .ZN(n7700)
         );
  AND4_X1 U5782 ( .A1(n5386), .A2(n5385), .A3(n5384), .A4(n5383), .ZN(n7634)
         );
  AND4_X1 U5783 ( .A1(n5367), .A2(n5366), .A3(n5365), .A4(n5364), .ZN(n7484)
         );
  AND4_X1 U5784 ( .A1(n5343), .A2(n5342), .A3(n5341), .A4(n5340), .ZN(n7498)
         );
  OR2_X1 U5785 ( .A1(n6709), .A2(n5167), .ZN(n5174) );
  INV_X1 U5786 ( .A(n9230), .ZN(n5833) );
  INV_X1 U5787 ( .A(n4783), .ZN(n4778) );
  AOI21_X1 U5788 ( .B1(n9368), .B2(n9367), .A(n5790), .ZN(n6116) );
  AND2_X1 U5789 ( .A1(n9081), .A2(n9072), .ZN(n9367) );
  NAND2_X1 U5790 ( .A1(n9078), .A2(n9195), .ZN(n9384) );
  NAND2_X1 U5791 ( .A1(n9433), .A2(n4655), .ZN(n9390) );
  OAI21_X1 U5792 ( .B1(n9449), .B2(n4767), .A(n4764), .ZN(n9397) );
  AOI21_X1 U5793 ( .B1(n4766), .B2(n4765), .A(n4572), .ZN(n4764) );
  INV_X1 U5794 ( .A(n4772), .ZN(n4765) );
  AND2_X1 U5795 ( .A1(n9145), .A2(n9189), .ZN(n9399) );
  INV_X1 U5796 ( .A(n9448), .ZN(n4736) );
  AND2_X1 U5797 ( .A1(n9517), .A2(n4645), .ZN(n9450) );
  AND2_X1 U5798 ( .A1(n4647), .A2(n4646), .ZN(n4645) );
  NAND2_X1 U5799 ( .A1(n9517), .A2(n4647), .ZN(n9468) );
  AND2_X1 U5800 ( .A1(n9536), .A2(n9703), .ZN(n9517) );
  NAND2_X1 U5801 ( .A1(n9517), .A2(n9699), .ZN(n9499) );
  NAND2_X1 U5802 ( .A1(n9547), .A2(n9548), .ZN(n9546) );
  OR2_X1 U5803 ( .A1(n5459), .A2(n8795), .ZN(n5477) );
  NAND2_X1 U5804 ( .A1(n4760), .A2(n4759), .ZN(n7870) );
  AOI21_X1 U5805 ( .B1(n4761), .B2(n4763), .A(n4570), .ZN(n4759) );
  NAND2_X1 U5806 ( .A1(n7705), .A2(n9103), .ZN(n7704) );
  NAND2_X1 U5807 ( .A1(n4755), .A2(n4754), .ZN(n7613) );
  AOI21_X1 U5808 ( .B1(n4756), .B2(n4758), .A(n4571), .ZN(n4754) );
  NAND2_X1 U5809 ( .A1(n5379), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n5419) );
  AND2_X1 U5810 ( .A1(n5361), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n5379) );
  NAND2_X1 U5811 ( .A1(n4751), .A2(n9166), .ZN(n7482) );
  INV_X1 U5812 ( .A(n7660), .ZN(n4641) );
  NAND2_X1 U5813 ( .A1(n7364), .A2(n4642), .ZN(n7504) );
  NAND2_X1 U5814 ( .A1(n7364), .A2(n9898), .ZN(n7474) );
  AND2_X1 U5815 ( .A1(n7243), .A2(n7353), .ZN(n7364) );
  NOR2_X1 U5816 ( .A1(n7218), .A2(n7219), .ZN(n7243) );
  NAND2_X1 U5817 ( .A1(n5263), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n5302) );
  AND2_X1 U5818 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n5263) );
  NOR2_X1 U5819 ( .A1(n4775), .A2(n7149), .ZN(n4774) );
  INV_X1 U5820 ( .A(n5238), .ZN(n4775) );
  NAND2_X1 U5821 ( .A1(n8966), .A2(n9152), .ZN(n9105) );
  NAND2_X1 U5822 ( .A1(n4739), .A2(n9549), .ZN(n4738) );
  OAI21_X1 U5823 ( .B1(n7489), .B2(n4758), .A(n4756), .ZN(n7629) );
  NAND2_X1 U5824 ( .A1(n7488), .A2(n5387), .ZN(n7630) );
  INV_X1 U5825 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n5163) );
  INV_X1 U5826 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n4795) );
  INV_X1 U5827 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5178) );
  XNOR2_X1 U5828 ( .A(n5710), .B(n5709), .ZN(n8162) );
  NAND2_X1 U5829 ( .A1(n5698), .A2(n5697), .ZN(n5710) );
  XNOR2_X1 U5830 ( .A(n5696), .B(n5695), .ZN(n8781) );
  INV_X1 U5831 ( .A(n4914), .ZN(n4912) );
  NAND2_X1 U5832 ( .A1(n5752), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5754) );
  OAI21_X1 U5833 ( .B1(n5574), .B2(n4971), .A(n4969), .ZN(n5603) );
  XNOR2_X1 U5834 ( .A(n5393), .B(n5388), .ZN(n6705) );
  NAND2_X1 U5835 ( .A1(n5370), .A2(n5369), .ZN(n5393) );
  NAND2_X1 U5836 ( .A1(n4720), .A2(n4719), .ZN(n5354) );
  INV_X1 U5837 ( .A(n5352), .ZN(n4719) );
  INV_X1 U5838 ( .A(n5353), .ZN(n4720) );
  NAND2_X1 U5839 ( .A1(n4962), .A2(n4963), .ZN(n5330) );
  NAND2_X1 U5840 ( .A1(n5314), .A2(n5313), .ZN(n5322) );
  NOR2_X1 U5841 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), .ZN(
        n5148) );
  NAND2_X1 U5842 ( .A1(n4715), .A2(n5274), .ZN(n5293) );
  NAND2_X1 U5843 ( .A1(n5271), .A2(n5270), .ZN(n4715) );
  NAND2_X1 U5844 ( .A1(n7936), .A2(n4565), .ZN(n5010) );
  AND3_X1 U5845 ( .A1(n5042), .A2(n4661), .A3(n5040), .ZN(n7088) );
  NAND2_X1 U5846 ( .A1(n7085), .A2(n5041), .ZN(n5040) );
  NOR2_X1 U5847 ( .A1(n5140), .A2(n5145), .ZN(n4661) );
  INV_X1 U5848 ( .A(n8702), .ZN(n8211) );
  NAND2_X1 U5849 ( .A1(n7623), .A2(n7622), .ZN(n7716) );
  NAND2_X1 U5850 ( .A1(n7001), .A2(n7000), .ZN(n7003) );
  INV_X1 U5851 ( .A(n8580), .ZN(n8554) );
  NAND2_X1 U5852 ( .A1(n7459), .A2(n7458), .ZN(n7572) );
  OR2_X1 U5853 ( .A1(n8250), .A2(n8239), .ZN(n4690) );
  OAI21_X1 U5854 ( .B1(n7623), .B2(n5073), .A(n5071), .ZN(n7911) );
  AOI21_X1 U5855 ( .B1(n5072), .B2(n5076), .A(n4529), .ZN(n5071) );
  NAND2_X1 U5856 ( .A1(n7912), .A2(n4663), .ZN(n7913) );
  OAI21_X1 U5857 ( .B1(n7911), .B2(n7910), .A(n8608), .ZN(n4663) );
  NAND2_X1 U5858 ( .A1(n7013), .A2(n7012), .ZN(n7015) );
  OR2_X1 U5859 ( .A1(n8221), .A2(n4697), .ZN(n4696) );
  OR2_X1 U5860 ( .A1(n5069), .A2(n5068), .ZN(n5065) );
  NAND2_X1 U5861 ( .A1(n8230), .A2(n4658), .ZN(n8270) );
  NOR2_X1 U5862 ( .A1(n8268), .A2(n4659), .ZN(n4658) );
  INV_X1 U5863 ( .A(n8178), .ZN(n4659) );
  NAND2_X1 U5864 ( .A1(n8230), .A2(n8178), .ZN(n8269) );
  NAND2_X1 U5865 ( .A1(n7439), .A2(n7457), .ZN(n7459) );
  NAND2_X1 U5866 ( .A1(n4672), .A2(n7438), .ZN(n7439) );
  NAND2_X1 U5867 ( .A1(n7437), .A2(n7436), .ZN(n4672) );
  INV_X1 U5868 ( .A(n7954), .ZN(n6968) );
  XNOR2_X1 U5869 ( .A(n7084), .B(n8315), .ZN(n7177) );
  NAND2_X1 U5870 ( .A1(n8250), .A2(n4684), .ZN(n4677) );
  OR2_X1 U5871 ( .A1(n8250), .A2(n4683), .ZN(n4678) );
  NAND2_X1 U5872 ( .A1(n5074), .A2(n7714), .ZN(n7718) );
  NAND2_X1 U5873 ( .A1(n5074), .A2(n5072), .ZN(n7838) );
  INV_X1 U5874 ( .A(n7123), .ZN(n6267) );
  OR2_X1 U5875 ( .A1(n6543), .A2(n6227), .ZN(n6233) );
  NAND2_X1 U5876 ( .A1(n4796), .A2(n4801), .ZN(n6786) );
  NAND2_X1 U5877 ( .A1(n4798), .A2(n4801), .ZN(n6764) );
  INV_X1 U5878 ( .A(n4805), .ZN(n10009) );
  OR2_X1 U5879 ( .A1(n7776), .A2(n7825), .ZN(n4809) );
  NAND2_X1 U5880 ( .A1(n4807), .A2(n4806), .ZN(n8346) );
  XNOR2_X1 U5881 ( .A(n8370), .B(n8371), .ZN(n8348) );
  INV_X1 U5882 ( .A(n9939), .ZN(n10084) );
  INV_X1 U5883 ( .A(n4813), .ZN(n8421) );
  OR2_X1 U5884 ( .A1(n6876), .A2(n6653), .ZN(n8428) );
  NAND2_X1 U5885 ( .A1(n8483), .A2(n6577), .ZN(n8094) );
  NAND2_X1 U5886 ( .A1(n8480), .A2(n8479), .ZN(n8481) );
  NAND2_X1 U5887 ( .A1(n8502), .A2(n8618), .ZN(n8479) );
  AOI21_X1 U5888 ( .B1(n8552), .B2(n8110), .A(n4519), .ZN(n8540) );
  NAND2_X1 U5889 ( .A1(n6462), .A2(n6461), .ZN(n8666) );
  NAND2_X1 U5890 ( .A1(n6452), .A2(n6451), .ZN(n8671) );
  NAND2_X1 U5891 ( .A1(n6367), .A2(n6366), .ZN(n8686) );
  NAND2_X1 U5892 ( .A1(n4867), .A2(n7983), .ZN(n7517) );
  NAND2_X1 U5893 ( .A1(n6566), .A2(n4868), .ZN(n4867) );
  NAND2_X1 U5894 ( .A1(n6566), .A2(n7986), .ZN(n7447) );
  NAND2_X1 U5895 ( .A1(n7287), .A2(n7975), .ZN(n7313) );
  AOI21_X1 U5896 ( .B1(n7810), .B2(n6655), .A(n4698), .ZN(n6292) );
  AND2_X1 U5897 ( .A1(n6460), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n4698) );
  OR2_X1 U5898 ( .A1(n6905), .A2(n6904), .ZN(n10097) );
  INV_X1 U5899 ( .A(n8610), .ZN(n10105) );
  NAND2_X1 U5900 ( .A1(n6861), .A2(n4857), .ZN(n6865) );
  AND2_X1 U5901 ( .A1(n7529), .A2(n7688), .ZN(n10147) );
  INV_X1 U5902 ( .A(n10105), .ZN(n10103) );
  NAND2_X1 U5903 ( .A1(n7941), .A2(n7940), .ZN(n8691) );
  NAND2_X1 U5904 ( .A1(n8077), .A2(n8076), .ZN(n8695) );
  XOR2_X1 U5905 ( .A(n8499), .B(n8501), .Z(n8711) );
  NAND2_X1 U5906 ( .A1(n8784), .A2(n6203), .ZN(n6509) );
  OAI21_X1 U5907 ( .B1(n8653), .B2(n4884), .A(n4881), .ZN(n8515) );
  NAND2_X1 U5908 ( .A1(n6206), .A2(n6205), .ZN(n8719) );
  INV_X1 U5909 ( .A(n5120), .ZN(n5113) );
  NAND2_X1 U5910 ( .A1(n4887), .A2(n8051), .ZN(n8519) );
  NAND2_X1 U5911 ( .A1(n8653), .A2(n4888), .ZN(n4887) );
  NAND2_X1 U5912 ( .A1(n5116), .A2(n5117), .ZN(n8532) );
  NAND2_X1 U5913 ( .A1(n8653), .A2(n8047), .ZN(n8530) );
  NAND2_X1 U5914 ( .A1(n6469), .A2(n6468), .ZN(n8736) );
  NAND2_X1 U5915 ( .A1(n6437), .A2(n6436), .ZN(n8750) );
  NAND2_X1 U5916 ( .A1(n6425), .A2(n6424), .ZN(n8757) );
  NAND2_X1 U5917 ( .A1(n6401), .A2(n6400), .ZN(n7887) );
  AND2_X1 U5918 ( .A1(n7739), .A2(n7738), .ZN(n7756) );
  NAND2_X1 U5919 ( .A1(n4901), .A2(n8001), .ZN(n7735) );
  NAND2_X1 U5920 ( .A1(n6379), .A2(n6378), .ZN(n8000) );
  XNOR2_X1 U5921 ( .A(n6596), .B(n6595), .ZN(n8786) );
  NAND2_X1 U5922 ( .A1(n6600), .A2(n6599), .ZN(n8166) );
  INV_X1 U5923 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n10268) );
  INV_X1 U5924 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n10368) );
  INV_X1 U5925 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6704) );
  INV_X1 U5926 ( .A(n7787), .ZN(n9989) );
  OR2_X1 U5927 ( .A1(n6291), .A2(n6290), .ZN(n9976) );
  INV_X1 U5928 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6661) );
  INV_X1 U5929 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6660) );
  MUX2_X1 U5930 ( .A(n6246), .B(n6245), .S(P2_IR_REG_3__SCAN_IN), .Z(n6247) );
  INV_X1 U5931 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6659) );
  INV_X1 U5932 ( .A(n4816), .ZN(n4815) );
  OAI21_X1 U5933 ( .B1(n6213), .B2(n4819), .A(n4817), .ZN(n4816) );
  NAND2_X1 U5934 ( .A1(n4827), .A2(n7189), .ZN(n7339) );
  NAND2_X1 U5935 ( .A1(n5629), .A2(n5628), .ZN(n9435) );
  NAND2_X1 U5936 ( .A1(n5912), .A2(n4854), .ZN(n7595) );
  OR2_X1 U5937 ( .A1(n8816), .A2(n4846), .ZN(n4843) );
  INV_X1 U5938 ( .A(n4853), .ZN(n8846) );
  NAND2_X1 U5939 ( .A1(n5662), .A2(n5661), .ZN(n9404) );
  NAND2_X1 U5940 ( .A1(n8784), .A2(n5295), .ZN(n5662) );
  NAND2_X1 U5941 ( .A1(n5515), .A2(n5514), .ZN(n9537) );
  NAND2_X1 U5942 ( .A1(n4847), .A2(n6008), .ZN(n8889) );
  OR2_X1 U5943 ( .A1(n8816), .A2(n6009), .ZN(n4847) );
  NAND2_X1 U5944 ( .A1(n8836), .A2(n8835), .ZN(n4837) );
  NAND2_X1 U5945 ( .A1(n5534), .A2(n5533), .ZN(n9519) );
  INV_X1 U5946 ( .A(n8942), .ZN(n9758) );
  INV_X1 U5947 ( .A(n9766), .ZN(n8958) );
  OR2_X1 U5948 ( .A1(n5687), .A2(n7108), .ZN(n5205) );
  AND2_X1 U5949 ( .A1(n5793), .A2(n9339), .ZN(n9351) );
  AND2_X1 U5950 ( .A1(n6114), .A2(n6113), .ZN(n9356) );
  NAND2_X1 U5951 ( .A1(n4782), .A2(n4780), .ZN(n6114) );
  NAND2_X1 U5952 ( .A1(n4782), .A2(n5708), .ZN(n6112) );
  NAND2_X1 U5953 ( .A1(n4768), .A2(n4769), .ZN(n9411) );
  NAND2_X1 U5954 ( .A1(n9449), .A2(n4772), .ZN(n4768) );
  OAI21_X1 U5955 ( .B1(n9449), .B2(n5615), .A(n5614), .ZN(n9426) );
  NAND2_X1 U5956 ( .A1(n4790), .A2(n5583), .ZN(n9459) );
  NAND2_X1 U5957 ( .A1(n4793), .A2(n4791), .ZN(n4790) );
  NAND2_X1 U5958 ( .A1(n4793), .A2(n5572), .ZN(n9483) );
  NAND2_X1 U5959 ( .A1(n4743), .A2(n4744), .ZN(n7698) );
  NAND2_X1 U5960 ( .A1(n5437), .A2(n5436), .ZN(n8901) );
  NAND2_X1 U5961 ( .A1(n5767), .A2(n8990), .ZN(n7240) );
  NAND2_X1 U5962 ( .A1(n4776), .A2(n5238), .ZN(n7151) );
  OR2_X1 U5963 ( .A1(n9857), .A2(n7103), .ZN(n9873) );
  INV_X1 U5964 ( .A(n9859), .ZN(n9877) );
  MUX2_X1 U5965 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n8961), .S(n5431), .Z(n8963) );
  AND2_X1 U5966 ( .A1(n9590), .A2(n9589), .ZN(n9666) );
  XNOR2_X1 U5967 ( .A(n5724), .B(n5723), .ZN(n9728) );
  INV_X1 U5968 ( .A(n9236), .ZN(n9099) );
  INV_X1 U5969 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6669) );
  INV_X1 U5970 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6666) );
  NAND2_X1 U5971 ( .A1(n5057), .A2(n8205), .ZN(n5056) );
  NAND2_X1 U5972 ( .A1(n4617), .A2(n4616), .ZN(n8158) );
  AOI211_X1 U5973 ( .C1(n8466), .C2(n10058), .A(n8465), .B(n8464), .ZN(n8467)
         );
  AOI21_X1 U5974 ( .B1(n8418), .B2(n4812), .A(n4810), .ZN(n8445) );
  OR2_X1 U5975 ( .A1(n8705), .A2(n8630), .ZN(n4630) );
  NAND2_X1 U5976 ( .A1(n6632), .A2(n8678), .ZN(n6634) );
  AND2_X1 U5977 ( .A1(n6658), .A2(n6700), .ZN(P1_U3973) );
  OAI21_X1 U5978 ( .B1(n4654), .B2(n9766), .A(n6137), .ZN(n6138) );
  AND2_X1 U5979 ( .A1(n6087), .A2(n8942), .ZN(n6109) );
  NAND2_X1 U5980 ( .A1(n4611), .A2(n4556), .ZN(n8950) );
  OAI21_X1 U5981 ( .B1(n9100), .B2(n4626), .A(n4624), .ZN(n9240) );
  OAI21_X1 U5982 ( .B1(n9666), .B2(n9916), .A(n4651), .ZN(P1_U3552) );
  INV_X1 U5983 ( .A(n4652), .ZN(n4651) );
  OAI22_X1 U5984 ( .A1(n4948), .A2(n9652), .B1(n9918), .B2(n5759), .ZN(n4652)
         );
  AOI21_X1 U5985 ( .B1(n9349), .B2(n6638), .A(n6637), .ZN(n6639) );
  NOR2_X1 U5986 ( .A1(n9918), .A2(n6636), .ZN(n6637) );
  NAND2_X2 U5987 ( .A1(n8962), .A2(n7936), .ZN(n5234) );
  NAND2_X1 U5988 ( .A1(n6065), .A2(n6064), .ZN(n4518) );
  NOR2_X1 U5989 ( .A1(n8175), .A2(n6486), .ZN(n4519) );
  OR2_X1 U5990 ( .A1(n5409), .A2(n4998), .ZN(n4520) );
  XNOR2_X1 U5991 ( .A(n6553), .B(P2_IR_REG_21__SCAN_IN), .ZN(n6888) );
  AND2_X1 U5992 ( .A1(n6557), .A2(n6556), .ZN(n8145) );
  NAND2_X1 U5993 ( .A1(n4632), .A2(n4631), .ZN(n4521) );
  INV_X1 U5994 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n6157) );
  AND2_X1 U5995 ( .A1(n8896), .A2(n4838), .ZN(n4522) );
  AND2_X1 U5996 ( .A1(n4844), .A2(n4842), .ZN(n4523) );
  AND2_X1 U5997 ( .A1(n8066), .A2(n8484), .ZN(n4524) );
  AND2_X1 U5998 ( .A1(n6008), .A2(n6009), .ZN(n4525) );
  AND2_X1 U5999 ( .A1(n9038), .A2(n8983), .ZN(n4526) );
  AND2_X1 U6000 ( .A1(n5117), .A2(n4561), .ZN(n4527) );
  INV_X1 U6001 ( .A(n7448), .ZN(n4860) );
  AND2_X1 U6002 ( .A1(n4520), .A2(n5427), .ZN(n4528) );
  AND2_X1 U6003 ( .A1(n7837), .A2(n8619), .ZN(n4529) );
  NAND2_X1 U6004 ( .A1(n9517), .A2(n4649), .ZN(n4650) );
  AND2_X1 U6005 ( .A1(n5058), .A2(n4573), .ZN(n4530) );
  NAND3_X1 U6006 ( .A1(n6595), .A2(n6597), .A3(n6617), .ZN(n4531) );
  INV_X1 U6007 ( .A(n5131), .ZN(n5128) );
  NAND2_X1 U6008 ( .A1(n8211), .A2(n8200), .ZN(n5131) );
  NOR2_X1 U6009 ( .A1(n7998), .A2(n8087), .ZN(n4532) );
  AND2_X1 U6010 ( .A1(n4856), .A2(n4855), .ZN(n4533) );
  OR3_X1 U6011 ( .A1(n9579), .A2(n9025), .A3(n9655), .ZN(n4534) );
  OR2_X1 U6012 ( .A1(n5453), .A2(P1_IR_REG_14__SCAN_IN), .ZN(n4535) );
  AND2_X1 U6013 ( .A1(n4737), .A2(n4609), .ZN(n4536) );
  NAND2_X1 U6014 ( .A1(n5494), .A2(n5493), .ZN(n9555) );
  INV_X1 U6015 ( .A(n9555), .ZN(n4639) );
  NAND2_X1 U6016 ( .A1(n6984), .A2(n8111), .ZN(n6985) );
  INV_X2 U6017 ( .A(n6263), .ZN(n6203) );
  INV_X2 U6018 ( .A(n5264), .ZN(n5244) );
  NOR2_X1 U6019 ( .A1(n8548), .A2(n5119), .ZN(n5118) );
  NAND2_X2 U6020 ( .A1(n6189), .A2(n6190), .ZN(n6229) );
  INV_X1 U6021 ( .A(n4515), .ZN(n6079) );
  OR2_X1 U6022 ( .A1(n8321), .A2(n8320), .ZN(n4537) );
  NAND2_X1 U6023 ( .A1(n8184), .A2(n8183), .ZN(n5083) );
  INV_X1 U6024 ( .A(n7457), .ZN(n5067) );
  NAND2_X1 U6025 ( .A1(n8171), .A2(n8597), .ZN(n4538) );
  NAND2_X1 U6026 ( .A1(n6689), .A2(n6916), .ZN(n5052) );
  INV_X1 U6027 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n5276) );
  AND3_X1 U6028 ( .A1(n6449), .A2(n6448), .A3(n6447), .ZN(n4539) );
  AND2_X1 U6029 ( .A1(n7394), .A2(n7985), .ZN(n8120) );
  NOR2_X1 U6030 ( .A1(n9209), .A2(n9213), .ZN(n4540) );
  NAND4_X2 U6031 ( .A1(n5205), .A2(n5204), .A3(n5203), .A4(n5202), .ZN(n5852)
         );
  XOR2_X1 U6032 ( .A(n5207), .B(n5208), .Z(n4541) );
  NAND2_X1 U6033 ( .A1(n4843), .A2(n4844), .ZN(n8827) );
  AND2_X1 U6034 ( .A1(n8257), .A2(n8222), .ZN(n4542) );
  OR2_X1 U6035 ( .A1(n9470), .A2(n9246), .ZN(n4543) );
  NOR2_X1 U6036 ( .A1(n9665), .A2(n9335), .ZN(n9218) );
  INV_X1 U6037 ( .A(n9218), .ZN(n4949) );
  NAND2_X1 U6038 ( .A1(n9094), .A2(n9093), .ZN(n9343) );
  INV_X1 U6039 ( .A(n9343), .ZN(n4948) );
  AND2_X1 U6040 ( .A1(n4690), .A2(n8238), .ZN(n4544) );
  AND2_X1 U6041 ( .A1(n9435), .A2(n9244), .ZN(n4545) );
  OR2_X1 U6042 ( .A1(n10146), .A2(n8311), .ZN(n4546) );
  INV_X1 U6043 ( .A(n7974), .ZN(n4872) );
  NAND2_X1 U6044 ( .A1(n5562), .A2(n5561), .ZN(n9502) );
  AND2_X1 U6045 ( .A1(n8887), .A2(n6014), .ZN(n4547) );
  NAND2_X1 U6046 ( .A1(n5649), .A2(n5648), .ZN(n9420) );
  OR2_X1 U6047 ( .A1(n8702), .A2(n8200), .ZN(n8066) );
  OR2_X1 U6048 ( .A1(n8204), .A2(n8203), .ZN(n4548) );
  NOR2_X1 U6049 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n5212) );
  AND2_X1 U6050 ( .A1(n7979), .A2(n8090), .ZN(n4549) );
  OR2_X1 U6051 ( .A1(n8671), .A2(n8607), .ZN(n4550) );
  XOR2_X1 U6052 ( .A(n9339), .B(n9343), .Z(n4551) );
  AND2_X1 U6053 ( .A1(n5161), .A2(n4795), .ZN(n4552) );
  AND2_X1 U6054 ( .A1(n6892), .A2(n7209), .ZN(n4553) );
  OR2_X1 U6055 ( .A1(n7927), .A2(n10141), .ZN(n4554) );
  OR2_X1 U6056 ( .A1(n5554), .A2(n5553), .ZN(n5574) );
  INV_X1 U6057 ( .A(n8113), .ZN(n4612) );
  AND2_X1 U6058 ( .A1(n8190), .A2(n8298), .ZN(n4555) );
  AND2_X1 U6059 ( .A1(n8943), .A2(n8942), .ZN(n4556) );
  AND2_X1 U6060 ( .A1(n6021), .A2(n6020), .ZN(n4557) );
  INV_X1 U6061 ( .A(n9470), .ZN(n5791) );
  NAND2_X1 U6062 ( .A1(n5590), .A2(n5589), .ZN(n9470) );
  AND2_X1 U6063 ( .A1(n4642), .A2(n4641), .ZN(n4558) );
  AND2_X1 U6064 ( .A1(n5096), .A2(n5097), .ZN(n4559) );
  AND2_X1 U6065 ( .A1(n5011), .A2(n4899), .ZN(n4560) );
  OR2_X1 U6066 ( .A1(n8725), .A2(n8541), .ZN(n4561) );
  NAND2_X1 U6067 ( .A1(n9433), .A2(n4656), .ZN(n4657) );
  AND2_X1 U6068 ( .A1(n9040), .A2(n9041), .ZN(n4562) );
  INV_X1 U6069 ( .A(n4987), .ZN(n4986) );
  NAND2_X1 U6070 ( .A1(n5488), .A2(n4563), .ZN(n4987) );
  OR2_X1 U6071 ( .A1(n5505), .A2(SI_16_), .ZN(n4563) );
  NAND2_X1 U6072 ( .A1(n9420), .A2(n8847), .ZN(n4564) );
  AND2_X1 U6073 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n4565) );
  INV_X1 U6074 ( .A(n5076), .ZN(n5075) );
  OR2_X1 U6075 ( .A1(n7715), .A2(n5077), .ZN(n5076) );
  AND2_X1 U6076 ( .A1(n4546), .A2(n6348), .ZN(n4566) );
  INV_X1 U6077 ( .A(n7993), .ZN(n4862) );
  NAND2_X1 U6078 ( .A1(n8985), .A2(n4907), .ZN(n4567) );
  AND2_X1 U6079 ( .A1(n4813), .A2(n4812), .ZN(n4568) );
  BUF_X1 U6080 ( .A(n5832), .Z(n5840) );
  INV_X1 U6081 ( .A(n5832), .ZN(n4752) );
  AND2_X1 U6082 ( .A1(n5956), .A2(n5955), .ZN(n4569) );
  NOR2_X1 U6083 ( .A1(n9655), .A2(n9253), .ZN(n4570) );
  NOR2_X1 U6084 ( .A1(n4622), .A2(n9256), .ZN(n4571) );
  NOR2_X1 U6085 ( .A1(n9420), .A2(n8847), .ZN(n4572) );
  OAI211_X1 U6086 ( .C1(n6587), .C2(n6744), .A(n4898), .B(n4897), .ZN(n6225)
         );
  NAND2_X1 U6087 ( .A1(n9202), .A2(n9200), .ZN(n9136) );
  INV_X1 U6088 ( .A(n9136), .ZN(n4740) );
  INV_X1 U6089 ( .A(n4946), .ZN(n4945) );
  NAND2_X1 U6090 ( .A1(n4950), .A2(n4947), .ZN(n4946) );
  OR2_X1 U6091 ( .A1(n8197), .A2(n8195), .ZN(n4573) );
  AND2_X1 U6092 ( .A1(n5505), .A2(SI_16_), .ZN(n4574) );
  AND2_X1 U6093 ( .A1(n5294), .A2(SI_5_), .ZN(n4575) );
  AND2_X1 U6094 ( .A1(n5323), .A2(SI_7_), .ZN(n4576) );
  AND2_X1 U6095 ( .A1(n4740), .A2(n4948), .ZN(n4577) );
  NAND2_X1 U6096 ( .A1(n8036), .A2(n8033), .ZN(n4578) );
  NAND2_X1 U6097 ( .A1(n4913), .A2(n4911), .ZN(n4579) );
  NAND2_X1 U6098 ( .A1(n6152), .A2(n6151), .ZN(n4580) );
  NOR2_X1 U6099 ( .A1(n8547), .A2(n8533), .ZN(n4581) );
  AND2_X1 U6100 ( .A1(n4541), .A2(n7936), .ZN(n4582) );
  OR2_X1 U6101 ( .A1(n8106), .A2(n8065), .ZN(n4583) );
  INV_X1 U6102 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n6153) );
  INV_X1 U6103 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n6154) );
  NAND2_X1 U6104 ( .A1(n6498), .A2(n6497), .ZN(n8725) );
  OR2_X1 U6105 ( .A1(n6224), .A2(n4509), .ZN(n7946) );
  INV_X1 U6106 ( .A(n5073), .ZN(n5072) );
  NAND2_X1 U6107 ( .A1(n5078), .A2(n7714), .ZN(n5073) );
  AND2_X1 U6108 ( .A1(n6015), .A2(n8886), .ZN(n4584) );
  AND2_X1 U6109 ( .A1(n5429), .A2(SI_12_), .ZN(n4585) );
  INV_X1 U6110 ( .A(n4767), .ZN(n4766) );
  NAND2_X1 U6111 ( .A1(n4769), .A2(n4564), .ZN(n4767) );
  AND2_X1 U6112 ( .A1(n5083), .A2(n8272), .ZN(n4586) );
  OR2_X1 U6113 ( .A1(n7188), .A2(n4831), .ZN(n4587) );
  INV_X1 U6114 ( .A(n8051), .ZN(n4886) );
  INV_X1 U6115 ( .A(n5127), .ZN(n5125) );
  NOR2_X1 U6116 ( .A1(n5128), .A2(n6527), .ZN(n5127) );
  INV_X1 U6117 ( .A(n8708), .ZN(n8304) );
  NAND2_X1 U6118 ( .A1(n6518), .A2(n6517), .ZN(n8708) );
  NAND2_X1 U6119 ( .A1(n8719), .A2(n8534), .ZN(n4588) );
  OR2_X1 U6120 ( .A1(n5132), .A2(n5129), .ZN(n4589) );
  OR2_X1 U6121 ( .A1(n5115), .A2(n5113), .ZN(n4590) );
  AND3_X1 U6122 ( .A1(n7980), .A2(n7981), .A3(n8120), .ZN(n4591) );
  NOR2_X1 U6123 ( .A1(n6387), .A2(n5107), .ZN(n4592) );
  AND2_X1 U6124 ( .A1(n8057), .A2(n8514), .ZN(n4593) );
  AND2_X1 U6125 ( .A1(n4996), .A2(n5427), .ZN(n4594) );
  INV_X1 U6126 ( .A(n4685), .ZN(n4684) );
  NAND2_X1 U6127 ( .A1(n8238), .A2(n8192), .ZN(n4685) );
  NAND2_X1 U6128 ( .A1(n7997), .A2(n7993), .ZN(n4595) );
  AND2_X1 U6129 ( .A1(n4941), .A2(n4949), .ZN(n4596) );
  NAND2_X1 U6130 ( .A1(n7996), .A2(n7995), .ZN(n4597) );
  INV_X1 U6131 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n4818) );
  INV_X1 U6132 ( .A(n9392), .ZN(n9674) );
  NAND2_X1 U6133 ( .A1(n5683), .A2(n5682), .ZN(n9392) );
  AND2_X1 U6134 ( .A1(n5090), .A2(n4566), .ZN(n4598) );
  INV_X1 U6135 ( .A(n5320), .ZN(n5321) );
  XNOR2_X1 U6136 ( .A(n5323), .B(SI_7_), .ZN(n5320) );
  NAND2_X1 U6137 ( .A1(n5704), .A2(n5703), .ZN(n9375) );
  INV_X1 U6138 ( .A(n9375), .ZN(n4654) );
  INV_X1 U6139 ( .A(n10017), .ZN(n4802) );
  NAND2_X1 U6140 ( .A1(n4959), .A2(n6539), .ZN(n6632) );
  AND2_X1 U6141 ( .A1(n8012), .A2(n8013), .ZN(n8011) );
  INV_X1 U6142 ( .A(n8011), .ZN(n5022) );
  INV_X1 U6143 ( .A(n8203), .ZN(n5064) );
  AND4_X1 U6144 ( .A1(n6362), .A2(n6361), .A3(n6360), .A4(n6359), .ZN(n7426)
         );
  INV_X1 U6145 ( .A(n9103), .ZN(n4742) );
  OR2_X1 U6146 ( .A1(n5602), .A2(SI_21_), .ZN(n4599) );
  NAND2_X1 U6147 ( .A1(n7704), .A2(n5446), .ZN(n9565) );
  NAND2_X1 U6148 ( .A1(n4521), .A2(n5091), .ZN(n7518) );
  INV_X1 U6149 ( .A(n6129), .ZN(n4610) );
  NAND2_X1 U6150 ( .A1(n6375), .A2(n6374), .ZN(n7673) );
  NAND2_X1 U6151 ( .A1(n4837), .A2(n5949), .ZN(n8895) );
  INV_X1 U6152 ( .A(n8568), .ZN(n5102) );
  AND2_X1 U6153 ( .A1(n6506), .A2(n6505), .ZN(n8272) );
  INV_X1 U6154 ( .A(n8272), .ZN(n8541) );
  NAND2_X1 U6155 ( .A1(n5928), .A2(n5932), .ZN(n9756) );
  AND3_X1 U6156 ( .A1(n5048), .A2(n5047), .A3(n6248), .ZN(n6307) );
  NOR3_X1 U6157 ( .A1(n9579), .A2(n9025), .A3(n4637), .ZN(n4640) );
  NAND2_X1 U6158 ( .A1(n4913), .A2(n4914), .ZN(n5512) );
  AND2_X1 U6159 ( .A1(n6119), .A2(n5722), .ZN(n4600) );
  AND2_X1 U6160 ( .A1(n5602), .A2(SI_21_), .ZN(n4601) );
  AND2_X1 U6161 ( .A1(n4696), .A2(n8222), .ZN(n4602) );
  OR2_X1 U6162 ( .A1(n6388), .A2(n5088), .ZN(n4603) );
  AND2_X1 U6163 ( .A1(n4809), .A2(n4537), .ZN(n4604) );
  NAND2_X1 U6164 ( .A1(n5609), .A2(n5608), .ZN(n9451) );
  INV_X1 U6165 ( .A(n9451), .ZN(n4646) );
  NAND2_X1 U6166 ( .A1(n5456), .A2(n5455), .ZN(n9655) );
  INV_X1 U6167 ( .A(n9655), .ZN(n4638) );
  NAND2_X1 U6168 ( .A1(n7013), .A2(n5043), .ZN(n7086) );
  NAND2_X1 U6169 ( .A1(n6254), .A2(n6253), .ZN(n7375) );
  NAND2_X1 U6170 ( .A1(n4832), .A2(n7141), .ZN(n7187) );
  NOR2_X1 U6171 ( .A1(n7176), .A2(n7177), .ZN(n4605) );
  NOR2_X1 U6172 ( .A1(n7385), .A2(n7413), .ZN(n4606) );
  NAND2_X1 U6173 ( .A1(n7364), .A2(n4558), .ZN(n4644) );
  OR2_X1 U6174 ( .A1(n6388), .A2(n5084), .ZN(n4607) );
  INV_X1 U6175 ( .A(n5007), .ZN(n5006) );
  OAI21_X1 U6176 ( .B1(n5697), .B2(n5008), .A(n5711), .ZN(n5007) );
  OR2_X1 U6177 ( .A1(n8350), .A2(n8333), .ZN(n4608) );
  INV_X1 U6178 ( .A(n9571), .ZN(n9549) );
  NAND2_X1 U6179 ( .A1(n5222), .A2(n5221), .ZN(n7276) );
  INV_X1 U6180 ( .A(n8112), .ZN(n4856) );
  OR2_X1 U6181 ( .A1(n9333), .A2(n9101), .ZN(n4609) );
  INV_X1 U6182 ( .A(n7188), .ZN(n4828) );
  NAND2_X1 U6183 ( .A1(n8918), .A2(n8919), .ZN(n8917) );
  NAND2_X1 U6184 ( .A1(n7048), .A2(n5872), .ZN(n5880) );
  NOR2_X2 U6185 ( .A1(n8905), .A2(n8907), .ZN(n8909) );
  OAI21_X2 U6186 ( .B1(n8941), .B2(n8940), .A(n8939), .ZN(n4611) );
  NAND2_X1 U6187 ( .A1(n4841), .A2(n4840), .ZN(n6028) );
  NAND2_X1 U6188 ( .A1(n5783), .A2(n9182), .ZN(n9479) );
  NAND2_X1 U6189 ( .A1(n4721), .A2(n5321), .ZN(n4962) );
  NAND2_X1 U6190 ( .A1(n4623), .A2(n4736), .ZN(n9445) );
  NAND3_X1 U6191 ( .A1(n5103), .A2(n6152), .A3(n6151), .ZN(n6602) );
  AND3_X2 U6192 ( .A1(n6307), .A2(n6234), .A3(n6143), .ZN(n6152) );
  NAND2_X1 U6193 ( .A1(n8009), .A2(n5018), .ZN(n5017) );
  NAND2_X1 U6194 ( .A1(n4722), .A2(n8038), .ZN(n5034) );
  NAND2_X1 U6195 ( .A1(n5032), .A2(n5030), .ZN(n8044) );
  AOI21_X1 U6196 ( .B1(n5028), .B2(n4593), .A(n4733), .ZN(n4732) );
  NOR2_X1 U6197 ( .A1(n7992), .A2(n4591), .ZN(n4730) );
  NAND2_X1 U6198 ( .A1(n4700), .A2(n4699), .ZN(n5029) );
  AOI21_X1 U6199 ( .B1(n8078), .B2(n5014), .A(n8087), .ZN(n4956) );
  NAND2_X1 U6200 ( .A1(n5403), .A2(n5402), .ZN(n8926) );
  INV_X1 U6201 ( .A(n9443), .ZN(n4623) );
  INV_X1 U6202 ( .A(n4748), .ZN(n4747) );
  NAND2_X1 U6203 ( .A1(n7633), .A2(n9006), .ZN(n4749) );
  NAND2_X2 U6204 ( .A1(n4743), .A2(n4619), .ZN(n9568) );
  XNOR2_X1 U6205 ( .A(n4741), .B(n4740), .ZN(n4739) );
  INV_X1 U6206 ( .A(n6602), .ZN(n4902) );
  NAND2_X1 U6207 ( .A1(n4896), .A2(n4524), .ZN(n8483) );
  NAND2_X2 U6208 ( .A1(n7395), .A2(n7984), .ZN(n6566) );
  NAND2_X2 U6209 ( .A1(n6587), .A2(n5011), .ZN(n8075) );
  NOR2_X2 U6210 ( .A1(n9991), .A2(n6312), .ZN(n9990) );
  NOR2_X1 U6211 ( .A1(n10025), .A2(n6341), .ZN(n10024) );
  NOR2_X1 U6212 ( .A1(n8372), .A2(n8373), .ZN(n8375) );
  NOR2_X1 U6213 ( .A1(n10042), .A2(n10041), .ZN(n10040) );
  OR2_X2 U6214 ( .A1(n5907), .A2(n5906), .ZN(n5912) );
  NOR2_X1 U6215 ( .A1(n6028), .A2(n6027), .ZN(n8905) );
  INV_X1 U6216 ( .A(n4913), .ZN(n5453) );
  AND2_X4 U6217 ( .A1(n5154), .A2(n5275), .ZN(n4913) );
  NAND2_X1 U6218 ( .A1(n4826), .A2(n4510), .ZN(n4823) );
  INV_X1 U6219 ( .A(n5207), .ZN(n4712) );
  NAND2_X1 U6220 ( .A1(n9400), .A2(n9399), .ZN(n9398) );
  NAND2_X1 U6221 ( .A1(n5785), .A2(n9186), .ZN(n9443) );
  NAND2_X1 U6222 ( .A1(n5795), .A2(n5794), .ZN(n5796) );
  INV_X1 U6223 ( .A(n5314), .ZN(n4721) );
  AOI21_X1 U6224 ( .B1(n6116), .B2(n9135), .A(n9197), .ZN(n4741) );
  NAND2_X1 U6225 ( .A1(n4990), .A2(n4988), .ZN(n5696) );
  NAND2_X1 U6226 ( .A1(n4712), .A2(n5208), .ZN(n5211) );
  NAND2_X1 U6227 ( .A1(n5449), .A2(n5448), .ZN(n5452) );
  OAI21_X1 U6228 ( .B1(n5618), .B2(n5617), .A(n5616), .ZN(n5626) );
  NAND2_X1 U6229 ( .A1(n5728), .A2(n5727), .ZN(n7929) );
  NAND2_X1 U6230 ( .A1(n4627), .A2(n8610), .ZN(n7925) );
  NAND2_X1 U6231 ( .A1(n6591), .A2(n6592), .ZN(n4627) );
  NOR2_X1 U6232 ( .A1(n10024), .A2(n7770), .ZN(n10042) );
  NAND2_X2 U6233 ( .A1(n9945), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n9964) );
  OAI21_X2 U6234 ( .B1(n8557), .B2(n6575), .A(n8048), .ZN(n8549) );
  NAND2_X2 U6235 ( .A1(n8549), .A2(n8548), .ZN(n8653) );
  NAND2_X1 U6236 ( .A1(n4878), .A2(n4875), .ZN(n8499) );
  OAI21_X2 U6237 ( .B1(n7878), .B2(n7877), .A(n8013), .ZN(n7900) );
  NAND2_X1 U6238 ( .A1(n6568), .A2(n6567), .ZN(n4901) );
  NAND2_X1 U6239 ( .A1(n6186), .A2(n6187), .ZN(n8767) );
  NOR2_X1 U6240 ( .A1(n8400), .A2(n10384), .ZN(n8418) );
  XNOR2_X1 U6241 ( .A(n6158), .B(n6157), .ZN(n6582) );
  NAND3_X1 U6242 ( .A1(n8498), .A2(n8497), .A3(n4630), .ZN(P2_U3206) );
  XNOR2_X2 U6243 ( .A(n6968), .B(n8318), .ZN(n8111) );
  NAND2_X1 U6244 ( .A1(n6375), .A2(n4592), .ZN(n5106) );
  NAND2_X1 U6245 ( .A1(n6270), .A2(n6269), .ZN(n7121) );
  INV_X1 U6246 ( .A(n4632), .ZN(n7316) );
  NOR2_X2 U6247 ( .A1(n7315), .A2(n8120), .ZN(n4632) );
  NAND2_X1 U6248 ( .A1(n5108), .A2(n8007), .ZN(n7879) );
  NAND2_X1 U6249 ( .A1(n6364), .A2(n6363), .ZN(n7665) );
  OR2_X1 U6250 ( .A1(n5842), .A2(n5841), .ZN(n5843) );
  NAND2_X2 U6251 ( .A1(n8163), .A2(n5757), .ZN(n8962) );
  OR2_X1 U6252 ( .A1(n5206), .A2(n4541), .ZN(n5187) );
  NOR2_X1 U6253 ( .A1(n9579), .A2(n9655), .ZN(n9577) );
  INV_X1 U6254 ( .A(n4640), .ZN(n9554) );
  INV_X1 U6255 ( .A(n4644), .ZN(n7503) );
  NAND3_X1 U6256 ( .A1(n4913), .A2(n4911), .A3(n5161), .ZN(n5803) );
  NAND3_X1 U6257 ( .A1(n4913), .A2(n4552), .A3(n4911), .ZN(n4753) );
  INV_X1 U6258 ( .A(n4650), .ZN(n9467) );
  NAND2_X1 U6259 ( .A1(n4551), .A2(n7872), .ZN(n9590) );
  INV_X1 U6260 ( .A(n4657), .ZN(n9403) );
  NAND2_X1 U6261 ( .A1(n7912), .A2(n4662), .ZN(n8167) );
  NAND3_X1 U6262 ( .A1(n4669), .A2(n5065), .A3(n4667), .ZN(n7621) );
  NAND2_X1 U6263 ( .A1(n7428), .A2(n4668), .ZN(n4667) );
  NAND2_X1 U6264 ( .A1(n7437), .A2(n4670), .ZN(n4669) );
  INV_X1 U6265 ( .A(n5066), .ZN(n4671) );
  NAND2_X1 U6266 ( .A1(n4902), .A2(n6154), .ZN(n6605) );
  NAND2_X1 U6267 ( .A1(n4902), .A2(n4673), .ZN(n4674) );
  NAND3_X1 U6268 ( .A1(n4676), .A2(n4675), .A3(n8293), .ZN(n8291) );
  NAND2_X1 U6269 ( .A1(n8250), .A2(n4679), .ZN(n4675) );
  NAND2_X1 U6270 ( .A1(n8250), .A2(n8238), .ZN(n4692) );
  NAND3_X1 U6271 ( .A1(n4678), .A2(n4677), .A3(n4681), .ZN(n8292) );
  NAND2_X1 U6272 ( .A1(n4692), .A2(n4691), .ZN(n8191) );
  INV_X1 U6273 ( .A(n4691), .ZN(n4687) );
  INV_X1 U6274 ( .A(n8192), .ZN(n4689) );
  NAND2_X1 U6275 ( .A1(n8221), .A2(n4542), .ZN(n4693) );
  NAND2_X1 U6276 ( .A1(n4693), .A2(n4694), .ZN(n8231) );
  INV_X1 U6277 ( .A(n4538), .ZN(n4697) );
  AOI21_X1 U6278 ( .B1(n8044), .B2(n4701), .A(n4702), .ZN(n4699) );
  NAND2_X1 U6279 ( .A1(n8046), .A2(n4704), .ZN(n4700) );
  AOI21_X1 U6280 ( .B1(n8044), .B2(n8043), .A(n8042), .ZN(n8050) );
  XNOR2_X1 U6281 ( .A(n5209), .B(SI_1_), .ZN(n5207) );
  NAND2_X1 U6282 ( .A1(n8029), .A2(n8087), .ZN(n4723) );
  NAND3_X1 U6283 ( .A1(n7987), .A2(n7986), .A3(n8087), .ZN(n4726) );
  NAND2_X1 U6284 ( .A1(n4727), .A2(n6567), .ZN(n8004) );
  NAND2_X1 U6285 ( .A1(n4729), .A2(n4728), .ZN(n4727) );
  OAI21_X1 U6286 ( .B1(n4730), .B2(n4595), .A(n5027), .ZN(n4728) );
  OAI21_X1 U6287 ( .B1(n4730), .B2(n4597), .A(n4532), .ZN(n4729) );
  AOI21_X2 U6288 ( .B1(n9445), .B2(n4735), .A(n4734), .ZN(n9413) );
  OR2_X2 U6289 ( .A1(n7632), .A2(n4748), .ZN(n4743) );
  OAI21_X1 U6290 ( .B1(n7632), .B2(n7633), .A(n9006), .ZN(n7603) );
  NAND2_X1 U6291 ( .A1(n5770), .A2(n4749), .ZN(n4748) );
  NAND2_X1 U6292 ( .A1(n5767), .A2(n4750), .ZN(n7357) );
  NAND2_X1 U6293 ( .A1(n7357), .A2(n9164), .ZN(n4751) );
  INV_X1 U6294 ( .A(n6958), .ZN(n9872) );
  OAI21_X2 U6295 ( .B1(n9383), .B2(n9384), .A(n9195), .ZN(n9368) );
  NAND2_X1 U6296 ( .A1(n7489), .A2(n4756), .ZN(n4755) );
  NAND2_X1 U6297 ( .A1(n7705), .A2(n4761), .ZN(n4760) );
  NAND2_X1 U6298 ( .A1(n7276), .A2(n9108), .ZN(n4776) );
  NAND2_X1 U6299 ( .A1(n4776), .A2(n4774), .ZN(n5262) );
  NAND2_X1 U6300 ( .A1(n5694), .A2(n4783), .ZN(n4782) );
  NAND2_X1 U6301 ( .A1(n5694), .A2(n5693), .ZN(n9366) );
  NAND3_X1 U6302 ( .A1(n4913), .A2(n4794), .A3(n4911), .ZN(n5175) );
  INV_X1 U6303 ( .A(n6763), .ZN(n4800) );
  INV_X1 U6304 ( .A(n4809), .ZN(n8322) );
  INV_X1 U6305 ( .A(n8419), .ZN(n4811) );
  INV_X1 U6306 ( .A(n8420), .ZN(n4812) );
  XNOR2_X2 U6307 ( .A(n4814), .B(n9989), .ZN(n9991) );
  NAND2_X2 U6308 ( .A1(n4820), .A2(n6657), .ZN(n5850) );
  AND2_X2 U6309 ( .A1(n5748), .A2(n5807), .ZN(n9236) );
  NAND3_X1 U6310 ( .A1(n4824), .A2(n4823), .A3(n4822), .ZN(n5903) );
  NAND2_X1 U6311 ( .A1(n7140), .A2(n4825), .ZN(n4824) );
  AND2_X1 U6312 ( .A1(n4829), .A2(n7142), .ZN(n4825) );
  NAND3_X1 U6313 ( .A1(n4832), .A2(n7141), .A3(n4828), .ZN(n4827) );
  INV_X1 U6314 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n4833) );
  NAND2_X1 U6315 ( .A1(n8836), .A2(n4522), .ZN(n4835) );
  NAND2_X1 U6316 ( .A1(n8816), .A2(n4523), .ZN(n4841) );
  NAND3_X1 U6317 ( .A1(n5928), .A2(n5932), .A3(n5931), .ZN(n9760) );
  NAND2_X1 U6318 ( .A1(n9760), .A2(n5932), .ZN(n8918) );
  NAND2_X1 U6319 ( .A1(n8880), .A2(n4852), .ZN(n4850) );
  NAND2_X1 U6320 ( .A1(n5907), .A2(n5906), .ZN(n4854) );
  INV_X1 U6321 ( .A(n6561), .ZN(n6562) );
  NOR2_X1 U6322 ( .A1(n6561), .A2(n7950), .ZN(n7951) );
  NAND2_X1 U6323 ( .A1(n6561), .A2(n5052), .ZN(n6867) );
  NOR2_X1 U6324 ( .A1(n6561), .A2(n8111), .ZN(n4855) );
  OR2_X1 U6325 ( .A1(n6561), .A2(n6862), .ZN(n4857) );
  NAND3_X1 U6326 ( .A1(n4859), .A2(n4858), .A3(n7666), .ZN(n7663) );
  NAND2_X1 U6327 ( .A1(n6566), .A2(n4861), .ZN(n4859) );
  OAI21_X1 U6328 ( .B1(n6566), .B2(n4864), .A(n4861), .ZN(n7664) );
  NAND2_X1 U6329 ( .A1(n7120), .A2(n4871), .ZN(n4870) );
  NAND2_X1 U6330 ( .A1(n8653), .A2(n4879), .ZN(n4878) );
  NAND2_X1 U6331 ( .A1(n8491), .A2(n8067), .ZN(n4896) );
  NAND2_X1 U6332 ( .A1(n4890), .A2(n4893), .ZN(n8099) );
  NAND2_X1 U6333 ( .A1(n8491), .A2(n4891), .ZN(n4890) );
  AND2_X1 U6334 ( .A1(n4896), .A2(n8066), .ZN(n8485) );
  INV_X1 U6335 ( .A(n4894), .ZN(n4893) );
  OAI21_X1 U6336 ( .B1(n4524), .B2(n4895), .A(n8093), .ZN(n4894) );
  INV_X1 U6337 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n4899) );
  NAND2_X1 U6338 ( .A1(n4901), .A2(n4900), .ZN(n6570) );
  AND2_X1 U6339 ( .A1(n5143), .A2(n8001), .ZN(n4900) );
  OR2_X2 U6340 ( .A1(n8588), .A2(n8591), .ZN(n8590) );
  NOR2_X2 U6341 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n6212) );
  NAND2_X1 U6342 ( .A1(n6605), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6158) );
  NAND2_X1 U6343 ( .A1(n8979), .A2(n9096), .ZN(n4908) );
  NAND2_X1 U6344 ( .A1(n8979), .A2(n4905), .ZN(n4904) );
  NAND2_X1 U6345 ( .A1(n9113), .A2(n8983), .ZN(n4909) );
  NOR2_X1 U6346 ( .A1(n9045), .A2(n9180), .ZN(n9044) );
  NOR2_X1 U6347 ( .A1(n4526), .A2(n4562), .ZN(n4910) );
  NOR2_X2 U6348 ( .A1(n5160), .A2(n4912), .ZN(n4911) );
  NAND2_X1 U6349 ( .A1(n9059), .A2(n4921), .ZN(n4916) );
  NAND2_X1 U6350 ( .A1(n4916), .A2(n4917), .ZN(n9077) );
  AOI21_X1 U6351 ( .B1(n9090), .B2(n4933), .A(n4931), .ZN(n9100) );
  OAI21_X1 U6352 ( .B1(n9089), .B2(n9343), .A(n4944), .ZN(n4943) );
  NAND2_X1 U6353 ( .A1(n9343), .A2(n8983), .ZN(n4944) );
  INV_X1 U6354 ( .A(n4955), .ZN(n4953) );
  NOR2_X1 U6355 ( .A1(n8081), .A2(n4956), .ZN(n4955) );
  INV_X1 U6356 ( .A(n5574), .ZN(n4965) );
  OAI21_X1 U6357 ( .B1(n4965), .B2(n4968), .A(n4966), .ZN(n5618) );
  NAND2_X1 U6358 ( .A1(n5490), .A2(n4977), .ZN(n4973) );
  NAND2_X1 U6359 ( .A1(n4973), .A2(n4974), .ZN(n5554) );
  NAND2_X1 U6360 ( .A1(n5645), .A2(n4991), .ZN(n4990) );
  NAND2_X1 U6361 ( .A1(n5370), .A2(n4594), .ZN(n4994) );
  NAND2_X1 U6362 ( .A1(n4994), .A2(n4995), .ZN(n5449) );
  INV_X1 U6363 ( .A(n5698), .ZN(n5003) );
  OAI21_X1 U6364 ( .B1(n5698), .B2(n5008), .A(n5006), .ZN(n5724) );
  OAI21_X1 U6365 ( .B1(n5003), .B2(n5007), .A(n5004), .ZN(n5728) );
  CLKBUF_X1 U6366 ( .A(n7936), .Z(n5009) );
  NAND2_X2 U6367 ( .A1(n5011), .A2(P2_U3151), .ZN(n8765) );
  NAND2_X1 U6368 ( .A1(n5197), .A2(n5010), .ZN(n5208) );
  NAND2_X1 U6369 ( .A1(n5011), .A2(n5183), .ZN(n5197) );
  MUX2_X1 U6370 ( .A(n6669), .B(n6660), .S(n7936), .Z(n5256) );
  MUX2_X1 U6371 ( .A(n6664), .B(n6661), .S(n7936), .Z(n5272) );
  MUX2_X1 U6372 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(P1_DATAO_REG_5__SCAN_IN), 
        .S(n7936), .Z(n5294) );
  MUX2_X1 U6373 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(P1_DATAO_REG_6__SCAN_IN), 
        .S(n7936), .Z(n5312) );
  MUX2_X1 U6374 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(P1_DATAO_REG_7__SCAN_IN), 
        .S(n7936), .Z(n5323) );
  MUX2_X1 U6375 ( .A(n5324), .B(n6688), .S(n7936), .Z(n5326) );
  MUX2_X1 U6376 ( .A(n5347), .B(n6704), .S(n7936), .Z(n5349) );
  MUX2_X1 U6377 ( .A(n5371), .B(n10368), .S(n5009), .Z(n5389) );
  MUX2_X1 U6378 ( .A(n5394), .B(n10268), .S(n5009), .Z(n5396) );
  MUX2_X1 U6379 ( .A(n10457), .B(n10382), .S(n5009), .Z(n5428) );
  MUX2_X1 U6380 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(P1_DATAO_REG_14__SCAN_IN), 
        .S(n5009), .Z(n5469) );
  MUX2_X1 U6381 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(P1_DATAO_REG_15__SCAN_IN), 
        .S(n5009), .Z(n5485) );
  MUX2_X1 U6382 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(P1_DATAO_REG_18__SCAN_IN), 
        .S(n5009), .Z(n5545) );
  MUX2_X1 U6383 ( .A(n7515), .B(n7512), .S(n5009), .Z(n5585) );
  MUX2_X1 U6384 ( .A(n7687), .B(n7690), .S(n5009), .Z(n5605) );
  MUX2_X1 U6385 ( .A(n5647), .B(n6204), .S(n5009), .Z(n5639) );
  MUX2_X1 U6386 ( .A(n9732), .B(n8782), .S(n5009), .Z(n5679) );
  MUX2_X1 U6387 ( .A(n9731), .B(n8777), .S(n5009), .Z(n5726) );
  OAI211_X1 U6388 ( .C1(n5022), .C2(n8010), .A(n5017), .B(n5015), .ZN(n8023)
         );
  NAND3_X1 U6389 ( .A1(n5046), .A2(n7085), .A3(n5045), .ZN(n5042) );
  NAND2_X1 U6390 ( .A1(n6893), .A2(n6894), .ZN(n6967) );
  NAND3_X1 U6391 ( .A1(n6891), .A2(n4509), .A3(n6892), .ZN(n5049) );
  NAND2_X1 U6392 ( .A1(n8204), .A2(n5055), .ZN(n5054) );
  OAI211_X1 U6393 ( .C1(n8204), .C2(n5056), .A(n5054), .B(n8202), .ZN(P2_U3160) );
  NAND2_X1 U6394 ( .A1(n8182), .A2(n5082), .ZN(n5081) );
  AND2_X1 U6395 ( .A1(n8248), .A2(n5083), .ZN(n8213) );
  AND3_X2 U6396 ( .A1(n6592), .A2(n6591), .A3(n4554), .ZN(n6652) );
  NOR2_X2 U6397 ( .A1(n6605), .A2(n5089), .ZN(n6186) );
  NAND2_X1 U6398 ( .A1(n4598), .A2(n4521), .ZN(n6364) );
  NAND3_X1 U6399 ( .A1(n6152), .A2(n6151), .A3(n6153), .ZN(n6593) );
  NAND2_X1 U6400 ( .A1(n5106), .A2(n5104), .ZN(n5108) );
  NAND2_X1 U6401 ( .A1(n8552), .A2(n5111), .ZN(n5110) );
  OAI21_X1 U6402 ( .B1(n8500), .B2(n5125), .A(n5126), .ZN(n8477) );
  INV_X1 U6403 ( .A(n5121), .ZN(n6549) );
  OAI21_X1 U6404 ( .B1(n8500), .B2(n5124), .A(n5122), .ZN(n5121) );
  NAND4_X1 U6405 ( .A1(n5174), .A2(n5173), .A3(n5172), .A4(n5171), .ZN(n5832)
         );
  AND2_X1 U6406 ( .A1(n7061), .A2(n5765), .ZN(n8965) );
  NAND2_X1 U6407 ( .A1(n5169), .A2(n5168), .ZN(n5336) );
  OR2_X1 U6408 ( .A1(n5244), .A2(n5243), .ZN(n5245) );
  NAND3_X2 U6409 ( .A1(n5188), .A2(n5187), .A3(n5186), .ZN(n6958) );
  NAND2_X1 U6410 ( .A1(n6570), .A2(n6569), .ZN(n7878) );
  NAND2_X1 U6411 ( .A1(n6888), .A2(n7513), .ZN(n6889) );
  NAND2_X1 U6412 ( .A1(n6562), .A2(n6866), .ZN(n6868) );
  OR2_X1 U6413 ( .A1(n7328), .A2(n7225), .ZN(n6210) );
  NAND4_X2 U6414 ( .A1(n5227), .A2(n5226), .A3(n5225), .A4(n5224), .ZN(n9264)
         );
  OR2_X1 U6415 ( .A1(n5244), .A2(n5223), .ZN(n5224) );
  NAND2_X1 U6416 ( .A1(n5718), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5227) );
  NAND2_X1 U6417 ( .A1(n8191), .A2(n4689), .ZN(n8193) );
  INV_X1 U6418 ( .A(n8145), .ZN(n7513) );
  OR3_X1 U6419 ( .A1(n8579), .A2(n8578), .A3(n8593), .ZN(n8582) );
  OAI21_X2 U6420 ( .B1(n8499), .B2(n8064), .A(n8062), .ZN(n8491) );
  AND2_X2 U6421 ( .A1(n9726), .A2(n5168), .ZN(n5264) );
  AND2_X1 U6422 ( .A1(n6088), .A2(n9223), .ZN(n7872) );
  OR2_X1 U6423 ( .A1(n6123), .A2(n7099), .ZN(n9916) );
  INV_X1 U6424 ( .A(n8306), .ZN(n6486) );
  AND2_X1 U6426 ( .A1(n6634), .A2(n6633), .ZN(n5136) );
  OR2_X1 U6427 ( .A1(n9360), .A2(n9652), .ZN(n5137) );
  OR2_X1 U6428 ( .A1(n9360), .A2(n9713), .ZN(n5138) );
  INV_X2 U6429 ( .A(n10149), .ZN(n10148) );
  NAND2_X1 U6430 ( .A1(n6516), .A2(n6515), .ZN(n8521) );
  INV_X1 U6431 ( .A(n10159), .ZN(n10157) );
  INV_X1 U6432 ( .A(n9652), .ZN(n6638) );
  NOR2_X1 U6433 ( .A1(n7083), .A2(n7172), .ZN(n5140) );
  INV_X1 U6434 ( .A(n5823), .ZN(n5824) );
  INV_X1 U6435 ( .A(n6632), .ZN(n7922) );
  INV_X1 U6436 ( .A(n8120), .ZN(n6320) );
  AND2_X1 U6437 ( .A1(n8666), .A2(n8569), .ZN(n5141) );
  OR2_X1 U6438 ( .A1(n9502), .A2(n9248), .ZN(n5142) );
  INV_X1 U6439 ( .A(n6119), .ZN(n9360) );
  OR2_X1 U6440 ( .A1(n8005), .A2(n7734), .ZN(n5143) );
  AND4_X2 U6441 ( .A1(n6210), .A2(n6209), .A3(n6208), .A4(n6207), .ZN(n6224)
         );
  AND2_X1 U6442 ( .A1(n7420), .A2(n7419), .ZN(n5144) );
  AND2_X1 U6443 ( .A1(n7084), .A2(n8315), .ZN(n5145) );
  AND2_X1 U6444 ( .A1(n9163), .A2(n8992), .ZN(n5146) );
  OR2_X1 U6445 ( .A1(n7640), .A2(n8842), .ZN(n5147) );
  NAND2_X1 U6446 ( .A1(n8984), .A2(n8983), .ZN(n8985) );
  AND2_X1 U6447 ( .A1(n9104), .A2(n9014), .ZN(n9015) );
  AOI21_X1 U6448 ( .B1(n9017), .B2(n9016), .A(n9015), .ZN(n9018) );
  OR2_X1 U6449 ( .A1(n9026), .A2(n9025), .ZN(n9027) );
  AND2_X1 U6450 ( .A1(n9027), .A2(n9034), .ZN(n9028) );
  INV_X1 U6451 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n6141) );
  NAND2_X1 U6452 ( .A1(n7421), .A2(n7417), .ZN(n7420) );
  OR2_X1 U6453 ( .A1(n8000), .A2(n8309), .ZN(n6386) );
  INV_X1 U6454 ( .A(n7375), .ZN(n6268) );
  NOR4_X1 U6455 ( .A1(n9088), .A2(n9087), .A3(n9086), .A4(n9085), .ZN(n9090)
         );
  INV_X1 U6456 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5161) );
  NAND2_X1 U6457 ( .A1(n6347), .A2(n6346), .ZN(n6348) );
  INV_X1 U6458 ( .A(n8161), .ZN(n6190) );
  INV_X1 U6459 ( .A(n6510), .ZN(n6181) );
  INV_X1 U6460 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n6398) );
  INV_X1 U6461 ( .A(n5497), .ZN(n5495) );
  INV_X1 U6462 ( .A(n5593), .ZN(n5591) );
  OR2_X1 U6463 ( .A1(n9375), .A2(n9241), .ZN(n5708) );
  INV_X1 U6464 ( .A(n5565), .ZN(n5563) );
  INV_X1 U6465 ( .A(n5439), .ZN(n5438) );
  INV_X1 U6466 ( .A(n7024), .ZN(n5722) );
  INV_X1 U6467 ( .A(n5544), .ZN(n5547) );
  INV_X1 U6468 ( .A(n6480), .ZN(n6177) );
  OR2_X1 U6469 ( .A1(n5536), .A2(n5535), .ZN(n5565) );
  AND2_X1 U6470 ( .A1(n9064), .A2(n9065), .ZN(n9131) );
  OR2_X1 U6471 ( .A1(n9485), .A2(n9247), .ZN(n5583) );
  OR2_X1 U6472 ( .A1(n5477), .A2(n5476), .ZN(n5497) );
  OR2_X1 U6473 ( .A1(n5419), .A2(n5418), .ZN(n5439) );
  INV_X1 U6474 ( .A(n9219), .ZN(n6698) );
  NAND2_X1 U6475 ( .A1(n5743), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5531) );
  NAND2_X1 U6476 ( .A1(n5396), .A2(n5395), .ZN(n5408) );
  OR2_X1 U6477 ( .A1(n5315), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n5375) );
  NAND2_X1 U6478 ( .A1(n5273), .A2(SI_4_), .ZN(n5274) );
  AND2_X1 U6479 ( .A1(n8194), .A2(n8502), .ZN(n8195) );
  NAND2_X1 U6480 ( .A1(n6177), .A2(n10315), .ZN(n6489) );
  OR2_X1 U6481 ( .A1(n6489), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6499) );
  INV_X1 U6482 ( .A(n8521), .ZN(n8298) );
  NAND2_X1 U6483 ( .A1(n8141), .A2(n7529), .ZN(n8142) );
  AND2_X1 U6484 ( .A1(n6202), .A2(n6201), .ZN(n8242) );
  NOR2_X1 U6485 ( .A1(n7767), .A2(n9990), .ZN(n10011) );
  INV_X1 U6486 ( .A(n8463), .ZN(n8444) );
  OR2_X1 U6487 ( .A1(n6530), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n7921) );
  OR2_X1 U6488 ( .A1(n6519), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n6521) );
  OR2_X1 U6489 ( .A1(n10119), .A2(n7942), .ZN(n8523) );
  OR2_X1 U6490 ( .A1(n8087), .A2(n6907), .ZN(n8598) );
  AND2_X1 U6491 ( .A1(n7942), .A2(n7688), .ZN(n6990) );
  AND2_X1 U6492 ( .A1(n8878), .A2(n6037), .ZN(n8800) );
  AND2_X1 U6493 ( .A1(n6698), .A2(n5757), .ZN(n8932) );
  AND2_X1 U6494 ( .A1(n6028), .A2(n6027), .ZN(n8904) );
  OR2_X1 U6495 ( .A1(n5630), .A2(n8803), .ZN(n5666) );
  OR2_X1 U6496 ( .A1(n5610), .A2(n8911), .ZN(n5630) );
  OR2_X1 U6497 ( .A1(n6826), .A2(n6825), .ZN(n6837) );
  AND2_X1 U6498 ( .A1(n9053), .A2(n9182), .ZN(n9497) );
  AND2_X1 U6499 ( .A1(n7357), .A2(n8992), .ZN(n7358) );
  INV_X1 U6500 ( .A(n8932), .ZN(n8946) );
  AND2_X1 U6501 ( .A1(n9099), .A2(n7530), .ZN(n6088) );
  AND2_X1 U6502 ( .A1(n5764), .A2(n9097), .ZN(n9571) );
  XNOR2_X1 U6503 ( .A(n5428), .B(SI_12_), .ZN(n5427) );
  AND2_X1 U6504 ( .A1(n6908), .A2(n6902), .ZN(n8300) );
  INV_X1 U6505 ( .A(n8082), .ZN(n8470) );
  AND2_X1 U6506 ( .A1(n6526), .A2(n6525), .ZN(n8293) );
  INV_X1 U6507 ( .A(n10051), .ZN(n10069) );
  NAND2_X1 U6508 ( .A1(n7205), .A2(n10097), .ZN(n8610) );
  INV_X1 U6509 ( .A(n8662), .ZN(n8678) );
  NAND2_X1 U6510 ( .A1(n8025), .A2(n8032), .ZN(n8606) );
  INV_X1 U6511 ( .A(n8733), .ZN(n8756) );
  OAI211_X1 U6512 ( .C1(n6587), .C2(n7780), .A(n6265), .B(n6264), .ZN(n10117)
         );
  INV_X1 U6513 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n6595) );
  INV_X1 U6514 ( .A(n6107), .ZN(n6108) );
  NAND2_X1 U6515 ( .A1(n6090), .A2(n9717), .ZN(n9869) );
  AND2_X1 U6516 ( .A1(n5717), .A2(n9347), .ZN(n9358) );
  AND4_X1 U6517 ( .A1(n5502), .A2(n5501), .A3(n5500), .A4(n5499), .ZN(n8869)
         );
  INV_X1 U6518 ( .A(n9832), .ZN(n10559) );
  INV_X1 U6519 ( .A(n9861), .ZN(n9535) );
  INV_X1 U6520 ( .A(n9873), .ZN(n9866) );
  NOR2_X1 U6521 ( .A1(n9586), .A2(n9585), .ZN(n9662) );
  XNOR2_X1 U6522 ( .A(n5272), .B(SI_4_), .ZN(n5270) );
  XNOR2_X1 U6523 ( .A(n5256), .B(SI_3_), .ZN(n5254) );
  OAI211_X1 U6524 ( .C1(n5064), .C2(n8206), .A(n8205), .B(n4548), .ZN(n8210)
         );
  INV_X1 U6525 ( .A(n8719), .ZN(n8524) );
  AND2_X1 U6526 ( .A1(n6899), .A2(n6898), .ZN(n8267) );
  INV_X1 U6527 ( .A(n8263), .ZN(n8303) );
  INV_X1 U6528 ( .A(n8293), .ZN(n8509) );
  INV_X1 U6529 ( .A(n7734), .ZN(n8308) );
  INV_X1 U6530 ( .A(n7426), .ZN(n8311) );
  OR2_X1 U6531 ( .A1(n9919), .A2(n8779), .ZN(n10089) );
  INV_X1 U6532 ( .A(n8562), .ZN(n8630) );
  AOI21_X1 U6533 ( .B1(n6632), .B2(n8756), .A(n6650), .ZN(n6651) );
  INV_X1 U6534 ( .A(n8175), .ZN(n8734) );
  AND2_X1 U6535 ( .A1(n6649), .A2(n6648), .ZN(n10149) );
  INV_X1 U6536 ( .A(n6691), .ZN(n6695) );
  INV_X1 U6537 ( .A(n6888), .ZN(n7529) );
  INV_X1 U6538 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n10382) );
  INV_X1 U6539 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6688) );
  AND2_X1 U6540 ( .A1(n6091), .A2(n9869), .ZN(n9766) );
  INV_X1 U6541 ( .A(n6056), .ZN(n9242) );
  INV_X1 U6542 ( .A(n10566), .ZN(n9853) );
  OR2_X1 U6543 ( .A1(n9857), .A2(n7102), .ZN(n9861) );
  NAND2_X1 U6544 ( .A1(n9918), .A2(n9656), .ZN(n9652) );
  INV_X2 U6545 ( .A(n9916), .ZN(n9918) );
  INV_X1 U6546 ( .A(n9420), .ZN(n9682) );
  NAND2_X1 U6547 ( .A1(n9911), .A2(n9656), .ZN(n9713) );
  OR2_X1 U6548 ( .A1(n6123), .A2(n5826), .ZN(n9910) );
  INV_X1 U6549 ( .A(n9883), .ZN(n9884) );
  INV_X1 U6550 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n10457) );
  INV_X1 U6551 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6664) );
  INV_X1 U6552 ( .A(n8428), .ZN(P2_U3893) );
  NAND4_X1 U6553 ( .A1(n5150), .A2(n5279), .A3(n5149), .A4(n5372), .ZN(n5153)
         );
  NOR2_X1 U6554 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n5151) );
  NAND2_X1 U6555 ( .A1(n5373), .A2(n5151), .ZN(n5152) );
  NOR3_X1 U6556 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_24__SCAN_IN), .A3(
        P1_IR_REG_23__SCAN_IN), .ZN(n5159) );
  NOR2_X1 U6557 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), .ZN(
        n5158) );
  NOR2_X1 U6558 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), .ZN(
        n5157) );
  NOR2_X1 U6559 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n5156) );
  NAND4_X1 U6560 ( .A1(n5159), .A2(n5158), .A3(n5157), .A4(n5156), .ZN(n5160)
         );
  NOR2_X2 U6561 ( .A1(n5175), .A2(P1_IR_REG_28__SCAN_IN), .ZN(n5164) );
  XNOR2_X2 U6562 ( .A(n5162), .B(n5163), .ZN(n9726) );
  NAND2_X1 U6563 ( .A1(n5164), .A2(n5163), .ZN(n9720) );
  INV_X1 U6564 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n5165) );
  XNOR2_X2 U6565 ( .A(n5166), .B(n5165), .ZN(n5168) );
  INV_X2 U6566 ( .A(n5168), .ZN(n5170) );
  NAND2_X4 U6567 ( .A1(n9726), .A2(n5170), .ZN(n6709) );
  INV_X1 U6568 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n5167) );
  NAND2_X1 U6569 ( .A1(n5732), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n5173) );
  NAND2_X1 U6570 ( .A1(n5264), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n5172) );
  NAND2_X4 U6571 ( .A1(n5170), .A2(n5169), .ZN(n5687) );
  INV_X1 U6572 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n6961) );
  NAND2_X1 U6573 ( .A1(n5175), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5177) );
  INV_X1 U6574 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5176) );
  AND2_X4 U6575 ( .A1(n5182), .A2(n5181), .ZN(n7936) );
  INV_X1 U6576 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6667) );
  OR2_X1 U6577 ( .A1(n5234), .A2(n6667), .ZN(n5188) );
  AND2_X1 U6578 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n5183) );
  INV_X1 U6579 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n5185) );
  NAND2_X1 U6580 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5184) );
  XNOR2_X1 U6581 ( .A(n5185), .B(n5184), .ZN(n6812) );
  OR2_X1 U6582 ( .A1(n8962), .A2(n6812), .ZN(n5186) );
  NAND2_X1 U6583 ( .A1(n5840), .A2(n9872), .ZN(n9153) );
  INV_X1 U6584 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n5189) );
  OR2_X1 U6585 ( .A1(n5244), .A2(n5189), .ZN(n5194) );
  INV_X1 U6586 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n6921) );
  OR2_X1 U6587 ( .A1(n6709), .A2(n6921), .ZN(n5193) );
  INV_X2 U6588 ( .A(n5336), .ZN(n5732) );
  NAND2_X1 U6589 ( .A1(n5732), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5192) );
  INV_X1 U6590 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n5190) );
  OR2_X1 U6591 ( .A1(n5687), .A2(n5190), .ZN(n5191) );
  INV_X1 U6592 ( .A(SI_0_), .ZN(n5196) );
  INV_X1 U6593 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5195) );
  OAI21_X1 U6594 ( .B1(n7936), .B2(n5196), .A(n5195), .ZN(n5198) );
  AND2_X1 U6595 ( .A1(n5198), .A2(n5197), .ZN(n9740) );
  MUX2_X1 U6596 ( .A(P1_IR_REG_0__SCAN_IN), .B(n9740), .S(n8962), .Z(n6976) );
  NAND2_X1 U6597 ( .A1(n7074), .A2(n6976), .ZN(n7060) );
  NAND2_X1 U6598 ( .A1(n9107), .A2(n7060), .ZN(n5200) );
  NAND2_X1 U6599 ( .A1(n4752), .A2(n9872), .ZN(n5199) );
  NAND2_X1 U6600 ( .A1(n5200), .A2(n5199), .ZN(n7097) );
  INV_X1 U6601 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n7108) );
  NAND2_X1 U6602 ( .A1(n5732), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5204) );
  INV_X1 U6603 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n5201) );
  OR2_X1 U6604 ( .A1(n5244), .A2(n5201), .ZN(n5203) );
  INV_X1 U6605 ( .A(n6709), .ZN(n5596) );
  NAND2_X1 U6606 ( .A1(n5596), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5202) );
  OR2_X1 U6607 ( .A1(n5234), .A2(n6666), .ZN(n5220) );
  NAND2_X1 U6608 ( .A1(n5209), .A2(SI_1_), .ZN(n5210) );
  NAND2_X1 U6609 ( .A1(n5211), .A2(n5210), .ZN(n5229) );
  MUX2_X1 U6610 ( .A(n6659), .B(n6666), .S(n5431), .Z(n5230) );
  XNOR2_X1 U6611 ( .A(n5230), .B(SI_2_), .ZN(n5228) );
  XNOR2_X1 U6612 ( .A(n5229), .B(n5228), .ZN(n6665) );
  OR2_X1 U6613 ( .A1(n5206), .A2(n6665), .ZN(n5219) );
  NOR2_X1 U6614 ( .A1(n5212), .A2(n5276), .ZN(n5213) );
  MUX2_X1 U6615 ( .A(n5276), .B(n5213), .S(P1_IR_REG_2__SCAN_IN), .Z(n5214) );
  INV_X1 U6616 ( .A(n5214), .ZN(n5217) );
  INV_X1 U6617 ( .A(n5215), .ZN(n5216) );
  NAND2_X1 U6618 ( .A1(n5217), .A2(n5216), .ZN(n6931) );
  OR2_X1 U6619 ( .A1(n8962), .A2(n6931), .ZN(n5218) );
  NAND2_X1 U6620 ( .A1(n7097), .A2(n9105), .ZN(n5222) );
  OR2_X1 U6621 ( .A1(n5852), .A2(n7112), .ZN(n5221) );
  NAND2_X1 U6622 ( .A1(n5732), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n5226) );
  OR2_X1 U6623 ( .A1(n5687), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n5225) );
  INV_X1 U6624 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n5223) );
  NAND2_X1 U6625 ( .A1(n5229), .A2(n5228), .ZN(n5233) );
  INV_X1 U6626 ( .A(n5230), .ZN(n5231) );
  NAND2_X1 U6627 ( .A1(n5231), .A2(SI_2_), .ZN(n5232) );
  NAND2_X1 U6628 ( .A1(n5233), .A2(n5232), .ZN(n5255) );
  XNOR2_X1 U6629 ( .A(n5255), .B(n5254), .ZN(n6668) );
  OR2_X1 U6630 ( .A1(n5206), .A2(n6668), .ZN(n5237) );
  OR2_X1 U6631 ( .A1(n5234), .A2(n6669), .ZN(n5236) );
  OR2_X1 U6632 ( .A1(n5215), .A2(n5276), .ZN(n5250) );
  INV_X1 U6633 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n5249) );
  XNOR2_X1 U6634 ( .A(n5250), .B(n5249), .ZN(n6815) );
  OR2_X1 U6635 ( .A1(n8962), .A2(n6815), .ZN(n5235) );
  NAND2_X1 U6636 ( .A1(n9264), .A2(n9893), .ZN(n8981) );
  NAND2_X1 U6637 ( .A1(n9155), .A2(n8981), .ZN(n9108) );
  INV_X1 U6638 ( .A(n9893), .ZN(n8812) );
  OR2_X1 U6639 ( .A1(n9264), .A2(n8812), .ZN(n5238) );
  NAND2_X1 U6640 ( .A1(n5732), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5248) );
  INV_X1 U6641 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6817) );
  OR2_X1 U6642 ( .A1(n6709), .A2(n6817), .ZN(n5247) );
  INV_X1 U6643 ( .A(n5263), .ZN(n5242) );
  INV_X1 U6644 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n5240) );
  INV_X1 U6645 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n5239) );
  NAND2_X1 U6646 ( .A1(n5240), .A2(n5239), .ZN(n5241) );
  NAND2_X1 U6647 ( .A1(n5242), .A2(n5241), .ZN(n9854) );
  OR2_X1 U6648 ( .A1(n5687), .A2(n9854), .ZN(n5246) );
  INV_X1 U6649 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n5243) );
  NAND2_X1 U6650 ( .A1(n5250), .A2(n5249), .ZN(n5251) );
  NAND2_X1 U6651 ( .A1(n5251), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5253) );
  INV_X1 U6652 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n5252) );
  XNOR2_X1 U6653 ( .A(n5253), .B(n5252), .ZN(n6949) );
  NAND2_X1 U6654 ( .A1(n5255), .A2(n5254), .ZN(n5259) );
  INV_X1 U6655 ( .A(n5256), .ZN(n5257) );
  NAND2_X1 U6656 ( .A1(n5257), .A2(SI_3_), .ZN(n5258) );
  XNOR2_X1 U6657 ( .A(n5271), .B(n5270), .ZN(n6663) );
  OR2_X1 U6658 ( .A1(n5206), .A2(n6663), .ZN(n5261) );
  OR2_X1 U6659 ( .A1(n5234), .A2(n6664), .ZN(n5260) );
  OAI211_X1 U6660 ( .C1(n8962), .C2(n6949), .A(n5261), .B(n5260), .ZN(n9865)
         );
  NOR2_X1 U6661 ( .A1(n9263), .A2(n9865), .ZN(n7149) );
  NAND2_X1 U6662 ( .A1(n9263), .A2(n9865), .ZN(n7148) );
  NAND2_X1 U6663 ( .A1(n5262), .A2(n7148), .ZN(n7213) );
  NAND2_X1 U6664 ( .A1(n5732), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5269) );
  NAND2_X1 U6665 ( .A1(n5718), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n5268) );
  OAI21_X1 U6666 ( .B1(n5263), .B2(P1_REG3_REG_5__SCAN_IN), .A(n5302), .ZN(
        n7220) );
  OR2_X1 U6667 ( .A1(n5595), .A2(n7220), .ZN(n5267) );
  INV_X1 U6668 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n5265) );
  OR2_X1 U6669 ( .A1(n5244), .A2(n5265), .ZN(n5266) );
  NAND4_X1 U6670 ( .A1(n5269), .A2(n5268), .A3(n5267), .A4(n5266), .ZN(n9262)
         );
  INV_X1 U6671 ( .A(n5272), .ZN(n5273) );
  XNOR2_X1 U6672 ( .A(n5293), .B(n5291), .ZN(n6670) );
  NAND2_X1 U6673 ( .A1(n5295), .A2(n6670), .ZN(n5283) );
  NOR2_X1 U6674 ( .A1(n5275), .A2(n5276), .ZN(n5277) );
  MUX2_X1 U6675 ( .A(n5276), .B(n5277), .S(P1_IR_REG_5__SCAN_IN), .Z(n5278) );
  INV_X1 U6676 ( .A(n5278), .ZN(n5280) );
  NAND2_X1 U6677 ( .A1(n5275), .A2(n5279), .ZN(n5315) );
  NAND2_X1 U6678 ( .A1(n5280), .A2(n5315), .ZN(n9279) );
  OR2_X1 U6679 ( .A1(n8962), .A2(n9279), .ZN(n5282) );
  INV_X1 U6680 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6671) );
  OR2_X1 U6681 ( .A1(n5234), .A2(n6671), .ZN(n5281) );
  NAND2_X1 U6682 ( .A1(n9262), .A2(n7409), .ZN(n9163) );
  NAND2_X1 U6683 ( .A1(n8990), .A2(n9163), .ZN(n7212) );
  NAND2_X1 U6684 ( .A1(n5732), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n5289) );
  INV_X1 U6685 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n7247) );
  OR2_X1 U6686 ( .A1(n6709), .A2(n7247), .ZN(n5288) );
  INV_X1 U6687 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n5284) );
  XNOR2_X1 U6688 ( .A(n5302), .B(n5284), .ZN(n7246) );
  OR2_X1 U6689 ( .A1(n5687), .A2(n7246), .ZN(n5287) );
  INV_X1 U6690 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n5285) );
  OR2_X1 U6691 ( .A1(n5244), .A2(n5285), .ZN(n5286) );
  NAND4_X1 U6692 ( .A1(n5289), .A2(n5288), .A3(n5287), .A4(n5286), .ZN(n9261)
         );
  NAND2_X1 U6693 ( .A1(n5315), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5290) );
  XNOR2_X1 U6694 ( .A(n5290), .B(P1_IR_REG_6__SCAN_IN), .ZN(n9296) );
  AOI22_X1 U6695 ( .A1(n5560), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n5559), .B2(
        n9296), .ZN(n5297) );
  XNOR2_X1 U6696 ( .A(n5311), .B(n5309), .ZN(n6677) );
  NAND2_X1 U6697 ( .A1(n6677), .A2(n5295), .ZN(n5296) );
  OR2_X1 U6698 ( .A1(n9261), .A2(n7353), .ZN(n9113) );
  NAND2_X1 U6699 ( .A1(n9261), .A2(n7353), .ZN(n8992) );
  NAND2_X1 U6700 ( .A1(n9113), .A2(n8992), .ZN(n7239) );
  NAND2_X1 U6701 ( .A1(n7238), .A2(n7239), .ZN(n7237) );
  INV_X1 U6702 ( .A(n9261), .ZN(n5298) );
  NAND2_X1 U6703 ( .A1(n5298), .A2(n7353), .ZN(n5299) );
  NAND2_X1 U6704 ( .A1(n7237), .A2(n5299), .ZN(n7363) );
  NAND2_X1 U6705 ( .A1(n5718), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n5308) );
  NAND2_X1 U6706 ( .A1(n5732), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n5307) );
  INV_X1 U6707 ( .A(n5302), .ZN(n5300) );
  AOI21_X1 U6708 ( .B1(n5300), .B2(P1_REG3_REG_6__SCAN_IN), .A(
        P1_REG3_REG_7__SCAN_IN), .ZN(n5303) );
  NAND2_X1 U6709 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_REG3_REG_7__SCAN_IN), 
        .ZN(n5301) );
  OR2_X1 U6710 ( .A1(n5303), .A2(n5337), .ZN(n7342) );
  OR2_X1 U6711 ( .A1(n5687), .A2(n7342), .ZN(n5306) );
  INV_X1 U6712 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n5304) );
  OR2_X1 U6713 ( .A1(n5244), .A2(n5304), .ZN(n5305) );
  NAND4_X1 U6714 ( .A1(n5308), .A2(n5307), .A3(n5306), .A4(n5305), .ZN(n9260)
         );
  NAND2_X1 U6715 ( .A1(n5311), .A2(n5310), .ZN(n5314) );
  NAND2_X1 U6716 ( .A1(n5312), .A2(SI_6_), .ZN(n5313) );
  XNOR2_X1 U6717 ( .A(n5322), .B(n5320), .ZN(n6681) );
  NAND2_X1 U6718 ( .A1(n6681), .A2(n5295), .ZN(n5317) );
  NAND2_X1 U6719 ( .A1(n5375), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5332) );
  XNOR2_X1 U6720 ( .A(n5332), .B(P1_IR_REG_7__SCAN_IN), .ZN(n9309) );
  AOI22_X1 U6721 ( .A1(n5560), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n5559), .B2(
        n9309), .ZN(n5316) );
  OR2_X1 U6722 ( .A1(n9260), .A2(n9898), .ZN(n7466) );
  NAND2_X1 U6723 ( .A1(n9898), .A2(n9260), .ZN(n8994) );
  NAND2_X1 U6724 ( .A1(n7466), .A2(n8994), .ZN(n8988) );
  NAND2_X1 U6725 ( .A1(n7363), .A2(n8988), .ZN(n7362) );
  INV_X1 U6726 ( .A(n9260), .ZN(n5318) );
  NAND2_X1 U6727 ( .A1(n5318), .A2(n9898), .ZN(n5319) );
  NAND2_X1 U6728 ( .A1(n7362), .A2(n5319), .ZN(n7473) );
  INV_X1 U6729 ( .A(SI_8_), .ZN(n5325) );
  INV_X1 U6730 ( .A(n5326), .ZN(n5327) );
  NAND2_X1 U6731 ( .A1(n5327), .A2(SI_8_), .ZN(n5328) );
  NAND2_X1 U6732 ( .A1(n5330), .A2(n5329), .ZN(n5331) );
  NAND2_X1 U6733 ( .A1(n5346), .A2(n5331), .ZN(n6685) );
  NAND2_X1 U6734 ( .A1(n6685), .A2(n5295), .ZN(n5335) );
  NAND2_X1 U6735 ( .A1(n5332), .A2(n5372), .ZN(n5333) );
  NAND2_X1 U6736 ( .A1(n5333), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5356) );
  XNOR2_X1 U6737 ( .A(n5356), .B(P1_IR_REG_8__SCAN_IN), .ZN(n9321) );
  AOI22_X1 U6738 ( .A1(n5560), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n5559), .B2(
        n9321), .ZN(n5334) );
  NAND2_X1 U6739 ( .A1(n5335), .A2(n5334), .ZN(n7601) );
  NAND2_X1 U6740 ( .A1(n5718), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n5343) );
  INV_X1 U6741 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n6805) );
  OR2_X1 U6742 ( .A1(n6712), .A2(n6805), .ZN(n5342) );
  NOR2_X1 U6743 ( .A1(n5337), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n5338) );
  OR2_X1 U6744 ( .A1(n5361), .A2(n5338), .ZN(n7594) );
  OR2_X1 U6745 ( .A1(n5595), .A2(n7594), .ZN(n5341) );
  INV_X1 U6746 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n5339) );
  OR2_X1 U6747 ( .A1(n5244), .A2(n5339), .ZN(n5340) );
  OR2_X1 U6748 ( .A1(n7601), .A2(n7498), .ZN(n8995) );
  NAND2_X1 U6749 ( .A1(n7601), .A2(n7498), .ZN(n8999) );
  NAND2_X1 U6750 ( .A1(n8995), .A2(n8999), .ZN(n7472) );
  NAND2_X1 U6751 ( .A1(n7473), .A2(n7472), .ZN(n7471) );
  INV_X1 U6752 ( .A(n7498), .ZN(n9259) );
  OR2_X1 U6753 ( .A1(n7601), .A2(n9259), .ZN(n5344) );
  NAND2_X1 U6754 ( .A1(n7471), .A2(n5344), .ZN(n7502) );
  INV_X1 U6755 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n5347) );
  INV_X1 U6756 ( .A(SI_9_), .ZN(n5348) );
  NAND2_X1 U6757 ( .A1(n5349), .A2(n5348), .ZN(n5369) );
  INV_X1 U6758 ( .A(n5349), .ZN(n5350) );
  NAND2_X1 U6759 ( .A1(n5350), .A2(SI_9_), .ZN(n5351) );
  NAND2_X1 U6760 ( .A1(n6696), .A2(n5295), .ZN(n5360) );
  INV_X1 U6761 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n5355) );
  NAND2_X1 U6762 ( .A1(n5356), .A2(n5355), .ZN(n5357) );
  NAND2_X1 U6763 ( .A1(n5357), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5358) );
  XNOR2_X1 U6764 ( .A(n5358), .B(P1_IR_REG_9__SCAN_IN), .ZN(n6843) );
  AOI22_X1 U6765 ( .A1(n5560), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n5559), .B2(
        n6843), .ZN(n5359) );
  NAND2_X1 U6766 ( .A1(n5731), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5367) );
  INV_X1 U6767 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n7506) );
  OR2_X1 U6768 ( .A1(n6709), .A2(n7506), .ZN(n5366) );
  NOR2_X1 U6769 ( .A1(n5361), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n5362) );
  OR2_X1 U6770 ( .A1(n5379), .A2(n5362), .ZN(n7658) );
  OR2_X1 U6771 ( .A1(n5687), .A2(n7658), .ZN(n5365) );
  INV_X1 U6772 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n5363) );
  OR2_X1 U6773 ( .A1(n6712), .A2(n5363), .ZN(n5364) );
  OR2_X1 U6774 ( .A1(n7660), .A2(n7484), .ZN(n9008) );
  NAND2_X1 U6775 ( .A1(n7660), .A2(n7484), .ZN(n9004) );
  NAND2_X1 U6776 ( .A1(n9008), .A2(n9004), .ZN(n7501) );
  NAND2_X1 U6777 ( .A1(n7502), .A2(n7501), .ZN(n7500) );
  INV_X1 U6778 ( .A(n7484), .ZN(n9258) );
  OR2_X1 U6779 ( .A1(n7660), .A2(n9258), .ZN(n5368) );
  NAND2_X1 U6780 ( .A1(n7500), .A2(n5368), .ZN(n7489) );
  INV_X1 U6781 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n5371) );
  NAND2_X1 U6782 ( .A1(n6705), .A2(n5295), .ZN(n5378) );
  NAND2_X1 U6783 ( .A1(n5373), .A2(n5372), .ZN(n5374) );
  NOR2_X1 U6784 ( .A1(n5375), .A2(n5374), .ZN(n5400) );
  OR2_X1 U6785 ( .A1(n5400), .A2(n5276), .ZN(n5376) );
  XNOR2_X1 U6786 ( .A(n5376), .B(P1_IR_REG_10__SCAN_IN), .ZN(n9748) );
  AOI22_X1 U6787 ( .A1(n5560), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n5559), .B2(
        n9748), .ZN(n5377) );
  NAND2_X1 U6788 ( .A1(n5731), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5386) );
  INV_X1 U6789 ( .A(n5379), .ZN(n5381) );
  INV_X1 U6790 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n5380) );
  NAND2_X1 U6791 ( .A1(n5381), .A2(n5380), .ZN(n5382) );
  NAND2_X1 U6792 ( .A1(n5419), .A2(n5382), .ZN(n9771) );
  OR2_X1 U6793 ( .A1(n5687), .A2(n9771), .ZN(n5385) );
  INV_X1 U6794 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n7490) );
  OR2_X1 U6795 ( .A1(n6709), .A2(n7490), .ZN(n5384) );
  INV_X1 U6796 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n6846) );
  OR2_X1 U6797 ( .A1(n6712), .A2(n6846), .ZN(n5383) );
  OR2_X1 U6798 ( .A1(n7538), .A2(n7634), .ZN(n9170) );
  NAND2_X1 U6799 ( .A1(n7538), .A2(n7634), .ZN(n9010) );
  INV_X1 U6800 ( .A(n7634), .ZN(n9257) );
  OR2_X1 U6801 ( .A1(n7538), .A2(n9257), .ZN(n5387) );
  INV_X1 U6802 ( .A(n5389), .ZN(n5390) );
  INV_X1 U6803 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n5394) );
  INV_X1 U6804 ( .A(SI_11_), .ZN(n5395) );
  INV_X1 U6805 ( .A(n5396), .ZN(n5397) );
  NAND2_X1 U6806 ( .A1(n5397), .A2(SI_11_), .ZN(n5398) );
  NAND2_X1 U6807 ( .A1(n6718), .A2(n5295), .ZN(n5403) );
  INV_X1 U6808 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n5399) );
  NAND2_X1 U6809 ( .A1(n5400), .A2(n5399), .ZN(n5411) );
  NAND2_X1 U6810 ( .A1(n5411), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5401) );
  XNOR2_X1 U6811 ( .A(n5401), .B(P1_IR_REG_11__SCAN_IN), .ZN(n9787) );
  AOI22_X1 U6812 ( .A1(n5560), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n5559), .B2(
        n9787), .ZN(n5402) );
  NAND2_X1 U6813 ( .A1(n5731), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5407) );
  INV_X1 U6814 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n5417) );
  XNOR2_X1 U6815 ( .A(n5419), .B(n5417), .ZN(n8924) );
  OR2_X1 U6816 ( .A1(n5595), .A2(n8924), .ZN(n5406) );
  INV_X1 U6817 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n7643) );
  OR2_X1 U6818 ( .A1(n6709), .A2(n7643), .ZN(n5405) );
  INV_X1 U6819 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n6847) );
  OR2_X1 U6820 ( .A1(n6712), .A2(n6847), .ZN(n5404) );
  OR2_X1 U6821 ( .A1(n8926), .A2(n7606), .ZN(n9006) );
  NAND2_X1 U6822 ( .A1(n8926), .A2(n7606), .ZN(n9013) );
  NAND2_X1 U6823 ( .A1(n9006), .A2(n9013), .ZN(n7633) );
  INV_X1 U6824 ( .A(n7606), .ZN(n9256) );
  XNOR2_X1 U6825 ( .A(n5430), .B(n5427), .ZN(n6833) );
  NAND2_X1 U6826 ( .A1(n6833), .A2(n5295), .ZN(n5414) );
  OR2_X1 U6827 ( .A1(n5411), .A2(P1_IR_REG_11__SCAN_IN), .ZN(n5412) );
  NAND2_X1 U6828 ( .A1(n5412), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5433) );
  XNOR2_X1 U6829 ( .A(n5433), .B(P1_IR_REG_12__SCAN_IN), .ZN(n7556) );
  AOI22_X1 U6830 ( .A1(n5560), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n5559), .B2(
        n7556), .ZN(n5413) );
  INV_X1 U6831 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n7614) );
  OR2_X1 U6832 ( .A1(n6709), .A2(n7614), .ZN(n5425) );
  INV_X1 U6833 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n5415) );
  OR2_X1 U6834 ( .A1(n5244), .A2(n5415), .ZN(n5424) );
  INV_X1 U6835 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n5416) );
  OAI21_X1 U6836 ( .B1(n5419), .B2(n5417), .A(n5416), .ZN(n5420) );
  NAND2_X1 U6837 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_REG3_REG_12__SCAN_IN), 
        .ZN(n5418) );
  NAND2_X1 U6838 ( .A1(n5420), .A2(n5439), .ZN(n8840) );
  OR2_X1 U6839 ( .A1(n5687), .A2(n8840), .ZN(n5423) );
  INV_X1 U6840 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n5421) );
  OR2_X1 U6841 ( .A1(n6712), .A2(n5421), .ZN(n5422) );
  NAND2_X1 U6842 ( .A1(n8842), .A2(n7700), .ZN(n9172) );
  NAND2_X1 U6843 ( .A1(n9014), .A2(n9172), .ZN(n7612) );
  NAND2_X1 U6844 ( .A1(n7613), .A2(n7612), .ZN(n7611) );
  INV_X1 U6845 ( .A(n7700), .ZN(n9255) );
  OR2_X1 U6846 ( .A1(n8842), .A2(n9255), .ZN(n5426) );
  NAND2_X1 U6847 ( .A1(n7611), .A2(n5426), .ZN(n7705) );
  INV_X1 U6848 ( .A(n5428), .ZN(n5429) );
  MUX2_X1 U6849 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n5011), .Z(n5450) );
  XNOR2_X1 U6850 ( .A(n5450), .B(SI_13_), .ZN(n5447) );
  XNOR2_X1 U6851 ( .A(n5449), .B(n5447), .ZN(n6914) );
  NAND2_X1 U6852 ( .A1(n6914), .A2(n5295), .ZN(n5437) );
  INV_X1 U6853 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n5432) );
  NAND2_X1 U6854 ( .A1(n5433), .A2(n5432), .ZN(n5434) );
  NAND2_X1 U6855 ( .A1(n5434), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5435) );
  XNOR2_X1 U6856 ( .A(n5435), .B(P1_IR_REG_13__SCAN_IN), .ZN(n9799) );
  AOI22_X1 U6857 ( .A1(n5560), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n5559), .B2(
        n9799), .ZN(n5436) );
  NAND2_X1 U6858 ( .A1(n5718), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n5445) );
  INV_X1 U6859 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n7551) );
  OR2_X1 U6860 ( .A1(n6712), .A2(n7551), .ZN(n5444) );
  NAND2_X1 U6861 ( .A1(n5438), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n5459) );
  INV_X1 U6862 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n10445) );
  NAND2_X1 U6863 ( .A1(n5439), .A2(n10445), .ZN(n5440) );
  NAND2_X1 U6864 ( .A1(n5459), .A2(n5440), .ZN(n8899) );
  OR2_X1 U6865 ( .A1(n5687), .A2(n8899), .ZN(n5443) );
  INV_X1 U6866 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n5441) );
  OR2_X1 U6867 ( .A1(n5244), .A2(n5441), .ZN(n5442) );
  OR2_X1 U6868 ( .A1(n8901), .A2(n7605), .ZN(n9031) );
  NAND2_X1 U6869 ( .A1(n8901), .A2(n7605), .ZN(n9567) );
  NAND2_X1 U6870 ( .A1(n9031), .A2(n9567), .ZN(n9103) );
  INV_X1 U6871 ( .A(n7605), .ZN(n9254) );
  OR2_X1 U6872 ( .A1(n8901), .A2(n9254), .ZN(n5446) );
  INV_X1 U6873 ( .A(n5447), .ZN(n5448) );
  NAND2_X1 U6874 ( .A1(n5450), .A2(SI_13_), .ZN(n5451) );
  XNOR2_X1 U6875 ( .A(n5469), .B(SI_14_), .ZN(n5466) );
  XNOR2_X1 U6876 ( .A(n5468), .B(n5466), .ZN(n6974) );
  NAND2_X1 U6877 ( .A1(n6974), .A2(n5295), .ZN(n5456) );
  NAND2_X1 U6878 ( .A1(n5453), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5454) );
  XNOR2_X1 U6879 ( .A(n5454), .B(P1_IR_REG_14__SCAN_IN), .ZN(n9811) );
  AOI22_X1 U6880 ( .A1(n5560), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n5559), .B2(
        n9811), .ZN(n5455) );
  INV_X1 U6881 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n5457) );
  OR2_X1 U6882 ( .A1(n6709), .A2(n5457), .ZN(n5464) );
  INV_X1 U6883 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n5458) );
  OR2_X1 U6884 ( .A1(n6712), .A2(n5458), .ZN(n5463) );
  INV_X1 U6885 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n8795) );
  NAND2_X1 U6886 ( .A1(n5459), .A2(n8795), .ZN(n5460) );
  NAND2_X1 U6887 ( .A1(n5477), .A2(n5460), .ZN(n8794) );
  OR2_X1 U6888 ( .A1(n5595), .A2(n8794), .ZN(n5462) );
  INV_X1 U6889 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n10367) );
  OR2_X1 U6890 ( .A1(n5244), .A2(n10367), .ZN(n5461) );
  NAND4_X1 U6891 ( .A1(n5464), .A2(n5463), .A3(n5462), .A4(n5461), .ZN(n9253)
         );
  NAND2_X1 U6892 ( .A1(n9655), .A2(n9253), .ZN(n5465) );
  INV_X1 U6893 ( .A(n5466), .ZN(n5467) );
  NAND2_X1 U6894 ( .A1(n5468), .A2(n5467), .ZN(n5471) );
  NAND2_X1 U6895 ( .A1(n5469), .A2(SI_14_), .ZN(n5470) );
  XNOR2_X1 U6896 ( .A(n5485), .B(SI_15_), .ZN(n5472) );
  XNOR2_X1 U6897 ( .A(n5490), .B(n5472), .ZN(n7038) );
  NAND2_X1 U6898 ( .A1(n7038), .A2(n5295), .ZN(n5475) );
  NAND2_X1 U6899 ( .A1(n4535), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5473) );
  XNOR2_X1 U6900 ( .A(n5473), .B(P1_IR_REG_15__SCAN_IN), .ZN(n9822) );
  AOI22_X1 U6901 ( .A1(n5560), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n5559), .B2(
        n9822), .ZN(n5474) );
  NAND2_X1 U6902 ( .A1(n5731), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n5482) );
  INV_X1 U6903 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n7871) );
  OR2_X1 U6904 ( .A1(n6709), .A2(n7871), .ZN(n5481) );
  INV_X1 U6905 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n9816) );
  OR2_X1 U6906 ( .A1(n6712), .A2(n9816), .ZN(n5480) );
  INV_X1 U6907 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n5476) );
  NAND2_X1 U6908 ( .A1(n5477), .A2(n5476), .ZN(n5478) );
  NAND2_X1 U6909 ( .A1(n5497), .A2(n5478), .ZN(n8956) );
  OR2_X1 U6910 ( .A1(n5687), .A2(n8956), .ZN(n5479) );
  NAND4_X1 U6911 ( .A1(n5482), .A2(n5481), .A3(n5480), .A4(n5479), .ZN(n9252)
         );
  NOR2_X1 U6912 ( .A1(n9025), .A2(n9252), .ZN(n5484) );
  NAND2_X1 U6913 ( .A1(n9025), .A2(n9252), .ZN(n5483) );
  OAI21_X1 U6914 ( .B1(n7870), .B2(n5484), .A(n5483), .ZN(n9545) );
  INV_X1 U6915 ( .A(n5485), .ZN(n5487) );
  INV_X1 U6916 ( .A(SI_15_), .ZN(n5486) );
  NAND2_X1 U6917 ( .A1(n5487), .A2(n5486), .ZN(n5488) );
  MUX2_X1 U6918 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(P2_DATAO_REG_16__SCAN_IN), 
        .S(n5011), .Z(n5505) );
  INV_X1 U6919 ( .A(SI_16_), .ZN(n10417) );
  XNOR2_X1 U6920 ( .A(n5505), .B(n10417), .ZN(n5491) );
  XNOR2_X1 U6921 ( .A(n5506), .B(n5491), .ZN(n7070) );
  NAND2_X1 U6922 ( .A1(n7070), .A2(n5295), .ZN(n5494) );
  NAND2_X1 U6923 ( .A1(n5512), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5492) );
  XNOR2_X1 U6924 ( .A(n5492), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9837) );
  AOI22_X1 U6925 ( .A1(n5560), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n5559), .B2(
        n9837), .ZN(n5493) );
  NAND2_X1 U6926 ( .A1(n5718), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n5502) );
  INV_X1 U6927 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n10430) );
  OR2_X1 U6928 ( .A1(n5244), .A2(n10430), .ZN(n5501) );
  NAND2_X1 U6929 ( .A1(n5495), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n5518) );
  INV_X1 U6930 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n5496) );
  NAND2_X1 U6931 ( .A1(n5497), .A2(n5496), .ZN(n5498) );
  NAND2_X1 U6932 ( .A1(n5518), .A2(n5498), .ZN(n9556) );
  OR2_X1 U6933 ( .A1(n5687), .A2(n9556), .ZN(n5500) );
  INV_X1 U6934 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n10443) );
  OR2_X1 U6935 ( .A1(n6712), .A2(n10443), .ZN(n5499) );
  OR2_X1 U6936 ( .A1(n9555), .A2(n8869), .ZN(n9034) );
  NAND2_X1 U6937 ( .A1(n9555), .A2(n8869), .ZN(n9527) );
  NAND2_X1 U6938 ( .A1(n9034), .A2(n9527), .ZN(n9123) );
  NAND2_X1 U6939 ( .A1(n9545), .A2(n9123), .ZN(n5504) );
  INV_X1 U6940 ( .A(n8869), .ZN(n9251) );
  NAND2_X1 U6941 ( .A1(n9555), .A2(n9251), .ZN(n5503) );
  NAND2_X1 U6942 ( .A1(n5504), .A2(n5503), .ZN(n9534) );
  INV_X1 U6943 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n7211) );
  INV_X1 U6944 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n5507) );
  MUX2_X1 U6945 ( .A(n7211), .B(n5507), .S(n5011), .Z(n5509) );
  INV_X1 U6946 ( .A(SI_17_), .ZN(n5508) );
  NAND2_X1 U6947 ( .A1(n5509), .A2(n5508), .ZN(n5527) );
  INV_X1 U6948 ( .A(n5509), .ZN(n5510) );
  NAND2_X1 U6949 ( .A1(n5510), .A2(SI_17_), .ZN(n5511) );
  NAND2_X1 U6950 ( .A1(n5527), .A2(n5511), .ZN(n5528) );
  XNOR2_X1 U6951 ( .A(n5529), .B(n5528), .ZN(n7159) );
  NAND2_X1 U6952 ( .A1(n7159), .A2(n5295), .ZN(n5515) );
  INV_X1 U6953 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n5513) );
  XNOR2_X1 U6954 ( .A(n5531), .B(P1_IR_REG_17__SCAN_IN), .ZN(n7851) );
  AOI22_X1 U6955 ( .A1(n5560), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n5559), .B2(
        n7851), .ZN(n5514) );
  NAND2_X1 U6956 ( .A1(n5731), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n5523) );
  INV_X1 U6957 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n9539) );
  OR2_X1 U6958 ( .A1(n6709), .A2(n9539), .ZN(n5522) );
  INV_X1 U6959 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n10324) );
  OR2_X1 U6960 ( .A1(n6712), .A2(n10324), .ZN(n5521) );
  INV_X1 U6961 ( .A(n5518), .ZN(n5516) );
  NAND2_X1 U6962 ( .A1(n5516), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n5536) );
  INV_X1 U6963 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n5517) );
  NAND2_X1 U6964 ( .A1(n5518), .A2(n5517), .ZN(n5519) );
  NAND2_X1 U6965 ( .A1(n5536), .A2(n5519), .ZN(n9538) );
  OR2_X1 U6966 ( .A1(n5595), .A2(n9538), .ZN(n5520) );
  NAND4_X1 U6967 ( .A1(n5523), .A2(n5522), .A3(n5521), .A4(n5520), .ZN(n9250)
         );
  OR2_X1 U6968 ( .A1(n9537), .A2(n9250), .ZN(n5524) );
  NAND2_X1 U6969 ( .A1(n9534), .A2(n5524), .ZN(n5526) );
  NAND2_X1 U6970 ( .A1(n9537), .A2(n9250), .ZN(n5525) );
  NAND2_X1 U6971 ( .A1(n5526), .A2(n5525), .ZN(n9510) );
  INV_X1 U6972 ( .A(SI_18_), .ZN(n5530) );
  XNOR2_X1 U6973 ( .A(n5545), .B(n5530), .ZN(n5544) );
  XNOR2_X1 U6974 ( .A(n5548), .B(n5544), .ZN(n7298) );
  NAND2_X1 U6975 ( .A1(n7298), .A2(n5295), .ZN(n5534) );
  INV_X1 U6976 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5741) );
  NAND2_X1 U6977 ( .A1(n5531), .A2(n5741), .ZN(n5532) );
  XNOR2_X1 U6978 ( .A(n5556), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9850) );
  AOI22_X1 U6979 ( .A1(n5560), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n5559), .B2(
        n9850), .ZN(n5533) );
  NAND2_X1 U6980 ( .A1(n5718), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n5541) );
  INV_X1 U6981 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9637) );
  OR2_X1 U6982 ( .A1(n6712), .A2(n9637), .ZN(n5540) );
  INV_X1 U6983 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n5535) );
  NAND2_X1 U6984 ( .A1(n5536), .A2(n5535), .ZN(n5537) );
  NAND2_X1 U6985 ( .A1(n5565), .A2(n5537), .ZN(n9520) );
  OR2_X1 U6986 ( .A1(n5595), .A2(n9520), .ZN(n5539) );
  INV_X1 U6987 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n9701) );
  OR2_X1 U6988 ( .A1(n5244), .A2(n9701), .ZN(n5538) );
  NAND4_X1 U6989 ( .A1(n5541), .A2(n5540), .A3(n5539), .A4(n5538), .ZN(n9249)
         );
  AND2_X1 U6990 ( .A1(n9519), .A2(n9249), .ZN(n5543) );
  OR2_X1 U6991 ( .A1(n9519), .A2(n9249), .ZN(n5542) );
  INV_X1 U6992 ( .A(n9498), .ZN(n5571) );
  NAND2_X1 U6993 ( .A1(n5545), .A2(SI_18_), .ZN(n5546) );
  INV_X1 U6994 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7373) );
  INV_X1 U6995 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7371) );
  MUX2_X1 U6996 ( .A(n7373), .B(n7371), .S(n5011), .Z(n5550) );
  INV_X1 U6997 ( .A(SI_19_), .ZN(n5549) );
  NAND2_X1 U6998 ( .A1(n5550), .A2(n5549), .ZN(n5573) );
  INV_X1 U6999 ( .A(n5550), .ZN(n5551) );
  NAND2_X1 U7000 ( .A1(n5551), .A2(SI_19_), .ZN(n5552) );
  NAND2_X1 U7001 ( .A1(n5573), .A2(n5552), .ZN(n5553) );
  NAND2_X1 U7002 ( .A1(n5554), .A2(n5553), .ZN(n5555) );
  NAND2_X1 U7003 ( .A1(n5574), .A2(n5555), .ZN(n7370) );
  NAND2_X1 U7004 ( .A1(n7370), .A2(n5295), .ZN(n5562) );
  INV_X1 U7005 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n5740) );
  NAND2_X1 U7006 ( .A1(n5556), .A2(n5740), .ZN(n5557) );
  INV_X1 U7007 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5739) );
  XNOR2_X2 U7008 ( .A(n5558), .B(n5739), .ZN(n9230) );
  AOI22_X1 U7009 ( .A1(n5560), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n5559), .B2(
        n4621), .ZN(n5561) );
  NAND2_X1 U7010 ( .A1(n5264), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n5570) );
  INV_X1 U7011 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n9632) );
  OR2_X1 U7012 ( .A1(n6712), .A2(n9632), .ZN(n5569) );
  INV_X1 U7013 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n9504) );
  OR2_X1 U7014 ( .A1(n6709), .A2(n9504), .ZN(n5568) );
  NAND2_X1 U7015 ( .A1(n5563), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n5578) );
  INV_X1 U7016 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n5564) );
  NAND2_X1 U7017 ( .A1(n5565), .A2(n5564), .ZN(n5566) );
  NAND2_X1 U7018 ( .A1(n5578), .A2(n5566), .ZN(n9503) );
  OR2_X1 U7019 ( .A1(n5687), .A2(n9503), .ZN(n5567) );
  NAND4_X1 U7020 ( .A1(n5570), .A2(n5569), .A3(n5568), .A4(n5567), .ZN(n9248)
         );
  NAND2_X1 U7021 ( .A1(n9502), .A2(n9248), .ZN(n5572) );
  INV_X1 U7022 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7512) );
  INV_X1 U7023 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7515) );
  XNOR2_X1 U7024 ( .A(n5585), .B(SI_20_), .ZN(n5575) );
  XNOR2_X1 U7025 ( .A(n5587), .B(n5575), .ZN(n7511) );
  NAND2_X1 U7026 ( .A1(n7511), .A2(n5295), .ZN(n5577) );
  OR2_X1 U7027 ( .A1(n5234), .A2(n7515), .ZN(n5576) );
  INV_X1 U7028 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n8890) );
  NAND2_X1 U7029 ( .A1(n5578), .A2(n8890), .ZN(n5579) );
  NAND2_X1 U7030 ( .A1(n5593), .A2(n5579), .ZN(n9486) );
  NAND2_X1 U7031 ( .A1(n5731), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n5580) );
  OAI21_X1 U7032 ( .B1(n9486), .B2(n5595), .A(n5580), .ZN(n5582) );
  INV_X1 U7033 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n10371) );
  INV_X1 U7034 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n9487) );
  OAI22_X1 U7035 ( .A1(n6712), .A2(n10371), .B1(n6709), .B2(n9487), .ZN(n5581)
         );
  OR2_X1 U7036 ( .A1(n5582), .A2(n5581), .ZN(n9247) );
  AND2_X1 U7037 ( .A1(n9485), .A2(n9247), .ZN(n5584) );
  INV_X1 U7038 ( .A(SI_20_), .ZN(n5586) );
  INV_X1 U7039 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7528) );
  INV_X1 U7040 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7532) );
  MUX2_X1 U7041 ( .A(n7528), .B(n7532), .S(n5011), .Z(n5601) );
  XNOR2_X1 U7042 ( .A(n5601), .B(SI_21_), .ZN(n5588) );
  XNOR2_X1 U7043 ( .A(n5603), .B(n5588), .ZN(n7527) );
  NAND2_X1 U7044 ( .A1(n7527), .A2(n5295), .ZN(n5590) );
  OR2_X1 U7045 ( .A1(n5234), .A2(n7532), .ZN(n5589) );
  INV_X1 U7046 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n10446) );
  NAND2_X1 U7047 ( .A1(n5591), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n5610) );
  INV_X1 U7048 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n5592) );
  NAND2_X1 U7049 ( .A1(n5593), .A2(n5592), .ZN(n5594) );
  NAND2_X1 U7050 ( .A1(n5610), .A2(n5594), .ZN(n9471) );
  OR2_X1 U7051 ( .A1(n9471), .A2(n5595), .ZN(n5598) );
  AOI22_X1 U7052 ( .A1(n5732), .A2(P1_REG1_REG_21__SCAN_IN), .B1(n5718), .B2(
        P1_REG2_REG_21__SCAN_IN), .ZN(n5597) );
  OAI211_X1 U7053 ( .C1(n5244), .C2(n10446), .A(n5598), .B(n5597), .ZN(n9246)
         );
  NAND2_X1 U7054 ( .A1(n9470), .A2(n9246), .ZN(n5599) );
  NAND2_X1 U7055 ( .A1(n5600), .A2(n5599), .ZN(n9449) );
  INV_X1 U7056 ( .A(n5601), .ZN(n5602) );
  INV_X1 U7057 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7690) );
  INV_X1 U7058 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7687) );
  INV_X1 U7059 ( .A(SI_22_), .ZN(n5604) );
  NAND2_X1 U7060 ( .A1(n5605), .A2(n5604), .ZN(n5616) );
  INV_X1 U7061 ( .A(n5605), .ZN(n5606) );
  NAND2_X1 U7062 ( .A1(n5606), .A2(SI_22_), .ZN(n5607) );
  NAND2_X1 U7063 ( .A1(n5616), .A2(n5607), .ZN(n5617) );
  XNOR2_X1 U7064 ( .A(n5618), .B(n5617), .ZN(n7686) );
  NAND2_X1 U7065 ( .A1(n7686), .A2(n5295), .ZN(n5609) );
  OR2_X1 U7066 ( .A1(n5234), .A2(n7687), .ZN(n5608) );
  INV_X1 U7067 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n8911) );
  NAND2_X1 U7068 ( .A1(n5610), .A2(n8911), .ZN(n5611) );
  NAND2_X1 U7069 ( .A1(n5630), .A2(n5611), .ZN(n9452) );
  AOI22_X1 U7070 ( .A1(n5732), .A2(P1_REG1_REG_22__SCAN_IN), .B1(n5718), .B2(
        P1_REG2_REG_22__SCAN_IN), .ZN(n5613) );
  NAND2_X1 U7071 ( .A1(n5731), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n5612) );
  OAI211_X1 U7072 ( .C1(n9452), .C2(n5687), .A(n5613), .B(n5612), .ZN(n9245)
         );
  AND2_X1 U7073 ( .A1(n9451), .A2(n9245), .ZN(n5615) );
  OR2_X1 U7074 ( .A1(n9451), .A2(n9245), .ZN(n5614) );
  INV_X1 U7075 ( .A(n5626), .ZN(n5623) );
  INV_X1 U7076 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n7748) );
  INV_X1 U7077 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n7752) );
  MUX2_X1 U7078 ( .A(n7748), .B(n7752), .S(n5011), .Z(n5620) );
  INV_X1 U7079 ( .A(SI_23_), .ZN(n5619) );
  NAND2_X1 U7080 ( .A1(n5620), .A2(n5619), .ZN(n5637) );
  INV_X1 U7081 ( .A(n5620), .ZN(n5621) );
  NAND2_X1 U7082 ( .A1(n5621), .A2(SI_23_), .ZN(n5622) );
  NAND2_X1 U7083 ( .A1(n5637), .A2(n5622), .ZN(n5624) );
  NAND2_X1 U7084 ( .A1(n5623), .A2(n5624), .ZN(n5627) );
  INV_X1 U7085 ( .A(n5624), .ZN(n5625) );
  NAND2_X1 U7086 ( .A1(n5627), .A2(n5638), .ZN(n7750) );
  NAND2_X1 U7087 ( .A1(n7750), .A2(n5295), .ZN(n5629) );
  OR2_X1 U7088 ( .A1(n5234), .A2(n7752), .ZN(n5628) );
  INV_X1 U7089 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n8803) );
  NAND2_X1 U7090 ( .A1(n5630), .A2(n8803), .ZN(n5631) );
  NAND2_X1 U7091 ( .A1(n5666), .A2(n5631), .ZN(n9436) );
  INV_X1 U7092 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n9613) );
  NAND2_X1 U7093 ( .A1(n5718), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n5633) );
  NAND2_X1 U7094 ( .A1(n5264), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n5632) );
  OAI211_X1 U7095 ( .C1(n6712), .C2(n9613), .A(n5633), .B(n5632), .ZN(n5634)
         );
  INV_X1 U7096 ( .A(n5634), .ZN(n5635) );
  OAI21_X1 U7097 ( .B1(n9436), .B2(n5687), .A(n5635), .ZN(n9244) );
  NOR2_X1 U7098 ( .A1(n9435), .A2(n9244), .ZN(n5636) );
  INV_X1 U7099 ( .A(n5645), .ZN(n5642) );
  INV_X1 U7100 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n6204) );
  INV_X1 U7101 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n5647) );
  INV_X1 U7102 ( .A(SI_24_), .ZN(n10428) );
  NAND2_X1 U7103 ( .A1(n5639), .A2(n10428), .ZN(n5655) );
  INV_X1 U7104 ( .A(n5639), .ZN(n5640) );
  NAND2_X1 U7105 ( .A1(n5640), .A2(SI_24_), .ZN(n5641) );
  NAND2_X1 U7106 ( .A1(n5655), .A2(n5641), .ZN(n5643) );
  NAND2_X1 U7107 ( .A1(n5642), .A2(n5643), .ZN(n5646) );
  INV_X1 U7108 ( .A(n5643), .ZN(n5644) );
  NAND2_X1 U7109 ( .A1(n5646), .A2(n5656), .ZN(n7906) );
  NAND2_X1 U7110 ( .A1(n7906), .A2(n5295), .ZN(n5649) );
  OR2_X1 U7111 ( .A1(n5234), .A2(n5647), .ZN(n5648) );
  XNOR2_X1 U7112 ( .A(n5666), .B(P1_REG3_REG_24__SCAN_IN), .ZN(n9416) );
  INV_X1 U7113 ( .A(n5595), .ZN(n5736) );
  NAND2_X1 U7114 ( .A1(n9416), .A2(n5736), .ZN(n5654) );
  INV_X1 U7115 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n10416) );
  NAND2_X1 U7116 ( .A1(n5718), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n5651) );
  NAND2_X1 U7117 ( .A1(n5264), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n5650) );
  OAI211_X1 U7118 ( .C1(n6712), .C2(n10416), .A(n5651), .B(n5650), .ZN(n5652)
         );
  INV_X1 U7119 ( .A(n5652), .ZN(n5653) );
  NAND2_X1 U7120 ( .A1(n5654), .A2(n5653), .ZN(n8847) );
  INV_X1 U7121 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n8785) );
  INV_X1 U7122 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n9736) );
  MUX2_X1 U7123 ( .A(n8785), .B(n9736), .S(n5011), .Z(n5658) );
  INV_X1 U7124 ( .A(SI_25_), .ZN(n5657) );
  NAND2_X1 U7125 ( .A1(n5658), .A2(n5657), .ZN(n5677) );
  INV_X1 U7126 ( .A(n5658), .ZN(n5659) );
  NAND2_X1 U7127 ( .A1(n5659), .A2(SI_25_), .ZN(n5660) );
  AND2_X1 U7128 ( .A1(n5677), .A2(n5660), .ZN(n5675) );
  OR2_X1 U7129 ( .A1(n5234), .A2(n9736), .ZN(n5661) );
  INV_X1 U7130 ( .A(n5666), .ZN(n5664) );
  AND2_X1 U7131 ( .A1(P1_REG3_REG_24__SCAN_IN), .A2(P1_REG3_REG_25__SCAN_IN), 
        .ZN(n5663) );
  NAND2_X1 U7132 ( .A1(n5664), .A2(n5663), .ZN(n5685) );
  INV_X1 U7133 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n8881) );
  INV_X1 U7134 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n5665) );
  OAI21_X1 U7135 ( .B1(n5666), .B2(n8881), .A(n5665), .ZN(n5667) );
  AND2_X1 U7136 ( .A1(n5685), .A2(n5667), .ZN(n9405) );
  NAND2_X1 U7137 ( .A1(n9405), .A2(n5736), .ZN(n5672) );
  INV_X1 U7138 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n9604) );
  NAND2_X1 U7139 ( .A1(n5718), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n5669) );
  NAND2_X1 U7140 ( .A1(n5264), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n5668) );
  OAI211_X1 U7141 ( .C1(n6712), .C2(n9604), .A(n5669), .B(n5668), .ZN(n5670)
         );
  INV_X1 U7142 ( .A(n5670), .ZN(n5671) );
  NAND2_X1 U7143 ( .A1(n5672), .A2(n5671), .ZN(n9243) );
  NOR2_X1 U7144 ( .A1(n9404), .A2(n9243), .ZN(n5674) );
  NAND2_X1 U7145 ( .A1(n9404), .A2(n9243), .ZN(n5673) );
  INV_X1 U7146 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n8782) );
  INV_X1 U7147 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n9732) );
  INV_X1 U7148 ( .A(SI_26_), .ZN(n5678) );
  NAND2_X1 U7149 ( .A1(n5679), .A2(n5678), .ZN(n5697) );
  INV_X1 U7150 ( .A(n5679), .ZN(n5680) );
  NAND2_X1 U7151 ( .A1(n5680), .A2(SI_26_), .ZN(n5681) );
  AND2_X1 U7152 ( .A1(n5697), .A2(n5681), .ZN(n5695) );
  NAND2_X1 U7153 ( .A1(n8781), .A2(n5295), .ZN(n5683) );
  OR2_X1 U7154 ( .A1(n5234), .A2(n9732), .ZN(n5682) );
  INV_X1 U7155 ( .A(n5685), .ZN(n5684) );
  NAND2_X1 U7156 ( .A1(n5684), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n5716) );
  INV_X1 U7157 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n10348) );
  NAND2_X1 U7158 ( .A1(n5685), .A2(n10348), .ZN(n5686) );
  NAND2_X1 U7159 ( .A1(n5716), .A2(n5686), .ZN(n9388) );
  OR2_X1 U7160 ( .A1(n9388), .A2(n5687), .ZN(n5692) );
  INV_X1 U7161 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n9599) );
  NAND2_X1 U7162 ( .A1(n5718), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n5689) );
  NAND2_X1 U7163 ( .A1(n5264), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n5688) );
  OAI211_X1 U7164 ( .C1(n9599), .C2(n6712), .A(n5689), .B(n5688), .ZN(n5690)
         );
  INV_X1 U7165 ( .A(n5690), .ZN(n5691) );
  NAND2_X1 U7166 ( .A1(n9382), .A2(n9384), .ZN(n5694) );
  NAND2_X1 U7167 ( .A1(n9392), .A2(n9242), .ZN(n5693) );
  INV_X1 U7168 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n8778) );
  INV_X1 U7169 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n8164) );
  MUX2_X1 U7170 ( .A(n8778), .B(n8164), .S(n5011), .Z(n5700) );
  INV_X1 U7171 ( .A(SI_27_), .ZN(n5699) );
  NAND2_X1 U7172 ( .A1(n5700), .A2(n5699), .ZN(n5711) );
  INV_X1 U7173 ( .A(n5700), .ZN(n5701) );
  NAND2_X1 U7174 ( .A1(n5701), .A2(SI_27_), .ZN(n5702) );
  AND2_X1 U7175 ( .A1(n5711), .A2(n5702), .ZN(n5709) );
  NAND2_X1 U7176 ( .A1(n8162), .A2(n5295), .ZN(n5704) );
  OR2_X1 U7177 ( .A1(n5234), .A2(n8164), .ZN(n5703) );
  XNOR2_X1 U7178 ( .A(n5716), .B(P1_REG3_REG_27__SCAN_IN), .ZN(n9376) );
  INV_X1 U7179 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n9594) );
  NAND2_X1 U7180 ( .A1(n5718), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n5706) );
  NAND2_X1 U7181 ( .A1(n5731), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n5705) );
  OAI211_X1 U7182 ( .C1(n9594), .C2(n6712), .A(n5706), .B(n5705), .ZN(n5707)
         );
  AOI21_X1 U7183 ( .B1(n9376), .B2(n5736), .A(n5707), .ZN(n8947) );
  NAND2_X1 U7184 ( .A1(n9375), .A2(n8947), .ZN(n9072) );
  INV_X1 U7185 ( .A(n8947), .ZN(n9241) );
  INV_X1 U7186 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n8777) );
  INV_X1 U7187 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n9731) );
  XNOR2_X1 U7188 ( .A(n5726), .B(SI_28_), .ZN(n5723) );
  NAND2_X1 U7189 ( .A1(n9728), .A2(n5295), .ZN(n5713) );
  OR2_X1 U7190 ( .A1(n5234), .A2(n9731), .ZN(n5712) );
  INV_X1 U7191 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n6134) );
  INV_X1 U7192 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n5714) );
  OAI21_X1 U7193 ( .B1(n5716), .B2(n6134), .A(n5714), .ZN(n5717) );
  NAND2_X1 U7194 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(P1_REG3_REG_28__SCAN_IN), 
        .ZN(n5715) );
  OR2_X1 U7195 ( .A1(n5716), .A2(n5715), .ZN(n9347) );
  INV_X1 U7196 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n6124) );
  NAND2_X1 U7197 ( .A1(n5718), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n5720) );
  NAND2_X1 U7198 ( .A1(n5731), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n5719) );
  OAI211_X1 U7199 ( .C1(n6712), .C2(n6124), .A(n5720), .B(n5719), .ZN(n5721)
         );
  AOI21_X1 U7200 ( .B1(n9358), .B2(n5736), .A(n5721), .ZN(n7024) );
  NAND2_X1 U7201 ( .A1(n6119), .A2(n7024), .ZN(n9073) );
  INV_X1 U7202 ( .A(SI_28_), .ZN(n5725) );
  NAND2_X1 U7203 ( .A1(n5726), .A2(n5725), .ZN(n5727) );
  INV_X1 U7204 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n9727) );
  INV_X1 U7205 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n8160) );
  MUX2_X1 U7206 ( .A(n9727), .B(n8160), .S(n7936), .Z(n7928) );
  NAND2_X1 U7207 ( .A1(n8159), .A2(n5295), .ZN(n5730) );
  OR2_X1 U7208 ( .A1(n5234), .A2(n9727), .ZN(n5729) );
  INV_X1 U7209 ( .A(n9347), .ZN(n5737) );
  INV_X1 U7210 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n9346) );
  NAND2_X1 U7211 ( .A1(n5731), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n5734) );
  NAND2_X1 U7212 ( .A1(n5732), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n5733) );
  OAI211_X1 U7213 ( .C1(n6709), .C2(n9346), .A(n5734), .B(n5733), .ZN(n5735)
         );
  AOI21_X1 U7214 ( .B1(n5737), .B2(n5736), .A(n5735), .ZN(n6939) );
  NAND2_X1 U7215 ( .A1(n9349), .A2(n6939), .ZN(n9200) );
  XNOR2_X1 U7216 ( .A(n5738), .B(n4740), .ZN(n9345) );
  NAND3_X1 U7217 ( .A1(n5741), .A2(n5740), .A3(n5739), .ZN(n5742) );
  NOR2_X2 U7218 ( .A1(n5743), .A2(n5742), .ZN(n5749) );
  INV_X1 U7219 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5744) );
  NAND2_X1 U7220 ( .A1(n5749), .A2(n5744), .ZN(n5752) );
  INV_X1 U7221 ( .A(n5752), .ZN(n5746) );
  INV_X1 U7222 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5745) );
  NAND2_X1 U7223 ( .A1(n5746), .A2(n5745), .ZN(n5800) );
  NAND2_X1 U7224 ( .A1(n5800), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5747) );
  INV_X1 U7225 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5798) );
  NAND2_X1 U7226 ( .A1(n5747), .A2(n5798), .ZN(n5807) );
  OR2_X1 U7227 ( .A1(n5747), .A2(n5798), .ZN(n5748) );
  INV_X1 U7228 ( .A(n5749), .ZN(n5750) );
  NAND2_X1 U7229 ( .A1(n5750), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5751) );
  MUX2_X1 U7230 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5751), .S(
        P1_IR_REG_20__SCAN_IN), .Z(n5753) );
  NAND2_X1 U7231 ( .A1(n5753), .A2(n5752), .ZN(n9223) );
  AND2_X2 U7232 ( .A1(n9223), .A2(n9230), .ZN(n9233) );
  INV_X1 U7233 ( .A(n9233), .ZN(n5827) );
  NAND2_X1 U7234 ( .A1(n5836), .A2(n5827), .ZN(n5755) );
  XNOR2_X2 U7235 ( .A(n5754), .B(P1_IR_REG_21__SCAN_IN), .ZN(n9150) );
  INV_X1 U7236 ( .A(n9150), .ZN(n7530) );
  INV_X1 U7237 ( .A(n6088), .ZN(n7132) );
  AND2_X1 U7238 ( .A1(n5755), .A2(n7132), .ZN(n5756) );
  NAND2_X1 U7239 ( .A1(n9236), .A2(n9150), .ZN(n9219) );
  NAND2_X1 U7240 ( .A1(n6698), .A2(n9233), .ZN(n7131) );
  NAND2_X1 U7241 ( .A1(n5756), .A2(n7131), .ZN(n9564) );
  NAND2_X1 U7242 ( .A1(n9096), .A2(n9223), .ZN(n9659) );
  INV_X1 U7243 ( .A(n5757), .ZN(n6923) );
  NAND2_X1 U7244 ( .A1(n6698), .A2(n6923), .ZN(n8944) );
  INV_X1 U7245 ( .A(n8163), .ZN(n9774) );
  NAND2_X1 U7246 ( .A1(n9774), .A2(P1_B_REG_SCAN_IN), .ZN(n5758) );
  NAND2_X1 U7247 ( .A1(n8932), .A2(n5758), .ZN(n9333) );
  INV_X1 U7248 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n5759) );
  OR2_X1 U7249 ( .A1(n6712), .A2(n5759), .ZN(n5763) );
  INV_X1 U7250 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n9341) );
  OR2_X1 U7251 ( .A1(n6709), .A2(n9341), .ZN(n5762) );
  INV_X1 U7252 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n5760) );
  OR2_X1 U7253 ( .A1(n5244), .A2(n5760), .ZN(n5761) );
  AND3_X1 U7254 ( .A1(n5763), .A2(n5762), .A3(n5761), .ZN(n9101) );
  NAND2_X1 U7255 ( .A1(n9236), .A2(n4621), .ZN(n5764) );
  NAND2_X1 U7256 ( .A1(n9224), .A2(n9150), .ZN(n9097) );
  INV_X1 U7257 ( .A(n6976), .ZN(n7138) );
  NOR2_X1 U7258 ( .A1(n7074), .A2(n7138), .ZN(n7075) );
  NAND2_X1 U7259 ( .A1(n7059), .A2(n7075), .ZN(n7061) );
  INV_X1 U7260 ( .A(n9865), .ZN(n8974) );
  NAND2_X1 U7261 ( .A1(n9263), .A2(n8974), .ZN(n8980) );
  NAND2_X1 U7262 ( .A1(n7152), .A2(n8980), .ZN(n5766) );
  OR2_X1 U7263 ( .A1(n9263), .A2(n8974), .ZN(n8986) );
  NAND2_X1 U7264 ( .A1(n5766), .A2(n8986), .ZN(n7214) );
  NAND2_X1 U7265 ( .A1(n7214), .A2(n9111), .ZN(n5767) );
  INV_X1 U7266 ( .A(n9113), .ZN(n9159) );
  NAND2_X1 U7267 ( .A1(n9008), .A2(n8995), .ZN(n9001) );
  NAND2_X1 U7268 ( .A1(n8994), .A2(n8992), .ZN(n5768) );
  NOR2_X1 U7269 ( .A1(n9001), .A2(n5768), .ZN(n9164) );
  AND2_X1 U7270 ( .A1(n8999), .A2(n7466), .ZN(n8987) );
  OR2_X1 U7271 ( .A1(n8987), .A2(n9001), .ZN(n5769) );
  AND2_X1 U7272 ( .A1(n5769), .A2(n9004), .ZN(n9166) );
  INV_X1 U7273 ( .A(n9115), .ZN(n7483) );
  NAND2_X1 U7274 ( .A1(n7482), .A2(n7483), .ZN(n7481) );
  NAND2_X1 U7275 ( .A1(n7481), .A2(n9010), .ZN(n7632) );
  INV_X1 U7276 ( .A(n7612), .ZN(n5770) );
  INV_X1 U7277 ( .A(n9253), .ZN(n5771) );
  OR2_X1 U7278 ( .A1(n9655), .A2(n5771), .ZN(n9020) );
  NAND2_X1 U7279 ( .A1(n9655), .A2(n5771), .ZN(n9021) );
  NAND2_X1 U7280 ( .A1(n9020), .A2(n9021), .ZN(n9573) );
  INV_X1 U7281 ( .A(n9567), .ZN(n5772) );
  NOR2_X1 U7282 ( .A1(n9573), .A2(n5772), .ZN(n9036) );
  NAND2_X1 U7283 ( .A1(n9568), .A2(n9036), .ZN(n9569) );
  INV_X1 U7284 ( .A(n9252), .ZN(n5773) );
  OR2_X1 U7285 ( .A1(n9025), .A2(n5773), .ZN(n9033) );
  NAND2_X1 U7286 ( .A1(n9025), .A2(n5773), .ZN(n9022) );
  NAND2_X1 U7287 ( .A1(n9033), .A2(n9022), .ZN(n9121) );
  INV_X1 U7288 ( .A(n9020), .ZN(n9035) );
  NOR2_X1 U7289 ( .A1(n9121), .A2(n9035), .ZN(n5774) );
  NAND2_X1 U7290 ( .A1(n9569), .A2(n5774), .ZN(n5775) );
  NAND2_X1 U7291 ( .A1(n5775), .A2(n9022), .ZN(n9547) );
  INV_X1 U7292 ( .A(n9123), .ZN(n9548) );
  INV_X1 U7293 ( .A(n9250), .ZN(n5776) );
  OR2_X1 U7294 ( .A1(n9537), .A2(n5776), .ZN(n9511) );
  NAND2_X1 U7295 ( .A1(n9537), .A2(n5776), .ZN(n9042) );
  NAND2_X1 U7296 ( .A1(n9511), .A2(n9042), .ZN(n9533) );
  INV_X1 U7297 ( .A(n9527), .ZN(n9023) );
  NOR2_X1 U7298 ( .A1(n9533), .A2(n9023), .ZN(n5777) );
  NAND2_X1 U7299 ( .A1(n9546), .A2(n5777), .ZN(n9528) );
  INV_X1 U7300 ( .A(n9249), .ZN(n5778) );
  OR2_X1 U7301 ( .A1(n9519), .A2(n5778), .ZN(n9046) );
  NAND2_X1 U7302 ( .A1(n9519), .A2(n5778), .ZN(n9047) );
  NAND2_X1 U7303 ( .A1(n9046), .A2(n9047), .ZN(n9513) );
  INV_X1 U7304 ( .A(n9511), .ZN(n5779) );
  NOR2_X1 U7305 ( .A1(n9513), .A2(n5779), .ZN(n5780) );
  NAND2_X1 U7306 ( .A1(n9528), .A2(n5780), .ZN(n5781) );
  NAND2_X1 U7307 ( .A1(n5781), .A2(n9047), .ZN(n9493) );
  INV_X1 U7308 ( .A(n9248), .ZN(n5782) );
  OR2_X1 U7309 ( .A1(n9502), .A2(n5782), .ZN(n9053) );
  NAND2_X1 U7310 ( .A1(n9502), .A2(n5782), .ZN(n9182) );
  NAND2_X1 U7311 ( .A1(n9493), .A2(n9497), .ZN(n5783) );
  INV_X1 U7312 ( .A(n9246), .ZN(n9128) );
  OR2_X1 U7313 ( .A1(n9470), .A2(n9128), .ZN(n9060) );
  INV_X1 U7314 ( .A(n9247), .ZN(n9102) );
  OR2_X1 U7315 ( .A1(n9485), .A2(n9102), .ZN(n9460) );
  AND2_X1 U7316 ( .A1(n9060), .A2(n9460), .ZN(n9146) );
  NAND2_X1 U7317 ( .A1(n9479), .A2(n9146), .ZN(n5785) );
  AND2_X1 U7318 ( .A1(n9485), .A2(n9102), .ZN(n9054) );
  NAND2_X1 U7319 ( .A1(n9060), .A2(n9054), .ZN(n5784) );
  NAND2_X1 U7320 ( .A1(n9470), .A2(n9128), .ZN(n9061) );
  AND2_X1 U7321 ( .A1(n5784), .A2(n9061), .ZN(n9186) );
  INV_X1 U7322 ( .A(n9245), .ZN(n5786) );
  OR2_X1 U7323 ( .A1(n9451), .A2(n5786), .ZN(n9427) );
  NAND2_X1 U7324 ( .A1(n9451), .A2(n5786), .ZN(n9063) );
  NAND2_X1 U7325 ( .A1(n9427), .A2(n9063), .ZN(n9448) );
  INV_X1 U7326 ( .A(n9244), .ZN(n5787) );
  OR2_X1 U7327 ( .A1(n9435), .A2(n5787), .ZN(n9064) );
  NAND2_X1 U7328 ( .A1(n9435), .A2(n5787), .ZN(n9065) );
  INV_X1 U7329 ( .A(n8847), .ZN(n5788) );
  OR2_X1 U7330 ( .A1(n9420), .A2(n5788), .ZN(n9142) );
  NAND2_X1 U7331 ( .A1(n9420), .A2(n5788), .ZN(n9188) );
  NAND2_X1 U7332 ( .A1(n9413), .A2(n9412), .ZN(n5789) );
  NAND2_X1 U7333 ( .A1(n5789), .A2(n9142), .ZN(n9400) );
  INV_X1 U7334 ( .A(n9243), .ZN(n8945) );
  NAND2_X1 U7335 ( .A1(n9404), .A2(n8945), .ZN(n9189) );
  INV_X1 U7336 ( .A(n9072), .ZN(n5790) );
  INV_X1 U7337 ( .A(n9080), .ZN(n9197) );
  INV_X1 U7338 ( .A(n9435), .ZN(n9686) );
  OR2_X1 U7339 ( .A1(n6958), .A2(n6976), .ZN(n7105) );
  NAND2_X1 U7340 ( .A1(n7278), .A2(n9893), .ZN(n7277) );
  OR2_X1 U7341 ( .A1(n7277), .A2(n9865), .ZN(n7218) );
  INV_X1 U7342 ( .A(n7538), .ZN(n9767) );
  INV_X1 U7343 ( .A(n4622), .ZN(n7733) );
  NAND2_X1 U7344 ( .A1(n7639), .A2(n7733), .ZN(n7640) );
  INV_X1 U7345 ( .A(n9025), .ZN(n9714) );
  INV_X1 U7346 ( .A(n9519), .ZN(n9703) );
  INV_X1 U7347 ( .A(n9502), .ZN(n9699) );
  AOI21_X1 U7348 ( .B1(n9349), .B2(n6120), .A(n9578), .ZN(n5793) );
  NAND2_X1 U7349 ( .A1(n4579), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5797) );
  XNOR2_X1 U7350 ( .A(n5797), .B(n5161), .ZN(n9739) );
  NAND2_X1 U7351 ( .A1(n9739), .A2(P1_B_REG_SCAN_IN), .ZN(n5802) );
  INV_X1 U7352 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n5808) );
  NAND2_X1 U7353 ( .A1(n5798), .A2(n5808), .ZN(n5799) );
  OAI21_X2 U7354 ( .B1(n5800), .B2(n5799), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n5801) );
  XNOR2_X2 U7355 ( .A(n5801), .B(P1_IR_REG_24__SCAN_IN), .ZN(n5823) );
  MUX2_X1 U7356 ( .A(n5802), .B(P1_B_REG_SCAN_IN), .S(n5823), .Z(n5805) );
  NAND2_X1 U7357 ( .A1(n5803), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5804) );
  XNOR2_X1 U7358 ( .A(n5804), .B(P1_IR_REG_26__SCAN_IN), .ZN(n5806) );
  NAND2_X1 U7359 ( .A1(n5805), .A2(n5806), .ZN(n9716) );
  NAND2_X1 U7360 ( .A1(n9734), .A2(n9739), .ZN(n9718) );
  OAI21_X1 U7361 ( .B1(n9716), .B2(P1_D_REG_1__SCAN_IN), .A(n9718), .ZN(n5822)
         );
  NAND2_X1 U7362 ( .A1(n5807), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5809) );
  XNOR2_X1 U7363 ( .A(n5809), .B(n5808), .ZN(n6700) );
  NAND2_X2 U7364 ( .A1(n5823), .A2(n5810), .ZN(n6657) );
  OAI211_X1 U7365 ( .C1(n9219), .C2(n9233), .A(n6700), .B(n6657), .ZN(n6097)
         );
  NOR2_X1 U7366 ( .A1(n6097), .A2(P1_U3086), .ZN(n7100) );
  NOR4_X1 U7367 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_17__SCAN_IN), .A3(
        P1_D_REG_18__SCAN_IN), .A4(P1_D_REG_19__SCAN_IN), .ZN(n5814) );
  NOR4_X1 U7368 ( .A1(P1_D_REG_14__SCAN_IN), .A2(P1_D_REG_12__SCAN_IN), .A3(
        P1_D_REG_13__SCAN_IN), .A4(P1_D_REG_15__SCAN_IN), .ZN(n5813) );
  NOR4_X1 U7369 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n5812) );
  NOR4_X1 U7370 ( .A1(P1_D_REG_20__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n5811) );
  NAND4_X1 U7371 ( .A1(n5814), .A2(n5813), .A3(n5812), .A4(n5811), .ZN(n5820)
         );
  NOR2_X1 U7372 ( .A1(P1_D_REG_8__SCAN_IN), .A2(P1_D_REG_21__SCAN_IN), .ZN(
        n5818) );
  NOR4_X1 U7373 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_23__SCAN_IN), .ZN(n5817) );
  NOR4_X1 U7374 ( .A1(P1_D_REG_7__SCAN_IN), .A2(P1_D_REG_9__SCAN_IN), .A3(
        P1_D_REG_10__SCAN_IN), .A4(P1_D_REG_11__SCAN_IN), .ZN(n5816) );
  NOR4_X1 U7375 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        P1_D_REG_5__SCAN_IN), .A4(P1_D_REG_6__SCAN_IN), .ZN(n5815) );
  NAND4_X1 U7376 ( .A1(n5818), .A2(n5817), .A3(n5816), .A4(n5815), .ZN(n5819)
         );
  NOR2_X1 U7377 ( .A1(n5820), .A2(n5819), .ZN(n6082) );
  OR2_X1 U7378 ( .A1(n9716), .A2(n6082), .ZN(n5821) );
  NAND2_X1 U7379 ( .A1(n7872), .A2(n4621), .ZN(n6095) );
  NAND4_X1 U7380 ( .A1(n5822), .A2(n7100), .A3(n5821), .A4(n6095), .ZN(n6123)
         );
  OR2_X1 U7381 ( .A1(n9716), .A2(P1_D_REG_0__SCAN_IN), .ZN(n5825) );
  NAND2_X1 U7382 ( .A1(n5824), .A2(n9734), .ZN(n9719) );
  NAND2_X1 U7383 ( .A1(n5825), .A2(n9719), .ZN(n7099) );
  INV_X1 U7384 ( .A(n7099), .ZN(n5826) );
  INV_X2 U7385 ( .A(n9910), .ZN(n9911) );
  INV_X1 U7386 ( .A(n9349), .ZN(n6635) );
  AND2_X1 U7387 ( .A1(n5827), .A2(n6088), .ZN(n9656) );
  NOR2_X1 U7388 ( .A1(n6635), .A2(n9713), .ZN(n5828) );
  INV_X1 U7389 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n5829) );
  NOR2_X1 U7390 ( .A1(n9911), .A2(n5829), .ZN(n5830) );
  NOR2_X1 U7391 ( .A1(n5828), .A2(n5830), .ZN(n5831) );
  OAI21_X1 U7392 ( .B1(n6640), .B2(n9910), .A(n5831), .ZN(P1_U3519) );
  NAND2_X1 U7393 ( .A1(n5832), .A2(n4513), .ZN(n5838) );
  NAND2_X1 U7394 ( .A1(n9099), .A2(n9233), .ZN(n5834) );
  NAND2_X1 U7395 ( .A1(n5861), .A2(n6958), .ZN(n5837) );
  NAND2_X1 U7396 ( .A1(n5838), .A2(n5837), .ZN(n5839) );
  INV_X2 U7397 ( .A(n5850), .ZN(n6075) );
  XNOR2_X1 U7398 ( .A(n5839), .B(n6075), .ZN(n5842) );
  NAND2_X1 U7399 ( .A1(n5842), .A2(n5841), .ZN(n7026) );
  NAND2_X1 U7400 ( .A1(n7074), .A2(n4514), .ZN(n5846) );
  INV_X1 U7401 ( .A(n6657), .ZN(n5847) );
  AOI22_X1 U7402 ( .A1(n5861), .A2(n6976), .B1(n5847), .B2(
        P1_REG1_REG_0__SCAN_IN), .ZN(n5845) );
  NAND2_X1 U7403 ( .A1(n5846), .A2(n5845), .ZN(n6920) );
  NAND2_X1 U7404 ( .A1(n7074), .A2(n4508), .ZN(n5849) );
  AOI22_X1 U7405 ( .A1(n6976), .A2(n6071), .B1(P1_IR_REG_0__SCAN_IN), .B2(
        n5847), .ZN(n5848) );
  NAND2_X1 U7406 ( .A1(n5849), .A2(n5848), .ZN(n6919) );
  NOR2_X1 U7407 ( .A1(n6976), .A2(n6066), .ZN(n5851) );
  AOI21_X1 U7408 ( .B1(n6920), .B2(n6919), .A(n5851), .ZN(n6954) );
  NAND2_X1 U7409 ( .A1(n7025), .A2(n7026), .ZN(n5859) );
  NAND2_X1 U7410 ( .A1(n5852), .A2(n6071), .ZN(n5854) );
  OR2_X1 U7411 ( .A1(n9888), .A2(n5895), .ZN(n5853) );
  NAND2_X1 U7412 ( .A1(n5854), .A2(n5853), .ZN(n5855) );
  XNOR2_X1 U7413 ( .A(n5855), .B(n6075), .ZN(n5857) );
  AOI22_X1 U7414 ( .A1(n5852), .A2(n6068), .B1(n7112), .B2(n4515), .ZN(n5856)
         );
  NAND2_X1 U7415 ( .A1(n5857), .A2(n5856), .ZN(n5860) );
  NAND2_X1 U7416 ( .A1(n5859), .A2(n7027), .ZN(n7030) );
  NAND2_X1 U7417 ( .A1(n9264), .A2(n4515), .ZN(n5863) );
  INV_X2 U7418 ( .A(n5861), .ZN(n5895) );
  INV_X4 U7419 ( .A(n5895), .ZN(n6077) );
  NAND2_X1 U7420 ( .A1(n8812), .A2(n6077), .ZN(n5862) );
  NAND2_X1 U7421 ( .A1(n5863), .A2(n5862), .ZN(n5864) );
  AOI22_X1 U7422 ( .A1(n9264), .A2(n6068), .B1(n8812), .B2(n4515), .ZN(n5870)
         );
  XNOR2_X1 U7423 ( .A(n5869), .B(n5870), .ZN(n8809) );
  NAND2_X1 U7424 ( .A1(n9263), .A2(n4515), .ZN(n5866) );
  NAND2_X1 U7425 ( .A1(n6077), .A2(n9865), .ZN(n5865) );
  NAND2_X1 U7426 ( .A1(n5866), .A2(n5865), .ZN(n5867) );
  XNOR2_X1 U7427 ( .A(n5867), .B(n6066), .ZN(n5875) );
  AND2_X1 U7428 ( .A1(n9865), .A2(n4515), .ZN(n5868) );
  XNOR2_X1 U7429 ( .A(n5875), .B(n5873), .ZN(n7049) );
  INV_X1 U7430 ( .A(n5869), .ZN(n5871) );
  NAND2_X1 U7431 ( .A1(n5871), .A2(n5870), .ZN(n7050) );
  AND2_X1 U7432 ( .A1(n7049), .A2(n7050), .ZN(n5872) );
  INV_X1 U7433 ( .A(n5873), .ZN(n5874) );
  NAND2_X1 U7434 ( .A1(n5875), .A2(n5874), .ZN(n5883) );
  NAND2_X1 U7435 ( .A1(n5880), .A2(n5883), .ZN(n5879) );
  NAND2_X1 U7436 ( .A1(n9262), .A2(n4515), .ZN(n5877) );
  NAND2_X1 U7437 ( .A1(n7219), .A2(n6077), .ZN(n5876) );
  NAND2_X1 U7438 ( .A1(n5877), .A2(n5876), .ZN(n5878) );
  XNOR2_X1 U7439 ( .A(n5878), .B(n6066), .ZN(n5881) );
  AOI22_X1 U7440 ( .A1(n9262), .A2(n6068), .B1(n7219), .B2(n4515), .ZN(n7142)
         );
  INV_X1 U7441 ( .A(n5881), .ZN(n5882) );
  AND2_X1 U7442 ( .A1(n5883), .A2(n5882), .ZN(n5884) );
  NAND2_X1 U7443 ( .A1(n9261), .A2(n4515), .ZN(n5886) );
  OR2_X1 U7444 ( .A1(n5895), .A2(n7353), .ZN(n5885) );
  NAND2_X1 U7445 ( .A1(n5886), .A2(n5885), .ZN(n5887) );
  XNOR2_X1 U7446 ( .A(n5887), .B(n6075), .ZN(n5890) );
  NAND2_X1 U7447 ( .A1(n9261), .A2(n6068), .ZN(n5889) );
  OR2_X1 U7448 ( .A1(n7353), .A2(n5844), .ZN(n5888) );
  AND2_X1 U7449 ( .A1(n5889), .A2(n5888), .ZN(n5891) );
  AND2_X1 U7450 ( .A1(n5890), .A2(n5891), .ZN(n7188) );
  INV_X1 U7451 ( .A(n5890), .ZN(n5893) );
  INV_X1 U7452 ( .A(n5891), .ZN(n5892) );
  NAND2_X1 U7453 ( .A1(n5893), .A2(n5892), .ZN(n7189) );
  NAND2_X1 U7454 ( .A1(n9260), .A2(n4515), .ZN(n5894) );
  OAI21_X1 U7455 ( .B1(n9898), .B2(n5895), .A(n5894), .ZN(n5896) );
  XNOR2_X1 U7456 ( .A(n5896), .B(n6075), .ZN(n7337) );
  OR2_X1 U7457 ( .A1(n9898), .A2(n5844), .ZN(n5898) );
  NAND2_X1 U7458 ( .A1(n9260), .A2(n6068), .ZN(n5897) );
  NAND2_X1 U7459 ( .A1(n7337), .A2(n7336), .ZN(n5899) );
  INV_X1 U7460 ( .A(n7337), .ZN(n5901) );
  INV_X1 U7461 ( .A(n7336), .ZN(n5900) );
  NAND2_X1 U7462 ( .A1(n5901), .A2(n5900), .ZN(n5902) );
  NAND2_X1 U7463 ( .A1(n5903), .A2(n5902), .ZN(n5907) );
  NAND2_X1 U7464 ( .A1(n7601), .A2(n6077), .ZN(n5904) );
  OAI21_X1 U7465 ( .B1(n7498), .B2(n6079), .A(n5904), .ZN(n5905) );
  XNOR2_X1 U7466 ( .A(n5905), .B(n6066), .ZN(n5906) );
  OR2_X1 U7467 ( .A1(n7498), .A2(n5908), .ZN(n5910) );
  NAND2_X1 U7468 ( .A1(n7601), .A2(n4515), .ZN(n5909) );
  NAND2_X1 U7469 ( .A1(n5910), .A2(n5909), .ZN(n7596) );
  INV_X1 U7470 ( .A(n7596), .ZN(n5911) );
  NAND2_X1 U7471 ( .A1(n7598), .A2(n5912), .ZN(n7651) );
  NAND2_X1 U7472 ( .A1(n7660), .A2(n6077), .ZN(n5914) );
  OR2_X1 U7473 ( .A1(n7484), .A2(n6079), .ZN(n5913) );
  NAND2_X1 U7474 ( .A1(n5914), .A2(n5913), .ZN(n5915) );
  XNOR2_X1 U7475 ( .A(n5915), .B(n6066), .ZN(n5917) );
  NOR2_X1 U7476 ( .A1(n7484), .A2(n5908), .ZN(n5916) );
  AOI21_X1 U7477 ( .B1(n7660), .B2(n4515), .A(n5916), .ZN(n5918) );
  XNOR2_X1 U7478 ( .A(n5917), .B(n5918), .ZN(n7652) );
  NAND2_X1 U7479 ( .A1(n7651), .A2(n7652), .ZN(n7650) );
  INV_X1 U7480 ( .A(n5917), .ZN(n5919) );
  NAND2_X1 U7481 ( .A1(n5919), .A2(n5918), .ZN(n5920) );
  INV_X1 U7482 ( .A(n5927), .ZN(n5925) );
  NAND2_X1 U7483 ( .A1(n7538), .A2(n6077), .ZN(n5922) );
  OR2_X1 U7484 ( .A1(n7634), .A2(n6079), .ZN(n5921) );
  NAND2_X1 U7485 ( .A1(n5922), .A2(n5921), .ZN(n5923) );
  XNOR2_X1 U7486 ( .A(n5923), .B(n6075), .ZN(n5926) );
  INV_X1 U7487 ( .A(n5926), .ZN(n5924) );
  NAND2_X1 U7488 ( .A1(n5925), .A2(n5924), .ZN(n5928) );
  NAND2_X1 U7489 ( .A1(n5927), .A2(n5926), .ZN(n5932) );
  NAND2_X1 U7490 ( .A1(n7538), .A2(n4515), .ZN(n5930) );
  OR2_X1 U7491 ( .A1(n7634), .A2(n6072), .ZN(n5929) );
  NAND2_X1 U7492 ( .A1(n5930), .A2(n5929), .ZN(n9757) );
  INV_X1 U7493 ( .A(n9757), .ZN(n5931) );
  NAND2_X1 U7494 ( .A1(n4622), .A2(n6077), .ZN(n5934) );
  OR2_X1 U7495 ( .A1(n7606), .A2(n6079), .ZN(n5933) );
  NAND2_X1 U7496 ( .A1(n5934), .A2(n5933), .ZN(n5935) );
  XNOR2_X1 U7497 ( .A(n5935), .B(n6066), .ZN(n5938) );
  NAND2_X1 U7498 ( .A1(n4622), .A2(n4515), .ZN(n5937) );
  OR2_X1 U7499 ( .A1(n7606), .A2(n6072), .ZN(n5936) );
  NAND2_X1 U7500 ( .A1(n5937), .A2(n5936), .ZN(n5939) );
  NAND2_X1 U7501 ( .A1(n5938), .A2(n5939), .ZN(n8919) );
  INV_X1 U7502 ( .A(n5938), .ZN(n5941) );
  INV_X1 U7503 ( .A(n5939), .ZN(n5940) );
  NAND2_X1 U7504 ( .A1(n5941), .A2(n5940), .ZN(n8921) );
  NAND2_X1 U7505 ( .A1(n8842), .A2(n6077), .ZN(n5943) );
  OR2_X1 U7506 ( .A1(n7700), .A2(n6079), .ZN(n5942) );
  NAND2_X1 U7507 ( .A1(n5943), .A2(n5942), .ZN(n5944) );
  XNOR2_X1 U7508 ( .A(n5944), .B(n6066), .ZN(n5946) );
  NOR2_X1 U7509 ( .A1(n7700), .A2(n6072), .ZN(n5945) );
  AOI21_X1 U7510 ( .B1(n8842), .B2(n4515), .A(n5945), .ZN(n5947) );
  XNOR2_X1 U7511 ( .A(n5946), .B(n5947), .ZN(n8835) );
  INV_X1 U7512 ( .A(n5946), .ZN(n5948) );
  NAND2_X1 U7513 ( .A1(n5948), .A2(n5947), .ZN(n5949) );
  NAND2_X1 U7514 ( .A1(n8901), .A2(n6077), .ZN(n5951) );
  OR2_X1 U7515 ( .A1(n7605), .A2(n6079), .ZN(n5950) );
  NAND2_X1 U7516 ( .A1(n5951), .A2(n5950), .ZN(n5952) );
  XNOR2_X1 U7517 ( .A(n5952), .B(n6066), .ZN(n5954) );
  NOR2_X1 U7518 ( .A1(n7605), .A2(n6072), .ZN(n5953) );
  AOI21_X1 U7519 ( .B1(n8901), .B2(n4515), .A(n5953), .ZN(n5955) );
  XNOR2_X1 U7520 ( .A(n5954), .B(n5955), .ZN(n8896) );
  INV_X1 U7521 ( .A(n5954), .ZN(n5956) );
  NAND2_X1 U7522 ( .A1(n9655), .A2(n6077), .ZN(n5958) );
  NAND2_X1 U7523 ( .A1(n9253), .A2(n4515), .ZN(n5957) );
  NAND2_X1 U7524 ( .A1(n5958), .A2(n5957), .ZN(n5959) );
  XNOR2_X1 U7525 ( .A(n5959), .B(n6066), .ZN(n5962) );
  AND2_X1 U7526 ( .A1(n9253), .A2(n6068), .ZN(n5960) );
  AOI21_X1 U7527 ( .B1(n9655), .B2(n4515), .A(n5960), .ZN(n8792) );
  INV_X1 U7528 ( .A(n5962), .ZN(n5963) );
  NAND2_X1 U7529 ( .A1(n5961), .A2(n5963), .ZN(n5964) );
  NAND2_X1 U7530 ( .A1(n9555), .A2(n6077), .ZN(n5966) );
  OR2_X1 U7531 ( .A1(n8869), .A2(n6079), .ZN(n5965) );
  NAND2_X1 U7532 ( .A1(n5966), .A2(n5965), .ZN(n5967) );
  XNOR2_X1 U7533 ( .A(n5967), .B(n6066), .ZN(n8854) );
  NAND2_X1 U7534 ( .A1(n9555), .A2(n4515), .ZN(n5969) );
  OR2_X1 U7535 ( .A1(n8869), .A2(n6072), .ZN(n5968) );
  NAND2_X1 U7536 ( .A1(n5969), .A2(n5968), .ZN(n8853) );
  NAND2_X1 U7537 ( .A1(n8854), .A2(n8853), .ZN(n8852) );
  NAND2_X1 U7538 ( .A1(n9025), .A2(n6077), .ZN(n5971) );
  NAND2_X1 U7539 ( .A1(n9252), .A2(n4515), .ZN(n5970) );
  NAND2_X1 U7540 ( .A1(n5971), .A2(n5970), .ZN(n5972) );
  XNOR2_X1 U7541 ( .A(n5972), .B(n6066), .ZN(n5977) );
  NAND2_X1 U7542 ( .A1(n9025), .A2(n4515), .ZN(n5974) );
  NAND2_X1 U7543 ( .A1(n9252), .A2(n6068), .ZN(n5973) );
  NAND2_X1 U7544 ( .A1(n5974), .A2(n5973), .ZN(n8952) );
  NAND2_X1 U7545 ( .A1(n5977), .A2(n8952), .ZN(n5975) );
  AND2_X1 U7546 ( .A1(n8852), .A2(n5975), .ZN(n5976) );
  NAND2_X1 U7547 ( .A1(n8855), .A2(n5976), .ZN(n5982) );
  INV_X1 U7548 ( .A(n8854), .ZN(n5980) );
  OAI21_X1 U7549 ( .B1(n5977), .B2(n8952), .A(n8853), .ZN(n5979) );
  NOR2_X1 U7550 ( .A1(n8853), .A2(n8952), .ZN(n5978) );
  INV_X1 U7551 ( .A(n5977), .ZN(n8856) );
  AOI22_X1 U7552 ( .A1(n5980), .A2(n5979), .B1(n5978), .B2(n8856), .ZN(n5981)
         );
  NAND2_X1 U7553 ( .A1(n5982), .A2(n5981), .ZN(n8865) );
  NAND2_X1 U7554 ( .A1(n9537), .A2(n6077), .ZN(n5984) );
  NAND2_X1 U7555 ( .A1(n9250), .A2(n4515), .ZN(n5983) );
  NAND2_X1 U7556 ( .A1(n5984), .A2(n5983), .ZN(n5985) );
  XNOR2_X1 U7557 ( .A(n5985), .B(n6066), .ZN(n5988) );
  NAND2_X1 U7558 ( .A1(n9537), .A2(n4514), .ZN(n5987) );
  NAND2_X1 U7559 ( .A1(n9250), .A2(n6068), .ZN(n5986) );
  NAND2_X1 U7560 ( .A1(n5987), .A2(n5986), .ZN(n5989) );
  NAND2_X1 U7561 ( .A1(n5988), .A2(n5989), .ZN(n8867) );
  NAND2_X1 U7562 ( .A1(n8865), .A2(n8867), .ZN(n5992) );
  INV_X1 U7563 ( .A(n5988), .ZN(n5991) );
  INV_X1 U7564 ( .A(n5989), .ZN(n5990) );
  NAND2_X1 U7565 ( .A1(n5991), .A2(n5990), .ZN(n8866) );
  NAND2_X1 U7566 ( .A1(n9502), .A2(n6077), .ZN(n5994) );
  NAND2_X1 U7567 ( .A1(n9248), .A2(n4515), .ZN(n5993) );
  NAND2_X1 U7568 ( .A1(n5994), .A2(n5993), .ZN(n5995) );
  XNOR2_X1 U7569 ( .A(n5995), .B(n6066), .ZN(n8819) );
  NAND2_X1 U7570 ( .A1(n9502), .A2(n4515), .ZN(n5997) );
  NAND2_X1 U7571 ( .A1(n9248), .A2(n6068), .ZN(n5996) );
  NAND2_X1 U7572 ( .A1(n5997), .A2(n5996), .ZN(n6004) );
  NAND2_X1 U7573 ( .A1(n9519), .A2(n6077), .ZN(n5999) );
  NAND2_X1 U7574 ( .A1(n9249), .A2(n4515), .ZN(n5998) );
  NAND2_X1 U7575 ( .A1(n5999), .A2(n5998), .ZN(n6000) );
  XNOR2_X1 U7576 ( .A(n6000), .B(n6066), .ZN(n6005) );
  NAND2_X1 U7577 ( .A1(n9519), .A2(n4515), .ZN(n6002) );
  NAND2_X1 U7578 ( .A1(n9249), .A2(n6068), .ZN(n6001) );
  NAND2_X1 U7579 ( .A1(n6002), .A2(n6001), .ZN(n8930) );
  OAI22_X1 U7580 ( .A1(n8819), .A2(n6004), .B1(n6005), .B2(n8930), .ZN(n6009)
         );
  INV_X1 U7581 ( .A(n6005), .ZN(n8817) );
  INV_X1 U7582 ( .A(n8930), .ZN(n6003) );
  INV_X1 U7583 ( .A(n6004), .ZN(n8818) );
  OAI21_X1 U7584 ( .B1(n8817), .B2(n6003), .A(n8818), .ZN(n6007) );
  AND2_X1 U7585 ( .A1(n6004), .A2(n8930), .ZN(n6006) );
  AOI22_X1 U7586 ( .A1(n8819), .A2(n6007), .B1(n6006), .B2(n6005), .ZN(n6008)
         );
  NAND2_X1 U7587 ( .A1(n9485), .A2(n6077), .ZN(n6011) );
  NAND2_X1 U7588 ( .A1(n9247), .A2(n4515), .ZN(n6010) );
  NAND2_X1 U7589 ( .A1(n6011), .A2(n6010), .ZN(n6012) );
  XNOR2_X1 U7590 ( .A(n6012), .B(n6075), .ZN(n8887) );
  AND2_X1 U7591 ( .A1(n9247), .A2(n6068), .ZN(n6013) );
  AOI21_X1 U7592 ( .B1(n9485), .B2(n4514), .A(n6013), .ZN(n6014) );
  INV_X1 U7593 ( .A(n8887), .ZN(n6015) );
  INV_X1 U7594 ( .A(n6014), .ZN(n8886) );
  NAND2_X1 U7595 ( .A1(n9470), .A2(n6077), .ZN(n6017) );
  NAND2_X1 U7596 ( .A1(n9246), .A2(n4515), .ZN(n6016) );
  NAND2_X1 U7597 ( .A1(n6017), .A2(n6016), .ZN(n6018) );
  XNOR2_X1 U7598 ( .A(n6018), .B(n6075), .ZN(n6021) );
  AND2_X1 U7599 ( .A1(n9246), .A2(n6068), .ZN(n6019) );
  AOI21_X1 U7600 ( .B1(n9470), .B2(n4515), .A(n6019), .ZN(n6020) );
  XNOR2_X1 U7601 ( .A(n6021), .B(n6020), .ZN(n8828) );
  NAND2_X1 U7602 ( .A1(n9451), .A2(n6077), .ZN(n6023) );
  NAND2_X1 U7603 ( .A1(n9245), .A2(n4515), .ZN(n6022) );
  NAND2_X1 U7604 ( .A1(n6023), .A2(n6022), .ZN(n6024) );
  XNOR2_X1 U7605 ( .A(n6024), .B(n6075), .ZN(n6027) );
  NAND2_X1 U7606 ( .A1(n9451), .A2(n6071), .ZN(n6026) );
  NAND2_X1 U7607 ( .A1(n9245), .A2(n6068), .ZN(n6025) );
  NAND2_X1 U7608 ( .A1(n6026), .A2(n6025), .ZN(n8907) );
  NAND2_X1 U7609 ( .A1(n9435), .A2(n6077), .ZN(n6030) );
  NAND2_X1 U7610 ( .A1(n9244), .A2(n4515), .ZN(n6029) );
  NAND2_X1 U7611 ( .A1(n6030), .A2(n6029), .ZN(n6031) );
  XNOR2_X1 U7612 ( .A(n6031), .B(n6075), .ZN(n6033) );
  AND2_X1 U7613 ( .A1(n9244), .A2(n6068), .ZN(n6032) );
  AOI21_X1 U7614 ( .B1(n9435), .B2(n4515), .A(n6032), .ZN(n6034) );
  NAND2_X1 U7615 ( .A1(n6033), .A2(n6034), .ZN(n8878) );
  INV_X1 U7616 ( .A(n6033), .ZN(n6036) );
  INV_X1 U7617 ( .A(n6034), .ZN(n6035) );
  NAND2_X1 U7618 ( .A1(n6036), .A2(n6035), .ZN(n6037) );
  NAND2_X1 U7619 ( .A1(n9420), .A2(n6077), .ZN(n6039) );
  NAND2_X1 U7620 ( .A1(n8847), .A2(n4515), .ZN(n6038) );
  NAND2_X1 U7621 ( .A1(n6039), .A2(n6038), .ZN(n6040) );
  XNOR2_X1 U7622 ( .A(n6040), .B(n6075), .ZN(n6042) );
  AND2_X1 U7623 ( .A1(n8847), .A2(n6068), .ZN(n6041) );
  AOI21_X1 U7624 ( .B1(n9420), .B2(n4514), .A(n6041), .ZN(n6043) );
  NAND2_X1 U7625 ( .A1(n6042), .A2(n6043), .ZN(n6047) );
  INV_X1 U7626 ( .A(n6042), .ZN(n6045) );
  INV_X1 U7627 ( .A(n6043), .ZN(n6044) );
  NAND2_X1 U7628 ( .A1(n6045), .A2(n6044), .ZN(n6046) );
  NAND2_X1 U7629 ( .A1(n6047), .A2(n6046), .ZN(n8877) );
  INV_X1 U7630 ( .A(n6047), .ZN(n6048) );
  AOI22_X1 U7631 ( .A1(n9404), .A2(n4515), .B1(n6068), .B2(n9243), .ZN(n6058)
         );
  NAND2_X1 U7632 ( .A1(n9404), .A2(n6077), .ZN(n6050) );
  NAND2_X1 U7633 ( .A1(n9243), .A2(n4514), .ZN(n6049) );
  NAND2_X1 U7634 ( .A1(n6050), .A2(n6049), .ZN(n6051) );
  XNOR2_X1 U7635 ( .A(n6051), .B(n6066), .ZN(n6060) );
  XOR2_X1 U7636 ( .A(n6058), .B(n6060), .Z(n8845) );
  NAND2_X1 U7637 ( .A1(n9392), .A2(n6077), .ZN(n6054) );
  NAND2_X1 U7638 ( .A1(n9242), .A2(n4515), .ZN(n6053) );
  NAND2_X1 U7639 ( .A1(n6054), .A2(n6053), .ZN(n6055) );
  XNOR2_X1 U7640 ( .A(n6055), .B(n6075), .ZN(n6062) );
  NOR2_X1 U7641 ( .A1(n6056), .A2(n6072), .ZN(n6057) );
  AOI21_X1 U7642 ( .B1(n9392), .B2(n4514), .A(n6057), .ZN(n6063) );
  XNOR2_X1 U7643 ( .A(n6062), .B(n6063), .ZN(n8939) );
  INV_X1 U7644 ( .A(n6058), .ZN(n6059) );
  NOR2_X1 U7645 ( .A1(n6060), .A2(n6059), .ZN(n8940) );
  INV_X1 U7646 ( .A(n6062), .ZN(n6065) );
  INV_X1 U7647 ( .A(n6063), .ZN(n6064) );
  AOI22_X1 U7648 ( .A1(n9375), .A2(n6077), .B1(n4515), .B2(n9241), .ZN(n6067)
         );
  XNOR2_X1 U7649 ( .A(n6067), .B(n6066), .ZN(n6070) );
  AOI22_X1 U7650 ( .A1(n9375), .A2(n4515), .B1(n6068), .B2(n9241), .ZN(n6069)
         );
  NAND2_X1 U7651 ( .A1(n6070), .A2(n6069), .ZN(n6103) );
  OAI21_X1 U7652 ( .B1(n6070), .B2(n6069), .A(n6103), .ZN(n6129) );
  NAND2_X1 U7653 ( .A1(n6119), .A2(n4515), .ZN(n6074) );
  OR2_X1 U7654 ( .A1(n7024), .A2(n6072), .ZN(n6073) );
  NAND2_X1 U7655 ( .A1(n6074), .A2(n6073), .ZN(n6076) );
  XNOR2_X1 U7656 ( .A(n6076), .B(n6075), .ZN(n6081) );
  NAND2_X1 U7657 ( .A1(n6119), .A2(n6077), .ZN(n6078) );
  OAI21_X1 U7658 ( .B1(n7024), .B2(n6079), .A(n6078), .ZN(n6080) );
  XNOR2_X1 U7659 ( .A(n6081), .B(n6080), .ZN(n6087) );
  INV_X1 U7660 ( .A(n6087), .ZN(n6104) );
  AND2_X1 U7661 ( .A1(n6082), .A2(P1_D_REG_1__SCAN_IN), .ZN(n6083) );
  OR2_X1 U7662 ( .A1(n9716), .A2(n6083), .ZN(n6084) );
  NAND2_X1 U7663 ( .A1(n6084), .A2(n9718), .ZN(n7098) );
  OR2_X1 U7664 ( .A1(n7099), .A2(n7098), .ZN(n6096) );
  NAND3_X1 U7665 ( .A1(n6657), .A2(P1_STATE_REG_SCAN_IN), .A3(n6700), .ZN(
        n6701) );
  NOR2_X1 U7666 ( .A1(n6096), .A2(n6701), .ZN(n6094) );
  NOR2_X1 U7667 ( .A1(n9656), .A2(n6698), .ZN(n6085) );
  NAND3_X1 U7668 ( .A1(n6104), .A2(n8942), .A3(n6103), .ZN(n6086) );
  OR2_X1 U7669 ( .A1(n6131), .A2(n6086), .ZN(n6111) );
  NAND2_X1 U7670 ( .A1(n6088), .A2(n9224), .ZN(n7103) );
  INV_X1 U7671 ( .A(n7103), .ZN(n6089) );
  NAND2_X1 U7672 ( .A1(n6094), .A2(n6089), .ZN(n6091) );
  INV_X1 U7673 ( .A(n6095), .ZN(n6090) );
  INV_X1 U7674 ( .A(n6701), .ZN(n9717) );
  OR2_X1 U7675 ( .A1(n8947), .A2(n8944), .ZN(n6093) );
  OR2_X1 U7676 ( .A1(n6939), .A2(n8946), .ZN(n6092) );
  NAND2_X1 U7677 ( .A1(n6093), .A2(n6092), .ZN(n6117) );
  INV_X1 U7678 ( .A(n6117), .ZN(n6102) );
  INV_X1 U7679 ( .A(n9764), .ZN(n8912) );
  NAND2_X1 U7680 ( .A1(n6096), .A2(n6095), .ZN(n6099) );
  INV_X1 U7681 ( .A(n6097), .ZN(n6098) );
  NAND2_X1 U7682 ( .A1(n6099), .A2(n6098), .ZN(n6100) );
  NAND2_X1 U7683 ( .A1(n6100), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9772) );
  INV_X1 U7684 ( .A(n9772), .ZN(n8883) );
  AOI22_X1 U7685 ( .A1(n9358), .A2(n8883), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3086), .ZN(n6101) );
  OAI21_X1 U7686 ( .B1(n6102), .B2(n8912), .A(n6101), .ZN(n6106) );
  NOR3_X1 U7687 ( .A1(n6104), .A2(n6103), .A3(n9758), .ZN(n6105) );
  AOI211_X1 U7688 ( .C1(n6119), .C2(n8958), .A(n6106), .B(n6105), .ZN(n6107)
         );
  AOI21_X1 U7689 ( .B1(n6131), .B2(n6109), .A(n6108), .ZN(n6110) );
  NAND2_X1 U7690 ( .A1(n6111), .A2(n6110), .ZN(P1_U3220) );
  NAND2_X1 U7691 ( .A1(n6112), .A2(n9135), .ZN(n6113) );
  INV_X1 U7692 ( .A(n9135), .ZN(n6115) );
  XNOR2_X1 U7693 ( .A(n6116), .B(n6115), .ZN(n6118) );
  AOI21_X1 U7694 ( .B1(n6119), .B2(n9373), .A(n9578), .ZN(n6121) );
  NAND2_X1 U7695 ( .A1(n6121), .A2(n6120), .ZN(n9357) );
  NAND2_X1 U7696 ( .A1(n9365), .A2(n9357), .ZN(n6122) );
  AOI21_X1 U7697 ( .B1(n9356), .B2(n9908), .A(n6122), .ZN(n6126) );
  MUX2_X1 U7698 ( .A(n6124), .B(n6126), .S(n9918), .Z(n6125) );
  NAND2_X1 U7699 ( .A1(n6125), .A2(n5137), .ZN(P1_U3550) );
  INV_X1 U7700 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n6127) );
  MUX2_X1 U7701 ( .A(n6127), .B(n6126), .S(n9911), .Z(n6128) );
  NAND2_X1 U7702 ( .A1(n6128), .A2(n5138), .ZN(P1_U3518) );
  AOI21_X1 U7703 ( .B1(n8943), .B2(n4518), .A(n4610), .ZN(n6130) );
  OAI21_X1 U7704 ( .B1(n6131), .B2(n6130), .A(n8942), .ZN(n6140) );
  OR2_X1 U7705 ( .A1(n7024), .A2(n8946), .ZN(n6133) );
  NAND2_X1 U7706 ( .A1(n9242), .A2(n9232), .ZN(n6132) );
  NAND2_X1 U7707 ( .A1(n6133), .A2(n6132), .ZN(n9370) );
  INV_X1 U7708 ( .A(n9376), .ZN(n6135) );
  OAI22_X1 U7709 ( .A1(n6135), .A2(n9772), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n6134), .ZN(n6136) );
  AOI21_X1 U7710 ( .B1(n9370), .B2(n9764), .A(n6136), .ZN(n6137) );
  INV_X1 U7711 ( .A(n6138), .ZN(n6139) );
  NAND2_X1 U7712 ( .A1(n6140), .A2(n6139), .ZN(P1_U3214) );
  NOR2_X1 U7713 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n6147) );
  NOR2_X1 U7714 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n6146) );
  INV_X1 U7715 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n6144) );
  NAND4_X1 U7716 ( .A1(n6147), .A2(n6146), .A3(n6145), .A4(n6144), .ZN(n6150)
         );
  INV_X1 U7717 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n6148) );
  NAND4_X1 U7718 ( .A1(n6550), .A2(n6398), .A3(n6447), .A4(n6148), .ZN(n6149)
         );
  INV_X1 U7719 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n6155) );
  NAND2_X1 U7720 ( .A1(n8162), .A2(n6203), .ZN(n6160) );
  OR2_X1 U7721 ( .A1(n8075), .A2(n8778), .ZN(n6159) );
  INV_X1 U7722 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n6167) );
  OR2_X2 U7723 ( .A1(n6357), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n6368) );
  OR2_X2 U7724 ( .A1(n6368), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6380) );
  INV_X1 U7725 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n10410) );
  INV_X1 U7726 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n6170) );
  OR2_X2 U7727 ( .A1(n6402), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n6414) );
  INV_X1 U7728 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n10299) );
  OR2_X2 U7729 ( .A1(n6426), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n6438) );
  INV_X1 U7730 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n6173) );
  OR2_X2 U7731 ( .A1(n6453), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n6463) );
  INV_X1 U7732 ( .A(n6463), .ZN(n6176) );
  INV_X1 U7733 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n6175) );
  OR2_X2 U7734 ( .A1(n6470), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n6480) );
  INV_X1 U7735 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n10315) );
  OR2_X2 U7736 ( .A1(n6499), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6501) );
  INV_X1 U7737 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n6178) );
  INV_X1 U7738 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n6180) );
  INV_X1 U7739 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n6182) );
  NAND2_X1 U7740 ( .A1(n6521), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n6184) );
  NAND2_X1 U7741 ( .A1(n6530), .A2(n6184), .ZN(n8496) );
  INV_X1 U7742 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n6187) );
  INV_X1 U7743 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n8764) );
  XNOR2_X2 U7745 ( .A(n6188), .B(n6187), .ZN(n8161) );
  NAND2_X1 U7746 ( .A1(n8496), .A2(n6540), .ZN(n6196) );
  INV_X1 U7747 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n8495) );
  NAND2_X1 U7748 ( .A1(n6532), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n6193) );
  NAND2_X1 U7749 ( .A1(n6491), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n6192) );
  OAI211_X1 U7750 ( .C1(n8495), .C2(n4507), .A(n6193), .B(n6192), .ZN(n6194)
         );
  INV_X1 U7751 ( .A(n6194), .ZN(n6195) );
  NAND2_X2 U7752 ( .A1(n6196), .A2(n6195), .ZN(n8502) );
  NAND2_X1 U7753 ( .A1(n6501), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n6197) );
  NAND2_X1 U7754 ( .A1(n6510), .A2(n6197), .ZN(n8526) );
  NAND2_X1 U7755 ( .A1(n8526), .A2(n6540), .ZN(n6202) );
  INV_X1 U7756 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n10408) );
  NAND2_X1 U7757 ( .A1(n6532), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n6199) );
  INV_X1 U7758 ( .A(n4507), .ZN(n6542) );
  NAND2_X1 U7759 ( .A1(n6542), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n6198) );
  OAI211_X1 U7760 ( .C1(n6543), .C2(n10408), .A(n6199), .B(n6198), .ZN(n6200)
         );
  INV_X1 U7761 ( .A(n6200), .ZN(n6201) );
  NAND2_X1 U7762 ( .A1(n7906), .A2(n6203), .ZN(n6206) );
  OR2_X1 U7763 ( .A1(n8075), .A2(n6204), .ZN(n6205) );
  INV_X1 U7764 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n7225) );
  INV_X1 U7765 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n10467) );
  OR2_X1 U7766 ( .A1(n6255), .A2(n10467), .ZN(n6209) );
  NAND2_X1 U7767 ( .A1(n6216), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n6208) );
  INV_X1 U7768 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n6912) );
  OR2_X1 U7769 ( .A1(n6229), .A2(n6912), .ZN(n6207) );
  NAND2_X1 U7770 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n6211) );
  MUX2_X1 U7771 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6211), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n6215) );
  INV_X1 U7772 ( .A(n6213), .ZN(n6214) );
  INV_X1 U7773 ( .A(n9935), .ZN(n6744) );
  NAND2_X1 U7774 ( .A1(n6224), .A2(n4509), .ZN(n7949) );
  NAND2_X1 U7775 ( .A1(n6216), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n6221) );
  INV_X1 U7776 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n6742) );
  OR2_X1 U7777 ( .A1(n6255), .A2(n6742), .ZN(n6220) );
  INV_X1 U7778 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n7207) );
  OR2_X1 U7779 ( .A1(n4507), .A2(n7207), .ZN(n6219) );
  INV_X1 U7780 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n6217) );
  OR2_X1 U7781 ( .A1(n6229), .A2(n6217), .ZN(n6218) );
  INV_X1 U7782 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n6729) );
  NAND2_X1 U7783 ( .A1(n7936), .A2(SI_0_), .ZN(n6223) );
  INV_X1 U7784 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n6222) );
  XNOR2_X1 U7785 ( .A(n6223), .B(n6222), .ZN(n8788) );
  MUX2_X1 U7786 ( .A(n6729), .B(n8788), .S(n6587), .Z(n7209) );
  OR2_X1 U7787 ( .A1(n6689), .A2(n7209), .ZN(n6862) );
  NAND2_X1 U7788 ( .A1(n6561), .A2(n6862), .ZN(n6861) );
  NAND2_X1 U7789 ( .A1(n6224), .A2(n6225), .ZN(n6226) );
  NAND2_X1 U7790 ( .A1(n6861), .A2(n6226), .ZN(n6984) );
  INV_X1 U7791 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n6227) );
  NAND2_X1 U7792 ( .A1(n4506), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6232) );
  INV_X1 U7793 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n6724) );
  OR2_X1 U7794 ( .A1(n4507), .A2(n6724), .ZN(n6231) );
  INV_X1 U7795 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n6228) );
  OR2_X1 U7796 ( .A1(n6229), .A2(n6228), .ZN(n6230) );
  INV_X1 U7797 ( .A(n6308), .ZN(n6235) );
  OR2_X1 U7798 ( .A1(n6263), .A2(n6665), .ZN(n6237) );
  OR2_X1 U7799 ( .A1(n8075), .A2(n6659), .ZN(n6236) );
  OAI211_X1 U7800 ( .C1(n6587), .C2(n6760), .A(n6237), .B(n6236), .ZN(n7954)
         );
  OR2_X1 U7801 ( .A1(n8318), .A2(n7954), .ZN(n6238) );
  NAND2_X1 U7802 ( .A1(n6985), .A2(n6238), .ZN(n7300) );
  NAND2_X1 U7803 ( .A1(n6532), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6244) );
  INV_X1 U7804 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n6239) );
  OR2_X1 U7805 ( .A1(n6543), .A2(n6239), .ZN(n6243) );
  INV_X1 U7806 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n6240) );
  OR2_X1 U7807 ( .A1(n4507), .A2(n6240), .ZN(n6242) );
  OR2_X1 U7808 ( .A1(n6229), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n6241) );
  NOR2_X1 U7809 ( .A1(n6308), .A2(n6246), .ZN(n6245) );
  INV_X1 U7810 ( .A(n6247), .ZN(n6249) );
  NAND2_X1 U7811 ( .A1(n6308), .A2(n6248), .ZN(n6279) );
  NAND2_X1 U7812 ( .A1(n6249), .A2(n6279), .ZN(n6779) );
  OR2_X1 U7813 ( .A1(n6263), .A2(n6668), .ZN(n6251) );
  OR2_X1 U7814 ( .A1(n8075), .A2(n6660), .ZN(n6250) );
  OAI211_X1 U7815 ( .C1(n6587), .C2(n6779), .A(n6251), .B(n6250), .ZN(n10109)
         );
  INV_X1 U7816 ( .A(n10109), .ZN(n6996) );
  OR2_X1 U7817 ( .A1(n7953), .A2(n6996), .ZN(n6252) );
  NAND2_X1 U7818 ( .A1(n7300), .A2(n6252), .ZN(n6254) );
  NAND2_X1 U7819 ( .A1(n7953), .A2(n6996), .ZN(n6253) );
  NAND2_X1 U7820 ( .A1(n6491), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n6260) );
  INV_X1 U7821 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n6777) );
  OR2_X1 U7822 ( .A1(n4517), .A2(n6777), .ZN(n6259) );
  NAND2_X1 U7823 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n6256) );
  AND2_X1 U7824 ( .A1(n6272), .A2(n6256), .ZN(n7019) );
  OR2_X1 U7825 ( .A1(n6229), .A2(n7019), .ZN(n6258) );
  INV_X1 U7826 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n7377) );
  OR2_X1 U7827 ( .A1(n4507), .A2(n7377), .ZN(n6257) );
  NAND2_X1 U7828 ( .A1(n7375), .A2(n7123), .ZN(n6266) );
  NAND2_X1 U7829 ( .A1(n6279), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6262) );
  INV_X1 U7830 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n6261) );
  OR2_X1 U7831 ( .A1(n6263), .A2(n6663), .ZN(n6265) );
  OR2_X1 U7832 ( .A1(n8075), .A2(n6661), .ZN(n6264) );
  NAND2_X1 U7833 ( .A1(n6266), .A2(n10117), .ZN(n6270) );
  NAND2_X1 U7834 ( .A1(n6268), .A2(n6267), .ZN(n6269) );
  NAND2_X1 U7835 ( .A1(n6491), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n6278) );
  INV_X1 U7836 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n6271) );
  OR2_X1 U7837 ( .A1(n4517), .A2(n6271), .ZN(n6277) );
  NAND2_X1 U7838 ( .A1(n6272), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n6273) );
  AND2_X1 U7839 ( .A1(n6295), .A2(n6273), .ZN(n7306) );
  OR2_X1 U7840 ( .A1(n6229), .A2(n7306), .ZN(n6276) );
  INV_X1 U7841 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n6274) );
  OR2_X1 U7842 ( .A1(n4507), .A2(n6274), .ZN(n6275) );
  NAND4_X1 U7843 ( .A1(n6278), .A2(n6277), .A3(n6276), .A4(n6275), .ZN(n8316)
         );
  NAND2_X1 U7844 ( .A1(n6286), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6281) );
  INV_X1 U7845 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n6280) );
  XNOR2_X1 U7846 ( .A(n6281), .B(n6280), .ZN(n9951) );
  NAND2_X1 U7847 ( .A1(n6670), .A2(n6203), .ZN(n6283) );
  INV_X1 U7848 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6673) );
  OR2_X1 U7849 ( .A1(n8075), .A2(n6673), .ZN(n6282) );
  OAI211_X1 U7850 ( .C1(n6587), .C2(n9951), .A(n6283), .B(n6282), .ZN(n7125)
         );
  AND2_X1 U7851 ( .A1(n8316), .A2(n7125), .ZN(n6285) );
  OR2_X1 U7852 ( .A1(n8316), .A2(n7125), .ZN(n6284) );
  NAND2_X1 U7853 ( .A1(n6677), .A2(n6203), .ZN(n6293) );
  NOR2_X1 U7854 ( .A1(n6286), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n6289) );
  NOR2_X1 U7855 ( .A1(n6289), .A2(n6246), .ZN(n6287) );
  MUX2_X1 U7856 ( .A(n6246), .B(n6287), .S(P2_IR_REG_6__SCAN_IN), .Z(n6291) );
  INV_X1 U7857 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n6288) );
  NAND2_X1 U7858 ( .A1(n6289), .A2(n6288), .ZN(n6305) );
  INV_X1 U7859 ( .A(n6305), .ZN(n6290) );
  INV_X1 U7860 ( .A(n9976), .ZN(n7810) );
  NAND2_X1 U7861 ( .A1(n7290), .A2(n10120), .ZN(n6301) );
  NAND2_X1 U7862 ( .A1(n6532), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6300) );
  INV_X1 U7863 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n6294) );
  OR2_X1 U7864 ( .A1(n6543), .A2(n6294), .ZN(n6299) );
  NAND2_X1 U7865 ( .A1(n6295), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n6296) );
  AND2_X1 U7866 ( .A1(n6313), .A2(n6296), .ZN(n7289) );
  OR2_X1 U7867 ( .A1(n6229), .A2(n7289), .ZN(n6298) );
  INV_X1 U7868 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n7764) );
  OR2_X1 U7869 ( .A1(n4507), .A2(n7764), .ZN(n6297) );
  NAND2_X1 U7870 ( .A1(n6301), .A2(n8315), .ZN(n6304) );
  INV_X1 U7871 ( .A(n7290), .ZN(n6302) );
  INV_X1 U7872 ( .A(n10120), .ZN(n7179) );
  NAND2_X1 U7873 ( .A1(n6302), .A2(n7179), .ZN(n6303) );
  NAND2_X1 U7874 ( .A1(n6304), .A2(n6303), .ZN(n7315) );
  NAND2_X1 U7875 ( .A1(n6681), .A2(n6203), .ZN(n6311) );
  NAND2_X1 U7876 ( .A1(n6305), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6306) );
  MUX2_X1 U7877 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6306), .S(
        P2_IR_REG_7__SCAN_IN), .Z(n6309) );
  NAND2_X1 U7878 ( .A1(n6308), .A2(n6307), .ZN(n6322) );
  AOI22_X1 U7879 ( .A1(n6460), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n6655), .B2(
        n7787), .ZN(n6310) );
  NAND2_X1 U7880 ( .A1(n6311), .A2(n6310), .ZN(n10128) );
  NAND2_X1 U7881 ( .A1(n6491), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n6319) );
  INV_X1 U7882 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n6312) );
  OR2_X1 U7883 ( .A1(n4507), .A2(n6312), .ZN(n6318) );
  NAND2_X1 U7884 ( .A1(n6313), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n6314) );
  AND2_X1 U7885 ( .A1(n6327), .A2(n6314), .ZN(n7321) );
  OR2_X1 U7886 ( .A1(n6229), .A2(n7321), .ZN(n6317) );
  INV_X1 U7887 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n6315) );
  OR2_X1 U7888 ( .A1(n4517), .A2(n6315), .ZN(n6316) );
  NAND4_X1 U7889 ( .A1(n6319), .A2(n6318), .A3(n6317), .A4(n6316), .ZN(n8314)
         );
  NAND2_X1 U7890 ( .A1(n10128), .A2(n7161), .ZN(n7985) );
  NAND2_X1 U7891 ( .A1(n6685), .A2(n6203), .ZN(n6325) );
  NAND2_X1 U7892 ( .A1(n6322), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6321) );
  MUX2_X1 U7893 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6321), .S(
        P2_IR_REG_8__SCAN_IN), .Z(n6323) );
  OR2_X1 U7894 ( .A1(n6322), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n6350) );
  AND2_X1 U7895 ( .A1(n6323), .A2(n6350), .ZN(n10004) );
  AOI22_X1 U7896 ( .A1(n6460), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n6655), .B2(
        n10004), .ZN(n6324) );
  NAND2_X1 U7897 ( .A1(n6325), .A2(n6324), .ZN(n10134) );
  NAND2_X1 U7898 ( .A1(n6491), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n6333) );
  INV_X1 U7899 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n6326) );
  OR2_X1 U7900 ( .A1(n4517), .A2(n6326), .ZN(n6332) );
  NAND2_X1 U7901 ( .A1(n6327), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n6328) );
  AND2_X1 U7902 ( .A1(n6339), .A2(n6328), .ZN(n7402) );
  OR2_X1 U7903 ( .A1(n6229), .A2(n7402), .ZN(n6331) );
  INV_X1 U7904 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n6329) );
  OR2_X1 U7905 ( .A1(n4507), .A2(n6329), .ZN(n6330) );
  NAND4_X1 U7906 ( .A1(n6333), .A2(n6332), .A3(n6331), .A4(n6330), .ZN(n8313)
         );
  INV_X1 U7907 ( .A(n8313), .ZN(n7382) );
  NAND2_X1 U7908 ( .A1(n10134), .A2(n7382), .ZN(n7986) );
  NAND2_X1 U7909 ( .A1(n7979), .A2(n7986), .ZN(n8118) );
  OR2_X1 U7910 ( .A1(n10128), .A2(n8314), .ZN(n7398) );
  AND2_X1 U7911 ( .A1(n8118), .A2(n7398), .ZN(n6334) );
  NAND2_X1 U7912 ( .A1(n10134), .A2(n8313), .ZN(n6335) );
  NAND2_X1 U7913 ( .A1(n6350), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6336) );
  XNOR2_X1 U7914 ( .A(n6336), .B(P2_IR_REG_9__SCAN_IN), .ZN(n10017) );
  AOI22_X1 U7915 ( .A1(n6460), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6655), .B2(
        n10017), .ZN(n6337) );
  NAND2_X1 U7916 ( .A1(n6491), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n6345) );
  INV_X1 U7917 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n6338) );
  OR2_X1 U7918 ( .A1(n4517), .A2(n6338), .ZN(n6344) );
  NAND2_X1 U7919 ( .A1(n6339), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n6340) );
  AND2_X1 U7920 ( .A1(n6357), .A2(n6340), .ZN(n7453) );
  OR2_X1 U7921 ( .A1(n6229), .A2(n7453), .ZN(n6343) );
  INV_X1 U7922 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n6341) );
  OR2_X1 U7923 ( .A1(n4507), .A2(n6341), .ZN(n6342) );
  NAND4_X1 U7924 ( .A1(n6345), .A2(n6344), .A3(n6343), .A4(n6342), .ZN(n8312)
         );
  AND2_X1 U7925 ( .A1(n10139), .A2(n8312), .ZN(n6349) );
  INV_X1 U7926 ( .A(n10139), .ZN(n6347) );
  NAND2_X1 U7927 ( .A1(n6705), .A2(n6203), .ZN(n6355) );
  OAI21_X1 U7928 ( .B1(n6350), .B2(P2_IR_REG_9__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n6352) );
  MUX2_X1 U7929 ( .A(n6352), .B(P2_IR_REG_31__SCAN_IN), .S(n6351), .Z(n6353)
         );
  AND2_X1 U7930 ( .A1(n6376), .A2(n6353), .ZN(n10031) );
  AOI22_X1 U7931 ( .A1(n6460), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6655), .B2(
        n10031), .ZN(n6354) );
  NAND2_X1 U7932 ( .A1(n6491), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n6362) );
  INV_X1 U7933 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n6356) );
  OR2_X1 U7934 ( .A1(n4517), .A2(n6356), .ZN(n6361) );
  NAND2_X1 U7935 ( .A1(n6357), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n6358) );
  AND2_X1 U7936 ( .A1(n6368), .A2(n6358), .ZN(n7523) );
  OR2_X1 U7937 ( .A1(n6229), .A2(n7523), .ZN(n6360) );
  INV_X1 U7938 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7773) );
  OR2_X1 U7939 ( .A1(n4507), .A2(n7773), .ZN(n6359) );
  NAND2_X1 U7940 ( .A1(n10146), .A2(n8311), .ZN(n6363) );
  NAND2_X1 U7941 ( .A1(n6718), .A2(n6203), .ZN(n6367) );
  NAND2_X1 U7942 ( .A1(n6376), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6365) );
  XNOR2_X1 U7943 ( .A(n6365), .B(P2_IR_REG_11__SCAN_IN), .ZN(n7819) );
  AOI22_X1 U7944 ( .A1(n6460), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n6655), .B2(
        n7819), .ZN(n6366) );
  NAND2_X1 U7945 ( .A1(n6491), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n6373) );
  INV_X1 U7946 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n7817) );
  OR2_X1 U7947 ( .A1(n4517), .A2(n7817), .ZN(n6372) );
  NAND2_X1 U7948 ( .A1(n6368), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6369) );
  AND2_X1 U7949 ( .A1(n6380), .A2(n6369), .ZN(n7440) );
  OR2_X1 U7950 ( .A1(n6229), .A2(n7440), .ZN(n6371) );
  INV_X1 U7951 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n7818) );
  OR2_X1 U7952 ( .A1(n4507), .A2(n7818), .ZN(n6370) );
  NAND2_X1 U7953 ( .A1(n8686), .A2(n7675), .ZN(n7997) );
  NAND2_X1 U7954 ( .A1(n7995), .A2(n7997), .ZN(n8124) );
  NAND2_X1 U7955 ( .A1(n7665), .A2(n8124), .ZN(n6375) );
  INV_X1 U7956 ( .A(n7675), .ZN(n8310) );
  NAND2_X1 U7957 ( .A1(n8686), .A2(n8310), .ZN(n6374) );
  NAND2_X1 U7958 ( .A1(n6833), .A2(n6203), .ZN(n6379) );
  NAND2_X1 U7959 ( .A1(n6388), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6377) );
  XNOR2_X1 U7960 ( .A(n6377), .B(P2_IR_REG_12__SCAN_IN), .ZN(n10068) );
  AOI22_X1 U7961 ( .A1(n6460), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n6655), .B2(
        n10068), .ZN(n6378) );
  NAND2_X1 U7962 ( .A1(n6491), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n6385) );
  INV_X1 U7963 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n7796) );
  OR2_X1 U7964 ( .A1(n4517), .A2(n7796), .ZN(n6384) );
  NAND2_X1 U7965 ( .A1(n6380), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n6381) );
  AND2_X1 U7966 ( .A1(n6392), .A2(n6381), .ZN(n7681) );
  OR2_X1 U7967 ( .A1(n6229), .A2(n7681), .ZN(n6383) );
  INV_X1 U7968 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n7775) );
  OR2_X1 U7969 ( .A1(n4507), .A2(n7775), .ZN(n6382) );
  NAND4_X1 U7970 ( .A1(n6385), .A2(n6384), .A3(n6383), .A4(n6382), .ZN(n8309)
         );
  AND2_X1 U7971 ( .A1(n8000), .A2(n8309), .ZN(n6387) );
  NAND2_X1 U7972 ( .A1(n6914), .A2(n6203), .ZN(n6391) );
  OR2_X1 U7973 ( .A1(n6399), .A2(n6246), .ZN(n6389) );
  XNOR2_X1 U7974 ( .A(n6389), .B(P2_IR_REG_13__SCAN_IN), .ZN(n8321) );
  AOI22_X1 U7975 ( .A1(n6460), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n6655), .B2(
        n8321), .ZN(n6390) );
  NAND2_X1 U7976 ( .A1(n6491), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n6397) );
  INV_X1 U7977 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n10413) );
  OR2_X1 U7978 ( .A1(n4517), .A2(n10413), .ZN(n6396) );
  NAND2_X1 U7979 ( .A1(n6392), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n6393) );
  AND2_X1 U7980 ( .A1(n6402), .A2(n6393), .ZN(n7742) );
  OR2_X1 U7981 ( .A1(n6229), .A2(n7742), .ZN(n6395) );
  INV_X1 U7982 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n7825) );
  OR2_X1 U7983 ( .A1(n4507), .A2(n7825), .ZN(n6394) );
  NOR2_X1 U7984 ( .A1(n8005), .A2(n8308), .ZN(n8008) );
  NAND2_X1 U7985 ( .A1(n8005), .A2(n8308), .ZN(n8007) );
  NAND2_X1 U7986 ( .A1(n6974), .A2(n6203), .ZN(n6401) );
  NAND2_X1 U7987 ( .A1(n4603), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6423) );
  XNOR2_X1 U7988 ( .A(n6423), .B(P2_IR_REG_14__SCAN_IN), .ZN(n8350) );
  AOI22_X1 U7989 ( .A1(n6460), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n6655), .B2(
        n8350), .ZN(n6400) );
  NAND2_X1 U7990 ( .A1(n6491), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n6407) );
  INV_X1 U7991 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n10395) );
  OR2_X1 U7992 ( .A1(n4517), .A2(n10395), .ZN(n6406) );
  NAND2_X1 U7993 ( .A1(n6402), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n6403) );
  AND2_X1 U7994 ( .A1(n6414), .A2(n6403), .ZN(n7888) );
  OR2_X1 U7995 ( .A1(n6229), .A2(n7888), .ZN(n6405) );
  INV_X1 U7996 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n8333) );
  OR2_X1 U7997 ( .A1(n4507), .A2(n8333), .ZN(n6404) );
  NAND4_X1 U7998 ( .A1(n6407), .A2(n6406), .A3(n6405), .A4(n6404), .ZN(n8307)
         );
  AND2_X1 U7999 ( .A1(n7887), .A2(n8307), .ZN(n6409) );
  OR2_X1 U8000 ( .A1(n7887), .A2(n8307), .ZN(n6408) );
  NAND2_X1 U8001 ( .A1(n7038), .A2(n6203), .ZN(n6413) );
  INV_X1 U8002 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n6421) );
  NAND2_X1 U8003 ( .A1(n6423), .A2(n6421), .ZN(n6410) );
  NAND2_X1 U8004 ( .A1(n6410), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6411) );
  XNOR2_X1 U8005 ( .A(n6411), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8371) );
  AOI22_X1 U8006 ( .A1(n6460), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n6655), .B2(
        n8371), .ZN(n6412) );
  NAND2_X1 U8007 ( .A1(n6414), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n6415) );
  NAND2_X1 U8008 ( .A1(n6426), .A2(n6415), .ZN(n7901) );
  NAND2_X1 U8009 ( .A1(n6540), .A2(n7901), .ZN(n6419) );
  INV_X1 U8010 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n10433) );
  OR2_X1 U8011 ( .A1(n6543), .A2(n10433), .ZN(n6418) );
  INV_X1 U8012 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n8355) );
  OR2_X1 U8013 ( .A1(n4517), .A2(n8355), .ZN(n6417) );
  INV_X1 U8014 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n8356) );
  OR2_X1 U8015 ( .A1(n4507), .A2(n8356), .ZN(n6416) );
  NAND4_X1 U8016 ( .A1(n6419), .A2(n6418), .A3(n6417), .A4(n6416), .ZN(n8619)
         );
  NAND2_X1 U8017 ( .A1(n8682), .A2(n8619), .ZN(n7896) );
  NOR2_X1 U8018 ( .A1(n8682), .A2(n8619), .ZN(n7898) );
  NAND2_X1 U8019 ( .A1(n7070), .A2(n6203), .ZN(n6425) );
  INV_X1 U8020 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n6420) );
  NAND2_X1 U8021 ( .A1(n6421), .A2(n6420), .ZN(n6446) );
  NAND2_X1 U8022 ( .A1(n6446), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6422) );
  NAND2_X1 U8023 ( .A1(n6423), .A2(n6422), .ZN(n6434) );
  XNOR2_X1 U8024 ( .A(n6434), .B(n6447), .ZN(n8402) );
  AOI22_X1 U8025 ( .A1(n6460), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n6655), .B2(
        n8402), .ZN(n6424) );
  NAND2_X1 U8026 ( .A1(n6426), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n6427) );
  NAND2_X1 U8027 ( .A1(n6438), .A2(n6427), .ZN(n8625) );
  NAND2_X1 U8028 ( .A1(n6540), .A2(n8625), .ZN(n6431) );
  INV_X1 U8029 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n8677) );
  OR2_X1 U8030 ( .A1(n4517), .A2(n8677), .ZN(n6430) );
  INV_X1 U8031 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n8755) );
  OR2_X1 U8032 ( .A1(n6543), .A2(n8755), .ZN(n6429) );
  INV_X1 U8033 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8624) );
  OR2_X1 U8034 ( .A1(n4507), .A2(n8624), .ZN(n6428) );
  NAND4_X1 U8035 ( .A1(n6431), .A2(n6430), .A3(n6429), .A4(n6428), .ZN(n8608)
         );
  INV_X1 U8036 ( .A(n8608), .ZN(n7916) );
  NAND2_X1 U8037 ( .A1(n8757), .A2(n7916), .ZN(n8027) );
  NAND2_X1 U8038 ( .A1(n8024), .A2(n8027), .ZN(n8614) );
  NAND2_X1 U8039 ( .A1(n8617), .A2(n8614), .ZN(n6433) );
  NAND2_X1 U8040 ( .A1(n8757), .A2(n8608), .ZN(n6432) );
  NAND2_X1 U8041 ( .A1(n6433), .A2(n6432), .ZN(n8605) );
  NAND2_X1 U8042 ( .A1(n7159), .A2(n6203), .ZN(n6437) );
  OAI21_X1 U8043 ( .B1(n6434), .B2(P2_IR_REG_16__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n6435) );
  XNOR2_X1 U8044 ( .A(n6435), .B(P2_IR_REG_17__SCAN_IN), .ZN(n8424) );
  AOI22_X1 U8045 ( .A1(n6460), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n6655), .B2(
        n8424), .ZN(n6436) );
  NAND2_X1 U8046 ( .A1(n6438), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n6439) );
  NAND2_X1 U8047 ( .A1(n6453), .A2(n6439), .ZN(n8611) );
  NAND2_X1 U8048 ( .A1(n8611), .A2(n6540), .ZN(n6444) );
  INV_X1 U8049 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n8749) );
  OR2_X1 U8050 ( .A1(n6543), .A2(n8749), .ZN(n6441) );
  INV_X1 U8051 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n8674) );
  OR2_X1 U8052 ( .A1(n4517), .A2(n8674), .ZN(n6440) );
  AND2_X1 U8053 ( .A1(n6441), .A2(n6440), .ZN(n6443) );
  INV_X1 U8054 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n10384) );
  OR2_X1 U8055 ( .A1(n4507), .A2(n10384), .ZN(n6442) );
  NAND2_X1 U8056 ( .A1(n8750), .A2(n8595), .ZN(n8032) );
  INV_X1 U8057 ( .A(n8595), .ZN(n8621) );
  AND2_X1 U8058 ( .A1(n8750), .A2(n8621), .ZN(n6445) );
  AOI21_X2 U8059 ( .B1(n8605), .B2(n8606), .A(n6445), .ZN(n8592) );
  NAND2_X1 U8060 ( .A1(n7298), .A2(n6203), .ZN(n6452) );
  INV_X1 U8061 ( .A(n6446), .ZN(n6449) );
  INV_X1 U8062 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n6448) );
  NAND2_X1 U8063 ( .A1(n4607), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6450) );
  XNOR2_X1 U8064 ( .A(n6450), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8447) );
  AOI22_X1 U8065 ( .A1(n6460), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n6655), .B2(
        n8447), .ZN(n6451) );
  INV_X1 U8066 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n10448) );
  NAND2_X1 U8067 ( .A1(n6453), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n6454) );
  NAND2_X1 U8068 ( .A1(n6463), .A2(n6454), .ZN(n8599) );
  NAND2_X1 U8069 ( .A1(n8599), .A2(n6540), .ZN(n6456) );
  AOI22_X1 U8070 ( .A1(n6532), .A2(P2_REG1_REG_18__SCAN_IN), .B1(n6491), .B2(
        P2_REG0_REG_18__SCAN_IN), .ZN(n6455) );
  OAI211_X1 U8071 ( .C1(n4507), .C2(n10448), .A(n6456), .B(n6455), .ZN(n8607)
         );
  NAND2_X1 U8072 ( .A1(n8671), .A2(n8607), .ZN(n6457) );
  NAND2_X1 U8073 ( .A1(n7370), .A2(n6203), .ZN(n6462) );
  INV_X1 U8074 ( .A(n6551), .ZN(n6458) );
  NAND2_X1 U8075 ( .A1(n6458), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6459) );
  AOI22_X1 U8076 ( .A1(n6460), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n8444), .B2(
        n6655), .ZN(n6461) );
  NAND2_X1 U8077 ( .A1(n6463), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n6464) );
  NAND2_X1 U8078 ( .A1(n6470), .A2(n6464), .ZN(n8583) );
  NAND2_X1 U8079 ( .A1(n8583), .A2(n6540), .ZN(n6467) );
  AOI22_X1 U8080 ( .A1(n6532), .A2(P2_REG1_REG_19__SCAN_IN), .B1(n6491), .B2(
        P2_REG0_REG_19__SCAN_IN), .ZN(n6466) );
  NAND2_X1 U8081 ( .A1(n6542), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n6465) );
  NAND2_X1 U8082 ( .A1(n8666), .A2(n8597), .ZN(n8036) );
  NAND2_X1 U8083 ( .A1(n8035), .A2(n8036), .ZN(n8576) );
  INV_X1 U8084 ( .A(n8597), .ZN(n8569) );
  NAND2_X1 U8085 ( .A1(n7511), .A2(n6203), .ZN(n6469) );
  OR2_X1 U8086 ( .A1(n8075), .A2(n7512), .ZN(n6468) );
  NAND2_X1 U8087 ( .A1(n6470), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n6471) );
  NAND2_X1 U8088 ( .A1(n6480), .A2(n6471), .ZN(n8566) );
  NAND2_X1 U8089 ( .A1(n8566), .A2(n6540), .ZN(n6476) );
  INV_X1 U8090 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n10432) );
  NAND2_X1 U8091 ( .A1(n6532), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n6473) );
  NAND2_X1 U8092 ( .A1(n6542), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n6472) );
  OAI211_X1 U8093 ( .C1(n6543), .C2(n10432), .A(n6473), .B(n6472), .ZN(n6474)
         );
  INV_X1 U8094 ( .A(n6474), .ZN(n6475) );
  NAND2_X1 U8095 ( .A1(n6476), .A2(n6475), .ZN(n8580) );
  NAND2_X1 U8096 ( .A1(n8736), .A2(n8554), .ZN(n8043) );
  NAND2_X1 U8097 ( .A1(n8039), .A2(n8043), .ZN(n8568) );
  NAND2_X1 U8098 ( .A1(n7527), .A2(n6203), .ZN(n6479) );
  OR2_X1 U8099 ( .A1(n8075), .A2(n7528), .ZN(n6478) );
  NAND2_X1 U8100 ( .A1(n6480), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n6481) );
  NAND2_X1 U8101 ( .A1(n6489), .A2(n6481), .ZN(n8558) );
  INV_X1 U8102 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n6484) );
  NAND2_X1 U8103 ( .A1(n6532), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n6483) );
  NAND2_X1 U8104 ( .A1(n6491), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n6482) );
  OAI211_X1 U8105 ( .C1(n6484), .C2(n4507), .A(n6483), .B(n6482), .ZN(n6485)
         );
  AOI21_X1 U8106 ( .B1(n8558), .B2(n6540), .A(n6485), .ZN(n8306) );
  NAND2_X1 U8107 ( .A1(n8175), .A2(n8306), .ZN(n8045) );
  NAND2_X1 U8108 ( .A1(n8048), .A2(n8045), .ZN(n8110) );
  NAND2_X1 U8109 ( .A1(n7686), .A2(n6203), .ZN(n6488) );
  OR2_X1 U8110 ( .A1(n8075), .A2(n7690), .ZN(n6487) );
  NAND2_X1 U8111 ( .A1(n6489), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6490) );
  NAND2_X1 U8112 ( .A1(n6499), .A2(n6490), .ZN(n8543) );
  NAND2_X1 U8113 ( .A1(n8543), .A2(n6540), .ZN(n6496) );
  INV_X1 U8114 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n8544) );
  NAND2_X1 U8115 ( .A1(n6491), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n6493) );
  INV_X1 U8116 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n10279) );
  OR2_X1 U8117 ( .A1(n4517), .A2(n10279), .ZN(n6492) );
  OAI211_X1 U8118 ( .C1(n4507), .C2(n8544), .A(n6493), .B(n6492), .ZN(n6494)
         );
  INV_X1 U8119 ( .A(n6494), .ZN(n6495) );
  NAND2_X1 U8120 ( .A1(n7750), .A2(n6203), .ZN(n6498) );
  OR2_X1 U8121 ( .A1(n8075), .A2(n7748), .ZN(n6497) );
  NAND2_X1 U8122 ( .A1(n6499), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6500) );
  NAND2_X1 U8123 ( .A1(n6501), .A2(n6500), .ZN(n8537) );
  NAND2_X1 U8124 ( .A1(n8537), .A2(n6540), .ZN(n6506) );
  INV_X1 U8125 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n8536) );
  NAND2_X1 U8126 ( .A1(n6491), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n6503) );
  INV_X1 U8127 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n10337) );
  OR2_X1 U8128 ( .A1(n4517), .A2(n10337), .ZN(n6502) );
  OAI211_X1 U8129 ( .C1(n8536), .C2(n4507), .A(n6503), .B(n6502), .ZN(n6504)
         );
  INV_X1 U8130 ( .A(n6504), .ZN(n6505) );
  INV_X1 U8131 ( .A(n8725), .ZN(n8220) );
  AOI21_X1 U8132 ( .B1(n8242), .B2(n8524), .A(n6507), .ZN(n8508) );
  OR2_X1 U8133 ( .A1(n8075), .A2(n8785), .ZN(n6508) );
  NAND2_X1 U8134 ( .A1(n6510), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n6511) );
  NAND2_X1 U8135 ( .A1(n6519), .A2(n6511), .ZN(n8511) );
  NAND2_X1 U8136 ( .A1(n8511), .A2(n6540), .ZN(n6516) );
  INV_X1 U8137 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n8516) );
  NAND2_X1 U8138 ( .A1(n6532), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n6513) );
  NAND2_X1 U8139 ( .A1(n6491), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n6512) );
  OAI211_X1 U8140 ( .C1(n8516), .C2(n4507), .A(n6513), .B(n6512), .ZN(n6514)
         );
  INV_X1 U8141 ( .A(n6514), .ZN(n6515) );
  NAND2_X1 U8142 ( .A1(n8781), .A2(n6203), .ZN(n6518) );
  OR2_X1 U8143 ( .A1(n8075), .A2(n8782), .ZN(n6517) );
  NAND2_X1 U8144 ( .A1(n6519), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n6520) );
  NAND2_X1 U8145 ( .A1(n6521), .A2(n6520), .ZN(n8505) );
  NAND2_X1 U8146 ( .A1(n8505), .A2(n6540), .ZN(n6526) );
  INV_X1 U8147 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n8504) );
  NAND2_X1 U8148 ( .A1(n6532), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n6523) );
  NAND2_X1 U8149 ( .A1(n6491), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n6522) );
  OAI211_X1 U8150 ( .C1(n8504), .C2(n4507), .A(n6523), .B(n6522), .ZN(n6524)
         );
  INV_X1 U8151 ( .A(n6524), .ZN(n6525) );
  NOR2_X1 U8152 ( .A1(n8708), .A2(n8509), .ZN(n6527) );
  NAND2_X1 U8153 ( .A1(n9728), .A2(n6203), .ZN(n6529) );
  OR2_X1 U8154 ( .A1(n8075), .A2(n8777), .ZN(n6528) );
  INV_X1 U8155 ( .A(n8635), .ZN(n8488) );
  NAND2_X1 U8156 ( .A1(n6530), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n6531) );
  NAND2_X1 U8157 ( .A1(n7921), .A2(n6531), .ZN(n8486) );
  NAND2_X1 U8158 ( .A1(n8486), .A2(n6540), .ZN(n6537) );
  INV_X1 U8159 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n10396) );
  NAND2_X1 U8160 ( .A1(n6532), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n6534) );
  NAND2_X1 U8161 ( .A1(n6542), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n6533) );
  OAI211_X1 U8162 ( .C1(n6543), .C2(n10396), .A(n6534), .B(n6533), .ZN(n6535)
         );
  INV_X1 U8163 ( .A(n6535), .ZN(n6536) );
  INV_X1 U8164 ( .A(n8494), .ZN(n8085) );
  NAND2_X1 U8165 ( .A1(n8488), .A2(n8085), .ZN(n6538) );
  OR2_X1 U8166 ( .A1(n8075), .A2(n8160), .ZN(n6539) );
  INV_X1 U8167 ( .A(n7921), .ZN(n6541) );
  NAND2_X1 U8168 ( .A1(n6541), .A2(n6540), .ZN(n7331) );
  INV_X1 U8169 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n10301) );
  NAND2_X1 U8170 ( .A1(n6542), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n6545) );
  INV_X1 U8171 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n10277) );
  OR2_X1 U8172 ( .A1(n6543), .A2(n10277), .ZN(n6544) );
  OAI211_X1 U8173 ( .C1(n10301), .C2(n4517), .A(n6545), .B(n6544), .ZN(n6546)
         );
  INV_X1 U8174 ( .A(n6546), .ZN(n6547) );
  NAND2_X1 U8175 ( .A1(n7331), .A2(n6547), .ZN(n8478) );
  INV_X1 U8176 ( .A(n8478), .ZN(n6548) );
  NAND2_X1 U8177 ( .A1(n6632), .A2(n6548), .ZN(n8084) );
  XNOR2_X1 U8178 ( .A(n6549), .B(n8105), .ZN(n6560) );
  NAND2_X1 U8179 ( .A1(n6551), .A2(n6550), .ZN(n6552) );
  NAND2_X1 U8180 ( .A1(n6552), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6555) );
  INV_X1 U8181 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n6554) );
  NAND2_X1 U8182 ( .A1(n6555), .A2(n6554), .ZN(n6557) );
  OR2_X1 U8183 ( .A1(n6555), .A2(n6554), .ZN(n6556) );
  NAND2_X1 U8184 ( .A1(n6888), .A2(n8145), .ZN(n6559) );
  NAND2_X1 U8185 ( .A1(n4580), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6558) );
  XNOR2_X1 U8186 ( .A(n6558), .B(P2_IR_REG_22__SCAN_IN), .ZN(n8155) );
  NAND2_X1 U8187 ( .A1(n8444), .A2(n8155), .ZN(n6644) );
  NAND2_X1 U8188 ( .A1(n6560), .A2(n8623), .ZN(n6592) );
  INV_X1 U8189 ( .A(n7209), .ZN(n6916) );
  AND2_X1 U8190 ( .A1(n6689), .A2(n6916), .ZN(n6866) );
  NAND2_X1 U8191 ( .A1(n6868), .A2(n7949), .ZN(n6982) );
  NAND2_X1 U8192 ( .A1(n6982), .A2(n6981), .ZN(n6563) );
  OR2_X1 U8193 ( .A1(n8318), .A2(n6968), .ZN(n7956) );
  NAND2_X1 U8194 ( .A1(n6563), .A2(n7956), .ZN(n7302) );
  XNOR2_X1 U8195 ( .A(n7953), .B(n6996), .ZN(n8114) );
  NAND2_X1 U8196 ( .A1(n7302), .A2(n8114), .ZN(n6564) );
  NAND2_X1 U8197 ( .A1(n7953), .A2(n10109), .ZN(n7969) );
  NAND2_X1 U8198 ( .A1(n6564), .A2(n7969), .ZN(n7374) );
  OR2_X1 U8199 ( .A1(n7123), .A2(n10117), .ZN(n7971) );
  NAND2_X1 U8200 ( .A1(n7374), .A2(n7971), .ZN(n6565) );
  NAND2_X1 U8201 ( .A1(n7123), .A2(n10117), .ZN(n7963) );
  NAND2_X1 U8202 ( .A1(n6565), .A2(n7963), .ZN(n7120) );
  NAND2_X1 U8203 ( .A1(n8316), .A2(n7307), .ZN(n7970) );
  OR2_X1 U8204 ( .A1(n10120), .A2(n8315), .ZN(n7965) );
  OR2_X1 U8205 ( .A1(n8316), .A2(n7307), .ZN(n7286) );
  NAND2_X1 U8206 ( .A1(n10120), .A2(n8315), .ZN(n7974) );
  AND2_X1 U8207 ( .A1(n7979), .A2(n7394), .ZN(n7984) );
  NAND2_X1 U8208 ( .A1(n7983), .A2(n7987), .ZN(n7448) );
  NOR2_X1 U8209 ( .A1(n10146), .A2(n7426), .ZN(n7982) );
  NAND2_X1 U8210 ( .A1(n10146), .A2(n7426), .ZN(n7993) );
  INV_X1 U8211 ( .A(n8124), .ZN(n7666) );
  NAND2_X1 U8212 ( .A1(n7663), .A2(n7997), .ZN(n7672) );
  INV_X1 U8213 ( .A(n7672), .ZN(n6568) );
  INV_X1 U8214 ( .A(n8309), .ZN(n7999) );
  XNOR2_X1 U8215 ( .A(n8000), .B(n7999), .ZN(n8125) );
  INV_X1 U8216 ( .A(n8125), .ZN(n6567) );
  OR2_X1 U8217 ( .A1(n8000), .A2(n7999), .ZN(n8001) );
  NAND2_X1 U8218 ( .A1(n8005), .A2(n7734), .ZN(n6569) );
  INV_X1 U8219 ( .A(n8307), .ZN(n7721) );
  AND2_X1 U8220 ( .A1(n7887), .A2(n7721), .ZN(n7877) );
  OR2_X1 U8221 ( .A1(n7887), .A2(n7721), .ZN(n8013) );
  INV_X1 U8222 ( .A(n8619), .ZN(n7841) );
  NOR2_X1 U8223 ( .A1(n8682), .A2(n7841), .ZN(n8015) );
  NAND2_X1 U8224 ( .A1(n8682), .A2(n7841), .ZN(n8017) );
  NAND2_X1 U8225 ( .A1(n6571), .A2(n8017), .ZN(n8615) );
  INV_X1 U8226 ( .A(n8027), .ZN(n8020) );
  OAI21_X1 U8227 ( .B1(n8615), .B2(n8020), .A(n8024), .ZN(n8604) );
  INV_X1 U8228 ( .A(n8025), .ZN(n6572) );
  INV_X1 U8229 ( .A(n8607), .ZN(n8225) );
  NAND2_X1 U8230 ( .A1(n8671), .A2(n8225), .ZN(n8033) );
  NAND2_X1 U8231 ( .A1(n8034), .A2(n8033), .ZN(n8591) );
  INV_X1 U8232 ( .A(n8035), .ZN(n6573) );
  NAND2_X1 U8233 ( .A1(n8565), .A2(n8039), .ZN(n6574) );
  NAND2_X1 U8234 ( .A1(n6574), .A2(n8043), .ZN(n8557) );
  INV_X1 U8235 ( .A(n8045), .ZN(n6575) );
  INV_X1 U8236 ( .A(n8533), .ZN(n8555) );
  OR2_X1 U8237 ( .A1(n8547), .A2(n8555), .ZN(n8047) );
  NOR2_X1 U8238 ( .A1(n8725), .A2(n8272), .ZN(n8109) );
  NAND2_X1 U8239 ( .A1(n8725), .A2(n8272), .ZN(n8051) );
  INV_X1 U8240 ( .A(n8060), .ZN(n6576) );
  NAND2_X1 U8241 ( .A1(n8702), .A2(n8200), .ZN(n8067) );
  NAND2_X1 U8242 ( .A1(n8635), .A2(n8085), .ZN(n6577) );
  XNOR2_X2 U8243 ( .A(n8094), .B(n8105), .ZN(n7927) );
  INV_X1 U8244 ( .A(n8155), .ZN(n7688) );
  NAND2_X1 U8245 ( .A1(n8145), .A2(n7688), .ZN(n6578) );
  NAND2_X1 U8246 ( .A1(n6578), .A2(n8463), .ZN(n6579) );
  NOR2_X1 U8247 ( .A1(n10147), .A2(n6579), .ZN(n6580) );
  NAND2_X2 U8248 ( .A1(n6888), .A2(n8155), .ZN(n8087) );
  NAND2_X1 U8249 ( .A1(n7513), .A2(n8463), .ZN(n6890) );
  OR2_X1 U8250 ( .A1(n8087), .A2(n6890), .ZN(n7201) );
  INV_X1 U8251 ( .A(n6581), .ZN(n8151) );
  XNOR2_X1 U8252 ( .A(n8151), .B(n8450), .ZN(n6902) );
  OR2_X1 U8253 ( .A1(n8087), .A2(n6902), .ZN(n8596) );
  INV_X1 U8254 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n8476) );
  NAND2_X1 U8255 ( .A1(n6491), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n6584) );
  INV_X1 U8256 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n8634) );
  OR2_X1 U8257 ( .A1(n4517), .A2(n8634), .ZN(n6583) );
  OAI211_X1 U8258 ( .C1(n4507), .C2(n8476), .A(n6584), .B(n6583), .ZN(n6585)
         );
  INV_X1 U8259 ( .A(n6585), .ZN(n6586) );
  NAND2_X1 U8260 ( .A1(n7331), .A2(n6586), .ZN(n8305) );
  INV_X1 U8261 ( .A(n6902), .ZN(n6907) );
  AND2_X1 U8262 ( .A1(n6587), .A2(P2_B_REG_SCAN_IN), .ZN(n6588) );
  NOR2_X1 U8263 ( .A1(n8598), .A2(n6588), .ZN(n8469) );
  AOI22_X1 U8264 ( .A1(n8618), .A2(n8494), .B1(n8305), .B2(n8469), .ZN(n6589)
         );
  OAI21_X1 U8265 ( .B1(n7927), .B2(n7520), .A(n6589), .ZN(n6590) );
  INV_X1 U8266 ( .A(n6590), .ZN(n6591) );
  INV_X1 U8267 ( .A(n6990), .ZN(n10141) );
  NAND2_X1 U8268 ( .A1(n6990), .A2(n7529), .ZN(n6905) );
  NAND2_X1 U8269 ( .A1(n6618), .A2(n6617), .ZN(n6594) );
  NAND2_X1 U8270 ( .A1(n6598), .A2(n6597), .ZN(n6600) );
  NAND2_X1 U8271 ( .A1(n6600), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6596) );
  OR2_X1 U8272 ( .A1(n6598), .A2(n6597), .ZN(n6599) );
  XNOR2_X1 U8273 ( .A(n8166), .B(P2_B_REG_SCAN_IN), .ZN(n6601) );
  NAND2_X1 U8274 ( .A1(n8786), .A2(n6601), .ZN(n6606) );
  NAND2_X1 U8275 ( .A1(n6602), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6603) );
  MUX2_X1 U8276 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6603), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n6604) );
  AND2_X1 U8277 ( .A1(n6605), .A2(n6604), .ZN(n6607) );
  INV_X1 U8278 ( .A(n6607), .ZN(n8783) );
  NAND2_X1 U8279 ( .A1(n8166), .A2(n8783), .ZN(n6692) );
  INV_X1 U8280 ( .A(n6886), .ZN(n7199) );
  NAND2_X1 U8281 ( .A1(n6905), .A2(n7199), .ZN(n6609) );
  NAND3_X1 U8282 ( .A1(n8145), .A2(n8155), .A3(n8463), .ZN(n6608) );
  NAND2_X1 U8283 ( .A1(n6609), .A2(n7198), .ZN(n6614) );
  INV_X1 U8284 ( .A(n7198), .ZN(n6612) );
  OR2_X1 U8285 ( .A1(n6674), .A2(P2_D_REG_1__SCAN_IN), .ZN(n6611) );
  NAND2_X1 U8286 ( .A1(n8786), .A2(n8783), .ZN(n6610) );
  NAND2_X1 U8287 ( .A1(n6611), .A2(n6610), .ZN(n7195) );
  NAND2_X1 U8288 ( .A1(n6612), .A2(n7195), .ZN(n6613) );
  AND2_X1 U8289 ( .A1(n6614), .A2(n6613), .ZN(n6631) );
  INV_X1 U8290 ( .A(n6890), .ZN(n8091) );
  OR2_X1 U8291 ( .A1(n8087), .A2(n8091), .ZN(n6877) );
  INV_X1 U8292 ( .A(n8786), .ZN(n6616) );
  NOR2_X1 U8293 ( .A1(n8166), .A2(n8783), .ZN(n6615) );
  NAND2_X1 U8294 ( .A1(n6616), .A2(n6615), .ZN(n6876) );
  XNOR2_X1 U8295 ( .A(n6618), .B(n6617), .ZN(n6875) );
  AND2_X1 U8296 ( .A1(n6875), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6694) );
  NAND2_X1 U8297 ( .A1(n6876), .A2(n6694), .ZN(n6904) );
  INV_X1 U8298 ( .A(n6904), .ZN(n6675) );
  NOR2_X1 U8299 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .ZN(
        n6622) );
  NOR4_X1 U8300 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_15__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n6621) );
  NOR4_X1 U8301 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_31__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n6620) );
  NOR4_X1 U8302 ( .A1(P2_D_REG_24__SCAN_IN), .A2(P2_D_REG_9__SCAN_IN), .A3(
        P2_D_REG_17__SCAN_IN), .A4(P2_D_REG_27__SCAN_IN), .ZN(n6619) );
  NAND4_X1 U8303 ( .A1(n6622), .A2(n6621), .A3(n6620), .A4(n6619), .ZN(n6628)
         );
  NOR4_X1 U8304 ( .A1(P2_D_REG_23__SCAN_IN), .A2(P2_D_REG_18__SCAN_IN), .A3(
        P2_D_REG_14__SCAN_IN), .A4(P2_D_REG_13__SCAN_IN), .ZN(n6626) );
  NOR4_X1 U8305 ( .A1(P2_D_REG_28__SCAN_IN), .A2(P2_D_REG_25__SCAN_IN), .A3(
        P2_D_REG_26__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n6625) );
  NOR4_X1 U8306 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n6624) );
  NOR4_X1 U8307 ( .A1(P2_D_REG_21__SCAN_IN), .A2(P2_D_REG_8__SCAN_IN), .A3(
        P2_D_REG_10__SCAN_IN), .A4(P2_D_REG_19__SCAN_IN), .ZN(n6623) );
  NAND4_X1 U8308 ( .A1(n6626), .A2(n6625), .A3(n6624), .A4(n6623), .ZN(n6627)
         );
  NOR2_X1 U8309 ( .A1(n6628), .A2(n6627), .ZN(n6629) );
  OR2_X1 U8310 ( .A1(n6674), .A2(n6629), .ZN(n6647) );
  AND2_X1 U8311 ( .A1(n6675), .A2(n6647), .ZN(n6630) );
  OR2_X1 U8312 ( .A1(n6886), .A2(n7195), .ZN(n6641) );
  AND2_X2 U8313 ( .A1(n6631), .A2(n7197), .ZN(n10159) );
  NAND2_X1 U8314 ( .A1(n10159), .A2(n10147), .ZN(n8662) );
  NAND2_X1 U8315 ( .A1(n10157), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n6633) );
  OAI21_X1 U8316 ( .B1(n6652), .B2(n10157), .A(n5136), .ZN(P2_U3488) );
  INV_X1 U8317 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n6636) );
  OAI21_X1 U8318 ( .B1(n6640), .B2(n9916), .A(n6639), .ZN(P1_U3551) );
  INV_X1 U8319 ( .A(n6641), .ZN(n6642) );
  NAND2_X1 U8320 ( .A1(n6642), .A2(n6647), .ZN(n6873) );
  INV_X1 U8321 ( .A(n6873), .ZN(n6643) );
  NAND2_X1 U8322 ( .A1(n6643), .A2(n6675), .ZN(n6903) );
  NOR2_X1 U8323 ( .A1(n6644), .A2(n7513), .ZN(n6645) );
  AND2_X1 U8324 ( .A1(n7529), .A2(n6645), .ZN(n6896) );
  INV_X1 U8325 ( .A(n6896), .ZN(n6880) );
  AND2_X1 U8326 ( .A1(n6880), .A2(n7201), .ZN(n6646) );
  OR2_X1 U8327 ( .A1(n6903), .A2(n6646), .ZN(n6649) );
  NAND3_X1 U8328 ( .A1(n6886), .A2(n7195), .A3(n6647), .ZN(n6883) );
  OR2_X1 U8329 ( .A1(n6883), .A2(n6904), .ZN(n6901) );
  INV_X1 U8330 ( .A(n6901), .ZN(n6897) );
  NAND2_X1 U8331 ( .A1(n6895), .A2(n8523), .ZN(n6874) );
  NAND2_X1 U8332 ( .A1(n6897), .A2(n6874), .ZN(n6648) );
  NAND2_X1 U8333 ( .A1(n10148), .A2(n10147), .ZN(n8733) );
  NOR2_X1 U8334 ( .A1(n10148), .A2(n10277), .ZN(n6650) );
  OAI21_X1 U8335 ( .B1(n6652), .B2(n10149), .A(n6651), .ZN(P2_U3456) );
  INV_X1 U8336 ( .A(n6694), .ZN(n6653) );
  INV_X1 U8337 ( .A(n6875), .ZN(n7746) );
  OR2_X1 U8338 ( .A1(n8087), .A2(n7746), .ZN(n6654) );
  OR2_X1 U8339 ( .A1(n6876), .A2(n7746), .ZN(n6720) );
  NAND2_X1 U8340 ( .A1(n6654), .A2(n6720), .ZN(n6723) );
  OR2_X1 U8341 ( .A1(n6723), .A2(n6655), .ZN(n6656) );
  NAND2_X1 U8342 ( .A1(n6656), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3150) );
  NOR2_X1 U8343 ( .A1(n6657), .A2(P1_U3086), .ZN(n6658) );
  XNOR2_X1 U8344 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  AND2_X1 U8345 ( .A1(n7936), .A2(P2_U3151), .ZN(n8774) );
  INV_X2 U8346 ( .A(n8774), .ZN(n8787) );
  OAI222_X1 U8347 ( .A1(n8765), .A2(n4899), .B1(n8787), .B2(n4541), .C1(
        P2_U3151), .C2(n9935), .ZN(P2_U3294) );
  OAI222_X1 U8348 ( .A1(n8765), .A2(n6659), .B1(n8787), .B2(n6665), .C1(
        P2_U3151), .C2(n6760), .ZN(P2_U3293) );
  OAI222_X1 U8349 ( .A1(n8765), .A2(n6660), .B1(n8787), .B2(n6668), .C1(
        P2_U3151), .C2(n6779), .ZN(P2_U3292) );
  OAI222_X1 U8350 ( .A1(n8765), .A2(n6661), .B1(n8787), .B2(n6663), .C1(
        P2_U3151), .C2(n7780), .ZN(P2_U3291) );
  NAND2_X1 U8351 ( .A1(n6904), .A2(P2_D_REG_1__SCAN_IN), .ZN(n6662) );
  OAI21_X1 U8352 ( .B1(n7195), .B2(n6904), .A(n6662), .ZN(P2_U3377) );
  AND2_X1 U8353 ( .A1(n7936), .A2(P1_U3086), .ZN(n9722) );
  INV_X1 U8354 ( .A(n9722), .ZN(n9735) );
  NAND2_X1 U8355 ( .A1(n5011), .A2(P1_U3086), .ZN(n9730) );
  OAI222_X1 U8356 ( .A1(n9735), .A2(n6664), .B1(n9730), .B2(n6663), .C1(
        P1_U3086), .C2(n6949), .ZN(P1_U3351) );
  OAI222_X1 U8357 ( .A1(n9735), .A2(n6666), .B1(n9730), .B2(n6665), .C1(
        P1_U3086), .C2(n6931), .ZN(P1_U3353) );
  OAI222_X1 U8358 ( .A1(n9735), .A2(n6667), .B1(n9730), .B2(n4541), .C1(
        P1_U3086), .C2(n6812), .ZN(P1_U3354) );
  OAI222_X1 U8359 ( .A1(n9735), .A2(n6669), .B1(n9730), .B2(n6668), .C1(
        P1_U3086), .C2(n6815), .ZN(P1_U3352) );
  INV_X1 U8360 ( .A(n6670), .ZN(n6672) );
  OAI222_X1 U8361 ( .A1(n9735), .A2(n6671), .B1(n9730), .B2(n6672), .C1(
        P1_U3086), .C2(n9279), .ZN(P1_U3350) );
  OAI222_X1 U8362 ( .A1(n8765), .A2(n6673), .B1(n8787), .B2(n6672), .C1(
        P2_U3151), .C2(n9951), .ZN(P2_U3290) );
  AND2_X1 U8363 ( .A1(n6675), .A2(n6674), .ZN(n6691) );
  INV_X1 U8364 ( .A(P2_D_REG_22__SCAN_IN), .ZN(n10258) );
  NOR2_X1 U8365 ( .A1(n6691), .A2(n10258), .ZN(P2_U3243) );
  INV_X1 U8366 ( .A(P2_D_REG_27__SCAN_IN), .ZN(n10466) );
  NOR2_X1 U8367 ( .A1(n6691), .A2(n10466), .ZN(P2_U3238) );
  INV_X1 U8368 ( .A(P2_D_REG_20__SCAN_IN), .ZN(n6676) );
  NOR2_X1 U8369 ( .A1(n6691), .A2(n6676), .ZN(P2_U3245) );
  INV_X1 U8370 ( .A(P2_D_REG_9__SCAN_IN), .ZN(n10373) );
  NOR2_X1 U8371 ( .A1(n6691), .A2(n10373), .ZN(P2_U3256) );
  INV_X1 U8372 ( .A(P2_D_REG_24__SCAN_IN), .ZN(n10316) );
  NOR2_X1 U8373 ( .A1(n6691), .A2(n10316), .ZN(P2_U3241) );
  INV_X1 U8374 ( .A(P2_D_REG_17__SCAN_IN), .ZN(n10397) );
  NOR2_X1 U8375 ( .A1(n6691), .A2(n10397), .ZN(P2_U3248) );
  INV_X1 U8376 ( .A(P2_D_REG_15__SCAN_IN), .ZN(n10283) );
  NOR2_X1 U8377 ( .A1(n6691), .A2(n10283), .ZN(P2_U3250) );
  INV_X1 U8378 ( .A(P2_D_REG_11__SCAN_IN), .ZN(n10326) );
  NOR2_X1 U8379 ( .A1(n6691), .A2(n10326), .ZN(P2_U3254) );
  INV_X1 U8380 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6678) );
  INV_X1 U8381 ( .A(n6677), .ZN(n6680) );
  OAI222_X1 U8382 ( .A1(n8765), .A2(n6678), .B1(n8787), .B2(n6680), .C1(
        P2_U3151), .C2(n9976), .ZN(P2_U3289) );
  INV_X1 U8383 ( .A(n9730), .ZN(n7749) );
  INV_X1 U8384 ( .A(n7749), .ZN(n9738) );
  AOI22_X1 U8385 ( .A1(n9296), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n9722), .ZN(n6679) );
  OAI21_X1 U8386 ( .B1(n6680), .B2(n9738), .A(n6679), .ZN(P1_U3349) );
  INV_X1 U8387 ( .A(n6681), .ZN(n6683) );
  AOI22_X1 U8388 ( .A1(n9309), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n9722), .ZN(n6682) );
  OAI21_X1 U8389 ( .B1(n6683), .B2(n9730), .A(n6682), .ZN(P1_U3348) );
  INV_X1 U8390 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6684) );
  OAI222_X1 U8391 ( .A1(n8765), .A2(n6684), .B1(n8787), .B2(n6683), .C1(
        P2_U3151), .C2(n9989), .ZN(P2_U3288) );
  INV_X1 U8392 ( .A(n6685), .ZN(n6687) );
  AOI22_X1 U8393 ( .A1(n9321), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n9722), .ZN(n6686) );
  OAI21_X1 U8394 ( .B1(n6687), .B2(n9738), .A(n6686), .ZN(P1_U3347) );
  INV_X1 U8395 ( .A(n10004), .ZN(n7778) );
  OAI222_X1 U8396 ( .A1(n8765), .A2(n6688), .B1(n8787), .B2(n6687), .C1(
        P2_U3151), .C2(n7778), .ZN(P2_U3287) );
  NAND2_X1 U8397 ( .A1(n8428), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n6690) );
  OAI21_X1 U8398 ( .B1(n6689), .B2(n8428), .A(n6690), .ZN(P2_U3491) );
  INV_X1 U8399 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n10370) );
  INV_X1 U8400 ( .A(n6692), .ZN(n6693) );
  AOI22_X1 U8401 ( .A1(n6695), .A2(n10370), .B1(n6694), .B2(n6693), .ZN(
        P2_U3376) );
  AND2_X1 U8402 ( .A1(n6695), .A2(P2_D_REG_5__SCAN_IN), .ZN(P2_U3260) );
  AND2_X1 U8403 ( .A1(n6695), .A2(P2_D_REG_14__SCAN_IN), .ZN(P2_U3251) );
  AND2_X1 U8404 ( .A1(n6695), .A2(P2_D_REG_30__SCAN_IN), .ZN(P2_U3235) );
  AND2_X1 U8405 ( .A1(n6695), .A2(P2_D_REG_12__SCAN_IN), .ZN(P2_U3253) );
  AND2_X1 U8406 ( .A1(n6695), .A2(P2_D_REG_8__SCAN_IN), .ZN(P2_U3257) );
  AND2_X1 U8407 ( .A1(n6695), .A2(P2_D_REG_13__SCAN_IN), .ZN(P2_U3252) );
  AND2_X1 U8408 ( .A1(n6695), .A2(P2_D_REG_3__SCAN_IN), .ZN(P2_U3262) );
  AND2_X1 U8409 ( .A1(n6695), .A2(P2_D_REG_26__SCAN_IN), .ZN(P2_U3239) );
  AND2_X1 U8410 ( .A1(n6695), .A2(P2_D_REG_2__SCAN_IN), .ZN(P2_U3263) );
  AND2_X1 U8411 ( .A1(n6695), .A2(P2_D_REG_7__SCAN_IN), .ZN(P2_U3258) );
  AND2_X1 U8412 ( .A1(n6695), .A2(P2_D_REG_23__SCAN_IN), .ZN(P2_U3242) );
  AND2_X1 U8413 ( .A1(n6695), .A2(P2_D_REG_6__SCAN_IN), .ZN(P2_U3259) );
  AND2_X1 U8414 ( .A1(n6695), .A2(P2_D_REG_21__SCAN_IN), .ZN(P2_U3244) );
  AND2_X1 U8415 ( .A1(n6695), .A2(P2_D_REG_4__SCAN_IN), .ZN(P2_U3261) );
  AND2_X1 U8416 ( .A1(n6695), .A2(P2_D_REG_25__SCAN_IN), .ZN(P2_U3240) );
  AND2_X1 U8417 ( .A1(n6695), .A2(P2_D_REG_19__SCAN_IN), .ZN(P2_U3246) );
  AND2_X1 U8418 ( .A1(n6695), .A2(P2_D_REG_18__SCAN_IN), .ZN(P2_U3247) );
  AND2_X1 U8419 ( .A1(n6695), .A2(P2_D_REG_29__SCAN_IN), .ZN(P2_U3236) );
  AND2_X1 U8420 ( .A1(n6695), .A2(P2_D_REG_28__SCAN_IN), .ZN(P2_U3237) );
  AND2_X1 U8421 ( .A1(n6695), .A2(P2_D_REG_16__SCAN_IN), .ZN(P2_U3249) );
  AND2_X1 U8422 ( .A1(n6695), .A2(P2_D_REG_10__SCAN_IN), .ZN(P2_U3255) );
  AND2_X1 U8423 ( .A1(n6695), .A2(P2_D_REG_31__SCAN_IN), .ZN(P2_U3234) );
  INV_X1 U8424 ( .A(n6696), .ZN(n6703) );
  AOI22_X1 U8425 ( .A1(n6843), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n9722), .ZN(n6697) );
  OAI21_X1 U8426 ( .B1(n6703), .B2(n9738), .A(n6697), .ZN(P1_U3346) );
  NAND2_X1 U8427 ( .A1(n6698), .A2(n6700), .ZN(n6699) );
  AND2_X1 U8428 ( .A1(n6699), .A2(n8962), .ZN(n6810) );
  INV_X1 U8429 ( .A(n6810), .ZN(n6702) );
  OR2_X1 U8430 ( .A1(n6700), .A2(P1_U3086), .ZN(n9235) );
  NAND2_X1 U8431 ( .A1(n6701), .A2(n9235), .ZN(n6811) );
  AND2_X1 U8432 ( .A1(n6702), .A2(n6811), .ZN(n10566) );
  NOR2_X1 U8433 ( .A1(n10566), .A2(P1_U3973), .ZN(P1_U3085) );
  OAI222_X1 U8434 ( .A1(n8765), .A2(n6704), .B1(n8787), .B2(n6703), .C1(
        P2_U3151), .C2(n4802), .ZN(P2_U3286) );
  INV_X1 U8435 ( .A(n6705), .ZN(n6707) );
  AOI22_X1 U8436 ( .A1(n9748), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n9722), .ZN(n6706) );
  OAI21_X1 U8437 ( .B1(n6707), .B2(n9738), .A(n6706), .ZN(P1_U3345) );
  INV_X1 U8438 ( .A(n10031), .ZN(n7777) );
  OAI222_X1 U8439 ( .A1(n8787), .A2(n6707), .B1(n7777), .B2(P2_U3151), .C1(
        n10368), .C2(n8765), .ZN(P2_U3285) );
  INV_X1 U8440 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n6714) );
  INV_X1 U8441 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n9587) );
  NAND2_X1 U8442 ( .A1(n5264), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n6711) );
  INV_X1 U8443 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n6708) );
  OR2_X1 U8444 ( .A1(n6709), .A2(n6708), .ZN(n6710) );
  OAI211_X1 U8445 ( .C1(n6712), .C2(n9587), .A(n6711), .B(n6710), .ZN(n9335)
         );
  NAND2_X1 U8446 ( .A1(n9335), .A2(P1_U3973), .ZN(n6713) );
  OAI21_X1 U8447 ( .B1(P1_U3973), .B2(n6714), .A(n6713), .ZN(P1_U3585) );
  NAND2_X1 U8448 ( .A1(n7074), .A2(P1_U3973), .ZN(n6715) );
  OAI21_X1 U8449 ( .B1(P1_U3973), .B2(n6222), .A(n6715), .ZN(P1_U3554) );
  INV_X1 U8450 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n8770) );
  INV_X1 U8451 ( .A(n9101), .ZN(n6716) );
  NAND2_X1 U8452 ( .A1(n6716), .A2(P1_U3973), .ZN(n6717) );
  OAI21_X1 U8453 ( .B1(n8770), .B2(P1_U3973), .A(n6717), .ZN(P1_U3584) );
  INV_X1 U8454 ( .A(n6718), .ZN(n6771) );
  AOI22_X1 U8455 ( .A1(n9787), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n9722), .ZN(n6719) );
  OAI21_X1 U8456 ( .B1(n6771), .B2(n9730), .A(n6719), .ZN(P1_U3344) );
  INV_X1 U8457 ( .A(n6720), .ZN(n6736) );
  NOR2_X1 U8459 ( .A1(n6723), .A2(n8779), .ZN(n6721) );
  MUX2_X1 U8460 ( .A(n6736), .B(n6721), .S(n6581), .Z(n6722) );
  NAND2_X1 U8461 ( .A1(n6722), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10051) );
  OR2_X1 U8462 ( .A1(n6581), .A2(P2_U3151), .ZN(n8775) );
  OR2_X1 U8463 ( .A1(n6723), .A2(n8775), .ZN(n9919) );
  INV_X1 U8464 ( .A(n10089), .ZN(n9969) );
  XNOR2_X1 U8465 ( .A(n6760), .B(n6724), .ZN(n6728) );
  AND2_X1 U8466 ( .A1(n6729), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6725) );
  NAND2_X1 U8467 ( .A1(n6213), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6726) );
  OAI21_X1 U8468 ( .B1(n9935), .B2(n6725), .A(n6726), .ZN(n9925) );
  NAND2_X1 U8469 ( .A1(n9927), .A2(n6726), .ZN(n6727) );
  NAND2_X1 U8470 ( .A1(n6728), .A2(n6727), .ZN(n6762) );
  OAI21_X1 U8471 ( .B1(n6728), .B2(n6727), .A(n6762), .ZN(n6740) );
  OR2_X1 U8472 ( .A1(n9919), .A2(n8450), .ZN(n9939) );
  NAND2_X1 U8473 ( .A1(n6213), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6733) );
  NAND2_X1 U8474 ( .A1(n9935), .A2(n6733), .ZN(n6732) );
  NAND2_X1 U8475 ( .A1(n6729), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6730) );
  OR2_X1 U8476 ( .A1(n6730), .A2(n6213), .ZN(n6731) );
  NAND2_X1 U8477 ( .A1(n6732), .A2(n6731), .ZN(n9937) );
  NAND2_X1 U8478 ( .A1(n9937), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n6734) );
  NAND2_X1 U8479 ( .A1(n6734), .A2(n6733), .ZN(n6755) );
  INV_X1 U8480 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n6992) );
  XNOR2_X1 U8481 ( .A(n6760), .B(n6992), .ZN(n6756) );
  XOR2_X1 U8482 ( .A(n6755), .B(n6756), .Z(n6735) );
  OAI22_X1 U8483 ( .A1(n9939), .A2(n6735), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6228), .ZN(n6739) );
  OR2_X1 U8484 ( .A1(P2_U3150), .A2(n6736), .ZN(n10049) );
  INV_X1 U8485 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n6737) );
  NOR2_X1 U8486 ( .A1(n10049), .A2(n6737), .ZN(n6738) );
  AOI211_X1 U8487 ( .C1(n9969), .C2(n6740), .A(n6739), .B(n6738), .ZN(n6748)
         );
  MUX2_X1 U8488 ( .A(P2_REG2_REG_1__SCAN_IN), .B(P2_REG1_REG_1__SCAN_IN), .S(
        n8779), .Z(n6741) );
  INV_X1 U8489 ( .A(n6741), .ZN(n6743) );
  XNOR2_X1 U8490 ( .A(n6741), .B(n6744), .ZN(n9932) );
  MUX2_X1 U8491 ( .A(n7207), .B(n6742), .S(n8779), .Z(n9920) );
  NAND2_X1 U8492 ( .A1(n9920), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n9931) );
  NAND2_X1 U8493 ( .A1(n9932), .A2(n9931), .ZN(n9930) );
  OAI21_X1 U8494 ( .B1(n6744), .B2(n6743), .A(n9930), .ZN(n6746) );
  MUX2_X1 U8495 ( .A(P2_REG2_REG_2__SCAN_IN), .B(P2_REG1_REG_2__SCAN_IN), .S(
        n8779), .Z(n6749) );
  XOR2_X1 U8496 ( .A(n6760), .B(n6749), .Z(n6745) );
  NAND2_X1 U8497 ( .A1(n6746), .A2(n6745), .ZN(n6750) );
  OR2_X1 U8498 ( .A1(n8428), .A2(n8151), .ZN(n10079) );
  INV_X1 U8499 ( .A(n10079), .ZN(n10058) );
  OAI211_X1 U8500 ( .C1(n6746), .C2(n6745), .A(n6750), .B(n10058), .ZN(n6747)
         );
  OAI211_X1 U8501 ( .C1(n10051), .C2(n6760), .A(n6748), .B(n6747), .ZN(
        P2_U3184) );
  MUX2_X1 U8502 ( .A(P2_REG2_REG_3__SCAN_IN), .B(P2_REG1_REG_3__SCAN_IN), .S(
        n8779), .Z(n6772) );
  XNOR2_X1 U8503 ( .A(n6772), .B(n6779), .ZN(n6754) );
  INV_X1 U8504 ( .A(n6760), .ZN(n6752) );
  INV_X1 U8505 ( .A(n6749), .ZN(n6751) );
  OAI21_X1 U8506 ( .B1(n6752), .B2(n6751), .A(n6750), .ZN(n6753) );
  NOR2_X1 U8507 ( .A1(n6753), .A2(n6754), .ZN(n6773) );
  AOI21_X1 U8508 ( .B1(n6754), .B2(n6753), .A(n6773), .ZN(n6770) );
  INV_X1 U8509 ( .A(n10049), .ZN(n10067) );
  NAND2_X1 U8510 ( .A1(n6756), .A2(n6755), .ZN(n6758) );
  NAND2_X1 U8511 ( .A1(n6760), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6757) );
  NAND2_X1 U8512 ( .A1(n6758), .A2(n6757), .ZN(n6780) );
  XNOR2_X1 U8513 ( .A(n6780), .B(n4799), .ZN(n6778) );
  INV_X1 U8514 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n10150) );
  XNOR2_X1 U8515 ( .A(n6778), .B(n10150), .ZN(n6759) );
  NAND2_X1 U8516 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_U3151), .ZN(n6994) );
  OAI21_X1 U8517 ( .B1(n9939), .B2(n6759), .A(n6994), .ZN(n6767) );
  NAND2_X1 U8518 ( .A1(n6760), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6761) );
  NAND2_X1 U8519 ( .A1(n6764), .A2(n6240), .ZN(n6765) );
  AOI21_X1 U8520 ( .B1(n6786), .B2(n6765), .A(n10089), .ZN(n6766) );
  AOI211_X1 U8521 ( .C1(P2_ADDR_REG_3__SCAN_IN), .C2(n10067), .A(n6767), .B(
        n6766), .ZN(n6769) );
  NAND2_X1 U8522 ( .A1(n10069), .A2(n4799), .ZN(n6768) );
  OAI211_X1 U8523 ( .C1(n6770), .C2(n10079), .A(n6769), .B(n6768), .ZN(
        P2_U3185) );
  INV_X1 U8524 ( .A(n7819), .ZN(n10050) );
  OAI222_X1 U8525 ( .A1(n8765), .A2(n10268), .B1(n8787), .B2(n6771), .C1(
        P2_U3151), .C2(n10050), .ZN(P2_U3284) );
  INV_X1 U8526 ( .A(n6772), .ZN(n6774) );
  AOI21_X1 U8527 ( .B1(n4799), .B2(n6774), .A(n6773), .ZN(n6776) );
  MUX2_X1 U8528 ( .A(P2_REG2_REG_4__SCAN_IN), .B(P2_REG1_REG_4__SCAN_IN), .S(
        n8779), .Z(n7801) );
  XOR2_X1 U8529 ( .A(n7780), .B(n7801), .Z(n6775) );
  NAND2_X1 U8530 ( .A1(n6776), .A2(n6775), .ZN(n7802) );
  OAI211_X1 U8531 ( .C1(n6776), .C2(n6775), .A(n7802), .B(n10058), .ZN(n6795)
         );
  INV_X1 U8532 ( .A(n7780), .ZN(n7804) );
  INV_X1 U8533 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n6792) );
  MUX2_X1 U8534 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n6777), .S(n7780), .Z(n6784)
         );
  NAND2_X1 U8535 ( .A1(n6778), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6782) );
  NAND2_X1 U8536 ( .A1(n6780), .A2(n6779), .ZN(n6781) );
  NAND2_X1 U8537 ( .A1(n6782), .A2(n6781), .ZN(n6783) );
  NAND2_X1 U8538 ( .A1(n6783), .A2(n6784), .ZN(n7782) );
  OAI21_X1 U8539 ( .B1(n6784), .B2(n6783), .A(n7782), .ZN(n6785) );
  AND2_X1 U8540 ( .A1(P2_U3151), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n7018) );
  AOI21_X1 U8541 ( .B1(n10084), .B2(n6785), .A(n7018), .ZN(n6791) );
  MUX2_X1 U8542 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n7377), .S(n7780), .Z(n6788)
         );
  NAND2_X1 U8543 ( .A1(n6787), .A2(n6788), .ZN(n7761) );
  OAI21_X1 U8544 ( .B1(n6788), .B2(n6787), .A(n7761), .ZN(n6789) );
  NAND2_X1 U8545 ( .A1(n9969), .A2(n6789), .ZN(n6790) );
  OAI211_X1 U8546 ( .C1(n6792), .C2(n10049), .A(n6791), .B(n6790), .ZN(n6793)
         );
  AOI21_X1 U8547 ( .B1(n7804), .B2(n10069), .A(n6793), .ZN(n6794) );
  NAND2_X1 U8548 ( .A1(n6795), .A2(n6794), .ZN(P2_U3186) );
  XNOR2_X1 U8549 ( .A(n6843), .B(P1_REG1_REG_9__SCAN_IN), .ZN(n6809) );
  INV_X1 U8550 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n9912) );
  MUX2_X1 U8551 ( .A(n9912), .B(P1_REG1_REG_2__SCAN_IN), .S(n6931), .Z(n6927)
         );
  XNOR2_X1 U8552 ( .A(n6812), .B(P1_REG1_REG_1__SCAN_IN), .ZN(n10565) );
  AND2_X1 U8553 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n10564) );
  NAND2_X1 U8554 ( .A1(n10565), .A2(n10564), .ZN(n10562) );
  INV_X1 U8555 ( .A(n6812), .ZN(n10567) );
  NAND2_X1 U8556 ( .A1(n10567), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6796) );
  NAND2_X1 U8557 ( .A1(n10562), .A2(n6796), .ZN(n6926) );
  NAND2_X1 U8558 ( .A1(n6927), .A2(n6926), .ZN(n6925) );
  OR2_X1 U8559 ( .A1(n6931), .A2(n9912), .ZN(n6797) );
  NAND2_X1 U8560 ( .A1(n6925), .A2(n6797), .ZN(n9271) );
  XNOR2_X1 U8561 ( .A(n6815), .B(P1_REG1_REG_3__SCAN_IN), .ZN(n9272) );
  NAND2_X1 U8562 ( .A1(n9271), .A2(n9272), .ZN(n9270) );
  INV_X1 U8563 ( .A(n6815), .ZN(n9269) );
  NAND2_X1 U8564 ( .A1(n9269), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6798) );
  NAND2_X1 U8565 ( .A1(n9270), .A2(n6798), .ZN(n6941) );
  XNOR2_X1 U8566 ( .A(n6949), .B(P1_REG1_REG_4__SCAN_IN), .ZN(n6942) );
  NAND2_X1 U8567 ( .A1(n6941), .A2(n6942), .ZN(n6940) );
  INV_X1 U8568 ( .A(n6949), .ZN(n6799) );
  NAND2_X1 U8569 ( .A1(n6799), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6800) );
  NAND2_X1 U8570 ( .A1(n6940), .A2(n6800), .ZN(n9285) );
  INV_X1 U8571 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n7234) );
  MUX2_X1 U8572 ( .A(n7234), .B(P1_REG1_REG_5__SCAN_IN), .S(n9279), .Z(n9286)
         );
  NAND2_X1 U8573 ( .A1(n9285), .A2(n9286), .ZN(n9284) );
  OR2_X1 U8574 ( .A1(n9279), .A2(n7234), .ZN(n6801) );
  NAND2_X1 U8575 ( .A1(n9284), .A2(n6801), .ZN(n9298) );
  INV_X1 U8576 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n10350) );
  MUX2_X1 U8577 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n10350), .S(n9296), .Z(n9299)
         );
  NAND2_X1 U8578 ( .A1(n9298), .A2(n9299), .ZN(n9297) );
  NAND2_X1 U8579 ( .A1(n9296), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6802) );
  NAND2_X1 U8580 ( .A1(n9297), .A2(n6802), .ZN(n9311) );
  INV_X1 U8581 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n6803) );
  XNOR2_X1 U8582 ( .A(n9309), .B(n6803), .ZN(n9312) );
  NAND2_X1 U8583 ( .A1(n9311), .A2(n9312), .ZN(n9310) );
  NAND2_X1 U8584 ( .A1(n9309), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6804) );
  NAND2_X1 U8585 ( .A1(n9310), .A2(n6804), .ZN(n9326) );
  XNOR2_X1 U8586 ( .A(n9321), .B(n6805), .ZN(n9327) );
  NAND2_X1 U8587 ( .A1(n9326), .A2(n9327), .ZN(n9325) );
  NAND2_X1 U8588 ( .A1(n9321), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6806) );
  NAND2_X1 U8589 ( .A1(n9325), .A2(n6806), .ZN(n6808) );
  OR2_X1 U8590 ( .A1(n6808), .A2(n6809), .ZN(n6845) );
  INV_X1 U8591 ( .A(n6845), .ZN(n6807) );
  AOI21_X1 U8592 ( .B1(n6809), .B2(n6808), .A(n6807), .ZN(n6832) );
  NAND2_X1 U8593 ( .A1(n6811), .A2(n6810), .ZN(n9777) );
  OR2_X1 U8594 ( .A1(n9777), .A2(n9774), .ZN(n9845) );
  OR2_X1 U8595 ( .A1(n9777), .A2(n6923), .ZN(n7858) );
  INV_X1 U8596 ( .A(n7858), .ZN(n10568) );
  INV_X1 U8597 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n7109) );
  MUX2_X1 U8598 ( .A(n7109), .B(P1_REG2_REG_2__SCAN_IN), .S(n6931), .Z(n6930)
         );
  XNOR2_X1 U8599 ( .A(n6812), .B(P1_REG2_REG_1__SCAN_IN), .ZN(n10561) );
  AND2_X1 U8600 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n10560) );
  NAND2_X1 U8601 ( .A1(n10561), .A2(n10560), .ZN(n10558) );
  NAND2_X1 U8602 ( .A1(n10567), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6813) );
  NAND2_X1 U8603 ( .A1(n10558), .A2(n6813), .ZN(n6929) );
  NAND2_X1 U8604 ( .A1(n6930), .A2(n6929), .ZN(n6928) );
  OR2_X1 U8605 ( .A1(n6931), .A2(n7109), .ZN(n6814) );
  NAND2_X1 U8606 ( .A1(n6928), .A2(n6814), .ZN(n9274) );
  XNOR2_X1 U8607 ( .A(n6815), .B(P1_REG2_REG_3__SCAN_IN), .ZN(n9275) );
  NAND2_X1 U8608 ( .A1(n9274), .A2(n9275), .ZN(n9273) );
  NAND2_X1 U8609 ( .A1(n9269), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6816) );
  NAND2_X1 U8610 ( .A1(n9273), .A2(n6816), .ZN(n6946) );
  XNOR2_X1 U8611 ( .A(n6949), .B(P1_REG2_REG_4__SCAN_IN), .ZN(n6947) );
  NAND2_X1 U8612 ( .A1(n6946), .A2(n6947), .ZN(n6945) );
  OR2_X1 U8613 ( .A1(n6949), .A2(n6817), .ZN(n6818) );
  NAND2_X1 U8614 ( .A1(n6945), .A2(n6818), .ZN(n9288) );
  INV_X1 U8615 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n6819) );
  MUX2_X1 U8616 ( .A(n6819), .B(P1_REG2_REG_5__SCAN_IN), .S(n9279), .Z(n9289)
         );
  NAND2_X1 U8617 ( .A1(n9288), .A2(n9289), .ZN(n9287) );
  OR2_X1 U8618 ( .A1(n9279), .A2(n6819), .ZN(n6820) );
  NAND2_X1 U8619 ( .A1(n9287), .A2(n6820), .ZN(n9301) );
  MUX2_X1 U8620 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n7247), .S(n9296), .Z(n9302)
         );
  NAND2_X1 U8621 ( .A1(n9301), .A2(n9302), .ZN(n9300) );
  NAND2_X1 U8622 ( .A1(n9296), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6821) );
  NAND2_X1 U8623 ( .A1(n9300), .A2(n6821), .ZN(n9314) );
  INV_X1 U8624 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n6822) );
  XNOR2_X1 U8625 ( .A(n9309), .B(n6822), .ZN(n9315) );
  NAND2_X1 U8626 ( .A1(n9314), .A2(n9315), .ZN(n9313) );
  NAND2_X1 U8627 ( .A1(n9309), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n6823) );
  NAND2_X1 U8628 ( .A1(n9313), .A2(n6823), .ZN(n9323) );
  INV_X1 U8629 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n7476) );
  XNOR2_X1 U8630 ( .A(n9321), .B(n7476), .ZN(n9324) );
  NAND2_X1 U8631 ( .A1(n9323), .A2(n9324), .ZN(n9322) );
  NAND2_X1 U8632 ( .A1(n9321), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6824) );
  NAND2_X1 U8633 ( .A1(n9322), .A2(n6824), .ZN(n6826) );
  XNOR2_X1 U8634 ( .A(n6843), .B(P1_REG2_REG_9__SCAN_IN), .ZN(n6825) );
  NAND2_X1 U8635 ( .A1(n6826), .A2(n6825), .ZN(n6828) );
  OR2_X1 U8636 ( .A1(n5757), .A2(n8163), .ZN(n6827) );
  OR2_X1 U8637 ( .A1(n9777), .A2(n6827), .ZN(n9832) );
  AOI21_X1 U8638 ( .B1(n6837), .B2(n6828), .A(n9832), .ZN(n6830) );
  INV_X1 U8639 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n10393) );
  NAND2_X1 U8640 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_U3086), .ZN(n7656) );
  OAI21_X1 U8641 ( .B1(n9853), .B2(n10393), .A(n7656), .ZN(n6829) );
  AOI211_X1 U8642 ( .C1(n10568), .C2(n6843), .A(n6830), .B(n6829), .ZN(n6831)
         );
  OAI21_X1 U8643 ( .B1(n6832), .B2(n9845), .A(n6831), .ZN(P1_U3252) );
  INV_X1 U8644 ( .A(n6833), .ZN(n6834) );
  INV_X1 U8645 ( .A(n10068), .ZN(n7822) );
  OAI222_X1 U8646 ( .A1(n8787), .A2(n6834), .B1(n7822), .B2(P2_U3151), .C1(
        n10382), .C2(n8765), .ZN(P2_U3283) );
  INV_X1 U8647 ( .A(n7556), .ZN(n6851) );
  OAI222_X1 U8648 ( .A1(n9735), .A2(n10457), .B1(n9730), .B2(n6834), .C1(n6851), .C2(P1_U3086), .ZN(P1_U3343) );
  NOR2_X1 U8649 ( .A1(P1_REG2_REG_12__SCAN_IN), .A2(n7556), .ZN(n6835) );
  AOI21_X1 U8650 ( .B1(n7556), .B2(P1_REG2_REG_12__SCAN_IN), .A(n6835), .ZN(
        n6841) );
  OR2_X1 U8651 ( .A1(n6843), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6836) );
  NAND2_X1 U8652 ( .A1(n6837), .A2(n6836), .ZN(n9745) );
  NAND2_X1 U8653 ( .A1(n9748), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6838) );
  OAI21_X1 U8654 ( .B1(n9748), .B2(P1_REG2_REG_10__SCAN_IN), .A(n6838), .ZN(
        n9744) );
  NOR2_X1 U8655 ( .A1(n9745), .A2(n9744), .ZN(n9747) );
  AOI21_X1 U8656 ( .B1(P1_REG2_REG_10__SCAN_IN), .B2(n9748), .A(n9747), .ZN(
        n9781) );
  NAND2_X1 U8657 ( .A1(n9787), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6839) );
  OAI21_X1 U8658 ( .B1(n9787), .B2(P1_REG2_REG_11__SCAN_IN), .A(n6839), .ZN(
        n9780) );
  NOR2_X1 U8659 ( .A1(n9781), .A2(n9780), .ZN(n9779) );
  AOI21_X1 U8660 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n9787), .A(n9779), .ZN(
        n6840) );
  NAND2_X1 U8661 ( .A1(n6841), .A2(n6840), .ZN(n7555) );
  OAI21_X1 U8662 ( .B1(n6841), .B2(n6840), .A(n7555), .ZN(n6842) );
  NAND2_X1 U8663 ( .A1(n6842), .A2(n10559), .ZN(n6855) );
  OR2_X1 U8664 ( .A1(n6843), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6844) );
  NAND2_X1 U8665 ( .A1(n6845), .A2(n6844), .ZN(n9742) );
  MUX2_X1 U8666 ( .A(n6846), .B(P1_REG1_REG_10__SCAN_IN), .S(n9748), .Z(n9741)
         );
  NOR2_X1 U8667 ( .A1(n9742), .A2(n9741), .ZN(n9752) );
  AOI21_X1 U8668 ( .B1(P1_REG1_REG_10__SCAN_IN), .B2(n9748), .A(n9752), .ZN(
        n9784) );
  MUX2_X1 U8669 ( .A(n6847), .B(P1_REG1_REG_11__SCAN_IN), .S(n9787), .Z(n9783)
         );
  NOR2_X1 U8670 ( .A1(n9784), .A2(n9783), .ZN(n9782) );
  AOI21_X1 U8671 ( .B1(P1_REG1_REG_11__SCAN_IN), .B2(n9787), .A(n9782), .ZN(
        n6849) );
  AOI22_X1 U8672 ( .A1(P1_REG1_REG_12__SCAN_IN), .A2(n7556), .B1(n6851), .B2(
        n5421), .ZN(n6848) );
  NAND2_X1 U8673 ( .A1(n6849), .A2(n6848), .ZN(n7550) );
  OAI21_X1 U8674 ( .B1(n6849), .B2(n6848), .A(n7550), .ZN(n6853) );
  INV_X1 U8675 ( .A(n9845), .ZN(n10563) );
  NAND2_X1 U8676 ( .A1(n10566), .A2(P1_ADDR_REG_12__SCAN_IN), .ZN(n6850) );
  NAND2_X1 U8677 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n8838) );
  OAI211_X1 U8678 ( .C1(n7858), .C2(n6851), .A(n6850), .B(n8838), .ZN(n6852)
         );
  AOI21_X1 U8679 ( .B1(n6853), .B2(n10563), .A(n6852), .ZN(n6854) );
  NAND2_X1 U8680 ( .A1(n6855), .A2(n6854), .ZN(P1_U3255) );
  INV_X1 U8681 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n6859) );
  NAND2_X1 U8682 ( .A1(n7520), .A2(n10141), .ZN(n10123) );
  OR2_X1 U8683 ( .A1(n6689), .A2(n6916), .ZN(n7943) );
  INV_X1 U8684 ( .A(n7943), .ZN(n7950) );
  OR2_X1 U8685 ( .A1(n7950), .A2(n6866), .ZN(n8112) );
  OAI21_X1 U8686 ( .B1(n8623), .B2(n10123), .A(n8112), .ZN(n6857) );
  NOR2_X1 U8687 ( .A1(n6224), .A2(n8598), .ZN(n7204) );
  INV_X1 U8688 ( .A(n7204), .ZN(n6856) );
  OAI211_X1 U8689 ( .C1(n7209), .C2(n10119), .A(n6857), .B(n6856), .ZN(n8690)
         );
  NAND2_X1 U8690 ( .A1(n8690), .A2(n10148), .ZN(n6858) );
  OAI21_X1 U8691 ( .B1(n6859), .B2(n10148), .A(n6858), .ZN(P2_U3390) );
  NAND2_X1 U8692 ( .A1(n8847), .A2(P1_U3973), .ZN(n6860) );
  OAI21_X1 U8693 ( .B1(n6204), .B2(P1_U3973), .A(n6860), .ZN(P1_U3578) );
  NAND2_X1 U8694 ( .A1(n8318), .A2(n8620), .ZN(n6863) );
  OAI21_X1 U8695 ( .B1(n6689), .B2(n8596), .A(n6863), .ZN(n6864) );
  AOI21_X1 U8696 ( .B1(n6865), .B2(n8623), .A(n6864), .ZN(n6870) );
  NAND2_X1 U8697 ( .A1(n6868), .A2(n6867), .ZN(n7224) );
  INV_X1 U8698 ( .A(n7520), .ZN(n6983) );
  NAND2_X1 U8699 ( .A1(n7224), .A2(n6983), .ZN(n6869) );
  AND2_X1 U8700 ( .A1(n6870), .A2(n6869), .ZN(n7226) );
  AOI22_X1 U8701 ( .A1(n7224), .A2(n6990), .B1(n10147), .B2(n4509), .ZN(n6871)
         );
  AND2_X1 U8702 ( .A1(n7226), .A2(n6871), .ZN(n10106) );
  MUX2_X1 U8703 ( .A(n10106), .B(n10467), .S(n10157), .Z(n6872) );
  INV_X1 U8704 ( .A(n6872), .ZN(P2_U3460) );
  INV_X1 U8705 ( .A(n6883), .ZN(n6881) );
  NAND2_X1 U8706 ( .A1(n6874), .A2(n6873), .ZN(n6879) );
  AND3_X1 U8707 ( .A1(n6877), .A2(n6876), .A3(n6875), .ZN(n6878) );
  OAI211_X1 U8708 ( .C1(n6881), .C2(n6880), .A(n6879), .B(n6878), .ZN(n6882)
         );
  NAND2_X1 U8709 ( .A1(n6882), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6885) );
  NOR2_X1 U8710 ( .A1(n7201), .A2(n6904), .ZN(n8152) );
  NAND2_X1 U8711 ( .A1(n8152), .A2(n6883), .ZN(n6884) );
  NAND2_X1 U8712 ( .A1(n6885), .A2(n6884), .ZN(n8295) );
  INV_X1 U8713 ( .A(n8295), .ZN(n8252) );
  NAND2_X1 U8714 ( .A1(n8252), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6971) );
  INV_X1 U8715 ( .A(n6971), .ZN(n6913) );
  NAND2_X1 U8716 ( .A1(n6887), .A2(n8145), .ZN(n6892) );
  OAI21_X1 U8717 ( .B1(n6894), .B2(n6893), .A(n6967), .ZN(n6900) );
  OR2_X1 U8718 ( .A1(n6903), .A2(n6895), .ZN(n6899) );
  NAND2_X1 U8719 ( .A1(n6897), .A2(n6896), .ZN(n6898) );
  NAND2_X1 U8720 ( .A1(n6900), .A2(n8205), .ZN(n6911) );
  NOR2_X1 U8721 ( .A1(n6901), .A2(n7201), .ZN(n6908) );
  OR2_X1 U8722 ( .A1(n6903), .A2(n10119), .ZN(n6906) );
  NAND2_X1 U8723 ( .A1(n6906), .A2(n10097), .ZN(n8263) );
  NAND2_X1 U8724 ( .A1(n6908), .A2(n6907), .ZN(n8297) );
  OAI22_X1 U8725 ( .A1(n8303), .A2(n6225), .B1(n6689), .B2(n8297), .ZN(n6909)
         );
  AOI21_X1 U8726 ( .B1(n8300), .B2(n8318), .A(n6909), .ZN(n6910) );
  OAI211_X1 U8727 ( .C1(n6913), .C2(n6912), .A(n6911), .B(n6910), .ZN(P2_U3162) );
  INV_X1 U8728 ( .A(n6914), .ZN(n6962) );
  AOI22_X1 U8729 ( .A1(n9799), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n9722), .ZN(n6915) );
  OAI21_X1 U8730 ( .B1(n6962), .B2(n9730), .A(n6915), .ZN(P1_U3342) );
  INV_X1 U8731 ( .A(n8300), .ZN(n8286) );
  AOI22_X1 U8732 ( .A1(n8205), .A2(n8112), .B1(n6916), .B2(n8263), .ZN(n6918)
         );
  NAND2_X1 U8733 ( .A1(n6971), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n6917) );
  OAI211_X1 U8734 ( .C1(n6224), .C2(n8286), .A(n6918), .B(n6917), .ZN(P2_U3172) );
  XNOR2_X1 U8735 ( .A(n6920), .B(n6919), .ZN(n6980) );
  MUX2_X1 U8736 ( .A(n6980), .B(n10560), .S(n9774), .Z(n6924) );
  AOI21_X1 U8737 ( .B1(n9774), .B2(n6921), .A(n5757), .ZN(n9773) );
  OAI21_X1 U8738 ( .B1(P1_IR_REG_0__SCAN_IN), .B2(n9773), .A(P1_U3973), .ZN(
        n6922) );
  AOI21_X1 U8739 ( .B1(n6924), .B2(n6923), .A(n6922), .ZN(n6952) );
  OAI211_X1 U8740 ( .C1(n6927), .C2(n6926), .A(n10563), .B(n6925), .ZN(n6936)
         );
  OAI211_X1 U8741 ( .C1(n6930), .C2(n6929), .A(n10559), .B(n6928), .ZN(n6935)
         );
  AOI22_X1 U8742 ( .A1(n10566), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n6934) );
  INV_X1 U8743 ( .A(n6931), .ZN(n6932) );
  NAND2_X1 U8744 ( .A1(n10568), .A2(n6932), .ZN(n6933) );
  NAND4_X1 U8745 ( .A1(n6936), .A2(n6935), .A3(n6934), .A4(n6933), .ZN(n6937)
         );
  OR2_X1 U8746 ( .A1(n6952), .A2(n6937), .ZN(P1_U3245) );
  INV_X1 U8747 ( .A(P1_U3973), .ZN(n9265) );
  NAND2_X1 U8748 ( .A1(n9265), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n6938) );
  OAI21_X1 U8749 ( .B1(n6939), .B2(n9265), .A(n6938), .ZN(P1_U3583) );
  INV_X1 U8750 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n6944) );
  OAI211_X1 U8751 ( .C1(n6942), .C2(n6941), .A(n10563), .B(n6940), .ZN(n6943)
         );
  NAND2_X1 U8752 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_U3086), .ZN(n7053) );
  OAI211_X1 U8753 ( .C1(n9853), .C2(n6944), .A(n6943), .B(n7053), .ZN(n6951)
         );
  OAI211_X1 U8754 ( .C1(n6947), .C2(n6946), .A(n10559), .B(n6945), .ZN(n6948)
         );
  OAI21_X1 U8755 ( .B1(n7858), .B2(n6949), .A(n6948), .ZN(n6950) );
  OR3_X1 U8756 ( .A1(n6952), .A2(n6951), .A3(n6950), .ZN(P1_U3247) );
  AND2_X1 U8757 ( .A1(n9772), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7037) );
  OAI21_X1 U8758 ( .B1(n6954), .B2(n6953), .A(n7025), .ZN(n6955) );
  NAND2_X1 U8759 ( .A1(n6955), .A2(n8942), .ZN(n6960) );
  INV_X1 U8760 ( .A(n5852), .ZN(n6957) );
  INV_X1 U8761 ( .A(n7074), .ZN(n6956) );
  OAI22_X1 U8762 ( .A1(n6957), .A2(n8946), .B1(n6956), .B2(n8944), .ZN(n7064)
         );
  AOI22_X1 U8763 ( .A1(n8958), .A2(n6958), .B1(n9764), .B2(n7064), .ZN(n6959)
         );
  OAI211_X1 U8764 ( .C1(n7037), .C2(n6961), .A(n6960), .B(n6959), .ZN(P1_U3222) );
  INV_X1 U8765 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6963) );
  INV_X1 U8766 ( .A(n8321), .ZN(n8325) );
  OAI222_X1 U8767 ( .A1(n8765), .A2(n6963), .B1(n8787), .B2(n6962), .C1(
        P2_U3151), .C2(n8325), .ZN(P2_U3282) );
  INV_X1 U8768 ( .A(n6964), .ZN(n6965) );
  NAND2_X1 U8769 ( .A1(n6965), .A2(n6224), .ZN(n6966) );
  NAND2_X1 U8770 ( .A1(n6967), .A2(n6966), .ZN(n6998) );
  XNOR2_X1 U8771 ( .A(n8189), .B(n7954), .ZN(n6999) );
  XNOR2_X1 U8772 ( .A(n6999), .B(n8318), .ZN(n6997) );
  XOR2_X1 U8773 ( .A(n6998), .B(n6997), .Z(n6973) );
  NOR2_X1 U8774 ( .A1(n8286), .A2(n7953), .ZN(n6970) );
  OAI22_X1 U8775 ( .A1(n8303), .A2(n6968), .B1(n6224), .B2(n8297), .ZN(n6969)
         );
  AOI211_X1 U8776 ( .C1(P2_REG3_REG_2__SCAN_IN), .C2(n6971), .A(n6970), .B(
        n6969), .ZN(n6972) );
  OAI21_X1 U8777 ( .B1(n6973), .B2(n8267), .A(n6972), .ZN(P2_U3177) );
  INV_X1 U8778 ( .A(n6974), .ZN(n7008) );
  AOI22_X1 U8779 ( .A1(n9811), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n9722), .ZN(n6975) );
  OAI21_X1 U8780 ( .B1(n7008), .B2(n9738), .A(n6975), .ZN(P1_U3341) );
  AND2_X1 U8781 ( .A1(n5840), .A2(n8932), .ZN(n7133) );
  AOI22_X1 U8782 ( .A1(n8958), .A2(n6976), .B1(n9764), .B2(n7133), .ZN(n6979)
         );
  INV_X1 U8783 ( .A(n7037), .ZN(n6977) );
  NAND2_X1 U8784 ( .A1(n6977), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n6978) );
  OAI211_X1 U8785 ( .C1(n6980), .C2(n9758), .A(n6979), .B(n6978), .ZN(P1_U3232) );
  XNOR2_X1 U8786 ( .A(n6982), .B(n6981), .ZN(n10101) );
  NAND2_X1 U8787 ( .A1(n10101), .A2(n6983), .ZN(n6989) );
  OAI21_X1 U8788 ( .B1(n8111), .B2(n6984), .A(n6985), .ZN(n6987) );
  OAI22_X1 U8789 ( .A1(n6224), .A2(n8596), .B1(n7953), .B2(n8598), .ZN(n6986)
         );
  AOI21_X1 U8790 ( .B1(n6987), .B2(n8623), .A(n6986), .ZN(n6988) );
  AND2_X1 U8791 ( .A1(n6989), .A2(n6988), .ZN(n10098) );
  AND2_X1 U8792 ( .A1(n7954), .A2(n10147), .ZN(n10095) );
  AOI21_X1 U8793 ( .B1(n10101), .B2(n6990), .A(n10095), .ZN(n6991) );
  AND2_X1 U8794 ( .A1(n10098), .A2(n6991), .ZN(n10108) );
  MUX2_X1 U8795 ( .A(n6992), .B(n10108), .S(n10159), .Z(n6993) );
  INV_X1 U8796 ( .A(n6993), .ZN(P2_U3461) );
  INV_X1 U8797 ( .A(n8297), .ZN(n8284) );
  AOI22_X1 U8798 ( .A1(n8284), .A2(n8318), .B1(n8300), .B2(n6267), .ZN(n6995)
         );
  OAI211_X1 U8799 ( .C1(n6996), .C2(n8303), .A(n6995), .B(n6994), .ZN(n7006)
         );
  XNOR2_X1 U8800 ( .A(n8189), .B(n10109), .ZN(n7010) );
  XNOR2_X1 U8801 ( .A(n7010), .B(n7953), .ZN(n7004) );
  NAND2_X1 U8802 ( .A1(n6998), .A2(n6997), .ZN(n7001) );
  INV_X1 U8803 ( .A(n8318), .ZN(n7955) );
  NAND2_X1 U8804 ( .A1(n6999), .A2(n7955), .ZN(n7000) );
  INV_X1 U8805 ( .A(n7013), .ZN(n7002) );
  AOI211_X1 U8806 ( .C1(n7004), .C2(n7003), .A(n8267), .B(n7002), .ZN(n7005)
         );
  AOI211_X1 U8807 ( .C1(n6161), .C2(n8295), .A(n7006), .B(n7005), .ZN(n7007)
         );
  INV_X1 U8808 ( .A(n7007), .ZN(P2_U3158) );
  INV_X1 U8809 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n7009) );
  INV_X1 U8810 ( .A(n8350), .ZN(n8347) );
  OAI222_X1 U8811 ( .A1(n8765), .A2(n7009), .B1(n8787), .B2(n7008), .C1(
        P2_U3151), .C2(n8347), .ZN(P2_U3281) );
  XNOR2_X1 U8812 ( .A(n8189), .B(n10117), .ZN(n7042) );
  XNOR2_X1 U8813 ( .A(n7042), .B(n7123), .ZN(n7016) );
  INV_X1 U8814 ( .A(n7010), .ZN(n7011) );
  INV_X1 U8815 ( .A(n7953), .ZN(n8317) );
  NAND2_X1 U8816 ( .A1(n7011), .A2(n8317), .ZN(n7012) );
  INV_X1 U8817 ( .A(n7086), .ZN(n7014) );
  AOI21_X1 U8818 ( .B1(n7016), .B2(n7015), .A(n7014), .ZN(n7022) );
  INV_X1 U8819 ( .A(n8316), .ZN(n7079) );
  OAI22_X1 U8820 ( .A1(n8286), .A2(n7079), .B1(n7953), .B2(n8297), .ZN(n7017)
         );
  AOI211_X1 U8821 ( .C1(n10117), .C2(n8263), .A(n7018), .B(n7017), .ZN(n7021)
         );
  INV_X1 U8822 ( .A(n7019), .ZN(n7378) );
  NAND2_X1 U8823 ( .A1(n8295), .A2(n7378), .ZN(n7020) );
  OAI211_X1 U8824 ( .C1(n7022), .C2(n8267), .A(n7021), .B(n7020), .ZN(P2_U3170) );
  NAND2_X1 U8825 ( .A1(n9265), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n7023) );
  OAI21_X1 U8826 ( .B1(n7024), .B2(n9265), .A(n7023), .ZN(P1_U3582) );
  INV_X1 U8827 ( .A(n7025), .ZN(n7029) );
  INV_X1 U8828 ( .A(n7026), .ZN(n7028) );
  NOR3_X1 U8829 ( .A1(n7029), .A2(n7028), .A3(n7027), .ZN(n7032) );
  INV_X1 U8830 ( .A(n7030), .ZN(n7031) );
  OAI21_X1 U8831 ( .B1(n7032), .B2(n7031), .A(n8942), .ZN(n7036) );
  NAND2_X1 U8832 ( .A1(n9264), .A2(n8932), .ZN(n7034) );
  NAND2_X1 U8833 ( .A1(n5840), .A2(n9232), .ZN(n7033) );
  NAND2_X1 U8834 ( .A1(n7034), .A2(n7033), .ZN(n7114) );
  AOI22_X1 U8835 ( .A1(n8958), .A2(n7112), .B1(n9764), .B2(n7114), .ZN(n7035)
         );
  OAI211_X1 U8836 ( .C1(n7037), .C2(n7108), .A(n7036), .B(n7035), .ZN(P1_U3237) );
  INV_X1 U8837 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n7039) );
  INV_X1 U8838 ( .A(n7038), .ZN(n7040) );
  INV_X1 U8839 ( .A(n8371), .ZN(n8377) );
  OAI222_X1 U8840 ( .A1(n8765), .A2(n7039), .B1(n8787), .B2(n7040), .C1(
        P2_U3151), .C2(n8377), .ZN(P2_U3280) );
  INV_X1 U8841 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n7041) );
  INV_X1 U8842 ( .A(n9822), .ZN(n7558) );
  OAI222_X1 U8843 ( .A1(n9735), .A2(n7041), .B1(n9738), .B2(n7040), .C1(
        P1_U3086), .C2(n7558), .ZN(P1_U3340) );
  NAND2_X1 U8844 ( .A1(n7042), .A2(n7123), .ZN(n7081) );
  NAND2_X1 U8845 ( .A1(n7086), .A2(n7081), .ZN(n7173) );
  XNOR2_X1 U8846 ( .A(n8189), .B(n7125), .ZN(n7080) );
  XNOR2_X1 U8847 ( .A(n7080), .B(n8316), .ZN(n7172) );
  XNOR2_X1 U8848 ( .A(n7173), .B(n7172), .ZN(n7046) );
  AOI22_X1 U8849 ( .A1(n8300), .A2(n8315), .B1(n8263), .B2(n7125), .ZN(n7044)
         );
  AND2_X1 U8850 ( .A1(P2_U3151), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n9948) );
  AOI21_X1 U8851 ( .B1(n8284), .B2(n6267), .A(n9948), .ZN(n7043) );
  OAI211_X1 U8852 ( .C1(n8252), .C2(n7306), .A(n7044), .B(n7043), .ZN(n7045)
         );
  AOI21_X1 U8853 ( .B1(n7046), .B2(n8205), .A(n7045), .ZN(n7047) );
  INV_X1 U8854 ( .A(n7047), .ZN(P2_U3167) );
  NAND2_X1 U8855 ( .A1(n4510), .A2(n8942), .ZN(n7058) );
  AOI21_X1 U8856 ( .B1(n7048), .B2(n7050), .A(n7049), .ZN(n7057) );
  INV_X1 U8857 ( .A(n9262), .ZN(n7052) );
  INV_X1 U8858 ( .A(n9264), .ZN(n7051) );
  OAI22_X1 U8859 ( .A1(n7052), .A2(n8946), .B1(n7051), .B2(n8944), .ZN(n7153)
         );
  INV_X1 U8860 ( .A(n7053), .ZN(n7055) );
  OAI22_X1 U8861 ( .A1(n9766), .A2(n8974), .B1(n9772), .B2(n9854), .ZN(n7054)
         );
  AOI211_X1 U8862 ( .C1(n9764), .C2(n7153), .A(n7055), .B(n7054), .ZN(n7056)
         );
  OAI21_X1 U8863 ( .B1(n7058), .B2(n7057), .A(n7056), .ZN(P1_U3230) );
  INV_X1 U8864 ( .A(n9659), .ZN(n7728) );
  XNOR2_X1 U8865 ( .A(n7059), .B(n7060), .ZN(n7062) );
  INV_X1 U8866 ( .A(n7062), .ZN(n9879) );
  INV_X1 U8867 ( .A(n9656), .ZN(n9905) );
  OAI211_X1 U8868 ( .C1(n7138), .C2(n9872), .A(n7872), .B(n7105), .ZN(n9875)
         );
  OAI21_X1 U8869 ( .B1(n9872), .B2(n9905), .A(n9875), .ZN(n7067) );
  OAI21_X1 U8870 ( .B1(n7059), .B2(n7075), .A(n7061), .ZN(n7065) );
  NOR2_X1 U8871 ( .A1(n7062), .A2(n9564), .ZN(n7063) );
  AOI211_X1 U8872 ( .C1(n9549), .C2(n7065), .A(n7064), .B(n7063), .ZN(n9882)
         );
  INV_X1 U8873 ( .A(n9882), .ZN(n7066) );
  AOI211_X1 U8874 ( .C1(n7728), .C2(n9879), .A(n7067), .B(n7066), .ZN(n9886)
         );
  NAND2_X1 U8875 ( .A1(n9916), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n7068) );
  OAI21_X1 U8876 ( .B1(n9886), .B2(n9916), .A(n7068), .ZN(P1_U3523) );
  NAND2_X1 U8877 ( .A1(n8534), .A2(P2_U3893), .ZN(n7069) );
  OAI21_X1 U8878 ( .B1(P2_U3893), .B2(n5647), .A(n7069), .ZN(P2_U3515) );
  INV_X1 U8879 ( .A(n9837), .ZN(n7554) );
  INV_X1 U8880 ( .A(n7070), .ZN(n7072) );
  INV_X1 U8881 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n7071) );
  OAI222_X1 U8882 ( .A1(P1_U3086), .A2(n7554), .B1(n9738), .B2(n7072), .C1(
        n7071), .C2(n9735), .ZN(P1_U3339) );
  INV_X1 U8883 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n7073) );
  INV_X1 U8884 ( .A(n8402), .ZN(n8399) );
  OAI222_X1 U8885 ( .A1(n8765), .A2(n7073), .B1(P2_U3151), .B2(n8399), .C1(
        n7072), .C2(n8787), .ZN(P2_U3279) );
  AND2_X1 U8886 ( .A1(n7074), .A2(n7138), .ZN(n9149) );
  OR2_X1 U8887 ( .A1(n9149), .A2(n7075), .ZN(n9106) );
  OAI21_X1 U8888 ( .B1(n9549), .B2(n9908), .A(n9106), .ZN(n7077) );
  INV_X1 U8889 ( .A(n7133), .ZN(n7076) );
  OAI211_X1 U8890 ( .C1(n7138), .C2(n7132), .A(n7077), .B(n7076), .ZN(n9661)
         );
  NAND2_X1 U8891 ( .A1(n9661), .A2(n9911), .ZN(n7078) );
  OAI21_X1 U8892 ( .B1(n9911), .B2(n5189), .A(n7078), .ZN(P1_U3453) );
  NAND2_X1 U8893 ( .A1(n7080), .A2(n7079), .ZN(n7174) );
  AND2_X1 U8894 ( .A1(n7081), .A2(n7082), .ZN(n7085) );
  INV_X1 U8895 ( .A(n7082), .ZN(n7083) );
  XNOR2_X1 U8896 ( .A(n10128), .B(n8189), .ZN(n7162) );
  XNOR2_X1 U8897 ( .A(n7162), .B(n8314), .ZN(n7087) );
  OAI21_X1 U8898 ( .B1(n7088), .B2(n7087), .A(n7424), .ZN(n7095) );
  AND2_X1 U8899 ( .A1(P2_U3151), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n9987) );
  AOI21_X1 U8900 ( .B1(n8284), .B2(n8315), .A(n9987), .ZN(n7093) );
  NAND2_X1 U8901 ( .A1(n8263), .A2(n10128), .ZN(n7092) );
  INV_X1 U8902 ( .A(n7321), .ZN(n7089) );
  NAND2_X1 U8903 ( .A1(n8295), .A2(n7089), .ZN(n7091) );
  NAND2_X1 U8904 ( .A1(n8300), .A2(n8313), .ZN(n7090) );
  NAND4_X1 U8905 ( .A1(n7093), .A2(n7092), .A3(n7091), .A4(n7090), .ZN(n7094)
         );
  AOI21_X1 U8906 ( .B1(n7095), .B2(n8205), .A(n7094), .ZN(n7096) );
  INV_X1 U8907 ( .A(n7096), .ZN(P2_U3153) );
  XNOR2_X1 U8908 ( .A(n7097), .B(n9105), .ZN(n9891) );
  INV_X1 U8909 ( .A(n9891), .ZN(n7119) );
  INV_X1 U8910 ( .A(n7098), .ZN(n7101) );
  NAND3_X1 U8911 ( .A1(n7101), .A2(n7100), .A3(n7099), .ZN(n7104) );
  AND2_X1 U8912 ( .A1(n9564), .A2(n7631), .ZN(n7102) );
  OR2_X1 U8913 ( .A1(n7104), .A2(n4621), .ZN(n9859) );
  INV_X1 U8914 ( .A(n7278), .ZN(n7107) );
  AOI21_X1 U8915 ( .B1(n7112), .B2(n7105), .A(n9578), .ZN(n7106) );
  NAND2_X1 U8916 ( .A1(n7107), .A2(n7106), .ZN(n9887) );
  OAI22_X1 U8917 ( .A1(n9859), .A2(n9887), .B1(n7108), .B2(n9869), .ZN(n7111)
         );
  NOR2_X1 U8918 ( .A1(n9561), .A2(n7109), .ZN(n7110) );
  AOI211_X1 U8919 ( .C1(n9866), .C2(n7112), .A(n7111), .B(n7110), .ZN(n7118)
         );
  XNOR2_X1 U8920 ( .A(n9105), .B(n8965), .ZN(n7113) );
  NAND2_X1 U8921 ( .A1(n7113), .A2(n9549), .ZN(n7116) );
  INV_X1 U8922 ( .A(n7114), .ZN(n7115) );
  NAND2_X1 U8923 ( .A1(n7116), .A2(n7115), .ZN(n9889) );
  NAND2_X1 U8924 ( .A1(n9889), .A2(n9561), .ZN(n7117) );
  OAI211_X1 U8925 ( .C1(n7119), .C2(n9861), .A(n7118), .B(n7117), .ZN(P1_U3291) );
  XNOR2_X1 U8926 ( .A(n8316), .B(n7125), .ZN(n8115) );
  XNOR2_X1 U8927 ( .A(n7120), .B(n8115), .ZN(n7311) );
  INV_X1 U8928 ( .A(n8315), .ZN(n7124) );
  INV_X1 U8929 ( .A(n8623), .ZN(n8593) );
  XOR2_X1 U8930 ( .A(n8115), .B(n7121), .Z(n7122) );
  OAI222_X1 U8931 ( .A1(n8598), .A2(n7124), .B1(n8596), .B2(n7123), .C1(n8593), 
        .C2(n7122), .ZN(n7308) );
  AOI21_X1 U8932 ( .B1(n10123), .B2(n7311), .A(n7308), .ZN(n7130) );
  AOI22_X1 U8933 ( .A1(n8678), .A2(n7125), .B1(n10157), .B2(
        P2_REG1_REG_5__SCAN_IN), .ZN(n7126) );
  OAI21_X1 U8934 ( .B1(n7130), .B2(n10157), .A(n7126), .ZN(P2_U3464) );
  INV_X1 U8935 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n7127) );
  OAI22_X1 U8936 ( .A1(n8733), .A2(n7307), .B1(n7127), .B2(n10148), .ZN(n7128)
         );
  INV_X1 U8937 ( .A(n7128), .ZN(n7129) );
  OAI21_X1 U8938 ( .B1(n7130), .B2(n10149), .A(n7129), .ZN(P2_U3405) );
  AOI21_X1 U8939 ( .B1(n9877), .B2(n7872), .A(n9866), .ZN(n7139) );
  NAND3_X1 U8940 ( .A1(n9106), .A2(n7132), .A3(n7131), .ZN(n7135) );
  INV_X1 U8941 ( .A(n9869), .ZN(n9855) );
  AOI21_X1 U8942 ( .B1(n9855), .B2(P1_REG3_REG_0__SCAN_IN), .A(n7133), .ZN(
        n7134) );
  AOI21_X1 U8943 ( .B1(n7135), .B2(n7134), .A(n9857), .ZN(n7136) );
  AOI21_X1 U8944 ( .B1(n9857), .B2(P1_REG2_REG_0__SCAN_IN), .A(n7136), .ZN(
        n7137) );
  OAI21_X1 U8945 ( .B1(n7139), .B2(n7138), .A(n7137), .ZN(P1_U3293) );
  NAND2_X1 U8946 ( .A1(n7140), .A2(n7141), .ZN(n7143) );
  XNOR2_X1 U8947 ( .A(n7143), .B(n7142), .ZN(n7147) );
  AOI22_X1 U8948 ( .A1(n8932), .A2(n9261), .B1(n9263), .B2(n9232), .ZN(n7215)
         );
  NOR2_X1 U8949 ( .A1(n8912), .A2(n7215), .ZN(n7145) );
  OAI22_X1 U8950 ( .A1(n9766), .A2(n7409), .B1(n9772), .B2(n7220), .ZN(n7144)
         );
  AOI211_X1 U8951 ( .C1(P1_REG3_REG_5__SCAN_IN), .C2(P1_U3086), .A(n7145), .B(
        n7144), .ZN(n7146) );
  OAI21_X1 U8952 ( .B1(n7147), .B2(n9758), .A(n7146), .ZN(P1_U3227) );
  INV_X1 U8953 ( .A(n9908), .ZN(n7583) );
  INV_X1 U8954 ( .A(n7148), .ZN(n7150) );
  OR2_X1 U8955 ( .A1(n7150), .A2(n7149), .ZN(n9109) );
  XNOR2_X1 U8956 ( .A(n7151), .B(n9109), .ZN(n9862) );
  XNOR2_X1 U8957 ( .A(n7152), .B(n9109), .ZN(n7154) );
  AOI21_X1 U8958 ( .B1(n7154), .B2(n9549), .A(n7153), .ZN(n9868) );
  INV_X1 U8959 ( .A(n7277), .ZN(n7155) );
  OAI211_X1 U8960 ( .C1(n7155), .C2(n8974), .A(n7872), .B(n7218), .ZN(n9860)
         );
  OAI211_X1 U8961 ( .C1(n7583), .C2(n9862), .A(n9868), .B(n9860), .ZN(n7407)
         );
  INV_X1 U8962 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n7156) );
  OAI22_X1 U8963 ( .A1(n9652), .A2(n8974), .B1(n9918), .B2(n7156), .ZN(n7157)
         );
  AOI21_X1 U8964 ( .B1(n7407), .B2(n9918), .A(n7157), .ZN(n7158) );
  INV_X1 U8965 ( .A(n7158), .ZN(P1_U3526) );
  INV_X1 U8966 ( .A(n7159), .ZN(n7210) );
  AOI22_X1 U8967 ( .A1(n7851), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n9722), .ZN(n7160) );
  OAI21_X1 U8968 ( .B1(n7210), .B2(n9730), .A(n7160), .ZN(P1_U3338) );
  NAND2_X1 U8969 ( .A1(n7162), .A2(n7161), .ZN(n7422) );
  NAND2_X1 U8970 ( .A1(n7424), .A2(n7422), .ZN(n7381) );
  XNOR2_X1 U8971 ( .A(n10134), .B(n8189), .ZN(n7383) );
  XNOR2_X1 U8972 ( .A(n7383), .B(n8313), .ZN(n7416) );
  XNOR2_X1 U8973 ( .A(n7381), .B(n7416), .ZN(n7170) );
  NAND2_X1 U8974 ( .A1(P2_U3151), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n10014) );
  INV_X1 U8975 ( .A(n10014), .ZN(n7163) );
  AOI21_X1 U8976 ( .B1(n8284), .B2(n8314), .A(n7163), .ZN(n7168) );
  NAND2_X1 U8977 ( .A1(n10134), .A2(n8263), .ZN(n7167) );
  INV_X1 U8978 ( .A(n7402), .ZN(n7164) );
  NAND2_X1 U8979 ( .A1(n8295), .A2(n7164), .ZN(n7166) );
  NAND2_X1 U8980 ( .A1(n8300), .A2(n8312), .ZN(n7165) );
  NAND4_X1 U8981 ( .A1(n7168), .A2(n7167), .A3(n7166), .A4(n7165), .ZN(n7169)
         );
  AOI21_X1 U8982 ( .B1(n7170), .B2(n8205), .A(n7169), .ZN(n7171) );
  INV_X1 U8983 ( .A(n7171), .ZN(P2_U3161) );
  NAND2_X1 U8984 ( .A1(n7173), .A2(n7172), .ZN(n7175) );
  NAND2_X1 U8985 ( .A1(n7175), .A2(n7174), .ZN(n7176) );
  AOI211_X1 U8986 ( .C1(n7177), .C2(n7176), .A(n8267), .B(n4605), .ZN(n7186)
         );
  INV_X1 U8987 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n7178) );
  NOR2_X1 U8988 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7178), .ZN(n9967) );
  AOI21_X1 U8989 ( .B1(n8284), .B2(n8316), .A(n9967), .ZN(n7184) );
  NAND2_X1 U8990 ( .A1(n8263), .A2(n7179), .ZN(n7183) );
  INV_X1 U8991 ( .A(n7289), .ZN(n7180) );
  NAND2_X1 U8992 ( .A1(n8295), .A2(n7180), .ZN(n7182) );
  NAND2_X1 U8993 ( .A1(n8300), .A2(n8314), .ZN(n7181) );
  NAND4_X1 U8994 ( .A1(n7184), .A2(n7183), .A3(n7182), .A4(n7181), .ZN(n7185)
         );
  OR2_X1 U8995 ( .A1(n7186), .A2(n7185), .ZN(P2_U3179) );
  NAND2_X1 U8996 ( .A1(n4828), .A2(n7189), .ZN(n7190) );
  XNOR2_X1 U8997 ( .A(n7187), .B(n7190), .ZN(n7194) );
  AOI22_X1 U8998 ( .A1(n8932), .A2(n9260), .B1(n9262), .B2(n9232), .ZN(n7241)
         );
  NOR2_X1 U8999 ( .A1(n8912), .A2(n7241), .ZN(n7192) );
  OAI22_X1 U9000 ( .A1(n9766), .A2(n7353), .B1(n9772), .B2(n7246), .ZN(n7191)
         );
  AOI211_X1 U9001 ( .C1(P1_REG3_REG_6__SCAN_IN), .C2(P1_U3086), .A(n7192), .B(
        n7191), .ZN(n7193) );
  OAI21_X1 U9002 ( .B1(n7194), .B2(n9758), .A(n7193), .ZN(P1_U3239) );
  NAND2_X1 U9003 ( .A1(n7198), .A2(n7195), .ZN(n7196) );
  OAI211_X1 U9004 ( .C1(n7199), .C2(n7198), .A(n7197), .B(n7196), .ZN(n7205)
         );
  INV_X1 U9005 ( .A(n7205), .ZN(n7200) );
  INV_X1 U9006 ( .A(n8523), .ZN(n8512) );
  NAND2_X1 U9007 ( .A1(n7200), .A2(n8512), .ZN(n8560) );
  INV_X1 U9008 ( .A(n10097), .ZN(n8626) );
  INV_X1 U9009 ( .A(n7201), .ZN(n7202) );
  NOR3_X1 U9010 ( .A1(n4856), .A2(n10147), .A3(n7202), .ZN(n7203) );
  AOI211_X1 U9011 ( .C1(n8626), .C2(P2_REG3_REG_0__SCAN_IN), .A(n7204), .B(
        n7203), .ZN(n7206) );
  MUX2_X1 U9012 ( .A(n7207), .B(n7206), .S(n10103), .Z(n7208) );
  OAI21_X1 U9013 ( .B1(n8560), .B2(n7209), .A(n7208), .ZN(P2_U3233) );
  INV_X1 U9014 ( .A(n8424), .ZN(n8430) );
  OAI222_X1 U9015 ( .A1(n8765), .A2(n7211), .B1(n8787), .B2(n7210), .C1(
        P2_U3151), .C2(n8430), .ZN(P2_U3278) );
  XNOR2_X1 U9016 ( .A(n7213), .B(n7212), .ZN(n7233) );
  XNOR2_X1 U9017 ( .A(n7214), .B(n9111), .ZN(n7217) );
  INV_X1 U9018 ( .A(n7215), .ZN(n7216) );
  AOI21_X1 U9019 ( .B1(n7217), .B2(n9549), .A(n7216), .ZN(n7232) );
  MUX2_X1 U9020 ( .A(n7232), .B(n6819), .S(n9857), .Z(n7223) );
  AOI211_X1 U9021 ( .C1(n7219), .C2(n7218), .A(n9578), .B(n7243), .ZN(n7230)
         );
  OAI22_X1 U9022 ( .A1(n9873), .A2(n7409), .B1(n9869), .B2(n7220), .ZN(n7221)
         );
  AOI21_X1 U9023 ( .B1(n7230), .B2(n9877), .A(n7221), .ZN(n7222) );
  OAI211_X1 U9024 ( .C1(n9861), .C2(n7233), .A(n7223), .B(n7222), .ZN(P1_U3288) );
  INV_X1 U9025 ( .A(n7224), .ZN(n7229) );
  AND2_X1 U9026 ( .A1(n6888), .A2(n7942), .ZN(n10102) );
  NAND2_X1 U9027 ( .A1(n10103), .A2(n10102), .ZN(n7926) );
  MUX2_X1 U9028 ( .A(n7226), .B(n7225), .S(n10105), .Z(n7228) );
  AOI22_X1 U9029 ( .A1(n8627), .A2(n4509), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        n8626), .ZN(n7227) );
  OAI211_X1 U9030 ( .C1(n7229), .C2(n7926), .A(n7228), .B(n7227), .ZN(P2_U3232) );
  INV_X1 U9031 ( .A(n7230), .ZN(n7231) );
  OAI211_X1 U9032 ( .C1(n7583), .C2(n7233), .A(n7232), .B(n7231), .ZN(n7411)
         );
  OAI22_X1 U9033 ( .A1(n9652), .A2(n7409), .B1(n9918), .B2(n7234), .ZN(n7235)
         );
  AOI21_X1 U9034 ( .B1(n7411), .B2(n9918), .A(n7235), .ZN(n7236) );
  INV_X1 U9035 ( .A(n7236), .ZN(P1_U3527) );
  OAI21_X1 U9036 ( .B1(n7238), .B2(n7239), .A(n7237), .ZN(n7350) );
  INV_X1 U9037 ( .A(n7350), .ZN(n7252) );
  XNOR2_X1 U9038 ( .A(n7240), .B(n7239), .ZN(n7242) );
  OAI21_X1 U9039 ( .B1(n7242), .B2(n9571), .A(n7241), .ZN(n7348) );
  NAND2_X1 U9040 ( .A1(n7348), .A2(n9561), .ZN(n7251) );
  INV_X1 U9041 ( .A(n7353), .ZN(n7245) );
  INV_X1 U9042 ( .A(n7243), .ZN(n7244) );
  AOI211_X1 U9043 ( .C1(n7245), .C2(n7244), .A(n9578), .B(n7364), .ZN(n7349)
         );
  NOR2_X1 U9044 ( .A1(n9873), .A2(n7353), .ZN(n7249) );
  OAI22_X1 U9045 ( .A1(n9561), .A2(n7247), .B1(n7246), .B2(n9869), .ZN(n7248)
         );
  AOI211_X1 U9046 ( .C1(n7349), .C2(n9877), .A(n7249), .B(n7248), .ZN(n7250)
         );
  OAI211_X1 U9047 ( .C1(n7252), .C2(n9861), .A(n7251), .B(n7250), .ZN(P1_U3287) );
  INV_X1 U9048 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n10166) );
  INV_X1 U9049 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n10456) );
  INV_X1 U9050 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n8406) );
  AOI22_X1 U9051 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .B1(n10456), .B2(n8406), .ZN(n10171) );
  INV_X1 U9052 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n10427) );
  INV_X1 U9053 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n8384) );
  AOI22_X1 U9054 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .B1(n10427), .B2(n8384), .ZN(n10174) );
  INV_X1 U9055 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n9826) );
  INV_X1 U9056 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n8354) );
  AOI22_X1 U9057 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .B1(n9826), .B2(n8354), .ZN(n10177) );
  NOR2_X1 U9058 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n7253) );
  AOI21_X1 U9059 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n7253), .ZN(n10180) );
  NOR2_X1 U9060 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n7254) );
  AOI21_X1 U9061 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n7254), .ZN(n10183) );
  NOR2_X1 U9062 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n7255) );
  AOI21_X1 U9063 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n7255), .ZN(n10186) );
  NOR2_X1 U9064 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n7256) );
  AOI21_X1 U9065 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n7256), .ZN(n10189) );
  NOR2_X1 U9066 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n7257) );
  AOI21_X1 U9067 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n7257), .ZN(n10192) );
  NOR2_X1 U9068 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n7258) );
  AOI21_X1 U9069 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(P2_ADDR_REG_9__SCAN_IN), 
        .A(n7258), .ZN(n10586) );
  NOR2_X1 U9070 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n7259) );
  AOI21_X1 U9071 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(P2_ADDR_REG_8__SCAN_IN), 
        .A(n7259), .ZN(n10589) );
  NOR2_X1 U9072 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n7260) );
  AOI21_X1 U9073 ( .B1(P1_ADDR_REG_7__SCAN_IN), .B2(P2_ADDR_REG_7__SCAN_IN), 
        .A(n7260), .ZN(n10583) );
  NOR2_X1 U9074 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(P1_ADDR_REG_6__SCAN_IN), 
        .ZN(n7261) );
  AOI21_X1 U9075 ( .B1(P1_ADDR_REG_6__SCAN_IN), .B2(P2_ADDR_REG_6__SCAN_IN), 
        .A(n7261), .ZN(n10577) );
  NOR2_X1 U9076 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n7262) );
  AOI21_X1 U9077 ( .B1(P1_ADDR_REG_5__SCAN_IN), .B2(P2_ADDR_REG_5__SCAN_IN), 
        .A(n7262), .ZN(n10580) );
  NAND2_X1 U9078 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .ZN(n10163) );
  INV_X1 U9079 ( .A(n10163), .ZN(n7263) );
  INV_X1 U9080 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10161) );
  NAND2_X1 U9081 ( .A1(n10163), .A2(n10161), .ZN(n10160) );
  AOI22_X1 U9082 ( .A1(n7263), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P2_ADDR_REG_1__SCAN_IN), .B2(n10160), .ZN(n10592) );
  NAND2_X1 U9083 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n7264) );
  OAI21_X1 U9084 ( .B1(P1_ADDR_REG_2__SCAN_IN), .B2(P2_ADDR_REG_2__SCAN_IN), 
        .A(n7264), .ZN(n10591) );
  NOR2_X1 U9085 ( .A1(n10592), .A2(n10591), .ZN(n10590) );
  AOI21_X1 U9086 ( .B1(P2_ADDR_REG_2__SCAN_IN), .B2(P1_ADDR_REG_2__SCAN_IN), 
        .A(n10590), .ZN(n10595) );
  NAND2_X1 U9087 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n7265) );
  OAI21_X1 U9088 ( .B1(P1_ADDR_REG_3__SCAN_IN), .B2(P2_ADDR_REG_3__SCAN_IN), 
        .A(n7265), .ZN(n10594) );
  NOR2_X1 U9089 ( .A1(n10595), .A2(n10594), .ZN(n10593) );
  AOI21_X1 U9090 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(P1_ADDR_REG_3__SCAN_IN), 
        .A(n10593), .ZN(n10598) );
  NOR2_X1 U9091 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n7266) );
  AOI21_X1 U9092 ( .B1(P2_ADDR_REG_4__SCAN_IN), .B2(P1_ADDR_REG_4__SCAN_IN), 
        .A(n7266), .ZN(n10597) );
  NAND2_X1 U9093 ( .A1(n10598), .A2(n10597), .ZN(n10596) );
  OAI21_X1 U9094 ( .B1(P1_ADDR_REG_4__SCAN_IN), .B2(P2_ADDR_REG_4__SCAN_IN), 
        .A(n10596), .ZN(n10579) );
  NAND2_X1 U9095 ( .A1(n10580), .A2(n10579), .ZN(n10578) );
  OAI21_X1 U9096 ( .B1(P2_ADDR_REG_5__SCAN_IN), .B2(P1_ADDR_REG_5__SCAN_IN), 
        .A(n10578), .ZN(n10576) );
  NAND2_X1 U9097 ( .A1(n10577), .A2(n10576), .ZN(n10575) );
  OAI21_X1 U9098 ( .B1(P2_ADDR_REG_6__SCAN_IN), .B2(P1_ADDR_REG_6__SCAN_IN), 
        .A(n10575), .ZN(n10582) );
  NAND2_X1 U9099 ( .A1(n10583), .A2(n10582), .ZN(n10581) );
  OAI21_X1 U9100 ( .B1(P2_ADDR_REG_7__SCAN_IN), .B2(P1_ADDR_REG_7__SCAN_IN), 
        .A(n10581), .ZN(n10588) );
  NAND2_X1 U9101 ( .A1(n10589), .A2(n10588), .ZN(n10587) );
  OAI21_X1 U9102 ( .B1(P2_ADDR_REG_8__SCAN_IN), .B2(P1_ADDR_REG_8__SCAN_IN), 
        .A(n10587), .ZN(n10585) );
  NAND2_X1 U9103 ( .A1(n10586), .A2(n10585), .ZN(n10584) );
  OAI21_X1 U9104 ( .B1(P2_ADDR_REG_9__SCAN_IN), .B2(P1_ADDR_REG_9__SCAN_IN), 
        .A(n10584), .ZN(n10191) );
  NAND2_X1 U9105 ( .A1(n10192), .A2(n10191), .ZN(n10190) );
  OAI21_X1 U9106 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n10190), .ZN(n10188) );
  NAND2_X1 U9107 ( .A1(n10189), .A2(n10188), .ZN(n10187) );
  OAI21_X1 U9108 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n10187), .ZN(n10185) );
  NAND2_X1 U9109 ( .A1(n10186), .A2(n10185), .ZN(n10184) );
  OAI21_X1 U9110 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10184), .ZN(n10182) );
  NAND2_X1 U9111 ( .A1(n10183), .A2(n10182), .ZN(n10181) );
  OAI21_X1 U9112 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n10181), .ZN(n10179) );
  NAND2_X1 U9113 ( .A1(n10180), .A2(n10179), .ZN(n10178) );
  OAI21_X1 U9114 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10178), .ZN(n10176) );
  NAND2_X1 U9115 ( .A1(n10177), .A2(n10176), .ZN(n10175) );
  OAI21_X1 U9116 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n10175), .ZN(n10173) );
  NAND2_X1 U9117 ( .A1(n10174), .A2(n10173), .ZN(n10172) );
  OAI21_X1 U9118 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n10172), .ZN(n10170) );
  NAND2_X1 U9119 ( .A1(n10171), .A2(n10170), .ZN(n10169) );
  OAI21_X1 U9120 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10169), .ZN(n10167) );
  NOR2_X1 U9121 ( .A1(n10166), .A2(n10167), .ZN(n7267) );
  NAND2_X1 U9122 ( .A1(n10166), .A2(n10167), .ZN(n10165) );
  OAI21_X1 U9123 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(n7267), .A(n10165), .ZN(
        n7271) );
  NOR2_X1 U9124 ( .A1(n7269), .A2(n7268), .ZN(n7270) );
  XNOR2_X1 U9125 ( .A(n7271), .B(n7270), .ZN(ADD_1068_U4) );
  XOR2_X1 U9126 ( .A(n9108), .B(n9156), .Z(n7275) );
  NAND2_X1 U9127 ( .A1(n5852), .A2(n9232), .ZN(n7273) );
  NAND2_X1 U9128 ( .A1(n9263), .A2(n8932), .ZN(n7272) );
  NAND2_X1 U9129 ( .A1(n7273), .A2(n7272), .ZN(n8811) );
  INV_X1 U9130 ( .A(n8811), .ZN(n7274) );
  OAI21_X1 U9131 ( .B1(n7275), .B2(n9571), .A(n7274), .ZN(n9894) );
  INV_X1 U9132 ( .A(n9894), .ZN(n7283) );
  XNOR2_X1 U9133 ( .A(n7276), .B(n9108), .ZN(n9896) );
  OAI211_X1 U9134 ( .C1(n7278), .C2(n9893), .A(n7277), .B(n7872), .ZN(n9892)
         );
  OAI22_X1 U9135 ( .A1(n9892), .A2(n9859), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        n9869), .ZN(n7279) );
  AOI21_X1 U9136 ( .B1(P1_REG2_REG_3__SCAN_IN), .B2(n9857), .A(n7279), .ZN(
        n7280) );
  OAI21_X1 U9137 ( .B1(n9893), .B2(n9873), .A(n7280), .ZN(n7281) );
  AOI21_X1 U9138 ( .B1(n9535), .B2(n9896), .A(n7281), .ZN(n7282) );
  OAI21_X1 U9139 ( .B1(n7283), .B2(n9857), .A(n7282), .ZN(P1_U3290) );
  INV_X1 U9140 ( .A(n10102), .ZN(n7284) );
  NAND2_X1 U9141 ( .A1(n7520), .A2(n7284), .ZN(n7285) );
  NAND2_X1 U9142 ( .A1(n7287), .A2(n7286), .ZN(n7288) );
  AND2_X1 U9143 ( .A1(n7965), .A2(n7974), .ZN(n8117) );
  XNOR2_X1 U9144 ( .A(n7288), .B(n8117), .ZN(n10124) );
  OAI22_X1 U9145 ( .A1(n8560), .A2(n10120), .B1(n7289), .B2(n10097), .ZN(n7296) );
  INV_X1 U9146 ( .A(n8117), .ZN(n7291) );
  XNOR2_X1 U9147 ( .A(n7290), .B(n7291), .ZN(n7292) );
  NAND2_X1 U9148 ( .A1(n7292), .A2(n8623), .ZN(n7294) );
  AOI22_X1 U9149 ( .A1(n8618), .A2(n8316), .B1(n8314), .B2(n8620), .ZN(n7293)
         );
  NAND2_X1 U9150 ( .A1(n7294), .A2(n7293), .ZN(n10121) );
  MUX2_X1 U9151 ( .A(n10121), .B(P2_REG2_REG_6__SCAN_IN), .S(n10105), .Z(n7295) );
  AOI211_X1 U9152 ( .C1(n8562), .C2(n10124), .A(n7296), .B(n7295), .ZN(n7297)
         );
  INV_X1 U9153 ( .A(n7297), .ZN(P2_U3227) );
  INV_X1 U9154 ( .A(n7298), .ZN(n7334) );
  AOI22_X1 U9155 ( .A1(n9850), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n9722), .ZN(n7299) );
  OAI21_X1 U9156 ( .B1(n7334), .B2(n9730), .A(n7299), .ZN(P1_U3337) );
  XOR2_X1 U9157 ( .A(n7300), .B(n8114), .Z(n7301) );
  AOI222_X1 U9158 ( .A1(n8623), .A2(n7301), .B1(n6267), .B2(n8620), .C1(n8318), 
        .C2(n8618), .ZN(n10112) );
  XNOR2_X1 U9159 ( .A(n7302), .B(n8114), .ZN(n10110) );
  AOI22_X1 U9160 ( .A1(n8627), .A2(n10109), .B1(n6161), .B2(n8626), .ZN(n7303)
         );
  OAI21_X1 U9161 ( .B1(n6240), .B2(n10103), .A(n7303), .ZN(n7304) );
  AOI21_X1 U9162 ( .B1(n10110), .B2(n8562), .A(n7304), .ZN(n7305) );
  OAI21_X1 U9163 ( .B1(n10112), .B2(n10105), .A(n7305), .ZN(P2_U3230) );
  OAI22_X1 U9164 ( .A1(n8560), .A2(n7307), .B1(n7306), .B2(n10097), .ZN(n7310)
         );
  MUX2_X1 U9165 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n7308), .S(n10103), .Z(n7309)
         );
  AOI211_X1 U9166 ( .C1(n7311), .C2(n8562), .A(n7310), .B(n7309), .ZN(n7312)
         );
  INV_X1 U9167 ( .A(n7312), .ZN(P2_U3228) );
  NAND3_X1 U9168 ( .A1(n7313), .A2(n6320), .A3(n7974), .ZN(n7314) );
  NAND2_X1 U9169 ( .A1(n7395), .A2(n7314), .ZN(n10125) );
  INV_X1 U9170 ( .A(n7315), .ZN(n7317) );
  OAI21_X1 U9171 ( .B1(n7317), .B2(n6320), .A(n7316), .ZN(n7318) );
  NAND2_X1 U9172 ( .A1(n7318), .A2(n8623), .ZN(n7320) );
  AOI22_X1 U9173 ( .A1(n8620), .A2(n8313), .B1(n8315), .B2(n8618), .ZN(n7319)
         );
  OAI211_X1 U9174 ( .C1(n7520), .C2(n10125), .A(n7320), .B(n7319), .ZN(n10126)
         );
  NAND2_X1 U9175 ( .A1(n10126), .A2(n10103), .ZN(n7324) );
  OAI22_X1 U9176 ( .A1(n10103), .A2(n6312), .B1(n7321), .B2(n10097), .ZN(n7322) );
  AOI21_X1 U9177 ( .B1(n8627), .B2(n10128), .A(n7322), .ZN(n7323) );
  OAI211_X1 U9178 ( .C1(n10125), .C2(n7926), .A(n7324), .B(n7323), .ZN(
        P2_U3226) );
  INV_X1 U9179 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n7333) );
  INV_X1 U9180 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n8473) );
  NAND2_X1 U9181 ( .A1(n6491), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n7327) );
  INV_X1 U9182 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n7325) );
  OR2_X1 U9183 ( .A1(n4517), .A2(n7325), .ZN(n7326) );
  OAI211_X1 U9184 ( .C1(n8473), .C2(n4507), .A(n7327), .B(n7326), .ZN(n7329)
         );
  INV_X1 U9185 ( .A(n7329), .ZN(n7330) );
  NAND2_X1 U9186 ( .A1(n8470), .A2(P2_U3893), .ZN(n7332) );
  OAI21_X1 U9187 ( .B1(P2_U3893), .B2(n7333), .A(n7332), .ZN(P2_U3522) );
  INV_X1 U9188 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n7335) );
  INV_X1 U9189 ( .A(n8447), .ZN(n8454) );
  OAI222_X1 U9190 ( .A1(n8765), .A2(n7335), .B1(n8454), .B2(P2_U3151), .C1(
        n8787), .C2(n7334), .ZN(P2_U3277) );
  XNOR2_X1 U9191 ( .A(n7337), .B(n7336), .ZN(n7338) );
  XNOR2_X1 U9192 ( .A(n7339), .B(n7338), .ZN(n7346) );
  OR2_X1 U9193 ( .A1(n7498), .A2(n8946), .ZN(n7341) );
  NAND2_X1 U9194 ( .A1(n9261), .A2(n9232), .ZN(n7340) );
  NAND2_X1 U9195 ( .A1(n7341), .A2(n7340), .ZN(n7360) );
  AOI22_X1 U9196 ( .A1(n9764), .A2(n7360), .B1(P1_REG3_REG_7__SCAN_IN), .B2(
        P1_U3086), .ZN(n7344) );
  INV_X1 U9197 ( .A(n7342), .ZN(n7365) );
  NAND2_X1 U9198 ( .A1(n8883), .A2(n7365), .ZN(n7343) );
  OAI211_X1 U9199 ( .C1(n9898), .C2(n9766), .A(n7344), .B(n7343), .ZN(n7345)
         );
  AOI21_X1 U9200 ( .B1(n7346), .B2(n8942), .A(n7345), .ZN(n7347) );
  INV_X1 U9201 ( .A(n7347), .ZN(P1_U3213) );
  AOI211_X1 U9202 ( .C1(n9908), .C2(n7350), .A(n7349), .B(n7348), .ZN(n7356)
         );
  OAI22_X1 U9203 ( .A1(n9652), .A2(n7353), .B1(n9918), .B2(n10350), .ZN(n7351)
         );
  INV_X1 U9204 ( .A(n7351), .ZN(n7352) );
  OAI21_X1 U9205 ( .B1(n7356), .B2(n9916), .A(n7352), .ZN(P1_U3528) );
  OAI22_X1 U9206 ( .A1(n9713), .A2(n7353), .B1(n9911), .B2(n5285), .ZN(n7354)
         );
  INV_X1 U9207 ( .A(n7354), .ZN(n7355) );
  OAI21_X1 U9208 ( .B1(n7356), .B2(n9910), .A(n7355), .ZN(P1_U3471) );
  INV_X1 U9209 ( .A(n8988), .ZN(n7359) );
  NAND2_X1 U9210 ( .A1(n7358), .A2(n7359), .ZN(n7467) );
  OAI21_X1 U9211 ( .B1(n7359), .B2(n7358), .A(n7467), .ZN(n7361) );
  AOI21_X1 U9212 ( .B1(n7361), .B2(n9549), .A(n7360), .ZN(n9899) );
  OAI21_X1 U9213 ( .B1(n7363), .B2(n8988), .A(n7362), .ZN(n9902) );
  OAI211_X1 U9214 ( .C1(n7364), .C2(n9898), .A(n7872), .B(n7474), .ZN(n9897)
         );
  NOR2_X1 U9215 ( .A1(n9897), .A2(n9859), .ZN(n7368) );
  AOI22_X1 U9216 ( .A1(n9857), .A2(P1_REG2_REG_7__SCAN_IN), .B1(n7365), .B2(
        n9855), .ZN(n7366) );
  OAI21_X1 U9217 ( .B1(n9873), .B2(n9898), .A(n7366), .ZN(n7367) );
  AOI211_X1 U9218 ( .C1(n9902), .C2(n9535), .A(n7368), .B(n7367), .ZN(n7369)
         );
  OAI21_X1 U9219 ( .B1(n9899), .B2(n9857), .A(n7369), .ZN(P1_U3286) );
  INV_X1 U9220 ( .A(n7370), .ZN(n7372) );
  OAI222_X1 U9221 ( .A1(n9735), .A2(n7371), .B1(n9738), .B2(n7372), .C1(
        P1_U3086), .C2(n9230), .ZN(P1_U3336) );
  OAI222_X1 U9222 ( .A1(n8765), .A2(n7373), .B1(n8787), .B2(n7372), .C1(n8463), 
        .C2(P2_U3151), .ZN(P2_U3276) );
  NAND2_X1 U9223 ( .A1(n7971), .A2(n7963), .ZN(n8113) );
  XNOR2_X1 U9224 ( .A(n7374), .B(n8113), .ZN(n10113) );
  XNOR2_X1 U9225 ( .A(n7375), .B(n8113), .ZN(n7376) );
  AOI222_X1 U9226 ( .A1(n8623), .A2(n7376), .B1(n8317), .B2(n8618), .C1(n8316), 
        .C2(n8620), .ZN(n10114) );
  MUX2_X1 U9227 ( .A(n7377), .B(n10114), .S(n8610), .Z(n7380) );
  AOI22_X1 U9228 ( .A1(n8627), .A2(n10117), .B1(n8626), .B2(n7378), .ZN(n7379)
         );
  OAI211_X1 U9229 ( .C1(n8630), .C2(n10113), .A(n7380), .B(n7379), .ZN(
        P2_U3229) );
  XNOR2_X1 U9230 ( .A(n7418), .B(n8312), .ZN(n7413) );
  NAND2_X1 U9231 ( .A1(n7381), .A2(n7416), .ZN(n7384) );
  NAND2_X1 U9232 ( .A1(n7383), .A2(n7382), .ZN(n7414) );
  NAND2_X1 U9233 ( .A1(n7384), .A2(n7414), .ZN(n7385) );
  AOI211_X1 U9234 ( .C1(n7413), .C2(n7385), .A(n8267), .B(n4606), .ZN(n7393)
         );
  NAND2_X1 U9235 ( .A1(n10139), .A2(n8263), .ZN(n7391) );
  NAND2_X1 U9236 ( .A1(P2_U3151), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n10028) );
  INV_X1 U9237 ( .A(n10028), .ZN(n7386) );
  AOI21_X1 U9238 ( .B1(n8284), .B2(n8313), .A(n7386), .ZN(n7390) );
  INV_X1 U9239 ( .A(n7453), .ZN(n7387) );
  NAND2_X1 U9240 ( .A1(n8295), .A2(n7387), .ZN(n7389) );
  NAND2_X1 U9241 ( .A1(n8300), .A2(n8311), .ZN(n7388) );
  NAND4_X1 U9242 ( .A1(n7391), .A2(n7390), .A3(n7389), .A4(n7388), .ZN(n7392)
         );
  OR2_X1 U9243 ( .A1(n7393), .A2(n7392), .ZN(P2_U3171) );
  NAND2_X1 U9244 ( .A1(n7395), .A2(n7394), .ZN(n7396) );
  XOR2_X1 U9245 ( .A(n8118), .B(n7396), .Z(n10131) );
  NAND2_X1 U9246 ( .A1(n7397), .A2(n8623), .ZN(n7401) );
  AOI21_X1 U9247 ( .B1(n7316), .B2(n7398), .A(n8118), .ZN(n7400) );
  AOI22_X1 U9248 ( .A1(n8618), .A2(n8314), .B1(n8312), .B2(n8620), .ZN(n7399)
         );
  OAI21_X1 U9249 ( .B1(n7401), .B2(n7400), .A(n7399), .ZN(n10132) );
  NAND2_X1 U9250 ( .A1(n10132), .A2(n10103), .ZN(n7405) );
  OAI22_X1 U9251 ( .A1(n10103), .A2(n6329), .B1(n7402), .B2(n10097), .ZN(n7403) );
  AOI21_X1 U9252 ( .B1(n8627), .B2(n10134), .A(n7403), .ZN(n7404) );
  OAI211_X1 U9253 ( .C1(n10131), .C2(n8630), .A(n7405), .B(n7404), .ZN(
        P2_U3225) );
  OAI22_X1 U9254 ( .A1(n9713), .A2(n8974), .B1(n9911), .B2(n5243), .ZN(n7406)
         );
  AOI21_X1 U9255 ( .B1(n7407), .B2(n9911), .A(n7406), .ZN(n7408) );
  INV_X1 U9256 ( .A(n7408), .ZN(P1_U3465) );
  OAI22_X1 U9257 ( .A1(n9713), .A2(n7409), .B1(n9911), .B2(n5265), .ZN(n7410)
         );
  AOI21_X1 U9258 ( .B1(n7411), .B2(n9911), .A(n7410), .ZN(n7412) );
  INV_X1 U9259 ( .A(n7412), .ZN(P1_U3468) );
  XNOR2_X1 U9260 ( .A(n10146), .B(n8196), .ZN(n7436) );
  INV_X1 U9261 ( .A(n7413), .ZN(n7415) );
  AND2_X1 U9262 ( .A1(n7415), .A2(n7414), .ZN(n7421) );
  INV_X1 U9263 ( .A(n7416), .ZN(n7417) );
  NAND2_X1 U9264 ( .A1(n7418), .A2(n8312), .ZN(n7419) );
  AND2_X1 U9265 ( .A1(n7422), .A2(n7421), .ZN(n7423) );
  NAND2_X1 U9266 ( .A1(n7427), .A2(n7426), .ZN(n7437) );
  INV_X1 U9267 ( .A(n7427), .ZN(n7428) );
  NAND2_X1 U9268 ( .A1(n7437), .A2(n7438), .ZN(n7429) );
  XOR2_X1 U9269 ( .A(n7436), .B(n7429), .Z(n7435) );
  INV_X1 U9270 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n7430) );
  NOR2_X1 U9271 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7430), .ZN(n10039) );
  NOR2_X1 U9272 ( .A1(n8297), .A2(n6346), .ZN(n7431) );
  AOI211_X1 U9273 ( .C1(n8300), .C2(n8310), .A(n10039), .B(n7431), .ZN(n7432)
         );
  OAI21_X1 U9274 ( .B1(n7523), .B2(n8252), .A(n7432), .ZN(n7433) );
  AOI21_X1 U9275 ( .B1(n10146), .B2(n8263), .A(n7433), .ZN(n7434) );
  OAI21_X1 U9276 ( .B1(n7435), .B2(n8267), .A(n7434), .ZN(P2_U3157) );
  INV_X1 U9277 ( .A(n8686), .ZN(n7446) );
  XNOR2_X1 U9278 ( .A(n8124), .B(n8196), .ZN(n7457) );
  OAI211_X1 U9279 ( .C1(n7439), .C2(n7457), .A(n7459), .B(n8205), .ZN(n7445)
         );
  INV_X1 U9280 ( .A(n7440), .ZN(n7668) );
  NAND2_X1 U9281 ( .A1(P2_U3151), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n10064) );
  INV_X1 U9282 ( .A(n10064), .ZN(n7441) );
  AOI21_X1 U9283 ( .B1(n8284), .B2(n8311), .A(n7441), .ZN(n7442) );
  OAI21_X1 U9284 ( .B1(n7999), .B2(n8286), .A(n7442), .ZN(n7443) );
  AOI21_X1 U9285 ( .B1(n7668), .B2(n8295), .A(n7443), .ZN(n7444) );
  OAI211_X1 U9286 ( .C1(n7446), .C2(n8303), .A(n7445), .B(n7444), .ZN(P2_U3176) );
  XNOR2_X1 U9287 ( .A(n7447), .B(n7448), .ZN(n10136) );
  XNOR2_X1 U9288 ( .A(n7449), .B(n4860), .ZN(n7450) );
  NAND2_X1 U9289 ( .A1(n7450), .A2(n8623), .ZN(n7452) );
  AOI22_X1 U9290 ( .A1(n8311), .A2(n8620), .B1(n8618), .B2(n8313), .ZN(n7451)
         );
  OAI211_X1 U9291 ( .C1(n7520), .C2(n10136), .A(n7452), .B(n7451), .ZN(n10137)
         );
  NAND2_X1 U9292 ( .A1(n10137), .A2(n8610), .ZN(n7456) );
  OAI22_X1 U9293 ( .A1(n10103), .A2(n6341), .B1(n7453), .B2(n10097), .ZN(n7454) );
  AOI21_X1 U9294 ( .B1(n8627), .B2(n10139), .A(n7454), .ZN(n7455) );
  OAI211_X1 U9295 ( .C1(n10136), .C2(n7926), .A(n7456), .B(n7455), .ZN(
        P2_U3224) );
  NAND2_X1 U9296 ( .A1(n5067), .A2(n8310), .ZN(n7458) );
  XNOR2_X1 U9297 ( .A(n8000), .B(n8196), .ZN(n7571) );
  XNOR2_X1 U9298 ( .A(n7571), .B(n7999), .ZN(n7460) );
  XNOR2_X1 U9299 ( .A(n7572), .B(n7460), .ZN(n7465) );
  NAND2_X1 U9300 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3151), .ZN(n10091) );
  OAI21_X1 U9301 ( .B1(n8297), .B2(n7675), .A(n10091), .ZN(n7461) );
  AOI21_X1 U9302 ( .B1(n8300), .B2(n8308), .A(n7461), .ZN(n7462) );
  OAI21_X1 U9303 ( .B1(n7681), .B2(n8252), .A(n7462), .ZN(n7463) );
  AOI21_X1 U9304 ( .B1(n8000), .B2(n8263), .A(n7463), .ZN(n7464) );
  OAI21_X1 U9305 ( .B1(n7465), .B2(n8267), .A(n7464), .ZN(P2_U3164) );
  NAND2_X1 U9306 ( .A1(n7467), .A2(n7466), .ZN(n7496) );
  XOR2_X1 U9307 ( .A(n7496), .B(n7472), .Z(n7470) );
  OR2_X1 U9308 ( .A1(n7484), .A2(n8946), .ZN(n7469) );
  NAND2_X1 U9309 ( .A1(n9260), .A2(n9232), .ZN(n7468) );
  NAND2_X1 U9310 ( .A1(n7469), .A2(n7468), .ZN(n7591) );
  AOI21_X1 U9311 ( .B1(n7470), .B2(n9549), .A(n7591), .ZN(n7543) );
  OAI21_X1 U9312 ( .B1(n7473), .B2(n7472), .A(n7471), .ZN(n7541) );
  AOI21_X1 U9313 ( .B1(n7474), .B2(n7601), .A(n9578), .ZN(n7475) );
  NAND2_X1 U9314 ( .A1(n7475), .A2(n7504), .ZN(n7542) );
  OAI22_X1 U9315 ( .A1(n9561), .A2(n7476), .B1(n7594), .B2(n9869), .ZN(n7477)
         );
  AOI21_X1 U9316 ( .B1(n9866), .B2(n7601), .A(n7477), .ZN(n7478) );
  OAI21_X1 U9317 ( .B1(n7542), .B2(n9859), .A(n7478), .ZN(n7479) );
  AOI21_X1 U9318 ( .B1(n7541), .B2(n9535), .A(n7479), .ZN(n7480) );
  OAI21_X1 U9319 ( .B1(n7543), .B2(n9857), .A(n7480), .ZN(P1_U3285) );
  OAI21_X1 U9320 ( .B1(n7483), .B2(n7482), .A(n7481), .ZN(n7487) );
  OR2_X1 U9321 ( .A1(n7484), .A2(n8944), .ZN(n7486) );
  OR2_X1 U9322 ( .A1(n7606), .A2(n8946), .ZN(n7485) );
  NAND2_X1 U9323 ( .A1(n7486), .A2(n7485), .ZN(n9763) );
  AOI21_X1 U9324 ( .B1(n7487), .B2(n9549), .A(n9763), .ZN(n7533) );
  OAI21_X1 U9325 ( .B1(n7489), .B2(n9115), .A(n7488), .ZN(n7536) );
  NAND2_X1 U9326 ( .A1(n7536), .A2(n9535), .ZN(n7494) );
  AOI211_X1 U9327 ( .C1(n7538), .C2(n4644), .A(n9578), .B(n7639), .ZN(n7535)
         );
  NOR2_X1 U9328 ( .A1(n9767), .A2(n9873), .ZN(n7492) );
  OAI22_X1 U9329 ( .A1(n9561), .A2(n7490), .B1(n9771), .B2(n9869), .ZN(n7491)
         );
  AOI211_X1 U9330 ( .C1(n7535), .C2(n9877), .A(n7492), .B(n7491), .ZN(n7493)
         );
  OAI211_X1 U9331 ( .C1(n9857), .C2(n7533), .A(n7494), .B(n7493), .ZN(P1_U3283) );
  INV_X1 U9332 ( .A(n8999), .ZN(n7495) );
  AOI21_X1 U9333 ( .B1(n7496), .B2(n8995), .A(n7495), .ZN(n7497) );
  XNOR2_X1 U9334 ( .A(n7497), .B(n7501), .ZN(n7499) );
  NOR2_X1 U9335 ( .A1(n7498), .A2(n8944), .ZN(n7655) );
  AOI21_X1 U9336 ( .B1(n7499), .B2(n9549), .A(n7655), .ZN(n7581) );
  OAI21_X1 U9337 ( .B1(n7502), .B2(n7501), .A(n7500), .ZN(n7579) );
  AOI211_X1 U9338 ( .C1(n7660), .C2(n7504), .A(n9578), .B(n7503), .ZN(n7505)
         );
  NOR2_X1 U9339 ( .A1(n7634), .A2(n8946), .ZN(n7654) );
  NOR2_X1 U9340 ( .A1(n7505), .A2(n7654), .ZN(n7580) );
  OAI22_X1 U9341 ( .A1(n9561), .A2(n7506), .B1(n7658), .B2(n9869), .ZN(n7507)
         );
  AOI21_X1 U9342 ( .B1(n9866), .B2(n7660), .A(n7507), .ZN(n7508) );
  OAI21_X1 U9343 ( .B1(n7580), .B2(n9859), .A(n7508), .ZN(n7509) );
  AOI21_X1 U9344 ( .B1(n7579), .B2(n9535), .A(n7509), .ZN(n7510) );
  OAI21_X1 U9345 ( .B1(n7581), .B2(n9857), .A(n7510), .ZN(P1_U3284) );
  INV_X1 U9346 ( .A(n7511), .ZN(n7514) );
  OAI222_X1 U9347 ( .A1(n8787), .A2(n7514), .B1(P2_U3151), .B2(n7513), .C1(
        n7512), .C2(n8765), .ZN(P2_U3275) );
  OAI222_X1 U9348 ( .A1(n9735), .A2(n7515), .B1(n9738), .B2(n7514), .C1(n9223), 
        .C2(P1_U3086), .ZN(P1_U3335) );
  OR2_X1 U9349 ( .A1(n7982), .A2(n4862), .ZN(n8123) );
  INV_X1 U9350 ( .A(n8123), .ZN(n7516) );
  XNOR2_X1 U9351 ( .A(n7517), .B(n7516), .ZN(n10142) );
  XNOR2_X1 U9352 ( .A(n7518), .B(n8123), .ZN(n7522) );
  AOI22_X1 U9353 ( .A1(n8310), .A2(n8620), .B1(n8618), .B2(n8312), .ZN(n7519)
         );
  OAI21_X1 U9354 ( .B1(n10142), .B2(n7520), .A(n7519), .ZN(n7521) );
  AOI21_X1 U9355 ( .B1(n7522), .B2(n8623), .A(n7521), .ZN(n10143) );
  MUX2_X1 U9356 ( .A(n7773), .B(n10143), .S(n8610), .Z(n7526) );
  INV_X1 U9357 ( .A(n7523), .ZN(n7524) );
  AOI22_X1 U9358 ( .A1(n10146), .A2(n8627), .B1(n8626), .B2(n7524), .ZN(n7525)
         );
  OAI211_X1 U9359 ( .C1(n10142), .C2(n7926), .A(n7526), .B(n7525), .ZN(
        P2_U3223) );
  INV_X1 U9360 ( .A(n7527), .ZN(n7531) );
  OAI222_X1 U9361 ( .A1(n8787), .A2(n7531), .B1(P2_U3151), .B2(n7529), .C1(
        n7528), .C2(n8765), .ZN(P2_U3274) );
  OAI222_X1 U9362 ( .A1(n9735), .A2(n7532), .B1(n9738), .B2(n7531), .C1(n7530), 
        .C2(P1_U3086), .ZN(P1_U3334) );
  INV_X1 U9363 ( .A(n7533), .ZN(n7534) );
  AOI211_X1 U9364 ( .C1(n9908), .C2(n7536), .A(n7535), .B(n7534), .ZN(n7540)
         );
  INV_X1 U9365 ( .A(n9713), .ZN(n7587) );
  AOI22_X1 U9366 ( .A1(n7538), .A2(n7587), .B1(n9910), .B2(
        P1_REG0_REG_10__SCAN_IN), .ZN(n7537) );
  OAI21_X1 U9367 ( .B1(n7540), .B2(n9910), .A(n7537), .ZN(P1_U3483) );
  AOI22_X1 U9368 ( .A1(n7538), .A2(n6638), .B1(n9916), .B2(
        P1_REG1_REG_10__SCAN_IN), .ZN(n7539) );
  OAI21_X1 U9369 ( .B1(n7540), .B2(n9916), .A(n7539), .ZN(P1_U3532) );
  INV_X1 U9370 ( .A(n7541), .ZN(n7544) );
  OAI211_X1 U9371 ( .C1(n7583), .C2(n7544), .A(n7543), .B(n7542), .ZN(n7547)
         );
  NAND2_X1 U9372 ( .A1(n7547), .A2(n9918), .ZN(n7546) );
  NAND2_X1 U9373 ( .A1(n6638), .A2(n7601), .ZN(n7545) );
  OAI211_X1 U9374 ( .C1(n9918), .C2(n6805), .A(n7546), .B(n7545), .ZN(P1_U3530) );
  NAND2_X1 U9375 ( .A1(n7547), .A2(n9911), .ZN(n7549) );
  NAND2_X1 U9376 ( .A1(n7587), .A2(n7601), .ZN(n7548) );
  OAI211_X1 U9377 ( .C1(n9911), .C2(n5339), .A(n7549), .B(n7548), .ZN(P1_U3477) );
  XNOR2_X1 U9378 ( .A(n7851), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n7846) );
  OAI21_X1 U9379 ( .B1(n7556), .B2(P1_REG1_REG_12__SCAN_IN), .A(n7550), .ZN(
        n9792) );
  MUX2_X1 U9380 ( .A(n7551), .B(P1_REG1_REG_13__SCAN_IN), .S(n9799), .Z(n9793)
         );
  NOR2_X1 U9381 ( .A1(n9792), .A2(n9793), .ZN(n9791) );
  AOI21_X1 U9382 ( .B1(P1_REG1_REG_13__SCAN_IN), .B2(n9799), .A(n9791), .ZN(
        n9808) );
  XNOR2_X1 U9383 ( .A(n9811), .B(P1_REG1_REG_14__SCAN_IN), .ZN(n9807) );
  NOR2_X1 U9384 ( .A1(n9808), .A2(n9807), .ZN(n9806) );
  AOI21_X1 U9385 ( .B1(n9811), .B2(P1_REG1_REG_14__SCAN_IN), .A(n9806), .ZN(
        n7552) );
  NOR2_X1 U9386 ( .A1(n7552), .A2(n7558), .ZN(n7553) );
  XNOR2_X1 U9387 ( .A(n7558), .B(n7552), .ZN(n9817) );
  NOR2_X1 U9388 ( .A1(n9816), .A2(n9817), .ZN(n9815) );
  NOR2_X1 U9389 ( .A1(n7553), .A2(n9815), .ZN(n9827) );
  XOR2_X1 U9390 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9837), .Z(n9828) );
  AOI22_X1 U9391 ( .A1(n9827), .A2(n9828), .B1(n7554), .B2(n10443), .ZN(n7847)
         );
  XOR2_X1 U9392 ( .A(n7846), .B(n7847), .Z(n7568) );
  XNOR2_X1 U9393 ( .A(n7851), .B(n9539), .ZN(n7563) );
  OAI21_X1 U9394 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(n7556), .A(n7555), .ZN(
        n9796) );
  XNOR2_X1 U9395 ( .A(n9799), .B(P1_REG2_REG_13__SCAN_IN), .ZN(n9795) );
  NOR2_X1 U9396 ( .A1(n9796), .A2(n9795), .ZN(n9794) );
  AOI21_X1 U9397 ( .B1(P1_REG2_REG_13__SCAN_IN), .B2(n9799), .A(n9794), .ZN(
        n9805) );
  NAND2_X1 U9398 ( .A1(P1_REG2_REG_14__SCAN_IN), .A2(n9811), .ZN(n7557) );
  OAI21_X1 U9399 ( .B1(P1_REG2_REG_14__SCAN_IN), .B2(n9811), .A(n7557), .ZN(
        n9804) );
  NOR2_X1 U9400 ( .A1(n9805), .A2(n9804), .ZN(n9803) );
  AOI21_X1 U9401 ( .B1(n9811), .B2(P1_REG2_REG_14__SCAN_IN), .A(n9803), .ZN(
        n7559) );
  NOR2_X1 U9402 ( .A1(n7559), .A2(n7558), .ZN(n7560) );
  XOR2_X1 U9403 ( .A(n9822), .B(n7559), .Z(n9819) );
  NOR2_X1 U9404 ( .A1(n7871), .A2(n9819), .ZN(n9818) );
  NOR2_X1 U9405 ( .A1(n7560), .A2(n9818), .ZN(n9834) );
  XNOR2_X1 U9406 ( .A(n9837), .B(P1_REG2_REG_16__SCAN_IN), .ZN(n9833) );
  OR2_X1 U9407 ( .A1(n9834), .A2(n9833), .ZN(n9830) );
  NAND2_X1 U9408 ( .A1(n9837), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n7561) );
  AND2_X1 U9409 ( .A1(n9830), .A2(n7561), .ZN(n7562) );
  NAND2_X1 U9410 ( .A1(n7562), .A2(n7563), .ZN(n7853) );
  OAI21_X1 U9411 ( .B1(n7563), .B2(n7562), .A(n7853), .ZN(n7564) );
  NAND2_X1 U9412 ( .A1(n7564), .A2(n10559), .ZN(n7567) );
  NAND2_X1 U9413 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n8872) );
  OAI21_X1 U9414 ( .B1(n9853), .B2(n10456), .A(n8872), .ZN(n7565) );
  AOI21_X1 U9415 ( .B1(n7851), .B2(n10568), .A(n7565), .ZN(n7566) );
  OAI211_X1 U9416 ( .C1(n9845), .C2(n7568), .A(n7567), .B(n7566), .ZN(P1_U3260) );
  XNOR2_X1 U9417 ( .A(n8005), .B(n8189), .ZN(n7570) );
  INV_X1 U9418 ( .A(n7570), .ZN(n7569) );
  NAND2_X1 U9419 ( .A1(n7569), .A2(n8308), .ZN(n7622) );
  NAND2_X1 U9420 ( .A1(n7570), .A2(n7734), .ZN(n7620) );
  NAND2_X1 U9421 ( .A1(n7622), .A2(n7620), .ZN(n7573) );
  XOR2_X1 U9422 ( .A(n7573), .B(n7621), .Z(n7578) );
  NAND2_X1 U9423 ( .A1(P2_U3151), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n7798) );
  OAI21_X1 U9424 ( .B1(n8286), .B2(n7721), .A(n7798), .ZN(n7574) );
  AOI21_X1 U9425 ( .B1(n8284), .B2(n8309), .A(n7574), .ZN(n7575) );
  OAI21_X1 U9426 ( .B1(n7742), .B2(n8252), .A(n7575), .ZN(n7576) );
  AOI21_X1 U9427 ( .B1(n8005), .B2(n8263), .A(n7576), .ZN(n7577) );
  OAI21_X1 U9428 ( .B1(n7578), .B2(n8267), .A(n7577), .ZN(P2_U3174) );
  INV_X1 U9429 ( .A(n7579), .ZN(n7582) );
  OAI211_X1 U9430 ( .C1(n7583), .C2(n7582), .A(n7581), .B(n7580), .ZN(n7586)
         );
  NAND2_X1 U9431 ( .A1(n7586), .A2(n9918), .ZN(n7585) );
  NAND2_X1 U9432 ( .A1(n6638), .A2(n7660), .ZN(n7584) );
  OAI211_X1 U9433 ( .C1(n9918), .C2(n5363), .A(n7585), .B(n7584), .ZN(P1_U3531) );
  INV_X1 U9434 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n7590) );
  NAND2_X1 U9435 ( .A1(n7586), .A2(n9911), .ZN(n7589) );
  NAND2_X1 U9436 ( .A1(n7587), .A2(n7660), .ZN(n7588) );
  OAI211_X1 U9437 ( .C1(n9911), .C2(n7590), .A(n7589), .B(n7588), .ZN(P1_U3480) );
  NAND2_X1 U9438 ( .A1(n9764), .A2(n7591), .ZN(n7593) );
  INV_X1 U9439 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n7592) );
  OR2_X1 U9440 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7592), .ZN(n9319) );
  OAI211_X1 U9441 ( .C1(n9772), .C2(n7594), .A(n7593), .B(n9319), .ZN(n7600)
         );
  NAND2_X1 U9442 ( .A1(n7595), .A2(n7596), .ZN(n7597) );
  AOI21_X1 U9443 ( .B1(n7598), .B2(n7597), .A(n9758), .ZN(n7599) );
  AOI211_X1 U9444 ( .C1(n7601), .C2(n8958), .A(n7600), .B(n7599), .ZN(n7602)
         );
  INV_X1 U9445 ( .A(n7602), .ZN(P1_U3221) );
  XNOR2_X1 U9446 ( .A(n7603), .B(n7612), .ZN(n7604) );
  NAND2_X1 U9447 ( .A1(n7604), .A2(n9549), .ZN(n7610) );
  OR2_X1 U9448 ( .A1(n7605), .A2(n8946), .ZN(n7608) );
  OR2_X1 U9449 ( .A1(n7606), .A2(n8944), .ZN(n7607) );
  NAND2_X1 U9450 ( .A1(n7608), .A2(n7607), .ZN(n8837) );
  INV_X1 U9451 ( .A(n8837), .ZN(n7609) );
  NAND2_X1 U9452 ( .A1(n7610), .A2(n7609), .ZN(n7691) );
  INV_X1 U9453 ( .A(n7691), .ZN(n7619) );
  OAI21_X1 U9454 ( .B1(n7613), .B2(n7612), .A(n7611), .ZN(n7693) );
  NAND2_X1 U9455 ( .A1(n7693), .A2(n9535), .ZN(n7618) );
  INV_X1 U9456 ( .A(n5147), .ZN(n7707) );
  AOI211_X1 U9457 ( .C1(n8842), .C2(n7640), .A(n9578), .B(n7707), .ZN(n7692)
         );
  INV_X1 U9458 ( .A(n8842), .ZN(n7697) );
  NOR2_X1 U9459 ( .A1(n7697), .A2(n9873), .ZN(n7616) );
  OAI22_X1 U9460 ( .A1(n9561), .A2(n7614), .B1(n8840), .B2(n9869), .ZN(n7615)
         );
  AOI211_X1 U9461 ( .C1(n7692), .C2(n9877), .A(n7616), .B(n7615), .ZN(n7617)
         );
  OAI211_X1 U9462 ( .C1(n9857), .C2(n7619), .A(n7618), .B(n7617), .ZN(P1_U3281) );
  NAND2_X1 U9463 ( .A1(n7621), .A2(n7620), .ZN(n7623) );
  XNOR2_X1 U9464 ( .A(n7887), .B(n8196), .ZN(n7712) );
  XNOR2_X1 U9465 ( .A(n7712), .B(n8307), .ZN(n7715) );
  XOR2_X1 U9466 ( .A(n7716), .B(n7715), .Z(n7628) );
  NAND2_X1 U9467 ( .A1(P2_U3151), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n8330) );
  OAI21_X1 U9468 ( .B1(n8286), .B2(n7841), .A(n8330), .ZN(n7624) );
  AOI21_X1 U9469 ( .B1(n8284), .B2(n8308), .A(n7624), .ZN(n7625) );
  OAI21_X1 U9470 ( .B1(n7888), .B2(n8252), .A(n7625), .ZN(n7626) );
  AOI21_X1 U9471 ( .B1(n7887), .B2(n8263), .A(n7626), .ZN(n7627) );
  OAI21_X1 U9472 ( .B1(n7628), .B2(n8267), .A(n7627), .ZN(P2_U3155) );
  OAI21_X1 U9473 ( .B1(n7630), .B2(n7633), .A(n7629), .ZN(n7727) );
  INV_X1 U9474 ( .A(n7727), .ZN(n7649) );
  NOR2_X1 U9475 ( .A1(n9857), .A2(n7631), .ZN(n9878) );
  INV_X1 U9476 ( .A(n9878), .ZN(n7648) );
  XOR2_X1 U9477 ( .A(n7633), .B(n7632), .Z(n7637) );
  OR2_X1 U9478 ( .A1(n7700), .A2(n8946), .ZN(n7636) );
  OR2_X1 U9479 ( .A1(n7634), .A2(n8944), .ZN(n7635) );
  NAND2_X1 U9480 ( .A1(n7636), .A2(n7635), .ZN(n8922) );
  AOI21_X1 U9481 ( .B1(n7637), .B2(n9549), .A(n8922), .ZN(n7638) );
  OAI21_X1 U9482 ( .B1(n7649), .B2(n9564), .A(n7638), .ZN(n7725) );
  NAND2_X1 U9483 ( .A1(n7725), .A2(n9561), .ZN(n7647) );
  INV_X1 U9484 ( .A(n7639), .ZN(n7642) );
  INV_X1 U9485 ( .A(n7640), .ZN(n7641) );
  AOI211_X1 U9486 ( .C1(n4622), .C2(n7642), .A(n9578), .B(n7641), .ZN(n7726)
         );
  NOR2_X1 U9487 ( .A1(n7733), .A2(n9873), .ZN(n7645) );
  OAI22_X1 U9488 ( .A1(n9561), .A2(n7643), .B1(n8924), .B2(n9869), .ZN(n7644)
         );
  AOI211_X1 U9489 ( .C1(n7726), .C2(n9877), .A(n7645), .B(n7644), .ZN(n7646)
         );
  OAI211_X1 U9490 ( .C1(n7649), .C2(n7648), .A(n7647), .B(n7646), .ZN(P1_U3282) );
  OAI21_X1 U9491 ( .B1(n7652), .B2(n7651), .A(n7650), .ZN(n7653) );
  NAND2_X1 U9492 ( .A1(n7653), .A2(n8942), .ZN(n7662) );
  OAI21_X1 U9493 ( .B1(n7655), .B2(n7654), .A(n9764), .ZN(n7657) );
  OAI211_X1 U9494 ( .C1(n9772), .C2(n7658), .A(n7657), .B(n7656), .ZN(n7659)
         );
  AOI21_X1 U9495 ( .B1(n7660), .B2(n8958), .A(n7659), .ZN(n7661) );
  NAND2_X1 U9496 ( .A1(n7662), .A2(n7661), .ZN(P1_U3231) );
  OAI21_X1 U9497 ( .B1(n7664), .B2(n7666), .A(n7663), .ZN(n8687) );
  INV_X1 U9498 ( .A(n8687), .ZN(n7671) );
  XNOR2_X1 U9499 ( .A(n7665), .B(n7666), .ZN(n7667) );
  AOI222_X1 U9500 ( .A1(n8623), .A2(n7667), .B1(n8309), .B2(n8620), .C1(n8311), 
        .C2(n8618), .ZN(n8689) );
  MUX2_X1 U9501 ( .A(n7818), .B(n8689), .S(n8610), .Z(n7670) );
  AOI22_X1 U9502 ( .A1(n8686), .A2(n8627), .B1(n8626), .B2(n7668), .ZN(n7669)
         );
  OAI211_X1 U9503 ( .C1(n7671), .C2(n8630), .A(n7670), .B(n7669), .ZN(P2_U3222) );
  XNOR2_X1 U9504 ( .A(n7672), .B(n8125), .ZN(n7685) );
  NAND2_X1 U9505 ( .A1(n10148), .A2(n10123), .ZN(n8760) );
  XNOR2_X1 U9506 ( .A(n7673), .B(n8125), .ZN(n7674) );
  OAI222_X1 U9507 ( .A1(n8598), .A2(n7734), .B1(n8596), .B2(n7675), .C1(n8593), 
        .C2(n7674), .ZN(n7680) );
  NAND2_X1 U9508 ( .A1(n7680), .A2(n10148), .ZN(n7677) );
  AOI22_X1 U9509 ( .A1(n8000), .A2(n8756), .B1(P2_REG0_REG_12__SCAN_IN), .B2(
        n10149), .ZN(n7676) );
  OAI211_X1 U9510 ( .C1(n7685), .C2(n8760), .A(n7677), .B(n7676), .ZN(P2_U3426) );
  NAND2_X1 U9511 ( .A1(n10159), .A2(n10123), .ZN(n8681) );
  NAND2_X1 U9512 ( .A1(n7680), .A2(n10159), .ZN(n7679) );
  AOI22_X1 U9513 ( .A1(n8000), .A2(n8678), .B1(P2_REG1_REG_12__SCAN_IN), .B2(
        n10157), .ZN(n7678) );
  OAI211_X1 U9514 ( .C1(n7685), .C2(n8681), .A(n7679), .B(n7678), .ZN(P2_U3471) );
  NAND2_X1 U9515 ( .A1(n7680), .A2(n8610), .ZN(n7684) );
  OAI22_X1 U9516 ( .A1(n10103), .A2(n7775), .B1(n7681), .B2(n10097), .ZN(n7682) );
  AOI21_X1 U9517 ( .B1(n8000), .B2(n8627), .A(n7682), .ZN(n7683) );
  OAI211_X1 U9518 ( .C1(n7685), .C2(n8630), .A(n7684), .B(n7683), .ZN(P2_U3221) );
  INV_X1 U9519 ( .A(n7686), .ZN(n7689) );
  OAI222_X1 U9520 ( .A1(n9735), .A2(n7687), .B1(n9738), .B2(n7689), .C1(
        P1_U3086), .C2(n9099), .ZN(P1_U3333) );
  OAI222_X1 U9521 ( .A1(n8765), .A2(n7690), .B1(n8787), .B2(n7689), .C1(n7688), 
        .C2(P2_U3151), .ZN(P2_U3273) );
  AOI211_X1 U9522 ( .C1(n7693), .C2(n9908), .A(n7692), .B(n7691), .ZN(n7695)
         );
  MUX2_X1 U9523 ( .A(n5421), .B(n7695), .S(n9918), .Z(n7694) );
  OAI21_X1 U9524 ( .B1(n7697), .B2(n9652), .A(n7694), .ZN(P1_U3534) );
  MUX2_X1 U9525 ( .A(n5415), .B(n7695), .S(n9911), .Z(n7696) );
  OAI21_X1 U9526 ( .B1(n7697), .B2(n9713), .A(n7696), .ZN(P1_U3489) );
  NAND2_X1 U9527 ( .A1(n7698), .A2(n9103), .ZN(n7699) );
  NAND2_X1 U9528 ( .A1(n9568), .A2(n7699), .ZN(n7703) );
  OR2_X1 U9529 ( .A1(n7700), .A2(n8944), .ZN(n7702) );
  NAND2_X1 U9530 ( .A1(n9253), .A2(n8932), .ZN(n7701) );
  NAND2_X1 U9531 ( .A1(n7702), .A2(n7701), .ZN(n8897) );
  AOI21_X1 U9532 ( .B1(n7703), .B2(n9549), .A(n8897), .ZN(n9904) );
  OAI21_X1 U9533 ( .B1(n7705), .B2(n9103), .A(n7704), .ZN(n9909) );
  NAND2_X1 U9534 ( .A1(n9909), .A2(n9535), .ZN(n7711) );
  INV_X1 U9535 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n7706) );
  OAI22_X1 U9536 ( .A1(n9561), .A2(n7706), .B1(n8899), .B2(n9869), .ZN(n7709)
         );
  INV_X1 U9537 ( .A(n8901), .ZN(n9906) );
  OAI211_X1 U9538 ( .C1(n7707), .C2(n9906), .A(n7872), .B(n9579), .ZN(n9903)
         );
  NOR2_X1 U9539 ( .A1(n9903), .A2(n9859), .ZN(n7708) );
  AOI211_X1 U9540 ( .C1(n9866), .C2(n8901), .A(n7709), .B(n7708), .ZN(n7710)
         );
  OAI211_X1 U9541 ( .C1(n9857), .C2(n9904), .A(n7711), .B(n7710), .ZN(P1_U3280) );
  INV_X1 U9542 ( .A(n8682), .ZN(n7903) );
  INV_X1 U9543 ( .A(n7712), .ZN(n7713) );
  NAND2_X1 U9544 ( .A1(n7713), .A2(n7721), .ZN(n7714) );
  XNOR2_X1 U9545 ( .A(n8682), .B(n8196), .ZN(n7837) );
  XNOR2_X1 U9546 ( .A(n7837), .B(n8619), .ZN(n7717) );
  AOI21_X1 U9547 ( .B1(n7718), .B2(n7717), .A(n8267), .ZN(n7719) );
  NAND2_X1 U9548 ( .A1(n7719), .A2(n7838), .ZN(n7724) );
  NAND2_X1 U9549 ( .A1(n8300), .A2(n8608), .ZN(n7720) );
  NAND2_X1 U9550 ( .A1(P2_U3151), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8352) );
  OAI211_X1 U9551 ( .C1(n7721), .C2(n8297), .A(n7720), .B(n8352), .ZN(n7722)
         );
  AOI21_X1 U9552 ( .B1(n7901), .B2(n8295), .A(n7722), .ZN(n7723) );
  OAI211_X1 U9553 ( .C1(n7903), .C2(n8303), .A(n7724), .B(n7723), .ZN(P2_U3181) );
  AOI211_X1 U9554 ( .C1(n7728), .C2(n7727), .A(n7726), .B(n7725), .ZN(n7730)
         );
  MUX2_X1 U9555 ( .A(n6847), .B(n7730), .S(n9918), .Z(n7729) );
  OAI21_X1 U9556 ( .B1(n7733), .B2(n9652), .A(n7729), .ZN(P1_U3533) );
  INV_X1 U9557 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n7731) );
  MUX2_X1 U9558 ( .A(n7731), .B(n7730), .S(n9911), .Z(n7732) );
  OAI21_X1 U9559 ( .B1(n7733), .B2(n9713), .A(n7732), .ZN(P1_U3486) );
  XNOR2_X1 U9560 ( .A(n8005), .B(n7734), .ZN(n8127) );
  XOR2_X1 U9561 ( .A(n8127), .B(n7735), .Z(n7759) );
  INV_X1 U9562 ( .A(n8005), .ZN(n7740) );
  XNOR2_X1 U9563 ( .A(n7736), .B(n8127), .ZN(n7737) );
  NAND2_X1 U9564 ( .A1(n7737), .A2(n8623), .ZN(n7739) );
  AOI22_X1 U9565 ( .A1(n8618), .A2(n8309), .B1(n8307), .B2(n8620), .ZN(n7738)
         );
  OAI21_X1 U9566 ( .B1(n7740), .B2(n8523), .A(n7756), .ZN(n7741) );
  NAND2_X1 U9567 ( .A1(n7741), .A2(n8610), .ZN(n7745) );
  INV_X1 U9568 ( .A(n7742), .ZN(n7743) );
  AOI22_X1 U9569 ( .A1(n10105), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n8626), .B2(
        n7743), .ZN(n7744) );
  OAI211_X1 U9570 ( .C1(n7759), .C2(n8630), .A(n7745), .B(n7744), .ZN(P2_U3220) );
  NAND2_X1 U9571 ( .A1(n7750), .A2(n8774), .ZN(n7747) );
  NAND2_X1 U9572 ( .A1(n7746), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8154) );
  OAI211_X1 U9573 ( .C1(n7748), .C2(n8765), .A(n7747), .B(n8154), .ZN(P2_U3272) );
  NAND2_X1 U9574 ( .A1(n7750), .A2(n7749), .ZN(n7751) );
  OAI211_X1 U9575 ( .C1(n7752), .C2(n9735), .A(n7751), .B(n9235), .ZN(P1_U3332) );
  INV_X1 U9576 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n7753) );
  MUX2_X1 U9577 ( .A(n7753), .B(n7756), .S(n10148), .Z(n7755) );
  NAND2_X1 U9578 ( .A1(n8005), .A2(n8756), .ZN(n7754) );
  OAI211_X1 U9579 ( .C1(n7759), .C2(n8760), .A(n7755), .B(n7754), .ZN(P2_U3429) );
  MUX2_X1 U9580 ( .A(n10413), .B(n7756), .S(n10159), .Z(n7758) );
  NAND2_X1 U9581 ( .A1(n8005), .A2(n8678), .ZN(n7757) );
  OAI211_X1 U9582 ( .C1(n8681), .C2(n7759), .A(n7758), .B(n7757), .ZN(P2_U3472) );
  NAND2_X1 U9583 ( .A1(n7780), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n7760) );
  NAND2_X1 U9584 ( .A1(n7761), .A2(n7760), .ZN(n7762) );
  NAND2_X1 U9585 ( .A1(n7762), .A2(n9951), .ZN(n9962) );
  AND2_X2 U9586 ( .A1(n7763), .A2(n9962), .ZN(n9945) );
  NAND2_X1 U9587 ( .A1(n9964), .A2(n9962), .ZN(n7765) );
  XNOR2_X1 U9588 ( .A(n9976), .B(n7764), .ZN(n9961) );
  NOR2_X1 U9589 ( .A1(n7787), .A2(n5139), .ZN(n7767) );
  NAND2_X1 U9590 ( .A1(P2_REG2_REG_8__SCAN_IN), .A2(n7778), .ZN(n7768) );
  OAI21_X1 U9591 ( .B1(n7778), .B2(P2_REG2_REG_8__SCAN_IN), .A(n7768), .ZN(
        n10010) );
  NOR2_X1 U9592 ( .A1(n10017), .A2(n7769), .ZN(n7770) );
  NAND2_X1 U9593 ( .A1(P2_REG2_REG_10__SCAN_IN), .A2(n7777), .ZN(n7771) );
  OAI21_X1 U9594 ( .B1(n7777), .B2(P2_REG2_REG_10__SCAN_IN), .A(n7771), .ZN(
        n10041) );
  INV_X1 U9595 ( .A(n10040), .ZN(n7772) );
  OAI21_X1 U9596 ( .B1(n10031), .B2(n7773), .A(n7772), .ZN(n7774) );
  XNOR2_X1 U9597 ( .A(n7774), .B(n10050), .ZN(n10061) );
  NOR2_X1 U9598 ( .A1(n10061), .A2(n7818), .ZN(n10060) );
  XNOR2_X1 U9599 ( .A(n10068), .B(n7775), .ZN(n10086) );
  AOI21_X2 U9600 ( .B1(P2_REG2_REG_12__SCAN_IN), .B2(n7822), .A(n10085), .ZN(
        n8320) );
  XNOR2_X1 U9601 ( .A(n8321), .B(n8320), .ZN(n7776) );
  AOI21_X1 U9602 ( .B1(n7825), .B2(n7776), .A(n8322), .ZN(n7836) );
  AOI22_X1 U9603 ( .A1(P2_REG1_REG_12__SCAN_IN), .A2(n7822), .B1(n10068), .B2(
        n7796), .ZN(n10072) );
  NAND2_X1 U9604 ( .A1(P2_REG1_REG_10__SCAN_IN), .A2(n7777), .ZN(n7793) );
  AOI22_X1 U9605 ( .A1(n10031), .A2(n6356), .B1(P2_REG1_REG_10__SCAN_IN), .B2(
        n7777), .ZN(n10036) );
  NAND2_X1 U9606 ( .A1(P2_REG1_REG_8__SCAN_IN), .A2(n7778), .ZN(n7790) );
  AOI22_X1 U9607 ( .A1(P2_REG1_REG_8__SCAN_IN), .A2(n7778), .B1(n10004), .B2(
        n6326), .ZN(n10003) );
  NAND2_X1 U9608 ( .A1(n9976), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n7786) );
  INV_X1 U9609 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n7779) );
  MUX2_X1 U9610 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n7779), .S(n9976), .Z(n9971)
         );
  NAND2_X1 U9611 ( .A1(n7780), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n7781) );
  INV_X1 U9612 ( .A(n9951), .ZN(n7807) );
  XNOR2_X1 U9613 ( .A(n7783), .B(n7807), .ZN(n9944) );
  NAND2_X1 U9614 ( .A1(n9944), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n7785) );
  NAND2_X1 U9615 ( .A1(n7783), .A2(n9951), .ZN(n7784) );
  NAND2_X1 U9616 ( .A1(n7785), .A2(n7784), .ZN(n9972) );
  NAND2_X1 U9617 ( .A1(n9971), .A2(n9972), .ZN(n9970) );
  NAND2_X1 U9618 ( .A1(n7786), .A2(n9970), .ZN(n7788) );
  NAND2_X1 U9619 ( .A1(n9989), .A2(n7788), .ZN(n7789) );
  XNOR2_X1 U9620 ( .A(n7788), .B(n7787), .ZN(n9986) );
  NAND2_X1 U9621 ( .A1(P2_REG1_REG_7__SCAN_IN), .A2(n9986), .ZN(n9985) );
  NAND2_X1 U9622 ( .A1(n7789), .A2(n9985), .ZN(n10002) );
  NAND2_X1 U9623 ( .A1(n4802), .A2(n7791), .ZN(n7792) );
  XNOR2_X1 U9624 ( .A(n7791), .B(n10017), .ZN(n10021) );
  NAND2_X1 U9625 ( .A1(P2_REG1_REG_9__SCAN_IN), .A2(n10021), .ZN(n10020) );
  NAND2_X1 U9626 ( .A1(n7792), .A2(n10020), .ZN(n10035) );
  NAND2_X1 U9627 ( .A1(n7794), .A2(n10050), .ZN(n7795) );
  XNOR2_X1 U9628 ( .A(n7794), .B(n7819), .ZN(n10056) );
  NAND2_X1 U9629 ( .A1(P2_REG1_REG_11__SCAN_IN), .A2(n10056), .ZN(n10055) );
  NAND2_X1 U9630 ( .A1(n7795), .A2(n10055), .ZN(n10071) );
  NAND2_X1 U9631 ( .A1(n10072), .A2(n10071), .ZN(n10070) );
  OAI21_X1 U9632 ( .B1(n10068), .B2(n7796), .A(n10070), .ZN(n8324) );
  OAI21_X1 U9633 ( .B1(P2_REG1_REG_13__SCAN_IN), .B2(n7797), .A(n8326), .ZN(
        n7834) );
  INV_X1 U9634 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n7800) );
  NAND2_X1 U9635 ( .A1(n10069), .A2(n8321), .ZN(n7799) );
  OAI211_X1 U9636 ( .C1(n10049), .C2(n7800), .A(n7799), .B(n7798), .ZN(n7833)
         );
  MUX2_X1 U9637 ( .A(P2_REG2_REG_6__SCAN_IN), .B(P2_REG1_REG_6__SCAN_IN), .S(
        n8779), .Z(n7808) );
  INV_X1 U9638 ( .A(n7808), .ZN(n7809) );
  MUX2_X1 U9639 ( .A(P2_REG2_REG_5__SCAN_IN), .B(P2_REG1_REG_5__SCAN_IN), .S(
        n8779), .Z(n7805) );
  INV_X1 U9640 ( .A(n7805), .ZN(n7806) );
  INV_X1 U9641 ( .A(n7801), .ZN(n7803) );
  OAI21_X1 U9642 ( .B1(n7804), .B2(n7803), .A(n7802), .ZN(n9954) );
  XOR2_X1 U9643 ( .A(n9951), .B(n7805), .Z(n9953) );
  NAND2_X1 U9644 ( .A1(n9954), .A2(n9953), .ZN(n9952) );
  OAI21_X1 U9645 ( .B1(n7807), .B2(n7806), .A(n9952), .ZN(n9979) );
  XNOR2_X1 U9646 ( .A(n7808), .B(n9976), .ZN(n9980) );
  NOR2_X1 U9647 ( .A1(n9979), .A2(n9980), .ZN(n9978) );
  AOI21_X1 U9648 ( .B1(n7810), .B2(n7809), .A(n9978), .ZN(n9997) );
  MUX2_X1 U9649 ( .A(P2_REG2_REG_7__SCAN_IN), .B(P2_REG1_REG_7__SCAN_IN), .S(
        n8779), .Z(n7811) );
  XNOR2_X1 U9650 ( .A(n7811), .B(n9989), .ZN(n9996) );
  OAI22_X1 U9651 ( .A1(n9997), .A2(n9996), .B1(n7811), .B2(n9989), .ZN(n10007)
         );
  MUX2_X1 U9652 ( .A(P2_REG2_REG_8__SCAN_IN), .B(P2_REG1_REG_8__SCAN_IN), .S(
        n8779), .Z(n7812) );
  XNOR2_X1 U9653 ( .A(n7812), .B(n10004), .ZN(n10006) );
  INV_X1 U9654 ( .A(n7812), .ZN(n7813) );
  AOI22_X1 U9655 ( .A1(n10007), .A2(n10006), .B1(n10004), .B2(n7813), .ZN(
        n10019) );
  MUX2_X1 U9656 ( .A(P2_REG2_REG_9__SCAN_IN), .B(P2_REG1_REG_9__SCAN_IN), .S(
        n8779), .Z(n7814) );
  XNOR2_X1 U9657 ( .A(n7814), .B(n4802), .ZN(n10018) );
  OAI22_X1 U9658 ( .A1(n10019), .A2(n10018), .B1(n7814), .B2(n4802), .ZN(
        n10033) );
  MUX2_X1 U9659 ( .A(P2_REG2_REG_10__SCAN_IN), .B(P2_REG1_REG_10__SCAN_IN), 
        .S(n8779), .Z(n7815) );
  XNOR2_X1 U9660 ( .A(n7815), .B(n10031), .ZN(n10032) );
  INV_X1 U9661 ( .A(n7815), .ZN(n7816) );
  AOI22_X1 U9662 ( .A1(n10033), .A2(n10032), .B1(n10031), .B2(n7816), .ZN(
        n10054) );
  MUX2_X1 U9663 ( .A(n7818), .B(n7817), .S(n8779), .Z(n7820) );
  XNOR2_X1 U9664 ( .A(n7820), .B(n7819), .ZN(n10053) );
  INV_X1 U9665 ( .A(n7820), .ZN(n7821) );
  OAI22_X1 U9666 ( .A1(n10054), .A2(n10053), .B1(n7821), .B2(n10050), .ZN(
        n10080) );
  MUX2_X1 U9667 ( .A(P2_REG2_REG_12__SCAN_IN), .B(P2_REG1_REG_12__SCAN_IN), 
        .S(n8779), .Z(n7823) );
  NAND2_X1 U9668 ( .A1(n7823), .A2(n7822), .ZN(n10074) );
  NAND2_X1 U9669 ( .A1(n10080), .A2(n10074), .ZN(n10075) );
  INV_X1 U9670 ( .A(n7823), .ZN(n7824) );
  NAND2_X1 U9671 ( .A1(n7824), .A2(n10068), .ZN(n10073) );
  MUX2_X1 U9672 ( .A(n7825), .B(n10413), .S(n8779), .Z(n7826) );
  NAND2_X1 U9673 ( .A1(n7826), .A2(n8321), .ZN(n8332) );
  INV_X1 U9674 ( .A(n7826), .ZN(n7827) );
  NAND2_X1 U9675 ( .A1(n7827), .A2(n8325), .ZN(n7828) );
  NAND2_X1 U9676 ( .A1(n8332), .A2(n7828), .ZN(n7829) );
  AOI21_X1 U9677 ( .B1(n10075), .B2(n10073), .A(n7829), .ZN(n8339) );
  INV_X1 U9678 ( .A(n8339), .ZN(n7831) );
  NAND3_X1 U9679 ( .A1(n10075), .A2(n10073), .A3(n7829), .ZN(n7830) );
  AOI21_X1 U9680 ( .B1(n7831), .B2(n7830), .A(n10079), .ZN(n7832) );
  AOI211_X1 U9681 ( .C1(n7834), .C2(n10084), .A(n7833), .B(n7832), .ZN(n7835)
         );
  OAI21_X1 U9682 ( .B1(n7836), .B2(n10089), .A(n7835), .ZN(P2_U3195) );
  XNOR2_X1 U9683 ( .A(n8757), .B(n8196), .ZN(n7910) );
  XNOR2_X1 U9684 ( .A(n7910), .B(n7916), .ZN(n7839) );
  XNOR2_X1 U9685 ( .A(n7911), .B(n7839), .ZN(n7845) );
  NAND2_X1 U9686 ( .A1(n8300), .A2(n8621), .ZN(n7840) );
  NAND2_X1 U9687 ( .A1(P2_U3151), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8382) );
  OAI211_X1 U9688 ( .C1(n7841), .C2(n8297), .A(n7840), .B(n8382), .ZN(n7842)
         );
  AOI21_X1 U9689 ( .B1(n8625), .B2(n8295), .A(n7842), .ZN(n7844) );
  NAND2_X1 U9690 ( .A1(n8757), .A2(n8263), .ZN(n7843) );
  OAI211_X1 U9691 ( .C1(n7845), .C2(n8267), .A(n7844), .B(n7843), .ZN(P2_U3166) );
  INV_X1 U9692 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n7865) );
  OAI22_X1 U9693 ( .A1(n7847), .A2(n7846), .B1(n7851), .B2(
        P1_REG1_REG_17__SCAN_IN), .ZN(n9846) );
  NAND2_X1 U9694 ( .A1(n9850), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n7848) );
  OAI21_X1 U9695 ( .B1(n9850), .B2(P1_REG1_REG_18__SCAN_IN), .A(n7848), .ZN(
        n9847) );
  NOR2_X1 U9696 ( .A1(n9846), .A2(n9847), .ZN(n9844) );
  INV_X1 U9697 ( .A(n7848), .ZN(n7849) );
  NOR2_X1 U9698 ( .A1(n9844), .A2(n7849), .ZN(n7850) );
  XNOR2_X1 U9699 ( .A(n7850), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n7859) );
  OR2_X1 U9700 ( .A1(n7851), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n7852) );
  AND2_X1 U9701 ( .A1(n7853), .A2(n7852), .ZN(n9842) );
  NAND2_X1 U9702 ( .A1(n9850), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n7855) );
  OR2_X1 U9703 ( .A1(n9850), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n7854) );
  AND2_X1 U9704 ( .A1(n7855), .A2(n7854), .ZN(n9841) );
  NAND2_X1 U9705 ( .A1(n9842), .A2(n9841), .ZN(n9840) );
  NAND2_X1 U9706 ( .A1(n9840), .A2(n7855), .ZN(n7856) );
  XNOR2_X1 U9707 ( .A(n7856), .B(P1_REG2_REG_19__SCAN_IN), .ZN(n7861) );
  INV_X1 U9708 ( .A(n7861), .ZN(n7857) );
  AOI22_X1 U9709 ( .A1(n10563), .A2(n7859), .B1(n7857), .B2(n10559), .ZN(n7863) );
  OAI21_X1 U9710 ( .B1(n7859), .B2(n9845), .A(n7858), .ZN(n7860) );
  AOI21_X1 U9711 ( .B1(n7861), .B2(n10559), .A(n7860), .ZN(n7862) );
  MUX2_X1 U9712 ( .A(n7863), .B(n7862), .S(n4621), .Z(n7864) );
  NAND2_X1 U9713 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n8822) );
  OAI211_X1 U9714 ( .C1(n7865), .C2(n9853), .A(n7864), .B(n8822), .ZN(P1_U3262) );
  NAND2_X1 U9715 ( .A1(n9569), .A2(n9020), .ZN(n7866) );
  XNOR2_X1 U9716 ( .A(n7866), .B(n9121), .ZN(n7869) );
  OR2_X1 U9717 ( .A1(n8869), .A2(n8946), .ZN(n7868) );
  NAND2_X1 U9718 ( .A1(n9253), .A2(n9232), .ZN(n7867) );
  NAND2_X1 U9719 ( .A1(n7868), .A2(n7867), .ZN(n8954) );
  AOI21_X1 U9720 ( .B1(n7869), .B2(n9549), .A(n8954), .ZN(n9648) );
  XNOR2_X1 U9721 ( .A(n7870), .B(n9121), .ZN(n9650) );
  NAND2_X1 U9722 ( .A1(n9650), .A2(n9535), .ZN(n7876) );
  OAI22_X1 U9723 ( .A1(n9561), .A2(n7871), .B1(n8956), .B2(n9869), .ZN(n7874)
         );
  OAI211_X1 U9724 ( .C1(n9577), .C2(n9714), .A(n4534), .B(n7872), .ZN(n9647)
         );
  NOR2_X1 U9725 ( .A1(n9647), .A2(n9859), .ZN(n7873) );
  AOI211_X1 U9726 ( .C1(n9866), .C2(n9025), .A(n7874), .B(n7873), .ZN(n7875)
         );
  OAI211_X1 U9727 ( .C1(n9857), .C2(n9648), .A(n7876), .B(n7875), .ZN(P1_U3278) );
  INV_X1 U9728 ( .A(n7877), .ZN(n8012) );
  XNOR2_X1 U9729 ( .A(n7878), .B(n5022), .ZN(n7894) );
  INV_X1 U9730 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n7881) );
  XNOR2_X1 U9731 ( .A(n7879), .B(n8011), .ZN(n7880) );
  AOI222_X1 U9732 ( .A1(n8623), .A2(n7880), .B1(n8619), .B2(n8620), .C1(n8308), 
        .C2(n8618), .ZN(n7886) );
  MUX2_X1 U9733 ( .A(n7881), .B(n7886), .S(n10148), .Z(n7883) );
  NAND2_X1 U9734 ( .A1(n7887), .A2(n8756), .ZN(n7882) );
  OAI211_X1 U9735 ( .C1(n7894), .C2(n8760), .A(n7883), .B(n7882), .ZN(P2_U3432) );
  MUX2_X1 U9736 ( .A(n10395), .B(n7886), .S(n10159), .Z(n7885) );
  NAND2_X1 U9737 ( .A1(n7887), .A2(n8678), .ZN(n7884) );
  OAI211_X1 U9738 ( .C1(n8681), .C2(n7894), .A(n7885), .B(n7884), .ZN(P2_U3473) );
  INV_X1 U9739 ( .A(n7886), .ZN(n7891) );
  INV_X1 U9740 ( .A(n7887), .ZN(n7889) );
  OAI22_X1 U9741 ( .A1(n7889), .A2(n8523), .B1(n7888), .B2(n10097), .ZN(n7890)
         );
  OAI21_X1 U9742 ( .B1(n7891), .B2(n7890), .A(n8610), .ZN(n7893) );
  NAND2_X1 U9743 ( .A1(n10105), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n7892) );
  OAI211_X1 U9744 ( .C1(n7894), .C2(n8630), .A(n7893), .B(n7892), .ZN(P2_U3219) );
  INV_X1 U9745 ( .A(n7896), .ZN(n7897) );
  OR2_X1 U9746 ( .A1(n7898), .A2(n7897), .ZN(n8128) );
  XOR2_X1 U9747 ( .A(n7895), .B(n8128), .Z(n7899) );
  AOI222_X1 U9748 ( .A1(n8623), .A2(n7899), .B1(n8608), .B2(n8620), .C1(n8307), 
        .C2(n8618), .ZN(n8685) );
  XOR2_X1 U9749 ( .A(n8128), .B(n7900), .Z(n8683) );
  AOI22_X1 U9750 ( .A1(n10105), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n8626), .B2(
        n7901), .ZN(n7902) );
  OAI21_X1 U9751 ( .B1(n7903), .B2(n8560), .A(n7902), .ZN(n7904) );
  AOI21_X1 U9752 ( .B1(n8683), .B2(n8562), .A(n7904), .ZN(n7905) );
  OAI21_X1 U9753 ( .B1(n8685), .B2(n10105), .A(n7905), .ZN(P2_U3218) );
  INV_X1 U9754 ( .A(n7906), .ZN(n8165) );
  OAI222_X1 U9755 ( .A1(P1_U3086), .A2(n5824), .B1(n9738), .B2(n8165), .C1(
        n9735), .C2(n5647), .ZN(P1_U3331) );
  XNOR2_X1 U9756 ( .A(n8750), .B(n8189), .ZN(n7907) );
  NAND2_X1 U9757 ( .A1(n7907), .A2(n8595), .ZN(n8277) );
  INV_X1 U9758 ( .A(n7907), .ZN(n7908) );
  NAND2_X1 U9759 ( .A1(n7908), .A2(n8621), .ZN(n7909) );
  NAND2_X1 U9760 ( .A1(n8277), .A2(n7909), .ZN(n7914) );
  NAND2_X1 U9761 ( .A1(n7911), .A2(n7910), .ZN(n7912) );
  INV_X1 U9762 ( .A(n8167), .ZN(n8280) );
  AOI21_X1 U9763 ( .B1(n7914), .B2(n7913), .A(n8280), .ZN(n7920) );
  NAND2_X1 U9764 ( .A1(n8300), .A2(n8607), .ZN(n7915) );
  NAND2_X1 U9765 ( .A1(P2_U3151), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n8404) );
  OAI211_X1 U9766 ( .C1(n7916), .C2(n8297), .A(n7915), .B(n8404), .ZN(n7917)
         );
  AOI21_X1 U9767 ( .B1(n8611), .B2(n8295), .A(n7917), .ZN(n7919) );
  NAND2_X1 U9768 ( .A1(n8750), .A2(n8263), .ZN(n7918) );
  OAI211_X1 U9769 ( .C1(n7920), .C2(n8267), .A(n7919), .B(n7918), .ZN(P2_U3168) );
  NOR2_X1 U9770 ( .A1(n7921), .A2(n10097), .ZN(n8471) );
  NOR2_X1 U9771 ( .A1(n7922), .A2(n8560), .ZN(n7923) );
  AOI211_X1 U9772 ( .C1(n10105), .C2(P2_REG2_REG_29__SCAN_IN), .A(n8471), .B(
        n7923), .ZN(n7924) );
  OAI211_X1 U9773 ( .C1(n7927), .C2(n7926), .A(n7925), .B(n7924), .ZN(P2_U3204) );
  NAND2_X1 U9774 ( .A1(n7929), .A2(n7928), .ZN(n7930) );
  INV_X1 U9775 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n9092) );
  MUX2_X1 U9776 ( .A(n9092), .B(n8770), .S(n7936), .Z(n7932) );
  INV_X1 U9777 ( .A(SI_30_), .ZN(n10339) );
  NAND2_X1 U9778 ( .A1(n7932), .A2(n10339), .ZN(n7935) );
  INV_X1 U9779 ( .A(n7932), .ZN(n7933) );
  NAND2_X1 U9780 ( .A1(n7933), .A2(SI_30_), .ZN(n7934) );
  AND2_X1 U9781 ( .A1(n7935), .A2(n7934), .ZN(n8071) );
  MUX2_X1 U9782 ( .A(n7333), .B(n6714), .S(n7936), .Z(n7937) );
  XNOR2_X1 U9783 ( .A(n7937), .B(SI_31_), .ZN(n7938) );
  NAND2_X1 U9784 ( .A1(n8961), .A2(n6203), .ZN(n7941) );
  OR2_X1 U9785 ( .A1(n8075), .A2(n6714), .ZN(n7940) );
  INV_X1 U9786 ( .A(n7942), .ZN(n10094) );
  NOR2_X1 U9787 ( .A1(n8146), .A2(n10094), .ZN(n8092) );
  NAND2_X1 U9788 ( .A1(n7943), .A2(n6888), .ZN(n7944) );
  NAND2_X1 U9789 ( .A1(n5052), .A2(n7944), .ZN(n7945) );
  NAND2_X1 U9790 ( .A1(n7945), .A2(n8087), .ZN(n7952) );
  INV_X1 U9791 ( .A(n7946), .ZN(n7947) );
  OAI21_X1 U9792 ( .B1(n7952), .B2(n7947), .A(n7949), .ZN(n7948) );
  MUX2_X1 U9793 ( .A(n7949), .B(n7948), .S(n8087), .Z(n7961) );
  AOI21_X1 U9794 ( .B1(n7952), .B2(n7951), .A(n8111), .ZN(n7960) );
  OAI21_X1 U9795 ( .B1(n7955), .B2(n7954), .A(n7962), .ZN(n7958) );
  NAND2_X1 U9796 ( .A1(n7969), .A2(n7956), .ZN(n7957) );
  MUX2_X1 U9797 ( .A(n7958), .B(n7957), .S(n8087), .Z(n7959) );
  INV_X1 U9798 ( .A(n7962), .ZN(n7964) );
  OAI211_X1 U9799 ( .C1(n7973), .C2(n7964), .A(n7975), .B(n7963), .ZN(n7968)
         );
  NAND2_X1 U9800 ( .A1(n7974), .A2(n7970), .ZN(n7966) );
  NAND2_X1 U9801 ( .A1(n7966), .A2(n7965), .ZN(n7967) );
  NAND2_X1 U9802 ( .A1(n7968), .A2(n7967), .ZN(n7978) );
  INV_X1 U9803 ( .A(n7969), .ZN(n7972) );
  OAI211_X1 U9804 ( .C1(n7973), .C2(n7972), .A(n7971), .B(n7970), .ZN(n7976)
         );
  AOI21_X1 U9805 ( .B1(n7976), .B2(n7975), .A(n4872), .ZN(n7977) );
  MUX2_X1 U9806 ( .A(n7978), .B(n7977), .S(n8090), .Z(n7980) );
  INV_X1 U9807 ( .A(n7981), .ZN(n7989) );
  INV_X1 U9808 ( .A(n7982), .ZN(n7996) );
  OAI211_X1 U9809 ( .C1(n7984), .C2(n7989), .A(n7996), .B(n7983), .ZN(n7991)
         );
  AND2_X1 U9810 ( .A1(n7986), .A2(n7985), .ZN(n7988) );
  OAI211_X1 U9811 ( .C1(n7989), .C2(n7988), .A(n7993), .B(n7987), .ZN(n7990)
         );
  MUX2_X1 U9812 ( .A(n7991), .B(n7990), .S(n8090), .Z(n7992) );
  INV_X1 U9813 ( .A(n7995), .ZN(n7994) );
  INV_X1 U9814 ( .A(n7997), .ZN(n7998) );
  NAND2_X1 U9815 ( .A1(n8000), .A2(n7999), .ZN(n8002) );
  MUX2_X1 U9816 ( .A(n8002), .B(n8001), .S(n8090), .Z(n8003) );
  NAND2_X1 U9817 ( .A1(n8004), .A2(n8003), .ZN(n8009) );
  MUX2_X1 U9818 ( .A(n8308), .B(n8005), .S(n8087), .Z(n8006) );
  NAND2_X1 U9819 ( .A1(n8009), .A2(n8008), .ZN(n8010) );
  MUX2_X1 U9820 ( .A(n8013), .B(n8012), .S(n8087), .Z(n8014) );
  INV_X1 U9821 ( .A(n8015), .ZN(n8016) );
  NAND2_X1 U9822 ( .A1(n8024), .A2(n8016), .ZN(n8019) );
  INV_X1 U9823 ( .A(n8017), .ZN(n8018) );
  MUX2_X1 U9824 ( .A(n8019), .B(n8018), .S(n8090), .Z(n8021) );
  NOR2_X1 U9825 ( .A1(n8021), .A2(n8020), .ZN(n8022) );
  NAND2_X1 U9826 ( .A1(n8028), .A2(n8024), .ZN(n8030) );
  NAND2_X1 U9827 ( .A1(n8034), .A2(n8025), .ZN(n8026) );
  AOI21_X1 U9828 ( .B1(n8028), .B2(n8027), .A(n8026), .ZN(n8029) );
  NAND2_X1 U9829 ( .A1(n8039), .A2(n8035), .ZN(n8031) );
  AND2_X1 U9830 ( .A1(n8035), .A2(n8034), .ZN(n8038) );
  INV_X1 U9831 ( .A(n8036), .ZN(n8037) );
  NAND2_X1 U9832 ( .A1(n8045), .A2(n8043), .ZN(n8041) );
  NAND2_X1 U9833 ( .A1(n8048), .A2(n8039), .ZN(n8040) );
  MUX2_X1 U9834 ( .A(n8041), .B(n8040), .S(n8090), .Z(n8042) );
  INV_X1 U9835 ( .A(n8050), .ZN(n8046) );
  INV_X1 U9836 ( .A(n8109), .ZN(n8052) );
  NAND2_X1 U9837 ( .A1(n8548), .A2(n8048), .ZN(n8049) );
  INV_X1 U9838 ( .A(n8547), .ZN(n8657) );
  AND2_X1 U9839 ( .A1(n8107), .A2(n8052), .ZN(n8054) );
  NOR2_X1 U9840 ( .A1(n8056), .A2(n4886), .ZN(n8053) );
  MUX2_X1 U9841 ( .A(n8054), .B(n8053), .S(n8090), .Z(n8055) );
  INV_X1 U9842 ( .A(n8056), .ZN(n8108) );
  MUX2_X1 U9843 ( .A(n8108), .B(n8107), .S(n8090), .Z(n8057) );
  INV_X1 U9844 ( .A(n8064), .ZN(n8058) );
  MUX2_X1 U9845 ( .A(n8060), .B(n8059), .S(n8090), .Z(n8061) );
  NAND2_X1 U9846 ( .A1(n8066), .A2(n8067), .ZN(n8106) );
  INV_X1 U9847 ( .A(n8062), .ZN(n8063) );
  MUX2_X1 U9848 ( .A(n8064), .B(n8063), .S(n8090), .Z(n8065) );
  MUX2_X1 U9849 ( .A(n8067), .B(n8066), .S(n8087), .Z(n8068) );
  INV_X1 U9850 ( .A(n8068), .ZN(n8069) );
  MUX2_X1 U9851 ( .A(n8085), .B(n8488), .S(n8087), .Z(n8079) );
  OR2_X1 U9852 ( .A1(n8105), .A2(n8079), .ZN(n8070) );
  NAND2_X1 U9853 ( .A1(n8080), .A2(n8070), .ZN(n8086) );
  NAND2_X1 U9854 ( .A1(n8086), .A2(n8488), .ZN(n8078) );
  NAND2_X1 U9855 ( .A1(n9091), .A2(n6203), .ZN(n8077) );
  OR2_X1 U9856 ( .A1(n8075), .A2(n8770), .ZN(n8076) );
  INV_X1 U9857 ( .A(n8305), .ZN(n8083) );
  NOR2_X1 U9858 ( .A1(n8080), .A2(n8079), .ZN(n8081) );
  NOR2_X1 U9859 ( .A1(n8691), .A2(n8082), .ZN(n8104) );
  NAND2_X1 U9860 ( .A1(n8695), .A2(n8083), .ZN(n8136) );
  NAND2_X1 U9861 ( .A1(n8136), .A2(n8084), .ZN(n8095) );
  AOI21_X1 U9862 ( .B1(n8086), .B2(n8085), .A(n8095), .ZN(n8089) );
  NAND2_X1 U9863 ( .A1(n8137), .A2(n8087), .ZN(n8088) );
  NOR2_X1 U9864 ( .A1(n8695), .A2(n8470), .ZN(n8096) );
  NOR2_X1 U9865 ( .A1(n8691), .A2(n8096), .ZN(n8097) );
  NOR2_X1 U9866 ( .A1(n8095), .A2(n8097), .ZN(n8098) );
  NAND2_X1 U9867 ( .A1(n8099), .A2(n8098), .ZN(n8102) );
  INV_X1 U9868 ( .A(n8137), .ZN(n8100) );
  NAND2_X1 U9869 ( .A1(n8100), .A2(n8691), .ZN(n8101) );
  NAND2_X1 U9870 ( .A1(n8102), .A2(n8101), .ZN(n8103) );
  NAND2_X1 U9871 ( .A1(n8103), .A2(n6888), .ZN(n8143) );
  INV_X1 U9872 ( .A(n8104), .ZN(n8140) );
  INV_X1 U9873 ( .A(n8105), .ZN(n8139) );
  INV_X1 U9874 ( .A(n8106), .ZN(n8492) );
  NAND2_X1 U9875 ( .A1(n8108), .A2(n8107), .ZN(n8520) );
  OR2_X1 U9876 ( .A1(n8109), .A2(n4886), .ZN(n8531) );
  INV_X1 U9877 ( .A(n8531), .ZN(n8529) );
  INV_X1 U9878 ( .A(n8110), .ZN(n8556) );
  INV_X1 U9879 ( .A(n8614), .ZN(n8616) );
  AND2_X1 U9880 ( .A1(n4612), .A2(n8114), .ZN(n8116) );
  NAND4_X1 U9881 ( .A1(n4533), .A2(n8117), .A3(n8116), .A4(n8115), .ZN(n8119)
         );
  NOR2_X1 U9882 ( .A1(n8119), .A2(n8118), .ZN(n8121) );
  NAND3_X1 U9883 ( .A1(n8121), .A2(n4860), .A3(n8120), .ZN(n8122) );
  OR4_X1 U9884 ( .A1(n8125), .A2(n8124), .A3(n8123), .A4(n8122), .ZN(n8126) );
  NOR3_X1 U9885 ( .A1(n5022), .A2(n8127), .A3(n8126), .ZN(n8129) );
  NAND3_X1 U9886 ( .A1(n8616), .A2(n8129), .A3(n8128), .ZN(n8130) );
  NOR4_X1 U9887 ( .A1(n8576), .A2(n8591), .A3(n8606), .A4(n8130), .ZN(n8131)
         );
  NAND4_X1 U9888 ( .A1(n8529), .A2(n8556), .A3(n5102), .A4(n8131), .ZN(n8133)
         );
  INV_X1 U9889 ( .A(n8548), .ZN(n8132) );
  NOR3_X1 U9890 ( .A1(n8520), .A2(n8133), .A3(n8132), .ZN(n8134) );
  AND4_X1 U9891 ( .A1(n8492), .A2(n8501), .A3(n8514), .A4(n8134), .ZN(n8135)
         );
  AND4_X1 U9892 ( .A1(n8137), .A2(n8136), .A3(n8135), .A4(n8484), .ZN(n8138)
         );
  NAND3_X1 U9893 ( .A1(n8140), .A2(n8139), .A3(n8138), .ZN(n8141) );
  NAND2_X1 U9894 ( .A1(n8143), .A2(n8142), .ZN(n8150) );
  INV_X1 U9895 ( .A(n8146), .ZN(n8144) );
  NAND3_X1 U9896 ( .A1(n8144), .A2(n8444), .A3(n8145), .ZN(n8149) );
  NAND3_X1 U9897 ( .A1(n8150), .A2(n8145), .A3(n8463), .ZN(n8148) );
  AOI21_X1 U9898 ( .B1(n8146), .B2(n8463), .A(n8154), .ZN(n8147) );
  OAI211_X1 U9899 ( .C1(n8150), .C2(n8149), .A(n8148), .B(n8147), .ZN(n8157)
         );
  NAND3_X1 U9900 ( .A1(n8152), .A2(n8151), .A3(n8779), .ZN(n8153) );
  OAI211_X1 U9901 ( .C1(n8155), .C2(n8154), .A(n8153), .B(P2_B_REG_SCAN_IN), 
        .ZN(n8156) );
  OAI21_X1 U9902 ( .B1(n8158), .B2(n8157), .A(n8156), .ZN(P2_U3296) );
  INV_X1 U9903 ( .A(n8159), .ZN(n9725) );
  OAI222_X1 U9904 ( .A1(n8787), .A2(n9725), .B1(n8161), .B2(P2_U3151), .C1(
        n8160), .C2(n8765), .ZN(P2_U3266) );
  INV_X1 U9905 ( .A(n8162), .ZN(n8780) );
  OAI222_X1 U9906 ( .A1(n9735), .A2(n8164), .B1(n9738), .B2(n8780), .C1(n8163), 
        .C2(P1_U3086), .ZN(P1_U3328) );
  OAI222_X1 U9907 ( .A1(P2_U3151), .A2(n8166), .B1(n8787), .B2(n8165), .C1(
        n8765), .C2(n6204), .ZN(P2_U3271) );
  INV_X1 U9908 ( .A(n9091), .ZN(n8771) );
  OAI222_X1 U9909 ( .A1(n9735), .A2(n9092), .B1(n9730), .B2(n8771), .C1(n5168), 
        .C2(P1_U3086), .ZN(P1_U3325) );
  NAND2_X1 U9910 ( .A1(n8167), .A2(n8277), .ZN(n8168) );
  XNOR2_X1 U9911 ( .A(n8671), .B(n8189), .ZN(n8169) );
  XNOR2_X1 U9912 ( .A(n8169), .B(n8607), .ZN(n8278) );
  NAND2_X1 U9913 ( .A1(n8168), .A2(n8278), .ZN(n8281) );
  NAND2_X1 U9914 ( .A1(n8169), .A2(n8225), .ZN(n8170) );
  NAND2_X1 U9915 ( .A1(n8281), .A2(n8170), .ZN(n8221) );
  XNOR2_X1 U9916 ( .A(n8666), .B(n8189), .ZN(n8171) );
  INV_X1 U9917 ( .A(n8171), .ZN(n8172) );
  NAND2_X1 U9918 ( .A1(n8172), .A2(n8569), .ZN(n8222) );
  XNOR2_X1 U9919 ( .A(n8736), .B(n8196), .ZN(n8173) );
  NAND2_X1 U9920 ( .A1(n8173), .A2(n8580), .ZN(n8257) );
  INV_X1 U9921 ( .A(n8173), .ZN(n8174) );
  NAND2_X1 U9922 ( .A1(n8174), .A2(n8554), .ZN(n8258) );
  XNOR2_X1 U9923 ( .A(n8175), .B(n8196), .ZN(n8176) );
  XNOR2_X1 U9924 ( .A(n8176), .B(n8306), .ZN(n8232) );
  NAND2_X1 U9925 ( .A1(n8231), .A2(n8232), .ZN(n8230) );
  INV_X1 U9926 ( .A(n8176), .ZN(n8177) );
  NAND2_X1 U9927 ( .A1(n8177), .A2(n8306), .ZN(n8178) );
  XNOR2_X1 U9928 ( .A(n8547), .B(n8196), .ZN(n8179) );
  XNOR2_X1 U9929 ( .A(n8179), .B(n8533), .ZN(n8268) );
  NAND2_X1 U9930 ( .A1(n8179), .A2(n8533), .ZN(n8180) );
  XNOR2_X1 U9931 ( .A(n8725), .B(n8196), .ZN(n8183) );
  INV_X1 U9932 ( .A(n8183), .ZN(n8181) );
  XNOR2_X1 U9933 ( .A(n8719), .B(n8189), .ZN(n8185) );
  NAND2_X1 U9934 ( .A1(n8185), .A2(n8242), .ZN(n8188) );
  INV_X1 U9935 ( .A(n8185), .ZN(n8186) );
  NAND2_X1 U9936 ( .A1(n8186), .A2(n8534), .ZN(n8187) );
  NAND2_X1 U9937 ( .A1(n8188), .A2(n8187), .ZN(n8247) );
  XNOR2_X1 U9938 ( .A(n8714), .B(n8189), .ZN(n8190) );
  XNOR2_X1 U9939 ( .A(n8190), .B(n8521), .ZN(n8238) );
  XNOR2_X1 U9940 ( .A(n8708), .B(n8196), .ZN(n8192) );
  NAND2_X1 U9941 ( .A1(n8291), .A2(n8193), .ZN(n8204) );
  XNOR2_X1 U9942 ( .A(n8702), .B(n8196), .ZN(n8194) );
  XNOR2_X1 U9943 ( .A(n8194), .B(n8502), .ZN(n8203) );
  XNOR2_X1 U9944 ( .A(n8484), .B(n8196), .ZN(n8197) );
  NAND2_X1 U9945 ( .A1(n8478), .A2(n8300), .ZN(n8199) );
  AOI22_X1 U9946 ( .A1(n8486), .A2(n8295), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3151), .ZN(n8198) );
  OAI211_X1 U9947 ( .C1(n8200), .C2(n8297), .A(n8199), .B(n8198), .ZN(n8201)
         );
  AOI21_X1 U9948 ( .B1(n8635), .B2(n8263), .A(n8201), .ZN(n8202) );
  INV_X1 U9949 ( .A(n8204), .ZN(n8206) );
  INV_X1 U9950 ( .A(n8267), .ZN(n8205) );
  AOI22_X1 U9951 ( .A1(n8496), .A2(n8295), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3151), .ZN(n8207) );
  OAI21_X1 U9952 ( .B1(n8293), .B2(n8297), .A(n8207), .ZN(n8208) );
  AOI21_X1 U9953 ( .B1(n8300), .B2(n8494), .A(n8208), .ZN(n8209) );
  OAI211_X1 U9954 ( .C1(n8211), .C2(n8303), .A(n8210), .B(n8209), .ZN(P2_U3154) );
  OAI21_X1 U9955 ( .B1(n8272), .B2(n8213), .A(n8212), .ZN(n8214) );
  NAND2_X1 U9956 ( .A1(n8214), .A2(n8205), .ZN(n8219) );
  INV_X1 U9957 ( .A(n8537), .ZN(n8216) );
  AOI22_X1 U9958 ( .A1(n8533), .A2(n8284), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3151), .ZN(n8215) );
  OAI21_X1 U9959 ( .B1(n8216), .B2(n8252), .A(n8215), .ZN(n8217) );
  AOI21_X1 U9960 ( .B1(n8534), .B2(n8300), .A(n8217), .ZN(n8218) );
  OAI211_X1 U9961 ( .C1(n8220), .C2(n8303), .A(n8219), .B(n8218), .ZN(P2_U3156) );
  NAND2_X1 U9962 ( .A1(n4538), .A2(n8222), .ZN(n8223) );
  XNOR2_X1 U9963 ( .A(n8221), .B(n8223), .ZN(n8229) );
  NAND2_X1 U9964 ( .A1(n8580), .A2(n8300), .ZN(n8224) );
  NAND2_X1 U9965 ( .A1(P2_U3151), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8461) );
  OAI211_X1 U9966 ( .C1(n8225), .C2(n8297), .A(n8224), .B(n8461), .ZN(n8226)
         );
  AOI21_X1 U9967 ( .B1(n8583), .B2(n8295), .A(n8226), .ZN(n8228) );
  NAND2_X1 U9968 ( .A1(n8666), .A2(n8263), .ZN(n8227) );
  OAI211_X1 U9969 ( .C1(n8229), .C2(n8267), .A(n8228), .B(n8227), .ZN(P2_U3159) );
  OAI21_X1 U9970 ( .B1(n8232), .B2(n8231), .A(n8230), .ZN(n8233) );
  NAND2_X1 U9971 ( .A1(n8233), .A2(n8205), .ZN(n8237) );
  AOI22_X1 U9972 ( .A1(n8533), .A2(n8300), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3151), .ZN(n8234) );
  OAI21_X1 U9973 ( .B1(n8554), .B2(n8297), .A(n8234), .ZN(n8235) );
  AOI21_X1 U9974 ( .B1(n8558), .B2(n8295), .A(n8235), .ZN(n8236) );
  OAI211_X1 U9975 ( .C1(n8734), .C2(n8303), .A(n8237), .B(n8236), .ZN(P2_U3163) );
  INV_X1 U9976 ( .A(n8714), .ZN(n8246) );
  NOR3_X1 U9977 ( .A1(n8250), .A2(n8239), .A3(n8238), .ZN(n8240) );
  OAI21_X1 U9978 ( .B1(n4544), .B2(n8240), .A(n8205), .ZN(n8245) );
  AOI22_X1 U9979 ( .A1(n8511), .A2(n8295), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3151), .ZN(n8241) );
  OAI21_X1 U9980 ( .B1(n8242), .B2(n8297), .A(n8241), .ZN(n8243) );
  AOI21_X1 U9981 ( .B1(n8509), .B2(n8300), .A(n8243), .ZN(n8244) );
  OAI211_X1 U9982 ( .C1(n8246), .C2(n8303), .A(n8245), .B(n8244), .ZN(P2_U3165) );
  AND3_X1 U9983 ( .A1(n8212), .A2(n8248), .A3(n8247), .ZN(n8249) );
  OAI21_X1 U9984 ( .B1(n8250), .B2(n8249), .A(n8205), .ZN(n8256) );
  INV_X1 U9985 ( .A(n8526), .ZN(n8253) );
  AOI22_X1 U9986 ( .A1(n8541), .A2(n8284), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3151), .ZN(n8251) );
  OAI21_X1 U9987 ( .B1(n8253), .B2(n8252), .A(n8251), .ZN(n8254) );
  AOI21_X1 U9988 ( .B1(n8300), .B2(n8521), .A(n8254), .ZN(n8255) );
  OAI211_X1 U9989 ( .C1(n8524), .C2(n8303), .A(n8256), .B(n8255), .ZN(P2_U3169) );
  NAND2_X1 U9990 ( .A1(n8258), .A2(n8257), .ZN(n8259) );
  XNOR2_X1 U9991 ( .A(n4602), .B(n8259), .ZN(n8266) );
  INV_X1 U9992 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n8260) );
  OAI22_X1 U9993 ( .A1(n8597), .A2(n8297), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8260), .ZN(n8262) );
  NOR2_X1 U9994 ( .A1(n8306), .A2(n8286), .ZN(n8261) );
  AOI211_X1 U9995 ( .C1(n8566), .C2(n8295), .A(n8262), .B(n8261), .ZN(n8265)
         );
  NAND2_X1 U9996 ( .A1(n8736), .A2(n8263), .ZN(n8264) );
  OAI211_X1 U9997 ( .C1(n8266), .C2(n8267), .A(n8265), .B(n8264), .ZN(P2_U3173) );
  AOI21_X1 U9998 ( .B1(n8269), .B2(n8268), .A(n8267), .ZN(n8271) );
  NAND2_X1 U9999 ( .A1(n8271), .A2(n8270), .ZN(n8276) );
  INV_X1 U10000 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n10281) );
  OAI22_X1 U10001 ( .A1(n8306), .A2(n8297), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10281), .ZN(n8274) );
  NOR2_X1 U10002 ( .A1(n8272), .A2(n8286), .ZN(n8273) );
  AOI211_X1 U10003 ( .C1(n8543), .C2(n8295), .A(n8274), .B(n8273), .ZN(n8275)
         );
  OAI211_X1 U10004 ( .C1(n8657), .C2(n8303), .A(n8276), .B(n8275), .ZN(
        P2_U3175) );
  INV_X1 U10005 ( .A(n8671), .ZN(n8290) );
  INV_X1 U10006 ( .A(n8277), .ZN(n8279) );
  NOR3_X1 U10007 ( .A1(n8280), .A2(n8279), .A3(n8278), .ZN(n8283) );
  INV_X1 U10008 ( .A(n8281), .ZN(n8282) );
  OAI21_X1 U10009 ( .B1(n8283), .B2(n8282), .A(n8205), .ZN(n8289) );
  NAND2_X1 U10010 ( .A1(n8284), .A2(n8621), .ZN(n8285) );
  NAND2_X1 U10011 ( .A1(P2_U3151), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8435) );
  OAI211_X1 U10012 ( .C1(n8597), .C2(n8286), .A(n8285), .B(n8435), .ZN(n8287)
         );
  AOI21_X1 U10013 ( .B1(n8599), .B2(n8295), .A(n8287), .ZN(n8288) );
  OAI211_X1 U10014 ( .C1(n8290), .C2(n8303), .A(n8289), .B(n8288), .ZN(
        P2_U3178) );
  OAI21_X1 U10015 ( .B1(n8293), .B2(n8292), .A(n8291), .ZN(n8294) );
  NAND2_X1 U10016 ( .A1(n8294), .A2(n8205), .ZN(n8302) );
  AOI22_X1 U10017 ( .A1(n8505), .A2(n8295), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3151), .ZN(n8296) );
  OAI21_X1 U10018 ( .B1(n8298), .B2(n8297), .A(n8296), .ZN(n8299) );
  AOI21_X1 U10019 ( .B1(n8300), .B2(n8502), .A(n8299), .ZN(n8301) );
  OAI211_X1 U10020 ( .C1(n8304), .C2(n8303), .A(n8302), .B(n8301), .ZN(
        P2_U3180) );
  MUX2_X1 U10021 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n8305), .S(P2_U3893), .Z(
        P2_U3521) );
  MUX2_X1 U10022 ( .A(n8478), .B(P2_DATAO_REG_29__SCAN_IN), .S(n8428), .Z(
        P2_U3520) );
  MUX2_X1 U10023 ( .A(n8494), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8428), .Z(
        P2_U3519) );
  MUX2_X1 U10024 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8502), .S(P2_U3893), .Z(
        P2_U3518) );
  MUX2_X1 U10025 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n8509), .S(P2_U3893), .Z(
        P2_U3517) );
  MUX2_X1 U10026 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n8521), .S(P2_U3893), .Z(
        P2_U3516) );
  MUX2_X1 U10027 ( .A(n8541), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8428), .Z(
        P2_U3514) );
  MUX2_X1 U10028 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8533), .S(P2_U3893), .Z(
        P2_U3513) );
  MUX2_X1 U10029 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n6486), .S(P2_U3893), .Z(
        P2_U3512) );
  MUX2_X1 U10030 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8580), .S(P2_U3893), .Z(
        P2_U3511) );
  MUX2_X1 U10031 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n8569), .S(P2_U3893), .Z(
        P2_U3510) );
  MUX2_X1 U10032 ( .A(n8607), .B(P2_DATAO_REG_18__SCAN_IN), .S(n8428), .Z(
        P2_U3509) );
  MUX2_X1 U10033 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8621), .S(P2_U3893), .Z(
        P2_U3508) );
  MUX2_X1 U10034 ( .A(n8608), .B(P2_DATAO_REG_16__SCAN_IN), .S(n8428), .Z(
        P2_U3507) );
  MUX2_X1 U10035 ( .A(n8619), .B(P2_DATAO_REG_15__SCAN_IN), .S(n8428), .Z(
        P2_U3506) );
  MUX2_X1 U10036 ( .A(n8307), .B(P2_DATAO_REG_14__SCAN_IN), .S(n8428), .Z(
        P2_U3505) );
  MUX2_X1 U10037 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n8308), .S(P2_U3893), .Z(
        P2_U3504) );
  MUX2_X1 U10038 ( .A(n8309), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8428), .Z(
        P2_U3503) );
  MUX2_X1 U10039 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n8310), .S(P2_U3893), .Z(
        P2_U3502) );
  MUX2_X1 U10040 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n8311), .S(P2_U3893), .Z(
        P2_U3501) );
  MUX2_X1 U10041 ( .A(n8312), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8428), .Z(
        P2_U3500) );
  MUX2_X1 U10042 ( .A(n8313), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8428), .Z(
        P2_U3499) );
  MUX2_X1 U10043 ( .A(n8314), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8428), .Z(
        P2_U3498) );
  MUX2_X1 U10044 ( .A(n8315), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8428), .Z(
        P2_U3497) );
  MUX2_X1 U10045 ( .A(n8316), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8428), .Z(
        P2_U3496) );
  MUX2_X1 U10046 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n6267), .S(P2_U3893), .Z(
        P2_U3495) );
  MUX2_X1 U10047 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(n8317), .S(P2_U3893), .Z(
        P2_U3494) );
  MUX2_X1 U10048 ( .A(n8318), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8428), .Z(
        P2_U3493) );
  INV_X1 U10049 ( .A(n6224), .ZN(n8319) );
  MUX2_X1 U10050 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n8319), .S(P2_U3893), .Z(
        P2_U3492) );
  AOI22_X1 U10051 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n8350), .B1(n8347), .B2(
        n8333), .ZN(n8323) );
  AOI21_X1 U10052 ( .B1(n4604), .B2(n8323), .A(n8346), .ZN(n8345) );
  AOI22_X1 U10053 ( .A1(P2_REG1_REG_14__SCAN_IN), .A2(n8347), .B1(n8350), .B2(
        n10395), .ZN(n8329) );
  NAND2_X1 U10054 ( .A1(n8325), .A2(n8324), .ZN(n8327) );
  NAND2_X1 U10055 ( .A1(n8327), .A2(n8326), .ZN(n8328) );
  NAND2_X1 U10056 ( .A1(n8329), .A2(n8328), .ZN(n8349) );
  OAI21_X1 U10057 ( .B1(n8329), .B2(n8328), .A(n8349), .ZN(n8343) );
  NAND2_X1 U10058 ( .A1(n10067), .A2(P2_ADDR_REG_14__SCAN_IN), .ZN(n8331) );
  OAI211_X1 U10059 ( .C1(n10051), .C2(n8347), .A(n8331), .B(n8330), .ZN(n8342)
         );
  INV_X1 U10060 ( .A(n8332), .ZN(n8338) );
  MUX2_X1 U10061 ( .A(n8333), .B(n10395), .S(n8779), .Z(n8334) );
  NAND2_X1 U10062 ( .A1(n8334), .A2(n8350), .ZN(n8361) );
  INV_X1 U10063 ( .A(n8334), .ZN(n8335) );
  NAND2_X1 U10064 ( .A1(n8335), .A2(n8347), .ZN(n8336) );
  AND2_X1 U10065 ( .A1(n8361), .A2(n8336), .ZN(n8337) );
  OAI21_X1 U10066 ( .B1(n8339), .B2(n8338), .A(n8337), .ZN(n8362) );
  OR3_X1 U10067 ( .A1(n8339), .A2(n8338), .A3(n8337), .ZN(n8340) );
  AOI21_X1 U10068 ( .B1(n8362), .B2(n8340), .A(n10079), .ZN(n8341) );
  AOI211_X1 U10069 ( .C1(n8343), .C2(n10084), .A(n8342), .B(n8341), .ZN(n8344)
         );
  OAI21_X1 U10070 ( .B1(n8345), .B2(n10089), .A(n8344), .ZN(P2_U3196) );
  NOR2_X1 U10071 ( .A1(n8356), .A2(n8348), .ZN(n8372) );
  AOI21_X1 U10072 ( .B1(n8356), .B2(n8348), .A(n8372), .ZN(n8369) );
  XNOR2_X1 U10073 ( .A(n8376), .B(n8371), .ZN(n8351) );
  NAND2_X1 U10074 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n8351), .ZN(n8378) );
  OAI21_X1 U10075 ( .B1(P2_REG1_REG_15__SCAN_IN), .B2(n8351), .A(n8378), .ZN(
        n8367) );
  NAND2_X1 U10076 ( .A1(n10069), .A2(n8371), .ZN(n8353) );
  OAI211_X1 U10077 ( .C1(n8354), .C2(n10049), .A(n8353), .B(n8352), .ZN(n8366)
         );
  MUX2_X1 U10078 ( .A(n8356), .B(n8355), .S(n8779), .Z(n8357) );
  NAND2_X1 U10079 ( .A1(n8357), .A2(n8371), .ZN(n8385) );
  INV_X1 U10080 ( .A(n8357), .ZN(n8358) );
  NAND2_X1 U10081 ( .A1(n8358), .A2(n8377), .ZN(n8359) );
  NAND2_X1 U10082 ( .A1(n8385), .A2(n8359), .ZN(n8360) );
  AOI21_X1 U10083 ( .B1(n8362), .B2(n8361), .A(n8360), .ZN(n8391) );
  INV_X1 U10084 ( .A(n8391), .ZN(n8364) );
  NAND3_X1 U10085 ( .A1(n8362), .A2(n8361), .A3(n8360), .ZN(n8363) );
  AOI21_X1 U10086 ( .B1(n8364), .B2(n8363), .A(n10079), .ZN(n8365) );
  AOI211_X1 U10087 ( .C1(n8367), .C2(n10084), .A(n8366), .B(n8365), .ZN(n8368)
         );
  OAI21_X1 U10088 ( .B1(n8369), .B2(n10089), .A(n8368), .ZN(P2_U3197) );
  NOR2_X1 U10089 ( .A1(n8371), .A2(n8370), .ZN(n8373) );
  AOI22_X1 U10090 ( .A1(P2_REG2_REG_16__SCAN_IN), .A2(n8402), .B1(n8399), .B2(
        n8624), .ZN(n8374) );
  NOR2_X1 U10091 ( .A1(n8375), .A2(n8374), .ZN(n8398) );
  AOI21_X1 U10092 ( .B1(n8375), .B2(n8374), .A(n8398), .ZN(n8397) );
  AOI22_X1 U10093 ( .A1(P2_REG1_REG_16__SCAN_IN), .A2(n8399), .B1(n8402), .B2(
        n8677), .ZN(n8381) );
  NAND2_X1 U10094 ( .A1(n8377), .A2(n8376), .ZN(n8379) );
  NAND2_X1 U10095 ( .A1(n8379), .A2(n8378), .ZN(n8380) );
  NAND2_X1 U10096 ( .A1(n8381), .A2(n8380), .ZN(n8401) );
  OAI21_X1 U10097 ( .B1(n8381), .B2(n8380), .A(n8401), .ZN(n8395) );
  NAND2_X1 U10098 ( .A1(n10069), .A2(n8402), .ZN(n8383) );
  OAI211_X1 U10099 ( .C1(n8384), .C2(n10049), .A(n8383), .B(n8382), .ZN(n8394)
         );
  INV_X1 U10100 ( .A(n8385), .ZN(n8390) );
  MUX2_X1 U10101 ( .A(n8624), .B(n8677), .S(n8779), .Z(n8386) );
  NAND2_X1 U10102 ( .A1(n8386), .A2(n8402), .ZN(n8407) );
  INV_X1 U10103 ( .A(n8386), .ZN(n8387) );
  NAND2_X1 U10104 ( .A1(n8387), .A2(n8399), .ZN(n8388) );
  AND2_X1 U10105 ( .A1(n8407), .A2(n8388), .ZN(n8389) );
  OAI21_X1 U10106 ( .B1(n8391), .B2(n8390), .A(n8389), .ZN(n8409) );
  OR3_X1 U10107 ( .A1(n8391), .A2(n8390), .A3(n8389), .ZN(n8392) );
  AOI21_X1 U10108 ( .B1(n8409), .B2(n8392), .A(n10079), .ZN(n8393) );
  AOI211_X1 U10109 ( .C1(n8395), .C2(n10084), .A(n8394), .B(n8393), .ZN(n8396)
         );
  OAI21_X1 U10110 ( .B1(n8397), .B2(n10089), .A(n8396), .ZN(P2_U3198) );
  XOR2_X1 U10111 ( .A(n8417), .B(n8430), .Z(n8400) );
  AOI21_X1 U10112 ( .B1(n10384), .B2(n8400), .A(n8418), .ZN(n8416) );
  NAND2_X1 U10113 ( .A1(P2_REG1_REG_17__SCAN_IN), .A2(n8403), .ZN(n8431) );
  OAI21_X1 U10114 ( .B1(P2_REG1_REG_17__SCAN_IN), .B2(n8403), .A(n8431), .ZN(
        n8414) );
  NAND2_X1 U10115 ( .A1(n10069), .A2(n8424), .ZN(n8405) );
  OAI211_X1 U10116 ( .C1(n8406), .C2(n10049), .A(n8405), .B(n8404), .ZN(n8413)
         );
  MUX2_X1 U10117 ( .A(n10384), .B(n8674), .S(n8779), .Z(n8423) );
  XNOR2_X1 U10118 ( .A(n8423), .B(n8424), .ZN(n8408) );
  AOI21_X1 U10119 ( .B1(n8409), .B2(n8407), .A(n8408), .ZN(n8422) );
  INV_X1 U10120 ( .A(n8422), .ZN(n8411) );
  NAND3_X1 U10121 ( .A1(n8409), .A2(n8408), .A3(n8407), .ZN(n8410) );
  AOI21_X1 U10122 ( .B1(n8411), .B2(n8410), .A(n10079), .ZN(n8412) );
  AOI211_X1 U10123 ( .C1(n8414), .C2(n10084), .A(n8413), .B(n8412), .ZN(n8415)
         );
  OAI21_X1 U10124 ( .B1(n8416), .B2(n10089), .A(n8415), .ZN(P2_U3199) );
  NOR2_X1 U10125 ( .A1(n8424), .A2(n8417), .ZN(n8419) );
  NAND2_X1 U10126 ( .A1(n8454), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n8443) );
  OAI21_X1 U10127 ( .B1(n8454), .B2(P2_REG2_REG_18__SCAN_IN), .A(n8443), .ZN(
        n8420) );
  AOI21_X1 U10128 ( .B1(n8421), .B2(n8420), .A(n4568), .ZN(n8442) );
  AOI21_X1 U10129 ( .B1(n8424), .B2(n8423), .A(n8422), .ZN(n8426) );
  MUX2_X1 U10130 ( .A(P2_REG2_REG_18__SCAN_IN), .B(P2_REG1_REG_18__SCAN_IN), 
        .S(n8779), .Z(n8425) );
  NOR2_X1 U10131 ( .A1(n8426), .A2(n8425), .ZN(n8448) );
  INV_X1 U10132 ( .A(n8448), .ZN(n8427) );
  NAND2_X1 U10133 ( .A1(n8426), .A2(n8425), .ZN(n8446) );
  NAND2_X1 U10134 ( .A1(n8427), .A2(n8446), .ZN(n8434) );
  OAI21_X1 U10135 ( .B1(n8434), .B2(n8428), .A(n10051), .ZN(n8440) );
  XNOR2_X1 U10136 ( .A(n8447), .B(P2_REG1_REG_18__SCAN_IN), .ZN(n8455) );
  NAND2_X1 U10137 ( .A1(n8430), .A2(n8429), .ZN(n8432) );
  NAND2_X1 U10138 ( .A1(n8432), .A2(n8431), .ZN(n8456) );
  XOR2_X1 U10139 ( .A(n8455), .B(n8456), .Z(n8433) );
  NOR2_X1 U10140 ( .A1(n8433), .A2(n9939), .ZN(n8439) );
  INV_X1 U10141 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n8437) );
  NAND3_X1 U10142 ( .A1(n8434), .A2(n10058), .A3(n8454), .ZN(n8436) );
  OAI211_X1 U10143 ( .C1(n10049), .C2(n8437), .A(n8436), .B(n8435), .ZN(n8438)
         );
  AOI211_X1 U10144 ( .C1(n8447), .C2(n8440), .A(n8439), .B(n8438), .ZN(n8441)
         );
  OAI21_X1 U10145 ( .B1(n8442), .B2(n10089), .A(n8441), .ZN(P2_U3200) );
  XNOR2_X1 U10146 ( .A(n8444), .B(P2_REG2_REG_19__SCAN_IN), .ZN(n8449) );
  XNOR2_X1 U10147 ( .A(n8445), .B(n8449), .ZN(n8468) );
  OAI21_X1 U10148 ( .B1(n8448), .B2(n8447), .A(n8446), .ZN(n8453) );
  XNOR2_X1 U10149 ( .A(n8463), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n8457) );
  INV_X1 U10150 ( .A(n8449), .ZN(n8451) );
  MUX2_X1 U10151 ( .A(n8457), .B(n8451), .S(n8450), .Z(n8452) );
  XNOR2_X1 U10152 ( .A(n8453), .B(n8452), .ZN(n8466) );
  AOI22_X1 U10153 ( .A1(n8456), .A2(n8455), .B1(P2_REG1_REG_18__SCAN_IN), .B2(
        n8454), .ZN(n8459) );
  INV_X1 U10154 ( .A(n8457), .ZN(n8458) );
  XNOR2_X1 U10155 ( .A(n8459), .B(n8458), .ZN(n8460) );
  NOR2_X1 U10156 ( .A1(n8460), .A2(n9939), .ZN(n8465) );
  NAND2_X1 U10157 ( .A1(n10067), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n8462) );
  OAI211_X1 U10158 ( .C1(n10051), .C2(n8463), .A(n8462), .B(n8461), .ZN(n8464)
         );
  OAI21_X1 U10159 ( .B1(n8468), .B2(n10089), .A(n8467), .ZN(P2_U3201) );
  NAND2_X1 U10160 ( .A1(n8691), .A2(n8627), .ZN(n8472) );
  AOI21_X1 U10161 ( .B1(n8692), .B2(n8610), .A(n8471), .ZN(n8474) );
  OAI211_X1 U10162 ( .C1(n10103), .C2(n8473), .A(n8472), .B(n8474), .ZN(
        P2_U3202) );
  NAND2_X1 U10163 ( .A1(n8695), .A2(n8627), .ZN(n8475) );
  OAI211_X1 U10164 ( .C1(n10103), .C2(n8476), .A(n8475), .B(n8474), .ZN(
        P2_U3203) );
  XNOR2_X1 U10165 ( .A(n8477), .B(n8484), .ZN(n8482) );
  NAND2_X1 U10166 ( .A1(n8478), .A2(n8620), .ZN(n8480) );
  OAI21_X1 U10167 ( .B1(n8485), .B2(n8484), .A(n8483), .ZN(n8636) );
  AOI22_X1 U10168 ( .A1(n8486), .A2(n8626), .B1(n10105), .B2(
        P2_REG2_REG_28__SCAN_IN), .ZN(n8487) );
  OAI21_X1 U10169 ( .B1(n8488), .B2(n8560), .A(n8487), .ZN(n8489) );
  AOI21_X1 U10170 ( .B1(n8636), .B2(n8562), .A(n8489), .ZN(n8490) );
  OAI21_X1 U10171 ( .B1(n8638), .B2(n10105), .A(n8490), .ZN(P2_U3205) );
  XNOR2_X1 U10172 ( .A(n8491), .B(n8492), .ZN(n8705) );
  MUX2_X1 U10173 ( .A(n8495), .B(n8700), .S(n8610), .Z(n8498) );
  AOI22_X1 U10174 ( .A1(n8702), .A2(n8627), .B1(n8626), .B2(n8496), .ZN(n8497)
         );
  XOR2_X1 U10175 ( .A(n8501), .B(n8500), .Z(n8503) );
  AOI222_X1 U10176 ( .A1(n8623), .A2(n8503), .B1(n8502), .B2(n8620), .C1(n8521), .C2(n8618), .ZN(n8706) );
  MUX2_X1 U10177 ( .A(n8504), .B(n8706), .S(n10103), .Z(n8507) );
  AOI22_X1 U10178 ( .A1(n8708), .A2(n8627), .B1(n8626), .B2(n8505), .ZN(n8506)
         );
  OAI211_X1 U10179 ( .C1(n8711), .C2(n8630), .A(n8507), .B(n8506), .ZN(
        P2_U3207) );
  XNOR2_X1 U10180 ( .A(n8508), .B(n8514), .ZN(n8510) );
  AOI222_X1 U10181 ( .A1(n8623), .A2(n8510), .B1(n8509), .B2(n8620), .C1(n8534), .C2(n8618), .ZN(n8712) );
  AOI22_X1 U10182 ( .A1(n8714), .A2(n8512), .B1(n8626), .B2(n8511), .ZN(n8513)
         );
  AOI21_X1 U10183 ( .B1(n8712), .B2(n8513), .A(n10105), .ZN(n8518) );
  XNOR2_X1 U10184 ( .A(n8515), .B(n8514), .ZN(n8717) );
  OAI22_X1 U10185 ( .A1(n8717), .A2(n8630), .B1(n8516), .B2(n10103), .ZN(n8517) );
  OR2_X1 U10186 ( .A1(n8518), .A2(n8517), .ZN(P2_U3208) );
  XNOR2_X1 U10187 ( .A(n8519), .B(n8520), .ZN(n8722) );
  XOR2_X1 U10188 ( .A(n8520), .B(n4590), .Z(n8522) );
  AOI222_X1 U10189 ( .A1(n8623), .A2(n8522), .B1(n8541), .B2(n8618), .C1(n8521), .C2(n8620), .ZN(n8718) );
  OAI21_X1 U10190 ( .B1(n8524), .B2(n8523), .A(n8718), .ZN(n8525) );
  NAND2_X1 U10191 ( .A1(n8525), .A2(n10103), .ZN(n8528) );
  AOI22_X1 U10192 ( .A1(n8526), .A2(n8626), .B1(n10105), .B2(
        P2_REG2_REG_24__SCAN_IN), .ZN(n8527) );
  OAI211_X1 U10193 ( .C1(n8722), .C2(n8630), .A(n8528), .B(n8527), .ZN(
        P2_U3209) );
  XNOR2_X1 U10194 ( .A(n8530), .B(n8529), .ZN(n8728) );
  XNOR2_X1 U10195 ( .A(n8532), .B(n8531), .ZN(n8535) );
  AOI222_X1 U10196 ( .A1(n8623), .A2(n8535), .B1(n8534), .B2(n8620), .C1(n8533), .C2(n8618), .ZN(n8723) );
  MUX2_X1 U10197 ( .A(n8536), .B(n8723), .S(n8610), .Z(n8539) );
  AOI22_X1 U10198 ( .A1(n8725), .A2(n8627), .B1(n8626), .B2(n8537), .ZN(n8538)
         );
  OAI211_X1 U10199 ( .C1(n8728), .C2(n8630), .A(n8539), .B(n8538), .ZN(
        P2_U3210) );
  XNOR2_X1 U10200 ( .A(n8540), .B(n8548), .ZN(n8542) );
  AOI222_X1 U10201 ( .A1(n8623), .A2(n8542), .B1(n6486), .B2(n8618), .C1(n8541), .C2(n8620), .ZN(n8656) );
  INV_X1 U10202 ( .A(n8543), .ZN(n8545) );
  OAI22_X1 U10203 ( .A1(n8545), .A2(n10097), .B1(n8610), .B2(n8544), .ZN(n8546) );
  AOI21_X1 U10204 ( .B1(n8547), .B2(n8627), .A(n8546), .ZN(n8551) );
  OR2_X1 U10205 ( .A1(n8549), .A2(n8548), .ZN(n8654) );
  NAND3_X1 U10206 ( .A1(n8654), .A2(n8562), .A3(n8653), .ZN(n8550) );
  OAI211_X1 U10207 ( .C1(n8656), .C2(n10105), .A(n8551), .B(n8550), .ZN(
        P2_U3211) );
  XNOR2_X1 U10208 ( .A(n8552), .B(n8556), .ZN(n8553) );
  OAI222_X1 U10209 ( .A1(n8598), .A2(n8555), .B1(n8596), .B2(n8554), .C1(n8593), .C2(n8553), .ZN(n8658) );
  INV_X1 U10210 ( .A(n8658), .ZN(n8564) );
  XNOR2_X1 U10211 ( .A(n8557), .B(n8556), .ZN(n8659) );
  AOI22_X1 U10212 ( .A1(n8558), .A2(n8626), .B1(n10105), .B2(
        P2_REG2_REG_21__SCAN_IN), .ZN(n8559) );
  OAI21_X1 U10213 ( .B1(n8734), .B2(n8560), .A(n8559), .ZN(n8561) );
  AOI21_X1 U10214 ( .B1(n8659), .B2(n8562), .A(n8561), .ZN(n8563) );
  OAI21_X1 U10215 ( .B1(n8564), .B2(n10105), .A(n8563), .ZN(P2_U3212) );
  XNOR2_X1 U10216 ( .A(n8565), .B(n8568), .ZN(n8739) );
  INV_X1 U10217 ( .A(n8566), .ZN(n8571) );
  OAI21_X1 U10218 ( .B1(n4559), .B2(n8568), .A(n8567), .ZN(n8570) );
  AOI222_X1 U10219 ( .A1(n8623), .A2(n8570), .B1(n6486), .B2(n8620), .C1(n8569), .C2(n8618), .ZN(n8735) );
  OAI21_X1 U10220 ( .B1(n8571), .B2(n10097), .A(n8735), .ZN(n8572) );
  NAND2_X1 U10221 ( .A1(n8572), .A2(n10103), .ZN(n8574) );
  AOI22_X1 U10222 ( .A1(n8736), .A2(n8627), .B1(P2_REG2_REG_20__SCAN_IN), .B2(
        n10105), .ZN(n8573) );
  OAI211_X1 U10223 ( .C1(n8739), .C2(n8630), .A(n8574), .B(n8573), .ZN(
        P2_U3213) );
  XOR2_X1 U10224 ( .A(n8575), .B(n8576), .Z(n8743) );
  NOR2_X1 U10225 ( .A1(n8577), .A2(n8576), .ZN(n8579) );
  AOI22_X1 U10226 ( .A1(n8580), .A2(n8620), .B1(n8618), .B2(n8607), .ZN(n8581)
         );
  NAND2_X1 U10227 ( .A1(n8582), .A2(n8581), .ZN(n8668) );
  INV_X1 U10228 ( .A(n8583), .ZN(n8584) );
  NOR2_X1 U10229 ( .A1(n8584), .A2(n10097), .ZN(n8585) );
  OAI21_X1 U10230 ( .B1(n8668), .B2(n8585), .A(n8610), .ZN(n8587) );
  AOI22_X1 U10231 ( .A1(n8666), .A2(n8627), .B1(P2_REG2_REG_19__SCAN_IN), .B2(
        n10105), .ZN(n8586) );
  OAI211_X1 U10232 ( .C1(n8743), .C2(n8630), .A(n8587), .B(n8586), .ZN(
        P2_U3214) );
  NAND2_X1 U10233 ( .A1(n8588), .A2(n8591), .ZN(n8589) );
  NAND2_X1 U10234 ( .A1(n8590), .A2(n8589), .ZN(n8747) );
  XOR2_X1 U10235 ( .A(n8592), .B(n8591), .Z(n8594) );
  OAI222_X1 U10236 ( .A1(n8598), .A2(n8597), .B1(n8596), .B2(n8595), .C1(n8594), .C2(n8593), .ZN(n8670) );
  NAND2_X1 U10237 ( .A1(n8670), .A2(n8610), .ZN(n8603) );
  INV_X1 U10238 ( .A(n8599), .ZN(n8600) );
  OAI22_X1 U10239 ( .A1(n8610), .A2(n10448), .B1(n8600), .B2(n10097), .ZN(
        n8601) );
  AOI21_X1 U10240 ( .B1(n8671), .B2(n8627), .A(n8601), .ZN(n8602) );
  OAI211_X1 U10241 ( .C1(n8747), .C2(n8630), .A(n8603), .B(n8602), .ZN(
        P2_U3215) );
  XOR2_X1 U10242 ( .A(n8604), .B(n8606), .Z(n8753) );
  XOR2_X1 U10243 ( .A(n8605), .B(n8606), .Z(n8609) );
  AOI222_X1 U10244 ( .A1(n8623), .A2(n8609), .B1(n8608), .B2(n8618), .C1(n8607), .C2(n8620), .ZN(n8748) );
  MUX2_X1 U10245 ( .A(n10384), .B(n8748), .S(n8610), .Z(n8613) );
  AOI22_X1 U10246 ( .A1(n8750), .A2(n8627), .B1(n8626), .B2(n8611), .ZN(n8612)
         );
  OAI211_X1 U10247 ( .C1(n8753), .C2(n8630), .A(n8613), .B(n8612), .ZN(
        P2_U3216) );
  XNOR2_X1 U10248 ( .A(n8615), .B(n8614), .ZN(n8761) );
  XNOR2_X1 U10249 ( .A(n8617), .B(n8616), .ZN(n8622) );
  AOI222_X1 U10250 ( .A1(n8623), .A2(n8622), .B1(n8621), .B2(n8620), .C1(n8619), .C2(n8618), .ZN(n8754) );
  MUX2_X1 U10251 ( .A(n8624), .B(n8754), .S(n10103), .Z(n8629) );
  AOI22_X1 U10252 ( .A1(n8757), .A2(n8627), .B1(n8626), .B2(n8625), .ZN(n8628)
         );
  OAI211_X1 U10253 ( .C1(n8761), .C2(n8630), .A(n8629), .B(n8628), .ZN(
        P2_U3217) );
  NAND2_X1 U10254 ( .A1(n8691), .A2(n8678), .ZN(n8631) );
  NAND2_X1 U10255 ( .A1(n8692), .A2(n10159), .ZN(n8632) );
  OAI211_X1 U10256 ( .C1(n10159), .C2(n7325), .A(n8631), .B(n8632), .ZN(
        P2_U3490) );
  NAND2_X1 U10257 ( .A1(n8695), .A2(n8678), .ZN(n8633) );
  OAI211_X1 U10258 ( .C1(n10159), .C2(n8634), .A(n8633), .B(n8632), .ZN(
        P2_U3489) );
  AOI22_X1 U10259 ( .A1(n8636), .A2(n10123), .B1(n10147), .B2(n8635), .ZN(
        n8637) );
  NAND2_X1 U10260 ( .A1(n8638), .A2(n8637), .ZN(n8699) );
  MUX2_X1 U10261 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n8699), .S(n10159), .Z(
        P2_U3487) );
  INV_X1 U10262 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n8639) );
  MUX2_X1 U10263 ( .A(n8639), .B(n8700), .S(n10159), .Z(n8641) );
  NAND2_X1 U10264 ( .A1(n8702), .A2(n8678), .ZN(n8640) );
  OAI211_X1 U10265 ( .C1(n8705), .C2(n8681), .A(n8641), .B(n8640), .ZN(
        P2_U3486) );
  INV_X1 U10266 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n8642) );
  MUX2_X1 U10267 ( .A(n8642), .B(n8706), .S(n10159), .Z(n8644) );
  NAND2_X1 U10268 ( .A1(n8708), .A2(n8678), .ZN(n8643) );
  OAI211_X1 U10269 ( .C1(n8681), .C2(n8711), .A(n8644), .B(n8643), .ZN(
        P2_U3485) );
  INV_X1 U10270 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n8645) );
  MUX2_X1 U10271 ( .A(n8645), .B(n8712), .S(n10159), .Z(n8647) );
  NAND2_X1 U10272 ( .A1(n8714), .A2(n8678), .ZN(n8646) );
  OAI211_X1 U10273 ( .C1(n8717), .C2(n8681), .A(n8647), .B(n8646), .ZN(
        P2_U3484) );
  INV_X1 U10274 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n8648) );
  MUX2_X1 U10275 ( .A(n8648), .B(n8718), .S(n10159), .Z(n8650) );
  NAND2_X1 U10276 ( .A1(n8719), .A2(n8678), .ZN(n8649) );
  OAI211_X1 U10277 ( .C1(n8681), .C2(n8722), .A(n8650), .B(n8649), .ZN(
        P2_U3483) );
  MUX2_X1 U10278 ( .A(n10337), .B(n8723), .S(n10159), .Z(n8652) );
  NAND2_X1 U10279 ( .A1(n8725), .A2(n8678), .ZN(n8651) );
  OAI211_X1 U10280 ( .C1(n8728), .C2(n8681), .A(n8652), .B(n8651), .ZN(
        P2_U3482) );
  NAND3_X1 U10281 ( .A1(n8654), .A2(n8653), .A3(n10123), .ZN(n8655) );
  OAI211_X1 U10282 ( .C1(n8657), .C2(n10119), .A(n8656), .B(n8655), .ZN(n8729)
         );
  MUX2_X1 U10283 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n8729), .S(n10159), .Z(
        P2_U3481) );
  INV_X1 U10284 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n8660) );
  AOI21_X1 U10285 ( .B1(n8659), .B2(n10123), .A(n8658), .ZN(n8730) );
  MUX2_X1 U10286 ( .A(n8660), .B(n8730), .S(n10159), .Z(n8661) );
  OAI21_X1 U10287 ( .B1(n8734), .B2(n8662), .A(n8661), .ZN(P2_U3480) );
  INV_X1 U10288 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n8663) );
  MUX2_X1 U10289 ( .A(n8663), .B(n8735), .S(n10159), .Z(n8665) );
  NAND2_X1 U10290 ( .A1(n8736), .A2(n8678), .ZN(n8664) );
  OAI211_X1 U10291 ( .C1(n8681), .C2(n8739), .A(n8665), .B(n8664), .ZN(
        P2_U3479) );
  INV_X1 U10292 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n10411) );
  AND2_X1 U10293 ( .A1(n8666), .A2(n10147), .ZN(n8667) );
  NOR2_X1 U10294 ( .A1(n8668), .A2(n8667), .ZN(n8740) );
  MUX2_X1 U10295 ( .A(n10411), .B(n8740), .S(n10159), .Z(n8669) );
  OAI21_X1 U10296 ( .B1(n8743), .B2(n8681), .A(n8669), .ZN(P2_U3478) );
  INV_X1 U10297 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8672) );
  AOI21_X1 U10298 ( .B1(n10147), .B2(n8671), .A(n8670), .ZN(n8744) );
  MUX2_X1 U10299 ( .A(n8672), .B(n8744), .S(n10159), .Z(n8673) );
  OAI21_X1 U10300 ( .B1(n8681), .B2(n8747), .A(n8673), .ZN(P2_U3477) );
  MUX2_X1 U10301 ( .A(n8674), .B(n8748), .S(n10159), .Z(n8676) );
  NAND2_X1 U10302 ( .A1(n8750), .A2(n8678), .ZN(n8675) );
  OAI211_X1 U10303 ( .C1(n8753), .C2(n8681), .A(n8676), .B(n8675), .ZN(
        P2_U3476) );
  MUX2_X1 U10304 ( .A(n8677), .B(n8754), .S(n10159), .Z(n8680) );
  NAND2_X1 U10305 ( .A1(n8757), .A2(n8678), .ZN(n8679) );
  OAI211_X1 U10306 ( .C1(n8681), .C2(n8761), .A(n8680), .B(n8679), .ZN(
        P2_U3475) );
  AOI22_X1 U10307 ( .A1(n8683), .A2(n10123), .B1(n10147), .B2(n8682), .ZN(
        n8684) );
  NAND2_X1 U10308 ( .A1(n8685), .A2(n8684), .ZN(n8762) );
  MUX2_X1 U10309 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n8762), .S(n10159), .Z(
        P2_U3474) );
  AOI22_X1 U10310 ( .A1(n8687), .A2(n10123), .B1(n10147), .B2(n8686), .ZN(
        n8688) );
  NAND2_X1 U10311 ( .A1(n8689), .A2(n8688), .ZN(n8763) );
  MUX2_X1 U10312 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n8763), .S(n10159), .Z(
        P2_U3470) );
  MUX2_X1 U10313 ( .A(n8690), .B(P2_REG1_REG_0__SCAN_IN), .S(n10157), .Z(
        P2_U3459) );
  INV_X1 U10314 ( .A(n8691), .ZN(n8694) );
  NAND2_X1 U10315 ( .A1(n10149), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n8693) );
  NAND2_X1 U10316 ( .A1(n8692), .A2(n10148), .ZN(n8696) );
  OAI211_X1 U10317 ( .C1(n8694), .C2(n8733), .A(n8693), .B(n8696), .ZN(
        P2_U3458) );
  INV_X1 U10318 ( .A(n8695), .ZN(n8698) );
  NAND2_X1 U10319 ( .A1(n10149), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n8697) );
  OAI211_X1 U10320 ( .C1(n8698), .C2(n8733), .A(n8697), .B(n8696), .ZN(
        P2_U3457) );
  MUX2_X1 U10321 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n8699), .S(n10148), .Z(
        P2_U3455) );
  INV_X1 U10322 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n8701) );
  MUX2_X1 U10323 ( .A(n8701), .B(n8700), .S(n10148), .Z(n8704) );
  NAND2_X1 U10324 ( .A1(n8702), .A2(n8756), .ZN(n8703) );
  OAI211_X1 U10325 ( .C1(n8705), .C2(n8760), .A(n8704), .B(n8703), .ZN(
        P2_U3454) );
  INV_X1 U10326 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n8707) );
  MUX2_X1 U10327 ( .A(n8707), .B(n8706), .S(n10148), .Z(n8710) );
  NAND2_X1 U10328 ( .A1(n8708), .A2(n8756), .ZN(n8709) );
  OAI211_X1 U10329 ( .C1(n8711), .C2(n8760), .A(n8710), .B(n8709), .ZN(
        P2_U3453) );
  INV_X1 U10330 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n8713) );
  MUX2_X1 U10331 ( .A(n8713), .B(n8712), .S(n10148), .Z(n8716) );
  NAND2_X1 U10332 ( .A1(n8714), .A2(n8756), .ZN(n8715) );
  OAI211_X1 U10333 ( .C1(n8717), .C2(n8760), .A(n8716), .B(n8715), .ZN(
        P2_U3452) );
  MUX2_X1 U10334 ( .A(n10408), .B(n8718), .S(n10148), .Z(n8721) );
  NAND2_X1 U10335 ( .A1(n8719), .A2(n8756), .ZN(n8720) );
  OAI211_X1 U10336 ( .C1(n8722), .C2(n8760), .A(n8721), .B(n8720), .ZN(
        P2_U3451) );
  INV_X1 U10337 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n8724) );
  MUX2_X1 U10338 ( .A(n8724), .B(n8723), .S(n10148), .Z(n8727) );
  NAND2_X1 U10339 ( .A1(n8725), .A2(n8756), .ZN(n8726) );
  OAI211_X1 U10340 ( .C1(n8728), .C2(n8760), .A(n8727), .B(n8726), .ZN(
        P2_U3450) );
  MUX2_X1 U10341 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n8729), .S(n10148), .Z(
        P2_U3449) );
  INV_X1 U10342 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n8731) );
  MUX2_X1 U10343 ( .A(n8731), .B(n8730), .S(n10148), .Z(n8732) );
  OAI21_X1 U10344 ( .B1(n8734), .B2(n8733), .A(n8732), .ZN(P2_U3448) );
  MUX2_X1 U10345 ( .A(n10432), .B(n8735), .S(n10148), .Z(n8738) );
  NAND2_X1 U10346 ( .A1(n8736), .A2(n8756), .ZN(n8737) );
  OAI211_X1 U10347 ( .C1(n8739), .C2(n8760), .A(n8738), .B(n8737), .ZN(
        P2_U3447) );
  INV_X1 U10348 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n8741) );
  MUX2_X1 U10349 ( .A(n8741), .B(n8740), .S(n10148), .Z(n8742) );
  OAI21_X1 U10350 ( .B1(n8743), .B2(n8760), .A(n8742), .ZN(P2_U3446) );
  INV_X1 U10351 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n8745) );
  MUX2_X1 U10352 ( .A(n8745), .B(n8744), .S(n10148), .Z(n8746) );
  OAI21_X1 U10353 ( .B1(n8747), .B2(n8760), .A(n8746), .ZN(P2_U3444) );
  MUX2_X1 U10354 ( .A(n8749), .B(n8748), .S(n10148), .Z(n8752) );
  NAND2_X1 U10355 ( .A1(n8750), .A2(n8756), .ZN(n8751) );
  OAI211_X1 U10356 ( .C1(n8753), .C2(n8760), .A(n8752), .B(n8751), .ZN(
        P2_U3441) );
  MUX2_X1 U10357 ( .A(n8755), .B(n8754), .S(n10148), .Z(n8759) );
  NAND2_X1 U10358 ( .A1(n8757), .A2(n8756), .ZN(n8758) );
  OAI211_X1 U10359 ( .C1(n8761), .C2(n8760), .A(n8759), .B(n8758), .ZN(
        P2_U3438) );
  MUX2_X1 U10360 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n8762), .S(n10148), .Z(
        P2_U3435) );
  MUX2_X1 U10361 ( .A(P2_REG0_REG_11__SCAN_IN), .B(n8763), .S(n10148), .Z(
        P2_U3423) );
  INV_X1 U10362 ( .A(n8961), .ZN(n9724) );
  NAND3_X1 U10363 ( .A1(n8764), .A2(P2_STATE_REG_SCAN_IN), .A3(
        P2_IR_REG_31__SCAN_IN), .ZN(n8766) );
  OAI22_X1 U10364 ( .A1(n8767), .A2(n8766), .B1(n6714), .B2(n8765), .ZN(n8768)
         );
  INV_X1 U10365 ( .A(n8768), .ZN(n8769) );
  OAI21_X1 U10366 ( .B1(n9724), .B2(n8787), .A(n8769), .ZN(P2_U3264) );
  OAI222_X1 U10367 ( .A1(n8773), .A2(P2_U3151), .B1(n8787), .B2(n8771), .C1(
        n8765), .C2(n8770), .ZN(P2_U3265) );
  NAND2_X1 U10368 ( .A1(n9728), .A2(n8774), .ZN(n8776) );
  OAI211_X1 U10369 ( .C1(n8765), .C2(n8777), .A(n8776), .B(n8775), .ZN(
        P2_U3267) );
  OAI222_X1 U10370 ( .A1(n8787), .A2(n8780), .B1(n8779), .B2(P2_U3151), .C1(
        n8778), .C2(n8765), .ZN(P2_U3268) );
  INV_X1 U10371 ( .A(n8781), .ZN(n9733) );
  OAI222_X1 U10372 ( .A1(n8787), .A2(n9733), .B1(P2_U3151), .B2(n8783), .C1(
        n8782), .C2(n8765), .ZN(P2_U3269) );
  INV_X1 U10373 ( .A(n8784), .ZN(n9737) );
  OAI222_X1 U10374 ( .A1(n8787), .A2(n9737), .B1(P2_U3151), .B2(n8786), .C1(
        n8785), .C2(n8765), .ZN(P2_U3270) );
  INV_X1 U10375 ( .A(n8788), .ZN(n8789) );
  MUX2_X1 U10376 ( .A(n8789), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  OAI21_X1 U10377 ( .B1(n8792), .B2(n8790), .A(n8791), .ZN(n8793) );
  NAND2_X1 U10378 ( .A1(n8793), .A2(n8942), .ZN(n8798) );
  INV_X1 U10379 ( .A(n8794), .ZN(n9580) );
  AOI22_X1 U10380 ( .A1(n9254), .A2(n9232), .B1(n8932), .B2(n9252), .ZN(n9566)
         );
  OAI22_X1 U10381 ( .A1(n8912), .A2(n9566), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8795), .ZN(n8796) );
  AOI21_X1 U10382 ( .B1(n9580), .B2(n8883), .A(n8796), .ZN(n8797) );
  OAI211_X1 U10383 ( .C1(n4638), .C2(n9766), .A(n8798), .B(n8797), .ZN(
        P1_U3215) );
  INV_X1 U10384 ( .A(n8799), .ZN(n8802) );
  NOR3_X1 U10385 ( .A1(n8909), .A2(n8904), .A3(n8800), .ZN(n8801) );
  OAI21_X1 U10386 ( .B1(n8802), .B2(n8801), .A(n8942), .ZN(n8807) );
  AOI22_X1 U10387 ( .A1(n8847), .A2(n8932), .B1(n9232), .B2(n9245), .ZN(n9431)
         );
  NOR2_X1 U10388 ( .A1(n9431), .A2(n8912), .ZN(n8805) );
  OAI22_X1 U10389 ( .A1(n9772), .A2(n9436), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8803), .ZN(n8804) );
  AOI211_X1 U10390 ( .C1(n9435), .C2(n8958), .A(n8805), .B(n8804), .ZN(n8806)
         );
  NAND2_X1 U10391 ( .A1(n8807), .A2(n8806), .ZN(P1_U3216) );
  OAI21_X1 U10392 ( .B1(n8809), .B2(n8808), .A(n7048), .ZN(n8810) );
  NAND2_X1 U10393 ( .A1(n8810), .A2(n8942), .ZN(n8815) );
  AOI22_X1 U10394 ( .A1(n9764), .A2(n8811), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        P1_U3086), .ZN(n8814) );
  AOI22_X1 U10395 ( .A1(n8958), .A2(n8812), .B1(n5240), .B2(n8883), .ZN(n8813)
         );
  NAND3_X1 U10396 ( .A1(n8815), .A2(n8814), .A3(n8813), .ZN(P1_U3218) );
  XNOR2_X1 U10397 ( .A(n8816), .B(n8817), .ZN(n8931) );
  NOR2_X1 U10398 ( .A1(n8931), .A2(n8930), .ZN(n8929) );
  AOI21_X1 U10399 ( .B1(n8817), .B2(n8816), .A(n8929), .ZN(n8821) );
  XNOR2_X1 U10400 ( .A(n8819), .B(n8818), .ZN(n8820) );
  XNOR2_X1 U10401 ( .A(n8821), .B(n8820), .ZN(n8826) );
  NOR2_X1 U10402 ( .A1(n9772), .A2(n9503), .ZN(n8824) );
  AOI22_X1 U10403 ( .A1(n9247), .A2(n8932), .B1(n9249), .B2(n9232), .ZN(n9495)
         );
  OAI21_X1 U10404 ( .B1(n8912), .B2(n9495), .A(n8822), .ZN(n8823) );
  AOI211_X1 U10405 ( .C1(n9502), .C2(n8958), .A(n8824), .B(n8823), .ZN(n8825)
         );
  OAI21_X1 U10406 ( .B1(n8826), .B2(n9758), .A(n8825), .ZN(P1_U3219) );
  XOR2_X1 U10407 ( .A(n8828), .B(n8827), .Z(n8834) );
  NAND2_X1 U10408 ( .A1(n9245), .A2(n8932), .ZN(n8830) );
  NAND2_X1 U10409 ( .A1(n9247), .A2(n9232), .ZN(n8829) );
  NAND2_X1 U10410 ( .A1(n8830), .A2(n8829), .ZN(n9464) );
  AOI22_X1 U10411 ( .A1(n9464), .A2(n9764), .B1(P1_REG3_REG_21__SCAN_IN), .B2(
        P1_U3086), .ZN(n8831) );
  OAI21_X1 U10412 ( .B1(n9471), .B2(n9772), .A(n8831), .ZN(n8832) );
  AOI21_X1 U10413 ( .B1(n9470), .B2(n8958), .A(n8832), .ZN(n8833) );
  OAI21_X1 U10414 ( .B1(n8834), .B2(n9758), .A(n8833), .ZN(P1_U3223) );
  XOR2_X1 U10415 ( .A(n8836), .B(n8835), .Z(n8844) );
  NAND2_X1 U10416 ( .A1(n9764), .A2(n8837), .ZN(n8839) );
  OAI211_X1 U10417 ( .C1(n9772), .C2(n8840), .A(n8839), .B(n8838), .ZN(n8841)
         );
  AOI21_X1 U10418 ( .B1(n8842), .B2(n8958), .A(n8841), .ZN(n8843) );
  OAI21_X1 U10419 ( .B1(n8844), .B2(n9758), .A(n8843), .ZN(P1_U3224) );
  AOI21_X1 U10420 ( .B1(n8846), .B2(n8845), .A(n8941), .ZN(n8851) );
  AOI22_X1 U10421 ( .A1(n9242), .A2(n8932), .B1(n9232), .B2(n8847), .ZN(n9401)
         );
  AOI22_X1 U10422 ( .A1(n8883), .A2(n9405), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3086), .ZN(n8848) );
  OAI21_X1 U10423 ( .B1(n9401), .B2(n8912), .A(n8848), .ZN(n8849) );
  AOI21_X1 U10424 ( .B1(n9404), .B2(n8958), .A(n8849), .ZN(n8850) );
  OAI21_X1 U10425 ( .B1(n8851), .B2(n9758), .A(n8850), .ZN(P1_U3225) );
  OAI21_X1 U10426 ( .B1(n8854), .B2(n8853), .A(n8852), .ZN(n8858) );
  XNOR2_X1 U10427 ( .A(n4511), .B(n8856), .ZN(n8953) );
  NOR2_X1 U10428 ( .A1(n8953), .A2(n8952), .ZN(n8951) );
  AOI21_X1 U10429 ( .B1(n8856), .B2(n4511), .A(n8951), .ZN(n8857) );
  XOR2_X1 U10430 ( .A(n8858), .B(n8857), .Z(n8864) );
  NAND2_X1 U10431 ( .A1(n9252), .A2(n9232), .ZN(n8860) );
  NAND2_X1 U10432 ( .A1(n9250), .A2(n8932), .ZN(n8859) );
  NAND2_X1 U10433 ( .A1(n8860), .A2(n8859), .ZN(n9551) );
  AOI22_X1 U10434 ( .A1(n9764), .A2(n9551), .B1(P1_REG3_REG_16__SCAN_IN), .B2(
        P1_U3086), .ZN(n8861) );
  OAI21_X1 U10435 ( .B1(n9556), .B2(n9772), .A(n8861), .ZN(n8862) );
  AOI21_X1 U10436 ( .B1(n9555), .B2(n8958), .A(n8862), .ZN(n8863) );
  OAI21_X1 U10437 ( .B1(n8864), .B2(n9758), .A(n8863), .ZN(P1_U3226) );
  NAND2_X1 U10438 ( .A1(n8867), .A2(n8866), .ZN(n8868) );
  XNOR2_X1 U10439 ( .A(n8865), .B(n8868), .ZN(n8876) );
  OR2_X1 U10440 ( .A1(n8869), .A2(n8944), .ZN(n8871) );
  NAND2_X1 U10441 ( .A1(n9249), .A2(n8932), .ZN(n8870) );
  NAND2_X1 U10442 ( .A1(n8871), .A2(n8870), .ZN(n9531) );
  NAND2_X1 U10443 ( .A1(n9764), .A2(n9531), .ZN(n8873) );
  OAI211_X1 U10444 ( .C1(n9772), .C2(n9538), .A(n8873), .B(n8872), .ZN(n8874)
         );
  AOI21_X1 U10445 ( .B1(n9537), .B2(n8958), .A(n8874), .ZN(n8875) );
  OAI21_X1 U10446 ( .B1(n8876), .B2(n9758), .A(n8875), .ZN(P1_U3228) );
  AND3_X1 U10447 ( .A1(n8799), .A2(n8878), .A3(n8877), .ZN(n8879) );
  OAI21_X1 U10448 ( .B1(n8880), .B2(n8879), .A(n8942), .ZN(n8885) );
  AOI22_X1 U10449 ( .A1(n9243), .A2(n8932), .B1(n9232), .B2(n9244), .ZN(n9414)
         );
  OAI22_X1 U10450 ( .A1(n9414), .A2(n8912), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8881), .ZN(n8882) );
  AOI21_X1 U10451 ( .B1(n9416), .B2(n8883), .A(n8882), .ZN(n8884) );
  OAI211_X1 U10452 ( .C1(n9682), .C2(n9766), .A(n8885), .B(n8884), .ZN(
        P1_U3229) );
  XNOR2_X1 U10453 ( .A(n8887), .B(n8886), .ZN(n8888) );
  XNOR2_X1 U10454 ( .A(n8889), .B(n8888), .ZN(n8894) );
  NOR2_X1 U10455 ( .A1(n9772), .A2(n9486), .ZN(n8892) );
  AOI22_X1 U10456 ( .A1(n9246), .A2(n8932), .B1(n9232), .B2(n9248), .ZN(n9481)
         );
  OAI22_X1 U10457 ( .A1(n8912), .A2(n9481), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8890), .ZN(n8891) );
  AOI211_X1 U10458 ( .C1(n9485), .C2(n8958), .A(n8892), .B(n8891), .ZN(n8893)
         );
  OAI21_X1 U10459 ( .B1(n8894), .B2(n9758), .A(n8893), .ZN(P1_U3233) );
  XOR2_X1 U10460 ( .A(n8895), .B(n8896), .Z(n8903) );
  AOI22_X1 U10461 ( .A1(n9764), .A2(n8897), .B1(P1_REG3_REG_13__SCAN_IN), .B2(
        P1_U3086), .ZN(n8898) );
  OAI21_X1 U10462 ( .B1(n8899), .B2(n9772), .A(n8898), .ZN(n8900) );
  AOI21_X1 U10463 ( .B1(n8901), .B2(n8958), .A(n8900), .ZN(n8902) );
  OAI21_X1 U10464 ( .B1(n8903), .B2(n9758), .A(n8902), .ZN(P1_U3234) );
  INV_X1 U10465 ( .A(n8904), .ZN(n8908) );
  OR2_X1 U10466 ( .A1(n8905), .A2(n8904), .ZN(n8906) );
  AOI22_X1 U10467 ( .A1(n8909), .A2(n8908), .B1(n8907), .B2(n8906), .ZN(n8916)
         );
  NOR2_X1 U10468 ( .A1(n9772), .A2(n9452), .ZN(n8914) );
  AND2_X1 U10469 ( .A1(n9246), .A2(n9232), .ZN(n8910) );
  AOI21_X1 U10470 ( .B1(n9244), .B2(n8932), .A(n8910), .ZN(n9446) );
  OAI22_X1 U10471 ( .A1(n9446), .A2(n8912), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8911), .ZN(n8913) );
  AOI211_X1 U10472 ( .C1(n9451), .C2(n8958), .A(n8914), .B(n8913), .ZN(n8915)
         );
  OAI21_X1 U10473 ( .B1(n8916), .B2(n9758), .A(n8915), .ZN(P1_U3235) );
  AOI21_X1 U10474 ( .B1(n8919), .B2(n8921), .A(n8918), .ZN(n8920) );
  AOI21_X1 U10475 ( .B1(n4512), .B2(n8921), .A(n8920), .ZN(n8928) );
  AOI22_X1 U10476 ( .A1(n9764), .A2(n8922), .B1(P1_REG3_REG_11__SCAN_IN), .B2(
        P1_U3086), .ZN(n8923) );
  OAI21_X1 U10477 ( .B1(n8924), .B2(n9772), .A(n8923), .ZN(n8925) );
  AOI21_X1 U10478 ( .B1(n4622), .B2(n8958), .A(n8925), .ZN(n8927) );
  OAI21_X1 U10479 ( .B1(n8928), .B2(n9758), .A(n8927), .ZN(P1_U3236) );
  AOI21_X1 U10480 ( .B1(n8931), .B2(n8930), .A(n8929), .ZN(n8938) );
  NAND2_X1 U10481 ( .A1(n9250), .A2(n9232), .ZN(n8934) );
  NAND2_X1 U10482 ( .A1(n9248), .A2(n8932), .ZN(n8933) );
  NAND2_X1 U10483 ( .A1(n8934), .A2(n8933), .ZN(n9514) );
  AOI22_X1 U10484 ( .A1(n9764), .A2(n9514), .B1(P1_REG3_REG_18__SCAN_IN), .B2(
        P1_U3086), .ZN(n8935) );
  OAI21_X1 U10485 ( .B1(n9520), .B2(n9772), .A(n8935), .ZN(n8936) );
  AOI21_X1 U10486 ( .B1(n9519), .B2(n8958), .A(n8936), .ZN(n8937) );
  OAI21_X1 U10487 ( .B1(n8938), .B2(n9758), .A(n8937), .ZN(P1_U3238) );
  OAI22_X1 U10488 ( .A1(n8947), .A2(n8946), .B1(n8945), .B2(n8944), .ZN(n9385)
         );
  OAI22_X1 U10489 ( .A1(n9388), .A2(n9772), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10348), .ZN(n8948) );
  AOI21_X1 U10490 ( .B1(n9385), .B2(n9764), .A(n8948), .ZN(n8949) );
  OAI211_X1 U10491 ( .C1(n9674), .C2(n9766), .A(n8950), .B(n8949), .ZN(
        P1_U3240) );
  AOI21_X1 U10492 ( .B1(n8953), .B2(n8952), .A(n8951), .ZN(n8960) );
  AOI22_X1 U10493 ( .A1(n9764), .A2(n8954), .B1(P1_REG3_REG_15__SCAN_IN), .B2(
        P1_U3086), .ZN(n8955) );
  OAI21_X1 U10494 ( .B1(n8956), .B2(n9772), .A(n8955), .ZN(n8957) );
  AOI21_X1 U10495 ( .B1(n9025), .B2(n8958), .A(n8957), .ZN(n8959) );
  OAI21_X1 U10496 ( .B1(n8960), .B2(n9758), .A(n8959), .ZN(P1_U3241) );
  INV_X1 U10497 ( .A(n9209), .ZN(n9220) );
  AOI21_X1 U10498 ( .B1(n9527), .B2(n9252), .A(n8983), .ZN(n9026) );
  INV_X1 U10499 ( .A(n9026), .ZN(n9041) );
  INV_X1 U10500 ( .A(n9034), .ZN(n8964) );
  OAI21_X1 U10501 ( .B1(n8964), .B2(n9022), .A(n9527), .ZN(n9040) );
  INV_X1 U10502 ( .A(n9263), .ZN(n8978) );
  INV_X1 U10503 ( .A(n8965), .ZN(n8971) );
  AND2_X1 U10504 ( .A1(n9152), .A2(n8983), .ZN(n8970) );
  NAND2_X1 U10505 ( .A1(n9155), .A2(n8966), .ZN(n8968) );
  NAND2_X1 U10506 ( .A1(n9152), .A2(n8981), .ZN(n8967) );
  MUX2_X1 U10507 ( .A(n8968), .B(n8967), .S(n9096), .Z(n8969) );
  INV_X1 U10508 ( .A(n9155), .ZN(n8972) );
  AOI21_X1 U10509 ( .B1(n8982), .B2(n8973), .A(n8972), .ZN(n8975) );
  INV_X1 U10510 ( .A(n8975), .ZN(n8977) );
  OAI21_X1 U10511 ( .B1(n8975), .B2(n9263), .A(n8974), .ZN(n8976) );
  OAI21_X1 U10512 ( .B1(n8978), .B2(n8977), .A(n8976), .ZN(n8979) );
  NAND2_X1 U10513 ( .A1(n8981), .A2(n8980), .ZN(n9158) );
  NOR2_X1 U10514 ( .A1(n8982), .A2(n9158), .ZN(n8984) );
  NAND2_X1 U10515 ( .A1(n8990), .A2(n8986), .ZN(n9162) );
  OAI22_X1 U10516 ( .A1(n8989), .A2(n8988), .B1(n9096), .B2(n8987), .ZN(n8998)
         );
  INV_X1 U10517 ( .A(n9163), .ZN(n9157) );
  OAI211_X1 U10518 ( .C1(n8991), .C2(n9157), .A(n8990), .B(n9113), .ZN(n8993)
         );
  NAND3_X1 U10519 ( .A1(n8993), .A2(n9096), .A3(n8992), .ZN(n8997) );
  NAND2_X1 U10520 ( .A1(n8995), .A2(n8994), .ZN(n8996) );
  AOI22_X1 U10521 ( .A1(n8998), .A2(n8997), .B1(n9096), .B2(n8996), .ZN(n9003)
         );
  NAND2_X1 U10522 ( .A1(n9004), .A2(n8999), .ZN(n9000) );
  MUX2_X1 U10523 ( .A(n9001), .B(n9000), .S(n9096), .Z(n9002) );
  NAND2_X1 U10524 ( .A1(n9009), .A2(n9004), .ZN(n9005) );
  NAND2_X1 U10525 ( .A1(n9013), .A2(n9010), .ZN(n9169) );
  AOI21_X1 U10526 ( .B1(n9005), .B2(n9170), .A(n9169), .ZN(n9007) );
  NAND2_X1 U10527 ( .A1(n9014), .A2(n9006), .ZN(n9173) );
  OAI21_X1 U10528 ( .B1(n9007), .B2(n9173), .A(n9172), .ZN(n9019) );
  NAND2_X1 U10529 ( .A1(n9009), .A2(n9008), .ZN(n9011) );
  NAND2_X1 U10530 ( .A1(n9011), .A2(n9010), .ZN(n9017) );
  INV_X1 U10531 ( .A(n9170), .ZN(n9012) );
  NOR2_X1 U10532 ( .A1(n9173), .A2(n9012), .ZN(n9016) );
  NAND2_X1 U10533 ( .A1(n9172), .A2(n9013), .ZN(n9104) );
  MUX2_X1 U10534 ( .A(n9019), .B(n9018), .S(n9096), .Z(n9032) );
  NAND2_X1 U10535 ( .A1(n9020), .A2(n9031), .ZN(n9148) );
  AOI21_X1 U10536 ( .B1(n9032), .B2(n9567), .A(n9148), .ZN(n9024) );
  NAND2_X1 U10537 ( .A1(n9022), .A2(n9021), .ZN(n9175) );
  NAND2_X1 U10538 ( .A1(n9029), .A2(n9028), .ZN(n9030) );
  NAND2_X1 U10539 ( .A1(n9030), .A2(n9096), .ZN(n9039) );
  NAND2_X1 U10540 ( .A1(n9032), .A2(n9031), .ZN(n9037) );
  NAND2_X1 U10541 ( .A1(n9034), .A2(n9033), .ZN(n9178) );
  AOI211_X1 U10542 ( .C1(n9037), .C2(n9036), .A(n9035), .B(n9178), .ZN(n9038)
         );
  NAND2_X1 U10543 ( .A1(n9047), .A2(n9042), .ZN(n9180) );
  NAND2_X1 U10544 ( .A1(n9053), .A2(n9046), .ZN(n9183) );
  INV_X1 U10545 ( .A(n9054), .ZN(n9043) );
  OAI211_X1 U10546 ( .C1(n9044), .C2(n9183), .A(n9043), .B(n9182), .ZN(n9052)
         );
  INV_X1 U10547 ( .A(n9045), .ZN(n9050) );
  AND2_X1 U10548 ( .A1(n9046), .A2(n9511), .ZN(n9125) );
  INV_X1 U10549 ( .A(n9047), .ZN(n9049) );
  INV_X1 U10550 ( .A(n9182), .ZN(n9048) );
  AOI211_X1 U10551 ( .C1(n9050), .C2(n9125), .A(n9049), .B(n9048), .ZN(n9051)
         );
  AOI21_X1 U10552 ( .B1(n9460), .B2(n9053), .A(n8983), .ZN(n9058) );
  INV_X1 U10553 ( .A(n9061), .ZN(n9055) );
  NOR2_X1 U10554 ( .A1(n9055), .A2(n9054), .ZN(n9056) );
  MUX2_X1 U10555 ( .A(n9146), .B(n9056), .S(n9096), .Z(n9057) );
  MUX2_X1 U10556 ( .A(n9061), .B(n9060), .S(n9096), .Z(n9062) );
  NAND2_X1 U10557 ( .A1(n9065), .A2(n9063), .ZN(n9185) );
  AND2_X1 U10558 ( .A1(n9064), .A2(n9185), .ZN(n9067) );
  NAND2_X1 U10559 ( .A1(n9064), .A2(n9427), .ZN(n9066) );
  AND2_X1 U10560 ( .A1(n9066), .A2(n9065), .ZN(n9140) );
  MUX2_X1 U10561 ( .A(n9067), .B(n9140), .S(n9096), .Z(n9068) );
  MUX2_X1 U10562 ( .A(n9188), .B(n9142), .S(n9096), .Z(n9069) );
  INV_X1 U10563 ( .A(n9078), .ZN(n9071) );
  INV_X1 U10564 ( .A(n9145), .ZN(n9070) );
  AOI211_X1 U10565 ( .C1(n9077), .C2(n9189), .A(n9071), .B(n9070), .ZN(n9074)
         );
  INV_X1 U10566 ( .A(n9195), .ZN(n9075) );
  NAND2_X1 U10567 ( .A1(n9073), .A2(n9072), .ZN(n9192) );
  NOR4_X1 U10568 ( .A1(n9074), .A2(n9075), .A3(n8983), .A4(n9192), .ZN(n9088)
         );
  INV_X1 U10569 ( .A(n9189), .ZN(n9076) );
  NAND2_X1 U10570 ( .A1(n9081), .A2(n9078), .ZN(n9198) );
  NAND2_X1 U10571 ( .A1(n9080), .A2(n8983), .ZN(n9084) );
  NOR3_X1 U10572 ( .A1(n9079), .A2(n9198), .A3(n9084), .ZN(n9087) );
  NOR2_X1 U10573 ( .A1(n9080), .A2(n8983), .ZN(n9086) );
  INV_X1 U10574 ( .A(n9081), .ZN(n9082) );
  AOI21_X1 U10575 ( .B1(n9096), .B2(n9082), .A(n9192), .ZN(n9083) );
  AOI21_X1 U10576 ( .B1(n9192), .B2(n9084), .A(n9083), .ZN(n9085) );
  MUX2_X1 U10577 ( .A(n9200), .B(n9202), .S(n9096), .Z(n9089) );
  NAND2_X1 U10578 ( .A1(n9091), .A2(n5295), .ZN(n9094) );
  OR2_X1 U10579 ( .A1(n5234), .A2(n9092), .ZN(n9093) );
  INV_X1 U10580 ( .A(n9335), .ZN(n9095) );
  NOR2_X1 U10581 ( .A1(n9095), .A2(n9101), .ZN(n9213) );
  NOR3_X1 U10582 ( .A1(n9235), .A2(n9236), .A3(n9097), .ZN(n9098) );
  OAI21_X1 U10583 ( .B1(n9100), .B2(n9099), .A(n9150), .ZN(n9139) );
  NOR2_X1 U10584 ( .A1(n9230), .A2(n9223), .ZN(n9227) );
  INV_X1 U10585 ( .A(n9235), .ZN(n9138) );
  OR2_X1 U10586 ( .A1(n9343), .A2(n9101), .ZN(n9204) );
  NAND2_X1 U10587 ( .A1(n9343), .A2(n9101), .ZN(n9206) );
  INV_X1 U10588 ( .A(n9384), .ZN(n9133) );
  XNOR2_X1 U10589 ( .A(n9485), .B(n9102), .ZN(n9484) );
  INV_X1 U10590 ( .A(n9180), .ZN(n9126) );
  INV_X1 U10591 ( .A(n9173), .ZN(n9119) );
  INV_X1 U10592 ( .A(n9104), .ZN(n9118) );
  NOR3_X1 U10593 ( .A1(n9106), .A2(n9105), .A3(n9150), .ZN(n9112) );
  NOR2_X1 U10594 ( .A1(n9108), .A2(n9107), .ZN(n9110) );
  AND4_X1 U10595 ( .A1(n9112), .A2(n9111), .A3(n9110), .A4(n9109), .ZN(n9114)
         );
  NAND4_X1 U10596 ( .A1(n9166), .A2(n9164), .A3(n9114), .A4(n9113), .ZN(n9116)
         );
  NOR2_X1 U10597 ( .A1(n9116), .A2(n9115), .ZN(n9117) );
  NAND4_X1 U10598 ( .A1(n4742), .A2(n9119), .A3(n9118), .A4(n9117), .ZN(n9120)
         );
  OR3_X1 U10599 ( .A1(n9121), .A2(n9120), .A3(n9573), .ZN(n9122) );
  NOR2_X1 U10600 ( .A1(n9123), .A2(n9122), .ZN(n9124) );
  NAND4_X1 U10601 ( .A1(n9497), .A2(n9126), .A3(n9125), .A4(n9124), .ZN(n9127)
         );
  NOR2_X1 U10602 ( .A1(n9484), .A2(n9127), .ZN(n9130) );
  XNOR2_X1 U10603 ( .A(n9470), .B(n9128), .ZN(n9461) );
  NOR2_X1 U10604 ( .A1(n9448), .A2(n9461), .ZN(n9129) );
  AND4_X1 U10605 ( .A1(n9412), .A2(n9131), .A3(n9130), .A4(n9129), .ZN(n9132)
         );
  AND4_X1 U10606 ( .A1(n9367), .A2(n9133), .A3(n9399), .A4(n9132), .ZN(n9134)
         );
  NAND4_X1 U10607 ( .A1(n9204), .A2(n9206), .A3(n9135), .A4(n9134), .ZN(n9137)
         );
  NAND4_X1 U10608 ( .A1(n9139), .A2(n9227), .A3(n9138), .A4(n9225), .ZN(n9239)
         );
  INV_X1 U10609 ( .A(n9140), .ZN(n9141) );
  NAND2_X1 U10610 ( .A1(n9142), .A2(n9141), .ZN(n9143) );
  NAND2_X1 U10611 ( .A1(n9143), .A2(n9188), .ZN(n9144) );
  NAND2_X1 U10612 ( .A1(n9145), .A2(n9144), .ZN(n9191) );
  INV_X1 U10613 ( .A(n9146), .ZN(n9147) );
  NOR2_X1 U10614 ( .A1(n9191), .A2(n9147), .ZN(n9212) );
  INV_X1 U10615 ( .A(n9148), .ZN(n9177) );
  INV_X1 U10616 ( .A(n9149), .ZN(n9151) );
  NAND4_X1 U10617 ( .A1(n9153), .A2(n9152), .A3(n9151), .A4(n9150), .ZN(n9154)
         );
  NAND3_X1 U10618 ( .A1(n9156), .A2(n9155), .A3(n9154), .ZN(n9161) );
  NOR2_X1 U10619 ( .A1(n9158), .A2(n9157), .ZN(n9160) );
  AOI21_X1 U10620 ( .B1(n9161), .B2(n9160), .A(n9159), .ZN(n9168) );
  INV_X1 U10621 ( .A(n9164), .ZN(n9167) );
  NAND3_X1 U10622 ( .A1(n9164), .A2(n9163), .A3(n9162), .ZN(n9165) );
  OAI211_X1 U10623 ( .C1(n9168), .C2(n9167), .A(n9166), .B(n9165), .ZN(n9171)
         );
  AOI21_X1 U10624 ( .B1(n9171), .B2(n9170), .A(n9169), .ZN(n9174) );
  OAI211_X1 U10625 ( .C1(n9174), .C2(n9173), .A(n9567), .B(n9172), .ZN(n9176)
         );
  AOI21_X1 U10626 ( .B1(n9177), .B2(n9176), .A(n9175), .ZN(n9179) );
  OAI21_X1 U10627 ( .B1(n9179), .B2(n9178), .A(n9527), .ZN(n9181) );
  AOI21_X1 U10628 ( .B1(n9511), .B2(n9181), .A(n9180), .ZN(n9184) );
  OAI21_X1 U10629 ( .B1(n9184), .B2(n9183), .A(n9182), .ZN(n9196) );
  INV_X1 U10630 ( .A(n9198), .ZN(n9194) );
  INV_X1 U10631 ( .A(n9185), .ZN(n9187) );
  AND3_X1 U10632 ( .A1(n9188), .A2(n9187), .A3(n9186), .ZN(n9190) );
  OAI21_X1 U10633 ( .B1(n9191), .B2(n9190), .A(n9189), .ZN(n9193) );
  AOI21_X1 U10634 ( .B1(n9194), .B2(n9193), .A(n9192), .ZN(n9199) );
  NAND3_X1 U10635 ( .A1(n9200), .A2(n9199), .A3(n9195), .ZN(n9211) );
  AOI21_X1 U10636 ( .B1(n9212), .B2(n9196), .A(n9211), .ZN(n9208) );
  AOI21_X1 U10637 ( .B1(n9199), .B2(n9198), .A(n9197), .ZN(n9203) );
  INV_X1 U10638 ( .A(n9200), .ZN(n9201) );
  AOI21_X1 U10639 ( .B1(n9203), .B2(n9202), .A(n9201), .ZN(n9215) );
  INV_X1 U10640 ( .A(n9215), .ZN(n9205) );
  NAND2_X1 U10641 ( .A1(n9205), .A2(n9204), .ZN(n9207) );
  OAI21_X1 U10642 ( .B1(n9208), .B2(n9207), .A(n9206), .ZN(n9210) );
  AOI21_X1 U10643 ( .B1(n9210), .B2(n4949), .A(n9209), .ZN(n9231) );
  INV_X1 U10644 ( .A(n9213), .ZN(n9217) );
  AOI21_X1 U10645 ( .B1(n9212), .B2(n9479), .A(n9211), .ZN(n9214) );
  OAI22_X1 U10646 ( .A1(n9215), .A2(n9214), .B1(n4948), .B2(n9213), .ZN(n9216)
         );
  OAI21_X1 U10647 ( .B1(n9217), .B2(n9343), .A(n9216), .ZN(n9221) );
  AOI211_X1 U10648 ( .C1(n9221), .C2(n9220), .A(n9219), .B(n9218), .ZN(n9222)
         );
  INV_X1 U10649 ( .A(n9222), .ZN(n9226) );
  INV_X1 U10650 ( .A(n9223), .ZN(n9224) );
  NAND3_X1 U10651 ( .A1(n9226), .A2(n9225), .A3(n9224), .ZN(n9229) );
  AOI211_X1 U10652 ( .C1(n9231), .C2(n9233), .A(n9227), .B(n9235), .ZN(n9228)
         );
  OAI211_X1 U10653 ( .C1(n9231), .C2(n9230), .A(n9229), .B(n9228), .ZN(n9238)
         );
  NAND4_X1 U10654 ( .A1(n9717), .A2(n9774), .A3(n9233), .A4(n9232), .ZN(n9234)
         );
  OAI211_X1 U10655 ( .C1(n9236), .C2(n9235), .A(n9234), .B(P1_B_REG_SCAN_IN), 
        .ZN(n9237) );
  NAND4_X1 U10656 ( .A1(n9240), .A2(n9239), .A3(n9238), .A4(n9237), .ZN(
        P1_U3242) );
  MUX2_X1 U10657 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9241), .S(P1_U3973), .Z(
        P1_U3581) );
  MUX2_X1 U10658 ( .A(n9242), .B(P1_DATAO_REG_26__SCAN_IN), .S(n9265), .Z(
        P1_U3580) );
  MUX2_X1 U10659 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9243), .S(P1_U3973), .Z(
        P1_U3579) );
  MUX2_X1 U10660 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9244), .S(P1_U3973), .Z(
        P1_U3577) );
  MUX2_X1 U10661 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9245), .S(P1_U3973), .Z(
        P1_U3576) );
  MUX2_X1 U10662 ( .A(n9246), .B(P1_DATAO_REG_21__SCAN_IN), .S(n9265), .Z(
        P1_U3575) );
  MUX2_X1 U10663 ( .A(n9247), .B(P1_DATAO_REG_20__SCAN_IN), .S(n9265), .Z(
        P1_U3574) );
  MUX2_X1 U10664 ( .A(n9248), .B(P1_DATAO_REG_19__SCAN_IN), .S(n9265), .Z(
        P1_U3573) );
  MUX2_X1 U10665 ( .A(n9249), .B(P1_DATAO_REG_18__SCAN_IN), .S(n9265), .Z(
        P1_U3572) );
  MUX2_X1 U10666 ( .A(n9250), .B(P1_DATAO_REG_17__SCAN_IN), .S(n9265), .Z(
        P1_U3571) );
  MUX2_X1 U10667 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9251), .S(P1_U3973), .Z(
        P1_U3570) );
  MUX2_X1 U10668 ( .A(n9252), .B(P1_DATAO_REG_15__SCAN_IN), .S(n9265), .Z(
        P1_U3569) );
  MUX2_X1 U10669 ( .A(n9253), .B(P1_DATAO_REG_14__SCAN_IN), .S(n9265), .Z(
        P1_U3568) );
  MUX2_X1 U10670 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9254), .S(P1_U3973), .Z(
        P1_U3567) );
  MUX2_X1 U10671 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n9255), .S(P1_U3973), .Z(
        P1_U3566) );
  MUX2_X1 U10672 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n9256), .S(P1_U3973), .Z(
        P1_U3565) );
  MUX2_X1 U10673 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n9257), .S(P1_U3973), .Z(
        P1_U3564) );
  MUX2_X1 U10674 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n9258), .S(P1_U3973), .Z(
        P1_U3563) );
  MUX2_X1 U10675 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n9259), .S(P1_U3973), .Z(
        P1_U3562) );
  MUX2_X1 U10676 ( .A(n9260), .B(P1_DATAO_REG_7__SCAN_IN), .S(n9265), .Z(
        P1_U3561) );
  MUX2_X1 U10677 ( .A(n9261), .B(P1_DATAO_REG_6__SCAN_IN), .S(n9265), .Z(
        P1_U3560) );
  MUX2_X1 U10678 ( .A(n9262), .B(P1_DATAO_REG_5__SCAN_IN), .S(n9265), .Z(
        P1_U3559) );
  MUX2_X1 U10679 ( .A(n9263), .B(P1_DATAO_REG_4__SCAN_IN), .S(n9265), .Z(
        P1_U3558) );
  MUX2_X1 U10680 ( .A(n9264), .B(P1_DATAO_REG_3__SCAN_IN), .S(n9265), .Z(
        P1_U3557) );
  MUX2_X1 U10681 ( .A(n5852), .B(P1_DATAO_REG_2__SCAN_IN), .S(n9265), .Z(
        P1_U3556) );
  MUX2_X1 U10682 ( .A(n5840), .B(P1_DATAO_REG_1__SCAN_IN), .S(n9265), .Z(
        P1_U3555) );
  INV_X1 U10683 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n9267) );
  NAND2_X1 U10684 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_U3086), .ZN(n9266) );
  OAI21_X1 U10685 ( .B1(n9853), .B2(n9267), .A(n9266), .ZN(n9268) );
  AOI21_X1 U10686 ( .B1(n9269), .B2(n10568), .A(n9268), .ZN(n9278) );
  OAI211_X1 U10687 ( .C1(n9272), .C2(n9271), .A(n10563), .B(n9270), .ZN(n9277)
         );
  OAI211_X1 U10688 ( .C1(n9275), .C2(n9274), .A(n10559), .B(n9273), .ZN(n9276)
         );
  NAND3_X1 U10689 ( .A1(n9278), .A2(n9277), .A3(n9276), .ZN(P1_U3246) );
  INV_X1 U10690 ( .A(n9279), .ZN(n9283) );
  INV_X1 U10691 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n9281) );
  NAND2_X1 U10692 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n9280) );
  OAI21_X1 U10693 ( .B1(n9853), .B2(n9281), .A(n9280), .ZN(n9282) );
  AOI21_X1 U10694 ( .B1(n9283), .B2(n10568), .A(n9282), .ZN(n9292) );
  OAI211_X1 U10695 ( .C1(n9286), .C2(n9285), .A(n10563), .B(n9284), .ZN(n9291)
         );
  OAI211_X1 U10696 ( .C1(n9289), .C2(n9288), .A(n10559), .B(n9287), .ZN(n9290)
         );
  NAND3_X1 U10697 ( .A1(n9292), .A2(n9291), .A3(n9290), .ZN(P1_U3248) );
  INV_X1 U10698 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n9294) );
  NAND2_X1 U10699 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_U3086), .ZN(n9293) );
  OAI21_X1 U10700 ( .B1(n9853), .B2(n9294), .A(n9293), .ZN(n9295) );
  AOI21_X1 U10701 ( .B1(n9296), .B2(n10568), .A(n9295), .ZN(n9305) );
  OAI211_X1 U10702 ( .C1(n9299), .C2(n9298), .A(n10563), .B(n9297), .ZN(n9304)
         );
  OAI211_X1 U10703 ( .C1(n9302), .C2(n9301), .A(n10559), .B(n9300), .ZN(n9303)
         );
  NAND3_X1 U10704 ( .A1(n9305), .A2(n9304), .A3(n9303), .ZN(P1_U3249) );
  INV_X1 U10705 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n9307) );
  NAND2_X1 U10706 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3086), .ZN(n9306) );
  OAI21_X1 U10707 ( .B1(n9853), .B2(n9307), .A(n9306), .ZN(n9308) );
  AOI21_X1 U10708 ( .B1(n9309), .B2(n10568), .A(n9308), .ZN(n9318) );
  OAI211_X1 U10709 ( .C1(n9312), .C2(n9311), .A(n10563), .B(n9310), .ZN(n9317)
         );
  OAI211_X1 U10710 ( .C1(n9315), .C2(n9314), .A(n10559), .B(n9313), .ZN(n9316)
         );
  NAND3_X1 U10711 ( .A1(n9318), .A2(n9317), .A3(n9316), .ZN(P1_U3250) );
  INV_X1 U10712 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n10454) );
  OAI21_X1 U10713 ( .B1(n9853), .B2(n10454), .A(n9319), .ZN(n9320) );
  AOI21_X1 U10714 ( .B1(n9321), .B2(n10568), .A(n9320), .ZN(n9330) );
  OAI211_X1 U10715 ( .C1(n9324), .C2(n9323), .A(n10559), .B(n9322), .ZN(n9329)
         );
  OAI211_X1 U10716 ( .C1(n9327), .C2(n9326), .A(n10563), .B(n9325), .ZN(n9328)
         );
  NAND3_X1 U10717 ( .A1(n9330), .A2(n9329), .A3(n9328), .ZN(P1_U3251) );
  NOR2_X1 U10718 ( .A1(n9339), .A2(n9343), .ZN(n9331) );
  XNOR2_X1 U10719 ( .A(n9665), .B(n9331), .ZN(n9332) );
  INV_X1 U10720 ( .A(n9333), .ZN(n9334) );
  AND2_X1 U10721 ( .A1(n9335), .A2(n9334), .ZN(n9585) );
  INV_X1 U10722 ( .A(n9585), .ZN(n9589) );
  OR2_X1 U10723 ( .A1(n9857), .A2(n9589), .ZN(n9340) );
  NAND2_X1 U10724 ( .A1(n9857), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n9336) );
  OAI211_X1 U10725 ( .C1(n9665), .C2(n9873), .A(n9340), .B(n9336), .ZN(n9337)
         );
  AOI21_X1 U10726 ( .B1(n9586), .B2(n9877), .A(n9337), .ZN(n9338) );
  INV_X1 U10727 ( .A(n9338), .ZN(P1_U3263) );
  OAI21_X1 U10728 ( .B1(n9561), .B2(n9341), .A(n9340), .ZN(n9342) );
  AOI21_X1 U10729 ( .B1(n9343), .B2(n9866), .A(n9342), .ZN(n9344) );
  OAI21_X1 U10730 ( .B1(n9590), .B2(n9859), .A(n9344), .ZN(P1_U3264) );
  NAND2_X1 U10731 ( .A1(n9345), .A2(n9535), .ZN(n9355) );
  OAI22_X1 U10732 ( .A1(n9347), .A2(n9869), .B1(n9561), .B2(n9346), .ZN(n9348)
         );
  AOI21_X1 U10733 ( .B1(n9349), .B2(n9866), .A(n9348), .ZN(n9354) );
  NAND2_X1 U10734 ( .A1(n9350), .A2(n9561), .ZN(n9353) );
  NAND2_X1 U10735 ( .A1(n9351), .A2(n9877), .ZN(n9352) );
  NAND4_X1 U10736 ( .A1(n9355), .A2(n9354), .A3(n9353), .A4(n9352), .ZN(
        P1_U3356) );
  NAND2_X1 U10737 ( .A1(n9356), .A2(n9535), .ZN(n9364) );
  INV_X1 U10738 ( .A(n9357), .ZN(n9362) );
  AOI22_X1 U10739 ( .A1(n9358), .A2(n9855), .B1(P1_REG2_REG_28__SCAN_IN), .B2(
        n9857), .ZN(n9359) );
  OAI21_X1 U10740 ( .B1(n9360), .B2(n9873), .A(n9359), .ZN(n9361) );
  AOI21_X1 U10741 ( .B1(n9362), .B2(n9877), .A(n9361), .ZN(n9363) );
  OAI211_X1 U10742 ( .C1(n9857), .C2(n9365), .A(n9364), .B(n9363), .ZN(
        P1_U3265) );
  XNOR2_X1 U10743 ( .A(n9366), .B(n9367), .ZN(n9593) );
  INV_X1 U10744 ( .A(n9593), .ZN(n9381) );
  XNOR2_X1 U10745 ( .A(n9368), .B(n9367), .ZN(n9369) );
  NAND2_X1 U10746 ( .A1(n9369), .A2(n9549), .ZN(n9372) );
  INV_X1 U10747 ( .A(n9370), .ZN(n9371) );
  NAND2_X1 U10748 ( .A1(n9372), .A2(n9371), .ZN(n9591) );
  INV_X1 U10749 ( .A(n9373), .ZN(n9374) );
  AOI211_X1 U10750 ( .C1(n9375), .C2(n9390), .A(n9578), .B(n9374), .ZN(n9592)
         );
  NAND2_X1 U10751 ( .A1(n9592), .A2(n9877), .ZN(n9378) );
  AOI22_X1 U10752 ( .A1(n9376), .A2(n9855), .B1(P1_REG2_REG_27__SCAN_IN), .B2(
        n9857), .ZN(n9377) );
  OAI211_X1 U10753 ( .C1(n4654), .C2(n9873), .A(n9378), .B(n9377), .ZN(n9379)
         );
  AOI21_X1 U10754 ( .B1(n9561), .B2(n9591), .A(n9379), .ZN(n9380) );
  OAI21_X1 U10755 ( .B1(n9381), .B2(n9861), .A(n9380), .ZN(P1_U3266) );
  XOR2_X1 U10756 ( .A(n9384), .B(n9382), .Z(n9598) );
  NAND2_X1 U10757 ( .A1(n9598), .A2(n9535), .ZN(n9396) );
  AOI22_X1 U10758 ( .A1(n9392), .A2(n9866), .B1(n9857), .B2(
        P1_REG2_REG_26__SCAN_IN), .ZN(n9395) );
  XOR2_X1 U10759 ( .A(n9384), .B(n9383), .Z(n9387) );
  INV_X1 U10760 ( .A(n9385), .ZN(n9386) );
  OAI21_X1 U10761 ( .B1(n9387), .B2(n9571), .A(n9386), .ZN(n9596) );
  NOR2_X1 U10762 ( .A1(n9388), .A2(n9869), .ZN(n9389) );
  OAI21_X1 U10763 ( .B1(n9596), .B2(n9389), .A(n9561), .ZN(n9394) );
  INV_X1 U10764 ( .A(n9390), .ZN(n9391) );
  AOI211_X1 U10765 ( .C1(n9392), .C2(n4657), .A(n9578), .B(n9391), .ZN(n9597)
         );
  NAND2_X1 U10766 ( .A1(n9597), .A2(n9877), .ZN(n9393) );
  NAND4_X1 U10767 ( .A1(n9396), .A2(n9395), .A3(n9394), .A4(n9393), .ZN(
        P1_U3267) );
  XOR2_X1 U10768 ( .A(n9397), .B(n9399), .Z(n9603) );
  INV_X1 U10769 ( .A(n9603), .ZN(n9410) );
  OAI211_X1 U10770 ( .C1(n9400), .C2(n9399), .A(n9398), .B(n9549), .ZN(n9402)
         );
  NAND2_X1 U10771 ( .A1(n9402), .A2(n9401), .ZN(n9601) );
  INV_X1 U10772 ( .A(n9404), .ZN(n9678) );
  AOI211_X1 U10773 ( .C1(n9404), .C2(n9417), .A(n9578), .B(n9403), .ZN(n9602)
         );
  NAND2_X1 U10774 ( .A1(n9602), .A2(n9877), .ZN(n9407) );
  AOI22_X1 U10775 ( .A1(n9405), .A2(n9855), .B1(n9857), .B2(
        P1_REG2_REG_25__SCAN_IN), .ZN(n9406) );
  OAI211_X1 U10776 ( .C1(n9678), .C2(n9873), .A(n9407), .B(n9406), .ZN(n9408)
         );
  AOI21_X1 U10777 ( .B1(n9561), .B2(n9601), .A(n9408), .ZN(n9409) );
  OAI21_X1 U10778 ( .B1(n9410), .B2(n9861), .A(n9409), .ZN(P1_U3268) );
  XNOR2_X1 U10779 ( .A(n9411), .B(n9412), .ZN(n9608) );
  XNOR2_X1 U10780 ( .A(n9413), .B(n9412), .ZN(n9415) );
  OAI21_X1 U10781 ( .B1(n9415), .B2(n9571), .A(n9414), .ZN(n9606) );
  AOI21_X1 U10782 ( .B1(n9416), .B2(n9855), .A(n9606), .ZN(n9423) );
  AOI22_X1 U10783 ( .A1(n9420), .A2(n9866), .B1(n9857), .B2(
        P1_REG2_REG_24__SCAN_IN), .ZN(n9422) );
  INV_X1 U10784 ( .A(n9433), .ZN(n9419) );
  INV_X1 U10785 ( .A(n9417), .ZN(n9418) );
  AOI211_X1 U10786 ( .C1(n9420), .C2(n9419), .A(n9578), .B(n9418), .ZN(n9607)
         );
  NAND2_X1 U10787 ( .A1(n9607), .A2(n9877), .ZN(n9421) );
  OAI211_X1 U10788 ( .C1(n9423), .C2(n9857), .A(n9422), .B(n9421), .ZN(n9424)
         );
  AOI21_X1 U10789 ( .B1(n9608), .B2(n9535), .A(n9424), .ZN(n9425) );
  INV_X1 U10790 ( .A(n9425), .ZN(P1_U3269) );
  XNOR2_X1 U10791 ( .A(n9426), .B(n9428), .ZN(n9612) );
  INV_X1 U10792 ( .A(n9612), .ZN(n9442) );
  NAND2_X1 U10793 ( .A1(n9445), .A2(n9427), .ZN(n9429) );
  XNOR2_X1 U10794 ( .A(n9429), .B(n9428), .ZN(n9430) );
  NAND2_X1 U10795 ( .A1(n9430), .A2(n9549), .ZN(n9432) );
  NAND2_X1 U10796 ( .A1(n9432), .A2(n9431), .ZN(n9610) );
  INV_X1 U10797 ( .A(n9450), .ZN(n9434) );
  AOI211_X1 U10798 ( .C1(n9435), .C2(n9434), .A(n9578), .B(n9433), .ZN(n9611)
         );
  NAND2_X1 U10799 ( .A1(n9611), .A2(n9877), .ZN(n9439) );
  INV_X1 U10800 ( .A(n9436), .ZN(n9437) );
  AOI22_X1 U10801 ( .A1(n9857), .A2(P1_REG2_REG_23__SCAN_IN), .B1(n9437), .B2(
        n9855), .ZN(n9438) );
  OAI211_X1 U10802 ( .C1(n9686), .C2(n9873), .A(n9439), .B(n9438), .ZN(n9440)
         );
  AOI21_X1 U10803 ( .B1(n9561), .B2(n9610), .A(n9440), .ZN(n9441) );
  OAI21_X1 U10804 ( .B1(n9442), .B2(n9861), .A(n9441), .ZN(P1_U3270) );
  NAND2_X1 U10805 ( .A1(n9443), .A2(n9448), .ZN(n9444) );
  NAND3_X1 U10806 ( .A1(n9445), .A2(n9549), .A3(n9444), .ZN(n9447) );
  NAND2_X1 U10807 ( .A1(n9447), .A2(n9446), .ZN(n9615) );
  INV_X1 U10808 ( .A(n9615), .ZN(n9458) );
  XOR2_X1 U10809 ( .A(n9449), .B(n9448), .Z(n9617) );
  NAND2_X1 U10810 ( .A1(n9617), .A2(n9535), .ZN(n9457) );
  AOI211_X1 U10811 ( .C1(n9451), .C2(n9468), .A(n9578), .B(n9450), .ZN(n9616)
         );
  NOR2_X1 U10812 ( .A1(n4646), .A2(n9873), .ZN(n9455) );
  INV_X1 U10813 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n9453) );
  OAI22_X1 U10814 ( .A1(n9561), .A2(n9453), .B1(n9452), .B2(n9869), .ZN(n9454)
         );
  AOI211_X1 U10815 ( .C1(n9616), .C2(n9877), .A(n9455), .B(n9454), .ZN(n9456)
         );
  OAI211_X1 U10816 ( .C1(n9857), .C2(n9458), .A(n9457), .B(n9456), .ZN(
        P1_U3271) );
  XNOR2_X1 U10817 ( .A(n9459), .B(n9461), .ZN(n9622) );
  INV_X1 U10818 ( .A(n9622), .ZN(n9477) );
  OAI21_X1 U10819 ( .B1(n9479), .B2(n9484), .A(n9460), .ZN(n9462) );
  XNOR2_X1 U10820 ( .A(n9462), .B(n9461), .ZN(n9463) );
  NAND2_X1 U10821 ( .A1(n9463), .A2(n9549), .ZN(n9466) );
  INV_X1 U10822 ( .A(n9464), .ZN(n9465) );
  NAND2_X1 U10823 ( .A1(n9466), .A2(n9465), .ZN(n9620) );
  INV_X1 U10824 ( .A(n9468), .ZN(n9469) );
  AOI211_X1 U10825 ( .C1(n9470), .C2(n4650), .A(n9578), .B(n9469), .ZN(n9621)
         );
  NAND2_X1 U10826 ( .A1(n9621), .A2(n9877), .ZN(n9474) );
  INV_X1 U10827 ( .A(n9471), .ZN(n9472) );
  AOI22_X1 U10828 ( .A1(n9857), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n9472), .B2(
        n9855), .ZN(n9473) );
  OAI211_X1 U10829 ( .C1(n5791), .C2(n9873), .A(n9474), .B(n9473), .ZN(n9475)
         );
  AOI21_X1 U10830 ( .B1(n9561), .B2(n9620), .A(n9475), .ZN(n9476) );
  OAI21_X1 U10831 ( .B1(n9477), .B2(n9861), .A(n9476), .ZN(P1_U3272) );
  INV_X1 U10832 ( .A(n9484), .ZN(n9478) );
  XNOR2_X1 U10833 ( .A(n9479), .B(n9478), .ZN(n9480) );
  NAND2_X1 U10834 ( .A1(n9480), .A2(n9549), .ZN(n9482) );
  NAND2_X1 U10835 ( .A1(n9482), .A2(n9481), .ZN(n9625) );
  INV_X1 U10836 ( .A(n9625), .ZN(n9492) );
  XOR2_X1 U10837 ( .A(n9484), .B(n9483), .Z(n9627) );
  NAND2_X1 U10838 ( .A1(n9627), .A2(n9535), .ZN(n9491) );
  AOI211_X1 U10839 ( .C1(n9485), .C2(n9499), .A(n9578), .B(n9467), .ZN(n9626)
         );
  INV_X1 U10840 ( .A(n9485), .ZN(n9695) );
  NOR2_X1 U10841 ( .A1(n9695), .A2(n9873), .ZN(n9489) );
  OAI22_X1 U10842 ( .A1(n9561), .A2(n9487), .B1(n9486), .B2(n9869), .ZN(n9488)
         );
  AOI211_X1 U10843 ( .C1(n9626), .C2(n9877), .A(n9489), .B(n9488), .ZN(n9490)
         );
  OAI211_X1 U10844 ( .C1(n9857), .C2(n9492), .A(n9491), .B(n9490), .ZN(
        P1_U3273) );
  XNOR2_X1 U10845 ( .A(n9493), .B(n9497), .ZN(n9494) );
  NAND2_X1 U10846 ( .A1(n9494), .A2(n9549), .ZN(n9496) );
  NAND2_X1 U10847 ( .A1(n9496), .A2(n9495), .ZN(n9629) );
  INV_X1 U10848 ( .A(n9629), .ZN(n9509) );
  XOR2_X1 U10849 ( .A(n9498), .B(n9497), .Z(n9631) );
  NAND2_X1 U10850 ( .A1(n9631), .A2(n9535), .ZN(n9508) );
  INV_X1 U10851 ( .A(n9517), .ZN(n9501) );
  INV_X1 U10852 ( .A(n9499), .ZN(n9500) );
  AOI211_X1 U10853 ( .C1(n9502), .C2(n9501), .A(n9578), .B(n9500), .ZN(n9630)
         );
  NOR2_X1 U10854 ( .A1(n9699), .A2(n9873), .ZN(n9506) );
  OAI22_X1 U10855 ( .A1(n9561), .A2(n9504), .B1(n9503), .B2(n9869), .ZN(n9505)
         );
  AOI211_X1 U10856 ( .C1(n9630), .C2(n9877), .A(n9506), .B(n9505), .ZN(n9507)
         );
  OAI211_X1 U10857 ( .C1(n9857), .C2(n9509), .A(n9508), .B(n9507), .ZN(
        P1_U3274) );
  XOR2_X1 U10858 ( .A(n9513), .B(n9510), .Z(n9636) );
  INV_X1 U10859 ( .A(n9636), .ZN(n9526) );
  NAND2_X1 U10860 ( .A1(n9528), .A2(n9511), .ZN(n9512) );
  XOR2_X1 U10861 ( .A(n9513), .B(n9512), .Z(n9516) );
  INV_X1 U10862 ( .A(n9514), .ZN(n9515) );
  OAI21_X1 U10863 ( .B1(n9516), .B2(n9571), .A(n9515), .ZN(n9634) );
  INV_X1 U10864 ( .A(n9536), .ZN(n9518) );
  AOI211_X1 U10865 ( .C1(n9519), .C2(n9518), .A(n9578), .B(n9517), .ZN(n9635)
         );
  NAND2_X1 U10866 ( .A1(n9635), .A2(n9877), .ZN(n9523) );
  INV_X1 U10867 ( .A(n9520), .ZN(n9521) );
  AOI22_X1 U10868 ( .A1(n9857), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9521), .B2(
        n9855), .ZN(n9522) );
  OAI211_X1 U10869 ( .C1(n9703), .C2(n9873), .A(n9523), .B(n9522), .ZN(n9524)
         );
  AOI21_X1 U10870 ( .B1(n9634), .B2(n9561), .A(n9524), .ZN(n9525) );
  OAI21_X1 U10871 ( .B1(n9526), .B2(n9861), .A(n9525), .ZN(P1_U3275) );
  NAND2_X1 U10872 ( .A1(n9546), .A2(n9527), .ZN(n9530) );
  INV_X1 U10873 ( .A(n9528), .ZN(n9529) );
  AOI211_X1 U10874 ( .C1(n9533), .C2(n9530), .A(n9571), .B(n9529), .ZN(n9532)
         );
  OR2_X1 U10875 ( .A1(n9532), .A2(n9531), .ZN(n9639) );
  INV_X1 U10876 ( .A(n9639), .ZN(n9544) );
  XOR2_X1 U10877 ( .A(n9534), .B(n9533), .Z(n9641) );
  NAND2_X1 U10878 ( .A1(n9641), .A2(n9535), .ZN(n9543) );
  AOI211_X1 U10879 ( .C1(n9537), .C2(n9554), .A(n9578), .B(n9536), .ZN(n9640)
         );
  INV_X1 U10880 ( .A(n9537), .ZN(n9707) );
  NOR2_X1 U10881 ( .A1(n9707), .A2(n9873), .ZN(n9541) );
  OAI22_X1 U10882 ( .A1(n9561), .A2(n9539), .B1(n9538), .B2(n9869), .ZN(n9540)
         );
  AOI211_X1 U10883 ( .C1(n9640), .C2(n9877), .A(n9541), .B(n9540), .ZN(n9542)
         );
  OAI211_X1 U10884 ( .C1(n9857), .C2(n9544), .A(n9543), .B(n9542), .ZN(
        P1_U3276) );
  XNOR2_X1 U10885 ( .A(n9545), .B(n9548), .ZN(n9645) );
  INV_X1 U10886 ( .A(n9645), .ZN(n9563) );
  OAI21_X1 U10887 ( .B1(n9548), .B2(n9547), .A(n9546), .ZN(n9550) );
  NAND2_X1 U10888 ( .A1(n9550), .A2(n9549), .ZN(n9553) );
  INV_X1 U10889 ( .A(n9551), .ZN(n9552) );
  NAND2_X1 U10890 ( .A1(n9553), .A2(n9552), .ZN(n9643) );
  AOI211_X1 U10891 ( .C1(n9555), .C2(n4534), .A(n9578), .B(n4640), .ZN(n9644)
         );
  NAND2_X1 U10892 ( .A1(n9644), .A2(n9877), .ZN(n9559) );
  INV_X1 U10893 ( .A(n9556), .ZN(n9557) );
  AOI22_X1 U10894 ( .A1(n9857), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n9557), .B2(
        n9855), .ZN(n9558) );
  OAI211_X1 U10895 ( .C1(n4639), .C2(n9873), .A(n9559), .B(n9558), .ZN(n9560)
         );
  AOI21_X1 U10896 ( .B1(n9643), .B2(n9561), .A(n9560), .ZN(n9562) );
  OAI21_X1 U10897 ( .B1(n9563), .B2(n9861), .A(n9562), .ZN(P1_U3277) );
  INV_X1 U10898 ( .A(n9564), .ZN(n9576) );
  XNOR2_X1 U10899 ( .A(n9565), .B(n9573), .ZN(n9653) );
  INV_X1 U10900 ( .A(n9566), .ZN(n9575) );
  NAND2_X1 U10901 ( .A1(n9568), .A2(n9567), .ZN(n9572) );
  INV_X1 U10902 ( .A(n9569), .ZN(n9570) );
  AOI211_X1 U10903 ( .C1(n9573), .C2(n9572), .A(n9571), .B(n9570), .ZN(n9574)
         );
  AOI211_X1 U10904 ( .C1(n9576), .C2(n9653), .A(n9575), .B(n9574), .ZN(n9658)
         );
  AOI211_X1 U10905 ( .C1(n9655), .C2(n9579), .A(n9578), .B(n9577), .ZN(n9654)
         );
  NAND2_X1 U10906 ( .A1(n9654), .A2(n9877), .ZN(n9582) );
  AOI22_X1 U10907 ( .A1(n9857), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n9580), .B2(
        n9855), .ZN(n9581) );
  OAI211_X1 U10908 ( .C1(n4638), .C2(n9873), .A(n9582), .B(n9581), .ZN(n9583)
         );
  AOI21_X1 U10909 ( .B1(n9653), .B2(n9878), .A(n9583), .ZN(n9584) );
  OAI21_X1 U10910 ( .B1(n9658), .B2(n9857), .A(n9584), .ZN(P1_U3279) );
  MUX2_X1 U10911 ( .A(n9587), .B(n9662), .S(n9918), .Z(n9588) );
  OAI21_X1 U10912 ( .B1(n9665), .B2(n9652), .A(n9588), .ZN(P1_U3553) );
  AOI211_X1 U10913 ( .C1(n9593), .C2(n9908), .A(n9592), .B(n9591), .ZN(n9668)
         );
  MUX2_X1 U10914 ( .A(n9594), .B(n9668), .S(n9918), .Z(n9595) );
  OAI21_X1 U10915 ( .B1(n4654), .B2(n9652), .A(n9595), .ZN(P1_U3549) );
  AOI211_X1 U10916 ( .C1(n9598), .C2(n9908), .A(n9597), .B(n9596), .ZN(n9671)
         );
  MUX2_X1 U10917 ( .A(n9599), .B(n9671), .S(n9918), .Z(n9600) );
  OAI21_X1 U10918 ( .B1(n9674), .B2(n9652), .A(n9600), .ZN(P1_U3548) );
  AOI211_X1 U10919 ( .C1(n9603), .C2(n9908), .A(n9602), .B(n9601), .ZN(n9675)
         );
  MUX2_X1 U10920 ( .A(n9604), .B(n9675), .S(n9918), .Z(n9605) );
  OAI21_X1 U10921 ( .B1(n9678), .B2(n9652), .A(n9605), .ZN(P1_U3547) );
  AOI211_X1 U10922 ( .C1(n9608), .C2(n9908), .A(n9607), .B(n9606), .ZN(n9679)
         );
  MUX2_X1 U10923 ( .A(n10416), .B(n9679), .S(n9918), .Z(n9609) );
  OAI21_X1 U10924 ( .B1(n9682), .B2(n9652), .A(n9609), .ZN(P1_U3546) );
  AOI211_X1 U10925 ( .C1(n9612), .C2(n9908), .A(n9611), .B(n9610), .ZN(n9683)
         );
  MUX2_X1 U10926 ( .A(n9613), .B(n9683), .S(n9918), .Z(n9614) );
  OAI21_X1 U10927 ( .B1(n9686), .B2(n9652), .A(n9614), .ZN(P1_U3545) );
  INV_X1 U10928 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n9618) );
  AOI211_X1 U10929 ( .C1(n9617), .C2(n9908), .A(n9616), .B(n9615), .ZN(n9687)
         );
  MUX2_X1 U10930 ( .A(n9618), .B(n9687), .S(n9918), .Z(n9619) );
  OAI21_X1 U10931 ( .B1(n4646), .B2(n9652), .A(n9619), .ZN(P1_U3544) );
  INV_X1 U10932 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n9623) );
  AOI211_X1 U10933 ( .C1(n9622), .C2(n9908), .A(n9621), .B(n9620), .ZN(n9690)
         );
  MUX2_X1 U10934 ( .A(n9623), .B(n9690), .S(n9918), .Z(n9624) );
  OAI21_X1 U10935 ( .B1(n5791), .B2(n9652), .A(n9624), .ZN(P1_U3543) );
  AOI211_X1 U10936 ( .C1(n9627), .C2(n9908), .A(n9626), .B(n9625), .ZN(n9692)
         );
  MUX2_X1 U10937 ( .A(n10371), .B(n9692), .S(n9918), .Z(n9628) );
  OAI21_X1 U10938 ( .B1(n9695), .B2(n9652), .A(n9628), .ZN(P1_U3542) );
  AOI211_X1 U10939 ( .C1(n9631), .C2(n9908), .A(n9630), .B(n9629), .ZN(n9696)
         );
  MUX2_X1 U10940 ( .A(n9632), .B(n9696), .S(n9918), .Z(n9633) );
  OAI21_X1 U10941 ( .B1(n9699), .B2(n9652), .A(n9633), .ZN(P1_U3541) );
  AOI211_X1 U10942 ( .C1(n9636), .C2(n9908), .A(n9635), .B(n9634), .ZN(n9700)
         );
  MUX2_X1 U10943 ( .A(n9637), .B(n9700), .S(n9918), .Z(n9638) );
  OAI21_X1 U10944 ( .B1(n9703), .B2(n9652), .A(n9638), .ZN(P1_U3540) );
  AOI211_X1 U10945 ( .C1(n9641), .C2(n9908), .A(n9640), .B(n9639), .ZN(n9704)
         );
  MUX2_X1 U10946 ( .A(n10324), .B(n9704), .S(n9918), .Z(n9642) );
  OAI21_X1 U10947 ( .B1(n9707), .B2(n9652), .A(n9642), .ZN(P1_U3539) );
  AOI211_X1 U10948 ( .C1(n9645), .C2(n9908), .A(n9644), .B(n9643), .ZN(n9708)
         );
  MUX2_X1 U10949 ( .A(n10443), .B(n9708), .S(n9918), .Z(n9646) );
  OAI21_X1 U10950 ( .B1(n4639), .B2(n9652), .A(n9646), .ZN(P1_U3538) );
  NAND2_X1 U10951 ( .A1(n9648), .A2(n9647), .ZN(n9649) );
  AOI21_X1 U10952 ( .B1(n9650), .B2(n9908), .A(n9649), .ZN(n9710) );
  MUX2_X1 U10953 ( .A(n9816), .B(n9710), .S(n9918), .Z(n9651) );
  OAI21_X1 U10954 ( .B1(n9714), .B2(n9652), .A(n9651), .ZN(P1_U3537) );
  INV_X1 U10955 ( .A(n9653), .ZN(n9660) );
  AOI21_X1 U10956 ( .B1(n9656), .B2(n9655), .A(n9654), .ZN(n9657) );
  OAI211_X1 U10957 ( .C1(n9660), .C2(n9659), .A(n9658), .B(n9657), .ZN(n9715)
         );
  MUX2_X1 U10958 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n9715), .S(n9918), .Z(
        P1_U3536) );
  MUX2_X1 U10959 ( .A(n9661), .B(P1_REG1_REG_0__SCAN_IN), .S(n9916), .Z(
        P1_U3522) );
  INV_X1 U10960 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n9663) );
  MUX2_X1 U10961 ( .A(n9663), .B(n9662), .S(n9911), .Z(n9664) );
  OAI21_X1 U10962 ( .B1(n9665), .B2(n9713), .A(n9664), .ZN(P1_U3521) );
  MUX2_X1 U10963 ( .A(n9666), .B(n5760), .S(n9910), .Z(n9667) );
  OAI21_X1 U10964 ( .B1(n4948), .B2(n9713), .A(n9667), .ZN(P1_U3520) );
  INV_X1 U10965 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n9669) );
  MUX2_X1 U10966 ( .A(n9669), .B(n9668), .S(n9911), .Z(n9670) );
  OAI21_X1 U10967 ( .B1(n4654), .B2(n9713), .A(n9670), .ZN(P1_U3517) );
  INV_X1 U10968 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n9672) );
  MUX2_X1 U10969 ( .A(n9672), .B(n9671), .S(n9911), .Z(n9673) );
  OAI21_X1 U10970 ( .B1(n9674), .B2(n9713), .A(n9673), .ZN(P1_U3516) );
  INV_X1 U10971 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n9676) );
  MUX2_X1 U10972 ( .A(n9676), .B(n9675), .S(n9911), .Z(n9677) );
  OAI21_X1 U10973 ( .B1(n9678), .B2(n9713), .A(n9677), .ZN(P1_U3515) );
  INV_X1 U10974 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n9680) );
  MUX2_X1 U10975 ( .A(n9680), .B(n9679), .S(n9911), .Z(n9681) );
  OAI21_X1 U10976 ( .B1(n9682), .B2(n9713), .A(n9681), .ZN(P1_U3514) );
  INV_X1 U10977 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n9684) );
  MUX2_X1 U10978 ( .A(n9684), .B(n9683), .S(n9911), .Z(n9685) );
  OAI21_X1 U10979 ( .B1(n9686), .B2(n9713), .A(n9685), .ZN(P1_U3513) );
  INV_X1 U10980 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n9688) );
  MUX2_X1 U10981 ( .A(n9688), .B(n9687), .S(n9911), .Z(n9689) );
  OAI21_X1 U10982 ( .B1(n4646), .B2(n9713), .A(n9689), .ZN(P1_U3512) );
  MUX2_X1 U10983 ( .A(n10446), .B(n9690), .S(n9911), .Z(n9691) );
  OAI21_X1 U10984 ( .B1(n5791), .B2(n9713), .A(n9691), .ZN(P1_U3511) );
  INV_X1 U10985 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n9693) );
  MUX2_X1 U10986 ( .A(n9693), .B(n9692), .S(n9911), .Z(n9694) );
  OAI21_X1 U10987 ( .B1(n9695), .B2(n9713), .A(n9694), .ZN(P1_U3510) );
  INV_X1 U10988 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n9697) );
  MUX2_X1 U10989 ( .A(n9697), .B(n9696), .S(n9911), .Z(n9698) );
  OAI21_X1 U10990 ( .B1(n9699), .B2(n9713), .A(n9698), .ZN(P1_U3509) );
  MUX2_X1 U10991 ( .A(n9701), .B(n9700), .S(n9911), .Z(n9702) );
  OAI21_X1 U10992 ( .B1(n9703), .B2(n9713), .A(n9702), .ZN(P1_U3507) );
  INV_X1 U10993 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n9705) );
  MUX2_X1 U10994 ( .A(n9705), .B(n9704), .S(n9911), .Z(n9706) );
  OAI21_X1 U10995 ( .B1(n9707), .B2(n9713), .A(n9706), .ZN(P1_U3504) );
  MUX2_X1 U10996 ( .A(n10430), .B(n9708), .S(n9911), .Z(n9709) );
  OAI21_X1 U10997 ( .B1(n4639), .B2(n9713), .A(n9709), .ZN(P1_U3501) );
  INV_X1 U10998 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n9711) );
  MUX2_X1 U10999 ( .A(n9711), .B(n9710), .S(n9911), .Z(n9712) );
  OAI21_X1 U11000 ( .B1(n9714), .B2(n9713), .A(n9712), .ZN(P1_U3498) );
  MUX2_X1 U11001 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n9715), .S(n9911), .Z(
        P1_U3495) );
  AND2_X1 U11002 ( .A1(n9717), .A2(n9716), .ZN(n9883) );
  MUX2_X1 U11003 ( .A(P1_D_REG_1__SCAN_IN), .B(n9718), .S(n9883), .Z(P1_U3440)
         );
  MUX2_X1 U11004 ( .A(P1_D_REG_0__SCAN_IN), .B(n9719), .S(n9883), .Z(P1_U3439)
         );
  NOR4_X1 U11005 ( .A1(n9720), .A2(P1_IR_REG_30__SCAN_IN), .A3(n5276), .A4(
        P1_U3086), .ZN(n9721) );
  AOI21_X1 U11006 ( .B1(n9722), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9721), .ZN(
        n9723) );
  OAI21_X1 U11007 ( .B1(n9724), .B2(n9730), .A(n9723), .ZN(P1_U3324) );
  OAI222_X1 U11008 ( .A1(n9735), .A2(n9727), .B1(P1_U3086), .B2(n9726), .C1(
        n9730), .C2(n9725), .ZN(P1_U3326) );
  INV_X1 U11009 ( .A(n9728), .ZN(n9729) );
  OAI222_X1 U11010 ( .A1(n9735), .A2(n9731), .B1(n9730), .B2(n9729), .C1(n5757), .C2(P1_U3086), .ZN(P1_U3327) );
  OAI222_X1 U11011 ( .A1(P1_U3086), .A2(n9734), .B1(n9738), .B2(n9733), .C1(
        n9732), .C2(n9735), .ZN(P1_U3329) );
  OAI222_X1 U11012 ( .A1(P1_U3086), .A2(n9739), .B1(n9738), .B2(n9737), .C1(
        n9736), .C2(n9735), .ZN(P1_U3330) );
  MUX2_X1 U11013 ( .A(n9740), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  INV_X1 U11014 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n9755) );
  NAND2_X1 U11015 ( .A1(n9742), .A2(n9741), .ZN(n9743) );
  NAND2_X1 U11016 ( .A1(n9743), .A2(n10563), .ZN(n9751) );
  AND2_X1 U11017 ( .A1(n9745), .A2(n9744), .ZN(n9746) );
  OR3_X1 U11018 ( .A1(n9747), .A2(n9832), .A3(n9746), .ZN(n9750) );
  NAND2_X1 U11019 ( .A1(n10568), .A2(n9748), .ZN(n9749) );
  OAI211_X1 U11020 ( .C1(n9752), .C2(n9751), .A(n9750), .B(n9749), .ZN(n9753)
         );
  INV_X1 U11021 ( .A(n9753), .ZN(n9754) );
  NAND2_X1 U11022 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n9761) );
  OAI211_X1 U11023 ( .C1(n9853), .C2(n9755), .A(n9754), .B(n9761), .ZN(
        P1_U3253) );
  NAND2_X1 U11024 ( .A1(n9756), .A2(n9757), .ZN(n9759) );
  AOI21_X1 U11025 ( .B1(n9760), .B2(n9759), .A(n9758), .ZN(n9769) );
  INV_X1 U11026 ( .A(n9761), .ZN(n9762) );
  AOI21_X1 U11027 ( .B1(n9764), .B2(n9763), .A(n9762), .ZN(n9765) );
  OAI21_X1 U11028 ( .B1(n9767), .B2(n9766), .A(n9765), .ZN(n9768) );
  NOR2_X1 U11029 ( .A1(n9769), .A2(n9768), .ZN(n9770) );
  OAI21_X1 U11030 ( .B1(n9772), .B2(n9771), .A(n9770), .ZN(P1_U3217) );
  XNOR2_X1 U11031 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  OAI21_X1 U11032 ( .B1(n9774), .B2(P1_REG1_REG_0__SCAN_IN), .A(n9773), .ZN(
        n9775) );
  XOR2_X1 U11033 ( .A(P1_IR_REG_0__SCAN_IN), .B(n9775), .Z(n9778) );
  AOI22_X1 U11034 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(n10566), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n9776) );
  OAI21_X1 U11035 ( .B1(n9778), .B2(n9777), .A(n9776), .ZN(P1_U3243) );
  INV_X1 U11036 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n9790) );
  AOI211_X1 U11037 ( .C1(n9781), .C2(n9780), .A(n9779), .B(n9832), .ZN(n9786)
         );
  AOI211_X1 U11038 ( .C1(n9784), .C2(n9783), .A(n9782), .B(n9845), .ZN(n9785)
         );
  AOI211_X1 U11039 ( .C1(n10568), .C2(n9787), .A(n9786), .B(n9785), .ZN(n9789)
         );
  NAND2_X1 U11040 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n9788) );
  OAI211_X1 U11041 ( .C1(n9853), .C2(n9790), .A(n9789), .B(n9788), .ZN(
        P1_U3254) );
  INV_X1 U11042 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n9802) );
  AOI211_X1 U11043 ( .C1(n9793), .C2(n9792), .A(n9845), .B(n9791), .ZN(n9798)
         );
  AOI211_X1 U11044 ( .C1(n9796), .C2(n9795), .A(n9832), .B(n9794), .ZN(n9797)
         );
  AOI211_X1 U11045 ( .C1(n10568), .C2(n9799), .A(n9798), .B(n9797), .ZN(n9801)
         );
  NAND2_X1 U11046 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3086), .ZN(n9800) );
  OAI211_X1 U11047 ( .C1(n9853), .C2(n9802), .A(n9801), .B(n9800), .ZN(
        P1_U3256) );
  INV_X1 U11048 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n9814) );
  AOI211_X1 U11049 ( .C1(n9805), .C2(n9804), .A(n9803), .B(n9832), .ZN(n9810)
         );
  AOI211_X1 U11050 ( .C1(n9808), .C2(n9807), .A(n9845), .B(n9806), .ZN(n9809)
         );
  AOI211_X1 U11051 ( .C1(n10568), .C2(n9811), .A(n9810), .B(n9809), .ZN(n9813)
         );
  NAND2_X1 U11052 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n9812) );
  OAI211_X1 U11053 ( .C1(n9853), .C2(n9814), .A(n9813), .B(n9812), .ZN(
        P1_U3257) );
  AOI211_X1 U11054 ( .C1(n9817), .C2(n9816), .A(n9815), .B(n9845), .ZN(n9821)
         );
  AOI211_X1 U11055 ( .C1(n9819), .C2(n7871), .A(n9818), .B(n9832), .ZN(n9820)
         );
  AOI211_X1 U11056 ( .C1(n10568), .C2(n9822), .A(n9821), .B(n9820), .ZN(n9825)
         );
  NAND2_X1 U11057 ( .A1(P1_REG3_REG_15__SCAN_IN), .A2(P1_U3086), .ZN(n9824) );
  OAI211_X1 U11058 ( .C1(n9853), .C2(n9826), .A(n9825), .B(n9824), .ZN(
        P1_U3258) );
  XOR2_X1 U11059 ( .A(n9828), .B(n9827), .Z(n9829) );
  NOR2_X1 U11060 ( .A1(n9829), .A2(n9845), .ZN(n9836) );
  INV_X1 U11061 ( .A(n9830), .ZN(n9831) );
  AOI211_X1 U11062 ( .C1(n9834), .C2(n9833), .A(n9832), .B(n9831), .ZN(n9835)
         );
  AOI211_X1 U11063 ( .C1(n10568), .C2(n9837), .A(n9836), .B(n9835), .ZN(n9839)
         );
  NAND2_X1 U11064 ( .A1(P1_REG3_REG_16__SCAN_IN), .A2(P1_U3086), .ZN(n9838) );
  OAI211_X1 U11065 ( .C1(n9853), .C2(n10427), .A(n9839), .B(n9838), .ZN(
        P1_U3259) );
  OAI211_X1 U11066 ( .C1(n9842), .C2(n9841), .A(n9840), .B(n10559), .ZN(n9843)
         );
  INV_X1 U11067 ( .A(n9843), .ZN(n9849) );
  AOI211_X1 U11068 ( .C1(n9847), .C2(n9846), .A(n9845), .B(n9844), .ZN(n9848)
         );
  AOI211_X1 U11069 ( .C1(n10568), .C2(n9850), .A(n9849), .B(n9848), .ZN(n9852)
         );
  NAND2_X1 U11070 ( .A1(P1_REG3_REG_18__SCAN_IN), .A2(P1_U3086), .ZN(n9851) );
  OAI211_X1 U11071 ( .C1(n9853), .C2(n10166), .A(n9852), .B(n9851), .ZN(
        P1_U3261) );
  INV_X1 U11072 ( .A(n9854), .ZN(n9856) );
  AOI22_X1 U11073 ( .A1(n9857), .A2(P1_REG2_REG_4__SCAN_IN), .B1(n9856), .B2(
        n9855), .ZN(n9858) );
  OAI21_X1 U11074 ( .B1(n9860), .B2(n9859), .A(n9858), .ZN(n9864) );
  NOR2_X1 U11075 ( .A1(n9862), .A2(n9861), .ZN(n9863) );
  AOI211_X1 U11076 ( .C1(n9866), .C2(n9865), .A(n9864), .B(n9863), .ZN(n9867)
         );
  OAI21_X1 U11077 ( .B1(n9857), .B2(n9868), .A(n9867), .ZN(P1_U3289) );
  NOR2_X1 U11078 ( .A1(n9869), .A2(n6961), .ZN(n9870) );
  AOI21_X1 U11079 ( .B1(n9857), .B2(P1_REG2_REG_1__SCAN_IN), .A(n9870), .ZN(
        n9871) );
  OAI21_X1 U11080 ( .B1(n9873), .B2(n9872), .A(n9871), .ZN(n9874) );
  INV_X1 U11081 ( .A(n9874), .ZN(n9881) );
  INV_X1 U11082 ( .A(n9875), .ZN(n9876) );
  AOI22_X1 U11083 ( .A1(n9879), .A2(n9878), .B1(n9877), .B2(n9876), .ZN(n9880)
         );
  OAI211_X1 U11084 ( .C1(n9857), .C2(n9882), .A(n9881), .B(n9880), .ZN(
        P1_U3292) );
  AND2_X1 U11085 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n9884), .ZN(P1_U3294) );
  AND2_X1 U11086 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n9884), .ZN(P1_U3295) );
  AND2_X1 U11087 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n9884), .ZN(P1_U3296) );
  AND2_X1 U11088 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n9884), .ZN(P1_U3297) );
  AND2_X1 U11089 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n9884), .ZN(P1_U3298) );
  AND2_X1 U11090 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n9884), .ZN(P1_U3299) );
  AND2_X1 U11091 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n9884), .ZN(P1_U3300) );
  AND2_X1 U11092 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n9884), .ZN(P1_U3301) );
  INV_X1 U11093 ( .A(P1_D_REG_23__SCAN_IN), .ZN(n10441) );
  NOR2_X1 U11094 ( .A1(n9883), .A2(n10441), .ZN(P1_U3302) );
  AND2_X1 U11095 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n9884), .ZN(P1_U3303) );
  INV_X1 U11096 ( .A(P1_D_REG_21__SCAN_IN), .ZN(n10385) );
  NOR2_X1 U11097 ( .A1(n9883), .A2(n10385), .ZN(P1_U3304) );
  AND2_X1 U11098 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n9884), .ZN(P1_U3305) );
  AND2_X1 U11099 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n9884), .ZN(P1_U3306) );
  AND2_X1 U11100 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n9884), .ZN(P1_U3307) );
  AND2_X1 U11101 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n9884), .ZN(P1_U3308) );
  AND2_X1 U11102 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n9884), .ZN(P1_U3309) );
  AND2_X1 U11103 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n9884), .ZN(P1_U3310) );
  AND2_X1 U11104 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n9884), .ZN(P1_U3311) );
  AND2_X1 U11105 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n9884), .ZN(P1_U3312) );
  AND2_X1 U11106 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n9884), .ZN(P1_U3313) );
  AND2_X1 U11107 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n9884), .ZN(P1_U3314) );
  AND2_X1 U11108 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n9884), .ZN(P1_U3315) );
  AND2_X1 U11109 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n9884), .ZN(P1_U3316) );
  INV_X1 U11110 ( .A(P1_D_REG_8__SCAN_IN), .ZN(n10381) );
  NOR2_X1 U11111 ( .A1(n9883), .A2(n10381), .ZN(P1_U3317) );
  AND2_X1 U11112 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n9884), .ZN(P1_U3318) );
  AND2_X1 U11113 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n9884), .ZN(P1_U3319) );
  AND2_X1 U11114 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n9884), .ZN(P1_U3320) );
  INV_X1 U11115 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n10407) );
  NOR2_X1 U11116 ( .A1(n9883), .A2(n10407), .ZN(P1_U3321) );
  AND2_X1 U11117 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n9884), .ZN(P1_U3322) );
  AND2_X1 U11118 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n9884), .ZN(P1_U3323) );
  INV_X1 U11119 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n9885) );
  AOI22_X1 U11120 ( .A1(n9911), .A2(n9886), .B1(n9885), .B2(n9910), .ZN(
        P1_U3456) );
  OAI21_X1 U11121 ( .B1(n9888), .B2(n9905), .A(n9887), .ZN(n9890) );
  AOI211_X1 U11122 ( .C1(n9908), .C2(n9891), .A(n9890), .B(n9889), .ZN(n9913)
         );
  AOI22_X1 U11123 ( .A1(n9911), .A2(n9913), .B1(n5201), .B2(n9910), .ZN(
        P1_U3459) );
  OAI21_X1 U11124 ( .B1(n9893), .B2(n9905), .A(n9892), .ZN(n9895) );
  AOI211_X1 U11125 ( .C1(n9908), .C2(n9896), .A(n9895), .B(n9894), .ZN(n9914)
         );
  AOI22_X1 U11126 ( .A1(n9911), .A2(n9914), .B1(n5223), .B2(n9910), .ZN(
        P1_U3462) );
  OAI21_X1 U11127 ( .B1(n9898), .B2(n9905), .A(n9897), .ZN(n9901) );
  INV_X1 U11128 ( .A(n9899), .ZN(n9900) );
  AOI211_X1 U11129 ( .C1(n9908), .C2(n9902), .A(n9901), .B(n9900), .ZN(n9915)
         );
  AOI22_X1 U11130 ( .A1(n9911), .A2(n9915), .B1(n5304), .B2(n9910), .ZN(
        P1_U3474) );
  OAI211_X1 U11131 ( .C1(n9906), .C2(n9905), .A(n9904), .B(n9903), .ZN(n9907)
         );
  AOI21_X1 U11132 ( .B1(n9909), .B2(n9908), .A(n9907), .ZN(n9917) );
  AOI22_X1 U11133 ( .A1(n9911), .A2(n9917), .B1(n5441), .B2(n9910), .ZN(
        P1_U3492) );
  AOI22_X1 U11134 ( .A1(n9918), .A2(n9913), .B1(n9912), .B2(n9916), .ZN(
        P1_U3524) );
  INV_X1 U11135 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n10290) );
  AOI22_X1 U11136 ( .A1(n9918), .A2(n9914), .B1(n10290), .B2(n9916), .ZN(
        P1_U3525) );
  AOI22_X1 U11137 ( .A1(n9918), .A2(n9915), .B1(n6803), .B2(n9916), .ZN(
        P1_U3529) );
  AOI22_X1 U11138 ( .A1(n9918), .A2(n9917), .B1(n7551), .B2(n9916), .ZN(
        P1_U3535) );
  AOI22_X1 U11139 ( .A1(n10069), .A2(P2_IR_REG_0__SCAN_IN), .B1(n10067), .B2(
        P2_ADDR_REG_0__SCAN_IN), .ZN(n9924) );
  INV_X1 U11140 ( .A(n9919), .ZN(n9922) );
  XNOR2_X1 U11141 ( .A(n9920), .B(P2_IR_REG_0__SCAN_IN), .ZN(n9921) );
  OAI21_X1 U11142 ( .B1(n9922), .B2(n10058), .A(n9921), .ZN(n9923) );
  OAI211_X1 U11143 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n6217), .A(n9924), .B(
        n9923), .ZN(P2_U3182) );
  NAND2_X1 U11144 ( .A1(n9925), .A2(n7225), .ZN(n9926) );
  NAND2_X1 U11145 ( .A1(n9927), .A2(n9926), .ZN(n9929) );
  AOI22_X1 U11146 ( .A1(n9969), .A2(n9929), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        P2_U3151), .ZN(n9934) );
  OAI211_X1 U11147 ( .C1(n9932), .C2(n9931), .A(n9930), .B(n10058), .ZN(n9933)
         );
  OAI211_X1 U11148 ( .C1(n10051), .C2(n9935), .A(n9934), .B(n9933), .ZN(n9936)
         );
  INV_X1 U11149 ( .A(n9936), .ZN(n9943) );
  INV_X1 U11150 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n9940) );
  XNOR2_X1 U11151 ( .A(n9937), .B(n10467), .ZN(n9938) );
  OAI22_X1 U11152 ( .A1(n10049), .A2(n9940), .B1(n9939), .B2(n9938), .ZN(n9941) );
  INV_X1 U11153 ( .A(n9941), .ZN(n9942) );
  NAND2_X1 U11154 ( .A1(n9943), .A2(n9942), .ZN(P2_U3183) );
  INV_X1 U11155 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n9960) );
  XNOR2_X1 U11156 ( .A(n9944), .B(P2_REG1_REG_5__SCAN_IN), .ZN(n9958) );
  INV_X1 U11157 ( .A(n9945), .ZN(n9946) );
  NAND2_X1 U11158 ( .A1(n9946), .A2(n6274), .ZN(n9947) );
  NAND2_X1 U11159 ( .A1(n9964), .A2(n9947), .ZN(n9949) );
  AOI21_X1 U11160 ( .B1(n9969), .B2(n9949), .A(n9948), .ZN(n9950) );
  OAI21_X1 U11161 ( .B1(n9951), .B2(n10051), .A(n9950), .ZN(n9957) );
  OAI211_X1 U11162 ( .C1(n9954), .C2(n9953), .A(n9952), .B(n10058), .ZN(n9955)
         );
  INV_X1 U11163 ( .A(n9955), .ZN(n9956) );
  AOI211_X1 U11164 ( .C1(n10084), .C2(n9958), .A(n9957), .B(n9956), .ZN(n9959)
         );
  OAI21_X1 U11165 ( .B1(n10049), .B2(n9960), .A(n9959), .ZN(P2_U3187) );
  INV_X1 U11166 ( .A(n9961), .ZN(n9963) );
  NAND3_X1 U11167 ( .A1(n9964), .A2(n9963), .A3(n9962), .ZN(n9965) );
  NAND2_X1 U11168 ( .A1(n9966), .A2(n9965), .ZN(n9968) );
  AOI21_X1 U11169 ( .B1(n9969), .B2(n9968), .A(n9967), .ZN(n9975) );
  OAI21_X1 U11170 ( .B1(n9972), .B2(n9971), .A(n9970), .ZN(n9973) );
  NAND2_X1 U11171 ( .A1(n10084), .A2(n9973), .ZN(n9974) );
  OAI211_X1 U11172 ( .C1(n10051), .C2(n9976), .A(n9975), .B(n9974), .ZN(n9977)
         );
  INV_X1 U11173 ( .A(n9977), .ZN(n9984) );
  AOI21_X1 U11174 ( .B1(n9980), .B2(n9979), .A(n9978), .ZN(n9981) );
  NOR2_X1 U11175 ( .A1(n9981), .A2(n10079), .ZN(n9982) );
  AOI21_X1 U11176 ( .B1(n10067), .B2(P2_ADDR_REG_6__SCAN_IN), .A(n9982), .ZN(
        n9983) );
  NAND2_X1 U11177 ( .A1(n9984), .A2(n9983), .ZN(P2_U3188) );
  OAI21_X1 U11178 ( .B1(P2_REG1_REG_7__SCAN_IN), .B2(n9986), .A(n9985), .ZN(
        n9995) );
  INV_X1 U11179 ( .A(n9987), .ZN(n9988) );
  OAI21_X1 U11180 ( .B1(n10051), .B2(n9989), .A(n9988), .ZN(n9994) );
  AOI21_X1 U11181 ( .B1(n6312), .B2(n9991), .A(n9990), .ZN(n9992) );
  NOR2_X1 U11182 ( .A1(n9992), .A2(n10089), .ZN(n9993) );
  AOI211_X1 U11183 ( .C1(n10084), .C2(n9995), .A(n9994), .B(n9993), .ZN(n10000) );
  XNOR2_X1 U11184 ( .A(n9997), .B(n9996), .ZN(n9998) );
  AOI22_X1 U11185 ( .A1(n9998), .A2(n10058), .B1(n10067), .B2(
        P2_ADDR_REG_7__SCAN_IN), .ZN(n9999) );
  NAND2_X1 U11186 ( .A1(n10000), .A2(n9999), .ZN(P2_U3189) );
  OAI21_X1 U11187 ( .B1(n10003), .B2(n10002), .A(n10001), .ZN(n10005) );
  AOI22_X1 U11188 ( .A1(n10005), .A2(n10084), .B1(n10004), .B2(n10069), .ZN(
        n10016) );
  XNOR2_X1 U11189 ( .A(n10007), .B(n10006), .ZN(n10008) );
  AOI22_X1 U11190 ( .A1(n10008), .A2(n10058), .B1(n10067), .B2(
        P2_ADDR_REG_8__SCAN_IN), .ZN(n10015) );
  AOI21_X1 U11191 ( .B1(n10011), .B2(n10010), .A(n10009), .ZN(n10012) );
  OR2_X1 U11192 ( .A1(n10012), .A2(n10089), .ZN(n10013) );
  NAND4_X1 U11193 ( .A1(n10016), .A2(n10015), .A3(n10014), .A4(n10013), .ZN(
        P2_U3190) );
  AOI22_X1 U11194 ( .A1(n10069), .A2(n10017), .B1(n10067), .B2(
        P2_ADDR_REG_9__SCAN_IN), .ZN(n10030) );
  XNOR2_X1 U11195 ( .A(n10019), .B(n10018), .ZN(n10023) );
  OAI21_X1 U11196 ( .B1(P2_REG1_REG_9__SCAN_IN), .B2(n10021), .A(n10020), .ZN(
        n10022) );
  AOI22_X1 U11197 ( .A1(n10023), .A2(n10058), .B1(n10084), .B2(n10022), .ZN(
        n10029) );
  AOI21_X1 U11198 ( .B1(n10025), .B2(n6341), .A(n10024), .ZN(n10026) );
  OR2_X1 U11199 ( .A1(n10089), .A2(n10026), .ZN(n10027) );
  NAND4_X1 U11200 ( .A1(n10030), .A2(n10029), .A3(n10028), .A4(n10027), .ZN(
        P2_U3191) );
  AOI22_X1 U11201 ( .A1(n10069), .A2(n10031), .B1(n10067), .B2(
        P2_ADDR_REG_10__SCAN_IN), .ZN(n10047) );
  XNOR2_X1 U11202 ( .A(n10033), .B(n10032), .ZN(n10038) );
  OAI21_X1 U11203 ( .B1(n10036), .B2(n10035), .A(n10034), .ZN(n10037) );
  AOI22_X1 U11204 ( .A1(n10038), .A2(n10058), .B1(n10084), .B2(n10037), .ZN(
        n10046) );
  INV_X1 U11205 ( .A(n10039), .ZN(n10045) );
  AOI21_X1 U11206 ( .B1(n10042), .B2(n10041), .A(n10040), .ZN(n10043) );
  OR2_X1 U11207 ( .A1(n10043), .A2(n10089), .ZN(n10044) );
  NAND4_X1 U11208 ( .A1(n10047), .A2(n10046), .A3(n10045), .A4(n10044), .ZN(
        P2_U3192) );
  INV_X1 U11209 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n10048) );
  OAI22_X1 U11210 ( .A1(n10051), .A2(n10050), .B1(n10049), .B2(n10048), .ZN(
        n10052) );
  INV_X1 U11211 ( .A(n10052), .ZN(n10066) );
  XNOR2_X1 U11212 ( .A(n10054), .B(n10053), .ZN(n10059) );
  OAI21_X1 U11213 ( .B1(n10056), .B2(P2_REG1_REG_11__SCAN_IN), .A(n10055), 
        .ZN(n10057) );
  AOI22_X1 U11214 ( .A1(n10059), .A2(n10058), .B1(n10084), .B2(n10057), .ZN(
        n10065) );
  AOI21_X1 U11215 ( .B1(n7818), .B2(n10061), .A(n10060), .ZN(n10062) );
  OR2_X1 U11216 ( .A1(n10089), .A2(n10062), .ZN(n10063) );
  NAND4_X1 U11217 ( .A1(n10066), .A2(n10065), .A3(n10064), .A4(n10063), .ZN(
        P2_U3193) );
  AOI22_X1 U11218 ( .A1(n10069), .A2(n10068), .B1(n10067), .B2(
        P2_ADDR_REG_12__SCAN_IN), .ZN(n10093) );
  OAI21_X1 U11219 ( .B1(n10072), .B2(n10071), .A(n10070), .ZN(n10083) );
  INV_X1 U11220 ( .A(n10073), .ZN(n10081) );
  AOI21_X1 U11221 ( .B1(n10074), .B2(n10073), .A(n10080), .ZN(n10077) );
  INV_X1 U11222 ( .A(n10075), .ZN(n10076) );
  NOR2_X1 U11223 ( .A1(n10077), .A2(n10076), .ZN(n10078) );
  AOI211_X1 U11224 ( .C1(n10081), .C2(n10080), .A(n10079), .B(n10078), .ZN(
        n10082) );
  AOI21_X1 U11225 ( .B1(n10084), .B2(n10083), .A(n10082), .ZN(n10092) );
  AOI21_X1 U11226 ( .B1(n10087), .B2(n10086), .A(n10085), .ZN(n10088) );
  OR2_X1 U11227 ( .A1(n10089), .A2(n10088), .ZN(n10090) );
  NAND4_X1 U11228 ( .A1(n10093), .A2(n10092), .A3(n10091), .A4(n10090), .ZN(
        P2_U3194) );
  NAND2_X1 U11229 ( .A1(n10095), .A2(n10094), .ZN(n10096) );
  OAI21_X1 U11230 ( .B1(n10097), .B2(n6228), .A(n10096), .ZN(n10100) );
  INV_X1 U11231 ( .A(n10098), .ZN(n10099) );
  AOI211_X1 U11232 ( .C1(n10102), .C2(n10101), .A(n10100), .B(n10099), .ZN(
        n10104) );
  AOI22_X1 U11233 ( .A1(n10105), .A2(n6724), .B1(n10104), .B2(n10103), .ZN(
        P2_U3231) );
  INV_X1 U11234 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n10107) );
  AOI22_X1 U11235 ( .A1(n10149), .A2(n10107), .B1(n10106), .B2(n10148), .ZN(
        P2_U3393) );
  AOI22_X1 U11236 ( .A1(n10149), .A2(n6227), .B1(n10108), .B2(n10148), .ZN(
        P2_U3396) );
  AOI22_X1 U11237 ( .A1(n10110), .A2(n10123), .B1(n10147), .B2(n10109), .ZN(
        n10111) );
  AND2_X1 U11238 ( .A1(n10112), .A2(n10111), .ZN(n10151) );
  AOI22_X1 U11239 ( .A1(n10149), .A2(n6239), .B1(n10151), .B2(n10148), .ZN(
        P2_U3399) );
  INV_X1 U11240 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n10118) );
  INV_X1 U11241 ( .A(n10123), .ZN(n10130) );
  NOR2_X1 U11242 ( .A1(n10113), .A2(n10130), .ZN(n10116) );
  INV_X1 U11243 ( .A(n10114), .ZN(n10115) );
  AOI211_X1 U11244 ( .C1(n10147), .C2(n10117), .A(n10116), .B(n10115), .ZN(
        n10152) );
  AOI22_X1 U11245 ( .A1(n10149), .A2(n10118), .B1(n10152), .B2(n10148), .ZN(
        P2_U3402) );
  NOR2_X1 U11246 ( .A1(n10120), .A2(n10119), .ZN(n10122) );
  AOI211_X1 U11247 ( .C1(n10124), .C2(n10123), .A(n10122), .B(n10121), .ZN(
        n10153) );
  AOI22_X1 U11248 ( .A1(n10149), .A2(n6294), .B1(n10153), .B2(n10148), .ZN(
        P2_U3408) );
  INV_X1 U11249 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n10129) );
  NOR2_X1 U11250 ( .A1(n10125), .A2(n10141), .ZN(n10127) );
  AOI211_X1 U11251 ( .C1(n10147), .C2(n10128), .A(n10127), .B(n10126), .ZN(
        n10154) );
  AOI22_X1 U11252 ( .A1(n10149), .A2(n10129), .B1(n10154), .B2(n10148), .ZN(
        P2_U3411) );
  INV_X1 U11253 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n10135) );
  NOR2_X1 U11254 ( .A1(n10131), .A2(n10130), .ZN(n10133) );
  AOI211_X1 U11255 ( .C1(n10147), .C2(n10134), .A(n10133), .B(n10132), .ZN(
        n10155) );
  AOI22_X1 U11256 ( .A1(n10149), .A2(n10135), .B1(n10155), .B2(n10148), .ZN(
        P2_U3414) );
  INV_X1 U11257 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n10140) );
  NOR2_X1 U11258 ( .A1(n10136), .A2(n10141), .ZN(n10138) );
  AOI211_X1 U11259 ( .C1(n10147), .C2(n10139), .A(n10138), .B(n10137), .ZN(
        n10156) );
  AOI22_X1 U11260 ( .A1(n10149), .A2(n10140), .B1(n10156), .B2(n10148), .ZN(
        P2_U3417) );
  INV_X1 U11261 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n10365) );
  NOR2_X1 U11262 ( .A1(n10142), .A2(n10141), .ZN(n10145) );
  INV_X1 U11263 ( .A(n10143), .ZN(n10144) );
  AOI211_X1 U11264 ( .C1(n10147), .C2(n10146), .A(n10145), .B(n10144), .ZN(
        n10158) );
  AOI22_X1 U11265 ( .A1(n10149), .A2(n10365), .B1(n10158), .B2(n10148), .ZN(
        P2_U3420) );
  AOI22_X1 U11266 ( .A1(n10159), .A2(n10151), .B1(n10150), .B2(n10157), .ZN(
        P2_U3462) );
  AOI22_X1 U11267 ( .A1(n10159), .A2(n10152), .B1(n6777), .B2(n10157), .ZN(
        P2_U3463) );
  AOI22_X1 U11268 ( .A1(n10159), .A2(n10153), .B1(n7779), .B2(n10157), .ZN(
        P2_U3465) );
  AOI22_X1 U11269 ( .A1(n10159), .A2(n10154), .B1(n6315), .B2(n10157), .ZN(
        P2_U3466) );
  AOI22_X1 U11270 ( .A1(n10159), .A2(n10155), .B1(n6326), .B2(n10157), .ZN(
        P2_U3467) );
  AOI22_X1 U11271 ( .A1(n10159), .A2(n10156), .B1(n6338), .B2(n10157), .ZN(
        P2_U3468) );
  AOI22_X1 U11272 ( .A1(n10159), .A2(n10158), .B1(n6356), .B2(n10157), .ZN(
        P2_U3469) );
  OAI21_X1 U11273 ( .B1(n10163), .B2(n10161), .A(n10160), .ZN(n10162) );
  XNOR2_X1 U11274 ( .A(n10162), .B(P2_ADDR_REG_1__SCAN_IN), .ZN(ADD_1068_U5)
         );
  OAI21_X1 U11275 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(P2_ADDR_REG_0__SCAN_IN), 
        .A(n10163), .ZN(n10164) );
  INV_X1 U11276 ( .A(n10164), .ZN(ADD_1068_U46) );
  OAI21_X1 U11277 ( .B1(n10167), .B2(n10166), .A(n10165), .ZN(n10168) );
  XNOR2_X1 U11278 ( .A(n10168), .B(P2_ADDR_REG_18__SCAN_IN), .ZN(ADD_1068_U55)
         );
  OAI21_X1 U11279 ( .B1(n10171), .B2(n10170), .A(n10169), .ZN(ADD_1068_U56) );
  OAI21_X1 U11280 ( .B1(n10174), .B2(n10173), .A(n10172), .ZN(ADD_1068_U57) );
  OAI21_X1 U11281 ( .B1(n10177), .B2(n10176), .A(n10175), .ZN(ADD_1068_U58) );
  OAI21_X1 U11282 ( .B1(n10180), .B2(n10179), .A(n10178), .ZN(ADD_1068_U59) );
  OAI21_X1 U11283 ( .B1(n10183), .B2(n10182), .A(n10181), .ZN(ADD_1068_U60) );
  OAI21_X1 U11284 ( .B1(n10186), .B2(n10185), .A(n10184), .ZN(ADD_1068_U61) );
  OAI21_X1 U11285 ( .B1(n10189), .B2(n10188), .A(n10187), .ZN(ADD_1068_U62) );
  OAI21_X1 U11286 ( .B1(n10192), .B2(n10191), .A(n10190), .ZN(ADD_1068_U63) );
  AOI22_X1 U11287 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(keyinput233), .B1(SI_16_), 
        .B2(keyinput145), .ZN(n10193) );
  OAI221_X1 U11288 ( .B1(P1_REG3_REG_8__SCAN_IN), .B2(keyinput233), .C1(SI_16_), .C2(keyinput145), .A(n10193), .ZN(n10200) );
  AOI22_X1 U11289 ( .A1(P2_DATAO_REG_12__SCAN_IN), .A2(keyinput207), .B1(
        P1_DATAO_REG_20__SCAN_IN), .B2(keyinput229), .ZN(n10194) );
  OAI221_X1 U11290 ( .B1(P2_DATAO_REG_12__SCAN_IN), .B2(keyinput207), .C1(
        P1_DATAO_REG_20__SCAN_IN), .C2(keyinput229), .A(n10194), .ZN(n10199)
         );
  AOI22_X1 U11291 ( .A1(P1_DATAO_REG_4__SCAN_IN), .A2(keyinput188), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(keyinput179), .ZN(n10195) );
  OAI221_X1 U11292 ( .B1(P1_DATAO_REG_4__SCAN_IN), .B2(keyinput188), .C1(
        P2_DATAO_REG_10__SCAN_IN), .C2(keyinput179), .A(n10195), .ZN(n10198)
         );
  AOI22_X1 U11293 ( .A1(P1_REG2_REG_19__SCAN_IN), .A2(keyinput250), .B1(
        P1_IR_REG_25__SCAN_IN), .B2(keyinput252), .ZN(n10196) );
  OAI221_X1 U11294 ( .B1(P1_REG2_REG_19__SCAN_IN), .B2(keyinput250), .C1(
        P1_IR_REG_25__SCAN_IN), .C2(keyinput252), .A(n10196), .ZN(n10197) );
  NOR4_X1 U11295 ( .A1(n10200), .A2(n10199), .A3(n10198), .A4(n10197), .ZN(
        n10228) );
  AOI22_X1 U11296 ( .A1(P2_REG1_REG_31__SCAN_IN), .A2(keyinput147), .B1(SI_18_), .B2(keyinput164), .ZN(n10201) );
  OAI221_X1 U11297 ( .B1(P2_REG1_REG_31__SCAN_IN), .B2(keyinput147), .C1(
        SI_18_), .C2(keyinput164), .A(n10201), .ZN(n10208) );
  AOI22_X1 U11298 ( .A1(P2_REG1_REG_14__SCAN_IN), .A2(keyinput243), .B1(SI_1_), 
        .B2(keyinput214), .ZN(n10202) );
  OAI221_X1 U11299 ( .B1(P2_REG1_REG_14__SCAN_IN), .B2(keyinput243), .C1(SI_1_), .C2(keyinput214), .A(n10202), .ZN(n10207) );
  AOI22_X1 U11300 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(keyinput246), .B1(
        P1_D_REG_23__SCAN_IN), .B2(keyinput154), .ZN(n10203) );
  OAI221_X1 U11301 ( .B1(P1_ADDR_REG_5__SCAN_IN), .B2(keyinput246), .C1(
        P1_D_REG_23__SCAN_IN), .C2(keyinput154), .A(n10203), .ZN(n10206) );
  AOI22_X1 U11302 ( .A1(P2_D_REG_20__SCAN_IN), .A2(keyinput199), .B1(
        P1_REG0_REG_21__SCAN_IN), .B2(keyinput167), .ZN(n10204) );
  OAI221_X1 U11303 ( .B1(P2_D_REG_20__SCAN_IN), .B2(keyinput199), .C1(
        P1_REG0_REG_21__SCAN_IN), .C2(keyinput167), .A(n10204), .ZN(n10205) );
  NOR4_X1 U11304 ( .A1(n10208), .A2(n10207), .A3(n10206), .A4(n10205), .ZN(
        n10227) );
  AOI22_X1 U11305 ( .A1(P1_REG1_REG_12__SCAN_IN), .A2(keyinput204), .B1(
        P1_IR_REG_0__SCAN_IN), .B2(keyinput182), .ZN(n10209) );
  OAI221_X1 U11306 ( .B1(P1_REG1_REG_12__SCAN_IN), .B2(keyinput204), .C1(
        P1_IR_REG_0__SCAN_IN), .C2(keyinput182), .A(n10209), .ZN(n10216) );
  AOI22_X1 U11307 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(keyinput128), .B1(
        P1_DATAO_REG_10__SCAN_IN), .B2(keyinput200), .ZN(n10210) );
  OAI221_X1 U11308 ( .B1(P2_ADDR_REG_5__SCAN_IN), .B2(keyinput128), .C1(
        P1_DATAO_REG_10__SCAN_IN), .C2(keyinput200), .A(n10210), .ZN(n10215)
         );
  AOI22_X1 U11309 ( .A1(P2_D_REG_9__SCAN_IN), .A2(keyinput175), .B1(
        P2_IR_REG_19__SCAN_IN), .B2(keyinput180), .ZN(n10211) );
  OAI221_X1 U11310 ( .B1(P2_D_REG_9__SCAN_IN), .B2(keyinput175), .C1(
        P2_IR_REG_19__SCAN_IN), .C2(keyinput180), .A(n10211), .ZN(n10214) );
  AOI22_X1 U11311 ( .A1(P2_IR_REG_30__SCAN_IN), .A2(keyinput251), .B1(
        P1_DATAO_REG_23__SCAN_IN), .B2(keyinput187), .ZN(n10212) );
  OAI221_X1 U11312 ( .B1(P2_IR_REG_30__SCAN_IN), .B2(keyinput251), .C1(
        P1_DATAO_REG_23__SCAN_IN), .C2(keyinput187), .A(n10212), .ZN(n10213)
         );
  NOR4_X1 U11313 ( .A1(n10216), .A2(n10215), .A3(n10214), .A4(n10213), .ZN(
        n10226) );
  AOI22_X1 U11314 ( .A1(P2_REG1_REG_1__SCAN_IN), .A2(keyinput181), .B1(
        P2_IR_REG_24__SCAN_IN), .B2(keyinput249), .ZN(n10217) );
  OAI221_X1 U11315 ( .B1(P2_REG1_REG_1__SCAN_IN), .B2(keyinput181), .C1(
        P2_IR_REG_24__SCAN_IN), .C2(keyinput249), .A(n10217), .ZN(n10224) );
  AOI22_X1 U11316 ( .A1(P2_REG3_REG_2__SCAN_IN), .A2(keyinput140), .B1(
        P2_REG2_REG_9__SCAN_IN), .B2(keyinput160), .ZN(n10218) );
  OAI221_X1 U11317 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(keyinput140), .C1(
        P2_REG2_REG_9__SCAN_IN), .C2(keyinput160), .A(n10218), .ZN(n10223) );
  AOI22_X1 U11318 ( .A1(P1_REG2_REG_20__SCAN_IN), .A2(keyinput152), .B1(
        P1_REG1_REG_23__SCAN_IN), .B2(keyinput162), .ZN(n10219) );
  OAI221_X1 U11319 ( .B1(P1_REG2_REG_20__SCAN_IN), .B2(keyinput152), .C1(
        P1_REG1_REG_23__SCAN_IN), .C2(keyinput162), .A(n10219), .ZN(n10222) );
  AOI22_X1 U11320 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(keyinput254), .B1(
        P2_REG2_REG_18__SCAN_IN), .B2(keyinput231), .ZN(n10220) );
  OAI221_X1 U11321 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(keyinput254), .C1(
        P2_REG2_REG_18__SCAN_IN), .C2(keyinput231), .A(n10220), .ZN(n10221) );
  NOR4_X1 U11322 ( .A1(n10224), .A2(n10223), .A3(n10222), .A4(n10221), .ZN(
        n10225) );
  NAND4_X1 U11323 ( .A1(n10228), .A2(n10227), .A3(n10226), .A4(n10225), .ZN(
        n10363) );
  AOI22_X1 U11324 ( .A1(P1_REG2_REG_22__SCAN_IN), .A2(keyinput206), .B1(
        P1_IR_REG_14__SCAN_IN), .B2(keyinput221), .ZN(n10229) );
  OAI221_X1 U11325 ( .B1(P1_REG2_REG_22__SCAN_IN), .B2(keyinput206), .C1(
        P1_IR_REG_14__SCAN_IN), .C2(keyinput221), .A(n10229), .ZN(n10236) );
  AOI22_X1 U11326 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(keyinput142), .B1(
        P1_REG1_REG_7__SCAN_IN), .B2(keyinput245), .ZN(n10230) );
  OAI221_X1 U11327 ( .B1(P2_REG3_REG_17__SCAN_IN), .B2(keyinput142), .C1(
        P1_REG1_REG_7__SCAN_IN), .C2(keyinput245), .A(n10230), .ZN(n10235) );
  AOI22_X1 U11328 ( .A1(P1_ADDR_REG_16__SCAN_IN), .A2(keyinput177), .B1(
        P1_REG2_REG_29__SCAN_IN), .B2(keyinput255), .ZN(n10231) );
  OAI221_X1 U11329 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(keyinput177), .C1(
        P1_REG2_REG_29__SCAN_IN), .C2(keyinput255), .A(n10231), .ZN(n10234) );
  AOI22_X1 U11330 ( .A1(P1_ADDR_REG_15__SCAN_IN), .A2(keyinput223), .B1(
        P2_REG0_REG_28__SCAN_IN), .B2(keyinput158), .ZN(n10232) );
  OAI221_X1 U11331 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(keyinput223), .C1(
        P2_REG0_REG_28__SCAN_IN), .C2(keyinput158), .A(n10232), .ZN(n10233) );
  NOR4_X1 U11332 ( .A1(n10236), .A2(n10235), .A3(n10234), .A4(n10233), .ZN(
        n10266) );
  AOI22_X1 U11333 ( .A1(P2_DATAO_REG_2__SCAN_IN), .A2(keyinput139), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(keyinput174), .ZN(n10237) );
  OAI221_X1 U11334 ( .B1(P2_DATAO_REG_2__SCAN_IN), .B2(keyinput139), .C1(
        P2_DATAO_REG_17__SCAN_IN), .C2(keyinput174), .A(n10237), .ZN(n10244)
         );
  AOI22_X1 U11335 ( .A1(P2_REG1_REG_13__SCAN_IN), .A2(keyinput209), .B1(
        P1_REG0_REG_14__SCAN_IN), .B2(keyinput132), .ZN(n10238) );
  OAI221_X1 U11336 ( .B1(P2_REG1_REG_13__SCAN_IN), .B2(keyinput209), .C1(
        P1_REG0_REG_14__SCAN_IN), .C2(keyinput132), .A(n10238), .ZN(n10243) );
  AOI22_X1 U11337 ( .A1(P2_ADDR_REG_19__SCAN_IN), .A2(keyinput170), .B1(
        P1_IR_REG_27__SCAN_IN), .B2(keyinput215), .ZN(n10239) );
  OAI221_X1 U11338 ( .B1(P2_ADDR_REG_19__SCAN_IN), .B2(keyinput170), .C1(
        P1_IR_REG_27__SCAN_IN), .C2(keyinput215), .A(n10239), .ZN(n10242) );
  AOI22_X1 U11339 ( .A1(P2_REG0_REG_15__SCAN_IN), .A2(keyinput183), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(keyinput194), .ZN(n10240) );
  OAI221_X1 U11340 ( .B1(P2_REG0_REG_15__SCAN_IN), .B2(keyinput183), .C1(
        P2_DATAO_REG_18__SCAN_IN), .C2(keyinput194), .A(n10240), .ZN(n10241)
         );
  NOR4_X1 U11341 ( .A1(n10244), .A2(n10243), .A3(n10242), .A4(n10241), .ZN(
        n10265) );
  AOI22_X1 U11342 ( .A1(P2_REG0_REG_18__SCAN_IN), .A2(keyinput129), .B1(
        P1_IR_REG_26__SCAN_IN), .B2(keyinput211), .ZN(n10245) );
  OAI221_X1 U11343 ( .B1(P2_REG0_REG_18__SCAN_IN), .B2(keyinput129), .C1(
        P1_IR_REG_26__SCAN_IN), .C2(keyinput211), .A(n10245), .ZN(n10252) );
  AOI22_X1 U11344 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(keyinput137), .B1(
        P2_REG3_REG_4__SCAN_IN), .B2(keyinput208), .ZN(n10246) );
  OAI221_X1 U11345 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(keyinput137), .C1(
        P2_REG3_REG_4__SCAN_IN), .C2(keyinput208), .A(n10246), .ZN(n10251) );
  AOI22_X1 U11346 ( .A1(P2_ADDR_REG_0__SCAN_IN), .A2(keyinput159), .B1(
        P2_REG0_REG_20__SCAN_IN), .B2(keyinput203), .ZN(n10247) );
  OAI221_X1 U11347 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(keyinput159), .C1(
        P2_REG0_REG_20__SCAN_IN), .C2(keyinput203), .A(n10247), .ZN(n10250) );
  AOI22_X1 U11348 ( .A1(P1_REG1_REG_27__SCAN_IN), .A2(keyinput210), .B1(
        P1_REG3_REG_7__SCAN_IN), .B2(keyinput230), .ZN(n10248) );
  OAI221_X1 U11349 ( .B1(P1_REG1_REG_27__SCAN_IN), .B2(keyinput210), .C1(
        P1_REG3_REG_7__SCAN_IN), .C2(keyinput230), .A(n10248), .ZN(n10249) );
  NOR4_X1 U11350 ( .A1(n10252), .A2(n10251), .A3(n10250), .A4(n10249), .ZN(
        n10264) );
  AOI22_X1 U11351 ( .A1(n5201), .A2(keyinput225), .B1(keyinput163), .B2(n10466), .ZN(n10253) );
  OAI221_X1 U11352 ( .B1(n5201), .B2(keyinput225), .C1(n10466), .C2(
        keyinput163), .A(n10253), .ZN(n10262) );
  INV_X1 U11353 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n10414) );
  AOI22_X1 U11354 ( .A1(n6326), .A2(keyinput235), .B1(n10414), .B2(keyinput171), .ZN(n10254) );
  OAI221_X1 U11355 ( .B1(n6326), .B2(keyinput235), .C1(n10414), .C2(
        keyinput171), .A(n10254), .ZN(n10261) );
  XNOR2_X1 U11356 ( .A(n10456), .B(keyinput212), .ZN(n10257) );
  XNOR2_X1 U11357 ( .A(P1_REG1_REG_1__SCAN_IN), .B(keyinput213), .ZN(n10256)
         );
  XNOR2_X1 U11358 ( .A(P1_REG2_REG_0__SCAN_IN), .B(keyinput237), .ZN(n10255)
         );
  NAND3_X1 U11359 ( .A1(n10257), .A2(n10256), .A3(n10255), .ZN(n10260) );
  XNOR2_X1 U11360 ( .A(n10258), .B(keyinput238), .ZN(n10259) );
  NOR4_X1 U11361 ( .A1(n10262), .A2(n10261), .A3(n10260), .A4(n10259), .ZN(
        n10263) );
  NAND4_X1 U11362 ( .A1(n10266), .A2(n10265), .A3(n10264), .A4(n10263), .ZN(
        n10362) );
  AOI22_X1 U11363 ( .A1(n10407), .A2(keyinput247), .B1(keyinput135), .B2(
        n10268), .ZN(n10267) );
  OAI221_X1 U11364 ( .B1(n10407), .B2(keyinput247), .C1(n10268), .C2(
        keyinput135), .A(n10267), .ZN(n10275) );
  AOI22_X1 U11365 ( .A1(n10410), .A2(keyinput161), .B1(n10381), .B2(
        keyinput217), .ZN(n10269) );
  OAI221_X1 U11366 ( .B1(n10410), .B2(keyinput161), .C1(n10381), .C2(
        keyinput217), .A(n10269), .ZN(n10274) );
  AOI22_X1 U11367 ( .A1(n10371), .A2(keyinput236), .B1(keyinput227), .B2(
        n10365), .ZN(n10270) );
  OAI221_X1 U11368 ( .B1(n10371), .B2(keyinput236), .C1(n10365), .C2(
        keyinput227), .A(n10270), .ZN(n10273) );
  AOI22_X1 U11369 ( .A1(n8476), .A2(keyinput153), .B1(n10443), .B2(keyinput228), .ZN(n10271) );
  OAI221_X1 U11370 ( .B1(n8476), .B2(keyinput153), .C1(n10443), .C2(
        keyinput228), .A(n10271), .ZN(n10272) );
  NOR4_X1 U11371 ( .A1(n10275), .A2(n10274), .A3(n10273), .A4(n10272), .ZN(
        n10311) );
  AOI22_X1 U11372 ( .A1(n10277), .A2(keyinput156), .B1(n5189), .B2(keyinput143), .ZN(n10276) );
  OAI221_X1 U11373 ( .B1(n10277), .B2(keyinput156), .C1(n5189), .C2(
        keyinput143), .A(n10276), .ZN(n10287) );
  AOI22_X1 U11374 ( .A1(n7247), .A2(keyinput226), .B1(keyinput149), .B2(n10279), .ZN(n10278) );
  OAI221_X1 U11375 ( .B1(n7247), .B2(keyinput226), .C1(n10279), .C2(
        keyinput149), .A(n10278), .ZN(n10286) );
  AOI22_X1 U11376 ( .A1(n10281), .A2(keyinput168), .B1(n5415), .B2(keyinput196), .ZN(n10280) );
  OAI221_X1 U11377 ( .B1(n10281), .B2(keyinput168), .C1(n5415), .C2(
        keyinput196), .A(n10280), .ZN(n10285) );
  AOI22_X1 U11378 ( .A1(n10283), .A2(keyinput133), .B1(keyinput150), .B2(
        n10411), .ZN(n10282) );
  OAI221_X1 U11379 ( .B1(n10283), .B2(keyinput133), .C1(n10411), .C2(
        keyinput150), .A(n10282), .ZN(n10284) );
  NOR4_X1 U11380 ( .A1(n10287), .A2(n10286), .A3(n10285), .A4(n10284), .ZN(
        n10310) );
  AOI22_X1 U11381 ( .A1(n10385), .A2(keyinput220), .B1(keyinput244), .B2(n8536), .ZN(n10288) );
  OAI221_X1 U11382 ( .B1(n10385), .B2(keyinput220), .C1(n8536), .C2(
        keyinput244), .A(n10288), .ZN(n10297) );
  AOI22_X1 U11383 ( .A1(n6227), .A2(keyinput134), .B1(n10290), .B2(keyinput136), .ZN(n10289) );
  OAI221_X1 U11384 ( .B1(n6227), .B2(keyinput134), .C1(n10290), .C2(
        keyinput136), .A(n10289), .ZN(n10296) );
  AOI22_X1 U11385 ( .A1(n10384), .A2(keyinput218), .B1(n5149), .B2(keyinput241), .ZN(n10291) );
  OAI221_X1 U11386 ( .B1(n10384), .B2(keyinput218), .C1(n5149), .C2(
        keyinput241), .A(n10291), .ZN(n10295) );
  XNOR2_X1 U11387 ( .A(P2_REG1_REG_2__SCAN_IN), .B(keyinput193), .ZN(n10293)
         );
  XNOR2_X1 U11388 ( .A(SI_29_), .B(keyinput172), .ZN(n10292) );
  NAND2_X1 U11389 ( .A1(n10293), .A2(n10292), .ZN(n10294) );
  NOR4_X1 U11390 ( .A1(n10297), .A2(n10296), .A3(n10295), .A4(n10294), .ZN(
        n10309) );
  AOI22_X1 U11391 ( .A1(n7706), .A2(keyinput222), .B1(keyinput253), .B2(n10299), .ZN(n10298) );
  OAI221_X1 U11392 ( .B1(n7706), .B2(keyinput222), .C1(n10299), .C2(
        keyinput253), .A(n10298), .ZN(n10307) );
  AOI22_X1 U11393 ( .A1(n10397), .A2(keyinput191), .B1(keyinput169), .B2(
        n10301), .ZN(n10300) );
  OAI221_X1 U11394 ( .B1(n10397), .B2(keyinput191), .C1(n10301), .C2(
        keyinput169), .A(n10300), .ZN(n10306) );
  AOI22_X1 U11395 ( .A1(n10428), .A2(keyinput186), .B1(keyinput141), .B2(
        n10416), .ZN(n10302) );
  OAI221_X1 U11396 ( .B1(n10428), .B2(keyinput186), .C1(n10416), .C2(
        keyinput141), .A(n10302), .ZN(n10305) );
  AOI22_X1 U11397 ( .A1(n10382), .A2(keyinput198), .B1(keyinput184), .B2(
        n10454), .ZN(n10303) );
  OAI221_X1 U11398 ( .B1(n10382), .B2(keyinput198), .C1(n10454), .C2(
        keyinput184), .A(n10303), .ZN(n10304) );
  NOR4_X1 U11399 ( .A1(n10307), .A2(n10306), .A3(n10305), .A4(n10304), .ZN(
        n10308) );
  NAND4_X1 U11400 ( .A1(n10311), .A2(n10310), .A3(n10309), .A4(n10308), .ZN(
        n10361) );
  AOI22_X1 U11401 ( .A1(n10408), .A2(keyinput248), .B1(n5741), .B2(keyinput242), .ZN(n10312) );
  OAI221_X1 U11402 ( .B1(n10408), .B2(keyinput248), .C1(n5741), .C2(
        keyinput242), .A(n10312), .ZN(n10322) );
  AOI22_X1 U11403 ( .A1(n10445), .A2(keyinput178), .B1(keyinput146), .B2(n5243), .ZN(n10313) );
  OAI221_X1 U11404 ( .B1(n10445), .B2(keyinput178), .C1(n5243), .C2(
        keyinput146), .A(n10313), .ZN(n10321) );
  AOI22_X1 U11405 ( .A1(n10316), .A2(keyinput224), .B1(keyinput157), .B2(
        n10315), .ZN(n10314) );
  OAI221_X1 U11406 ( .B1(n10316), .B2(keyinput224), .C1(n10315), .C2(
        keyinput157), .A(n10314), .ZN(n10320) );
  XOR2_X1 U11407 ( .A(n6294), .B(keyinput144), .Z(n10318) );
  XNOR2_X1 U11408 ( .A(P1_IR_REG_12__SCAN_IN), .B(keyinput185), .ZN(n10317) );
  NAND2_X1 U11409 ( .A1(n10318), .A2(n10317), .ZN(n10319) );
  NOR4_X1 U11410 ( .A1(n10322), .A2(n10321), .A3(n10320), .A4(n10319), .ZN(
        n10359) );
  INV_X1 U11411 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n10398) );
  AOI22_X1 U11412 ( .A1(n10324), .A2(keyinput201), .B1(keyinput197), .B2(
        n10398), .ZN(n10323) );
  OAI221_X1 U11413 ( .B1(n10324), .B2(keyinput201), .C1(n10398), .C2(
        keyinput197), .A(n10323), .ZN(n10333) );
  AOI22_X1 U11414 ( .A1(n10326), .A2(keyinput166), .B1(keyinput148), .B2(n8544), .ZN(n10325) );
  OAI221_X1 U11415 ( .B1(n10326), .B2(keyinput166), .C1(n8544), .C2(
        keyinput148), .A(n10325), .ZN(n10332) );
  XNOR2_X1 U11416 ( .A(P2_IR_REG_9__SCAN_IN), .B(keyinput189), .ZN(n10330) );
  XNOR2_X1 U11417 ( .A(P2_D_REG_0__SCAN_IN), .B(keyinput155), .ZN(n10329) );
  XNOR2_X1 U11418 ( .A(P2_IR_REG_18__SCAN_IN), .B(keyinput151), .ZN(n10328) );
  XNOR2_X1 U11419 ( .A(P1_IR_REG_3__SCAN_IN), .B(keyinput173), .ZN(n10327) );
  NAND4_X1 U11420 ( .A1(n10330), .A2(n10329), .A3(n10328), .A4(n10327), .ZN(
        n10331) );
  NOR3_X1 U11421 ( .A1(n10333), .A2(n10332), .A3(n10331), .ZN(n10358) );
  INV_X1 U11422 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n10335) );
  AOI22_X1 U11423 ( .A1(n10335), .A2(keyinput232), .B1(keyinput195), .B2(n6271), .ZN(n10334) );
  OAI221_X1 U11424 ( .B1(n10335), .B2(keyinput232), .C1(n6271), .C2(
        keyinput195), .A(n10334), .ZN(n10345) );
  AOI22_X1 U11425 ( .A1(n6217), .A2(keyinput219), .B1(n10337), .B2(keyinput190), .ZN(n10336) );
  OAI221_X1 U11426 ( .B1(n6217), .B2(keyinput219), .C1(n10337), .C2(
        keyinput190), .A(n10336), .ZN(n10344) );
  AOI22_X1 U11427 ( .A1(n6329), .A2(keyinput240), .B1(keyinput192), .B2(n10339), .ZN(n10338) );
  OAI221_X1 U11428 ( .B1(n6329), .B2(keyinput240), .C1(n10339), .C2(
        keyinput192), .A(n10338), .ZN(n10343) );
  XOR2_X1 U11429 ( .A(n5355), .B(keyinput202), .Z(n10341) );
  XNOR2_X1 U11430 ( .A(P1_RD_REG_SCAN_IN), .B(keyinput138), .ZN(n10340) );
  NAND2_X1 U11431 ( .A1(n10341), .A2(n10340), .ZN(n10342) );
  NOR4_X1 U11432 ( .A1(n10345), .A2(n10344), .A3(n10343), .A4(n10342), .ZN(
        n10357) );
  INV_X1 U11433 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n10379) );
  AOI22_X1 U11434 ( .A1(n6595), .A2(keyinput176), .B1(keyinput205), .B2(n10379), .ZN(n10346) );
  OAI221_X1 U11435 ( .B1(n6595), .B2(keyinput176), .C1(n10379), .C2(
        keyinput205), .A(n10346), .ZN(n10355) );
  AOI22_X1 U11436 ( .A1(n10348), .A2(keyinput216), .B1(keyinput165), .B2(n6239), .ZN(n10347) );
  OAI221_X1 U11437 ( .B1(n10348), .B2(keyinput216), .C1(n6239), .C2(
        keyinput165), .A(n10347), .ZN(n10354) );
  AOI22_X1 U11438 ( .A1(n10430), .A2(keyinput239), .B1(keyinput234), .B2(
        n10350), .ZN(n10349) );
  OAI221_X1 U11439 ( .B1(n10430), .B2(keyinput239), .C1(n10350), .C2(
        keyinput234), .A(n10349), .ZN(n10353) );
  AOI22_X1 U11440 ( .A1(n10393), .A2(keyinput131), .B1(n6421), .B2(keyinput130), .ZN(n10351) );
  OAI221_X1 U11441 ( .B1(n10393), .B2(keyinput131), .C1(n6421), .C2(
        keyinput130), .A(n10351), .ZN(n10352) );
  NOR4_X1 U11442 ( .A1(n10355), .A2(n10354), .A3(n10353), .A4(n10352), .ZN(
        n10356) );
  NAND4_X1 U11443 ( .A1(n10359), .A2(n10358), .A3(n10357), .A4(n10356), .ZN(
        n10360) );
  NOR4_X1 U11444 ( .A1(n10363), .A2(n10362), .A3(n10361), .A4(n10360), .ZN(
        n10557) );
  AOI22_X1 U11445 ( .A1(n10365), .A2(keyinput99), .B1(keyinput19), .B2(n7325), 
        .ZN(n10364) );
  OAI221_X1 U11446 ( .B1(n10365), .B2(keyinput99), .C1(n7325), .C2(keyinput19), 
        .A(n10364), .ZN(n10377) );
  AOI22_X1 U11447 ( .A1(n10368), .A2(keyinput72), .B1(keyinput4), .B2(n10367), 
        .ZN(n10366) );
  OAI221_X1 U11448 ( .B1(n10368), .B2(keyinput72), .C1(n10367), .C2(keyinput4), 
        .A(n10366), .ZN(n10376) );
  AOI22_X1 U11449 ( .A1(n10371), .A2(keyinput108), .B1(keyinput27), .B2(n10370), .ZN(n10369) );
  OAI221_X1 U11450 ( .B1(n10371), .B2(keyinput108), .C1(n10370), .C2(
        keyinput27), .A(n10369), .ZN(n10375) );
  AOI22_X1 U11451 ( .A1(n8764), .A2(keyinput123), .B1(n10373), .B2(keyinput47), 
        .ZN(n10372) );
  OAI221_X1 U11452 ( .B1(n8764), .B2(keyinput123), .C1(n10373), .C2(keyinput47), .A(n10372), .ZN(n10374) );
  NOR4_X1 U11453 ( .A1(n10377), .A2(n10376), .A3(n10375), .A4(n10374), .ZN(
        n10425) );
  AOI22_X1 U11454 ( .A1(n6271), .A2(keyinput67), .B1(n10379), .B2(keyinput77), 
        .ZN(n10378) );
  OAI221_X1 U11455 ( .B1(n6271), .B2(keyinput67), .C1(n10379), .C2(keyinput77), 
        .A(n10378), .ZN(n10391) );
  AOI22_X1 U11456 ( .A1(n10382), .A2(keyinput70), .B1(n10381), .B2(keyinput89), 
        .ZN(n10380) );
  OAI221_X1 U11457 ( .B1(n10382), .B2(keyinput70), .C1(n10381), .C2(keyinput89), .A(n10380), .ZN(n10390) );
  AOI22_X1 U11458 ( .A1(n10385), .A2(keyinput92), .B1(keyinput90), .B2(n10384), 
        .ZN(n10383) );
  OAI221_X1 U11459 ( .B1(n10385), .B2(keyinput92), .C1(n10384), .C2(keyinput90), .A(n10383), .ZN(n10389) );
  XNOR2_X1 U11460 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(keyinput11), .ZN(n10387)
         );
  XNOR2_X1 U11461 ( .A(P1_REG1_REG_27__SCAN_IN), .B(keyinput82), .ZN(n10386)
         );
  NAND2_X1 U11462 ( .A1(n10387), .A2(n10386), .ZN(n10388) );
  NOR4_X1 U11463 ( .A1(n10391), .A2(n10390), .A3(n10389), .A4(n10388), .ZN(
        n10424) );
  AOI22_X1 U11464 ( .A1(n6161), .A2(keyinput9), .B1(keyinput3), .B2(n10393), 
        .ZN(n10392) );
  OAI221_X1 U11465 ( .B1(n6161), .B2(keyinput9), .C1(n10393), .C2(keyinput3), 
        .A(n10392), .ZN(n10405) );
  AOI22_X1 U11466 ( .A1(n10396), .A2(keyinput30), .B1(keyinput115), .B2(n10395), .ZN(n10394) );
  OAI221_X1 U11467 ( .B1(n10396), .B2(keyinput30), .C1(n10395), .C2(
        keyinput115), .A(n10394), .ZN(n10404) );
  XNOR2_X1 U11468 ( .A(n10397), .B(keyinput63), .ZN(n10403) );
  XOR2_X1 U11469 ( .A(n10398), .B(keyinput69), .Z(n10401) );
  XNOR2_X1 U11470 ( .A(P2_IR_REG_18__SCAN_IN), .B(keyinput23), .ZN(n10400) );
  XNOR2_X1 U11471 ( .A(P2_IR_REG_19__SCAN_IN), .B(keyinput52), .ZN(n10399) );
  NAND3_X1 U11472 ( .A1(n10401), .A2(n10400), .A3(n10399), .ZN(n10402) );
  NOR4_X1 U11473 ( .A1(n10405), .A2(n10404), .A3(n10403), .A4(n10402), .ZN(
        n10423) );
  AOI22_X1 U11474 ( .A1(n10408), .A2(keyinput120), .B1(n10407), .B2(
        keyinput119), .ZN(n10406) );
  OAI221_X1 U11475 ( .B1(n10408), .B2(keyinput120), .C1(n10407), .C2(
        keyinput119), .A(n10406), .ZN(n10421) );
  AOI22_X1 U11476 ( .A1(n10411), .A2(keyinput22), .B1(n10410), .B2(keyinput33), 
        .ZN(n10409) );
  OAI221_X1 U11477 ( .B1(n10411), .B2(keyinput22), .C1(n10410), .C2(keyinput33), .A(n10409), .ZN(n10420) );
  AOI22_X1 U11478 ( .A1(n10414), .A2(keyinput43), .B1(keyinput81), .B2(n10413), 
        .ZN(n10412) );
  OAI221_X1 U11479 ( .B1(n10414), .B2(keyinput43), .C1(n10413), .C2(keyinput81), .A(n10412), .ZN(n10419) );
  AOI22_X1 U11480 ( .A1(n10417), .A2(keyinput17), .B1(keyinput13), .B2(n10416), 
        .ZN(n10415) );
  OAI221_X1 U11481 ( .B1(n10417), .B2(keyinput17), .C1(n10416), .C2(keyinput13), .A(n10415), .ZN(n10418) );
  NOR4_X1 U11482 ( .A1(n10421), .A2(n10420), .A3(n10419), .A4(n10418), .ZN(
        n10422) );
  NAND4_X1 U11483 ( .A1(n10425), .A2(n10424), .A3(n10423), .A4(n10422), .ZN(
        n10556) );
  AOI22_X1 U11484 ( .A1(n10428), .A2(keyinput58), .B1(keyinput49), .B2(n10427), 
        .ZN(n10426) );
  OAI221_X1 U11485 ( .B1(n10428), .B2(keyinput58), .C1(n10427), .C2(keyinput49), .A(n10426), .ZN(n10439) );
  AOI22_X1 U11486 ( .A1(n8476), .A2(keyinput25), .B1(n10430), .B2(keyinput111), 
        .ZN(n10429) );
  OAI221_X1 U11487 ( .B1(n8476), .B2(keyinput25), .C1(n10430), .C2(keyinput111), .A(n10429), .ZN(n10438) );
  AOI22_X1 U11488 ( .A1(n10433), .A2(keyinput55), .B1(n10432), .B2(keyinput75), 
        .ZN(n10431) );
  OAI221_X1 U11489 ( .B1(n10433), .B2(keyinput55), .C1(n10432), .C2(keyinput75), .A(n10431), .ZN(n10437) );
  XNOR2_X1 U11490 ( .A(P1_IR_REG_27__SCAN_IN), .B(keyinput87), .ZN(n10435) );
  XNOR2_X1 U11491 ( .A(P2_REG3_REG_21__SCAN_IN), .B(keyinput29), .ZN(n10434)
         );
  NAND2_X1 U11492 ( .A1(n10435), .A2(n10434), .ZN(n10436) );
  NOR4_X1 U11493 ( .A1(n10439), .A2(n10438), .A3(n10437), .A4(n10436), .ZN(
        n10479) );
  AOI22_X1 U11494 ( .A1(n7706), .A2(keyinput94), .B1(n10441), .B2(keyinput26), 
        .ZN(n10440) );
  OAI221_X1 U11495 ( .B1(n7706), .B2(keyinput94), .C1(n10441), .C2(keyinput26), 
        .A(n10440), .ZN(n10452) );
  AOI22_X1 U11496 ( .A1(n10443), .A2(keyinput100), .B1(keyinput2), .B2(n6421), 
        .ZN(n10442) );
  OAI221_X1 U11497 ( .B1(n10443), .B2(keyinput100), .C1(n6421), .C2(keyinput2), 
        .A(n10442), .ZN(n10451) );
  AOI22_X1 U11498 ( .A1(n10446), .A2(keyinput39), .B1(n10445), .B2(keyinput50), 
        .ZN(n10444) );
  OAI221_X1 U11499 ( .B1(n10446), .B2(keyinput39), .C1(n10445), .C2(keyinput50), .A(n10444), .ZN(n10450) );
  AOI22_X1 U11500 ( .A1(n6228), .A2(keyinput12), .B1(n10448), .B2(keyinput103), 
        .ZN(n10447) );
  OAI221_X1 U11501 ( .B1(n6228), .B2(keyinput12), .C1(n10448), .C2(keyinput103), .A(n10447), .ZN(n10449) );
  NOR4_X1 U11502 ( .A1(n10452), .A2(n10451), .A3(n10450), .A4(n10449), .ZN(
        n10478) );
  AOI22_X1 U11503 ( .A1(n6217), .A2(keyinput91), .B1(keyinput56), .B2(n10454), 
        .ZN(n10453) );
  OAI221_X1 U11504 ( .B1(n6217), .B2(keyinput91), .C1(n10454), .C2(keyinput56), 
        .A(n10453), .ZN(n10464) );
  AOI22_X1 U11505 ( .A1(n10457), .A2(keyinput79), .B1(keyinput84), .B2(n10456), 
        .ZN(n10455) );
  OAI221_X1 U11506 ( .B1(n10457), .B2(keyinput79), .C1(n10456), .C2(keyinput84), .A(n10455), .ZN(n10463) );
  XNOR2_X1 U11507 ( .A(P1_IR_REG_0__SCAN_IN), .B(keyinput54), .ZN(n10461) );
  XNOR2_X1 U11508 ( .A(P1_REG3_REG_8__SCAN_IN), .B(keyinput105), .ZN(n10460)
         );
  XNOR2_X1 U11509 ( .A(P1_RD_REG_SCAN_IN), .B(keyinput10), .ZN(n10459) );
  XNOR2_X1 U11510 ( .A(P2_REG3_REG_22__SCAN_IN), .B(keyinput40), .ZN(n10458)
         );
  NAND4_X1 U11511 ( .A1(n10461), .A2(n10460), .A3(n10459), .A4(n10458), .ZN(
        n10462) );
  NOR3_X1 U11512 ( .A1(n10464), .A2(n10463), .A3(n10462), .ZN(n10477) );
  AOI22_X1 U11513 ( .A1(n6227), .A2(keyinput6), .B1(n10466), .B2(keyinput35), 
        .ZN(n10465) );
  OAI221_X1 U11514 ( .B1(n6227), .B2(keyinput6), .C1(n10466), .C2(keyinput35), 
        .A(n10465), .ZN(n10475) );
  XNOR2_X1 U11515 ( .A(n10467), .B(keyinput53), .ZN(n10474) );
  XNOR2_X1 U11516 ( .A(keyinput78), .B(n9453), .ZN(n10473) );
  XNOR2_X1 U11517 ( .A(P2_REG1_REG_2__SCAN_IN), .B(keyinput65), .ZN(n10471) );
  XNOR2_X1 U11518 ( .A(P1_IR_REG_25__SCAN_IN), .B(keyinput124), .ZN(n10470) );
  XNOR2_X1 U11519 ( .A(P1_REG2_REG_0__SCAN_IN), .B(keyinput109), .ZN(n10469)
         );
  XNOR2_X1 U11520 ( .A(P2_REG1_REG_23__SCAN_IN), .B(keyinput62), .ZN(n10468)
         );
  NAND4_X1 U11521 ( .A1(n10471), .A2(n10470), .A3(n10469), .A4(n10468), .ZN(
        n10472) );
  NOR4_X1 U11522 ( .A1(n10475), .A2(n10474), .A3(n10473), .A4(n10472), .ZN(
        n10476) );
  NAND4_X1 U11523 ( .A1(n10479), .A2(n10478), .A3(n10477), .A4(n10476), .ZN(
        n10555) );
  OAI22_X1 U11524 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(keyinput113), .B1(
        P2_D_REG_15__SCAN_IN), .B2(keyinput5), .ZN(n10480) );
  AOI221_X1 U11525 ( .B1(P1_IR_REG_6__SCAN_IN), .B2(keyinput113), .C1(
        keyinput5), .C2(P2_D_REG_15__SCAN_IN), .A(n10480), .ZN(n10487) );
  OAI22_X1 U11526 ( .A1(P2_REG0_REG_29__SCAN_IN), .A2(keyinput28), .B1(
        keyinput118), .B2(P1_ADDR_REG_5__SCAN_IN), .ZN(n10481) );
  AOI221_X1 U11527 ( .B1(P2_REG0_REG_29__SCAN_IN), .B2(keyinput28), .C1(
        P1_ADDR_REG_5__SCAN_IN), .C2(keyinput118), .A(n10481), .ZN(n10486) );
  OAI22_X1 U11528 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(keyinput93), .B1(keyinput1), .B2(P2_REG0_REG_18__SCAN_IN), .ZN(n10482) );
  AOI221_X1 U11529 ( .B1(P1_IR_REG_14__SCAN_IN), .B2(keyinput93), .C1(
        P2_REG0_REG_18__SCAN_IN), .C2(keyinput1), .A(n10482), .ZN(n10485) );
  OAI22_X1 U11530 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(keyinput57), .B1(keyinput8), .B2(P1_REG1_REG_3__SCAN_IN), .ZN(n10483) );
  AOI221_X1 U11531 ( .B1(P1_IR_REG_12__SCAN_IN), .B2(keyinput57), .C1(
        P1_REG1_REG_3__SCAN_IN), .C2(keyinput8), .A(n10483), .ZN(n10484) );
  NAND4_X1 U11532 ( .A1(n10487), .A2(n10486), .A3(n10485), .A4(n10484), .ZN(
        n10515) );
  OAI22_X1 U11533 ( .A1(P2_REG1_REG_22__SCAN_IN), .A2(keyinput21), .B1(
        P2_ADDR_REG_0__SCAN_IN), .B2(keyinput31), .ZN(n10488) );
  AOI221_X1 U11534 ( .B1(P2_REG1_REG_22__SCAN_IN), .B2(keyinput21), .C1(
        keyinput31), .C2(P2_ADDR_REG_0__SCAN_IN), .A(n10488), .ZN(n10495) );
  OAI22_X1 U11535 ( .A1(P2_D_REG_22__SCAN_IN), .A2(keyinput110), .B1(
        keyinput107), .B2(P2_REG1_REG_8__SCAN_IN), .ZN(n10489) );
  AOI221_X1 U11536 ( .B1(P2_D_REG_22__SCAN_IN), .B2(keyinput110), .C1(
        P2_REG1_REG_8__SCAN_IN), .C2(keyinput107), .A(n10489), .ZN(n10494) );
  OAI22_X1 U11537 ( .A1(P2_ADDR_REG_19__SCAN_IN), .A2(keyinput42), .B1(
        keyinput32), .B2(P2_REG2_REG_9__SCAN_IN), .ZN(n10490) );
  AOI221_X1 U11538 ( .B1(P2_ADDR_REG_19__SCAN_IN), .B2(keyinput42), .C1(
        P2_REG2_REG_9__SCAN_IN), .C2(keyinput32), .A(n10490), .ZN(n10493) );
  OAI22_X1 U11539 ( .A1(P2_IR_REG_24__SCAN_IN), .A2(keyinput121), .B1(SI_29_), 
        .B2(keyinput44), .ZN(n10491) );
  AOI221_X1 U11540 ( .B1(P2_IR_REG_24__SCAN_IN), .B2(keyinput121), .C1(
        keyinput44), .C2(SI_29_), .A(n10491), .ZN(n10492) );
  NAND4_X1 U11541 ( .A1(n10495), .A2(n10494), .A3(n10493), .A4(n10492), .ZN(
        n10514) );
  OAI22_X1 U11542 ( .A1(P2_REG3_REG_15__SCAN_IN), .A2(keyinput125), .B1(
        keyinput112), .B2(P2_REG2_REG_8__SCAN_IN), .ZN(n10496) );
  AOI221_X1 U11543 ( .B1(P2_REG3_REG_15__SCAN_IN), .B2(keyinput125), .C1(
        P2_REG2_REG_8__SCAN_IN), .C2(keyinput112), .A(n10496), .ZN(n10503) );
  OAI22_X1 U11544 ( .A1(P1_REG1_REG_23__SCAN_IN), .A2(keyinput34), .B1(
        P1_REG1_REG_1__SCAN_IN), .B2(keyinput85), .ZN(n10497) );
  AOI221_X1 U11545 ( .B1(P1_REG1_REG_23__SCAN_IN), .B2(keyinput34), .C1(
        keyinput85), .C2(P1_REG1_REG_1__SCAN_IN), .A(n10497), .ZN(n10502) );
  OAI22_X1 U11546 ( .A1(n6803), .A2(keyinput117), .B1(keyinput74), .B2(
        P1_IR_REG_8__SCAN_IN), .ZN(n10498) );
  AOI221_X1 U11547 ( .B1(n6803), .B2(keyinput117), .C1(P1_IR_REG_8__SCAN_IN), 
        .C2(keyinput74), .A(n10498), .ZN(n10501) );
  OAI22_X1 U11548 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(keyinput102), .B1(
        keyinput104), .B2(P2_REG3_REG_26__SCAN_IN), .ZN(n10499) );
  AOI221_X1 U11549 ( .B1(P1_REG3_REG_7__SCAN_IN), .B2(keyinput102), .C1(
        P2_REG3_REG_26__SCAN_IN), .C2(keyinput104), .A(n10499), .ZN(n10500) );
  NAND4_X1 U11550 ( .A1(n10503), .A2(n10502), .A3(n10501), .A4(n10500), .ZN(
        n10513) );
  OAI22_X1 U11551 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(keyinput80), .B1(
        P2_REG2_REG_22__SCAN_IN), .B2(keyinput20), .ZN(n10504) );
  AOI221_X1 U11552 ( .B1(P2_REG3_REG_4__SCAN_IN), .B2(keyinput80), .C1(
        keyinput20), .C2(P2_REG2_REG_22__SCAN_IN), .A(n10504), .ZN(n10511) );
  OAI22_X1 U11553 ( .A1(P1_REG3_REG_26__SCAN_IN), .A2(keyinput88), .B1(
        keyinput16), .B2(P2_REG0_REG_6__SCAN_IN), .ZN(n10505) );
  AOI221_X1 U11554 ( .B1(P1_REG3_REG_26__SCAN_IN), .B2(keyinput88), .C1(
        P2_REG0_REG_6__SCAN_IN), .C2(keyinput16), .A(n10505), .ZN(n10510) );
  OAI22_X1 U11555 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(keyinput45), .B1(keyinput86), .B2(SI_1_), .ZN(n10506) );
  AOI221_X1 U11556 ( .B1(P1_IR_REG_3__SCAN_IN), .B2(keyinput45), .C1(SI_1_), 
        .C2(keyinput86), .A(n10506), .ZN(n10509) );
  OAI22_X1 U11557 ( .A1(P2_D_REG_20__SCAN_IN), .A2(keyinput71), .B1(
        P2_D_REG_24__SCAN_IN), .B2(keyinput96), .ZN(n10507) );
  AOI221_X1 U11558 ( .B1(P2_D_REG_20__SCAN_IN), .B2(keyinput71), .C1(
        keyinput96), .C2(P2_D_REG_24__SCAN_IN), .A(n10507), .ZN(n10508) );
  NAND4_X1 U11559 ( .A1(n10511), .A2(n10510), .A3(n10509), .A4(n10508), .ZN(
        n10512) );
  NOR4_X1 U11560 ( .A1(n10515), .A2(n10514), .A3(n10513), .A4(n10512), .ZN(
        n10553) );
  OAI22_X1 U11561 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(keyinput83), .B1(
        P2_D_REG_11__SCAN_IN), .B2(keyinput38), .ZN(n10516) );
  AOI221_X1 U11562 ( .B1(P1_IR_REG_26__SCAN_IN), .B2(keyinput83), .C1(
        keyinput38), .C2(P2_D_REG_11__SCAN_IN), .A(n10516), .ZN(n10523) );
  OAI22_X1 U11563 ( .A1(P1_REG1_REG_12__SCAN_IN), .A2(keyinput76), .B1(
        P1_REG0_REG_2__SCAN_IN), .B2(keyinput97), .ZN(n10517) );
  AOI221_X1 U11564 ( .B1(P1_REG1_REG_12__SCAN_IN), .B2(keyinput76), .C1(
        keyinput97), .C2(P1_REG0_REG_2__SCAN_IN), .A(n10517), .ZN(n10522) );
  OAI22_X1 U11565 ( .A1(SI_18_), .A2(keyinput36), .B1(keyinput14), .B2(
        P2_REG3_REG_17__SCAN_IN), .ZN(n10518) );
  AOI221_X1 U11566 ( .B1(SI_18_), .B2(keyinput36), .C1(P2_REG3_REG_17__SCAN_IN), .C2(keyinput14), .A(n10518), .ZN(n10521) );
  OAI22_X1 U11567 ( .A1(P1_REG2_REG_6__SCAN_IN), .A2(keyinput98), .B1(
        P2_REG1_REG_29__SCAN_IN), .B2(keyinput41), .ZN(n10519) );
  AOI221_X1 U11568 ( .B1(P1_REG2_REG_6__SCAN_IN), .B2(keyinput98), .C1(
        keyinput41), .C2(P2_REG1_REG_29__SCAN_IN), .A(n10519), .ZN(n10520) );
  NAND4_X1 U11569 ( .A1(n10523), .A2(n10522), .A3(n10521), .A4(n10520), .ZN(
        n10551) );
  OAI22_X1 U11570 ( .A1(P2_DATAO_REG_17__SCAN_IN), .A2(keyinput46), .B1(
        P1_ADDR_REG_15__SCAN_IN), .B2(keyinput95), .ZN(n10524) );
  AOI221_X1 U11571 ( .B1(P2_DATAO_REG_17__SCAN_IN), .B2(keyinput46), .C1(
        keyinput95), .C2(P1_ADDR_REG_15__SCAN_IN), .A(n10524), .ZN(n10531) );
  OAI22_X1 U11572 ( .A1(P1_REG2_REG_19__SCAN_IN), .A2(keyinput122), .B1(
        keyinput0), .B2(P2_ADDR_REG_5__SCAN_IN), .ZN(n10525) );
  AOI221_X1 U11573 ( .B1(P1_REG2_REG_19__SCAN_IN), .B2(keyinput122), .C1(
        P2_ADDR_REG_5__SCAN_IN), .C2(keyinput0), .A(n10525), .ZN(n10530) );
  OAI22_X1 U11574 ( .A1(P1_DATAO_REG_23__SCAN_IN), .A2(keyinput59), .B1(
        keyinput127), .B2(P1_REG2_REG_29__SCAN_IN), .ZN(n10526) );
  AOI221_X1 U11575 ( .B1(P1_DATAO_REG_23__SCAN_IN), .B2(keyinput59), .C1(
        P1_REG2_REG_29__SCAN_IN), .C2(keyinput127), .A(n10526), .ZN(n10529) );
  OAI22_X1 U11576 ( .A1(P1_REG0_REG_12__SCAN_IN), .A2(keyinput68), .B1(
        keyinput64), .B2(SI_30_), .ZN(n10527) );
  AOI221_X1 U11577 ( .B1(P1_REG0_REG_12__SCAN_IN), .B2(keyinput68), .C1(SI_30_), .C2(keyinput64), .A(n10527), .ZN(n10528) );
  NAND4_X1 U11578 ( .A1(n10531), .A2(n10530), .A3(n10529), .A4(n10528), .ZN(
        n10550) );
  OAI22_X1 U11579 ( .A1(P2_IR_REG_25__SCAN_IN), .A2(keyinput48), .B1(
        keyinput116), .B2(P2_REG2_REG_23__SCAN_IN), .ZN(n10532) );
  AOI221_X1 U11580 ( .B1(P2_IR_REG_25__SCAN_IN), .B2(keyinput48), .C1(
        P2_REG2_REG_23__SCAN_IN), .C2(keyinput116), .A(n10532), .ZN(n10539) );
  OAI22_X1 U11581 ( .A1(P1_DATAO_REG_4__SCAN_IN), .A2(keyinput60), .B1(
        keyinput37), .B2(P2_REG0_REG_3__SCAN_IN), .ZN(n10533) );
  AOI221_X1 U11582 ( .B1(P1_DATAO_REG_4__SCAN_IN), .B2(keyinput60), .C1(
        P2_REG0_REG_3__SCAN_IN), .C2(keyinput37), .A(n10533), .ZN(n10538) );
  OAI22_X1 U11583 ( .A1(P1_REG0_REG_4__SCAN_IN), .A2(keyinput18), .B1(
        P1_REG0_REG_0__SCAN_IN), .B2(keyinput15), .ZN(n10534) );
  AOI221_X1 U11584 ( .B1(P1_REG0_REG_4__SCAN_IN), .B2(keyinput18), .C1(
        keyinput15), .C2(P1_REG0_REG_0__SCAN_IN), .A(n10534), .ZN(n10537) );
  OAI22_X1 U11585 ( .A1(P2_DATAO_REG_10__SCAN_IN), .A2(keyinput51), .B1(
        keyinput73), .B2(P1_REG1_REG_17__SCAN_IN), .ZN(n10535) );
  AOI221_X1 U11586 ( .B1(P2_DATAO_REG_10__SCAN_IN), .B2(keyinput51), .C1(
        P1_REG1_REG_17__SCAN_IN), .C2(keyinput73), .A(n10535), .ZN(n10536) );
  NAND4_X1 U11587 ( .A1(n10539), .A2(n10538), .A3(n10537), .A4(n10536), .ZN(
        n10549) );
  OAI22_X1 U11588 ( .A1(P1_REG2_REG_20__SCAN_IN), .A2(keyinput24), .B1(
        keyinput126), .B2(P2_ADDR_REG_11__SCAN_IN), .ZN(n10540) );
  AOI221_X1 U11589 ( .B1(P1_REG2_REG_20__SCAN_IN), .B2(keyinput24), .C1(
        P2_ADDR_REG_11__SCAN_IN), .C2(keyinput126), .A(n10540), .ZN(n10547) );
  OAI22_X1 U11590 ( .A1(P1_DATAO_REG_11__SCAN_IN), .A2(keyinput7), .B1(
        P1_REG1_REG_6__SCAN_IN), .B2(keyinput106), .ZN(n10541) );
  AOI221_X1 U11591 ( .B1(P1_DATAO_REG_11__SCAN_IN), .B2(keyinput7), .C1(
        keyinput106), .C2(P1_REG1_REG_6__SCAN_IN), .A(n10541), .ZN(n10546) );
  OAI22_X1 U11592 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(keyinput114), .B1(
        keyinput61), .B2(P2_IR_REG_9__SCAN_IN), .ZN(n10542) );
  AOI221_X1 U11593 ( .B1(P1_IR_REG_17__SCAN_IN), .B2(keyinput114), .C1(
        P2_IR_REG_9__SCAN_IN), .C2(keyinput61), .A(n10542), .ZN(n10545) );
  OAI22_X1 U11594 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(keyinput101), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(keyinput66), .ZN(n10543) );
  AOI221_X1 U11595 ( .B1(P1_DATAO_REG_20__SCAN_IN), .B2(keyinput101), .C1(
        keyinput66), .C2(P2_DATAO_REG_18__SCAN_IN), .A(n10543), .ZN(n10544) );
  NAND4_X1 U11596 ( .A1(n10547), .A2(n10546), .A3(n10545), .A4(n10544), .ZN(
        n10548) );
  NOR4_X1 U11597 ( .A1(n10551), .A2(n10550), .A3(n10549), .A4(n10548), .ZN(
        n10552) );
  NAND2_X1 U11598 ( .A1(n10553), .A2(n10552), .ZN(n10554) );
  NOR4_X1 U11599 ( .A1(n10557), .A2(n10556), .A3(n10555), .A4(n10554), .ZN(
        n10574) );
  OAI211_X1 U11600 ( .C1(n10561), .C2(n10560), .A(n10559), .B(n10558), .ZN(
        n10572) );
  OAI211_X1 U11601 ( .C1(n10565), .C2(n10564), .A(n10563), .B(n10562), .ZN(
        n10571) );
  AOI22_X1 U11602 ( .A1(n10566), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n10570) );
  NAND2_X1 U11603 ( .A1(n10568), .A2(n10567), .ZN(n10569) );
  NAND4_X1 U11604 ( .A1(n10572), .A2(n10571), .A3(n10570), .A4(n10569), .ZN(
        n10573) );
  XOR2_X1 U11605 ( .A(n10574), .B(n10573), .Z(P1_U3244) );
  OAI21_X1 U11606 ( .B1(n10577), .B2(n10576), .A(n10575), .ZN(ADD_1068_U50) );
  OAI21_X1 U11607 ( .B1(n10580), .B2(n10579), .A(n10578), .ZN(ADD_1068_U51) );
  OAI21_X1 U11608 ( .B1(n10583), .B2(n10582), .A(n10581), .ZN(ADD_1068_U49) );
  OAI21_X1 U11609 ( .B1(n10586), .B2(n10585), .A(n10584), .ZN(ADD_1068_U47) );
  OAI21_X1 U11610 ( .B1(n10589), .B2(n10588), .A(n10587), .ZN(ADD_1068_U48) );
  AOI21_X1 U11611 ( .B1(n10592), .B2(n10591), .A(n10590), .ZN(ADD_1068_U54) );
  AOI21_X1 U11612 ( .B1(n10595), .B2(n10594), .A(n10593), .ZN(ADD_1068_U53) );
  OAI21_X1 U11613 ( .B1(n10598), .B2(n10597), .A(n10596), .ZN(ADD_1068_U52) );
  CLKBUF_X1 U5041 ( .A(n5336), .Z(n6712) );
  AND3_X1 U6425 ( .A1(n6232), .A2(n6231), .A3(n6230), .ZN(n5135) );
  OR2_X1 U7744 ( .A1(n6186), .A2(n6246), .ZN(n6188) );
  INV_X2 U8458 ( .A(n8450), .ZN(n8779) );
endmodule

