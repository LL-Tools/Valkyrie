

module b15_C_2inp_gates_syn ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, 
        READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, 
        CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, 
        REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, 
        FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, U3445, U3446, U3447, U3448, 
        U3213, U3212, U3211, U3210, U3209, U3208, U3207, U3206, U3205, U3204, 
        U3203, U3202, U3201, U3200, U3199, U3198, U3197, U3196, U3195, U3194, 
        U3193, U3192, U3191, U3190, U3189, U3188, U3187, U3186, U3185, U3184, 
        U3183, U3182, U3181, U3451, U3452, U3180, U3179, U3178, U3177, U3176, 
        U3175, U3174, U3173, U3172, U3171, U3170, U3169, U3168, U3167, U3166, 
        U3165, U3164, U3163, U3162, U3161, U3160, U3159, U3158, U3157, U3156, 
        U3155, U3154, U3153, U3152, U3151, U3453, U3150, U3149, U3148, U3147, 
        U3146, U3145, U3144, U3143, U3142, U3141, U3140, U3139, U3138, U3137, 
        U3136, U3135, U3134, U3133, U3132, U3131, U3130, U3129, U3128, U3127, 
        U3126, U3125, U3124, U3123, U3122, U3121, U3120, U3119, U3118, U3117, 
        U3116, U3115, U3114, U3113, U3112, U3111, U3110, U3109, U3108, U3107, 
        U3106, U3105, U3104, U3103, U3102, U3101, U3100, U3099, U3098, U3097, 
        U3096, U3095, U3094, U3093, U3092, U3091, U3090, U3089, U3088, U3087, 
        U3086, U3085, U3084, U3083, U3082, U3081, U3080, U3079, U3078, U3077, 
        U3076, U3075, U3074, U3073, U3072, U3071, U3070, U3069, U3068, U3067, 
        U3066, U3065, U3064, U3063, U3062, U3061, U3060, U3059, U3058, U3057, 
        U3056, U3055, U3054, U3053, U3052, U3051, U3050, U3049, U3048, U3047, 
        U3046, U3045, U3044, U3043, U3042, U3041, U3040, U3039, U3038, U3037, 
        U3036, U3035, U3034, U3033, U3032, U3031, U3030, U3029, U3028, U3027, 
        U3026, U3025, U3024, U3023, U3022, U3021, U3020, U3455, U3456, U3459, 
        U3460, U3461, U3019, U3462, U3463, U3464, U3465, U3018, U3017, U3016, 
        U3015, U3014, U3013, U3012, U3011, U3010, U3009, U3008, U3007, U3006, 
        U3005, U3004, U3003, U3002, U3001, U3000, U2999, U2998, U2997, U2996, 
        U2995, U2994, U2993, U2992, U2991, U2990, U2989, U2988, U2987, U2986, 
        U2985, U2984, U2983, U2982, U2981, U2980, U2979, U2978, U2977, U2976, 
        U2975, U2974, U2973, U2972, U2971, U2970, U2969, U2968, U2967, U2966, 
        U2965, U2964, U2963, U2962, U2961, U2960, U2959, U2958, U2957, U2956, 
        U2955, U2954, U2953, U2952, U2951, U2950, U2949, U2948, U2947, U2946, 
        U2945, U2944, U2943, U2942, U2941, U2940, U2939, U2938, U2937, U2936, 
        U2935, U2934, U2933, U2932, U2931, U2930, U2929, U2928, U2927, U2926, 
        U2925, U2924, U2923, U2922, U2921, U2920, U2919, U2918, U2917, U2916, 
        U2915, U2914, U2913, U2912, U2911, U2910, U2909, U2908, U2907, U2906, 
        U2905, U2904, U2903, U2902, U2901, U2900, U2899, U2898, U2897, U2896, 
        U2895, U2894, U2893, U2892, U2891, U2890, U2889, U2888, U2887, U2886, 
        U2885, U2884, U2883, U2882, U2881, U2880, U2879, U2878, U2877, U2876, 
        U2875, U2874, U2873, U2872, U2871, U2870, U2869, U2868, U2867, U2866, 
        U2865, U2864, U2863, U2862, U2861, U2860, U2859, U2858, U2857, U2856, 
        U2855, U2854, U2853, U2852, U2851, U2850, U2849, U2848, U2847, U2846, 
        U2845, U2844, U2843, U2842, U2841, U2840, U2839, U2838, U2837, U2836, 
        U2835, U2834, U2833, U2832, U2831, U2830, U2829, U2828, U2827, U2826, 
        U2825, U2824, U2823, U2822, U2821, U2820, U2819, U2818, U2817, U2816, 
        U2815, U2814, U2813, U2812, U2811, U2810, U2809, U2808, U2807, U2806, 
        U2805, U2804, U2803, U2802, U2801, U2800, U2799, U2798, U2797, U2796, 
        U2795, U3468, U2794, U3469, U3470, U2793, U3471, U2792, U3472, U2791, 
        U3473, U2790, U2789, U3474, U2788, keyinput63, keyinput62, keyinput61, 
        keyinput60, keyinput59, keyinput58, keyinput57, keyinput56, keyinput55, 
        keyinput54, keyinput53, keyinput52, keyinput51, keyinput50, keyinput49, 
        keyinput48, keyinput47, keyinput46, keyinput45, keyinput44, keyinput43, 
        keyinput42, keyinput41, keyinput40, keyinput39, keyinput38, keyinput37, 
        keyinput36, keyinput35, keyinput34, keyinput33, keyinput32, keyinput31, 
        keyinput30, keyinput29, keyinput28, keyinput27, keyinput26, keyinput25, 
        keyinput24, keyinput23, keyinput22, keyinput21, keyinput20, keyinput19, 
        keyinput18, keyinput17, keyinput16, keyinput15, keyinput14, keyinput13, 
        keyinput12, keyinput11, keyinput10, keyinput9, keyinput8, keyinput7, 
        keyinput6, keyinput5, keyinput4, keyinput3, keyinput2, keyinput1, 
        keyinput0 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
         READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
         M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
         STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
         W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput63, keyinput62,
         keyinput61, keyinput60, keyinput59, keyinput58, keyinput57,
         keyinput56, keyinput55, keyinput54, keyinput53, keyinput52,
         keyinput51, keyinput50, keyinput49, keyinput48, keyinput47,
         keyinput46, keyinput45, keyinput44, keyinput43, keyinput42,
         keyinput41, keyinput40, keyinput39, keyinput38, keyinput37,
         keyinput36, keyinput35, keyinput34, keyinput33, keyinput32,
         keyinput31, keyinput30, keyinput29, keyinput28, keyinput27,
         keyinput26, keyinput25, keyinput24, keyinput23, keyinput22,
         keyinput21, keyinput20, keyinput19, keyinput18, keyinput17,
         keyinput16, keyinput15, keyinput14, keyinput13, keyinput12,
         keyinput11, keyinput10, keyinput9, keyinput8, keyinput7, keyinput6,
         keyinput5, keyinput4, keyinput3, keyinput2, keyinput1, keyinput0;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971,
         n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981,
         n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991,
         n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001,
         n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011,
         n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021,
         n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031,
         n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041,
         n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051,
         n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061,
         n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071,
         n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081,
         n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091,
         n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101,
         n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111,
         n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121,
         n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131,
         n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141,
         n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151,
         n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161,
         n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171,
         n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181,
         n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191,
         n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201,
         n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211,
         n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221,
         n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231,
         n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241,
         n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251,
         n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261,
         n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271,
         n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281,
         n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291,
         n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301,
         n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311,
         n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321,
         n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331,
         n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341,
         n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351,
         n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361,
         n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371,
         n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381,
         n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391,
         n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401,
         n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411,
         n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421,
         n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431,
         n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441,
         n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451,
         n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461,
         n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471,
         n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481,
         n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491,
         n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501,
         n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511,
         n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521,
         n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531,
         n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541,
         n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551,
         n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561,
         n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571,
         n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581,
         n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591,
         n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601,
         n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611,
         n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621,
         n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631,
         n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641,
         n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651,
         n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661,
         n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671,
         n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681,
         n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691,
         n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701,
         n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711,
         n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721,
         n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731,
         n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741,
         n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751,
         n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761,
         n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771,
         n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781,
         n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791,
         n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801,
         n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811,
         n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821,
         n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831,
         n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841,
         n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851,
         n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861,
         n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871,
         n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881,
         n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891,
         n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901,
         n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911,
         n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921,
         n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931,
         n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941,
         n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951,
         n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961,
         n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971,
         n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981,
         n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991,
         n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001,
         n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011,
         n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021,
         n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031,
         n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041,
         n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051,
         n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061,
         n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071,
         n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081,
         n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091,
         n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101,
         n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111,
         n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121,
         n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131,
         n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141,
         n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151,
         n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161,
         n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171,
         n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181,
         n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191,
         n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201,
         n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4210, n4211, n4213,
         n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223,
         n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233,
         n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243,
         n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253,
         n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263,
         n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273,
         n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283,
         n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293,
         n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303,
         n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313,
         n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323,
         n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333,
         n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343,
         n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353,
         n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363,
         n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373,
         n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383,
         n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393,
         n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403,
         n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413,
         n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423,
         n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433,
         n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443,
         n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453,
         n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463,
         n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473,
         n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483,
         n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493,
         n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503,
         n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513,
         n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523,
         n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533,
         n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543,
         n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553,
         n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563,
         n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573,
         n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583,
         n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593,
         n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603,
         n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613,
         n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623,
         n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633,
         n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643,
         n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653,
         n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663,
         n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673,
         n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683,
         n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693,
         n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703,
         n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713,
         n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723,
         n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733,
         n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743,
         n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753,
         n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763,
         n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773,
         n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783,
         n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793,
         n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803,
         n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813,
         n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823,
         n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833,
         n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843,
         n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853,
         n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863,
         n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873,
         n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883,
         n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893,
         n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903,
         n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913,
         n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923,
         n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933,
         n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943,
         n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953,
         n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963,
         n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973,
         n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983,
         n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993,
         n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003,
         n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013,
         n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023,
         n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033,
         n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043,
         n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053,
         n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063,
         n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073,
         n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083,
         n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093,
         n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103,
         n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113,
         n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123,
         n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133,
         n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143,
         n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153,
         n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163,
         n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173,
         n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183,
         n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193,
         n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203,
         n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213,
         n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223,
         n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233,
         n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243,
         n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253,
         n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263,
         n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273,
         n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283,
         n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293,
         n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303,
         n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313,
         n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323,
         n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333,
         n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343,
         n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353,
         n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363,
         n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373,
         n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383,
         n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393,
         n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403,
         n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413,
         n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423,
         n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433,
         n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443,
         n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453,
         n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463,
         n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473,
         n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483,
         n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493,
         n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503,
         n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513,
         n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523,
         n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533,
         n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543,
         n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553,
         n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563,
         n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573,
         n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583,
         n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593,
         n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603,
         n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613,
         n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623,
         n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633,
         n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643,
         n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653,
         n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663,
         n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673,
         n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683,
         n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693,
         n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703,
         n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713,
         n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723,
         n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733,
         n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743,
         n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753,
         n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763,
         n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773,
         n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783,
         n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793,
         n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803,
         n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813,
         n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823,
         n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833,
         n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843,
         n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853,
         n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863,
         n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873,
         n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883,
         n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893,
         n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903,
         n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913,
         n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923,
         n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933,
         n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943,
         n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953,
         n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963,
         n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973,
         n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983,
         n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993,
         n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003,
         n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013,
         n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023,
         n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033,
         n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043,
         n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053,
         n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063,
         n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073,
         n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083,
         n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093,
         n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103,
         n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113,
         n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123,
         n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133,
         n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143,
         n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153,
         n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163,
         n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173,
         n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183,
         n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193,
         n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203,
         n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213,
         n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223,
         n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233,
         n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243,
         n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253,
         n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263,
         n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273,
         n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283,
         n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293,
         n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303,
         n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313,
         n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323,
         n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333,
         n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343,
         n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353,
         n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363,
         n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373,
         n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383,
         n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393,
         n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403,
         n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413,
         n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423,
         n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433,
         n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443,
         n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453,
         n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463,
         n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473,
         n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483,
         n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493,
         n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503,
         n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513,
         n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523,
         n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533,
         n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543,
         n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553,
         n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563,
         n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573,
         n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583,
         n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593,
         n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603,
         n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613,
         n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623,
         n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633,
         n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643,
         n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653,
         n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663,
         n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673,
         n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683,
         n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693,
         n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703,
         n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713,
         n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723,
         n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733,
         n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743,
         n6744;

  AND2_X1 U3410 ( .A1(n5319), .A2(n3626), .ZN(n3641) );
  OAI21_X1 U3411 ( .B1(n5785), .B2(STATE2_REG_0__SCAN_IN), .A(n3214), .ZN(
        n3344) );
  CLKBUF_X2 U3412 ( .A(n4151), .Z(n4224) );
  CLKBUF_X2 U3413 ( .A(n3224), .Z(n3232) );
  NAND4_X2 U3415 ( .A1(n3102), .A2(n3101), .A3(n3100), .A4(n3099), .ZN(n3518)
         );
  AND2_X1 U3416 ( .A1(n2988), .A2(n2986), .ZN(n3218) );
  CLKBUF_X1 U3417 ( .A(n3266), .Z(n2962) );
  AND2_X1 U3418 ( .A1(n4381), .A2(n2992), .ZN(n3266) );
  CLKBUF_X2 U3420 ( .A(n3081), .Z(n4211) );
  OR2_X1 U3421 ( .A1(n3148), .A2(n3518), .ZN(n3652) );
  NAND2_X1 U3422 ( .A1(n4473), .A2(n3511), .ZN(n3642) );
  OR2_X1 U3423 ( .A1(n4332), .A2(n5249), .ZN(n3638) );
  NAND2_X1 U3424 ( .A1(n3292), .A2(n3291), .ZN(n4624) );
  AND4_X2 U3426 ( .A1(n3047), .A2(n3046), .A3(n3045), .A4(n3044), .ZN(n3231)
         );
  NAND2_X1 U3427 ( .A1(n3518), .A2(n3517), .ZN(n3539) );
  OR2_X1 U3428 ( .A1(n4977), .A2(n3767), .ZN(n3768) );
  NAND2_X1 U3429 ( .A1(n3389), .A2(n3388), .ZN(n3749) );
  XNOR2_X1 U3430 ( .A(n4624), .B(n4623), .ZN(n4505) );
  NAND2_X1 U3431 ( .A1(n3358), .A2(n3357), .ZN(n3715) );
  NAND2_X1 U3433 ( .A1(n5392), .A2(n3631), .ZN(n4255) );
  CLKBUF_X2 U3434 ( .A(n3539), .Z(n2964) );
  AOI21_X1 U3435 ( .B1(n3749), .B2(n2965), .A(n3748), .ZN(n4977) );
  AND2_X2 U3437 ( .A1(n3509), .A2(n3518), .ZN(n4294) );
  INV_X1 U3438 ( .A(n5995), .ZN(n6698) );
  NAND2_X1 U3439 ( .A1(n5314), .A2(n5313), .ZN(n5465) );
  INV_X1 U3440 ( .A(n6077), .ZN(n6702) );
  BUF_X1 U3441 ( .A(n3015), .Z(n4225) );
  AOI21_X4 U3443 ( .B1(n5659), .B2(n6160), .A(n3437), .ZN(n5520) );
  NAND2_X1 U3444 ( .A1(n5348), .A2(n5347), .ZN(n5349) );
  NOR3_X1 U34450 ( .A1(n3438), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .A3(n5346), .ZN(n3439) );
  CLKBUF_X1 U34460 ( .A(n5501), .Z(n5513) );
  NAND2_X1 U34470 ( .A1(n5443), .A2(n5442), .ZN(n5388) );
  NOR2_X2 U34480 ( .A1(n5401), .A2(n5402), .ZN(n5443) );
  NAND2_X1 U3449 ( .A1(n4103), .A2(n4102), .ZN(n5401) );
  INV_X1 U3450 ( .A(n5453), .ZN(n4103) );
  NAND2_X1 U34510 ( .A1(n5553), .A2(n5454), .ZN(n5453) );
  NAND2_X1 U34520 ( .A1(n4255), .A2(n5319), .ZN(n4256) );
  INV_X2 U34530 ( .A(n2967), .ZN(n2963) );
  XNOR2_X1 U3454 ( .A(n3367), .B(n3375), .ZN(n3723) );
  AOI21_X1 U34550 ( .B1(n4505), .B2(n6443), .A(n3311), .ZN(n3365) );
  CLKBUF_X1 U34560 ( .A(n4417), .Z(n5783) );
  NAND2_X1 U3457 ( .A1(n3198), .A2(n3197), .ZN(n3200) );
  XNOR2_X1 U3458 ( .A(n3345), .B(n3344), .ZN(n4417) );
  NAND2_X2 U34590 ( .A1(n5472), .A2(n4405), .ZN(n5914) );
  AND2_X1 U34600 ( .A1(n3344), .A2(n3258), .ZN(n3327) );
  INV_X1 U34610 ( .A(n3290), .ZN(n3292) );
  XNOR2_X1 U34620 ( .A(n3343), .B(n3342), .ZN(n3345) );
  NAND2_X1 U34630 ( .A1(n3564), .A2(n3563), .ZN(n5190) );
  OAI21_X1 U34640 ( .B1(n4837), .B2(n3465), .A(n3338), .ZN(n4349) );
  NAND2_X1 U34650 ( .A1(n3252), .A2(n3325), .ZN(n3343) );
  INV_X2 U3466 ( .A(n4429), .ZN(n4572) );
  NAND2_X1 U3467 ( .A1(n3215), .A2(n3217), .ZN(n3202) );
  OR2_X1 U34680 ( .A1(n3173), .A2(n3172), .ZN(n3215) );
  CLKBUF_X1 U34690 ( .A(n3516), .Z(n4336) );
  CLKBUF_X1 U34700 ( .A(n3490), .Z(n4299) );
  INV_X1 U34710 ( .A(n3551), .ZN(n3622) );
  CLKBUF_X1 U34720 ( .A(n3551), .Z(n3625) );
  BUF_X2 U34730 ( .A(n3537), .Z(n3626) );
  NAND2_X2 U3475 ( .A1(n3133), .A2(n3123), .ZN(n3126) );
  INV_X1 U3476 ( .A(n3511), .ZN(n3124) );
  OR2_X1 U3477 ( .A1(n3230), .A2(n3229), .ZN(n3410) );
  CLKBUF_X1 U3478 ( .A(n3123), .Z(n4477) );
  NAND4_X2 U3479 ( .A1(n3013), .A2(n3012), .A3(n3011), .A4(n3010), .ZN(n3141)
         );
  OR2_X1 U3480 ( .A1(n3242), .A2(n3241), .ZN(n3346) );
  OR2_X2 U3481 ( .A1(n3025), .A2(n3024), .ZN(n3146) );
  AND4_X1 U3482 ( .A1(n3029), .A2(n3028), .A3(n3027), .A4(n3026), .ZN(n3047)
         );
  AND4_X1 U3483 ( .A1(n3038), .A2(n3037), .A3(n3036), .A4(n3035), .ZN(n3045)
         );
  AND4_X1 U3484 ( .A1(n3076), .A2(n3075), .A3(n3074), .A4(n3073), .ZN(n3077)
         );
  AND4_X1 U3485 ( .A1(n2997), .A2(n2996), .A3(n2995), .A4(n2994), .ZN(n3013)
         );
  AND4_X1 U3486 ( .A1(n3009), .A2(n3008), .A3(n3007), .A4(n3006), .ZN(n3010)
         );
  AND4_X1 U3487 ( .A1(n3106), .A2(n3105), .A3(n3104), .A4(n3103), .ZN(n3122)
         );
  AND4_X1 U3488 ( .A1(n3034), .A2(n3033), .A3(n3032), .A4(n3031), .ZN(n3046)
         );
  AND4_X1 U3489 ( .A1(n3072), .A2(n3071), .A3(n3070), .A4(n3069), .ZN(n3078)
         );
  BUF_X2 U3490 ( .A(n3189), .Z(n4219) );
  BUF_X2 U3491 ( .A(n4210), .Z(n4173) );
  BUF_X2 U3493 ( .A(n3218), .Z(n4214) );
  INV_X2 U3494 ( .A(n6248), .ZN(n3668) );
  CLKBUF_X1 U3495 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .Z(n4607) );
  AOI211_X2 U3496 ( .C1(n3667), .C2(n6280), .A(n5339), .B(n3666), .ZN(n3683)
         );
  XNOR2_X2 U3497 ( .A(n3363), .B(n6272), .ZN(n4726) );
  OAI22_X2 U3498 ( .A1(n3715), .A2(n3465), .B1(n6559), .B2(n3362), .ZN(n3363)
         );
  NOR2_X2 U3499 ( .A1(n4661), .A2(n4924), .ZN(n4921) );
  AND2_X4 U3500 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n2986) );
  NAND2_X1 U3501 ( .A1(n3328), .A2(n3327), .ZN(n3366) );
  AND2_X2 U3502 ( .A1(n5261), .A2(n4409), .ZN(n3551) );
  NAND2_X1 U3503 ( .A1(n3155), .A2(n3154), .ZN(n3649) );
  NAND2_X1 U3504 ( .A1(n5520), .A2(n5519), .ZN(n5501) );
  NAND2_X1 U3505 ( .A1(n4199), .A2(n4200), .ZN(n5334) );
  NAND2_X1 U3506 ( .A1(n4320), .A2(n6440), .ZN(n4308) );
  CLKBUF_X1 U3507 ( .A(n3060), .Z(n4078) );
  AND2_X1 U3508 ( .A1(n3140), .A2(n3146), .ZN(n3646) );
  OR2_X1 U3509 ( .A1(n3139), .A2(n4486), .ZN(n3140) );
  CLKBUF_X1 U3510 ( .A(n3177), .Z(n3178) );
  NOR2_X2 U3511 ( .A1(n5937), .A2(n5247), .ZN(n5246) );
  INV_X1 U3512 ( .A(n3704), .ZN(n4237) );
  OR2_X1 U3513 ( .A1(n3424), .A2(n2970), .ZN(n5576) );
  OR2_X1 U3514 ( .A1(n5624), .A2(n3423), .ZN(n3424) );
  AND2_X1 U3515 ( .A1(n5603), .A2(n2971), .ZN(n5577) );
  AND2_X1 U3516 ( .A1(n6158), .A2(n3419), .ZN(n3420) );
  NAND2_X1 U3517 ( .A1(n2967), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n3419) );
  NAND2_X1 U3518 ( .A1(n3622), .A2(n3534), .ZN(n3536) );
  NAND2_X1 U3519 ( .A1(n2975), .A2(n3166), .ZN(n3887) );
  NAND2_X1 U3520 ( .A1(n3299), .A2(n3298), .ZN(n4623) );
  AND4_X1 U3521 ( .A1(n3089), .A2(n3088), .A3(n3087), .A4(n3086), .ZN(n3101)
         );
  AND4_X1 U3522 ( .A1(n3110), .A2(n3109), .A3(n3108), .A4(n3107), .ZN(n3121)
         );
  AND2_X1 U3523 ( .A1(n6074), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5207) );
  INV_X1 U3524 ( .A(n4008), .ZN(n4009) );
  NAND2_X1 U3525 ( .A1(n5528), .A2(n5518), .ZN(n5512) );
  OAI21_X1 U3526 ( .B1(n5570), .B2(n2979), .A(n2967), .ZN(n3435) );
  BUF_X1 U3527 ( .A(n3437), .Z(n5528) );
  NOR2_X2 U3528 ( .A1(n5051), .A2(n5034), .ZN(n5064) );
  NOR2_X2 U3529 ( .A1(n5197), .A2(n5038), .ZN(n5059) );
  NOR2_X2 U3530 ( .A1(n4449), .A2(n3543), .ZN(n4577) );
  NAND2_X1 U3531 ( .A1(n3489), .A2(n3488), .ZN(n4320) );
  OR2_X1 U3532 ( .A1(n3487), .A2(n3486), .ZN(n3488) );
  BUF_X1 U3534 ( .A(n4505), .Z(n6059) );
  AND2_X1 U3535 ( .A1(n5472), .A2(n5250), .ZN(n6104) );
  INV_X1 U3536 ( .A(n5472), .ZN(n6103) );
  OR2_X1 U3537 ( .A1(n5390), .A2(n4200), .ZN(n4201) );
  XNOR2_X1 U3538 ( .A(n4027), .B(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5332)
         );
  NAND2_X1 U3539 ( .A1(n4026), .A2(n4025), .ZN(n4027) );
  OR2_X1 U3540 ( .A1(n4467), .A2(n6443), .ZN(n3260) );
  INV_X1 U3541 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n2980) );
  CLKBUF_X1 U3542 ( .A(n3223), .Z(n4221) );
  CLKBUF_X1 U3543 ( .A(n3266), .Z(n3888) );
  CLKBUF_X1 U3544 ( .A(n4112), .Z(n3961) );
  CLKBUF_X1 U3545 ( .A(n4176), .Z(n4213) );
  OR2_X1 U3546 ( .A1(n5576), .A2(n5597), .ZN(n3425) );
  OR2_X1 U3547 ( .A1(n4486), .A2(n6443), .ZN(n3259) );
  INV_X1 U3548 ( .A(n3475), .ZN(n3460) );
  OR2_X1 U3549 ( .A1(n3213), .A2(n3212), .ZN(n3347) );
  NOR2_X1 U3550 ( .A1(n3366), .A2(n3365), .ZN(n3376) );
  NAND2_X1 U3551 ( .A1(n3260), .A2(n3259), .ZN(n3483) );
  AND2_X1 U3552 ( .A1(n3132), .A2(n3153), .ZN(n3490) );
  NOR2_X1 U3553 ( .A1(n3151), .A2(n3652), .ZN(n3132) );
  NOR2_X2 U3554 ( .A1(n5388), .A2(n5391), .ZN(n4199) );
  NAND2_X1 U3555 ( .A1(n3853), .A2(n3852), .ZN(n4661) );
  INV_X1 U3556 ( .A(n4664), .ZN(n3852) );
  INV_X1 U3557 ( .A(n4662), .ZN(n3853) );
  NOR2_X1 U3558 ( .A1(n3717), .A2(n4728), .ZN(n3727) );
  OR2_X1 U3559 ( .A1(n3196), .A2(n3195), .ZN(n3359) );
  NOR2_X1 U3560 ( .A1(n2978), .A2(n3630), .ZN(n3631) );
  NOR2_X1 U3561 ( .A1(n5529), .A2(n5530), .ZN(n3437) );
  INV_X1 U3562 ( .A(n3632), .ZN(n3602) );
  OR2_X1 U3563 ( .A1(n4337), .A2(n3656), .ZN(n3658) );
  NAND2_X1 U3564 ( .A1(n4577), .A2(n4576), .ZN(n4575) );
  INV_X1 U3565 ( .A(n3642), .ZN(n3492) );
  AND2_X1 U3566 ( .A1(n4481), .A2(n4494), .ZN(n3441) );
  INV_X1 U3567 ( .A(n3148), .ZN(n3520) );
  OR2_X1 U3568 ( .A1(n3328), .A2(n3327), .ZN(n3329) );
  INV_X1 U3569 ( .A(n3215), .ZN(n3216) );
  NOR2_X2 U3570 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n2987) );
  AND2_X1 U3571 ( .A1(n3482), .A2(n3481), .ZN(n3504) );
  NAND2_X1 U3572 ( .A1(n3475), .A2(n3441), .ZN(n3487) );
  NAND2_X1 U3573 ( .A1(n3490), .A2(n3509), .ZN(n3516) );
  INV_X1 U3574 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6612) );
  INV_X1 U3575 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4830) );
  AND4_X1 U3576 ( .A1(n3043), .A2(n3042), .A3(n3041), .A4(n3040), .ZN(n3044)
         );
  AND4_X1 U3577 ( .A1(n3068), .A2(n3067), .A3(n3066), .A4(n3065), .ZN(n3079)
         );
  CLKBUF_X1 U3578 ( .A(n4457), .Z(n4652) );
  AND2_X1 U3579 ( .A1(n4060), .A2(n4059), .ZN(n5551) );
  AND2_X1 U3580 ( .A1(n5317), .A2(n3599), .ZN(n5468) );
  AND2_X2 U3581 ( .A1(n4061), .A2(n5551), .ZN(n5553) );
  NOR2_X1 U3583 ( .A1(n4142), .A2(n5524), .ZN(n4143) );
  NAND2_X1 U3584 ( .A1(n4143), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n4191)
         );
  CLKBUF_X1 U3585 ( .A(n5388), .Z(n5389) );
  OR2_X1 U3586 ( .A1(n4095), .A2(n5541), .ZN(n4097) );
  OR2_X1 U3587 ( .A1(n4097), .A2(n4096), .ZN(n4142) );
  BUF_X1 U3588 ( .A(n5401), .Z(n5411) );
  NOR2_X1 U3589 ( .A1(n4056), .A2(n4055), .ZN(n4057) );
  NAND2_X1 U3590 ( .A1(n4057), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n4095)
         );
  OR2_X1 U3591 ( .A1(n3988), .A2(n3987), .ZN(n4056) );
  CLKBUF_X1 U3592 ( .A(n4010), .Z(n3992) );
  INV_X1 U3593 ( .A(n5303), .ZN(n3956) );
  NAND2_X1 U3594 ( .A1(PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n3918), .ZN(n3950)
         );
  CLKBUF_X1 U3595 ( .A(n5066), .Z(n5067) );
  NOR2_X1 U3596 ( .A1(n3884), .A2(n6723), .ZN(n3918) );
  NAND2_X1 U3597 ( .A1(n3869), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n3883)
         );
  CLKBUF_X1 U3598 ( .A(n4921), .Z(n4922) );
  OR2_X1 U3599 ( .A1(n3837), .A2(n5437), .ZN(n3854) );
  NAND2_X1 U3600 ( .A1(n3788), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3837)
         );
  CLKBUF_X1 U3601 ( .A(n4662), .Z(n4663) );
  AND2_X1 U3602 ( .A1(n3802), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3788)
         );
  NOR2_X1 U3603 ( .A1(n3751), .A2(n6567), .ZN(n3802) );
  AND2_X1 U3604 ( .A1(n3750), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3827)
         );
  NAND2_X1 U3605 ( .A1(n3769), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3743)
         );
  INV_X1 U3606 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3742) );
  OR2_X1 U3607 ( .A1(n4968), .A2(n4967), .ZN(n5426) );
  CLKBUF_X1 U3608 ( .A(n4471), .Z(n4968) );
  NAND2_X1 U3609 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3717) );
  OR2_X1 U3610 ( .A1(n6542), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4013) );
  BUF_X1 U3612 ( .A(n5461), .Z(n5679) );
  NAND2_X1 U3613 ( .A1(n3687), .A2(n3686), .ZN(n5558) );
  OR2_X1 U3614 ( .A1(n6160), .A2(n3685), .ZN(n3686) );
  NOR2_X2 U3615 ( .A1(n5944), .A2(n5307), .ZN(n5317) );
  OR2_X1 U3616 ( .A1(n6160), .A2(n3431), .ZN(n3432) );
  CLKBUF_X1 U3617 ( .A(n5574), .Z(n5931) );
  XNOR2_X1 U3619 ( .A(n6160), .B(n5744), .ZN(n5597) );
  AND2_X1 U3620 ( .A1(n5578), .A2(n5577), .ZN(n5596) );
  AND2_X1 U3621 ( .A1(n5625), .A2(n3426), .ZN(n5603) );
  OR2_X1 U3622 ( .A1(n3422), .A2(n5616), .ZN(n5604) );
  NAND2_X1 U3623 ( .A1(n3578), .A2(n3577), .ZN(n5049) );
  INV_X1 U3624 ( .A(n4666), .ZN(n3578) );
  CLKBUF_X1 U3625 ( .A(n5575), .Z(n5628) );
  AND3_X1 U3626 ( .A1(n3566), .A2(n3607), .A3(n3565), .ZN(n5189) );
  OR2_X1 U3627 ( .A1(n2963), .A2(n3418), .ZN(n6158) );
  INV_X1 U3628 ( .A(n5061), .ZN(n3564) );
  NAND2_X1 U3629 ( .A1(n3550), .A2(n3549), .ZN(n5195) );
  INV_X1 U3630 ( .A(n4716), .ZN(n3549) );
  INV_X1 U3631 ( .A(n4575), .ZN(n3550) );
  AND2_X1 U3632 ( .A1(n3555), .A2(n3554), .ZN(n5196) );
  NOR2_X1 U3633 ( .A1(n3658), .A2(n3657), .ZN(n4295) );
  NAND2_X1 U3634 ( .A1(n3536), .A2(n3535), .ZN(n3542) );
  INV_X1 U3635 ( .A(n6276), .ZN(n5771) );
  CLKBUF_X1 U3636 ( .A(n3508), .Z(n4334) );
  OR2_X1 U3637 ( .A1(n3136), .A2(n4607), .ZN(n3137) );
  CLKBUF_X1 U3638 ( .A(n4456), .Z(n4732) );
  INV_X1 U3639 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3160) );
  AND2_X2 U3640 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4620) );
  AND2_X1 U3641 ( .A1(n5783), .A2(n4837), .ZN(n4744) );
  NAND2_X1 U3642 ( .A1(n4399), .A2(n4289), .ZN(n6557) );
  CLKBUF_X1 U3643 ( .A(n4330), .Z(n5208) );
  AND2_X1 U3644 ( .A1(n5207), .A2(n4259), .ZN(n6697) );
  NAND2_X1 U3645 ( .A1(n4264), .A2(n4263), .ZN(n6695) );
  BUF_X1 U3646 ( .A(n5354), .Z(n5324) );
  INV_X1 U3647 ( .A(n5364), .ZN(n5479) );
  NAND2_X1 U3648 ( .A1(n4551), .A2(n4404), .ZN(n5472) );
  AND2_X1 U3649 ( .A1(n4310), .A2(n4313), .ZN(n6132) );
  CLKBUF_X1 U3650 ( .A(n6117), .Z(n6553) );
  XNOR2_X1 U3651 ( .A(n4249), .B(n4248), .ZN(n5341) );
  OR2_X1 U3652 ( .A1(n4247), .A2(n5362), .ZN(n4249) );
  XOR2_X1 U3653 ( .A(n5333), .B(n5334), .Z(n5364) );
  INV_X1 U3654 ( .A(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n4728) );
  NAND2_X1 U3655 ( .A1(n5504), .A2(n5503), .ZN(n5506) );
  NAND2_X1 U3656 ( .A1(n5512), .A2(n5502), .ZN(n5503) );
  OR2_X1 U3657 ( .A1(n5707), .A2(n3662), .ZN(n5698) );
  INV_X1 U3658 ( .A(n5780), .ZN(n6282) );
  INV_X1 U3659 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n4929) );
  INV_X1 U3660 ( .A(n4732), .ZN(n5788) );
  AND2_X2 U3661 ( .A1(n3160), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4384)
         );
  NAND2_X1 U3662 ( .A1(STATE2_REG_3__SCAN_IN), .A2(n4320), .ZN(n6533) );
  OR2_X1 U3663 ( .A1(n5095), .A2(n5094), .ZN(n5120) );
  NOR2_X1 U3664 ( .A1(n4838), .A2(n4837), .ZN(n5801) );
  INV_X1 U3665 ( .A(n5801), .ZN(n5843) );
  OAI21_X1 U3666 ( .B1(n4998), .B2(n6717), .A(n4994), .ZN(n5020) );
  INV_X1 U3667 ( .A(n6341), .ZN(n4917) );
  NOR2_X1 U3668 ( .A1(n4809), .A2(n4808), .ZN(n4859) );
  INV_X1 U3669 ( .A(n4962), .ZN(n6367) );
  INV_X1 U3670 ( .A(n6388), .ZN(n4794) );
  INV_X1 U3671 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n6443) );
  INV_X1 U3672 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n6536) );
  INV_X1 U3673 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n6717) );
  NAND2_X1 U3674 ( .A1(n4205), .A2(n4204), .ZN(n4206) );
  INV_X1 U3675 ( .A(n4021), .ZN(n4022) );
  AND2_X1 U3676 ( .A1(n3691), .A2(STATE2_REG_2__SCAN_IN), .ZN(n2965) );
  INV_X1 U3677 ( .A(n2967), .ZN(n6160) );
  NAND2_X1 U3678 ( .A1(n3139), .A2(n3146), .ZN(n4405) );
  AND4_X1 U3679 ( .A1(n2985), .A2(n2984), .A3(n2983), .A4(n2982), .ZN(n2966)
         );
  NAND2_X1 U3680 ( .A1(n3386), .A2(n3387), .ZN(n3400) );
  AND2_X1 U3681 ( .A1(n3400), .A2(n3326), .ZN(n2967) );
  AND2_X1 U3682 ( .A1(n3835), .A2(n3834), .ZN(n2968) );
  NAND2_X1 U3683 ( .A1(n2963), .A2(n5579), .ZN(n2969) );
  NOR2_X1 U3684 ( .A1(n2963), .A2(n5606), .ZN(n2970) );
  OAI21_X1 U3685 ( .B1(n3293), .B2(n3180), .A(n3184), .ZN(n3291) );
  NAND2_X1 U3686 ( .A1(n2963), .A2(n5606), .ZN(n2971) );
  NAND2_X1 U3687 ( .A1(n2963), .A2(n6202), .ZN(n2972) );
  AND4_X1 U3688 ( .A1(n3064), .A2(n3063), .A3(n3062), .A4(n3061), .ZN(n2973)
         );
  AND3_X1 U3689 ( .A1(n2991), .A2(n2990), .A3(n2989), .ZN(n2974) );
  AND2_X1 U3690 ( .A1(n4481), .A2(n4486), .ZN(n2975) );
  INV_X1 U3691 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n6567) );
  OR2_X1 U3692 ( .A1(n2967), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n2976)
         );
  NOR2_X1 U3693 ( .A1(n5796), .A2(n4989), .ZN(n2977) );
  NOR2_X1 U3694 ( .A1(n4351), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n2978)
         );
  OR3_X1 U3695 ( .A1(n3434), .A2(INSTADDRPOINTER_REG_24__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n2979) );
  NOR2_X1 U3696 ( .A1(n3146), .A2(n6661), .ZN(n5336) );
  NAND2_X1 U3697 ( .A1(n3691), .A2(n3146), .ZN(n3655) );
  AND2_X1 U3698 ( .A1(n3327), .A2(n3288), .ZN(n3289) );
  INV_X1 U3699 ( .A(n3231), .ZN(n3127) );
  NAND2_X1 U3700 ( .A1(n3328), .A2(n3289), .ZN(n3312) );
  NAND2_X1 U3701 ( .A1(n3691), .A2(n3127), .ZN(n3128) );
  AND2_X1 U3702 ( .A1(n4929), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3456)
         );
  INV_X1 U3703 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3716) );
  NAND2_X1 U3704 ( .A1(n3149), .A2(n4331), .ZN(n3162) );
  INV_X1 U3705 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n2981) );
  INV_X1 U3706 ( .A(n3310), .ZN(n3311) );
  OR2_X1 U3707 ( .A1(n3343), .A2(n3342), .ZN(n3258) );
  INV_X1 U3708 ( .A(n3141), .ZN(n3133) );
  AND2_X1 U3709 ( .A1(n4192), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n4193)
         );
  INV_X1 U3710 ( .A(n3123), .ZN(n3691) );
  NAND2_X1 U3711 ( .A1(n4420), .A2(n3700), .ZN(n3701) );
  INV_X1 U3712 ( .A(EBX_REG_2__SCAN_IN), .ZN(n3534) );
  INV_X1 U3713 ( .A(n3162), .ZN(n3163) );
  AND2_X1 U3714 ( .A1(n4467), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3446) );
  INV_X1 U3715 ( .A(n4405), .ZN(n3048) );
  NOR2_X1 U3716 ( .A1(n2964), .A2(EBX_REG_29__SCAN_IN), .ZN(n3630) );
  AOI22_X1 U3717 ( .A1(n3266), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3060), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3019) );
  CLKBUF_X1 U3718 ( .A(n3716), .Z(n4617) );
  NAND2_X1 U3719 ( .A1(n4193), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4247)
         );
  INV_X1 U3720 ( .A(n5413), .ZN(n4102) );
  NAND2_X1 U3721 ( .A1(n3692), .A2(n4074), .ZN(n3711) );
  NAND2_X1 U3722 ( .A1(n3626), .A2(EBX_REG_2__SCAN_IN), .ZN(n3535) );
  AND2_X1 U3723 ( .A1(n3446), .A2(n4486), .ZN(n3475) );
  OR2_X1 U3724 ( .A1(n3642), .A2(n4477), .ZN(n3080) );
  NAND2_X1 U3725 ( .A1(n3986), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n3988)
         );
  INV_X1 U3726 ( .A(n4668), .ZN(n3577) );
  INV_X1 U3727 ( .A(n5046), .ZN(n3563) );
  INV_X1 U3728 ( .A(n4187), .ZN(n4239) );
  NOR2_X1 U3729 ( .A1(n3950), .A2(n5581), .ZN(n3951) );
  NOR2_X1 U3730 ( .A1(n3854), .A2(n5230), .ZN(n3869) );
  AOI21_X1 U3731 ( .B1(n3741), .B2(n2965), .A(n3740), .ZN(n5030) );
  NAND2_X1 U3732 ( .A1(n3141), .A2(n3231), .ZN(n3148) );
  INV_X1 U3733 ( .A(n5346), .ZN(n5347) );
  OR2_X1 U3734 ( .A1(n2963), .A2(n6225), .ZN(n5240) );
  AND2_X1 U3735 ( .A1(n3533), .A2(n3532), .ZN(n4450) );
  NAND2_X1 U3736 ( .A1(n3694), .A2(n6443), .ZN(n3332) );
  AND2_X1 U3737 ( .A1(n3329), .A2(n3366), .ZN(n4456) );
  AND2_X1 U3738 ( .A1(n4466), .A2(n4465), .ZN(n4499) );
  AND2_X1 U3739 ( .A1(n5385), .A2(REIP_REG_30__SCAN_IN), .ZN(n4285) );
  AND2_X1 U3740 ( .A1(n5341), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4260) );
  NAND2_X1 U3741 ( .A1(n5207), .A2(n4269), .ZN(n6018) );
  INV_X1 U3742 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n6400) );
  AND2_X1 U3743 ( .A1(n3951), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n3986)
         );
  OR2_X1 U3744 ( .A1(n3883), .A2(n5292), .ZN(n3884) );
  NAND2_X1 U3745 ( .A1(n3827), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3751)
         );
  AND2_X1 U3746 ( .A1(PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n3727), .ZN(n3769)
         );
  INV_X1 U3747 ( .A(n6186), .ZN(n5618) );
  INV_X1 U3748 ( .A(n3689), .ZN(n3690) );
  NAND2_X1 U3749 ( .A1(n5564), .A2(n2976), .ZN(n3687) );
  OR2_X1 U3750 ( .A1(n5596), .A2(n5597), .ZN(n5586) );
  NAND2_X1 U3751 ( .A1(n3542), .A2(n3541), .ZN(n4451) );
  INV_X1 U3752 ( .A(n3441), .ZN(n3465) );
  OAI21_X1 U3753 ( .B1(n6560), .B2(n4629), .A(n6533), .ZN(n4465) );
  OR2_X1 U3754 ( .A1(n4829), .A2(n5783), .ZN(n4838) );
  INV_X1 U3755 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6419) );
  OR2_X1 U3756 ( .A1(n4516), .A2(n4837), .ZN(n6391) );
  NAND2_X1 U3757 ( .A1(n3508), .A2(n4467), .ZN(n4296) );
  INV_X1 U3758 ( .A(n4013), .ZN(n6556) );
  OR2_X1 U3759 ( .A1(n4285), .A2(n4284), .ZN(n4286) );
  NOR2_X1 U3760 ( .A1(n5680), .A2(n5455), .ZN(n5456) );
  OR2_X1 U3761 ( .A1(n6688), .A2(n4277), .ZN(n5895) );
  NOR2_X1 U3762 ( .A1(n6018), .A2(n4271), .ZN(n6002) );
  OR2_X1 U3763 ( .A1(n6557), .A2(n4246), .ZN(n6074) );
  AND2_X1 U3764 ( .A1(n6074), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6078) );
  AND2_X1 U3765 ( .A1(n5456), .A2(n5415), .ZN(n5417) );
  OR2_X1 U3766 ( .A1(n5062), .A2(n5941), .ZN(n5944) );
  OR2_X1 U3767 ( .A1(n5049), .A2(n5048), .ZN(n5051) );
  CLKBUF_X1 U3768 ( .A(n4575), .Z(n4717) );
  NAND2_X1 U3769 ( .A1(n5334), .A2(n4201), .ZN(n5367) );
  INV_X1 U3770 ( .A(n5246), .ZN(n5304) );
  AND2_X1 U3771 ( .A1(n5472), .A2(n3048), .ZN(n5499) );
  OAI21_X1 U3772 ( .B1(n5874), .B2(n5634), .A(n4020), .ZN(n4021) );
  CLKBUF_X1 U3773 ( .A(n4661), .Z(n4923) );
  AND2_X1 U3774 ( .A1(n5041), .A2(n4983), .ZN(n5087) );
  NOR2_X1 U3775 ( .A1(n3743), .A2(n3742), .ZN(n3750) );
  INV_X1 U3776 ( .A(n6195), .ZN(n6164) );
  AND2_X1 U3777 ( .A1(n6169), .A2(n4015), .ZN(n6186) );
  NAND2_X1 U3778 ( .A1(n5350), .A2(n5349), .ZN(n5351) );
  XNOR2_X1 U3779 ( .A(n5539), .B(n3690), .ZN(n5689) );
  NOR2_X1 U3780 ( .A1(n5558), .A2(n5559), .ZN(n5557) );
  INV_X1 U3781 ( .A(n5586), .ZN(n5595) );
  INV_X1 U3782 ( .A(n6249), .ZN(n6280) );
  NAND2_X1 U3783 ( .A1(n3515), .A2(n3514), .ZN(n3669) );
  NAND2_X1 U3784 ( .A1(n6443), .A2(n4465), .ZN(n4991) );
  INV_X1 U3785 ( .A(n6391), .ZN(n5124) );
  INV_X1 U3786 ( .A(n4838), .ZN(n4831) );
  INV_X1 U3787 ( .A(n6308), .ZN(n5841) );
  INV_X1 U3788 ( .A(n4920), .ZN(n6318) );
  OR2_X1 U3789 ( .A1(n4655), .A2(n5783), .ZN(n4464) );
  INV_X1 U3790 ( .A(n4858), .ZN(n6336) );
  INV_X1 U3791 ( .A(n5128), .ZN(n5185) );
  INV_X1 U3792 ( .A(n6373), .ZN(n5129) );
  NOR2_X1 U3793 ( .A1(n4743), .A2(n4732), .ZN(n4803) );
  INV_X1 U3794 ( .A(n4837), .ZN(n4808) );
  OR2_X1 U3795 ( .A1(n4308), .A2(n4296), .ZN(n4399) );
  NOR2_X1 U3796 ( .A1(n4287), .A2(n4286), .ZN(n4288) );
  INV_X1 U3797 ( .A(n6078), .ZN(n6693) );
  NAND2_X1 U3798 ( .A1(n6074), .A2(n4250), .ZN(n5995) );
  INV_X1 U3799 ( .A(n6697), .ZN(n6085) );
  INV_X1 U3800 ( .A(n5087), .ZN(n5228) );
  INV_X1 U3801 ( .A(n5499), .ZN(n5203) );
  OR2_X1 U3802 ( .A1(n6132), .A2(n6117), .ZN(n6119) );
  INV_X1 U3803 ( .A(n6132), .ZN(n6138) );
  NOR2_X1 U3804 ( .A1(n4207), .A2(n4206), .ZN(n4208) );
  OR2_X1 U3805 ( .A1(n6186), .A2(n4423), .ZN(n6195) );
  NAND2_X1 U3806 ( .A1(n5689), .A2(n6282), .ZN(n5694) );
  NOR2_X1 U3807 ( .A1(n5732), .A2(n5770), .ZN(n6196) );
  NAND2_X1 U3808 ( .A1(n4831), .A2(n4837), .ZN(n5127) );
  NAND2_X1 U3809 ( .A1(n4745), .A2(n4744), .ZN(n6308) );
  OR2_X1 U3810 ( .A1(n4464), .A2(n4808), .ZN(n5026) );
  OR2_X1 U3811 ( .A1(n4464), .A2(n4837), .ZN(n4920) );
  INV_X1 U3812 ( .A(n4859), .ZN(n4895) );
  NAND2_X1 U3813 ( .A1(n4799), .A2(n4808), .ZN(n5128) );
  NAND2_X1 U3814 ( .A1(n4803), .A2(n4744), .ZN(n6373) );
  NAND2_X1 U3815 ( .A1(n4670), .A2(n4808), .ZN(n4797) );
  OAI21_X1 U3816 ( .B1(n5479), .B2(n5995), .A(n4288), .ZN(U2797) );
  INV_X1 U3817 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5659) );
  AND2_X2 U3818 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n2980), .ZN(n2992)
         );
  AND2_X2 U3819 ( .A1(n2992), .A2(n4384), .ZN(n3279) );
  BUF_X4 U3820 ( .A(n3279), .Z(n4112) );
  AND2_X2 U3821 ( .A1(n4384), .A2(n4620), .ZN(n3189) );
  AOI22_X1 U3822 ( .A1(n4112), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3189), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n2985) );
  NOR2_X4 U3823 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4621) );
  AND2_X2 U3824 ( .A1(n2992), .A2(n4621), .ZN(n3039) );
  BUF_X4 U3825 ( .A(n3039), .Z(n4150) );
  CLKBUF_X3 U3826 ( .A(n2987), .Z(n4610) );
  AND2_X2 U3827 ( .A1(n4384), .A2(n4610), .ZN(n3223) );
  AOI22_X1 U3828 ( .A1(n4150), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3223), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n2984) );
  AND2_X2 U3829 ( .A1(n2987), .A2(n4621), .ZN(n3094) );
  AND2_X2 U3830 ( .A1(n4620), .A2(n2986), .ZN(n3190) );
  AOI22_X1 U3831 ( .A1(n3094), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n3190), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n2983) );
  AND2_X2 U3832 ( .A1(n2981), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4381)
         );
  AND2_X2 U3833 ( .A1(n3716), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n2988)
         );
  AND2_X2 U3834 ( .A1(n4381), .A2(n2988), .ZN(n3224) );
  AND2_X2 U3835 ( .A1(n4621), .A2(n4620), .ZN(n3015) );
  AOI22_X1 U3836 ( .A1(n3224), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3015), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n2982) );
  AND2_X2 U3837 ( .A1(n2992), .A2(n2986), .ZN(n3049) );
  AND2_X2 U3838 ( .A1(n2988), .A2(n4621), .ZN(n4174) );
  AOI22_X1 U3839 ( .A1(n3049), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4174), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n2991) );
  AND2_X2 U3840 ( .A1(n2987), .A2(n2986), .ZN(n3030) );
  AOI22_X1 U3841 ( .A1(n3218), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3030), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n2990) );
  AND2_X2 U3842 ( .A1(n4384), .A2(n2988), .ZN(n3081) );
  AND2_X2 U3843 ( .A1(n4381), .A2(n4610), .ZN(n4210) );
  AOI22_X1 U3844 ( .A1(n3081), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n4210), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n2989) );
  AND2_X2 U3845 ( .A1(n4381), .A2(n4620), .ZN(n3060) );
  AOI22_X1 U3846 ( .A1(n3266), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3060), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n2993) );
  NAND3_X2 U3847 ( .A1(n2966), .A2(n2974), .A3(n2993), .ZN(n3123) );
  INV_X1 U3848 ( .A(n3123), .ZN(n3014) );
  NAND2_X1 U3849 ( .A1(n3081), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n2997) );
  NAND2_X1 U3850 ( .A1(n4210), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n2996) );
  NAND2_X1 U3851 ( .A1(n3049), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n2995)
         );
  NAND2_X1 U3852 ( .A1(n4174), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n2994) );
  NAND2_X1 U3853 ( .A1(n3060), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3001)
         );
  NAND2_X1 U3854 ( .A1(n3266), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3000)
         );
  NAND2_X1 U3855 ( .A1(n3218), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n2999) );
  NAND2_X1 U3856 ( .A1(n3030), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n2998) );
  NAND2_X1 U3858 ( .A1(n3224), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3005) );
  NAND2_X1 U3859 ( .A1(n4150), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3004) );
  NAND2_X1 U3860 ( .A1(n3223), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3003) );
  NAND2_X1 U3861 ( .A1(n3015), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3002)
         );
  NAND2_X1 U3863 ( .A1(n3279), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3009) );
  NAND2_X1 U3864 ( .A1(n3189), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3008)
         );
  NAND2_X1 U3865 ( .A1(n3094), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3007) );
  NAND2_X1 U3866 ( .A1(n3190), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3006)
         );
  NAND2_X2 U3867 ( .A1(n3014), .A2(n3141), .ZN(n3139) );
  AOI22_X1 U3868 ( .A1(n4210), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3049), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3018) );
  AOI22_X1 U3869 ( .A1(n3189), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4174), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3017) );
  AOI22_X1 U3870 ( .A1(n3223), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3015), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3016) );
  NAND4_X1 U3871 ( .A1(n3019), .A2(n3018), .A3(n3017), .A4(n3016), .ZN(n3025)
         );
  BUF_X2 U3872 ( .A(n3279), .Z(n4220) );
  AOI22_X1 U3873 ( .A1(n4220), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3081), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3023) );
  BUF_X2 U3874 ( .A(n3039), .Z(n4131) );
  AOI22_X1 U3875 ( .A1(n3224), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n4131), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3022) );
  BUF_X4 U3876 ( .A(n3030), .Z(n4157) );
  AOI22_X1 U3877 ( .A1(n3218), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4157), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3021) );
  AOI22_X1 U3878 ( .A1(n3094), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n3190), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3020) );
  NAND4_X1 U3879 ( .A1(n3023), .A2(n3022), .A3(n3021), .A4(n3020), .ZN(n3024)
         );
  NAND2_X1 U3880 ( .A1(n3081), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3029) );
  NAND2_X1 U3881 ( .A1(n4210), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3028) );
  NAND2_X1 U3882 ( .A1(n3049), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3027)
         );
  NAND2_X1 U3883 ( .A1(n4174), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3026) );
  NAND2_X1 U3884 ( .A1(n3060), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3034)
         );
  NAND2_X1 U3885 ( .A1(n3266), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3033)
         );
  NAND2_X1 U3886 ( .A1(n3218), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3032) );
  BUF_X2 U3887 ( .A(n3030), .Z(n4176) );
  NAND2_X1 U3888 ( .A1(n4176), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3031) );
  NAND2_X1 U3889 ( .A1(n4112), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3038) );
  NAND2_X1 U3890 ( .A1(n3189), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3037)
         );
  CLKBUF_X3 U3891 ( .A(n3094), .Z(n4151) );
  NAND2_X1 U3892 ( .A1(n4151), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3036) );
  NAND2_X1 U3893 ( .A1(n3190), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3035)
         );
  NAND2_X1 U3894 ( .A1(n3224), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3043) );
  NAND2_X1 U3895 ( .A1(n3039), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3042) );
  NAND2_X1 U3896 ( .A1(n3223), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3041) );
  NAND2_X1 U3897 ( .A1(n3015), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3040)
         );
  NAND2_X1 U3898 ( .A1(n3126), .A2(n3231), .ZN(n3147) );
  NAND2_X1 U3899 ( .A1(n3048), .A2(n3125), .ZN(n3495) );
  AOI22_X1 U3900 ( .A1(n3266), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3060), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3053) );
  AOI22_X1 U3901 ( .A1(n3081), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n4210), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3052) );
  AOI22_X1 U3902 ( .A1(n3049), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4174), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3051) );
  AOI22_X1 U3903 ( .A1(n3218), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4157), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3050) );
  NAND4_X1 U3904 ( .A1(n3053), .A2(n3052), .A3(n3051), .A4(n3050), .ZN(n3059)
         );
  AOI22_X1 U3905 ( .A1(n4220), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3189), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3057) );
  AOI22_X1 U3906 ( .A1(n4150), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3223), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3056) );
  AOI22_X1 U3907 ( .A1(n3094), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3190), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3055) );
  AOI22_X1 U3908 ( .A1(n3224), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3015), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3054) );
  NAND4_X1 U3909 ( .A1(n3057), .A2(n3056), .A3(n3055), .A4(n3054), .ZN(n3058)
         );
  NAND2_X1 U3911 ( .A1(n3060), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3064)
         );
  NAND2_X1 U3912 ( .A1(n3266), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3063)
         );
  NAND2_X1 U3913 ( .A1(n3049), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3062)
         );
  NAND2_X1 U3914 ( .A1(n4210), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3061) );
  NAND2_X1 U3915 ( .A1(n3189), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3068)
         );
  NAND2_X1 U3916 ( .A1(n4150), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3067) );
  NAND2_X1 U3917 ( .A1(n3224), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3066) );
  NAND2_X1 U3918 ( .A1(n3094), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3065) );
  NAND2_X1 U3919 ( .A1(n3218), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3072) );
  NAND2_X1 U3920 ( .A1(n3081), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3071) );
  NAND2_X1 U3921 ( .A1(n4174), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3070) );
  NAND2_X1 U3922 ( .A1(n4176), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3069) );
  NAND2_X1 U3923 ( .A1(n4112), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3076) );
  NAND2_X1 U3924 ( .A1(n3223), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3075) );
  NAND2_X1 U3925 ( .A1(n3190), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3074)
         );
  NAND2_X1 U3926 ( .A1(n3015), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3073)
         );
  AND4_X2 U3927 ( .A1(n2973), .A2(n3079), .A3(n3078), .A4(n3077), .ZN(n3511)
         );
  NOR2_X2 U3928 ( .A1(n3495), .A2(n3080), .ZN(n3508) );
  NAND2_X1 U3929 ( .A1(n3060), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3085)
         );
  NAND2_X1 U3930 ( .A1(n3266), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3084)
         );
  NAND2_X1 U3931 ( .A1(n3081), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3083) );
  NAND2_X1 U3932 ( .A1(n4176), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3082) );
  AND4_X2 U3933 ( .A1(n3085), .A2(n3084), .A3(n3083), .A4(n3082), .ZN(n3102)
         );
  NAND2_X1 U3934 ( .A1(n4210), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3089) );
  NAND2_X1 U3935 ( .A1(n3218), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3088) );
  NAND2_X1 U3936 ( .A1(n3049), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3087)
         );
  NAND2_X1 U3937 ( .A1(n4174), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3086) );
  NAND2_X1 U3938 ( .A1(n3189), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3093)
         );
  NAND2_X1 U3939 ( .A1(n4150), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3092) );
  NAND2_X1 U3940 ( .A1(n3224), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3091) );
  NAND2_X1 U3941 ( .A1(n3190), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3090)
         );
  NAND2_X1 U3943 ( .A1(n4112), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3098) );
  NAND2_X1 U3944 ( .A1(n3223), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3097) );
  NAND2_X1 U3945 ( .A1(n3094), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3096) );
  NAND2_X1 U3946 ( .A1(n3015), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3095)
         );
  AND4_X2 U3947 ( .A1(n3098), .A2(n3097), .A3(n3096), .A4(n3095), .ZN(n3099)
         );
  BUF_X4 U3948 ( .A(n3518), .Z(n4467) );
  NAND2_X1 U3949 ( .A1(n3081), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3106) );
  NAND2_X1 U3950 ( .A1(n4210), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3105) );
  NAND2_X1 U3951 ( .A1(n3049), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3104)
         );
  NAND2_X1 U3952 ( .A1(n4174), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3103) );
  NAND2_X1 U3953 ( .A1(n3224), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3110) );
  NAND2_X1 U3954 ( .A1(n4150), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3109) );
  NAND2_X1 U3955 ( .A1(n3223), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3108) );
  NAND2_X1 U3956 ( .A1(n3015), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3107)
         );
  NAND2_X1 U3957 ( .A1(n3060), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3114)
         );
  NAND2_X1 U3958 ( .A1(n3266), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3113)
         );
  NAND2_X1 U3959 ( .A1(n3218), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3112) );
  NAND2_X1 U3960 ( .A1(n4157), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3111) );
  AND4_X2 U3961 ( .A1(n3114), .A2(n3113), .A3(n3112), .A4(n3111), .ZN(n3120)
         );
  NAND2_X1 U3962 ( .A1(n4112), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3118) );
  NAND2_X1 U3963 ( .A1(n3189), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3117)
         );
  NAND2_X1 U3964 ( .A1(n4151), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3116) );
  NAND2_X1 U3965 ( .A1(n3190), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3115)
         );
  AND4_X2 U3966 ( .A1(n3118), .A2(n3117), .A3(n3116), .A4(n3115), .ZN(n3119)
         );
  NAND4_X4 U3967 ( .A1(n3122), .A2(n3121), .A3(n3120), .A4(n3119), .ZN(n3517)
         );
  INV_X1 U3968 ( .A(STATE_REG_1__SCAN_IN), .ZN(n6462) );
  XNOR2_X1 U3969 ( .A(n6462), .B(STATE_REG_2__SCAN_IN), .ZN(n3498) );
  NOR2_X1 U3970 ( .A1(n3517), .A2(n3498), .ZN(n3142) );
  NAND2_X1 U3971 ( .A1(n3139), .A2(n4473), .ZN(n3168) );
  NAND2_X1 U3972 ( .A1(n3168), .A2(n3146), .ZN(n3151) );
  INV_X1 U3973 ( .A(n3147), .ZN(n3125) );
  NAND3_X1 U3974 ( .A1(n3125), .A2(n3655), .A3(n3124), .ZN(n3131) );
  NAND2_X1 U3975 ( .A1(n3126), .A2(n3128), .ZN(n3129) );
  NAND2_X1 U3976 ( .A1(n3129), .A2(n3511), .ZN(n3130) );
  NAND2_X1 U3977 ( .A1(n3131), .A2(n3130), .ZN(n3153) );
  INV_X2 U3978 ( .A(n3517), .ZN(n3509) );
  NOR2_X4 U3979 ( .A1(n4467), .A2(n3517), .ZN(n3154) );
  NOR2_X2 U3980 ( .A1(n3124), .A2(n4473), .ZN(n3167) );
  NAND3_X1 U3981 ( .A1(n3154), .A2(n3133), .A3(n3167), .ZN(n4332) );
  NAND2_X1 U3982 ( .A1(n4477), .A2(n3146), .ZN(n5249) );
  OAI211_X1 U3983 ( .C1(n4296), .C2(n3142), .A(n3516), .B(n3638), .ZN(n3134)
         );
  NAND2_X1 U3984 ( .A1(n3134), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3159) );
  INV_X1 U3985 ( .A(n3159), .ZN(n3138) );
  NAND2_X1 U3986 ( .A1(n6536), .A2(n6717), .ZN(n6542) );
  XNOR2_X1 U3987 ( .A(n4929), .B(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n5796)
         );
  AND2_X1 U3988 ( .A1(n6536), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3506) );
  INV_X1 U3989 ( .A(n3506), .ZN(n6429) );
  AND2_X1 U3990 ( .A1(n6429), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3135)
         );
  AOI21_X1 U3991 ( .B1(n6556), .B2(n5796), .A(n3135), .ZN(n3158) );
  INV_X1 U3992 ( .A(n3158), .ZN(n3136) );
  NAND2_X1 U3993 ( .A1(n3138), .A2(n3137), .ZN(n3161) );
  NAND2_X1 U3994 ( .A1(n3139), .A2(n4467), .ZN(n3493) );
  INV_X2 U3995 ( .A(n3231), .ZN(n4486) );
  INV_X1 U3996 ( .A(n3518), .ZN(n3650) );
  NAND2_X1 U3997 ( .A1(n3650), .A2(n3517), .ZN(n4293) );
  BUF_X2 U3998 ( .A(n3141), .Z(n4481) );
  NAND2_X1 U3999 ( .A1(n4293), .A2(n4481), .ZN(n3144) );
  INV_X1 U4000 ( .A(n3142), .ZN(n3143) );
  AOI21_X1 U4001 ( .B1(n3144), .B2(n3143), .A(n3642), .ZN(n3145) );
  OAI211_X1 U4002 ( .C1(n3231), .C2(n3493), .A(n3646), .B(n3145), .ZN(n3150)
         );
  INV_X1 U4003 ( .A(n3146), .ZN(n5473) );
  OAI21_X1 U4004 ( .B1(n3147), .B2(n5473), .A(n4294), .ZN(n3149) );
  AND2_X4 U4005 ( .A1(n4473), .A2(n3517), .ZN(n5261) );
  NAND2_X1 U4006 ( .A1(n3520), .A2(n5261), .ZN(n4331) );
  NOR2_X1 U4007 ( .A1(n3150), .A2(n3162), .ZN(n3156) );
  INV_X1 U4008 ( .A(n3151), .ZN(n3152) );
  NAND2_X1 U4009 ( .A1(n3153), .A2(n3152), .ZN(n3155) );
  NAND2_X1 U4010 ( .A1(n3156), .A2(n3649), .ZN(n3157) );
  NAND2_X2 U4011 ( .A1(n3157), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3293) );
  OAI211_X1 U4012 ( .C1(n3293), .C2(n3160), .A(n3159), .B(n3158), .ZN(n3177)
         );
  NAND2_X1 U4013 ( .A1(n3161), .A2(n3177), .ZN(n3201) );
  INV_X1 U4014 ( .A(n3201), .ZN(n3176) );
  NAND2_X1 U4015 ( .A1(n3649), .A2(n3163), .ZN(n3173) );
  NAND2_X1 U4016 ( .A1(n3495), .A2(n3887), .ZN(n3164) );
  NAND2_X1 U4017 ( .A1(n3164), .A2(n4473), .ZN(n3165) );
  NAND2_X1 U4018 ( .A1(n3165), .A2(n4494), .ZN(n3171) );
  OR2_X1 U4019 ( .A1(n6542), .A2(n6443), .ZN(n6446) );
  AOI21_X1 U4020 ( .B1(n3166), .B2(n3167), .A(n6446), .ZN(n3170) );
  INV_X1 U4021 ( .A(n3154), .ZN(n4400) );
  OAI211_X1 U4022 ( .C1(n3650), .C2(n3124), .A(n3652), .B(n4400), .ZN(n3644)
         );
  NAND2_X1 U4023 ( .A1(n3168), .A2(n4294), .ZN(n3169) );
  NAND4_X1 U4024 ( .A1(n3171), .A2(n3170), .A3(n3644), .A4(n3169), .ZN(n3172)
         );
  MUX2_X1 U4025 ( .A(n6429), .B(n6556), .S(n4929), .Z(n3174) );
  INV_X1 U4026 ( .A(n3174), .ZN(n3175) );
  NAND2_X1 U4028 ( .A1(n3176), .A2(n3202), .ZN(n3179) );
  NAND2_X2 U4029 ( .A1(n3179), .A2(n3178), .ZN(n3290) );
  INV_X1 U4030 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3180) );
  AND2_X1 U4031 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3181) );
  NAND2_X1 U4032 ( .A1(n3181), .A2(n4830), .ZN(n4737) );
  INV_X1 U4033 ( .A(n3181), .ZN(n3182) );
  NAND2_X1 U4034 ( .A1(n3182), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3183) );
  NAND2_X1 U4035 ( .A1(n4737), .A2(n3183), .ZN(n4766) );
  AOI22_X1 U4036 ( .A1(n6556), .A2(n4766), .B1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n6429), .ZN(n3184) );
  XNOR2_X1 U4037 ( .A(n3290), .B(n3291), .ZN(n4330) );
  NAND2_X1 U4038 ( .A1(n4330), .A2(n6443), .ZN(n3198) );
  INV_X1 U4039 ( .A(n3259), .ZN(n4392) );
  AOI22_X1 U4040 ( .A1(n2962), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3060), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3188) );
  AOI22_X1 U4041 ( .A1(n4211), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n4173), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3187) );
  AOI22_X1 U4042 ( .A1(n3049), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4156), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3186) );
  AOI22_X1 U4043 ( .A1(n4214), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4157), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3185) );
  NAND4_X1 U4044 ( .A1(n3188), .A2(n3187), .A3(n3186), .A4(n3185), .ZN(n3196)
         );
  AOI22_X1 U4045 ( .A1(n4220), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4219), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3194) );
  BUF_X1 U4046 ( .A(n4131), .Z(n4222) );
  INV_X1 U4047 ( .A(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n6677) );
  BUF_X1 U4048 ( .A(n3223), .Z(n4107) );
  AOI22_X1 U4049 ( .A1(n4222), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4107), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3193) );
  INV_X1 U4050 ( .A(n3190), .ZN(n3261) );
  AOI22_X1 U4051 ( .A1(n4224), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n4223), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3192) );
  AOI22_X1 U4052 ( .A1(n3232), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n4225), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3191) );
  NAND4_X1 U4053 ( .A1(n3194), .A2(n3193), .A3(n3192), .A4(n3191), .ZN(n3195)
         );
  NAND2_X1 U4054 ( .A1(n4392), .A2(n3359), .ZN(n3197) );
  INV_X1 U4055 ( .A(n3260), .ZN(n3254) );
  AOI22_X1 U4056 ( .A1(n3475), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3254), 
        .B2(n3359), .ZN(n3199) );
  XNOR2_X2 U4057 ( .A(n3200), .B(n3199), .ZN(n3328) );
  AOI22_X1 U4059 ( .A1(n4220), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4175), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3207) );
  AOI22_X1 U4060 ( .A1(n4222), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4107), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3206) );
  AOI22_X1 U4061 ( .A1(n4078), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n4214), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3205) );
  AOI22_X1 U4062 ( .A1(n3232), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n4225), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3204) );
  NAND4_X1 U4063 ( .A1(n3207), .A2(n3206), .A3(n3205), .A4(n3204), .ZN(n3213)
         );
  AOI22_X1 U4064 ( .A1(n4211), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n4173), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3211) );
  AOI22_X1 U4065 ( .A1(n4219), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n4156), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3210) );
  AOI22_X1 U4066 ( .A1(n3888), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4157), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3209) );
  AOI22_X1 U4067 ( .A1(n4224), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n4223), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3208) );
  NAND4_X1 U4068 ( .A1(n3211), .A2(n3210), .A3(n3209), .A4(n3208), .ZN(n3212)
         );
  NAND2_X1 U4069 ( .A1(n4392), .A2(n3347), .ZN(n3214) );
  XNOR2_X1 U4070 ( .A(n3217), .B(n3216), .ZN(n3694) );
  AOI22_X1 U4071 ( .A1(n2962), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3060), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3222) );
  AOI22_X1 U4072 ( .A1(n4211), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n4173), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3221) );
  AOI22_X1 U4073 ( .A1(n3049), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4156), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3220) );
  AOI22_X1 U4074 ( .A1(n4214), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n4157), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3219) );
  NAND4_X1 U4075 ( .A1(n3222), .A2(n3221), .A3(n3220), .A4(n3219), .ZN(n3230)
         );
  AOI22_X1 U4076 ( .A1(n4220), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4219), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3228) );
  AOI22_X1 U4077 ( .A1(n4222), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4221), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3227) );
  AOI22_X1 U4078 ( .A1(n4224), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n4223), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3226) );
  AOI22_X1 U4079 ( .A1(n3232), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4225), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3225) );
  NAND4_X1 U4080 ( .A1(n3228), .A2(n3227), .A3(n3226), .A4(n3225), .ZN(n3229)
         );
  NOR2_X1 U4081 ( .A1(n3259), .A2(n3410), .ZN(n3253) );
  NAND2_X1 U4082 ( .A1(n3231), .A2(n3410), .ZN(n3247) );
  NOR2_X1 U4083 ( .A1(n3247), .A2(n6443), .ZN(n3251) );
  AOI22_X1 U4084 ( .A1(n3888), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3060), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3236) );
  AOI22_X1 U4085 ( .A1(n3232), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n4131), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3235) );
  AOI22_X1 U4086 ( .A1(n3049), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4156), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3234) );
  AOI22_X1 U4087 ( .A1(n4220), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n4151), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3233) );
  NAND4_X1 U4088 ( .A1(n3236), .A2(n3235), .A3(n3234), .A4(n3233), .ZN(n3242)
         );
  AOI22_X1 U4089 ( .A1(n3081), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n4173), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3240) );
  AOI22_X1 U4090 ( .A1(n4214), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n4157), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3239) );
  AOI22_X1 U4091 ( .A1(n4221), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n4225), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3238) );
  AOI22_X1 U4092 ( .A1(n4219), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n4223), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3237) );
  NAND4_X1 U4093 ( .A1(n3240), .A2(n3239), .A3(n3238), .A4(n3237), .ZN(n3241)
         );
  INV_X1 U4094 ( .A(n3346), .ZN(n3243) );
  MUX2_X1 U4095 ( .A(n3253), .B(n3251), .S(n3243), .Z(n3333) );
  INV_X1 U4096 ( .A(n3333), .ZN(n3244) );
  NAND2_X1 U4097 ( .A1(n3332), .A2(n3244), .ZN(n3250) );
  NAND2_X1 U4098 ( .A1(n3475), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3249) );
  INV_X1 U4099 ( .A(n3446), .ZN(n3245) );
  OAI21_X1 U4100 ( .B1(n3346), .B2(n6443), .A(n3245), .ZN(n3246) );
  AND2_X1 U4101 ( .A1(n3247), .A2(n3246), .ZN(n3248) );
  NAND2_X1 U4102 ( .A1(n3249), .A2(n3248), .ZN(n3334) );
  NAND2_X1 U4103 ( .A1(n3250), .A2(n3334), .ZN(n3252) );
  INV_X1 U4104 ( .A(n3251), .ZN(n3325) );
  INV_X1 U4105 ( .A(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3257) );
  INV_X1 U4106 ( .A(n3253), .ZN(n3256) );
  NAND2_X1 U4107 ( .A1(n3254), .A2(n3347), .ZN(n3255) );
  OAI211_X1 U4108 ( .C1(n3460), .C2(n3257), .A(n3256), .B(n3255), .ZN(n3342)
         );
  INV_X1 U4109 ( .A(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3274) );
  AOI22_X1 U4110 ( .A1(n4173), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n4214), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3265) );
  AOI22_X1 U4111 ( .A1(n4211), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n4175), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3264) );
  AOI22_X1 U4112 ( .A1(n3961), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4156), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3263) );
  AOI22_X1 U4113 ( .A1(n4222), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4223), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3262) );
  NAND4_X1 U4114 ( .A1(n3265), .A2(n3264), .A3(n3263), .A4(n3262), .ZN(n3272)
         );
  AOI22_X1 U4115 ( .A1(n2962), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3060), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3270) );
  AOI22_X1 U4116 ( .A1(n3232), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n4107), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3269) );
  AOI22_X1 U4117 ( .A1(n4219), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n4157), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3268) );
  AOI22_X1 U4118 ( .A1(n4224), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n4225), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3267) );
  NAND4_X1 U4119 ( .A1(n3270), .A2(n3269), .A3(n3268), .A4(n3267), .ZN(n3271)
         );
  OR2_X1 U4120 ( .A1(n3272), .A2(n3271), .ZN(n3390) );
  NAND2_X1 U4121 ( .A1(n3483), .A2(n3390), .ZN(n3273) );
  OAI21_X1 U4122 ( .B1(n3460), .B2(n3274), .A(n3273), .ZN(n3377) );
  INV_X1 U4123 ( .A(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3287) );
  AOI22_X1 U4124 ( .A1(n3888), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3060), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3278) );
  AOI22_X1 U4125 ( .A1(INSTQUEUE_REG_3__4__SCAN_IN), .A2(n4173), .B1(n4211), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3277) );
  AOI22_X1 U4126 ( .A1(n3049), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4156), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3276) );
  AOI22_X1 U4127 ( .A1(n4214), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n4157), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3275) );
  NAND4_X1 U4128 ( .A1(n3278), .A2(n3277), .A3(n3276), .A4(n3275), .ZN(n3285)
         );
  AOI22_X1 U4129 ( .A1(INSTQUEUE_REG_10__4__SCAN_IN), .A2(n3961), .B1(n4219), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3283) );
  AOI22_X1 U4130 ( .A1(INSTQUEUE_REG_2__4__SCAN_IN), .A2(n4107), .B1(n4131), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3282) );
  AOI22_X1 U4131 ( .A1(n4224), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n4223), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3281) );
  AOI22_X1 U4132 ( .A1(n3232), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n4225), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3280) );
  NAND4_X1 U4133 ( .A1(n3283), .A2(n3282), .A3(n3281), .A4(n3280), .ZN(n3284)
         );
  OR2_X1 U4134 ( .A1(n3285), .A2(n3284), .ZN(n3391) );
  NAND2_X1 U4135 ( .A1(n3483), .A2(n3391), .ZN(n3286) );
  OAI21_X1 U4136 ( .B1(n3460), .B2(n3287), .A(n3286), .ZN(n3375) );
  AND2_X1 U4137 ( .A1(n3377), .A2(n3375), .ZN(n3288) );
  INV_X1 U4138 ( .A(n3293), .ZN(n3294) );
  NAND2_X1 U4139 ( .A1(n3294), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3299) );
  NAND2_X1 U4140 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6711) );
  OR2_X1 U4141 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6711), .ZN(n4898)
         );
  INV_X1 U4142 ( .A(n4898), .ZN(n3295) );
  NAND2_X1 U4143 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n3295), .ZN(n6324) );
  NAND2_X1 U4144 ( .A1(n6419), .A2(n6324), .ZN(n3296) );
  NAND3_X1 U4145 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .ZN(n4760) );
  INV_X1 U4146 ( .A(n4760), .ZN(n4513) );
  NAND2_X1 U4147 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4513), .ZN(n4580) );
  NAND2_X1 U4148 ( .A1(n3296), .A2(n4580), .ZN(n4989) );
  OAI22_X1 U4149 ( .A1(n4013), .A2(n4989), .B1(n3506), .B2(n6419), .ZN(n3297)
         );
  INV_X1 U4150 ( .A(n3297), .ZN(n3298) );
  AOI22_X1 U4151 ( .A1(n2962), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4214), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3303) );
  AOI22_X1 U4152 ( .A1(n4222), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4107), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3302) );
  AOI22_X1 U4153 ( .A1(n4211), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n4156), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3301) );
  AOI22_X1 U4154 ( .A1(n4225), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4223), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3300) );
  NAND4_X1 U4155 ( .A1(n3303), .A2(n3302), .A3(n3301), .A4(n3300), .ZN(n3309)
         );
  AOI22_X1 U4156 ( .A1(n4173), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n4175), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3307) );
  AOI22_X1 U4157 ( .A1(n4220), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4219), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3306) );
  AOI22_X1 U4158 ( .A1(n4078), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n4157), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3305) );
  AOI22_X1 U4159 ( .A1(n3232), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4151), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3304) );
  NAND4_X1 U4160 ( .A1(n3307), .A2(n3306), .A3(n3305), .A4(n3304), .ZN(n3308)
         );
  OR2_X1 U4161 ( .A1(n3309), .A2(n3308), .ZN(n3368) );
  AOI22_X1 U4162 ( .A1(n3475), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3483), 
        .B2(n3368), .ZN(n3310) );
  NOR2_X2 U4163 ( .A1(n3312), .A2(n4457), .ZN(n3386) );
  INV_X1 U4164 ( .A(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3324) );
  AOI22_X1 U4165 ( .A1(n3888), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3060), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3316) );
  AOI22_X1 U4166 ( .A1(n4211), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4173), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3315) );
  AOI22_X1 U4167 ( .A1(n3049), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4156), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3314) );
  AOI22_X1 U4168 ( .A1(n4214), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4213), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3313) );
  NAND4_X1 U4169 ( .A1(n3316), .A2(n3315), .A3(n3314), .A4(n3313), .ZN(n3322)
         );
  AOI22_X1 U4170 ( .A1(n3961), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4219), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3320) );
  AOI22_X1 U4171 ( .A1(n4222), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4107), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3319) );
  AOI22_X1 U4172 ( .A1(n4224), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n4223), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3318) );
  AOI22_X1 U4173 ( .A1(n3232), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n4225), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3317) );
  NAND4_X1 U4174 ( .A1(n3320), .A2(n3319), .A3(n3318), .A4(n3317), .ZN(n3321)
         );
  OR2_X1 U4175 ( .A1(n3322), .A2(n3321), .ZN(n3402) );
  NAND2_X1 U4176 ( .A1(n3483), .A2(n3402), .ZN(n3323) );
  OAI21_X1 U4177 ( .B1(n3460), .B2(n3324), .A(n3323), .ZN(n3387) );
  NOR2_X1 U4178 ( .A1(n3325), .A2(n3465), .ZN(n3326) );
  NAND2_X1 U4179 ( .A1(n3347), .A2(n3346), .ZN(n3361) );
  XNOR2_X1 U4180 ( .A(n3361), .B(n3359), .ZN(n3330) );
  INV_X1 U4181 ( .A(n4294), .ZN(n6559) );
  NAND2_X1 U4182 ( .A1(n3650), .A2(n4473), .ZN(n3336) );
  OAI21_X1 U4183 ( .B1(n3330), .B2(n6559), .A(n3336), .ZN(n3331) );
  AOI21_X1 U4184 ( .B1(n4456), .B2(n3441), .A(n3331), .ZN(n6187) );
  NAND2_X1 U4185 ( .A1(n3332), .A2(n3334), .ZN(n3335) );
  MUX2_X2 U4186 ( .A(n3335), .B(n3334), .S(n3333), .Z(n4837) );
  OAI21_X1 U4187 ( .B1(n6559), .B2(n3346), .A(n3336), .ZN(n3337) );
  INV_X1 U4188 ( .A(n3337), .ZN(n3338) );
  NAND2_X1 U4189 ( .A1(n4349), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n3339)
         );
  INV_X1 U4190 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4413) );
  NAND2_X1 U4191 ( .A1(n3339), .A2(n4413), .ZN(n3341) );
  AND2_X1 U4192 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n3340) );
  NAND2_X1 U4193 ( .A1(n4349), .A2(n3340), .ZN(n3352) );
  AND2_X1 U4194 ( .A1(n3341), .A2(n3352), .ZN(n4406) );
  NAND2_X1 U4195 ( .A1(n4417), .A2(n3441), .ZN(n3351) );
  XNOR2_X1 U4196 ( .A(n3347), .B(n3346), .ZN(n3348) );
  OAI211_X1 U4197 ( .C1(n3348), .C2(n6559), .A(n3492), .B(n4481), .ZN(n3349)
         );
  INV_X1 U4198 ( .A(n3349), .ZN(n3350) );
  NAND2_X1 U4199 ( .A1(n3351), .A2(n3350), .ZN(n4407) );
  NAND2_X1 U4200 ( .A1(n4406), .A2(n4407), .ZN(n3353) );
  NAND2_X1 U4201 ( .A1(n3353), .A2(n3352), .ZN(n6188) );
  NAND2_X1 U4202 ( .A1(n6188), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3354)
         );
  NAND2_X1 U4203 ( .A1(n6187), .A2(n3354), .ZN(n3356) );
  OR2_X1 U4204 ( .A1(n6188), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3355)
         );
  AND2_X1 U4205 ( .A1(n3356), .A2(n3355), .ZN(n4725) );
  INV_X1 U4206 ( .A(n3376), .ZN(n3358) );
  NAND2_X1 U4207 ( .A1(n3366), .A2(n4457), .ZN(n3357) );
  INV_X1 U4208 ( .A(n3359), .ZN(n3360) );
  NAND2_X1 U4209 ( .A1(n3361), .A2(n3360), .ZN(n3369) );
  XNOR2_X1 U4210 ( .A(n3369), .B(n3368), .ZN(n3362) );
  INV_X1 U4211 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n6272) );
  NAND2_X1 U4212 ( .A1(n4725), .A2(n4726), .ZN(n4724) );
  NAND2_X1 U4213 ( .A1(n3363), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n3364)
         );
  NAND2_X1 U4214 ( .A1(n4724), .A2(n3364), .ZN(n6180) );
  OR2_X1 U4215 ( .A1(n3366), .A2(n3365), .ZN(n3367) );
  NAND2_X1 U4216 ( .A1(n3723), .A2(n3441), .ZN(n3372) );
  NAND2_X1 U4217 ( .A1(n3369), .A2(n3368), .ZN(n3393) );
  XNOR2_X1 U4218 ( .A(n3393), .B(n3391), .ZN(n3370) );
  NAND2_X1 U4219 ( .A1(n3370), .A2(n4294), .ZN(n3371) );
  NAND2_X1 U4220 ( .A1(n3372), .A2(n3371), .ZN(n3373) );
  INV_X1 U4221 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n6646) );
  XNOR2_X1 U4222 ( .A(n3373), .B(n6646), .ZN(n6179) );
  NAND2_X1 U4223 ( .A1(n6180), .A2(n6179), .ZN(n6178) );
  NAND2_X1 U4224 ( .A1(n3373), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n3374)
         );
  NAND2_X1 U4225 ( .A1(n6178), .A2(n3374), .ZN(n4707) );
  NAND2_X1 U4226 ( .A1(n3376), .A2(n3375), .ZN(n3378) );
  XNOR2_X1 U4227 ( .A(n3378), .B(n3377), .ZN(n3773) );
  NAND2_X1 U4228 ( .A1(n3773), .A2(n3441), .ZN(n3383) );
  INV_X1 U4229 ( .A(n3391), .ZN(n3379) );
  OR2_X1 U4230 ( .A1(n3393), .A2(n3379), .ZN(n3380) );
  XNOR2_X1 U4231 ( .A(n3380), .B(n3390), .ZN(n3381) );
  NAND2_X1 U4232 ( .A1(n3381), .A2(n4294), .ZN(n3382) );
  NAND2_X1 U4233 ( .A1(n3383), .A2(n3382), .ZN(n3384) );
  INV_X1 U4234 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4713) );
  XNOR2_X1 U4235 ( .A(n3384), .B(n4713), .ZN(n4706) );
  NAND2_X1 U4236 ( .A1(n4707), .A2(n4706), .ZN(n4705) );
  NAND2_X1 U4237 ( .A1(n3384), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n3385)
         );
  NAND2_X1 U4238 ( .A1(n4705), .A2(n3385), .ZN(n6172) );
  INV_X1 U4239 ( .A(n3386), .ZN(n3389) );
  INV_X1 U4240 ( .A(n3387), .ZN(n3388) );
  NAND3_X1 U4241 ( .A1(n3400), .A2(n3441), .A3(n3749), .ZN(n3396) );
  NAND2_X1 U4242 ( .A1(n3391), .A2(n3390), .ZN(n3392) );
  OR2_X1 U4243 ( .A1(n3393), .A2(n3392), .ZN(n3401) );
  XNOR2_X1 U4244 ( .A(n3401), .B(n3402), .ZN(n3394) );
  NAND2_X1 U4245 ( .A1(n3394), .A2(n4294), .ZN(n3395) );
  NAND2_X1 U4246 ( .A1(n3396), .A2(n3395), .ZN(n3397) );
  INV_X1 U4247 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n6254) );
  XNOR2_X1 U4248 ( .A(n3397), .B(n6254), .ZN(n6171) );
  NAND2_X1 U4249 ( .A1(n6172), .A2(n6171), .ZN(n6170) );
  NAND2_X1 U4250 ( .A1(n3397), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n3398)
         );
  NAND2_X1 U4251 ( .A1(n6170), .A2(n3398), .ZN(n5029) );
  AOI22_X1 U4252 ( .A1(n3475), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n3483), 
        .B2(n3410), .ZN(n3399) );
  XNOR2_X1 U4253 ( .A(n3400), .B(n3399), .ZN(n3736) );
  OR2_X1 U4254 ( .A1(n3736), .A2(n3465), .ZN(n3406) );
  INV_X1 U4255 ( .A(n3401), .ZN(n3403) );
  NAND2_X1 U4256 ( .A1(n3403), .A2(n3402), .ZN(n3409) );
  XNOR2_X1 U4257 ( .A(n3409), .B(n3410), .ZN(n3404) );
  NAND2_X1 U4258 ( .A1(n3404), .A2(n4294), .ZN(n3405) );
  NAND2_X1 U4259 ( .A1(n3406), .A2(n3405), .ZN(n3407) );
  INV_X1 U4260 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n6598) );
  XNOR2_X1 U4261 ( .A(n3407), .B(n6598), .ZN(n5028) );
  NAND2_X1 U4262 ( .A1(n5029), .A2(n5028), .ZN(n5027) );
  NAND2_X1 U4263 ( .A1(n3407), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n3408)
         );
  NAND2_X1 U4264 ( .A1(n5027), .A2(n3408), .ZN(n5084) );
  INV_X1 U4265 ( .A(n3409), .ZN(n3411) );
  NAND3_X1 U4266 ( .A1(n3411), .A2(n4294), .A3(n3410), .ZN(n3412) );
  NAND2_X1 U4267 ( .A1(n2963), .A2(n3412), .ZN(n3414) );
  INV_X1 U4268 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n3413) );
  XNOR2_X1 U4269 ( .A(n3414), .B(n3413), .ZN(n5083) );
  NAND2_X1 U4270 ( .A1(n5084), .A2(n5083), .ZN(n5082) );
  NAND2_X1 U4271 ( .A1(n3414), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n3415)
         );
  NAND2_X1 U4272 ( .A1(n5082), .A2(n3415), .ZN(n5242) );
  INV_X1 U4273 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n6225) );
  NAND2_X1 U4274 ( .A1(n2963), .A2(n6225), .ZN(n5239) );
  NAND2_X1 U4275 ( .A1(n5242), .A2(n5239), .ZN(n3416) );
  NAND2_X1 U4276 ( .A1(n3416), .A2(n5240), .ZN(n6157) );
  INV_X1 U4277 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n6202) );
  INV_X1 U4278 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n3418) );
  NAND2_X1 U4279 ( .A1(n2963), .A2(n3418), .ZN(n6156) );
  AND2_X1 U4280 ( .A1(n2972), .A2(n6156), .ZN(n3417) );
  NAND2_X1 U4281 ( .A1(n6157), .A2(n3417), .ZN(n3421) );
  NAND2_X1 U4282 ( .A1(n3421), .A2(n3420), .ZN(n5575) );
  INV_X1 U4283 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n5772) );
  NOR2_X1 U4284 ( .A1(n6160), .A2(n5772), .ZN(n5624) );
  NAND2_X1 U4285 ( .A1(n2963), .A2(n5950), .ZN(n3426) );
  INV_X1 U4286 ( .A(n3426), .ZN(n3422) );
  XNOR2_X1 U4287 ( .A(n2963), .B(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5616)
         );
  INV_X1 U4288 ( .A(n5604), .ZN(n3423) );
  INV_X1 U4289 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5606) );
  INV_X1 U4290 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5744) );
  NOR2_X1 U4291 ( .A1(n5575), .A2(n3425), .ZN(n3429) );
  NAND2_X1 U4292 ( .A1(n2963), .A2(n5772), .ZN(n5625) );
  INV_X1 U4293 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5579) );
  NAND2_X1 U4294 ( .A1(n2963), .A2(n5744), .ZN(n5585) );
  AND2_X1 U4295 ( .A1(n2969), .A2(n5585), .ZN(n3427) );
  NAND2_X1 U4296 ( .A1(n5577), .A2(n3427), .ZN(n3428) );
  NOR2_X1 U4297 ( .A1(n3429), .A2(n3428), .ZN(n5574) );
  AND2_X1 U4298 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n3660) );
  OR2_X1 U4299 ( .A1(n2967), .A2(n3660), .ZN(n3430) );
  NAND2_X1 U4300 ( .A1(n5574), .A2(n3430), .ZN(n3433) );
  NOR3_X1 U4301 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_18__SCAN_IN), .A3(INSTADDRPOINTER_REG_16__SCAN_IN), 
        .ZN(n3431) );
  NAND2_X2 U4302 ( .A1(n3433), .A2(n3432), .ZN(n5570) );
  AND2_X1 U4303 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n3661) );
  NAND2_X1 U4304 ( .A1(INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5683) );
  NAND2_X1 U4305 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n3676) );
  NOR2_X1 U4306 ( .A1(n5683), .A2(n3676), .ZN(n3663) );
  NAND3_X1 U4307 ( .A1(n5570), .A2(n3661), .A3(n3663), .ZN(n3436) );
  OR4_X1 U4308 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .A3(INSTADDRPOINTER_REG_22__SCAN_IN), 
        .A4(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n3434) );
  NAND2_X1 U4309 ( .A1(n3436), .A2(n3435), .ZN(n5529) );
  XOR2_X1 U4310 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .B(n2963), .Z(n5530) );
  INV_X1 U4311 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n3618) );
  NOR2_X1 U4312 ( .A1(n2967), .A2(n3618), .ZN(n5519) );
  NAND2_X1 U4313 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5635) );
  NOR2_X2 U4314 ( .A1(n5501), .A2(n5635), .ZN(n5345) );
  AND2_X1 U4315 ( .A1(INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n3680) );
  INV_X1 U4316 ( .A(n5528), .ZN(n3438) );
  AND2_X1 U4317 ( .A1(n2967), .A2(n3618), .ZN(n5518) );
  NOR2_X1 U4318 ( .A1(INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5637) );
  INV_X1 U4319 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n6625) );
  NAND3_X1 U4320 ( .A1(n5518), .A2(n5637), .A3(n6625), .ZN(n5346) );
  AOI21_X1 U4321 ( .B1(n5345), .B2(n3680), .A(n3439), .ZN(n3440) );
  INV_X1 U4322 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n4326) );
  XNOR2_X1 U4323 ( .A(n3440), .B(n4326), .ZN(n5344) );
  XNOR2_X1 U4324 ( .A(n4607), .B(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3455)
         );
  XOR2_X1 U4325 ( .A(n3455), .B(n3456), .Z(n3501) );
  INV_X1 U4326 ( .A(n3483), .ZN(n3442) );
  OAI21_X1 U4327 ( .B1(n3442), .B2(n3509), .A(n4481), .ZN(n3452) );
  AND2_X1 U4328 ( .A1(n3509), .A2(n4481), .ZN(n3443) );
  NOR2_X1 U4329 ( .A1(n3154), .A2(n3443), .ZN(n3467) );
  INV_X1 U4330 ( .A(n3456), .ZN(n3445) );
  NAND2_X1 U4331 ( .A1(n6400), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n3444) );
  NAND2_X1 U4332 ( .A1(n3445), .A2(n3444), .ZN(n3447) );
  OAI21_X1 U4333 ( .B1(n3520), .B2(n3447), .A(n3446), .ZN(n3450) );
  INV_X1 U4334 ( .A(n3447), .ZN(n3448) );
  NAND2_X1 U4335 ( .A1(n3483), .A2(n3448), .ZN(n3449) );
  AOI22_X1 U4336 ( .A1(n3467), .A2(n3450), .B1(n3487), .B2(n3449), .ZN(n3451)
         );
  OAI21_X1 U4337 ( .B1(n3501), .B2(n3452), .A(n3451), .ZN(n3454) );
  NAND3_X1 U4338 ( .A1(n3452), .A2(STATE2_REG_0__SCAN_IN), .A3(n3501), .ZN(
        n3453) );
  OAI211_X1 U4339 ( .C1(n3501), .C2(n3487), .A(n3454), .B(n3453), .ZN(n3470)
         );
  NAND2_X1 U4340 ( .A1(n3456), .A2(n3455), .ZN(n3458) );
  NAND2_X1 U4341 ( .A1(n6612), .A2(n4607), .ZN(n3457) );
  NAND2_X1 U4342 ( .A1(n3458), .A2(n3457), .ZN(n3462) );
  XNOR2_X1 U4343 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3461) );
  INV_X1 U4344 ( .A(n3461), .ZN(n3459) );
  XNOR2_X1 U4345 ( .A(n3462), .B(n3459), .ZN(n3500) );
  NAND2_X1 U4346 ( .A1(n3483), .A2(n3500), .ZN(n3466) );
  OAI211_X1 U4347 ( .C1(n3460), .C2(n3500), .A(n3467), .B(n3466), .ZN(n3469)
         );
  XNOR2_X1 U4348 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3471) );
  NAND2_X1 U4349 ( .A1(n3462), .A2(n3461), .ZN(n3464) );
  NAND2_X1 U4350 ( .A1(n4830), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3463) );
  NAND2_X1 U4351 ( .A1(n3464), .A2(n3463), .ZN(n3472) );
  XOR2_X1 U4352 ( .A(n3471), .B(n3472), .Z(n3499) );
  OAI22_X1 U4353 ( .A1(n3467), .A2(n3466), .B1(n3499), .B2(n3465), .ZN(n3468)
         );
  AOI21_X1 U4354 ( .B1(n3470), .B2(n3469), .A(n3468), .ZN(n3477) );
  NAND2_X1 U4355 ( .A1(n3472), .A2(n3471), .ZN(n3474) );
  NAND2_X1 U4356 ( .A1(n6419), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3473) );
  NAND2_X1 U4357 ( .A1(n3474), .A2(n3473), .ZN(n3480) );
  NAND2_X1 U4358 ( .A1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n5963), .ZN(n3481) );
  OR2_X1 U4359 ( .A1(n3480), .A2(n3481), .ZN(n3502) );
  AOI21_X1 U4360 ( .B1(n3499), .B2(n3502), .A(n3475), .ZN(n3476) );
  OAI22_X1 U4361 ( .A1(n3477), .A2(n3476), .B1(n3487), .B2(n3502), .ZN(n3478)
         );
  AOI21_X1 U4362 ( .B1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n6443), .A(n3478), 
        .ZN(n3485) );
  INV_X1 U4363 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n6417) );
  AND2_X1 U4364 ( .A1(n6417), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n3479)
         );
  OR2_X1 U4365 ( .A1(n3480), .A2(n3479), .ZN(n3482) );
  NAND2_X1 U4366 ( .A1(n3483), .A2(n3504), .ZN(n3484) );
  NAND2_X1 U4367 ( .A1(n3485), .A2(n3484), .ZN(n3489) );
  INV_X1 U4368 ( .A(n3504), .ZN(n3486) );
  INV_X1 U4369 ( .A(n3887), .ZN(n6401) );
  NAND2_X1 U4370 ( .A1(n6401), .A2(n4494), .ZN(n3657) );
  INV_X1 U4371 ( .A(n4299), .ZN(n3497) );
  NAND2_X1 U4372 ( .A1(n3887), .A2(n3650), .ZN(n3491) );
  AND3_X1 U4373 ( .A1(n3646), .A2(n3492), .A3(n3491), .ZN(n3521) );
  NAND2_X1 U4374 ( .A1(n6559), .A2(n3493), .ZN(n3494) );
  NAND2_X1 U4375 ( .A1(n3495), .A2(n3494), .ZN(n3645) );
  NAND2_X1 U4376 ( .A1(n3521), .A2(n3645), .ZN(n3496) );
  NAND2_X1 U4377 ( .A1(n3497), .A2(n3496), .ZN(n4318) );
  INV_X1 U4378 ( .A(STATE_REG_0__SCAN_IN), .ZN(n6466) );
  NAND2_X1 U4379 ( .A1(n3498), .A2(n6466), .ZN(n6461) );
  INV_X1 U4380 ( .A(n6461), .ZN(n4313) );
  AND3_X1 U4381 ( .A1(n3501), .A2(n3500), .A3(n3499), .ZN(n3503) );
  OAI21_X1 U4382 ( .B1(n3504), .B2(n3503), .A(n3502), .ZN(n4297) );
  INV_X1 U4383 ( .A(READY_N), .ZN(n6554) );
  AND2_X1 U4384 ( .A1(n4297), .A2(n6554), .ZN(n4321) );
  OAI211_X1 U4385 ( .C1(n3509), .C2(n4313), .A(n3124), .B(n4321), .ZN(n3505)
         );
  OAI211_X1 U4386 ( .C1(n4320), .C2(n3657), .A(n4318), .B(n3505), .ZN(n3507)
         );
  AND2_X1 U4387 ( .A1(n3506), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6440) );
  NAND2_X1 U4388 ( .A1(n3507), .A2(n6440), .ZN(n3515) );
  NAND2_X1 U4389 ( .A1(n3509), .A2(n6461), .ZN(n4268) );
  NAND3_X1 U4390 ( .A1(n4334), .A2(n6554), .A3(n4268), .ZN(n3510) );
  NAND3_X1 U4391 ( .A1(n3510), .A2(n4467), .A3(n5249), .ZN(n3512) );
  NAND2_X1 U4392 ( .A1(n3512), .A2(n3511), .ZN(n3513) );
  OR2_X1 U4393 ( .A1(n4308), .A2(n3513), .ZN(n3514) );
  AND2_X1 U4394 ( .A1(n3521), .A2(n3154), .ZN(n4319) );
  INV_X1 U4395 ( .A(n4319), .ZN(n4327) );
  INV_X4 U4396 ( .A(n3539), .ZN(n4409) );
  INV_X1 U4397 ( .A(n3638), .ZN(n3519) );
  AOI22_X1 U4398 ( .A1(n4334), .A2(n4409), .B1(n3519), .B2(n4486), .ZN(n3522)
         );
  NAND2_X1 U4399 ( .A1(n3521), .A2(n3520), .ZN(n6396) );
  NAND4_X1 U4400 ( .A1(n4336), .A2(n4327), .A3(n3522), .A4(n6396), .ZN(n3523)
         );
  NAND2_X1 U4401 ( .A1(n3669), .A2(n3523), .ZN(n5780) );
  INV_X1 U4402 ( .A(EBX_REG_1__SCAN_IN), .ZN(n3525) );
  NAND2_X1 U4403 ( .A1(n3551), .A2(n3525), .ZN(n3529) );
  INV_X1 U4404 ( .A(n4473), .ZN(n3524) );
  NAND2_X1 U4405 ( .A1(n3524), .A2(n4467), .ZN(n3537) );
  NAND2_X1 U4406 ( .A1(n3537), .A2(n4413), .ZN(n3527) );
  INV_X4 U4407 ( .A(n5261), .ZN(n5319) );
  NAND2_X1 U4408 ( .A1(n4409), .A2(n3525), .ZN(n3526) );
  NAND3_X1 U4409 ( .A1(n3527), .A2(n5319), .A3(n3526), .ZN(n3528) );
  NAND2_X1 U4410 ( .A1(n3529), .A2(n3528), .ZN(n3531) );
  NAND2_X1 U4411 ( .A1(n3537), .A2(EBX_REG_0__SCAN_IN), .ZN(n3530) );
  OAI21_X1 U4412 ( .B1(n5261), .B2(EBX_REG_0__SCAN_IN), .A(n3530), .ZN(n4350)
         );
  XNOR2_X1 U4413 ( .A(n3531), .B(n4350), .ZN(n4410) );
  NAND2_X1 U4414 ( .A1(n4410), .A2(n4409), .ZN(n4411) );
  NAND2_X1 U4415 ( .A1(n4411), .A2(n3531), .ZN(n4449) );
  NAND2_X2 U4416 ( .A1(n5319), .A2(n4409), .ZN(n3632) );
  MUX2_X1 U4417 ( .A(n3632), .B(n5319), .S(EBX_REG_3__SCAN_IN), .Z(n3533) );
  NAND2_X1 U4418 ( .A1(n6272), .A2(n3641), .ZN(n3532) );
  INV_X1 U4419 ( .A(n3537), .ZN(n3538) );
  NAND2_X1 U4420 ( .A1(n3538), .A2(n2964), .ZN(n3607) );
  NAND2_X1 U4421 ( .A1(n2964), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3540)
         );
  AND2_X1 U4422 ( .A1(n3607), .A2(n3540), .ZN(n3541) );
  NAND2_X1 U4423 ( .A1(n4450), .A2(n4451), .ZN(n3543) );
  MUX2_X1 U4424 ( .A(n3622), .B(n3626), .S(EBX_REG_4__SCAN_IN), .Z(n3546) );
  NAND2_X1 U4425 ( .A1(n2964), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n3544)
         );
  AND2_X1 U4426 ( .A1(n3607), .A2(n3544), .ZN(n3545) );
  NAND2_X1 U4427 ( .A1(n3546), .A2(n3545), .ZN(n4576) );
  NAND2_X1 U4428 ( .A1(n4713), .A2(n3641), .ZN(n3548) );
  MUX2_X1 U4429 ( .A(n3632), .B(n5319), .S(EBX_REG_5__SCAN_IN), .Z(n3547) );
  NAND2_X1 U4430 ( .A1(n3548), .A2(n3547), .ZN(n4716) );
  INV_X1 U4431 ( .A(EBX_REG_6__SCAN_IN), .ZN(n5200) );
  NAND2_X1 U4432 ( .A1(n3625), .A2(n5200), .ZN(n3555) );
  NAND2_X1 U4433 ( .A1(n3626), .A2(n6254), .ZN(n3553) );
  NAND2_X1 U4434 ( .A1(n4409), .A2(n5200), .ZN(n3552) );
  NAND3_X1 U4435 ( .A1(n3553), .A2(n5319), .A3(n3552), .ZN(n3554) );
  OR2_X2 U4436 ( .A1(n5195), .A2(n5196), .ZN(n5197) );
  NAND2_X1 U4437 ( .A1(n6598), .A2(n3641), .ZN(n3557) );
  MUX2_X1 U4438 ( .A(n3632), .B(n5319), .S(EBX_REG_7__SCAN_IN), .Z(n3556) );
  NAND2_X1 U4439 ( .A1(n3557), .A2(n3556), .ZN(n5038) );
  MUX2_X1 U4440 ( .A(n3622), .B(n3626), .S(EBX_REG_8__SCAN_IN), .Z(n3560) );
  NAND2_X1 U4441 ( .A1(n2964), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n3558)
         );
  AND2_X1 U4442 ( .A1(n3607), .A2(n3558), .ZN(n3559) );
  NAND2_X1 U4443 ( .A1(n3560), .A2(n3559), .ZN(n5058) );
  NAND2_X1 U4444 ( .A1(n5059), .A2(n5058), .ZN(n5061) );
  NAND2_X1 U4445 ( .A1(n6225), .A2(n3641), .ZN(n3562) );
  MUX2_X1 U4446 ( .A(n3632), .B(n5319), .S(EBX_REG_9__SCAN_IN), .Z(n3561) );
  NAND2_X1 U4447 ( .A1(n3562), .A2(n3561), .ZN(n5046) );
  MUX2_X1 U4448 ( .A(n3622), .B(n3626), .S(EBX_REG_10__SCAN_IN), .Z(n3566) );
  NAND2_X1 U4449 ( .A1(n2964), .A2(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n3565) );
  NOR2_X2 U4450 ( .A1(n5190), .A2(n5189), .ZN(n6013) );
  INV_X1 U4451 ( .A(EBX_REG_11__SCAN_IN), .ZN(n6097) );
  NAND2_X1 U4452 ( .A1(n3602), .A2(n6097), .ZN(n3569) );
  NAND2_X1 U4453 ( .A1(n4409), .A2(n6097), .ZN(n3567) );
  OAI211_X1 U4454 ( .C1(n5261), .C2(n6202), .A(n3567), .B(n3626), .ZN(n3568)
         );
  AND2_X1 U4455 ( .A1(n3569), .A2(n3568), .ZN(n6012) );
  AND2_X2 U4456 ( .A1(n6013), .A2(n6012), .ZN(n6015) );
  MUX2_X1 U4457 ( .A(n3622), .B(n3626), .S(EBX_REG_12__SCAN_IN), .Z(n3572) );
  NAND2_X1 U4458 ( .A1(n2964), .A2(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n3570) );
  AND2_X1 U4459 ( .A1(n3607), .A2(n3570), .ZN(n3571) );
  NAND2_X1 U4460 ( .A1(n3572), .A2(n3571), .ZN(n5430) );
  NAND2_X1 U4461 ( .A1(n6015), .A2(n5430), .ZN(n4666) );
  INV_X1 U4462 ( .A(EBX_REG_13__SCAN_IN), .ZN(n3573) );
  NAND2_X1 U4463 ( .A1(n3602), .A2(n3573), .ZN(n3576) );
  INV_X1 U4464 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5950) );
  NAND2_X1 U4465 ( .A1(n4409), .A2(n3573), .ZN(n3574) );
  OAI211_X1 U4466 ( .C1(n5261), .C2(n5950), .A(n3574), .B(n3626), .ZN(n3575)
         );
  NAND2_X1 U4467 ( .A1(n3576), .A2(n3575), .ZN(n4668) );
  MUX2_X1 U4468 ( .A(n3622), .B(n3626), .S(EBX_REG_14__SCAN_IN), .Z(n3580) );
  NAND2_X1 U4469 ( .A1(n2964), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n3579) );
  AND3_X1 U4470 ( .A1(n3580), .A2(n3607), .A3(n3579), .ZN(n5048) );
  INV_X1 U4471 ( .A(EBX_REG_15__SCAN_IN), .ZN(n5036) );
  NAND2_X1 U4472 ( .A1(n3602), .A2(n5036), .ZN(n3583) );
  NAND2_X1 U4473 ( .A1(n4409), .A2(n5036), .ZN(n3581) );
  OAI211_X1 U4474 ( .C1(n5261), .C2(n5744), .A(n3581), .B(n3626), .ZN(n3582)
         );
  NAND2_X1 U4475 ( .A1(n3583), .A2(n3582), .ZN(n5034) );
  MUX2_X1 U4476 ( .A(n3622), .B(n3626), .S(EBX_REG_16__SCAN_IN), .Z(n3586) );
  NAND2_X1 U4477 ( .A1(n2964), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n3584) );
  AND2_X1 U4478 ( .A1(n3607), .A2(n3584), .ZN(n3585) );
  NAND2_X1 U4479 ( .A1(n3586), .A2(n3585), .ZN(n5063) );
  NAND2_X1 U4480 ( .A1(n5064), .A2(n5063), .ZN(n5062) );
  INV_X1 U4481 ( .A(EBX_REG_17__SCAN_IN), .ZN(n6090) );
  NAND2_X1 U4482 ( .A1(n3602), .A2(n6090), .ZN(n3589) );
  INV_X1 U4483 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5948) );
  NAND2_X1 U4484 ( .A1(n4409), .A2(n6090), .ZN(n3587) );
  OAI211_X1 U4485 ( .C1(n5261), .C2(n5948), .A(n3587), .B(n3626), .ZN(n3588)
         );
  NAND2_X1 U4486 ( .A1(n3589), .A2(n3588), .ZN(n5941) );
  INV_X1 U4487 ( .A(EBX_REG_19__SCAN_IN), .ZN(n5901) );
  NAND2_X1 U4488 ( .A1(n3625), .A2(n5901), .ZN(n3593) );
  INV_X1 U4489 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n6641) );
  NAND2_X1 U4490 ( .A1(n3626), .A2(n6641), .ZN(n3591) );
  NAND2_X1 U4491 ( .A1(n4409), .A2(n5901), .ZN(n3590) );
  NAND3_X1 U4492 ( .A1(n3591), .A2(n5319), .A3(n3590), .ZN(n3592) );
  AND2_X1 U4493 ( .A1(n3593), .A2(n3592), .ZN(n5307) );
  INV_X1 U4494 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n3685) );
  NOR2_X1 U4495 ( .A1(n2964), .A2(EBX_REG_20__SCAN_IN), .ZN(n3594) );
  AOI21_X1 U4496 ( .B1(n3641), .B2(n3685), .A(n3594), .ZN(n5320) );
  INV_X1 U4497 ( .A(n3641), .ZN(n4351) );
  OR2_X1 U4498 ( .A1(n4351), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n3595)
         );
  INV_X1 U4499 ( .A(EBX_REG_18__SCAN_IN), .ZN(n5991) );
  NAND2_X1 U4500 ( .A1(n4409), .A2(n5991), .ZN(n5262) );
  NAND2_X1 U4501 ( .A1(n3595), .A2(n5262), .ZN(n5318) );
  NAND2_X1 U4502 ( .A1(n5261), .A2(EBX_REG_20__SCAN_IN), .ZN(n3597) );
  NAND2_X1 U4503 ( .A1(n5318), .A2(n5319), .ZN(n3596) );
  OAI211_X1 U4504 ( .C1(n5320), .C2(n5318), .A(n3597), .B(n3596), .ZN(n3598)
         );
  INV_X1 U4505 ( .A(n3598), .ZN(n3599) );
  MUX2_X1 U4506 ( .A(n3602), .B(n5261), .S(EBX_REG_21__SCAN_IN), .Z(n3601) );
  NOR2_X1 U4507 ( .A1(n4351), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n3600)
         );
  NOR2_X1 U4508 ( .A1(n3601), .A2(n3600), .ZN(n5467) );
  NAND2_X1 U4509 ( .A1(n5468), .A2(n5467), .ZN(n5461) );
  INV_X1 U4510 ( .A(EBX_REG_23__SCAN_IN), .ZN(n6657) );
  NAND2_X1 U4511 ( .A1(n3602), .A2(n6657), .ZN(n3605) );
  INV_X1 U4512 ( .A(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5669) );
  NAND2_X1 U4513 ( .A1(n4409), .A2(n6657), .ZN(n3603) );
  OAI211_X1 U4514 ( .C1(n5261), .C2(n5669), .A(n3603), .B(n3626), .ZN(n3604)
         );
  AND2_X1 U4515 ( .A1(n3605), .A2(n3604), .ZN(n5676) );
  MUX2_X1 U4516 ( .A(n3622), .B(n3626), .S(EBX_REG_22__SCAN_IN), .Z(n3609) );
  NAND2_X1 U4517 ( .A1(n2964), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n3606) );
  AND2_X1 U4518 ( .A1(n3607), .A2(n3606), .ZN(n3608) );
  NAND2_X1 U4519 ( .A1(n3609), .A2(n3608), .ZN(n5675) );
  NAND2_X1 U4520 ( .A1(n5676), .A2(n5675), .ZN(n3610) );
  OR2_X2 U4521 ( .A1(n5461), .A2(n3610), .ZN(n5680) );
  INV_X1 U4522 ( .A(EBX_REG_24__SCAN_IN), .ZN(n5458) );
  NAND2_X1 U4523 ( .A1(n3625), .A2(n5458), .ZN(n3615) );
  INV_X1 U4524 ( .A(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n3611) );
  NAND2_X1 U4525 ( .A1(n3626), .A2(n3611), .ZN(n3613) );
  NAND2_X1 U4526 ( .A1(n4409), .A2(n5458), .ZN(n3612) );
  NAND3_X1 U4527 ( .A1(n3613), .A2(n5319), .A3(n3612), .ZN(n3614) );
  AND2_X1 U4528 ( .A1(n3615), .A2(n3614), .ZN(n5455) );
  MUX2_X1 U4529 ( .A(n3632), .B(n5319), .S(EBX_REG_25__SCAN_IN), .Z(n3617) );
  NAND2_X1 U4530 ( .A1(n3641), .A2(n5659), .ZN(n3616) );
  AND2_X1 U4531 ( .A1(n3617), .A2(n3616), .ZN(n5415) );
  NAND2_X1 U4532 ( .A1(n3626), .A2(n3618), .ZN(n3620) );
  INV_X1 U4533 ( .A(EBX_REG_26__SCAN_IN), .ZN(n6732) );
  NAND2_X1 U4534 ( .A1(n4409), .A2(n6732), .ZN(n3619) );
  NAND3_X1 U4535 ( .A1(n3620), .A2(n5319), .A3(n3619), .ZN(n3621) );
  OAI21_X1 U4536 ( .B1(n3622), .B2(EBX_REG_26__SCAN_IN), .A(n3621), .ZN(n5404)
         );
  NAND2_X1 U4537 ( .A1(n5417), .A2(n5404), .ZN(n5403) );
  MUX2_X1 U4538 ( .A(n3632), .B(n5319), .S(EBX_REG_27__SCAN_IN), .Z(n3623) );
  OAI21_X1 U4539 ( .B1(INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n4351), .A(n3623), 
        .ZN(n5448) );
  OR2_X2 U4540 ( .A1(n5403), .A2(n5448), .ZN(n5445) );
  INV_X1 U4541 ( .A(EBX_REG_28__SCAN_IN), .ZN(n3624) );
  NAND2_X1 U4542 ( .A1(n3625), .A2(n3624), .ZN(n3629) );
  INV_X1 U4543 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5505) );
  NAND2_X1 U4544 ( .A1(n3626), .A2(n5505), .ZN(n3627) );
  OAI211_X1 U4545 ( .C1(EBX_REG_28__SCAN_IN), .C2(n2964), .A(n3627), .B(n5319), 
        .ZN(n3628) );
  AND2_X1 U4546 ( .A1(n3629), .A2(n3628), .ZN(n5393) );
  NOR2_X4 U4547 ( .A1(n5445), .A2(n5393), .ZN(n5392) );
  AOI22_X1 U4548 ( .A1(n4351), .A2(EBX_REG_30__SCAN_IN), .B1(
        INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n2964), .ZN(n4252) );
  MUX2_X1 U4549 ( .A(EBX_REG_29__SCAN_IN), .B(n2978), .S(n5319), .Z(n3634) );
  NOR2_X1 U4550 ( .A1(n3632), .A2(EBX_REG_29__SCAN_IN), .ZN(n3633) );
  NOR2_X1 U4551 ( .A1(n3634), .A2(n3633), .ZN(n5326) );
  NAND3_X1 U4552 ( .A1(n5392), .A2(n4252), .A3(n5326), .ZN(n3635) );
  NAND2_X1 U4553 ( .A1(n4256), .A2(n3635), .ZN(n3637) );
  OAI22_X1 U4554 ( .A1(n4351), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        EBX_REG_31__SCAN_IN), .B2(n2964), .ZN(n3636) );
  XNOR2_X2 U4555 ( .A(n3637), .B(n3636), .ZN(n5383) );
  INV_X1 U4556 ( .A(n5383), .ZN(n3667) );
  NAND2_X1 U4557 ( .A1(n4334), .A2(n4294), .ZN(n6427) );
  OAI21_X1 U4558 ( .B1(n3638), .B2(n4486), .A(n6427), .ZN(n3639) );
  NAND2_X1 U4559 ( .A1(n3669), .A2(n3639), .ZN(n6249) );
  NOR2_X1 U4560 ( .A1(STATE2_REG_0__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n6454) );
  INV_X1 U4561 ( .A(n6454), .ZN(n3640) );
  OR2_X1 U4562 ( .A1(n6542), .A2(n3640), .ZN(n6248) );
  INV_X1 U4563 ( .A(REIP_REG_31__SCAN_IN), .ZN(n6524) );
  NOR2_X1 U4564 ( .A1(n6248), .A2(n6524), .ZN(n5339) );
  NAND2_X1 U4565 ( .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n5755) );
  NOR2_X1 U4566 ( .A1(n5950), .A2(n5755), .ZN(n5761) );
  NAND2_X1 U4567 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n5761), .ZN(n5743) );
  NAND2_X1 U4568 ( .A1(INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5739) );
  NOR2_X1 U4569 ( .A1(n5743), .A2(n5739), .ZN(n3671) );
  INV_X1 U4570 ( .A(n3671), .ZN(n3673) );
  OR2_X1 U4571 ( .A1(n4293), .A2(n3124), .ZN(n4317) );
  NAND2_X1 U4572 ( .A1(n3641), .A2(n4317), .ZN(n3643) );
  NAND2_X1 U4573 ( .A1(n3643), .A2(n3642), .ZN(n3647) );
  AND4_X1 U4574 ( .A1(n3647), .A2(n3646), .A3(n3645), .A4(n3644), .ZN(n3648)
         );
  NAND2_X1 U4575 ( .A1(n3649), .A2(n3648), .ZN(n4337) );
  AND2_X1 U4576 ( .A1(n3167), .A2(n3650), .ZN(n3651) );
  NAND2_X1 U4577 ( .A1(n6401), .A2(n3651), .ZN(n4612) );
  INV_X1 U4578 ( .A(n3652), .ZN(n3653) );
  NAND2_X1 U4579 ( .A1(n3653), .A2(n5261), .ZN(n3654) );
  OAI211_X1 U4580 ( .C1(n4332), .C2(n3655), .A(n4612), .B(n3654), .ZN(n3656)
         );
  NAND2_X1 U4581 ( .A1(n3669), .A2(n4295), .ZN(n6276) );
  INV_X1 U4582 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6275) );
  INV_X1 U4583 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n6285) );
  OAI21_X1 U4584 ( .B1(n4413), .B2(n6275), .A(n6285), .ZN(n6259) );
  NAND3_X1 U4585 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .A3(n6259), .ZN(n4712) );
  NOR2_X1 U4586 ( .A1(n4713), .A2(n4712), .ZN(n6246) );
  INV_X1 U4587 ( .A(n6246), .ZN(n4711) );
  NOR2_X1 U4588 ( .A1(n6254), .A2(n4711), .ZN(n6214) );
  NAND2_X1 U4589 ( .A1(n5771), .A2(n6214), .ZN(n6208) );
  NAND2_X1 U4590 ( .A1(INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n6227) );
  NAND2_X1 U4591 ( .A1(INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n6215) );
  OR2_X1 U4592 ( .A1(n6227), .A2(n6215), .ZN(n3659) );
  NOR2_X1 U4593 ( .A1(n6208), .A2(n3659), .ZN(n5732) );
  NAND2_X1 U4594 ( .A1(n3669), .A2(n3658), .ZN(n5754) );
  AND2_X1 U4595 ( .A1(n4299), .A2(n4494), .ZN(n6404) );
  NAND2_X1 U4596 ( .A1(n3669), .A2(n6404), .ZN(n5758) );
  NAND2_X1 U4597 ( .A1(n5754), .A2(n5758), .ZN(n6206) );
  NAND2_X1 U4598 ( .A1(n5758), .A2(n6275), .ZN(n4408) );
  NAND2_X1 U4599 ( .A1(n6206), .A2(n4408), .ZN(n6284) );
  NAND2_X1 U4600 ( .A1(INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n6261) );
  NOR2_X1 U4601 ( .A1(n6285), .A2(n4413), .ZN(n4709) );
  INV_X1 U4602 ( .A(n4709), .ZN(n6274) );
  NOR2_X1 U4603 ( .A1(n6261), .A2(n6274), .ZN(n4714) );
  NAND3_X1 U4604 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_5__SCAN_IN), .A3(n4714), .ZN(n6205) );
  OR2_X1 U4605 ( .A1(n3659), .A2(n6205), .ZN(n5733) );
  NOR2_X1 U4606 ( .A1(n6284), .A2(n5733), .ZN(n5770) );
  NOR2_X1 U4607 ( .A1(n3673), .A2(n6196), .ZN(n5940) );
  NAND2_X1 U4608 ( .A1(n5940), .A2(n3660), .ZN(n5707) );
  INV_X1 U4609 ( .A(n3661), .ZN(n3662) );
  INV_X1 U4610 ( .A(n3663), .ZN(n3664) );
  NOR2_X1 U4611 ( .A1(n5698), .A2(n3664), .ZN(n5660) );
  AND2_X1 U4612 ( .A1(INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n3679) );
  NAND2_X1 U4613 ( .A1(n5660), .A2(n3679), .ZN(n5646) );
  OR2_X1 U4614 ( .A1(n5646), .A2(n5635), .ZN(n5353) );
  INV_X1 U4615 ( .A(n3680), .ZN(n3665) );
  NOR3_X1 U4616 ( .A1(n5353), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .A3(n3665), 
        .ZN(n3666) );
  OR2_X1 U4617 ( .A1(n6206), .A2(n5771), .ZN(n6210) );
  INV_X1 U4618 ( .A(n6210), .ZN(n5735) );
  NOR2_X1 U4619 ( .A1(n3669), .A2(n3668), .ZN(n4356) );
  INV_X1 U4620 ( .A(n5754), .ZN(n3670) );
  NOR2_X1 U4621 ( .A1(n5771), .A2(n3670), .ZN(n5756) );
  NOR2_X1 U4622 ( .A1(INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n5756), .ZN(n4353)
         );
  NOR2_X1 U4623 ( .A1(n4356), .A2(n4353), .ZN(n4708) );
  NAND2_X1 U4624 ( .A1(n6276), .A2(n4708), .ZN(n6207) );
  NAND4_X1 U4625 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_17__SCAN_IN), .A3(INSTADDRPOINTER_REG_19__SCAN_IN), 
        .A4(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n3672) );
  NAND2_X1 U4626 ( .A1(n5732), .A2(n3671), .ZN(n5708) );
  AOI222_X1 U4627 ( .A1(n6207), .A2(n3672), .B1(n6207), .B2(n5708), .C1(n3672), 
        .C2(n6206), .ZN(n3674) );
  OAI21_X1 U4628 ( .B1(n5733), .B2(n3673), .A(n6206), .ZN(n5709) );
  AND2_X1 U4629 ( .A1(n3674), .A2(n5709), .ZN(n5696) );
  NAND2_X1 U4630 ( .A1(n6210), .A2(n5683), .ZN(n3675) );
  NAND2_X1 U4631 ( .A1(n5696), .A2(n3675), .ZN(n5686) );
  INV_X1 U4632 ( .A(n3676), .ZN(n3677) );
  AOI21_X1 U4633 ( .B1(n6284), .B2(n6276), .A(n3677), .ZN(n3678) );
  NOR2_X1 U4634 ( .A1(n5686), .A2(n3678), .ZN(n5651) );
  OAI21_X1 U4635 ( .B1(n5735), .B2(n3679), .A(n5651), .ZN(n5648) );
  AOI21_X1 U4636 ( .B1(n5635), .B2(n6210), .A(n5648), .ZN(n5352) );
  OAI21_X1 U4637 ( .B1(n3680), .B2(n5735), .A(n5352), .ZN(n3681) );
  NAND2_X1 U4638 ( .A1(n3681), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n3682) );
  AND2_X1 U4639 ( .A1(n3683), .A2(n3682), .ZN(n3684) );
  OAI21_X1 U4640 ( .B1(n5344), .B2(n5780), .A(n3684), .ZN(U2987) );
  OAI21_X1 U4641 ( .B1(n2967), .B2(INSTADDRPOINTER_REG_19__SCAN_IN), .A(n5570), 
        .ZN(n5549) );
  OAI21_X1 U4642 ( .B1(n6641), .B2(n6160), .A(n5549), .ZN(n5564) );
  XNOR2_X1 U4643 ( .A(n2967), .B(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5559)
         );
  INV_X1 U4644 ( .A(n5557), .ZN(n3688) );
  OAI21_X1 U4645 ( .B1(n2967), .B2(INSTADDRPOINTER_REG_21__SCAN_IN), .A(n3688), 
        .ZN(n5539) );
  NOR2_X1 U4646 ( .A1(n6160), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5537)
         );
  AOI21_X1 U4647 ( .B1(INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n6160), .A(n5537), 
        .ZN(n3689) );
  OR2_X2 U4648 ( .A1(n4308), .A2(n6396), .ZN(n6169) );
  INV_X1 U4649 ( .A(n6169), .ZN(n6191) );
  NAND2_X1 U4650 ( .A1(n5689), .A2(n6191), .ZN(n4023) );
  NAND2_X1 U4651 ( .A1(n4456), .A2(n2965), .ZN(n3692) );
  INV_X2 U4652 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n6661) );
  NAND2_X1 U4653 ( .A1(n6661), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4074) );
  NOR2_X1 U4654 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATEBS16_REG_SCAN_IN), .ZN(
        n4241) );
  INV_X1 U4656 ( .A(n5249), .ZN(n3693) );
  AND2_X1 U4657 ( .A1(n3693), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3703) );
  INV_X1 U4658 ( .A(n3703), .ZN(n3726) );
  NAND2_X1 U4659 ( .A1(n6403), .A2(n2965), .ZN(n3696) );
  AOI22_X1 U4660 ( .A1(n5336), .A2(EAX_REG_0__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n6661), .ZN(n3695) );
  OAI211_X1 U4661 ( .C1(n3726), .C2(n6400), .A(n3696), .B(n3695), .ZN(n4396)
         );
  MUX2_X1 U4662 ( .A(n4241), .B(n4397), .S(n4396), .Z(n4420) );
  AND2_X1 U4663 ( .A1(n2965), .A2(n4420), .ZN(n3697) );
  NAND2_X1 U4664 ( .A1(n4417), .A2(n3697), .ZN(n3702) );
  AOI22_X1 U4665 ( .A1(n5336), .A2(EAX_REG_1__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n6661), .ZN(n3699) );
  NAND2_X1 U4666 ( .A1(n3703), .A2(n4607), .ZN(n3698) );
  AND2_X1 U4667 ( .A1(n3699), .A2(n3698), .ZN(n4418) );
  INV_X1 U4668 ( .A(n4418), .ZN(n3700) );
  NAND2_X1 U4669 ( .A1(n3702), .A2(n3701), .ZN(n3712) );
  NAND2_X1 U4670 ( .A1(n3711), .A2(n3712), .ZN(n3710) );
  NAND2_X1 U4671 ( .A1(n3703), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3709) );
  INV_X1 U4672 ( .A(n5336), .ZN(n3704) );
  INV_X1 U4673 ( .A(PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3706) );
  INV_X1 U4674 ( .A(n4241), .ZN(n4235) );
  INV_X1 U4675 ( .A(n4235), .ZN(n4196) );
  OAI21_X1 U4676 ( .B1(PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .A(n3717), .ZN(n6194) );
  NAND2_X1 U4677 ( .A1(n4196), .A2(n6194), .ZN(n3705) );
  OAI21_X1 U4678 ( .B1(n4074), .B2(n3706), .A(n3705), .ZN(n3707) );
  AOI21_X1 U4679 ( .B1(n4237), .B2(EAX_REG_2__SCAN_IN), .A(n3707), .ZN(n3708)
         );
  AND2_X1 U4680 ( .A1(n3709), .A2(n3708), .ZN(n4438) );
  NAND2_X1 U4681 ( .A1(n3710), .A2(n4438), .ZN(n3714) );
  INV_X1 U4682 ( .A(n3711), .ZN(n4439) );
  NAND2_X1 U4683 ( .A1(n4439), .A2(n4437), .ZN(n3713) );
  NAND2_X1 U4684 ( .A1(n3714), .A2(n3713), .ZN(n4436) );
  INV_X1 U4685 ( .A(n4743), .ZN(n3722) );
  INV_X1 U4686 ( .A(n3717), .ZN(n3718) );
  INV_X1 U4687 ( .A(n3727), .ZN(n3728) );
  OAI21_X1 U4688 ( .B1(PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n3718), .A(n3728), 
        .ZN(n4727) );
  INV_X1 U4689 ( .A(n4074), .ZN(n5335) );
  AOI22_X1 U4690 ( .A1(n4196), .A2(n4727), .B1(n5335), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3720) );
  NAND2_X1 U4691 ( .A1(n4237), .A2(EAX_REG_3__SCAN_IN), .ZN(n3719) );
  OAI211_X1 U4692 ( .C1(n3726), .C2(n4617), .A(n3720), .B(n3719), .ZN(n3721)
         );
  AOI21_X1 U4693 ( .B1(n3722), .B2(n2965), .A(n3721), .ZN(n4446) );
  NOR2_X2 U4694 ( .A1(n4436), .A2(n4446), .ZN(n4447) );
  NAND2_X1 U4695 ( .A1(n3723), .A2(n2965), .ZN(n3735) );
  NAND2_X1 U4696 ( .A1(n6661), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3725)
         );
  NAND2_X1 U4697 ( .A1(n4237), .A2(EAX_REG_4__SCAN_IN), .ZN(n3724) );
  OAI211_X1 U4698 ( .C1(n3726), .C2(n5963), .A(n3725), .B(n3724), .ZN(n3733)
         );
  INV_X1 U4699 ( .A(n3769), .ZN(n3731) );
  INV_X1 U4700 ( .A(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3729) );
  NAND2_X1 U4701 ( .A1(n3729), .A2(n3728), .ZN(n3730) );
  NAND2_X1 U4702 ( .A1(n3731), .A2(n3730), .ZN(n6185) );
  AND2_X1 U4703 ( .A1(n6185), .A2(n4241), .ZN(n3732) );
  AOI21_X1 U4704 ( .B1(n3733), .B2(n4235), .A(n3732), .ZN(n3734) );
  NAND2_X1 U4705 ( .A1(n3735), .A2(n3734), .ZN(n4472) );
  NAND2_X1 U4706 ( .A1(n4447), .A2(n4472), .ZN(n4471) );
  INV_X1 U4707 ( .A(n4471), .ZN(n3836) );
  INV_X1 U4708 ( .A(n3736), .ZN(n3741) );
  INV_X1 U4709 ( .A(EAX_REG_7__SCAN_IN), .ZN(n3739) );
  XNOR2_X1 U4710 ( .A(n3750), .B(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n5070) );
  INV_X1 U4711 ( .A(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n5073) );
  NOR2_X1 U4712 ( .A1(n4074), .A2(n5073), .ZN(n3737) );
  AOI21_X1 U4713 ( .B1(n5070), .B2(n4241), .A(n3737), .ZN(n3738) );
  OAI21_X1 U4714 ( .B1(n3704), .B2(n3739), .A(n3738), .ZN(n3740) );
  NAND2_X1 U4715 ( .A1(n4237), .A2(EAX_REG_6__SCAN_IN), .ZN(n3747) );
  INV_X1 U4716 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n5973) );
  OAI21_X1 U4717 ( .B1(n5973), .B2(PHYADDRPOINTER_REG_6__SCAN_IN), .A(n6661), 
        .ZN(n3746) );
  AND2_X1 U4718 ( .A1(n3743), .A2(n3742), .ZN(n3744) );
  OR2_X1 U4719 ( .A1(n3744), .A2(n3750), .ZN(n6177) );
  NOR2_X1 U4720 ( .A1(n6177), .A2(n4235), .ZN(n3745) );
  AOI21_X1 U4721 ( .B1(n3747), .B2(n3746), .A(n3745), .ZN(n3748) );
  AOI21_X1 U4722 ( .B1(n3751), .B2(n6567), .A(n3802), .ZN(n6030) );
  OR2_X1 U4723 ( .A1(n6030), .A2(n4235), .ZN(n3766) );
  AOI22_X1 U4724 ( .A1(n3888), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4214), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3755) );
  AOI22_X1 U4725 ( .A1(n4211), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n4173), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3754) );
  AOI22_X1 U4726 ( .A1(n3961), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4156), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3753) );
  AOI22_X1 U4727 ( .A1(n4222), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4224), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3752) );
  NAND4_X1 U4728 ( .A1(n3755), .A2(n3754), .A3(n3753), .A4(n3752), .ZN(n3761)
         );
  CLKBUF_X1 U4729 ( .A(n3049), .Z(n4175) );
  AOI22_X1 U4730 ( .A1(n4175), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4219), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3759) );
  AOI22_X1 U4731 ( .A1(n3232), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4107), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3758) );
  AOI22_X1 U4732 ( .A1(n4078), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n4213), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3757) );
  AOI22_X1 U4733 ( .A1(n4225), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n4223), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3756) );
  NAND4_X1 U4734 ( .A1(n3759), .A2(n3758), .A3(n3757), .A4(n3756), .ZN(n3760)
         );
  OAI21_X1 U4735 ( .B1(n3761), .B2(n3760), .A(n2965), .ZN(n3764) );
  NAND2_X1 U4736 ( .A1(n4237), .A2(EAX_REG_9__SCAN_IN), .ZN(n3763) );
  NAND2_X1 U4737 ( .A1(n5335), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3762)
         );
  AND3_X1 U4738 ( .A1(n3764), .A2(n3763), .A3(n3762), .ZN(n3765) );
  NAND2_X1 U4739 ( .A1(n3766), .A2(n3765), .ZN(n5043) );
  INV_X1 U4740 ( .A(n5043), .ZN(n3767) );
  NOR2_X2 U4741 ( .A1(n5030), .A2(n3768), .ZN(n5428) );
  INV_X1 U4742 ( .A(EAX_REG_5__SCAN_IN), .ZN(n3771) );
  XNOR2_X1 U4743 ( .A(n3769), .B(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n5265) );
  AOI22_X1 U4744 ( .A1(n5265), .A2(n4241), .B1(n5335), .B2(
        PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3770) );
  OAI21_X1 U4745 ( .B1(n3704), .B2(n3771), .A(n3770), .ZN(n3772) );
  AOI21_X1 U4746 ( .B1(n3773), .B2(n2965), .A(n3772), .ZN(n4967) );
  INV_X1 U4747 ( .A(n4967), .ZN(n3835) );
  INV_X1 U4748 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n5437) );
  XNOR2_X1 U4749 ( .A(n3837), .B(n5437), .ZN(n5629) );
  AOI21_X1 U4750 ( .B1(STATEBS16_REG_SCAN_IN), .B2(n5437), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3775) );
  AND2_X1 U4751 ( .A1(n4237), .A2(EAX_REG_12__SCAN_IN), .ZN(n3774) );
  OAI22_X1 U4752 ( .A1(n5629), .A2(n4235), .B1(n3775), .B2(n3774), .ZN(n3787)
         );
  AOI22_X1 U4753 ( .A1(INSTQUEUE_REG_3__4__SCAN_IN), .A2(n4107), .B1(n3232), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3779) );
  AOI22_X1 U4754 ( .A1(n4078), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n4214), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3778) );
  AOI22_X1 U4755 ( .A1(n4173), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n4213), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3777) );
  AOI22_X1 U4756 ( .A1(n4175), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n4223), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3776) );
  NAND4_X1 U4757 ( .A1(n3779), .A2(n3778), .A3(n3777), .A4(n3776), .ZN(n3785)
         );
  AOI22_X1 U4758 ( .A1(n2962), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4211), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3783) );
  AOI22_X1 U4759 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n3961), .B1(n4156), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3782) );
  AOI22_X1 U4760 ( .A1(n4219), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n4151), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3781) );
  AOI22_X1 U4761 ( .A1(INSTQUEUE_REG_10__4__SCAN_IN), .A2(n4222), .B1(n4225), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3780) );
  NAND4_X1 U4762 ( .A1(n3783), .A2(n3782), .A3(n3781), .A4(n3780), .ZN(n3784)
         );
  OAI21_X1 U4763 ( .B1(n3785), .B2(n3784), .A(n2965), .ZN(n3786) );
  NAND2_X1 U4764 ( .A1(n3787), .A2(n3786), .ZN(n5429) );
  INV_X1 U4765 ( .A(n5429), .ZN(n3833) );
  XOR2_X1 U4766 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .B(n3788), .Z(n6163) );
  AOI22_X1 U4767 ( .A1(n2962), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4078), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3792) );
  AOI22_X1 U4768 ( .A1(n3232), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4107), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3791) );
  AOI22_X1 U4769 ( .A1(n4173), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n4214), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3790) );
  AOI22_X1 U4770 ( .A1(n4174), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n4225), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3789) );
  NAND4_X1 U4771 ( .A1(n3792), .A2(n3791), .A3(n3790), .A4(n3789), .ZN(n3798)
         );
  AOI22_X1 U4772 ( .A1(n3961), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4175), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3796) );
  AOI22_X1 U4773 ( .A1(n4211), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4213), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3795) );
  AOI22_X1 U4774 ( .A1(n4222), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4151), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3794) );
  AOI22_X1 U4775 ( .A1(n4219), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n4223), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3793) );
  NAND4_X1 U4776 ( .A1(n3796), .A2(n3795), .A3(n3794), .A4(n3793), .ZN(n3797)
         );
  OR2_X1 U4777 ( .A1(n3798), .A2(n3797), .ZN(n3799) );
  AOI22_X1 U4778 ( .A1(n2965), .A2(n3799), .B1(n5335), .B2(
        PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3801) );
  NAND2_X1 U4779 ( .A1(n4237), .A2(EAX_REG_11__SCAN_IN), .ZN(n3800) );
  OAI211_X1 U4780 ( .C1(n6163), .C2(n4235), .A(n3801), .B(n3800), .ZN(n5495)
         );
  INV_X1 U4781 ( .A(n5495), .ZN(n3832) );
  XNOR2_X1 U4782 ( .A(n3802), .B(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n5298)
         );
  AOI22_X1 U4783 ( .A1(n4078), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n4214), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3806) );
  AOI22_X1 U4784 ( .A1(n3961), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4219), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3805) );
  AOI22_X1 U4785 ( .A1(n4211), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n4156), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3804) );
  AOI22_X1 U4786 ( .A1(n3232), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4225), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3803) );
  NAND4_X1 U4787 ( .A1(n3806), .A2(n3805), .A3(n3804), .A4(n3803), .ZN(n3812)
         );
  AOI22_X1 U4788 ( .A1(n4173), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n4175), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3810) );
  AOI22_X1 U4789 ( .A1(n4222), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4107), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3809) );
  AOI22_X1 U4790 ( .A1(n2962), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4213), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3808) );
  AOI22_X1 U4791 ( .A1(n4224), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n4223), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3807) );
  NAND4_X1 U4792 ( .A1(n3810), .A2(n3809), .A3(n3808), .A4(n3807), .ZN(n3811)
         );
  OAI21_X1 U4793 ( .B1(n3812), .B2(n3811), .A(n2965), .ZN(n3815) );
  NAND2_X1 U4794 ( .A1(n5336), .A2(EAX_REG_10__SCAN_IN), .ZN(n3814) );
  NAND2_X1 U4795 ( .A1(n5335), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3813)
         );
  NAND3_X1 U4796 ( .A1(n3815), .A2(n3814), .A3(n3813), .ZN(n3816) );
  AOI21_X1 U4797 ( .B1(n5298), .B2(n4241), .A(n3816), .ZN(n5056) );
  AOI22_X1 U4798 ( .A1(n4078), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n4173), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3820) );
  AOI22_X1 U4799 ( .A1(n4222), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n4107), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3819) );
  AOI22_X1 U4800 ( .A1(n3049), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4156), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3818) );
  AOI22_X1 U4801 ( .A1(n4225), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n4223), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3817) );
  NAND4_X1 U4802 ( .A1(n3820), .A2(n3819), .A3(n3818), .A4(n3817), .ZN(n3826)
         );
  AOI22_X1 U4803 ( .A1(n3961), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4219), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3824) );
  AOI22_X1 U4804 ( .A1(n3888), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4214), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3823) );
  AOI22_X1 U4805 ( .A1(n4211), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n4213), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3822) );
  AOI22_X1 U4806 ( .A1(n3232), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n4151), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3821) );
  NAND4_X1 U4807 ( .A1(n3824), .A2(n3823), .A3(n3822), .A4(n3821), .ZN(n3825)
         );
  OAI21_X1 U4808 ( .B1(n3826), .B2(n3825), .A(n2965), .ZN(n3831) );
  NAND2_X1 U4809 ( .A1(n5336), .A2(EAX_REG_8__SCAN_IN), .ZN(n3830) );
  XNOR2_X1 U4810 ( .A(n3827), .B(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n5221) );
  NAND2_X1 U4811 ( .A1(n5221), .A2(n4241), .ZN(n3829) );
  NAND2_X1 U4812 ( .A1(n5335), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3828)
         );
  NAND4_X1 U4813 ( .A1(n3831), .A2(n3830), .A3(n3829), .A4(n3828), .ZN(n4981)
         );
  INV_X1 U4814 ( .A(n4981), .ZN(n4978) );
  OR2_X1 U4815 ( .A1(n5056), .A2(n4978), .ZN(n5053) );
  OR2_X1 U4816 ( .A1(n3832), .A2(n5053), .ZN(n5425) );
  NOR2_X1 U4817 ( .A1(n3833), .A2(n5425), .ZN(n3834) );
  NAND3_X1 U4818 ( .A1(n3836), .A2(n5428), .A3(n2968), .ZN(n4662) );
  INV_X1 U4819 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n5230) );
  XOR2_X1 U4820 ( .A(n5230), .B(n3854), .Z(n5620) );
  INV_X1 U4821 ( .A(n5620), .ZN(n5235) );
  AOI22_X1 U4822 ( .A1(n4211), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n4173), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3841) );
  AOI22_X1 U4823 ( .A1(n4222), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4107), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3840) );
  AOI22_X1 U4824 ( .A1(n4214), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4213), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3839) );
  AOI22_X1 U4825 ( .A1(n4175), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4224), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3838) );
  NAND4_X1 U4826 ( .A1(n3841), .A2(n3840), .A3(n3839), .A4(n3838), .ZN(n3847)
         );
  AOI22_X1 U4827 ( .A1(n3888), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4078), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3845) );
  AOI22_X1 U4828 ( .A1(n4220), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4156), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3844) );
  AOI22_X1 U4829 ( .A1(n4219), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n4223), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3843) );
  AOI22_X1 U4830 ( .A1(n3232), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4225), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3842) );
  NAND4_X1 U4831 ( .A1(n3845), .A2(n3844), .A3(n3843), .A4(n3842), .ZN(n3846)
         );
  OAI21_X1 U4832 ( .B1(n3847), .B2(n3846), .A(n2965), .ZN(n3850) );
  NAND2_X1 U4833 ( .A1(n4237), .A2(EAX_REG_13__SCAN_IN), .ZN(n3849) );
  NAND2_X1 U4834 ( .A1(n5335), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3848)
         );
  NAND3_X1 U4835 ( .A1(n3850), .A2(n3849), .A3(n3848), .ZN(n3851) );
  AOI21_X1 U4836 ( .B1(n5235), .B2(n4196), .A(n3851), .ZN(n4664) );
  XNOR2_X1 U4837 ( .A(n3869), .B(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n5611)
         );
  AOI22_X1 U4838 ( .A1(n2962), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4078), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3858) );
  AOI22_X1 U4839 ( .A1(n4211), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n4173), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3857) );
  AOI22_X1 U4840 ( .A1(n3232), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4107), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3856) );
  AOI22_X1 U4841 ( .A1(n4175), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4151), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3855) );
  NAND4_X1 U4842 ( .A1(n3858), .A2(n3857), .A3(n3856), .A4(n3855), .ZN(n3864)
         );
  AOI22_X1 U4843 ( .A1(n3961), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4156), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3862) );
  AOI22_X1 U4844 ( .A1(n4214), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4213), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3861) );
  AOI22_X1 U4845 ( .A1(n4222), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4225), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3860) );
  AOI22_X1 U4846 ( .A1(n4219), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n4223), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3859) );
  NAND4_X1 U4847 ( .A1(n3862), .A2(n3861), .A3(n3860), .A4(n3859), .ZN(n3863)
         );
  OAI21_X1 U4848 ( .B1(n3864), .B2(n3863), .A(n2965), .ZN(n3867) );
  NAND2_X1 U4849 ( .A1(n4237), .A2(EAX_REG_14__SCAN_IN), .ZN(n3866) );
  NAND2_X1 U4850 ( .A1(n5335), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n3865)
         );
  NAND3_X1 U4851 ( .A1(n3867), .A2(n3866), .A3(n3865), .ZN(n3868) );
  AOI21_X1 U4852 ( .B1(n5611), .B2(n4196), .A(n3868), .ZN(n4924) );
  INV_X1 U4853 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n5292) );
  XOR2_X1 U4854 ( .A(n5292), .B(n3883), .Z(n5601) );
  AOI22_X1 U4855 ( .A1(n3888), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4078), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3873) );
  AOI22_X1 U4856 ( .A1(n4222), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4107), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3872) );
  AOI22_X1 U4857 ( .A1(n4175), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4156), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3871) );
  AOI22_X1 U4858 ( .A1(n3961), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4151), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3870) );
  NAND4_X1 U4859 ( .A1(n3873), .A2(n3872), .A3(n3871), .A4(n3870), .ZN(n3879)
         );
  AOI22_X1 U4860 ( .A1(n4211), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4173), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3877) );
  AOI22_X1 U4861 ( .A1(n4214), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4213), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3876) );
  AOI22_X1 U4862 ( .A1(n3232), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n4225), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3875) );
  AOI22_X1 U4863 ( .A1(n4219), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n4223), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3874) );
  NAND4_X1 U4864 ( .A1(n3877), .A2(n3876), .A3(n3875), .A4(n3874), .ZN(n3878)
         );
  OR2_X1 U4865 ( .A1(n3879), .A2(n3878), .ZN(n3880) );
  AOI22_X1 U4866 ( .A1(n2965), .A2(n3880), .B1(n5335), .B2(
        PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3882) );
  NAND2_X1 U4867 ( .A1(n4237), .A2(EAX_REG_15__SCAN_IN), .ZN(n3881) );
  OAI211_X1 U4868 ( .C1(n5601), .C2(n4235), .A(n3882), .B(n3881), .ZN(n4964)
         );
  AND2_X2 U4869 ( .A1(n4921), .A2(n4964), .ZN(n4963) );
  INV_X1 U4870 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n6723) );
  NAND2_X1 U4871 ( .A1(n3884), .A2(n6723), .ZN(n3886) );
  INV_X1 U4872 ( .A(n3918), .ZN(n3885) );
  NAND2_X1 U4873 ( .A1(n3886), .A2(n3885), .ZN(n6007) );
  NAND2_X1 U4874 ( .A1(n6007), .A2(n4196), .ZN(n3903) );
  NOR2_X1 U4875 ( .A1(n3887), .A2(n6443), .ZN(n4187) );
  AOI22_X1 U4876 ( .A1(n2962), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n3060), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3892) );
  AOI22_X1 U4877 ( .A1(n4211), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n4175), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3891) );
  AOI22_X1 U4878 ( .A1(n4173), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n4214), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3890) );
  AOI22_X1 U4879 ( .A1(n4219), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n4224), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3889) );
  NAND4_X1 U4880 ( .A1(n3892), .A2(n3891), .A3(n3890), .A4(n3889), .ZN(n3898)
         );
  AOI22_X1 U4881 ( .A1(n4222), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4107), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3896) );
  AOI22_X1 U4882 ( .A1(n4174), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n4213), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3895) );
  AOI22_X1 U4883 ( .A1(n3232), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3015), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3894) );
  AOI22_X1 U4884 ( .A1(n3961), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4223), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3893) );
  NAND4_X1 U4885 ( .A1(n3896), .A2(n3895), .A3(n3894), .A4(n3893), .ZN(n3897)
         );
  OR2_X1 U4886 ( .A1(n3898), .A2(n3897), .ZN(n3901) );
  INV_X1 U4887 ( .A(EAX_REG_16__SCAN_IN), .ZN(n3899) );
  OAI22_X1 U4888 ( .A1(n3704), .A2(n3899), .B1(n4074), .B2(n6723), .ZN(n3900)
         );
  AOI21_X1 U4889 ( .B1(n4187), .B2(n3901), .A(n3900), .ZN(n3902) );
  NAND2_X1 U4890 ( .A1(n3903), .A2(n3902), .ZN(n5068) );
  NAND2_X1 U4891 ( .A1(n4963), .A2(n5068), .ZN(n5066) );
  AOI22_X1 U4892 ( .A1(n4211), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4214), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3907) );
  AOI22_X1 U4893 ( .A1(n3232), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4131), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3906) );
  AOI22_X1 U4894 ( .A1(n4219), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n4156), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3905) );
  AOI22_X1 U4895 ( .A1(n4224), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n4223), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3904) );
  NAND4_X1 U4896 ( .A1(n3907), .A2(n3906), .A3(n3905), .A4(n3904), .ZN(n3913)
         );
  AOI22_X1 U4897 ( .A1(n3888), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4078), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3911) );
  AOI22_X1 U4898 ( .A1(n3961), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4175), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3910) );
  AOI22_X1 U4899 ( .A1(n4173), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n4176), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3909) );
  AOI22_X1 U4900 ( .A1(n4107), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n3015), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3908) );
  NAND4_X1 U4901 ( .A1(n3911), .A2(n3910), .A3(n3909), .A4(n3908), .ZN(n3912)
         );
  NOR2_X1 U4902 ( .A1(n3913), .A2(n3912), .ZN(n3917) );
  OAI21_X1 U4903 ( .B1(PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n5973), .A(n6661), 
        .ZN(n3914) );
  INV_X1 U4904 ( .A(n3914), .ZN(n3915) );
  AOI21_X1 U4905 ( .B1(n4237), .B2(EAX_REG_17__SCAN_IN), .A(n3915), .ZN(n3916)
         );
  OAI21_X1 U4906 ( .B1(n4239), .B2(n3917), .A(n3916), .ZN(n3920) );
  OAI21_X1 U4907 ( .B1(PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n3918), .A(n3950), 
        .ZN(n6703) );
  OR2_X1 U4908 ( .A1(n6703), .A2(n4235), .ZN(n3919) );
  NAND2_X1 U4909 ( .A1(n3920), .A2(n3919), .ZN(n5935) );
  OR2_X2 U4910 ( .A1(n5066), .A2(n5935), .ZN(n5937) );
  AOI22_X1 U4911 ( .A1(n2962), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4078), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3924) );
  AOI22_X1 U4912 ( .A1(n4211), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4173), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3923) );
  AOI22_X1 U4913 ( .A1(n4175), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4156), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3922) );
  AOI22_X1 U4914 ( .A1(n4214), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4176), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3921) );
  NAND4_X1 U4915 ( .A1(n3924), .A2(n3923), .A3(n3922), .A4(n3921), .ZN(n3930)
         );
  AOI22_X1 U4916 ( .A1(n3961), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4219), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3928) );
  AOI22_X1 U4917 ( .A1(n4222), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4107), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3927) );
  AOI22_X1 U4918 ( .A1(n4224), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n4223), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3926) );
  AOI22_X1 U4919 ( .A1(n3232), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3015), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3925) );
  NAND4_X1 U4920 ( .A1(n3928), .A2(n3927), .A3(n3926), .A4(n3925), .ZN(n3929)
         );
  NOR2_X1 U4921 ( .A1(n3930), .A2(n3929), .ZN(n3933) );
  INV_X1 U4922 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n5581) );
  AOI21_X1 U4923 ( .B1(n5581), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3931) );
  AOI21_X1 U4924 ( .B1(n4237), .B2(EAX_REG_18__SCAN_IN), .A(n3931), .ZN(n3932)
         );
  OAI21_X1 U4925 ( .B1(n4239), .B2(n3933), .A(n3932), .ZN(n3935) );
  XNOR2_X1 U4926 ( .A(n3950), .B(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n5998)
         );
  NAND2_X1 U4927 ( .A1(n5998), .A2(n4196), .ZN(n3934) );
  NAND2_X1 U4928 ( .A1(n3935), .A2(n3934), .ZN(n5247) );
  AOI22_X1 U4929 ( .A1(n3888), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4078), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3939) );
  AOI22_X1 U4930 ( .A1(n3961), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4211), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3938) );
  AOI22_X1 U4931 ( .A1(n4173), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n4214), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3937) );
  AOI22_X1 U4932 ( .A1(n4224), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n3015), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3936) );
  NAND4_X1 U4933 ( .A1(n3939), .A2(n3938), .A3(n3937), .A4(n3936), .ZN(n3945)
         );
  AOI22_X1 U4934 ( .A1(n4222), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4107), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3943) );
  AOI22_X1 U4935 ( .A1(n4219), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n4156), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3942) );
  AOI22_X1 U4936 ( .A1(n4175), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4213), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3941) );
  AOI22_X1 U4937 ( .A1(n3232), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4223), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3940) );
  NAND4_X1 U4938 ( .A1(n3943), .A2(n3942), .A3(n3941), .A4(n3940), .ZN(n3944)
         );
  NOR2_X1 U4939 ( .A1(n3945), .A2(n3944), .ZN(n3949) );
  OAI21_X1 U4940 ( .B1(PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n5973), .A(n6661), 
        .ZN(n3946) );
  INV_X1 U4941 ( .A(n3946), .ZN(n3947) );
  AOI21_X1 U4942 ( .B1(n4237), .B2(EAX_REG_19__SCAN_IN), .A(n3947), .ZN(n3948)
         );
  OAI21_X1 U4943 ( .B1(n4239), .B2(n3949), .A(n3948), .ZN(n3955) );
  NOR2_X1 U4944 ( .A1(n3951), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n3952)
         );
  OR2_X1 U4945 ( .A1(n3986), .A2(n3952), .ZN(n5900) );
  INV_X1 U4946 ( .A(n5900), .ZN(n3953) );
  NAND2_X1 U4947 ( .A1(n3953), .A2(n4241), .ZN(n3954) );
  NAND2_X1 U4948 ( .A1(n3955), .A2(n3954), .ZN(n5303) );
  AND2_X2 U4949 ( .A1(n5246), .A2(n3956), .ZN(n5314) );
  AOI22_X1 U4950 ( .A1(n2962), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n4078), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3960) );
  AOI22_X1 U4951 ( .A1(n4211), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n4173), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3959) );
  AOI22_X1 U4952 ( .A1(INSTQUEUE_REG_14__4__SCAN_IN), .A2(n4175), .B1(n4174), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3958) );
  AOI22_X1 U4953 ( .A1(INSTQUEUE_REG_10__4__SCAN_IN), .A2(n4214), .B1(n4176), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3957) );
  NAND4_X1 U4954 ( .A1(n3960), .A2(n3959), .A3(n3958), .A4(n3957), .ZN(n3967)
         );
  AOI22_X1 U4955 ( .A1(n3961), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4219), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3965) );
  AOI22_X1 U4956 ( .A1(INSTQUEUE_REG_4__4__SCAN_IN), .A2(n4107), .B1(n4131), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3964) );
  AOI22_X1 U4957 ( .A1(n4224), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n3190), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3963) );
  AOI22_X1 U4958 ( .A1(n3224), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n4225), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3962) );
  NAND4_X1 U4959 ( .A1(n3965), .A2(n3964), .A3(n3963), .A4(n3962), .ZN(n3966)
         );
  NOR2_X1 U4960 ( .A1(n3967), .A2(n3966), .ZN(n3970) );
  INV_X1 U4961 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n5898) );
  AOI21_X1 U4962 ( .B1(n5898), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3968) );
  AOI21_X1 U4963 ( .B1(n4237), .B2(EAX_REG_20__SCAN_IN), .A(n3968), .ZN(n3969)
         );
  OAI21_X1 U4964 ( .B1(n4239), .B2(n3970), .A(n3969), .ZN(n3972) );
  XNOR2_X1 U4965 ( .A(n3986), .B(n5898), .ZN(n5890) );
  NAND2_X1 U4966 ( .A1(n5890), .A2(n4241), .ZN(n3971) );
  AND2_X1 U4967 ( .A1(n3972), .A2(n3971), .ZN(n5313) );
  AOI22_X1 U4968 ( .A1(n3961), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4173), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3976) );
  AOI22_X1 U4969 ( .A1(n3224), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4131), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3975) );
  AOI22_X1 U4970 ( .A1(n3888), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4176), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3974) );
  AOI22_X1 U4971 ( .A1(n4219), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n3190), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3973) );
  NAND4_X1 U4972 ( .A1(n3976), .A2(n3975), .A3(n3974), .A4(n3973), .ZN(n3982)
         );
  AOI22_X1 U4973 ( .A1(n4211), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4175), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3980) );
  AOI22_X1 U4974 ( .A1(n4078), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n4214), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3979) );
  AOI22_X1 U4975 ( .A1(n4174), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n4224), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3978) );
  AOI22_X1 U4976 ( .A1(n4107), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n4225), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3977) );
  NAND4_X1 U4977 ( .A1(n3980), .A2(n3979), .A3(n3978), .A4(n3977), .ZN(n3981)
         );
  NOR2_X1 U4978 ( .A1(n3982), .A2(n3981), .ZN(n3985) );
  INV_X1 U4979 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n3987) );
  OAI21_X1 U4980 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n3987), .A(n4235), .ZN(
        n3983) );
  AOI21_X1 U4981 ( .B1(n4237), .B2(EAX_REG_21__SCAN_IN), .A(n3983), .ZN(n3984)
         );
  OAI21_X1 U4982 ( .B1(n4239), .B2(n3985), .A(n3984), .ZN(n3991) );
  NAND2_X1 U4983 ( .A1(n3988), .A2(n3987), .ZN(n3989) );
  NAND2_X1 U4984 ( .A1(n4056), .A2(n3989), .ZN(n5881) );
  OR2_X1 U4985 ( .A1(n5881), .A2(n4235), .ZN(n3990) );
  NAND2_X1 U4986 ( .A1(n3991), .A2(n3990), .ZN(n5466) );
  NOR2_X2 U4987 ( .A1(n5465), .A2(n5466), .ZN(n4010) );
  INV_X1 U4988 ( .A(n3992), .ZN(n5464) );
  AOI22_X1 U4989 ( .A1(n2962), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4078), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3996) );
  AOI22_X1 U4990 ( .A1(n4211), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4173), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3995) );
  AOI22_X1 U4991 ( .A1(n4175), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4174), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3994) );
  AOI22_X1 U4992 ( .A1(n4214), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4176), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3993) );
  NAND4_X1 U4993 ( .A1(n3996), .A2(n3995), .A3(n3994), .A4(n3993), .ZN(n4002)
         );
  AOI22_X1 U4994 ( .A1(n3961), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4219), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4000) );
  AOI22_X1 U4995 ( .A1(n4222), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4221), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3999) );
  AOI22_X1 U4996 ( .A1(n4224), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n3190), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3998) );
  AOI22_X1 U4997 ( .A1(n3224), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4225), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3997) );
  NAND4_X1 U4998 ( .A1(n4000), .A2(n3999), .A3(n3998), .A4(n3997), .ZN(n4001)
         );
  NOR2_X1 U4999 ( .A1(n4002), .A2(n4001), .ZN(n4005) );
  INV_X1 U5000 ( .A(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n4055) );
  AOI21_X1 U5001 ( .B1(n4055), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4003) );
  AOI21_X1 U5002 ( .B1(n4237), .B2(EAX_REG_22__SCAN_IN), .A(n4003), .ZN(n4004)
         );
  OAI21_X1 U5003 ( .B1(n4239), .B2(n4005), .A(n4004), .ZN(n4007) );
  XNOR2_X1 U5004 ( .A(n4056), .B(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5873)
         );
  NAND2_X1 U5005 ( .A1(n5873), .A2(n4241), .ZN(n4006) );
  NAND2_X1 U5006 ( .A1(n4007), .A2(n4006), .ZN(n4008) );
  AND2_X1 U5007 ( .A1(n5464), .A2(n4008), .ZN(n4011) );
  AND2_X2 U5008 ( .A1(n4010), .A2(n4009), .ZN(n4061) );
  OR2_X1 U5009 ( .A1(n4011), .A2(n4061), .ZN(n5874) );
  NAND3_X1 U5010 ( .A1(n6443), .A2(STATEBS16_REG_SCAN_IN), .A3(
        STATE2_REG_1__SCAN_IN), .ZN(n6452) );
  INV_X1 U5011 ( .A(n6452), .ZN(n4012) );
  NOR2_X1 U5012 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATE2_REG_3__SCAN_IN), .ZN(
        n5089) );
  AND2_X1 U5013 ( .A1(n4012), .A2(n5089), .ZN(n5593) );
  INV_X1 U5014 ( .A(n5593), .ZN(n5634) );
  INV_X1 U5015 ( .A(n5089), .ZN(n5791) );
  NAND2_X1 U5016 ( .A1(n5791), .A2(n4013), .ZN(n4014) );
  NAND2_X1 U5017 ( .A1(n4014), .A2(n6443), .ZN(n4015) );
  NAND2_X1 U5018 ( .A1(n6443), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4017) );
  NAND2_X1 U5019 ( .A1(n5973), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4016) );
  AND2_X1 U5020 ( .A1(n4017), .A2(n4016), .ZN(n4423) );
  INV_X1 U5021 ( .A(REIP_REG_22__SCAN_IN), .ZN(n4018) );
  NOR2_X1 U5022 ( .A1(n6248), .A2(n4018), .ZN(n5692) );
  NOR2_X1 U5023 ( .A1(n5618), .A2(n4055), .ZN(n4019) );
  AOI211_X1 U5024 ( .C1(n6164), .C2(n5873), .A(n5692), .B(n4019), .ZN(n4020)
         );
  NAND2_X1 U5025 ( .A1(n4023), .A2(n4022), .ZN(U2964) );
  INV_X1 U5026 ( .A(n5345), .ZN(n4026) );
  NAND2_X1 U5027 ( .A1(n5518), .A2(n5637), .ZN(n4024) );
  OR2_X1 U5028 ( .A1(n5520), .A2(n4024), .ZN(n4025) );
  AOI22_X1 U5029 ( .A1(n3888), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n4078), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4031) );
  AOI22_X1 U5030 ( .A1(n4211), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n4173), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n4030) );
  INV_X1 U5031 ( .A(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n6710) );
  AOI22_X1 U5032 ( .A1(n4175), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n4156), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n4029) );
  AOI22_X1 U5033 ( .A1(n4214), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4213), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n4028) );
  NAND4_X1 U5034 ( .A1(n4031), .A2(n4030), .A3(n4029), .A4(n4028), .ZN(n4037)
         );
  AOI22_X1 U5035 ( .A1(n4112), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4219), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n4035) );
  AOI22_X1 U5036 ( .A1(n4150), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4107), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n4034) );
  AOI22_X1 U5037 ( .A1(n4224), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n4223), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4033) );
  AOI22_X1 U5038 ( .A1(n3232), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3015), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4032) );
  NAND4_X1 U5039 ( .A1(n4035), .A2(n4034), .A3(n4033), .A4(n4032), .ZN(n4036)
         );
  OR2_X1 U5040 ( .A1(n4037), .A2(n4036), .ZN(n4050) );
  AOI22_X1 U5041 ( .A1(n2962), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4078), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4041) );
  AOI22_X1 U5042 ( .A1(n4211), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n4173), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4040) );
  AOI22_X1 U5043 ( .A1(n4175), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n4156), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4039) );
  AOI22_X1 U5044 ( .A1(n4214), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4213), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4038) );
  NAND4_X1 U5045 ( .A1(n4041), .A2(n4040), .A3(n4039), .A4(n4038), .ZN(n4047)
         );
  AOI22_X1 U5046 ( .A1(n4112), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4219), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4045) );
  AOI22_X1 U5047 ( .A1(n4150), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4107), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4044) );
  AOI22_X1 U5048 ( .A1(n4224), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n4223), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4043) );
  AOI22_X1 U5049 ( .A1(n3232), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3015), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4042) );
  NAND4_X1 U5050 ( .A1(n4045), .A2(n4044), .A3(n4043), .A4(n4042), .ZN(n4046)
         );
  OR2_X1 U5051 ( .A1(n4047), .A2(n4046), .ZN(n4049) );
  AND2_X1 U5052 ( .A1(n4049), .A2(n4050), .ZN(n4089) );
  INV_X1 U5053 ( .A(n4089), .ZN(n4048) );
  OAI21_X1 U5054 ( .B1(n4050), .B2(n4049), .A(n4048), .ZN(n4054) );
  NAND2_X1 U5055 ( .A1(n6661), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n4051)
         );
  NAND2_X1 U5056 ( .A1(n4235), .A2(n4051), .ZN(n4052) );
  AOI21_X1 U5057 ( .B1(n4237), .B2(EAX_REG_23__SCAN_IN), .A(n4052), .ZN(n4053)
         );
  OAI21_X1 U5058 ( .B1(n4239), .B2(n4054), .A(n4053), .ZN(n4060) );
  OR2_X1 U5059 ( .A1(n4057), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n4058)
         );
  NAND2_X1 U5060 ( .A1(n4095), .A2(n4058), .ZN(n5864) );
  OR2_X1 U5061 ( .A1(n5864), .A2(n4235), .ZN(n4059) );
  XNOR2_X1 U5062 ( .A(n4095), .B(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5853)
         );
  AOI22_X1 U5063 ( .A1(n2962), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n4078), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4065) );
  AOI22_X1 U5064 ( .A1(n4211), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4173), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n4064) );
  AOI22_X1 U5065 ( .A1(n4175), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n4174), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n4063) );
  AOI22_X1 U5066 ( .A1(n4214), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4176), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n4062) );
  NAND4_X1 U5067 ( .A1(n4065), .A2(n4064), .A3(n4063), .A4(n4062), .ZN(n4071)
         );
  AOI22_X1 U5068 ( .A1(n4112), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4219), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n4069) );
  AOI22_X1 U5069 ( .A1(n4150), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4107), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n4068) );
  AOI22_X1 U5070 ( .A1(n4224), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n4223), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4067) );
  AOI22_X1 U5071 ( .A1(n3232), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3015), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4066) );
  NAND4_X1 U5072 ( .A1(n4069), .A2(n4068), .A3(n4067), .A4(n4066), .ZN(n4070)
         );
  OR2_X1 U5073 ( .A1(n4071), .A2(n4070), .ZN(n4090) );
  INV_X1 U5074 ( .A(n4090), .ZN(n4072) );
  XNOR2_X1 U5075 ( .A(n4089), .B(n4072), .ZN(n4073) );
  NAND2_X1 U5076 ( .A1(n4187), .A2(n4073), .ZN(n4077) );
  INV_X1 U5077 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5541) );
  NOR2_X1 U5078 ( .A1(n4074), .A2(n5541), .ZN(n4075) );
  AOI21_X1 U5079 ( .B1(n4237), .B2(EAX_REG_24__SCAN_IN), .A(n4075), .ZN(n4076)
         );
  OAI211_X1 U5080 ( .C1(n5853), .C2(n4235), .A(n4077), .B(n4076), .ZN(n5454)
         );
  AOI22_X1 U5081 ( .A1(n4078), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n4211), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n4082) );
  AOI22_X1 U5082 ( .A1(n3888), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4131), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n4081) );
  AOI22_X1 U5083 ( .A1(n3232), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4225), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4080) );
  AOI22_X1 U5084 ( .A1(n4221), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n4213), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n4079) );
  NAND4_X1 U5085 ( .A1(n4082), .A2(n4081), .A3(n4080), .A4(n4079), .ZN(n4088)
         );
  AOI22_X1 U5086 ( .A1(n4112), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4173), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n4086) );
  AOI22_X1 U5087 ( .A1(n3049), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n4156), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n4085) );
  AOI22_X1 U5088 ( .A1(n4214), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4223), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4084) );
  AOI22_X1 U5089 ( .A1(n4219), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n4151), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4083) );
  NAND4_X1 U5090 ( .A1(n4086), .A2(n4085), .A3(n4084), .A4(n4083), .ZN(n4087)
         );
  OR2_X1 U5091 ( .A1(n4088), .A2(n4087), .ZN(n4104) );
  NAND2_X1 U5092 ( .A1(n4090), .A2(n4089), .ZN(n4106) );
  INV_X1 U5093 ( .A(n4106), .ZN(n4091) );
  XNOR2_X1 U5094 ( .A(n4104), .B(n4091), .ZN(n4094) );
  INV_X1 U5095 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n4096) );
  OAI21_X1 U5096 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n4096), .A(n4235), .ZN(
        n4092) );
  AOI21_X1 U5097 ( .B1(n4237), .B2(EAX_REG_25__SCAN_IN), .A(n4092), .ZN(n4093)
         );
  OAI21_X1 U5098 ( .B1(n4239), .B2(n4094), .A(n4093), .ZN(n4101) );
  NAND2_X1 U5099 ( .A1(n4097), .A2(n4096), .ZN(n4098) );
  NAND2_X1 U5100 ( .A1(n4142), .A2(n4098), .ZN(n5533) );
  INV_X1 U5101 ( .A(n5533), .ZN(n4099) );
  NAND2_X1 U5102 ( .A1(n4099), .A2(n4196), .ZN(n4100) );
  NAND2_X1 U5103 ( .A1(n4101), .A2(n4100), .ZN(n5413) );
  INV_X1 U5104 ( .A(n4104), .ZN(n4105) );
  OR2_X1 U5105 ( .A1(n4106), .A2(n4105), .ZN(n4125) );
  AOI22_X1 U5106 ( .A1(n3888), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4078), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4111) );
  AOI22_X1 U5107 ( .A1(n4175), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n4219), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n4110) );
  AOI22_X1 U5108 ( .A1(n4173), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n4214), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n4109) );
  AOI22_X1 U5109 ( .A1(n4107), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3190), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4108) );
  NAND4_X1 U5110 ( .A1(n4111), .A2(n4110), .A3(n4109), .A4(n4108), .ZN(n4118)
         );
  AOI22_X1 U5111 ( .A1(n3224), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4131), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n4116) );
  AOI22_X1 U5112 ( .A1(n4112), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4156), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n4115) );
  AOI22_X1 U5113 ( .A1(n4211), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4213), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n4114) );
  AOI22_X1 U5114 ( .A1(n4224), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n4225), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4113) );
  NAND4_X1 U5115 ( .A1(n4116), .A2(n4115), .A3(n4114), .A4(n4113), .ZN(n4117)
         );
  NOR2_X1 U5116 ( .A1(n4118), .A2(n4117), .ZN(n4126) );
  XOR2_X1 U5117 ( .A(n4125), .B(n4126), .Z(n4119) );
  NAND2_X1 U5118 ( .A1(n4119), .A2(n4187), .ZN(n4122) );
  INV_X1 U5119 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n5524) );
  OAI21_X1 U5120 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n5524), .A(n4235), .ZN(
        n4120) );
  AOI21_X1 U5121 ( .B1(n4237), .B2(EAX_REG_26__SCAN_IN), .A(n4120), .ZN(n4121)
         );
  NAND2_X1 U5122 ( .A1(n4122), .A2(n4121), .ZN(n4124) );
  XNOR2_X1 U5123 ( .A(n4142), .B(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n5522)
         );
  NAND2_X1 U5124 ( .A1(n5522), .A2(n4196), .ZN(n4123) );
  NAND2_X1 U5125 ( .A1(n4124), .A2(n4123), .ZN(n5402) );
  NOR2_X1 U5126 ( .A1(n4126), .A2(n4125), .ZN(n4165) );
  AOI22_X1 U5127 ( .A1(INSTQUEUE_REG_14__4__SCAN_IN), .A2(n3888), .B1(n3060), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4130) );
  AOI22_X1 U5128 ( .A1(n4211), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n4173), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n4129) );
  AOI22_X1 U5129 ( .A1(n4175), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n4156), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n4128) );
  AOI22_X1 U5130 ( .A1(n4214), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4157), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4127) );
  NAND4_X1 U5131 ( .A1(n4130), .A2(n4129), .A3(n4128), .A4(n4127), .ZN(n4137)
         );
  AOI22_X1 U5132 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n3961), .B1(n4219), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n4135) );
  AOI22_X1 U5133 ( .A1(INSTQUEUE_REG_5__4__SCAN_IN), .A2(n4221), .B1(n4131), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n4134) );
  AOI22_X1 U5134 ( .A1(n4224), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n3190), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4133) );
  AOI22_X1 U5135 ( .A1(n3224), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4225), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4132) );
  NAND4_X1 U5136 ( .A1(n4135), .A2(n4134), .A3(n4133), .A4(n4132), .ZN(n4136)
         );
  OR2_X1 U5137 ( .A1(n4137), .A2(n4136), .ZN(n4164) );
  INV_X1 U5138 ( .A(n4164), .ZN(n4138) );
  XNOR2_X1 U5139 ( .A(n4165), .B(n4138), .ZN(n4139) );
  NAND2_X1 U5140 ( .A1(n4139), .A2(n4187), .ZN(n4149) );
  NAND2_X1 U5141 ( .A1(n6661), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n4140)
         );
  NAND2_X1 U5142 ( .A1(n4235), .A2(n4140), .ZN(n4141) );
  AOI21_X1 U5143 ( .B1(n4237), .B2(EAX_REG_27__SCAN_IN), .A(n4141), .ZN(n4148)
         );
  INV_X1 U5144 ( .A(n4143), .ZN(n4145) );
  INV_X1 U5145 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n4144) );
  NAND2_X1 U5146 ( .A1(n4145), .A2(n4144), .ZN(n4146) );
  NAND2_X1 U5147 ( .A1(n4191), .A2(n4146), .ZN(n5845) );
  NOR2_X1 U5148 ( .A1(n5845), .A2(n4235), .ZN(n4147) );
  AOI21_X1 U5149 ( .B1(n4149), .B2(n4148), .A(n4147), .ZN(n5442) );
  INV_X1 U5150 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5394) );
  XNOR2_X1 U5151 ( .A(n4191), .B(n5394), .ZN(n5508) );
  INV_X1 U5152 ( .A(EAX_REG_28__SCAN_IN), .ZN(n4169) );
  AOI22_X1 U5153 ( .A1(n2962), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n4078), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4155) );
  AOI22_X1 U5154 ( .A1(n4220), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4219), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n4154) );
  AOI22_X1 U5155 ( .A1(n4150), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4221), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4153) );
  AOI22_X1 U5156 ( .A1(n3224), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4151), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4152) );
  NAND4_X1 U5157 ( .A1(n4155), .A2(n4154), .A3(n4153), .A4(n4152), .ZN(n4163)
         );
  AOI22_X1 U5158 ( .A1(n4211), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4173), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4161) );
  AOI22_X1 U5159 ( .A1(n4175), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n4156), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n4160) );
  AOI22_X1 U5160 ( .A1(n4214), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4157), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4159) );
  AOI22_X1 U5161 ( .A1(n4225), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n3190), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4158) );
  NAND4_X1 U5162 ( .A1(n4161), .A2(n4160), .A3(n4159), .A4(n4158), .ZN(n4162)
         );
  NOR2_X1 U5163 ( .A1(n4163), .A2(n4162), .ZN(n4172) );
  NAND2_X1 U5164 ( .A1(n4165), .A2(n4164), .ZN(n4171) );
  XOR2_X1 U5165 ( .A(n4172), .B(n4171), .Z(n4166) );
  NAND2_X1 U5166 ( .A1(n4166), .A2(n4187), .ZN(n4168) );
  AOI21_X1 U5167 ( .B1(PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n6661), .A(n4241), 
        .ZN(n4167) );
  OAI211_X1 U5168 ( .C1(n3704), .C2(n4169), .A(n4168), .B(n4167), .ZN(n4170)
         );
  OAI21_X1 U5169 ( .B1(n4235), .B2(n5508), .A(n4170), .ZN(n5391) );
  NOR2_X1 U5170 ( .A1(n4172), .A2(n4171), .ZN(n4189) );
  AOI22_X1 U5171 ( .A1(n3888), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4078), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4180) );
  AOI22_X1 U5172 ( .A1(n4211), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4173), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n4179) );
  AOI22_X1 U5173 ( .A1(n4175), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n4174), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n4178) );
  AOI22_X1 U5174 ( .A1(n4214), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4176), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4177) );
  NAND4_X1 U5175 ( .A1(n4180), .A2(n4179), .A3(n4178), .A4(n4177), .ZN(n4186)
         );
  AOI22_X1 U5176 ( .A1(n3961), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4219), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4184) );
  AOI22_X1 U5177 ( .A1(n4222), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4221), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4183) );
  AOI22_X1 U5178 ( .A1(n4224), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3190), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4182) );
  AOI22_X1 U5179 ( .A1(n3224), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4225), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4181) );
  NAND4_X1 U5180 ( .A1(n4184), .A2(n4183), .A3(n4182), .A4(n4181), .ZN(n4185)
         );
  OR2_X1 U5181 ( .A1(n4186), .A2(n4185), .ZN(n4188) );
  NAND2_X1 U5182 ( .A1(n4189), .A2(n4188), .ZN(n4233) );
  OAI211_X1 U5183 ( .C1(n4189), .C2(n4188), .A(n4233), .B(n4187), .ZN(n4198)
         );
  INV_X1 U5184 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4202) );
  NOR2_X1 U5185 ( .A1(n4202), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4190) );
  AOI211_X1 U5186 ( .C1(n4237), .C2(EAX_REG_29__SCAN_IN), .A(n4190), .B(n4196), 
        .ZN(n4197) );
  INV_X1 U5187 ( .A(n4191), .ZN(n4192) );
  INV_X1 U5188 ( .A(n4193), .ZN(n4194) );
  NAND2_X1 U5189 ( .A1(n4194), .A2(n4202), .ZN(n4195) );
  AND2_X1 U5190 ( .A1(n4247), .A2(n4195), .ZN(n5370) );
  AOI22_X1 U5191 ( .A1(n4198), .A2(n4197), .B1(n5370), .B2(n4196), .ZN(n4200)
         );
  NOR2_X1 U5192 ( .A1(n5367), .A2(n5634), .ZN(n4207) );
  NAND2_X1 U5193 ( .A1(n5370), .A2(n6164), .ZN(n4205) );
  NAND2_X1 U5194 ( .A1(n3668), .A2(REIP_REG_29__SCAN_IN), .ZN(n5327) );
  OAI21_X1 U5195 ( .B1(n5618), .B2(n4202), .A(n5327), .ZN(n4203) );
  INV_X1 U5196 ( .A(n4203), .ZN(n4204) );
  OAI21_X1 U5197 ( .B1(n5332), .B2(n6169), .A(n4208), .ZN(U2957) );
  AOI22_X1 U5198 ( .A1(n2962), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3060), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4218) );
  AOI22_X1 U5199 ( .A1(n4211), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4210), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4217) );
  AOI22_X1 U5200 ( .A1(n3049), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n4156), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n4216) );
  AOI22_X1 U5201 ( .A1(n4214), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4213), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4215) );
  NAND4_X1 U5202 ( .A1(n4218), .A2(n4217), .A3(n4216), .A4(n4215), .ZN(n4231)
         );
  AOI22_X1 U5203 ( .A1(n4220), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4219), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4229) );
  AOI22_X1 U5204 ( .A1(n4222), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4221), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4228) );
  AOI22_X1 U5205 ( .A1(n4224), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n4223), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4227) );
  AOI22_X1 U5206 ( .A1(n3224), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4225), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4226) );
  NAND4_X1 U5207 ( .A1(n4229), .A2(n4228), .A3(n4227), .A4(n4226), .ZN(n4230)
         );
  NOR2_X1 U5208 ( .A1(n4231), .A2(n4230), .ZN(n4232) );
  XNOR2_X1 U5209 ( .A(n4233), .B(n4232), .ZN(n4240) );
  NAND2_X1 U5210 ( .A1(n6661), .A2(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n4234)
         );
  NAND2_X1 U5211 ( .A1(n4235), .A2(n4234), .ZN(n4236) );
  AOI21_X1 U5212 ( .B1(n4237), .B2(EAX_REG_30__SCAN_IN), .A(n4236), .ZN(n4238)
         );
  OAI21_X1 U5213 ( .B1(n4240), .B2(n4239), .A(n4238), .ZN(n4243) );
  XNOR2_X1 U5214 ( .A(n4247), .B(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5359)
         );
  NAND2_X1 U5215 ( .A1(n5359), .A2(n4241), .ZN(n4242) );
  NAND2_X1 U5216 ( .A1(n4243), .A2(n4242), .ZN(n5333) );
  AND2_X1 U5217 ( .A1(n4299), .A2(n4297), .ZN(n4291) );
  NAND2_X1 U5218 ( .A1(n4291), .A2(n6440), .ZN(n4289) );
  NOR2_X1 U5219 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATE2_REG_1__SCAN_IN), .ZN(
        n6560) );
  INV_X1 U5220 ( .A(n6560), .ZN(n6451) );
  NOR3_X1 U5221 ( .A1(n6443), .A2(n6717), .A3(n6451), .ZN(n6438) );
  AND3_X1 U5222 ( .A1(n5973), .A2(n6454), .A3(STATE2_REG_1__SCAN_IN), .ZN(
        n6450) );
  INV_X1 U5223 ( .A(n6450), .ZN(n4244) );
  NAND2_X1 U5224 ( .A1(n6248), .A2(n4244), .ZN(n4245) );
  OR2_X1 U5225 ( .A1(n6438), .A2(n4245), .ZN(n4246) );
  INV_X1 U5226 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5362) );
  INV_X1 U5227 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4248) );
  NOR2_X1 U5228 ( .A1(n5341), .A2(n6536), .ZN(n4250) );
  INV_X1 U5229 ( .A(n4252), .ZN(n4251) );
  AOI21_X1 U5230 ( .B1(n4255), .B2(n5392), .A(n4251), .ZN(n4257) );
  INV_X1 U5231 ( .A(n5392), .ZN(n4253) );
  AOI21_X1 U5232 ( .B1(n4253), .B2(n5261), .A(n4252), .ZN(n4254) );
  AOI22_X1 U5233 ( .A1(n4257), .A2(n4256), .B1(n4255), .B2(n4254), .ZN(n5354)
         );
  NOR2_X1 U5234 ( .A1(READY_N), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4267) );
  INV_X1 U5235 ( .A(EBX_REG_31__SCAN_IN), .ZN(n5325) );
  OR2_X1 U5236 ( .A1(n4267), .A2(n5325), .ZN(n4258) );
  NOR2_X1 U5237 ( .A1(n2964), .A2(n4258), .ZN(n4259) );
  AND2_X2 U5238 ( .A1(n6074), .A2(n4260), .ZN(n6077) );
  AOI22_X1 U5239 ( .A1(PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n6078), .B1(n6077), 
        .B2(n5359), .ZN(n4266) );
  OR3_X1 U5240 ( .A1(READY_N), .A2(STATEBS16_REG_SCAN_IN), .A3(n6461), .ZN(
        n6426) );
  AND2_X1 U5241 ( .A1(n4294), .A2(n6426), .ZN(n4261) );
  AND2_X1 U5242 ( .A1(n5207), .A2(n4261), .ZN(n5378) );
  INV_X1 U5243 ( .A(n5378), .ZN(n4264) );
  NOR2_X1 U5244 ( .A1(n4267), .A2(EBX_REG_31__SCAN_IN), .ZN(n4262) );
  NAND3_X1 U5245 ( .A1(n5207), .A2(n4262), .A3(n4467), .ZN(n4263) );
  NAND2_X1 U5246 ( .A1(n6695), .A2(EBX_REG_30__SCAN_IN), .ZN(n4265) );
  OAI211_X1 U5247 ( .C1(n5324), .C2(n6085), .A(n4266), .B(n4265), .ZN(n4287)
         );
  NAND3_X1 U5248 ( .A1(REIP_REG_23__SCAN_IN), .A2(REIP_REG_22__SCAN_IN), .A3(
        REIP_REG_21__SCAN_IN), .ZN(n4278) );
  INV_X1 U5249 ( .A(REIP_REG_19__SCAN_IN), .ZN(n6501) );
  INV_X1 U5250 ( .A(REIP_REG_18__SCAN_IN), .ZN(n6499) );
  NOR2_X1 U5251 ( .A1(n6501), .A2(n6499), .ZN(n4275) );
  INV_X1 U5252 ( .A(n4275), .ZN(n4270) );
  INV_X1 U5253 ( .A(REIP_REG_16__SCAN_IN), .ZN(n6496) );
  AND3_X1 U5254 ( .A1(n4268), .A2(n4267), .A3(n4467), .ZN(n4269) );
  NAND3_X1 U5255 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_3__SCAN_IN), .A3(
        REIP_REG_2__SCAN_IN), .ZN(n6042) );
  INV_X1 U5256 ( .A(REIP_REG_4__SCAN_IN), .ZN(n6477) );
  INV_X1 U5257 ( .A(REIP_REG_5__SCAN_IN), .ZN(n6724) );
  NOR3_X1 U5258 ( .A1(n6042), .A2(n6477), .A3(n6724), .ZN(n5078) );
  NAND4_X1 U5259 ( .A1(n5078), .A2(REIP_REG_7__SCAN_IN), .A3(
        REIP_REG_6__SCAN_IN), .A4(REIP_REG_8__SCAN_IN), .ZN(n5219) );
  INV_X1 U5260 ( .A(REIP_REG_9__SCAN_IN), .ZN(n6484) );
  NOR2_X1 U5261 ( .A1(n5219), .A2(n6484), .ZN(n5273) );
  NAND2_X1 U5262 ( .A1(n5273), .A2(REIP_REG_10__SCAN_IN), .ZN(n6017) );
  INV_X1 U5263 ( .A(REIP_REG_11__SCAN_IN), .ZN(n6488) );
  NOR2_X1 U5264 ( .A1(n6017), .A2(n6488), .ZN(n5231) );
  NAND2_X1 U5265 ( .A1(n5231), .A2(REIP_REG_12__SCAN_IN), .ZN(n5232) );
  INV_X1 U5266 ( .A(REIP_REG_13__SCAN_IN), .ZN(n6492) );
  NOR2_X1 U5267 ( .A1(n5232), .A2(n6492), .ZN(n5284) );
  NAND2_X1 U5268 ( .A1(n5284), .A2(REIP_REG_14__SCAN_IN), .ZN(n4271) );
  NAND2_X1 U5269 ( .A1(REIP_REG_15__SCAN_IN), .A2(n6002), .ZN(n6005) );
  NOR2_X1 U5270 ( .A1(n6496), .A2(n6005), .ZN(n6689) );
  NAND2_X1 U5271 ( .A1(REIP_REG_17__SCAN_IN), .A2(n6689), .ZN(n5906) );
  NOR2_X1 U5272 ( .A1(n4270), .A2(n5906), .ZN(n5894) );
  NAND2_X1 U5273 ( .A1(REIP_REG_20__SCAN_IN), .A2(n5894), .ZN(n5876) );
  NOR2_X1 U5274 ( .A1(n4278), .A2(n5876), .ZN(n5418) );
  NAND4_X1 U5275 ( .A1(n5418), .A2(REIP_REG_24__SCAN_IN), .A3(
        REIP_REG_26__SCAN_IN), .A4(REIP_REG_25__SCAN_IN), .ZN(n5852) );
  NAND2_X1 U5276 ( .A1(REIP_REG_28__SCAN_IN), .A2(REIP_REG_27__SCAN_IN), .ZN(
        n4282) );
  NOR2_X1 U5277 ( .A1(n5852), .A2(n4282), .ZN(n5380) );
  INV_X1 U5278 ( .A(REIP_REG_29__SCAN_IN), .ZN(n6520) );
  NAND2_X1 U5279 ( .A1(n5380), .A2(n6520), .ZN(n5375) );
  INV_X1 U5280 ( .A(n6018), .ZN(n6069) );
  INV_X1 U5281 ( .A(REIP_REG_24__SCAN_IN), .ZN(n6506) );
  INV_X1 U5282 ( .A(REIP_REG_26__SCAN_IN), .ZN(n6511) );
  INV_X1 U5283 ( .A(REIP_REG_25__SCAN_IN), .ZN(n6508) );
  NOR3_X1 U5284 ( .A1(n6506), .A2(n6511), .A3(n6508), .ZN(n4281) );
  AND2_X1 U5285 ( .A1(n6018), .A2(n6074), .ZN(n5253) );
  INV_X1 U5286 ( .A(n4271), .ZN(n4272) );
  OAI21_X1 U5287 ( .B1(n6018), .B2(n4272), .A(n6074), .ZN(n6001) );
  AND3_X1 U5288 ( .A1(REIP_REG_17__SCAN_IN), .A2(REIP_REG_15__SCAN_IN), .A3(
        REIP_REG_16__SCAN_IN), .ZN(n4273) );
  NOR2_X1 U5289 ( .A1(n6018), .A2(n4273), .ZN(n4274) );
  OR2_X1 U5290 ( .A1(n6001), .A2(n4274), .ZN(n6688) );
  AND2_X1 U5291 ( .A1(n4275), .A2(REIP_REG_20__SCAN_IN), .ZN(n4276) );
  NOR2_X1 U5292 ( .A1(n5253), .A2(n4276), .ZN(n4277) );
  INV_X1 U5293 ( .A(n4278), .ZN(n4279) );
  NOR2_X1 U5294 ( .A1(n6018), .A2(n4279), .ZN(n4280) );
  NOR2_X1 U5295 ( .A1(n5895), .A2(n4280), .ZN(n5871) );
  OAI21_X1 U5296 ( .B1(n4281), .B2(n5253), .A(n5871), .ZN(n5847) );
  AOI21_X1 U5297 ( .B1(n4282), .B2(n6069), .A(n5847), .ZN(n5397) );
  NAND2_X1 U5298 ( .A1(n5375), .A2(n5397), .ZN(n5385) );
  INV_X1 U5299 ( .A(n5380), .ZN(n4283) );
  NOR3_X1 U5300 ( .A1(n4283), .A2(REIP_REG_30__SCAN_IN), .A3(n6520), .ZN(n4284) );
  NOR2_X1 U5301 ( .A1(n5791), .A2(STATE2_REG_1__SCAN_IN), .ZN(n5071) );
  AOI21_X1 U5302 ( .B1(n4289), .B2(MEMORYFETCH_REG_SCAN_IN), .A(n5071), .ZN(
        n4290) );
  NAND2_X1 U5303 ( .A1(n4399), .A2(n4290), .ZN(U2788) );
  INV_X1 U5304 ( .A(n4296), .ZN(n4292) );
  OAI22_X1 U5305 ( .A1(n4320), .A2(n3154), .B1(n4292), .B2(n4291), .ZN(n5967)
         );
  INV_X1 U5306 ( .A(n4293), .ZN(n5206) );
  OR2_X1 U5307 ( .A1(n5206), .A2(n4294), .ZN(n4306) );
  AOI21_X1 U5308 ( .B1(n4306), .B2(n6461), .A(READY_N), .ZN(n6558) );
  NOR2_X1 U5309 ( .A1(n5967), .A2(n6558), .ZN(n6425) );
  INV_X1 U5310 ( .A(n6440), .ZN(n6447) );
  NOR2_X1 U5311 ( .A1(n6425), .A2(n6447), .ZN(n5974) );
  INV_X1 U5312 ( .A(MORE_REG_SCAN_IN), .ZN(n4304) );
  INV_X1 U5313 ( .A(n4320), .ZN(n4302) );
  INV_X1 U5314 ( .A(n4295), .ZN(n4328) );
  NAND3_X1 U5315 ( .A1(n4327), .A2(n4296), .A3(n6396), .ZN(n4300) );
  INV_X1 U5316 ( .A(n4297), .ZN(n4298) );
  AOI22_X1 U5317 ( .A1(n4302), .A2(n4300), .B1(n4299), .B2(n4298), .ZN(n4301)
         );
  OAI21_X1 U5318 ( .B1(n4302), .B2(n4328), .A(n4301), .ZN(n6397) );
  NAND2_X1 U5319 ( .A1(n5974), .A2(n6397), .ZN(n4303) );
  OAI21_X1 U5320 ( .B1(n5974), .B2(n4304), .A(n4303), .ZN(U3471) );
  INV_X1 U5321 ( .A(n6557), .ZN(n4307) );
  OAI21_X1 U5322 ( .B1(n5071), .B2(READREQUEST_REG_SCAN_IN), .A(n4307), .ZN(
        n4305) );
  OAI21_X1 U5323 ( .B1(n4307), .B2(n4306), .A(n4305), .ZN(U3474) );
  OR2_X1 U5324 ( .A1(n4308), .A2(n6427), .ZN(n4429) );
  INV_X1 U5325 ( .A(n6404), .ZN(n4614) );
  OR2_X1 U5326 ( .A1(n4308), .A2(n4614), .ZN(n4309) );
  NAND2_X1 U5327 ( .A1(n4429), .A2(n4309), .ZN(n4310) );
  NOR2_X1 U5328 ( .A1(n6661), .A2(n6536), .ZN(n4629) );
  NAND2_X1 U5329 ( .A1(n6443), .A2(n4629), .ZN(n6110) );
  INV_X1 U5330 ( .A(n6110), .ZN(n6117) );
  INV_X1 U5331 ( .A(DATAO_REG_16__SCAN_IN), .ZN(n6596) );
  NAND2_X1 U5332 ( .A1(n6132), .A2(n4467), .ZN(n4378) );
  INV_X1 U5333 ( .A(UWORD_REG_0__SCAN_IN), .ZN(n6649) );
  OAI222_X1 U5334 ( .A1(n6119), .A2(n6596), .B1(n4378), .B2(n3899), .C1(n6649), 
        .C2(n6110), .ZN(U2907) );
  INV_X1 U5335 ( .A(DATAO_REG_28__SCAN_IN), .ZN(n4312) );
  INV_X1 U5336 ( .A(n4378), .ZN(n6108) );
  AOI22_X1 U5337 ( .A1(n6108), .A2(EAX_REG_28__SCAN_IN), .B1(n6553), .B2(
        UWORD_REG_12__SCAN_IN), .ZN(n4311) );
  OAI21_X1 U5338 ( .B1(n6119), .B2(n4312), .A(n4311), .ZN(U2895) );
  OR2_X1 U5339 ( .A1(n4320), .A2(n4328), .ZN(n4390) );
  OAI21_X1 U5340 ( .B1(n4313), .B2(n4409), .A(n4334), .ZN(n4314) );
  OAI21_X1 U5341 ( .B1(n4614), .B2(n6461), .A(n4314), .ZN(n4315) );
  NAND3_X1 U5342 ( .A1(n4320), .A2(n6554), .A3(n4315), .ZN(n4316) );
  NAND4_X1 U5343 ( .A1(n4390), .A2(n4318), .A3(n4317), .A4(n4316), .ZN(n4324)
         );
  NAND2_X1 U5344 ( .A1(n4320), .A2(n4319), .ZN(n4323) );
  INV_X1 U5345 ( .A(n4336), .ZN(n5960) );
  NAND2_X1 U5346 ( .A1(n5960), .A2(n4321), .ZN(n4322) );
  NAND2_X1 U5347 ( .A1(n4323), .A2(n4322), .ZN(n4403) );
  OR2_X1 U5348 ( .A1(n4324), .A2(n4403), .ZN(n4622) );
  INV_X1 U5349 ( .A(FLUSH_REG_SCAN_IN), .ZN(n6647) );
  NAND2_X1 U5350 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n4629), .ZN(n6529) );
  NOR2_X1 U5351 ( .A1(n6647), .A2(n6529), .ZN(n4325) );
  AOI21_X1 U5352 ( .B1(n6440), .B2(n4622), .A(n4325), .ZN(n5965) );
  NAND2_X1 U5353 ( .A1(n6443), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6530) );
  NAND2_X1 U5354 ( .A1(n5965), .A2(n6530), .ZN(n6540) );
  OAI21_X1 U5355 ( .B1(n2986), .B2(n6533), .A(n6540), .ZN(n4347) );
  OAI22_X1 U5356 ( .A1(n4413), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .B1(n4326), .B2(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4386) );
  INV_X1 U5357 ( .A(n4386), .ZN(n4345) );
  NAND2_X1 U5358 ( .A1(STATE2_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4385) );
  NAND2_X1 U5359 ( .A1(n4328), .A2(n4327), .ZN(n4604) );
  XNOR2_X1 U5360 ( .A(n2986), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4341)
         );
  XNOR2_X1 U5361 ( .A(n4607), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4329)
         );
  OAI22_X1 U5362 ( .A1(n4614), .A2(n4329), .B1(n4612), .B2(n4341), .ZN(n4340)
         );
  INV_X1 U5363 ( .A(n5208), .ZN(n5790) );
  NAND2_X1 U5364 ( .A1(n4332), .A2(n4331), .ZN(n4333) );
  NOR2_X1 U5365 ( .A1(n4334), .A2(n4333), .ZN(n4335) );
  NAND2_X1 U5366 ( .A1(n4336), .A2(n4335), .ZN(n4338) );
  NOR2_X1 U5367 ( .A1(n4338), .A2(n4337), .ZN(n4380) );
  NOR2_X1 U5368 ( .A1(n5790), .A2(n4380), .ZN(n4339) );
  AOI211_X1 U5369 ( .C1(n4604), .C2(n4341), .A(n4340), .B(n4339), .ZN(n4603)
         );
  OR2_X1 U5370 ( .A1(n4603), .A2(n6542), .ZN(n4344) );
  INV_X1 U5371 ( .A(n6533), .ZN(n4342) );
  NAND3_X1 U5372 ( .A1(n2986), .A2(n3180), .A3(n4342), .ZN(n4343) );
  OAI211_X1 U5373 ( .C1(n4345), .C2(n4385), .A(n4344), .B(n4343), .ZN(n4346)
         );
  AOI22_X1 U5374 ( .A1(n4347), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(n6540), .B2(n4346), .ZN(n4348) );
  INV_X1 U5375 ( .A(n4348), .ZN(U3459) );
  XNOR2_X1 U5376 ( .A(n4349), .B(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4428)
         );
  OAI21_X1 U5377 ( .B1(n4351), .B2(INSTADDRPOINTER_REG_0__SCAN_IN), .A(n4350), 
        .ZN(n5255) );
  INV_X1 U5378 ( .A(n5255), .ZN(n4354) );
  INV_X1 U5379 ( .A(REIP_REG_0__SCAN_IN), .ZN(n6549) );
  NOR2_X1 U5380 ( .A1(n6248), .A2(n6549), .ZN(n4352) );
  AOI211_X1 U5381 ( .C1(n6280), .C2(n4354), .A(n4353), .B(n4352), .ZN(n4358)
         );
  INV_X1 U5382 ( .A(n5758), .ZN(n4355) );
  OAI21_X1 U5383 ( .B1(n4356), .B2(n4355), .A(INSTADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n4357) );
  OAI211_X1 U5384 ( .C1(n4428), .C2(n5780), .A(n4358), .B(n4357), .ZN(U3018)
         );
  INV_X1 U5385 ( .A(EAX_REG_25__SCAN_IN), .ZN(n4360) );
  INV_X2 U5386 ( .A(n6119), .ZN(n6136) );
  AOI22_X1 U5387 ( .A1(UWORD_REG_9__SCAN_IN), .A2(n6117), .B1(n6136), .B2(
        DATAO_REG_25__SCAN_IN), .ZN(n4359) );
  OAI21_X1 U5388 ( .B1(n4360), .B2(n4378), .A(n4359), .ZN(U2898) );
  INV_X1 U5389 ( .A(EAX_REG_22__SCAN_IN), .ZN(n6580) );
  AOI22_X1 U5390 ( .A1(UWORD_REG_6__SCAN_IN), .A2(n6117), .B1(n6136), .B2(
        DATAO_REG_22__SCAN_IN), .ZN(n4361) );
  OAI21_X1 U5391 ( .B1(n6580), .B2(n4378), .A(n4361), .ZN(U2901) );
  INV_X1 U5392 ( .A(EAX_REG_20__SCAN_IN), .ZN(n4363) );
  AOI22_X1 U5393 ( .A1(UWORD_REG_4__SCAN_IN), .A2(n6553), .B1(n6136), .B2(
        DATAO_REG_20__SCAN_IN), .ZN(n4362) );
  OAI21_X1 U5394 ( .B1(n4363), .B2(n4378), .A(n4362), .ZN(U2903) );
  INV_X1 U5395 ( .A(EAX_REG_21__SCAN_IN), .ZN(n4365) );
  AOI22_X1 U5396 ( .A1(UWORD_REG_5__SCAN_IN), .A2(n6117), .B1(n6136), .B2(
        DATAO_REG_21__SCAN_IN), .ZN(n4364) );
  OAI21_X1 U5397 ( .B1(n4365), .B2(n4378), .A(n4364), .ZN(U2902) );
  INV_X1 U5398 ( .A(EAX_REG_24__SCAN_IN), .ZN(n4367) );
  AOI22_X1 U5399 ( .A1(UWORD_REG_8__SCAN_IN), .A2(n6117), .B1(n6136), .B2(
        DATAO_REG_24__SCAN_IN), .ZN(n4366) );
  OAI21_X1 U5400 ( .B1(n4367), .B2(n4378), .A(n4366), .ZN(U2899) );
  INV_X1 U5401 ( .A(EAX_REG_17__SCAN_IN), .ZN(n4369) );
  AOI22_X1 U5402 ( .A1(UWORD_REG_1__SCAN_IN), .A2(n6553), .B1(n6136), .B2(
        DATAO_REG_17__SCAN_IN), .ZN(n4368) );
  OAI21_X1 U5403 ( .B1(n4369), .B2(n4378), .A(n4368), .ZN(U2906) );
  INV_X1 U5404 ( .A(EAX_REG_18__SCAN_IN), .ZN(n6599) );
  AOI22_X1 U5405 ( .A1(UWORD_REG_2__SCAN_IN), .A2(n6553), .B1(n6136), .B2(
        DATAO_REG_18__SCAN_IN), .ZN(n4370) );
  OAI21_X1 U5406 ( .B1(n6599), .B2(n4378), .A(n4370), .ZN(U2905) );
  INV_X1 U5407 ( .A(EAX_REG_19__SCAN_IN), .ZN(n4372) );
  AOI22_X1 U5408 ( .A1(UWORD_REG_3__SCAN_IN), .A2(n6117), .B1(n6136), .B2(
        DATAO_REG_19__SCAN_IN), .ZN(n4371) );
  OAI21_X1 U5409 ( .B1(n4372), .B2(n4378), .A(n4371), .ZN(U2904) );
  INV_X1 U5410 ( .A(EAX_REG_30__SCAN_IN), .ZN(n4374) );
  AOI22_X1 U5411 ( .A1(UWORD_REG_14__SCAN_IN), .A2(n6553), .B1(n6136), .B2(
        DATAO_REG_30__SCAN_IN), .ZN(n4373) );
  OAI21_X1 U5412 ( .B1(n4374), .B2(n4378), .A(n4373), .ZN(U2893) );
  INV_X1 U5413 ( .A(EAX_REG_26__SCAN_IN), .ZN(n4376) );
  AOI22_X1 U5414 ( .A1(UWORD_REG_10__SCAN_IN), .A2(n6553), .B1(n6136), .B2(
        DATAO_REG_26__SCAN_IN), .ZN(n4375) );
  OAI21_X1 U5415 ( .B1(n4376), .B2(n4378), .A(n4375), .ZN(U2897) );
  INV_X1 U5416 ( .A(EAX_REG_29__SCAN_IN), .ZN(n4379) );
  AOI22_X1 U5417 ( .A1(UWORD_REG_13__SCAN_IN), .A2(n6117), .B1(n6136), .B2(
        DATAO_REG_29__SCAN_IN), .ZN(n4377) );
  OAI21_X1 U5418 ( .B1(n4379), .B2(n4378), .A(n4377), .ZN(U2894) );
  INV_X1 U5419 ( .A(n5785), .ZN(n6070) );
  INV_X1 U5420 ( .A(n4380), .ZN(n6402) );
  OAI21_X1 U5421 ( .B1(n4381), .B2(n4384), .A(n6401), .ZN(n4382) );
  OAI21_X1 U5422 ( .B1(n4614), .B2(n4607), .A(n4382), .ZN(n4383) );
  AOI21_X1 U5423 ( .B1(n6070), .B2(n6402), .A(n4383), .ZN(n6406) );
  INV_X1 U5424 ( .A(n4384), .ZN(n4387) );
  OAI222_X1 U5425 ( .A1(n6542), .A2(n6406), .B1(n4387), .B2(n6533), .C1(n4386), 
        .C2(n4385), .ZN(n4388) );
  OAI21_X1 U5426 ( .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n6533), .A(n6540), 
        .ZN(n6538) );
  AOI22_X1 U5427 ( .A1(n6540), .A2(n4388), .B1(n4607), .B2(n6538), .ZN(n4389)
         );
  INV_X1 U5428 ( .A(n4389), .ZN(U3460) );
  NOR2_X1 U5429 ( .A1(n4390), .A2(n6447), .ZN(n4395) );
  INV_X1 U5430 ( .A(n3126), .ZN(n4393) );
  NOR2_X1 U5431 ( .A1(n3146), .A2(n6429), .ZN(n4391) );
  NAND4_X1 U5432 ( .A1(n4393), .A2(n4392), .A3(n3167), .A4(n4391), .ZN(n4401)
         );
  NOR2_X1 U5433 ( .A1(n4401), .A2(n2964), .ZN(n4394) );
  OR2_X2 U5434 ( .A1(n4395), .A2(n4394), .ZN(n6096) );
  NAND2_X1 U5435 ( .A1(n6096), .A2(n5473), .ZN(n6091) );
  AND2_X1 U5436 ( .A1(n6096), .A2(n3146), .ZN(n6088) );
  INV_X2 U5437 ( .A(n6088), .ZN(n6092) );
  XNOR2_X1 U5438 ( .A(n4397), .B(n4396), .ZN(n5260) );
  INV_X1 U5439 ( .A(EBX_REG_0__SCAN_IN), .ZN(n4398) );
  OAI222_X1 U5440 ( .A1(n5255), .A2(n6091), .B1(n6092), .B2(n5260), .C1(n4398), 
        .C2(n6096), .ZN(U2859) );
  NOR2_X1 U5441 ( .A1(n4399), .A2(READY_N), .ZN(n4430) );
  NAND2_X1 U5442 ( .A1(n4430), .A2(n4494), .ZN(n4551) );
  NOR2_X1 U5443 ( .A1(n4401), .A2(n4400), .ZN(n4402) );
  AOI21_X1 U5444 ( .B1(n4403), .B2(n6440), .A(n4402), .ZN(n4404) );
  INV_X1 U5445 ( .A(DATAI_0_), .ZN(n6656) );
  INV_X1 U5446 ( .A(EAX_REG_0__SCAN_IN), .ZN(n6673) );
  OAI222_X1 U5447 ( .A1(n5914), .A2(n5260), .B1(n5203), .B2(n6656), .C1(n5472), 
        .C2(n6673), .ZN(U2891) );
  XNOR2_X1 U5448 ( .A(n4407), .B(n4406), .ZN(n4445) );
  NAND3_X1 U5449 ( .A1(n6210), .A2(n4413), .A3(n4408), .ZN(n4416) );
  OR2_X1 U5450 ( .A1(n4410), .A2(n4409), .ZN(n4412) );
  AND2_X1 U5451 ( .A1(n4412), .A2(n4411), .ZN(n6086) );
  INV_X1 U5452 ( .A(n6086), .ZN(n4433) );
  INV_X1 U5453 ( .A(REIP_REG_1__SCAN_IN), .ZN(n6573) );
  OAI22_X1 U5454 ( .A1(n6248), .A2(n6573), .B1(n4708), .B2(n4413), .ZN(n4414)
         );
  AOI21_X1 U5455 ( .B1(n6280), .B2(n4433), .A(n4414), .ZN(n4415) );
  OAI211_X1 U5456 ( .C1(n4445), .C2(n5780), .A(n4416), .B(n4415), .ZN(U3017)
         );
  NAND2_X1 U5457 ( .A1(n5783), .A2(n2965), .ZN(n4419) );
  NAND2_X1 U5458 ( .A1(n4419), .A2(n4418), .ZN(n4421) );
  NOR2_X1 U5459 ( .A1(n4421), .A2(n4420), .ZN(n4422) );
  NOR2_X1 U5460 ( .A1(n3712), .A2(n4422), .ZN(n6072) );
  INV_X1 U5461 ( .A(n6072), .ZN(n4435) );
  INV_X1 U5462 ( .A(DATAI_1_), .ZN(n4493) );
  INV_X1 U5463 ( .A(EAX_REG_1__SCAN_IN), .ZN(n6135) );
  OAI222_X1 U5464 ( .A1(n4435), .A2(n5914), .B1(n5203), .B2(n4493), .C1(n5472), 
        .C2(n6135), .ZN(U2890) );
  NAND2_X1 U5465 ( .A1(n5618), .A2(n4423), .ZN(n4424) );
  AOI22_X1 U5466 ( .A1(n4424), .A2(PHYADDRPOINTER_REG_0__SCAN_IN), .B1(n3668), 
        .B2(REIP_REG_0__SCAN_IN), .ZN(n4427) );
  INV_X1 U5467 ( .A(n5260), .ZN(n4425) );
  INV_X1 U5468 ( .A(n5634), .ZN(n6165) );
  NAND2_X1 U5469 ( .A1(n4425), .A2(n6165), .ZN(n4426) );
  OAI211_X1 U5470 ( .C1(n4428), .C2(n6169), .A(n4427), .B(n4426), .ZN(U2986)
         );
  OR2_X1 U5471 ( .A1(n4430), .A2(n4572), .ZN(n6146) );
  INV_X1 U5472 ( .A(LWORD_REG_15__SCAN_IN), .ZN(n4432) );
  INV_X1 U5473 ( .A(n4551), .ZN(n6143) );
  AOI22_X1 U5474 ( .A1(n6143), .A2(DATAI_15_), .B1(EAX_REG_15__SCAN_IN), .B2(
        n4572), .ZN(n4431) );
  OAI21_X1 U5475 ( .B1(n6146), .B2(n4432), .A(n4431), .ZN(U2954) );
  INV_X1 U5476 ( .A(n6091), .ZN(n6087) );
  INV_X1 U5477 ( .A(n6096), .ZN(n5462) );
  AOI22_X1 U5478 ( .A1(n6087), .A2(n4433), .B1(n5462), .B2(EBX_REG_1__SCAN_IN), 
        .ZN(n4434) );
  OAI21_X1 U5479 ( .B1(n4435), .B2(n6092), .A(n4434), .ZN(U2858) );
  INV_X1 U5480 ( .A(n3712), .ZN(n4437) );
  NAND3_X1 U5481 ( .A1(n4439), .A2(n4438), .A3(n4437), .ZN(n4440) );
  AND2_X1 U5482 ( .A1(n4436), .A2(n4440), .ZN(n6190) );
  INV_X1 U5483 ( .A(n6190), .ZN(n5216) );
  XNOR2_X1 U5484 ( .A(n4449), .B(n4451), .ZN(n6279) );
  AOI22_X1 U5485 ( .A1(n6087), .A2(n6279), .B1(n5462), .B2(EBX_REG_2__SCAN_IN), 
        .ZN(n4441) );
  OAI21_X1 U5486 ( .B1(n5216), .B2(n6092), .A(n4441), .ZN(U2857) );
  AOI22_X1 U5487 ( .A1(n6186), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .B1(n3668), 
        .B2(REIP_REG_1__SCAN_IN), .ZN(n4442) );
  OAI21_X1 U5488 ( .B1(n6195), .B2(PHYADDRPOINTER_REG_1__SCAN_IN), .A(n4442), 
        .ZN(n4443) );
  AOI21_X1 U5489 ( .B1(n6072), .B2(n6165), .A(n4443), .ZN(n4444) );
  OAI21_X1 U5490 ( .B1(n4445), .B2(n6169), .A(n4444), .ZN(U2985) );
  AND2_X1 U5491 ( .A1(n4446), .A2(n4436), .ZN(n4448) );
  OR2_X1 U5492 ( .A1(n4448), .A2(n4447), .ZN(n6057) );
  INV_X1 U5493 ( .A(n4449), .ZN(n4452) );
  AOI21_X1 U5494 ( .B1(n4452), .B2(n4451), .A(n4450), .ZN(n4453) );
  NOR2_X1 U5495 ( .A1(n4453), .A2(n4577), .ZN(n6266) );
  AOI22_X1 U5496 ( .A1(n6087), .A2(n6266), .B1(n5462), .B2(EBX_REG_3__SCAN_IN), 
        .ZN(n4454) );
  OAI21_X1 U5497 ( .B1(n6057), .B2(n6092), .A(n4454), .ZN(U2856) );
  AOI22_X1 U5498 ( .A1(n5499), .A2(DATAI_2_), .B1(n6103), .B2(
        EAX_REG_2__SCAN_IN), .ZN(n4455) );
  OAI21_X1 U5499 ( .B1(n5216), .B2(n5914), .A(n4455), .ZN(U2889) );
  NAND2_X1 U5500 ( .A1(n4732), .A2(n4652), .ZN(n4655) );
  INV_X1 U5501 ( .A(n4655), .ZN(n4589) );
  NOR2_X1 U5502 ( .A1(n5783), .A2(n5973), .ZN(n4802) );
  AOI21_X1 U5503 ( .B1(n4589), .B2(n4802), .A(n5791), .ZN(n4462) );
  NAND2_X1 U5504 ( .A1(n5208), .A2(n5785), .ZN(n4933) );
  OR2_X1 U5505 ( .A1(n4933), .A2(n4623), .ZN(n4987) );
  INV_X1 U5506 ( .A(n6403), .ZN(n5254) );
  OR2_X1 U5507 ( .A1(n4987), .A2(n5254), .ZN(n4458) );
  NAND3_X1 U5508 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n6419), .A3(n6612), .ZN(n4985) );
  OR2_X1 U5509 ( .A1(n4929), .A2(n4985), .ZN(n4500) );
  NAND2_X1 U5510 ( .A1(n4458), .A2(n4500), .ZN(n4460) );
  INV_X1 U5511 ( .A(n4985), .ZN(n4459) );
  AOI22_X1 U5512 ( .A1(n4462), .A2(n4460), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n4459), .ZN(n4504) );
  NOR2_X1 U5513 ( .A1(n6656), .A2(n4991), .ZN(n6376) );
  INV_X1 U5514 ( .A(n6376), .ZN(n5807) );
  AOI21_X1 U5515 ( .B1(n4929), .B2(STATE2_REG_3__SCAN_IN), .A(n4991), .ZN(
        n4833) );
  INV_X1 U5516 ( .A(n4460), .ZN(n4461) );
  AOI22_X1 U5517 ( .A1(n4462), .A2(n4461), .B1(n4985), .B2(n5791), .ZN(n4463)
         );
  NAND2_X1 U5518 ( .A1(n4833), .A2(n4463), .ZN(n4498) );
  NAND2_X1 U5519 ( .A1(n4498), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n4470) );
  INV_X1 U5520 ( .A(n5026), .ZN(n4986) );
  AND2_X1 U5521 ( .A1(n5593), .A2(DATAI_24_), .ZN(n6310) );
  NAND2_X1 U5522 ( .A1(n5593), .A2(DATAI_16_), .ZN(n6379) );
  INV_X1 U5523 ( .A(n6530), .ZN(n4466) );
  NAND2_X1 U5524 ( .A1(n4499), .A2(n4467), .ZN(n5173) );
  OAI22_X1 U5525 ( .A1(n4920), .A2(n6379), .B1(n5173), .B2(n4500), .ZN(n4468)
         );
  AOI21_X1 U5526 ( .B1(n4986), .B2(n6310), .A(n4468), .ZN(n4469) );
  OAI211_X1 U5527 ( .C1(n4504), .C2(n5807), .A(n4470), .B(n4469), .ZN(U3060)
         );
  OAI21_X1 U5528 ( .B1(n4447), .B2(n4472), .A(n4968), .ZN(n6046) );
  INV_X1 U5529 ( .A(DATAI_4_), .ZN(n4485) );
  INV_X1 U5530 ( .A(EAX_REG_4__SCAN_IN), .ZN(n6129) );
  OAI222_X1 U5531 ( .A1(n6046), .A2(n5914), .B1(n5203), .B2(n4485), .C1(n5472), 
        .C2(n6129), .ZN(U2887) );
  INV_X1 U5532 ( .A(DATAI_3_), .ZN(n4538) );
  NOR2_X1 U5533 ( .A1(n4538), .A2(n4991), .ZN(n6348) );
  INV_X1 U5534 ( .A(n6348), .ZN(n5820) );
  NAND2_X1 U5535 ( .A1(n4498), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4476) );
  NAND2_X1 U5536 ( .A1(n5593), .A2(DATAI_19_), .ZN(n5150) );
  INV_X1 U5537 ( .A(n5150), .ZN(n6347) );
  NAND2_X1 U5538 ( .A1(n5593), .A2(DATAI_27_), .ZN(n6351) );
  NAND2_X1 U5539 ( .A1(n4499), .A2(n4473), .ZN(n5149) );
  OAI22_X1 U5540 ( .A1(n5026), .A2(n6351), .B1(n5149), .B2(n4500), .ZN(n4474)
         );
  AOI21_X1 U5541 ( .B1(n6347), .B2(n6318), .A(n4474), .ZN(n4475) );
  OAI211_X1 U5542 ( .C1(n4504), .C2(n5820), .A(n4476), .B(n4475), .ZN(U3063)
         );
  INV_X1 U5543 ( .A(DATAI_6_), .ZN(n6733) );
  NOR2_X1 U5544 ( .A1(n6733), .A2(n4991), .ZN(n6360) );
  INV_X1 U5545 ( .A(n6360), .ZN(n5832) );
  NAND2_X1 U5546 ( .A1(n4498), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4480) );
  NAND2_X1 U5547 ( .A1(n5593), .A2(DATAI_22_), .ZN(n5162) );
  INV_X1 U5548 ( .A(n5162), .ZN(n6359) );
  NAND2_X1 U5549 ( .A1(n5593), .A2(DATAI_30_), .ZN(n6363) );
  NAND2_X1 U5550 ( .A1(n4499), .A2(n4477), .ZN(n5161) );
  OAI22_X1 U5551 ( .A1(n5026), .A2(n6363), .B1(n5161), .B2(n4500), .ZN(n4478)
         );
  AOI21_X1 U5552 ( .B1(n6359), .B2(n6318), .A(n4478), .ZN(n4479) );
  OAI211_X1 U5553 ( .C1(n4504), .C2(n5832), .A(n4480), .B(n4479), .ZN(U3066)
         );
  INV_X1 U5554 ( .A(DATAI_5_), .ZN(n4973) );
  NOR2_X1 U5555 ( .A1(n4973), .A2(n4991), .ZN(n6354) );
  INV_X1 U5556 ( .A(n6354), .ZN(n5828) );
  NAND2_X1 U5557 ( .A1(n4498), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4484) );
  NAND2_X1 U5558 ( .A1(n5593), .A2(DATAI_21_), .ZN(n5156) );
  INV_X1 U5559 ( .A(n5156), .ZN(n6353) );
  NAND2_X1 U5560 ( .A1(n5593), .A2(DATAI_29_), .ZN(n6357) );
  NAND2_X1 U5561 ( .A1(n4499), .A2(n4481), .ZN(n5155) );
  OAI22_X1 U5562 ( .A1(n5026), .A2(n6357), .B1(n5155), .B2(n4500), .ZN(n4482)
         );
  AOI21_X1 U5563 ( .B1(n6353), .B2(n6318), .A(n4482), .ZN(n4483) );
  OAI211_X1 U5564 ( .C1(n4504), .C2(n5828), .A(n4484), .B(n4483), .ZN(U3065)
         );
  NOR2_X1 U5565 ( .A1(n4485), .A2(n4991), .ZN(n6298) );
  INV_X1 U5566 ( .A(n6298), .ZN(n5824) );
  NAND2_X1 U5567 ( .A1(n4498), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4489) );
  NAND2_X1 U5568 ( .A1(n5593), .A2(DATAI_20_), .ZN(n5144) );
  INV_X1 U5569 ( .A(n5144), .ZN(n6297) );
  NAND2_X1 U5570 ( .A1(n5593), .A2(DATAI_28_), .ZN(n6301) );
  NAND2_X1 U5571 ( .A1(n4499), .A2(n4486), .ZN(n5143) );
  OAI22_X1 U5572 ( .A1(n5026), .A2(n6301), .B1(n5143), .B2(n4500), .ZN(n4487)
         );
  AOI21_X1 U5573 ( .B1(n6297), .B2(n6318), .A(n4487), .ZN(n4488) );
  OAI211_X1 U5574 ( .C1(n4504), .C2(n5824), .A(n4489), .B(n4488), .ZN(U3064)
         );
  INV_X1 U5575 ( .A(DATAI_2_), .ZN(n4542) );
  NOR2_X1 U5576 ( .A1(n4542), .A2(n4991), .ZN(n6327) );
  INV_X1 U5577 ( .A(n6327), .ZN(n5816) );
  NAND2_X1 U5578 ( .A1(n4498), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4492) );
  NAND2_X1 U5579 ( .A1(n5593), .A2(DATAI_18_), .ZN(n6323) );
  INV_X1 U5580 ( .A(n6323), .ZN(n6326) );
  NAND2_X1 U5581 ( .A1(n5593), .A2(DATAI_26_), .ZN(n6330) );
  NAND2_X1 U5582 ( .A1(n4499), .A2(n3124), .ZN(n5183) );
  OAI22_X1 U5583 ( .A1(n5026), .A2(n6330), .B1(n5183), .B2(n4500), .ZN(n4490)
         );
  AOI21_X1 U5584 ( .B1(n6326), .B2(n6318), .A(n4490), .ZN(n4491) );
  OAI211_X1 U5585 ( .C1(n4504), .C2(n5816), .A(n4492), .B(n4491), .ZN(U3062)
         );
  NOR2_X1 U5586 ( .A1(n4493), .A2(n4991), .ZN(n6386) );
  INV_X1 U5587 ( .A(n6386), .ZN(n5812) );
  NAND2_X1 U5588 ( .A1(n4498), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n4497) );
  NAND2_X1 U5589 ( .A1(n5593), .A2(DATAI_17_), .ZN(n6390) );
  INV_X1 U5590 ( .A(n6390), .ZN(n6343) );
  NAND2_X1 U5591 ( .A1(n5593), .A2(DATAI_25_), .ZN(n6387) );
  NAND2_X1 U5592 ( .A1(n4499), .A2(n4494), .ZN(n5177) );
  OAI22_X1 U5593 ( .A1(n5026), .A2(n6387), .B1(n5177), .B2(n4500), .ZN(n4495)
         );
  AOI21_X1 U5594 ( .B1(n6343), .B2(n6318), .A(n4495), .ZN(n4496) );
  OAI211_X1 U5595 ( .C1(n4504), .C2(n5812), .A(n4497), .B(n4496), .ZN(U3061)
         );
  INV_X1 U5596 ( .A(DATAI_7_), .ZN(n6632) );
  NOR2_X1 U5597 ( .A1(n6632), .A2(n4991), .ZN(n6369) );
  INV_X1 U5598 ( .A(n6369), .ZN(n5839) );
  NAND2_X1 U5599 ( .A1(n4498), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4503) );
  NAND2_X1 U5600 ( .A1(n5593), .A2(DATAI_23_), .ZN(n5168) );
  INV_X1 U5601 ( .A(n5168), .ZN(n6366) );
  NAND2_X1 U5602 ( .A1(n5593), .A2(DATAI_31_), .ZN(n6374) );
  NAND2_X1 U5603 ( .A1(n4499), .A2(n3146), .ZN(n5167) );
  OAI22_X1 U5604 ( .A1(n5026), .A2(n6374), .B1(n5167), .B2(n4500), .ZN(n4501)
         );
  AOI21_X1 U5605 ( .B1(n6366), .B2(n6318), .A(n4501), .ZN(n4502) );
  OAI211_X1 U5606 ( .C1(n4504), .C2(n5839), .A(n4503), .B(n4502), .ZN(U3067)
         );
  AND2_X1 U5607 ( .A1(n6059), .A2(n6403), .ZN(n4801) );
  NAND2_X1 U5608 ( .A1(n5208), .A2(n6070), .ZN(n4765) );
  INV_X1 U5609 ( .A(n4765), .ZN(n4506) );
  INV_X1 U5610 ( .A(n4580), .ZN(n6384) );
  AOI21_X1 U5611 ( .B1(n4801), .B2(n4506), .A(n6384), .ZN(n4512) );
  INV_X1 U5612 ( .A(n4652), .ZN(n4507) );
  AND2_X1 U5613 ( .A1(n4507), .A2(n5783), .ZN(n4508) );
  NAND2_X1 U5614 ( .A1(n4732), .A2(n4508), .ZN(n4516) );
  INV_X1 U5615 ( .A(n4516), .ZN(n4509) );
  INV_X1 U5616 ( .A(n5791), .ZN(n5797) );
  NAND2_X1 U5617 ( .A1(n5797), .A2(n5973), .ZN(n5800) );
  OAI21_X1 U5618 ( .B1(n4509), .B2(n5634), .A(n5800), .ZN(n4511) );
  NOR2_X1 U5619 ( .A1(n5797), .A2(n4513), .ZN(n4510) );
  INV_X1 U5620 ( .A(n4833), .ZN(n4739) );
  AOI211_X1 U5621 ( .C1(n4512), .C2(n4511), .A(n4510), .B(n4739), .ZN(n6395)
         );
  INV_X1 U5622 ( .A(n6395), .ZN(n4536) );
  OR2_X1 U5623 ( .A1(n4512), .A2(n5791), .ZN(n4515) );
  NAND2_X1 U5624 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n4513), .ZN(n4514) );
  NAND2_X1 U5625 ( .A1(n4515), .A2(n4514), .ZN(n6385) );
  INV_X1 U5626 ( .A(n5143), .ZN(n6296) );
  AOI22_X1 U5627 ( .A1(n6298), .A2(n6385), .B1(n6384), .B2(n6296), .ZN(n4518)
         );
  OR2_X1 U5628 ( .A1(n4516), .A2(n4808), .ZN(n6388) );
  INV_X1 U5629 ( .A(n6301), .ZN(n5146) );
  NAND2_X1 U5630 ( .A1(n4794), .A2(n5146), .ZN(n4517) );
  OAI211_X1 U5631 ( .C1(n6391), .C2(n5144), .A(n4518), .B(n4517), .ZN(n4519)
         );
  AOI21_X1 U5632 ( .B1(n4536), .B2(INSTQUEUE_REG_15__4__SCAN_IN), .A(n4519), 
        .ZN(n4520) );
  INV_X1 U5633 ( .A(n4520), .ZN(U3144) );
  INV_X1 U5634 ( .A(n5155), .ZN(n6352) );
  AOI22_X1 U5635 ( .A1(n6354), .A2(n6385), .B1(n6384), .B2(n6352), .ZN(n4522)
         );
  INV_X1 U5636 ( .A(n6357), .ZN(n5158) );
  NAND2_X1 U5637 ( .A1(n4794), .A2(n5158), .ZN(n4521) );
  OAI211_X1 U5638 ( .C1(n6391), .C2(n5156), .A(n4522), .B(n4521), .ZN(n4523)
         );
  AOI21_X1 U5639 ( .B1(n4536), .B2(INSTQUEUE_REG_15__5__SCAN_IN), .A(n4523), 
        .ZN(n4524) );
  INV_X1 U5640 ( .A(n4524), .ZN(U3145) );
  INV_X1 U5641 ( .A(n5161), .ZN(n6358) );
  AOI22_X1 U5642 ( .A1(n6360), .A2(n6385), .B1(n6384), .B2(n6358), .ZN(n4526)
         );
  INV_X1 U5643 ( .A(n6363), .ZN(n5164) );
  NAND2_X1 U5644 ( .A1(n4794), .A2(n5164), .ZN(n4525) );
  OAI211_X1 U5645 ( .C1(n6391), .C2(n5162), .A(n4526), .B(n4525), .ZN(n4527)
         );
  AOI21_X1 U5646 ( .B1(n4536), .B2(INSTQUEUE_REG_15__6__SCAN_IN), .A(n4527), 
        .ZN(n4528) );
  INV_X1 U5647 ( .A(n4528), .ZN(U3146) );
  INV_X1 U5648 ( .A(n5149), .ZN(n6346) );
  AOI22_X1 U5649 ( .A1(n6348), .A2(n6385), .B1(n6384), .B2(n6346), .ZN(n4530)
         );
  INV_X1 U5650 ( .A(n6351), .ZN(n5152) );
  NAND2_X1 U5651 ( .A1(n4794), .A2(n5152), .ZN(n4529) );
  OAI211_X1 U5652 ( .C1(n6391), .C2(n5150), .A(n4530), .B(n4529), .ZN(n4531)
         );
  AOI21_X1 U5653 ( .B1(n4536), .B2(INSTQUEUE_REG_15__3__SCAN_IN), .A(n4531), 
        .ZN(n4532) );
  INV_X1 U5654 ( .A(n4532), .ZN(U3143) );
  INV_X1 U5655 ( .A(n5167), .ZN(n6365) );
  AOI22_X1 U5656 ( .A1(n6369), .A2(n6385), .B1(n6384), .B2(n6365), .ZN(n4534)
         );
  INV_X1 U5657 ( .A(n6374), .ZN(n5170) );
  NAND2_X1 U5658 ( .A1(n4794), .A2(n5170), .ZN(n4533) );
  OAI211_X1 U5659 ( .C1(n6391), .C2(n5168), .A(n4534), .B(n4533), .ZN(n4535)
         );
  AOI21_X1 U5660 ( .B1(n4536), .B2(INSTQUEUE_REG_15__7__SCAN_IN), .A(n4535), 
        .ZN(n4537) );
  INV_X1 U5661 ( .A(n4537), .ZN(U3147) );
  INV_X1 U5662 ( .A(EAX_REG_3__SCAN_IN), .ZN(n6131) );
  OAI222_X1 U5663 ( .A1(n6057), .A2(n5914), .B1(n5203), .B2(n4538), .C1(n5472), 
        .C2(n6131), .ZN(U2888) );
  INV_X2 U5664 ( .A(n6146), .ZN(n6153) );
  AOI22_X1 U5665 ( .A1(n6153), .A2(LWORD_REG_7__SCAN_IN), .B1(
        EAX_REG_7__SCAN_IN), .B2(n4572), .ZN(n4539) );
  NAND2_X1 U5666 ( .A1(n6143), .A2(DATAI_7_), .ZN(n4556) );
  NAND2_X1 U5667 ( .A1(n4539), .A2(n4556), .ZN(U2946) );
  AOI22_X1 U5668 ( .A1(n6153), .A2(UWORD_REG_5__SCAN_IN), .B1(
        EAX_REG_21__SCAN_IN), .B2(n4572), .ZN(n4540) );
  NAND2_X1 U5669 ( .A1(n6143), .A2(DATAI_5_), .ZN(n4548) );
  NAND2_X1 U5670 ( .A1(n4540), .A2(n4548), .ZN(U2929) );
  AOI22_X1 U5671 ( .A1(n6153), .A2(UWORD_REG_13__SCAN_IN), .B1(
        EAX_REG_29__SCAN_IN), .B2(n4572), .ZN(n4541) );
  INV_X1 U5672 ( .A(DATAI_13_), .ZN(n4704) );
  OR2_X1 U5673 ( .A1(n4551), .A2(n4704), .ZN(n4562) );
  NAND2_X1 U5674 ( .A1(n4541), .A2(n4562), .ZN(U2937) );
  AOI22_X1 U5675 ( .A1(n6153), .A2(UWORD_REG_2__SCAN_IN), .B1(
        EAX_REG_18__SCAN_IN), .B2(n4572), .ZN(n4543) );
  OR2_X1 U5676 ( .A1(n4551), .A2(n4542), .ZN(n4570) );
  NAND2_X1 U5677 ( .A1(n4543), .A2(n4570), .ZN(U2926) );
  AOI22_X1 U5678 ( .A1(n6153), .A2(UWORD_REG_9__SCAN_IN), .B1(
        EAX_REG_25__SCAN_IN), .B2(n4572), .ZN(n4544) );
  NAND2_X1 U5679 ( .A1(n6143), .A2(DATAI_9_), .ZN(n4545) );
  NAND2_X1 U5680 ( .A1(n4544), .A2(n4545), .ZN(U2933) );
  AOI22_X1 U5681 ( .A1(n6153), .A2(LWORD_REG_9__SCAN_IN), .B1(
        EAX_REG_9__SCAN_IN), .B2(n4572), .ZN(n4546) );
  NAND2_X1 U5682 ( .A1(n4546), .A2(n4545), .ZN(U2948) );
  AOI22_X1 U5683 ( .A1(n6153), .A2(LWORD_REG_4__SCAN_IN), .B1(
        EAX_REG_4__SCAN_IN), .B2(n4572), .ZN(n4547) );
  NAND2_X1 U5684 ( .A1(n6143), .A2(DATAI_4_), .ZN(n4554) );
  NAND2_X1 U5685 ( .A1(n4547), .A2(n4554), .ZN(U2943) );
  AOI22_X1 U5686 ( .A1(n6153), .A2(LWORD_REG_5__SCAN_IN), .B1(
        EAX_REG_5__SCAN_IN), .B2(n4572), .ZN(n4549) );
  NAND2_X1 U5687 ( .A1(n4549), .A2(n4548), .ZN(U2944) );
  AOI22_X1 U5688 ( .A1(n6153), .A2(LWORD_REG_6__SCAN_IN), .B1(
        EAX_REG_6__SCAN_IN), .B2(n4572), .ZN(n4550) );
  NAND2_X1 U5689 ( .A1(n6143), .A2(DATAI_6_), .ZN(n4558) );
  NAND2_X1 U5690 ( .A1(n4550), .A2(n4558), .ZN(U2945) );
  AOI22_X1 U5691 ( .A1(n6153), .A2(LWORD_REG_14__SCAN_IN), .B1(
        EAX_REG_14__SCAN_IN), .B2(n4572), .ZN(n4552) );
  INV_X1 U5692 ( .A(DATAI_14_), .ZN(n4925) );
  OR2_X1 U5693 ( .A1(n4551), .A2(n4925), .ZN(n4565) );
  NAND2_X1 U5694 ( .A1(n4552), .A2(n4565), .ZN(U2953) );
  AOI22_X1 U5695 ( .A1(n6153), .A2(UWORD_REG_3__SCAN_IN), .B1(
        EAX_REG_19__SCAN_IN), .B2(n4572), .ZN(n4553) );
  NAND2_X1 U5696 ( .A1(n6143), .A2(DATAI_3_), .ZN(n4560) );
  NAND2_X1 U5697 ( .A1(n4553), .A2(n4560), .ZN(U2927) );
  AOI22_X1 U5698 ( .A1(n6153), .A2(UWORD_REG_4__SCAN_IN), .B1(
        EAX_REG_20__SCAN_IN), .B2(n4572), .ZN(n4555) );
  NAND2_X1 U5699 ( .A1(n4555), .A2(n4554), .ZN(U2928) );
  AOI22_X1 U5700 ( .A1(n6153), .A2(UWORD_REG_7__SCAN_IN), .B1(
        EAX_REG_23__SCAN_IN), .B2(n4572), .ZN(n4557) );
  NAND2_X1 U5701 ( .A1(n4557), .A2(n4556), .ZN(U2931) );
  AOI22_X1 U5702 ( .A1(n6153), .A2(UWORD_REG_6__SCAN_IN), .B1(
        EAX_REG_22__SCAN_IN), .B2(n4572), .ZN(n4559) );
  NAND2_X1 U5703 ( .A1(n4559), .A2(n4558), .ZN(U2930) );
  AOI22_X1 U5704 ( .A1(n6153), .A2(LWORD_REG_3__SCAN_IN), .B1(
        EAX_REG_3__SCAN_IN), .B2(n4572), .ZN(n4561) );
  NAND2_X1 U5705 ( .A1(n4561), .A2(n4560), .ZN(U2942) );
  AOI22_X1 U5706 ( .A1(n6153), .A2(LWORD_REG_13__SCAN_IN), .B1(
        EAX_REG_13__SCAN_IN), .B2(n4572), .ZN(n4563) );
  NAND2_X1 U5707 ( .A1(n4563), .A2(n4562), .ZN(U2952) );
  AOI22_X1 U5708 ( .A1(n6153), .A2(UWORD_REG_0__SCAN_IN), .B1(
        EAX_REG_16__SCAN_IN), .B2(n4572), .ZN(n4564) );
  NAND2_X1 U5709 ( .A1(n6143), .A2(DATAI_0_), .ZN(n4568) );
  NAND2_X1 U5710 ( .A1(n4564), .A2(n4568), .ZN(U2924) );
  AOI22_X1 U5711 ( .A1(n6153), .A2(UWORD_REG_14__SCAN_IN), .B1(
        EAX_REG_30__SCAN_IN), .B2(n4572), .ZN(n4566) );
  NAND2_X1 U5712 ( .A1(n4566), .A2(n4565), .ZN(U2938) );
  AOI22_X1 U5713 ( .A1(n6153), .A2(LWORD_REG_1__SCAN_IN), .B1(
        EAX_REG_1__SCAN_IN), .B2(n4572), .ZN(n4567) );
  NAND2_X1 U5714 ( .A1(n6143), .A2(DATAI_1_), .ZN(n4573) );
  NAND2_X1 U5715 ( .A1(n4567), .A2(n4573), .ZN(U2940) );
  AOI22_X1 U5716 ( .A1(n6153), .A2(LWORD_REG_0__SCAN_IN), .B1(
        EAX_REG_0__SCAN_IN), .B2(n4572), .ZN(n4569) );
  NAND2_X1 U5717 ( .A1(n4569), .A2(n4568), .ZN(U2939) );
  AOI22_X1 U5718 ( .A1(n6153), .A2(LWORD_REG_2__SCAN_IN), .B1(
        EAX_REG_2__SCAN_IN), .B2(n4572), .ZN(n4571) );
  NAND2_X1 U5719 ( .A1(n4571), .A2(n4570), .ZN(U2941) );
  AOI22_X1 U5720 ( .A1(n6153), .A2(UWORD_REG_1__SCAN_IN), .B1(
        EAX_REG_17__SCAN_IN), .B2(n4572), .ZN(n4574) );
  NAND2_X1 U5721 ( .A1(n4574), .A2(n4573), .ZN(U2925) );
  OAI21_X1 U5722 ( .B1(n4577), .B2(n4576), .A(n4717), .ZN(n6256) );
  INV_X1 U5723 ( .A(EBX_REG_4__SCAN_IN), .ZN(n6581) );
  OAI222_X1 U5724 ( .A1(n6256), .A2(n6091), .B1(n6096), .B2(n6581), .C1(n6092), 
        .C2(n6046), .ZN(U2855) );
  INV_X1 U5725 ( .A(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4583) );
  INV_X1 U5726 ( .A(n6330), .ZN(n6319) );
  NAND2_X1 U5727 ( .A1(n6327), .A2(n6385), .ZN(n4579) );
  NAND2_X1 U5728 ( .A1(n5124), .A2(n6326), .ZN(n4578) );
  OAI211_X1 U5729 ( .C1(n5183), .C2(n4580), .A(n4579), .B(n4578), .ZN(n4581)
         );
  AOI21_X1 U5730 ( .B1(n6319), .B2(n4794), .A(n4581), .ZN(n4582) );
  OAI21_X1 U5731 ( .B1(n6395), .B2(n4583), .A(n4582), .ZN(U3142) );
  NAND2_X1 U5732 ( .A1(n5783), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5787) );
  NAND2_X1 U5733 ( .A1(n5787), .A2(n5797), .ZN(n4635) );
  INV_X1 U5734 ( .A(n4635), .ZN(n5782) );
  AOI21_X1 U5735 ( .B1(n5797), .B2(n4655), .A(n5782), .ZN(n4585) );
  OR2_X1 U5736 ( .A1(n4765), .A2(n4623), .ZN(n4896) );
  OR2_X1 U5737 ( .A1(n4896), .A2(n5254), .ZN(n4584) );
  AND2_X1 U5738 ( .A1(n4584), .A2(n6324), .ZN(n4586) );
  OAI22_X1 U5739 ( .A1(n4585), .A2(n4586), .B1(n4898), .B2(n6661), .ZN(n6337)
         );
  INV_X1 U5740 ( .A(n6337), .ZN(n4602) );
  INV_X1 U5741 ( .A(n4585), .ZN(n4587) );
  AOI22_X1 U5742 ( .A1(n4587), .A2(n4586), .B1(n4898), .B2(n5791), .ZN(n4588)
         );
  NAND2_X1 U5743 ( .A1(n4833), .A2(n4588), .ZN(n6338) );
  NAND2_X1 U5744 ( .A1(n6338), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4592) );
  NAND2_X1 U5745 ( .A1(n4589), .A2(n4744), .ZN(n6341) );
  NAND2_X1 U5746 ( .A1(n5783), .A2(n4808), .ZN(n4746) );
  OR2_X1 U5747 ( .A1(n4655), .A2(n4746), .ZN(n4858) );
  OAI22_X1 U5748 ( .A1(n4858), .A2(n5144), .B1(n5143), .B2(n6324), .ZN(n4590)
         );
  AOI21_X1 U5749 ( .B1(n5146), .B2(n4917), .A(n4590), .ZN(n4591) );
  OAI211_X1 U5750 ( .C1(n4602), .C2(n5824), .A(n4592), .B(n4591), .ZN(U3080)
         );
  NAND2_X1 U5751 ( .A1(n6338), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n4595) );
  OAI22_X1 U5752 ( .A1(n4858), .A2(n6379), .B1(n5173), .B2(n6324), .ZN(n4593)
         );
  AOI21_X1 U5753 ( .B1(n6310), .B2(n4917), .A(n4593), .ZN(n4594) );
  OAI211_X1 U5754 ( .C1(n4602), .C2(n5807), .A(n4595), .B(n4594), .ZN(U3076)
         );
  NAND2_X1 U5755 ( .A1(n6338), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4598) );
  OAI22_X1 U5756 ( .A1(n4858), .A2(n5168), .B1(n5167), .B2(n6324), .ZN(n4596)
         );
  AOI21_X1 U5757 ( .B1(n5170), .B2(n4917), .A(n4596), .ZN(n4597) );
  OAI211_X1 U5758 ( .C1(n4602), .C2(n5839), .A(n4598), .B(n4597), .ZN(U3083)
         );
  NAND2_X1 U5759 ( .A1(n6338), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n4601) );
  INV_X1 U5760 ( .A(n6387), .ZN(n6313) );
  OAI22_X1 U5761 ( .A1(n4858), .A2(n6390), .B1(n5177), .B2(n6324), .ZN(n4599)
         );
  AOI21_X1 U5762 ( .B1(n6313), .B2(n4917), .A(n4599), .ZN(n4600) );
  OAI211_X1 U5763 ( .C1(n4602), .C2(n5812), .A(n4601), .B(n4600), .ZN(U3077)
         );
  NAND2_X1 U5764 ( .A1(n6647), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4626) );
  INV_X1 U5765 ( .A(n4626), .ZN(n4619) );
  MUX2_X1 U5766 ( .A(n3180), .B(n4603), .S(n4622), .Z(n6411) );
  INV_X1 U5767 ( .A(n4604), .ZN(n4606) );
  MUX2_X1 U5768 ( .A(n4610), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(n2986), 
        .Z(n4605) );
  NOR3_X1 U5769 ( .A1(n4606), .A2(n4620), .A3(n4605), .ZN(n4616) );
  NAND2_X1 U5770 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n4607), .ZN(n4609) );
  INV_X1 U5771 ( .A(n4609), .ZN(n4608) );
  MUX2_X1 U5772 ( .A(n4609), .B(n4608), .S(INSTQUEUERD_ADDR_REG_3__SCAN_IN), 
        .Z(n4613) );
  INV_X1 U5773 ( .A(n4610), .ZN(n4611) );
  OAI211_X1 U5774 ( .C1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .C2(n2986), .A(n3261), .B(n4611), .ZN(n6532) );
  OAI22_X1 U5775 ( .A1(n4614), .A2(n4613), .B1(n4612), .B2(n6532), .ZN(n4615)
         );
  AOI211_X1 U5776 ( .C1(n6059), .C2(n6402), .A(n4616), .B(n4615), .ZN(n6534)
         );
  MUX2_X1 U5777 ( .A(n4617), .B(n6534), .S(n4622), .Z(n6416) );
  NOR3_X1 U5778 ( .A1(n6411), .A2(n6416), .A3(STATE2_REG_1__SCAN_IN), .ZN(
        n4618) );
  AOI21_X1 U5779 ( .B1(n4620), .B2(n4619), .A(n4618), .ZN(n6423) );
  NOR2_X1 U5780 ( .A1(n6423), .A2(n4621), .ZN(n4631) );
  INV_X1 U5781 ( .A(n4622), .ZN(n6407) );
  INV_X1 U5782 ( .A(n4623), .ZN(n4927) );
  NOR2_X1 U5783 ( .A1(n4624), .A2(n4927), .ZN(n4625) );
  XNOR2_X1 U5784 ( .A(n4625), .B(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n6049)
         );
  INV_X1 U5785 ( .A(n6049), .ZN(n5962) );
  AOI22_X1 U5786 ( .A1(n6407), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B1(n5960), .B2(n5962), .ZN(n4627) );
  INV_X1 U5787 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n5963) );
  OAI22_X1 U5788 ( .A1(n4627), .A2(STATE2_REG_1__SCAN_IN), .B1(n4626), .B2(
        n5963), .ZN(n6399) );
  NOR3_X1 U5789 ( .A1(n4631), .A2(n6399), .A3(FLUSH_REG_SCAN_IN), .ZN(n4628)
         );
  OAI21_X1 U5790 ( .B1(n4628), .B2(n6529), .A(n4991), .ZN(n6291) );
  INV_X1 U5791 ( .A(n4629), .ZN(n4630) );
  OR3_X1 U5792 ( .A1(n4631), .A2(n6399), .A3(n4630), .ZN(n6442) );
  INV_X1 U5793 ( .A(n6442), .ZN(n4633) );
  AND2_X1 U5794 ( .A1(n6717), .A2(STATE2_REG_1__SCAN_IN), .ZN(n5789) );
  OAI22_X1 U5795 ( .A1(n4837), .A2(n5791), .B1(n5254), .B2(n5789), .ZN(n4632)
         );
  OAI21_X1 U5796 ( .B1(n4633), .B2(n4632), .A(n6291), .ZN(n4634) );
  OAI21_X1 U5797 ( .B1(n6291), .B2(n4929), .A(n4634), .ZN(U3465) );
  OR2_X1 U5798 ( .A1(n4803), .A2(n5791), .ZN(n4636) );
  NAND2_X1 U5799 ( .A1(n4636), .A2(n4635), .ZN(n4645) );
  OR2_X1 U5800 ( .A1(n5208), .A2(n5785), .ZN(n4736) );
  INV_X1 U5801 ( .A(n4736), .ZN(n4637) );
  NAND2_X1 U5802 ( .A1(n4637), .A2(n6059), .ZN(n5131) );
  OR2_X1 U5803 ( .A1(n5131), .A2(n5254), .ZN(n4639) );
  INV_X1 U5804 ( .A(n4737), .ZN(n4638) );
  NAND2_X1 U5805 ( .A1(n4638), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6342) );
  NAND2_X1 U5806 ( .A1(n4639), .A2(n6342), .ZN(n4643) );
  NAND2_X1 U5807 ( .A1(n4645), .A2(n4643), .ZN(n4642) );
  NAND3_X1 U5808 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n4830), .ZN(n5135) );
  INV_X1 U5809 ( .A(n5135), .ZN(n4640) );
  NAND2_X1 U5810 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n4640), .ZN(n4641) );
  NAND2_X1 U5811 ( .A1(n4642), .A2(n4641), .ZN(n6368) );
  INV_X1 U5812 ( .A(n6368), .ZN(n4688) );
  INV_X1 U5813 ( .A(n4643), .ZN(n4644) );
  AOI22_X1 U5814 ( .A1(n4645), .A2(n4644), .B1(n5135), .B2(n5791), .ZN(n4646)
         );
  NAND2_X1 U5815 ( .A1(n4833), .A2(n4646), .ZN(n6370) );
  NAND2_X1 U5816 ( .A1(n6370), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n4651)
         );
  INV_X1 U5817 ( .A(n4746), .ZN(n4647) );
  NAND2_X1 U5818 ( .A1(n4803), .A2(n4647), .ZN(n4962) );
  OAI22_X1 U5819 ( .A1(n4962), .A2(n6379), .B1(n5173), .B2(n6342), .ZN(n4649)
         );
  INV_X1 U5820 ( .A(n6310), .ZN(n6377) );
  NOR2_X1 U5821 ( .A1(n6373), .A2(n6377), .ZN(n4648) );
  NOR2_X1 U5822 ( .A1(n4649), .A2(n4648), .ZN(n4650) );
  OAI211_X1 U5823 ( .C1(n4688), .C2(n5807), .A(n4651), .B(n4650), .ZN(U3108)
         );
  INV_X1 U5824 ( .A(n6291), .ZN(n4660) );
  INV_X1 U5825 ( .A(n4803), .ZN(n4654) );
  NOR2_X1 U5826 ( .A1(n5783), .A2(n4652), .ZN(n4653) );
  NAND2_X1 U5827 ( .A1(n4732), .A2(n4653), .ZN(n4677) );
  OR2_X1 U5828 ( .A1(n4677), .A2(n5973), .ZN(n4673) );
  AND2_X1 U5829 ( .A1(n4654), .A2(n4673), .ZN(n4734) );
  OAI21_X1 U5830 ( .B1(n4655), .B2(n5787), .A(n4734), .ZN(n4657) );
  INV_X1 U5831 ( .A(n6059), .ZN(n4996) );
  OAI22_X1 U5832 ( .A1(n4743), .A2(n5800), .B1(n4996), .B2(n5789), .ZN(n4656)
         );
  AOI21_X1 U5833 ( .B1(n4657), .B2(n5089), .A(n4656), .ZN(n4659) );
  NAND2_X1 U5834 ( .A1(n4660), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4658) );
  OAI21_X1 U5835 ( .B1(n4660), .B2(n4659), .A(n4658), .ZN(U3462) );
  NAND2_X1 U5836 ( .A1(n4663), .A2(n4664), .ZN(n4665) );
  NAND2_X1 U5837 ( .A1(n4923), .A2(n4665), .ZN(n5623) );
  CLKBUF_X1 U5838 ( .A(n4666), .Z(n5432) );
  INV_X1 U5839 ( .A(n5049), .ZN(n4667) );
  AOI21_X1 U5840 ( .B1(n4668), .B2(n5432), .A(n4667), .ZN(n5954) );
  AOI22_X1 U5841 ( .A1(n5954), .A2(n6087), .B1(n5462), .B2(EBX_REG_13__SCAN_IN), .ZN(n4669) );
  OAI21_X1 U5842 ( .B1(n5623), .B2(n6092), .A(n4669), .ZN(U2846) );
  INV_X1 U5843 ( .A(n4677), .ZN(n4670) );
  NOR3_X1 U5844 ( .A1(n4830), .A2(n6419), .A3(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .ZN(n4928) );
  INV_X1 U5845 ( .A(n4933), .ZN(n4671) );
  INV_X1 U5846 ( .A(n4928), .ZN(n4674) );
  NOR2_X1 U5847 ( .A1(n4929), .A2(n4674), .ZN(n4701) );
  AOI21_X1 U5848 ( .B1(n4801), .B2(n4671), .A(n4701), .ZN(n4676) );
  NAND3_X1 U5849 ( .A1(n5797), .A2(n4676), .A3(n4673), .ZN(n4672) );
  OAI211_X1 U5850 ( .C1(n5797), .C2(n4928), .A(n4833), .B(n4672), .ZN(n4700)
         );
  NAND2_X1 U5851 ( .A1(n5797), .A2(n4673), .ZN(n4675) );
  OAI22_X1 U5852 ( .A1(n4676), .A2(n4675), .B1(n6661), .B2(n4674), .ZN(n4699)
         );
  AOI22_X1 U5853 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n4700), .B1(n6298), 
        .B2(n4699), .ZN(n4679) );
  NOR2_X2 U5854 ( .A1(n4677), .A2(n4808), .ZN(n4959) );
  AOI22_X1 U5855 ( .A1(n4959), .A2(n5146), .B1(n6296), .B2(n4701), .ZN(n4678)
         );
  OAI211_X1 U5856 ( .C1(n5144), .C2(n4797), .A(n4679), .B(n4678), .ZN(U3128)
         );
  AOI22_X1 U5857 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(n4700), .B1(n6376), 
        .B2(n4699), .ZN(n4681) );
  INV_X1 U5858 ( .A(n5173), .ZN(n6375) );
  AOI22_X1 U5859 ( .A1(n4959), .A2(n6310), .B1(n6375), .B2(n4701), .ZN(n4680)
         );
  OAI211_X1 U5860 ( .C1(n6379), .C2(n4797), .A(n4681), .B(n4680), .ZN(U3124)
         );
  NAND2_X1 U5861 ( .A1(n6370), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n4684)
         );
  OAI22_X1 U5862 ( .A1(n4962), .A2(n6323), .B1(n5183), .B2(n6342), .ZN(n4682)
         );
  AOI21_X1 U5863 ( .B1(n6319), .B2(n5129), .A(n4682), .ZN(n4683) );
  OAI211_X1 U5864 ( .C1(n4688), .C2(n5816), .A(n4684), .B(n4683), .ZN(U3110)
         );
  NAND2_X1 U5865 ( .A1(n6370), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n4687)
         );
  OAI22_X1 U5866 ( .A1(n4962), .A2(n5144), .B1(n5143), .B2(n6342), .ZN(n4685)
         );
  AOI21_X1 U5867 ( .B1(n5146), .B2(n5129), .A(n4685), .ZN(n4686) );
  OAI211_X1 U5868 ( .C1(n4688), .C2(n5824), .A(n4687), .B(n4686), .ZN(U3112)
         );
  AOI22_X1 U5869 ( .A1(INSTQUEUE_REG_13__7__SCAN_IN), .A2(n4700), .B1(n6369), 
        .B2(n4699), .ZN(n4690) );
  AOI22_X1 U5870 ( .A1(n4959), .A2(n5170), .B1(n6365), .B2(n4701), .ZN(n4689)
         );
  OAI211_X1 U5871 ( .C1(n5168), .C2(n4797), .A(n4690), .B(n4689), .ZN(U3131)
         );
  AOI22_X1 U5872 ( .A1(INSTQUEUE_REG_13__6__SCAN_IN), .A2(n4700), .B1(n6360), 
        .B2(n4699), .ZN(n4692) );
  AOI22_X1 U5873 ( .A1(n4959), .A2(n5164), .B1(n6358), .B2(n4701), .ZN(n4691)
         );
  OAI211_X1 U5874 ( .C1(n5162), .C2(n4797), .A(n4692), .B(n4691), .ZN(U3130)
         );
  AOI22_X1 U5875 ( .A1(INSTQUEUE_REG_13__5__SCAN_IN), .A2(n4700), .B1(n6354), 
        .B2(n4699), .ZN(n4694) );
  AOI22_X1 U5876 ( .A1(n4959), .A2(n5158), .B1(n6352), .B2(n4701), .ZN(n4693)
         );
  OAI211_X1 U5877 ( .C1(n5156), .C2(n4797), .A(n4694), .B(n4693), .ZN(U3129)
         );
  AOI22_X1 U5878 ( .A1(INSTQUEUE_REG_13__1__SCAN_IN), .A2(n4700), .B1(n6386), 
        .B2(n4699), .ZN(n4696) );
  INV_X1 U5879 ( .A(n5177), .ZN(n6383) );
  AOI22_X1 U5880 ( .A1(n4959), .A2(n6313), .B1(n6383), .B2(n4701), .ZN(n4695)
         );
  OAI211_X1 U5881 ( .C1(n6390), .C2(n4797), .A(n4696), .B(n4695), .ZN(U3125)
         );
  AOI22_X1 U5882 ( .A1(INSTQUEUE_REG_13__3__SCAN_IN), .A2(n4700), .B1(n6348), 
        .B2(n4699), .ZN(n4698) );
  AOI22_X1 U5883 ( .A1(n4959), .A2(n5152), .B1(n6346), .B2(n4701), .ZN(n4697)
         );
  OAI211_X1 U5884 ( .C1(n5150), .C2(n4797), .A(n4698), .B(n4697), .ZN(U3127)
         );
  AOI22_X1 U5885 ( .A1(INSTQUEUE_REG_13__2__SCAN_IN), .A2(n4700), .B1(n6327), 
        .B2(n4699), .ZN(n4703) );
  INV_X1 U5886 ( .A(n5183), .ZN(n6325) );
  AOI22_X1 U5887 ( .A1(n4959), .A2(n6319), .B1(n6325), .B2(n4701), .ZN(n4702)
         );
  OAI211_X1 U5888 ( .C1(n6323), .C2(n4797), .A(n4703), .B(n4702), .ZN(U3126)
         );
  INV_X1 U5889 ( .A(EAX_REG_13__SCAN_IN), .ZN(n6725) );
  OAI222_X1 U5890 ( .A1(n5623), .A2(n5914), .B1(n5203), .B2(n4704), .C1(n5472), 
        .C2(n6725), .ZN(U2878) );
  OAI21_X1 U5891 ( .B1(n4707), .B2(n4706), .A(n4705), .ZN(n4972) );
  INV_X1 U5892 ( .A(n6206), .ZN(n4710) );
  OAI22_X1 U5893 ( .A1(n4710), .A2(n4709), .B1(n5771), .B2(n4708), .ZN(n6281)
         );
  AOI21_X1 U5894 ( .B1(n4711), .B2(n6210), .A(n6281), .ZN(n6253) );
  INV_X1 U5895 ( .A(n6253), .ZN(n4722) );
  OAI21_X1 U5896 ( .B1(n6276), .B2(n4712), .A(n4713), .ZN(n4721) );
  NAND2_X1 U5897 ( .A1(n4714), .A2(n4713), .ZN(n4715) );
  NOR2_X1 U5898 ( .A1(n6284), .A2(n4715), .ZN(n4720) );
  NAND2_X1 U5899 ( .A1(n4717), .A2(n4716), .ZN(n4718) );
  AND2_X1 U5900 ( .A1(n5195), .A2(n4718), .ZN(n5266) );
  INV_X1 U5901 ( .A(n5266), .ZN(n4974) );
  OAI22_X1 U5902 ( .A1(n6249), .A2(n4974), .B1(n6724), .B2(n6248), .ZN(n4719)
         );
  AOI211_X1 U5903 ( .C1(n4722), .C2(n4721), .A(n4720), .B(n4719), .ZN(n4723)
         );
  OAI21_X1 U5904 ( .B1(n5780), .B2(n4972), .A(n4723), .ZN(U3013) );
  OAI21_X1 U5905 ( .B1(n4726), .B2(n4725), .A(n4724), .ZN(n6267) );
  INV_X1 U5906 ( .A(n4727), .ZN(n6058) );
  NAND2_X1 U5907 ( .A1(n3668), .A2(REIP_REG_3__SCAN_IN), .ZN(n6264) );
  OAI21_X1 U5908 ( .B1(n5618), .B2(n4728), .A(n6264), .ZN(n4730) );
  NOR2_X1 U5909 ( .A1(n6057), .A2(n5634), .ZN(n4729) );
  AOI211_X1 U5910 ( .C1(n6164), .C2(n6058), .A(n4730), .B(n4729), .ZN(n4731)
         );
  OAI21_X1 U5911 ( .B1(n6169), .B2(n6267), .A(n4731), .ZN(U2983) );
  INV_X1 U5912 ( .A(n5787), .ZN(n4733) );
  NAND3_X1 U5913 ( .A1(n4734), .A2(n4733), .A3(n5788), .ZN(n4735) );
  NAND2_X1 U5914 ( .A1(n4735), .A2(n5797), .ZN(n4742) );
  NOR2_X1 U5915 ( .A1(n6059), .A2(n4736), .ZN(n5799) );
  NOR2_X1 U5916 ( .A1(n4737), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6302)
         );
  AOI21_X1 U5917 ( .B1(n5799), .B2(n6403), .A(n6302), .ZN(n4738) );
  NAND3_X1 U5918 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n6419), .A3(n4830), .ZN(n5798) );
  OAI22_X1 U5919 ( .A1(n4742), .A2(n4738), .B1(n5798), .B2(n6661), .ZN(n6304)
         );
  INV_X1 U5920 ( .A(n6304), .ZN(n4759) );
  INV_X1 U5921 ( .A(n4738), .ZN(n4741) );
  AOI21_X1 U5922 ( .B1(n5798), .B2(n5791), .A(n4739), .ZN(n4740) );
  OAI21_X1 U5923 ( .B1(n4742), .B2(n4741), .A(n4740), .ZN(n6305) );
  NAND2_X1 U5924 ( .A1(n5788), .A2(n4743), .ZN(n4829) );
  INV_X1 U5925 ( .A(n4829), .ZN(n4745) );
  NOR2_X2 U5926 ( .A1(n4829), .A2(n4746), .ZN(n6303) );
  AOI22_X1 U5927 ( .A1(n6303), .A2(n6359), .B1(n6358), .B2(n6302), .ZN(n4747)
         );
  OAI21_X1 U5928 ( .B1(n6363), .B2(n6308), .A(n4747), .ZN(n4748) );
  AOI21_X1 U5929 ( .B1(n6305), .B2(INSTQUEUE_REG_3__6__SCAN_IN), .A(n4748), 
        .ZN(n4749) );
  OAI21_X1 U5930 ( .B1(n4759), .B2(n5832), .A(n4749), .ZN(U3050) );
  INV_X1 U5931 ( .A(n6379), .ZN(n5809) );
  AOI22_X1 U5932 ( .A1(n6303), .A2(n5809), .B1(n6375), .B2(n6302), .ZN(n4750)
         );
  OAI21_X1 U5933 ( .B1(n6377), .B2(n6308), .A(n4750), .ZN(n4751) );
  AOI21_X1 U5934 ( .B1(n6305), .B2(INSTQUEUE_REG_3__0__SCAN_IN), .A(n4751), 
        .ZN(n4752) );
  OAI21_X1 U5935 ( .B1(n4759), .B2(n5807), .A(n4752), .ZN(U3044) );
  AOI22_X1 U5936 ( .A1(n6303), .A2(n6353), .B1(n6352), .B2(n6302), .ZN(n4753)
         );
  OAI21_X1 U5937 ( .B1(n6357), .B2(n6308), .A(n4753), .ZN(n4754) );
  AOI21_X1 U5938 ( .B1(n6305), .B2(INSTQUEUE_REG_3__5__SCAN_IN), .A(n4754), 
        .ZN(n4755) );
  OAI21_X1 U5939 ( .B1(n4759), .B2(n5828), .A(n4755), .ZN(U3049) );
  AOI22_X1 U5940 ( .A1(n6303), .A2(n6343), .B1(n6383), .B2(n6302), .ZN(n4756)
         );
  OAI21_X1 U5941 ( .B1(n6387), .B2(n6308), .A(n4756), .ZN(n4757) );
  AOI21_X1 U5942 ( .B1(n6305), .B2(INSTQUEUE_REG_3__1__SCAN_IN), .A(n4757), 
        .ZN(n4758) );
  OAI21_X1 U5943 ( .B1(n4759), .B2(n5812), .A(n4758), .ZN(U3045) );
  NOR2_X1 U5944 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4760), .ZN(n4768)
         );
  INV_X1 U5945 ( .A(n4991), .ZN(n4864) );
  OAI21_X1 U5946 ( .B1(n5796), .B2(n6661), .A(n4864), .ZN(n5137) );
  NOR2_X1 U5947 ( .A1(n4766), .A2(n6661), .ZN(n5132) );
  NOR3_X1 U5948 ( .A1(n5137), .A2(n6419), .A3(n5132), .ZN(n4764) );
  INV_X1 U5949 ( .A(n4797), .ZN(n4761) );
  OAI21_X1 U5950 ( .B1(n4761), .B2(n4794), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n4762) );
  NAND3_X1 U5951 ( .A1(n4765), .A2(n5797), .A3(n4762), .ZN(n4763) );
  OAI211_X1 U5952 ( .C1(n4768), .C2(n6717), .A(n4764), .B(n4763), .ZN(n4790)
         );
  NAND2_X1 U5953 ( .A1(n4790), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4771)
         );
  NOR2_X1 U5954 ( .A1(n4765), .A2(n5791), .ZN(n4902) );
  AND2_X1 U5955 ( .A1(n4766), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5138) );
  INV_X1 U5956 ( .A(n5138), .ZN(n5093) );
  NOR2_X1 U5957 ( .A1(n5093), .A2(n6419), .ZN(n4767) );
  AOI22_X1 U5958 ( .A1(n4902), .A2(n6059), .B1(n5796), .B2(n4767), .ZN(n4792)
         );
  INV_X1 U5959 ( .A(n4768), .ZN(n4791) );
  OAI22_X1 U5960 ( .A1(n5828), .A2(n4792), .B1(n5155), .B2(n4791), .ZN(n4769)
         );
  AOI21_X1 U5961 ( .B1(n6353), .B2(n4794), .A(n4769), .ZN(n4770) );
  OAI211_X1 U5962 ( .C1(n4797), .C2(n6357), .A(n4771), .B(n4770), .ZN(U3137)
         );
  NAND2_X1 U5963 ( .A1(n4790), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n4774)
         );
  OAI22_X1 U5964 ( .A1(n5812), .A2(n4792), .B1(n5177), .B2(n4791), .ZN(n4772)
         );
  AOI21_X1 U5965 ( .B1(n6343), .B2(n4794), .A(n4772), .ZN(n4773) );
  OAI211_X1 U5966 ( .C1(n4797), .C2(n6387), .A(n4774), .B(n4773), .ZN(U3133)
         );
  NAND2_X1 U5967 ( .A1(n4790), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4777)
         );
  OAI22_X1 U5968 ( .A1(n5824), .A2(n4792), .B1(n5143), .B2(n4791), .ZN(n4775)
         );
  AOI21_X1 U5969 ( .B1(n6297), .B2(n4794), .A(n4775), .ZN(n4776) );
  OAI211_X1 U5970 ( .C1(n4797), .C2(n6301), .A(n4777), .B(n4776), .ZN(U3136)
         );
  NAND2_X1 U5971 ( .A1(n4790), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4780)
         );
  OAI22_X1 U5972 ( .A1(n5807), .A2(n4792), .B1(n5173), .B2(n4791), .ZN(n4778)
         );
  AOI21_X1 U5973 ( .B1(n5809), .B2(n4794), .A(n4778), .ZN(n4779) );
  OAI211_X1 U5974 ( .C1(n4797), .C2(n6377), .A(n4780), .B(n4779), .ZN(U3132)
         );
  NAND2_X1 U5975 ( .A1(n4790), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4783)
         );
  OAI22_X1 U5976 ( .A1(n5839), .A2(n4792), .B1(n5167), .B2(n4791), .ZN(n4781)
         );
  AOI21_X1 U5977 ( .B1(n6366), .B2(n4794), .A(n4781), .ZN(n4782) );
  OAI211_X1 U5978 ( .C1(n4797), .C2(n6374), .A(n4783), .B(n4782), .ZN(U3139)
         );
  NAND2_X1 U5979 ( .A1(n4790), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4786)
         );
  OAI22_X1 U5980 ( .A1(n5816), .A2(n4792), .B1(n5183), .B2(n4791), .ZN(n4784)
         );
  AOI21_X1 U5981 ( .B1(n6326), .B2(n4794), .A(n4784), .ZN(n4785) );
  OAI211_X1 U5982 ( .C1(n4797), .C2(n6330), .A(n4786), .B(n4785), .ZN(U3134)
         );
  NAND2_X1 U5983 ( .A1(n4790), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4789)
         );
  OAI22_X1 U5984 ( .A1(n5820), .A2(n4792), .B1(n5149), .B2(n4791), .ZN(n4787)
         );
  AOI21_X1 U5985 ( .B1(n6347), .B2(n4794), .A(n4787), .ZN(n4788) );
  OAI211_X1 U5986 ( .C1(n4797), .C2(n6351), .A(n4789), .B(n4788), .ZN(U3135)
         );
  NAND2_X1 U5987 ( .A1(n4790), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4796)
         );
  OAI22_X1 U5988 ( .A1(n5832), .A2(n4792), .B1(n5161), .B2(n4791), .ZN(n4793)
         );
  AOI21_X1 U5989 ( .B1(n6359), .B2(n4794), .A(n4793), .ZN(n4795) );
  OAI211_X1 U5990 ( .C1(n4797), .C2(n6363), .A(n4796), .B(n4795), .ZN(U3138)
         );
  INV_X1 U5991 ( .A(n5783), .ZN(n4798) );
  NAND2_X1 U5992 ( .A1(n4803), .A2(n4798), .ZN(n4809) );
  INV_X1 U5993 ( .A(n4809), .ZN(n4799) );
  OR2_X1 U5994 ( .A1(n5208), .A2(n6070), .ZN(n4862) );
  INV_X1 U5995 ( .A(n4862), .ZN(n4800) );
  NAND3_X1 U5996 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n4830), .A3(n6612), .ZN(n4863) );
  NOR2_X1 U5997 ( .A1(n4929), .A2(n4863), .ZN(n4826) );
  AOI21_X1 U5998 ( .B1(n4801), .B2(n4800), .A(n4826), .ZN(n4807) );
  AOI21_X1 U5999 ( .B1(n4803), .B2(n4802), .A(n5791), .ZN(n4805) );
  AOI22_X1 U6000 ( .A1(n4807), .A2(n4805), .B1(n5791), .B2(n4863), .ZN(n4804)
         );
  NAND2_X1 U6001 ( .A1(n4833), .A2(n4804), .ZN(n4825) );
  INV_X1 U6002 ( .A(n4805), .ZN(n4806) );
  OAI22_X1 U6003 ( .A1(n4807), .A2(n4806), .B1(n6661), .B2(n4863), .ZN(n4824)
         );
  AOI22_X1 U6004 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n4825), .B1(n6298), 
        .B2(n4824), .ZN(n4811) );
  AOI22_X1 U6005 ( .A1(n4859), .A2(n5146), .B1(n6296), .B2(n4826), .ZN(n4810)
         );
  OAI211_X1 U6006 ( .C1(n5144), .C2(n5128), .A(n4811), .B(n4810), .ZN(U3096)
         );
  AOI22_X1 U6007 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n4825), .B1(n6376), 
        .B2(n4824), .ZN(n4813) );
  AOI22_X1 U6008 ( .A1(n4859), .A2(n6310), .B1(n6375), .B2(n4826), .ZN(n4812)
         );
  OAI211_X1 U6009 ( .C1(n6379), .C2(n5128), .A(n4813), .B(n4812), .ZN(U3092)
         );
  AOI22_X1 U6010 ( .A1(INSTQUEUE_REG_9__6__SCAN_IN), .A2(n4825), .B1(n6360), 
        .B2(n4824), .ZN(n4815) );
  AOI22_X1 U6011 ( .A1(n4859), .A2(n5164), .B1(n6358), .B2(n4826), .ZN(n4814)
         );
  OAI211_X1 U6012 ( .C1(n5162), .C2(n5128), .A(n4815), .B(n4814), .ZN(U3098)
         );
  AOI22_X1 U6013 ( .A1(INSTQUEUE_REG_9__7__SCAN_IN), .A2(n4825), .B1(n6369), 
        .B2(n4824), .ZN(n4817) );
  AOI22_X1 U6014 ( .A1(n4859), .A2(n5170), .B1(n6365), .B2(n4826), .ZN(n4816)
         );
  OAI211_X1 U6015 ( .C1(n5168), .C2(n5128), .A(n4817), .B(n4816), .ZN(U3099)
         );
  AOI22_X1 U6016 ( .A1(INSTQUEUE_REG_9__5__SCAN_IN), .A2(n4825), .B1(n6354), 
        .B2(n4824), .ZN(n4819) );
  AOI22_X1 U6017 ( .A1(n4859), .A2(n5158), .B1(n6352), .B2(n4826), .ZN(n4818)
         );
  OAI211_X1 U6018 ( .C1(n5156), .C2(n5128), .A(n4819), .B(n4818), .ZN(U3097)
         );
  AOI22_X1 U6019 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(n4825), .B1(n6386), 
        .B2(n4824), .ZN(n4821) );
  AOI22_X1 U6020 ( .A1(n4859), .A2(n6313), .B1(n6383), .B2(n4826), .ZN(n4820)
         );
  OAI211_X1 U6021 ( .C1(n6390), .C2(n5128), .A(n4821), .B(n4820), .ZN(U3093)
         );
  AOI22_X1 U6022 ( .A1(INSTQUEUE_REG_9__3__SCAN_IN), .A2(n4825), .B1(n6348), 
        .B2(n4824), .ZN(n4823) );
  AOI22_X1 U6023 ( .A1(n4859), .A2(n5152), .B1(n6346), .B2(n4826), .ZN(n4822)
         );
  OAI211_X1 U6024 ( .C1(n5150), .C2(n5128), .A(n4823), .B(n4822), .ZN(U3095)
         );
  AOI22_X1 U6025 ( .A1(INSTQUEUE_REG_9__2__SCAN_IN), .A2(n4825), .B1(n6327), 
        .B2(n4824), .ZN(n4828) );
  AOI22_X1 U6026 ( .A1(n4859), .A2(n6319), .B1(n6325), .B2(n4826), .ZN(n4827)
         );
  OAI211_X1 U6027 ( .C1(n6323), .C2(n5128), .A(n4828), .B(n4827), .ZN(U3094)
         );
  NOR2_X1 U6028 ( .A1(n6059), .A2(n4862), .ZN(n5097) );
  NAND3_X1 U6029 ( .A1(n6419), .A2(n4830), .A3(n6612), .ZN(n5091) );
  NOR2_X1 U6030 ( .A1(n4929), .A2(n5091), .ZN(n4855) );
  AOI21_X1 U6031 ( .B1(n5097), .B2(n6403), .A(n4855), .ZN(n4836) );
  AOI21_X1 U6032 ( .B1(n4831), .B2(STATEBS16_REG_SCAN_IN), .A(n5791), .ZN(
        n4834) );
  AOI22_X1 U6033 ( .A1(n4836), .A2(n4834), .B1(n5791), .B2(n5091), .ZN(n4832)
         );
  NAND2_X1 U6034 ( .A1(n4833), .A2(n4832), .ZN(n4854) );
  INV_X1 U6035 ( .A(n4834), .ZN(n4835) );
  OAI22_X1 U6036 ( .A1(n4836), .A2(n4835), .B1(n6661), .B2(n5091), .ZN(n4853)
         );
  AOI22_X1 U6037 ( .A1(INSTQUEUE_REG_1__6__SCAN_IN), .A2(n4854), .B1(n6360), 
        .B2(n4853), .ZN(n4840) );
  AOI22_X1 U6038 ( .A1(n5801), .A2(n6359), .B1(n6358), .B2(n4855), .ZN(n4839)
         );
  OAI211_X1 U6039 ( .C1(n6363), .C2(n5127), .A(n4840), .B(n4839), .ZN(U3034)
         );
  AOI22_X1 U6040 ( .A1(INSTQUEUE_REG_1__3__SCAN_IN), .A2(n4854), .B1(n6348), 
        .B2(n4853), .ZN(n4842) );
  AOI22_X1 U6041 ( .A1(n5801), .A2(n6347), .B1(n6346), .B2(n4855), .ZN(n4841)
         );
  OAI211_X1 U6042 ( .C1(n6351), .C2(n5127), .A(n4842), .B(n4841), .ZN(U3031)
         );
  AOI22_X1 U6043 ( .A1(INSTQUEUE_REG_1__7__SCAN_IN), .A2(n4854), .B1(n6369), 
        .B2(n4853), .ZN(n4844) );
  AOI22_X1 U6044 ( .A1(n5801), .A2(n6366), .B1(n6365), .B2(n4855), .ZN(n4843)
         );
  OAI211_X1 U6045 ( .C1(n6374), .C2(n5127), .A(n4844), .B(n4843), .ZN(U3035)
         );
  AOI22_X1 U6046 ( .A1(INSTQUEUE_REG_1__1__SCAN_IN), .A2(n4854), .B1(n6386), 
        .B2(n4853), .ZN(n4846) );
  AOI22_X1 U6047 ( .A1(n5801), .A2(n6343), .B1(n6383), .B2(n4855), .ZN(n4845)
         );
  OAI211_X1 U6048 ( .C1(n6387), .C2(n5127), .A(n4846), .B(n4845), .ZN(U3029)
         );
  AOI22_X1 U6049 ( .A1(INSTQUEUE_REG_1__4__SCAN_IN), .A2(n4854), .B1(n6298), 
        .B2(n4853), .ZN(n4848) );
  AOI22_X1 U6050 ( .A1(n5801), .A2(n6297), .B1(n6296), .B2(n4855), .ZN(n4847)
         );
  OAI211_X1 U6051 ( .C1(n6301), .C2(n5127), .A(n4848), .B(n4847), .ZN(U3032)
         );
  AOI22_X1 U6052 ( .A1(INSTQUEUE_REG_1__5__SCAN_IN), .A2(n4854), .B1(n6354), 
        .B2(n4853), .ZN(n4850) );
  AOI22_X1 U6053 ( .A1(n5801), .A2(n6353), .B1(n6352), .B2(n4855), .ZN(n4849)
         );
  OAI211_X1 U6054 ( .C1(n6357), .C2(n5127), .A(n4850), .B(n4849), .ZN(U3033)
         );
  AOI22_X1 U6055 ( .A1(INSTQUEUE_REG_1__0__SCAN_IN), .A2(n4854), .B1(n6376), 
        .B2(n4853), .ZN(n4852) );
  AOI22_X1 U6056 ( .A1(n5801), .A2(n5809), .B1(n6375), .B2(n4855), .ZN(n4851)
         );
  OAI211_X1 U6057 ( .C1(n6377), .C2(n5127), .A(n4852), .B(n4851), .ZN(U3028)
         );
  AOI22_X1 U6058 ( .A1(INSTQUEUE_REG_1__2__SCAN_IN), .A2(n4854), .B1(n6327), 
        .B2(n4853), .ZN(n4857) );
  AOI22_X1 U6059 ( .A1(n5801), .A2(n6326), .B1(n6325), .B2(n4855), .ZN(n4856)
         );
  OAI211_X1 U6060 ( .C1(n6330), .C2(n5127), .A(n4857), .B(n4856), .ZN(U3030)
         );
  NOR3_X1 U6061 ( .A1(n4859), .A2(n6336), .A3(n5791), .ZN(n4861) );
  INV_X1 U6062 ( .A(n5800), .ZN(n4860) );
  NOR2_X1 U6063 ( .A1(n4861), .A2(n4860), .ZN(n4866) );
  NOR2_X1 U6064 ( .A1(n4996), .A2(n4862), .ZN(n4867) );
  OR2_X1 U6065 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4863), .ZN(n4890)
         );
  OAI21_X1 U6066 ( .B1(n2977), .B2(n6661), .A(n4864), .ZN(n4930) );
  AOI211_X1 U6067 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n4890), .A(n5138), .B(
        n4930), .ZN(n4865) );
  OAI21_X1 U6068 ( .B1(n4866), .B2(n4867), .A(n4865), .ZN(n4889) );
  NAND2_X1 U6069 ( .A1(n4889), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n4870) );
  AOI22_X1 U6070 ( .A1(n4867), .A2(n5797), .B1(n5132), .B2(n2977), .ZN(n4891)
         );
  OAI22_X1 U6071 ( .A1(n5828), .A2(n4891), .B1(n5155), .B2(n4890), .ZN(n4868)
         );
  AOI21_X1 U6072 ( .B1(n5158), .B2(n6336), .A(n4868), .ZN(n4869) );
  OAI211_X1 U6073 ( .C1(n4895), .C2(n5156), .A(n4870), .B(n4869), .ZN(U3089)
         );
  NAND2_X1 U6074 ( .A1(n4889), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n4873) );
  OAI22_X1 U6075 ( .A1(n5807), .A2(n4891), .B1(n5173), .B2(n4890), .ZN(n4871)
         );
  AOI21_X1 U6076 ( .B1(n6310), .B2(n6336), .A(n4871), .ZN(n4872) );
  OAI211_X1 U6077 ( .C1(n4895), .C2(n6379), .A(n4873), .B(n4872), .ZN(U3084)
         );
  NAND2_X1 U6078 ( .A1(n4889), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n4876) );
  OAI22_X1 U6079 ( .A1(n5812), .A2(n4891), .B1(n5177), .B2(n4890), .ZN(n4874)
         );
  AOI21_X1 U6080 ( .B1(n6313), .B2(n6336), .A(n4874), .ZN(n4875) );
  OAI211_X1 U6081 ( .C1(n4895), .C2(n6390), .A(n4876), .B(n4875), .ZN(U3085)
         );
  NAND2_X1 U6082 ( .A1(n4889), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n4879) );
  OAI22_X1 U6083 ( .A1(n5816), .A2(n4891), .B1(n5183), .B2(n4890), .ZN(n4877)
         );
  AOI21_X1 U6084 ( .B1(n6319), .B2(n6336), .A(n4877), .ZN(n4878) );
  OAI211_X1 U6085 ( .C1(n4895), .C2(n6323), .A(n4879), .B(n4878), .ZN(U3086)
         );
  NAND2_X1 U6086 ( .A1(n4889), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n4882) );
  OAI22_X1 U6087 ( .A1(n5824), .A2(n4891), .B1(n5143), .B2(n4890), .ZN(n4880)
         );
  AOI21_X1 U6088 ( .B1(n5146), .B2(n6336), .A(n4880), .ZN(n4881) );
  OAI211_X1 U6089 ( .C1(n4895), .C2(n5144), .A(n4882), .B(n4881), .ZN(U3088)
         );
  NAND2_X1 U6090 ( .A1(n4889), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n4885) );
  OAI22_X1 U6091 ( .A1(n5832), .A2(n4891), .B1(n5161), .B2(n4890), .ZN(n4883)
         );
  AOI21_X1 U6092 ( .B1(n5164), .B2(n6336), .A(n4883), .ZN(n4884) );
  OAI211_X1 U6093 ( .C1(n4895), .C2(n5162), .A(n4885), .B(n4884), .ZN(U3090)
         );
  NAND2_X1 U6094 ( .A1(n4889), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n4888) );
  OAI22_X1 U6095 ( .A1(n5839), .A2(n4891), .B1(n5167), .B2(n4890), .ZN(n4886)
         );
  AOI21_X1 U6096 ( .B1(n5170), .B2(n6336), .A(n4886), .ZN(n4887) );
  OAI211_X1 U6097 ( .C1(n4895), .C2(n5168), .A(n4888), .B(n4887), .ZN(U3091)
         );
  NAND2_X1 U6098 ( .A1(n4889), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n4894) );
  OAI22_X1 U6099 ( .A1(n5820), .A2(n4891), .B1(n5149), .B2(n4890), .ZN(n4892)
         );
  AOI21_X1 U6100 ( .B1(n5152), .B2(n6336), .A(n4892), .ZN(n4893) );
  OAI211_X1 U6101 ( .C1(n4895), .C2(n5150), .A(n4894), .B(n4893), .ZN(U3087)
         );
  OAI21_X1 U6102 ( .B1(n6318), .B2(n4917), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n4897) );
  NAND3_X1 U6103 ( .A1(n4897), .A2(n5089), .A3(n4896), .ZN(n4900) );
  NOR2_X1 U6104 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4898), .ZN(n6316)
         );
  INV_X1 U6105 ( .A(n6316), .ZN(n4915) );
  AOI211_X1 U6106 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n4915), .A(n5132), .B(
        n5137), .ZN(n4899) );
  NAND3_X1 U6107 ( .A1(n4900), .A2(n4899), .A3(n6419), .ZN(n6320) );
  NAND2_X1 U6108 ( .A1(n6320), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n4905) );
  NOR2_X1 U6109 ( .A1(n5093), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4901)
         );
  AOI22_X1 U6110 ( .A1(n4902), .A2(n4996), .B1(n5796), .B2(n4901), .ZN(n6309)
         );
  OAI22_X1 U6111 ( .A1(n5824), .A2(n6309), .B1(n5143), .B2(n4915), .ZN(n4903)
         );
  AOI21_X1 U6112 ( .B1(n6297), .B2(n4917), .A(n4903), .ZN(n4904) );
  OAI211_X1 U6113 ( .C1(n4920), .C2(n6301), .A(n4905), .B(n4904), .ZN(U3072)
         );
  NAND2_X1 U6114 ( .A1(n6320), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n4908) );
  OAI22_X1 U6115 ( .A1(n5820), .A2(n6309), .B1(n5149), .B2(n4915), .ZN(n4906)
         );
  AOI21_X1 U6116 ( .B1(n6347), .B2(n4917), .A(n4906), .ZN(n4907) );
  OAI211_X1 U6117 ( .C1(n4920), .C2(n6351), .A(n4908), .B(n4907), .ZN(U3071)
         );
  NAND2_X1 U6118 ( .A1(n6320), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n4911) );
  OAI22_X1 U6119 ( .A1(n5832), .A2(n6309), .B1(n5161), .B2(n4915), .ZN(n4909)
         );
  AOI21_X1 U6120 ( .B1(n6359), .B2(n4917), .A(n4909), .ZN(n4910) );
  OAI211_X1 U6121 ( .C1(n4920), .C2(n6363), .A(n4911), .B(n4910), .ZN(U3074)
         );
  NAND2_X1 U6122 ( .A1(n6320), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4914) );
  OAI22_X1 U6123 ( .A1(n5828), .A2(n6309), .B1(n5155), .B2(n4915), .ZN(n4912)
         );
  AOI21_X1 U6124 ( .B1(n6353), .B2(n4917), .A(n4912), .ZN(n4913) );
  OAI211_X1 U6125 ( .C1(n4920), .C2(n6357), .A(n4914), .B(n4913), .ZN(U3073)
         );
  NAND2_X1 U6126 ( .A1(n6320), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4919) );
  OAI22_X1 U6127 ( .A1(n5839), .A2(n6309), .B1(n5167), .B2(n4915), .ZN(n4916)
         );
  AOI21_X1 U6128 ( .B1(n6366), .B2(n4917), .A(n4916), .ZN(n4918) );
  OAI211_X1 U6129 ( .C1(n4920), .C2(n6374), .A(n4919), .B(n4918), .ZN(U3075)
         );
  AOI21_X1 U6130 ( .B1(n4924), .B2(n4923), .A(n4922), .ZN(n5613) );
  INV_X1 U6131 ( .A(n5613), .ZN(n5052) );
  INV_X1 U6132 ( .A(EAX_REG_14__SCAN_IN), .ZN(n6610) );
  OAI222_X1 U6133 ( .A1(n5052), .A2(n5914), .B1(n5203), .B2(n4925), .C1(n5472), 
        .C2(n6610), .ZN(U2877) );
  OAI21_X1 U6134 ( .B1(n6367), .B2(n4959), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n4926) );
  OAI211_X1 U6135 ( .C1(n4927), .C2(n4933), .A(n4926), .B(n5797), .ZN(n4932)
         );
  NAND2_X1 U6136 ( .A1(n4929), .A2(n4928), .ZN(n4956) );
  AOI211_X1 U6137 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n4956), .A(n5132), .B(
        n4930), .ZN(n4931) );
  NAND2_X1 U6138 ( .A1(n4932), .A2(n4931), .ZN(n4955) );
  NAND2_X1 U6139 ( .A1(n4955), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n4936)
         );
  NOR2_X1 U6140 ( .A1(n4933), .A2(n5791), .ZN(n4997) );
  AOI22_X1 U6141 ( .A1(n4997), .A2(n6059), .B1(n2977), .B2(n5138), .ZN(n4957)
         );
  OAI22_X1 U6142 ( .A1(n5816), .A2(n4957), .B1(n5183), .B2(n4956), .ZN(n4934)
         );
  AOI21_X1 U6143 ( .B1(n6326), .B2(n4959), .A(n4934), .ZN(n4935) );
  OAI211_X1 U6144 ( .C1(n4962), .C2(n6330), .A(n4936), .B(n4935), .ZN(U3118)
         );
  NAND2_X1 U6145 ( .A1(n4955), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n4939)
         );
  OAI22_X1 U6146 ( .A1(n5812), .A2(n4957), .B1(n5177), .B2(n4956), .ZN(n4937)
         );
  AOI21_X1 U6147 ( .B1(n6343), .B2(n4959), .A(n4937), .ZN(n4938) );
  OAI211_X1 U6148 ( .C1(n4962), .C2(n6387), .A(n4939), .B(n4938), .ZN(U3117)
         );
  NAND2_X1 U6149 ( .A1(n4955), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n4942)
         );
  OAI22_X1 U6150 ( .A1(n5839), .A2(n4957), .B1(n5167), .B2(n4956), .ZN(n4940)
         );
  AOI21_X1 U6151 ( .B1(n6366), .B2(n4959), .A(n4940), .ZN(n4941) );
  OAI211_X1 U6152 ( .C1(n4962), .C2(n6374), .A(n4942), .B(n4941), .ZN(U3123)
         );
  NAND2_X1 U6153 ( .A1(n4955), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n4945)
         );
  OAI22_X1 U6154 ( .A1(n5820), .A2(n4957), .B1(n5149), .B2(n4956), .ZN(n4943)
         );
  AOI21_X1 U6155 ( .B1(n6347), .B2(n4959), .A(n4943), .ZN(n4944) );
  OAI211_X1 U6156 ( .C1(n4962), .C2(n6351), .A(n4945), .B(n4944), .ZN(U3119)
         );
  NAND2_X1 U6157 ( .A1(n4955), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n4948)
         );
  OAI22_X1 U6158 ( .A1(n5832), .A2(n4957), .B1(n5161), .B2(n4956), .ZN(n4946)
         );
  AOI21_X1 U6159 ( .B1(n6359), .B2(n4959), .A(n4946), .ZN(n4947) );
  OAI211_X1 U6160 ( .C1(n4962), .C2(n6363), .A(n4948), .B(n4947), .ZN(U3122)
         );
  NAND2_X1 U6161 ( .A1(n4955), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n4951)
         );
  OAI22_X1 U6162 ( .A1(n5824), .A2(n4957), .B1(n5143), .B2(n4956), .ZN(n4949)
         );
  AOI21_X1 U6163 ( .B1(n6297), .B2(n4959), .A(n4949), .ZN(n4950) );
  OAI211_X1 U6164 ( .C1(n4962), .C2(n6301), .A(n4951), .B(n4950), .ZN(U3120)
         );
  NAND2_X1 U6165 ( .A1(n4955), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n4954)
         );
  OAI22_X1 U6166 ( .A1(n5828), .A2(n4957), .B1(n5155), .B2(n4956), .ZN(n4952)
         );
  AOI21_X1 U6167 ( .B1(n6353), .B2(n4959), .A(n4952), .ZN(n4953) );
  OAI211_X1 U6168 ( .C1(n4962), .C2(n6357), .A(n4954), .B(n4953), .ZN(U3121)
         );
  NAND2_X1 U6169 ( .A1(n4955), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n4961)
         );
  OAI22_X1 U6170 ( .A1(n5807), .A2(n4957), .B1(n5173), .B2(n4956), .ZN(n4958)
         );
  AOI21_X1 U6171 ( .B1(n5809), .B2(n4959), .A(n4958), .ZN(n4960) );
  OAI211_X1 U6172 ( .C1(n4962), .C2(n6377), .A(n4961), .B(n4960), .ZN(U3116)
         );
  NOR2_X1 U6173 ( .A1(n4922), .A2(n4964), .ZN(n4965) );
  OR2_X1 U6174 ( .A1(n4963), .A2(n4965), .ZN(n5598) );
  AOI22_X1 U6175 ( .A1(n5499), .A2(DATAI_15_), .B1(n6103), .B2(
        EAX_REG_15__SCAN_IN), .ZN(n4966) );
  OAI21_X1 U6176 ( .B1(n5598), .B2(n5914), .A(n4966), .ZN(U2876) );
  INV_X1 U6177 ( .A(n5426), .ZN(n4979) );
  AOI21_X1 U6178 ( .B1(n4967), .B2(n4968), .A(n4979), .ZN(n5271) );
  AOI22_X1 U6179 ( .A1(n6186), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .B1(n3668), 
        .B2(REIP_REG_5__SCAN_IN), .ZN(n4969) );
  OAI21_X1 U6180 ( .B1(n6195), .B2(n5265), .A(n4969), .ZN(n4970) );
  AOI21_X1 U6181 ( .B1(n5271), .B2(n6165), .A(n4970), .ZN(n4971) );
  OAI21_X1 U6182 ( .B1(n6169), .B2(n4972), .A(n4971), .ZN(U2981) );
  INV_X1 U6183 ( .A(n5271), .ZN(n4976) );
  OAI222_X1 U6184 ( .A1(n4976), .A2(n5914), .B1(n5203), .B2(n4973), .C1(n5472), 
        .C2(n3771), .ZN(U2886) );
  INV_X1 U6185 ( .A(EBX_REG_5__SCAN_IN), .ZN(n4975) );
  OAI222_X1 U6186 ( .A1(n4976), .A2(n6092), .B1(n6096), .B2(n4975), .C1(n4974), 
        .C2(n6091), .ZN(U2854) );
  NOR2_X1 U6187 ( .A1(n5030), .A2(n4977), .ZN(n4980) );
  NOR2_X1 U6188 ( .A1(n5426), .A2(n4978), .ZN(n5042) );
  NAND2_X1 U6189 ( .A1(n4980), .A2(n5042), .ZN(n5041) );
  AND2_X1 U6190 ( .A1(n4980), .A2(n4979), .ZN(n4982) );
  OR2_X1 U6191 ( .A1(n4982), .A2(n4981), .ZN(n4983) );
  AOI22_X1 U6192 ( .A1(n5499), .A2(DATAI_8_), .B1(n6103), .B2(
        EAX_REG_8__SCAN_IN), .ZN(n4984) );
  OAI21_X1 U6193 ( .B1(n5228), .B2(n5914), .A(n4984), .ZN(U2883) );
  NOR2_X1 U6194 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4985), .ZN(n4998)
         );
  OAI21_X1 U6195 ( .B1(n4986), .B2(n6303), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n4988) );
  AND2_X1 U6196 ( .A1(n4988), .A2(n4987), .ZN(n4993) );
  INV_X1 U6197 ( .A(n4989), .ZN(n4990) );
  OR2_X1 U6198 ( .A1(n5796), .A2(n4990), .ZN(n4995) );
  AOI21_X1 U6199 ( .B1(n4995), .B2(STATE2_REG_2__SCAN_IN), .A(n4991), .ZN(
        n5092) );
  INV_X1 U6200 ( .A(n5092), .ZN(n4992) );
  AOI211_X1 U6201 ( .C1(n5797), .C2(n4993), .A(n5132), .B(n4992), .ZN(n4994)
         );
  NAND2_X1 U6202 ( .A1(n5020), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n5001) );
  INV_X1 U6203 ( .A(n4995), .ZN(n5096) );
  AOI22_X1 U6204 ( .A1(n4997), .A2(n4996), .B1(n5138), .B2(n5096), .ZN(n5022)
         );
  INV_X1 U6205 ( .A(n4998), .ZN(n5021) );
  OAI22_X1 U6206 ( .A1(n5816), .A2(n5022), .B1(n5183), .B2(n5021), .ZN(n4999)
         );
  AOI21_X1 U6207 ( .B1(n6303), .B2(n6319), .A(n4999), .ZN(n5000) );
  OAI211_X1 U6208 ( .C1(n5026), .C2(n6323), .A(n5001), .B(n5000), .ZN(U3054)
         );
  NAND2_X1 U6209 ( .A1(n5020), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n5004) );
  OAI22_X1 U6210 ( .A1(n5812), .A2(n5022), .B1(n5177), .B2(n5021), .ZN(n5002)
         );
  AOI21_X1 U6211 ( .B1(n6303), .B2(n6313), .A(n5002), .ZN(n5003) );
  OAI211_X1 U6212 ( .C1(n6390), .C2(n5026), .A(n5004), .B(n5003), .ZN(U3053)
         );
  NAND2_X1 U6213 ( .A1(n5020), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n5007) );
  OAI22_X1 U6214 ( .A1(n5824), .A2(n5022), .B1(n5143), .B2(n5021), .ZN(n5005)
         );
  AOI21_X1 U6215 ( .B1(n6303), .B2(n5146), .A(n5005), .ZN(n5006) );
  OAI211_X1 U6216 ( .C1(n5026), .C2(n5144), .A(n5007), .B(n5006), .ZN(U3056)
         );
  NAND2_X1 U6217 ( .A1(n5020), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n5010) );
  OAI22_X1 U6218 ( .A1(n5828), .A2(n5022), .B1(n5155), .B2(n5021), .ZN(n5008)
         );
  AOI21_X1 U6219 ( .B1(n6303), .B2(n5158), .A(n5008), .ZN(n5009) );
  OAI211_X1 U6220 ( .C1(n5026), .C2(n5156), .A(n5010), .B(n5009), .ZN(U3057)
         );
  NAND2_X1 U6221 ( .A1(n5020), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n5013) );
  OAI22_X1 U6222 ( .A1(n5807), .A2(n5022), .B1(n5173), .B2(n5021), .ZN(n5011)
         );
  AOI21_X1 U6223 ( .B1(n6303), .B2(n6310), .A(n5011), .ZN(n5012) );
  OAI211_X1 U6224 ( .C1(n5026), .C2(n6379), .A(n5013), .B(n5012), .ZN(U3052)
         );
  NAND2_X1 U6225 ( .A1(n5020), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n5016) );
  OAI22_X1 U6226 ( .A1(n5832), .A2(n5022), .B1(n5161), .B2(n5021), .ZN(n5014)
         );
  AOI21_X1 U6227 ( .B1(n6303), .B2(n5164), .A(n5014), .ZN(n5015) );
  OAI211_X1 U6228 ( .C1(n5026), .C2(n5162), .A(n5016), .B(n5015), .ZN(U3058)
         );
  NAND2_X1 U6229 ( .A1(n5020), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n5019) );
  OAI22_X1 U6230 ( .A1(n5839), .A2(n5022), .B1(n5167), .B2(n5021), .ZN(n5017)
         );
  AOI21_X1 U6231 ( .B1(n6303), .B2(n5170), .A(n5017), .ZN(n5018) );
  OAI211_X1 U6232 ( .C1(n5026), .C2(n5168), .A(n5019), .B(n5018), .ZN(U3059)
         );
  NAND2_X1 U6233 ( .A1(n5020), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n5025) );
  OAI22_X1 U6234 ( .A1(n5820), .A2(n5022), .B1(n5149), .B2(n5021), .ZN(n5023)
         );
  AOI21_X1 U6235 ( .B1(n6303), .B2(n5152), .A(n5023), .ZN(n5024) );
  OAI211_X1 U6236 ( .C1(n5026), .C2(n5150), .A(n5025), .B(n5024), .ZN(U3055)
         );
  OAI21_X1 U6237 ( .B1(n5029), .B2(n5028), .A(n5027), .ZN(n6240) );
  OR2_X1 U6238 ( .A1(n5426), .A2(n4977), .ZN(n5193) );
  XOR2_X1 U6239 ( .A(n5030), .B(n5193), .Z(n5037) );
  NAND2_X1 U6240 ( .A1(n3668), .A2(REIP_REG_7__SCAN_IN), .ZN(n6237) );
  NAND2_X1 U6241 ( .A1(n6186), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n5031)
         );
  OAI211_X1 U6242 ( .C1(n6195), .C2(n5070), .A(n6237), .B(n5031), .ZN(n5032)
         );
  AOI21_X1 U6243 ( .B1(n5037), .B2(n6165), .A(n5032), .ZN(n5033) );
  OAI21_X1 U6244 ( .B1(n6240), .B2(n6169), .A(n5033), .ZN(U2979) );
  AND2_X1 U6245 ( .A1(n5051), .A2(n5034), .ZN(n5035) );
  OR2_X1 U6246 ( .A1(n5035), .A2(n5064), .ZN(n5748) );
  OAI222_X1 U6247 ( .A1(n5598), .A2(n6092), .B1(n6096), .B2(n5036), .C1(n5748), 
        .C2(n6091), .ZN(U2844) );
  INV_X1 U6248 ( .A(n5037), .ZN(n5081) );
  AND2_X1 U6249 ( .A1(n5197), .A2(n5038), .ZN(n5039) );
  NOR2_X1 U6250 ( .A1(n5059), .A2(n5039), .ZN(n6239) );
  AOI22_X1 U6251 ( .A1(n6087), .A2(n6239), .B1(EBX_REG_7__SCAN_IN), .B2(n5462), 
        .ZN(n5040) );
  OAI21_X1 U6252 ( .B1(n5081), .B2(n6092), .A(n5040), .ZN(U2852) );
  INV_X1 U6253 ( .A(n5041), .ZN(n5044) );
  NAND2_X1 U6254 ( .A1(n5042), .A2(n5428), .ZN(n5055) );
  OAI21_X1 U6255 ( .B1(n5044), .B2(n5043), .A(n5055), .ZN(n6029) );
  INV_X1 U6256 ( .A(n5190), .ZN(n5045) );
  AOI21_X1 U6257 ( .B1(n5046), .B2(n5061), .A(n5045), .ZN(n6220) );
  AOI22_X1 U6258 ( .A1(n6087), .A2(n6220), .B1(EBX_REG_9__SCAN_IN), .B2(n5462), 
        .ZN(n5047) );
  OAI21_X1 U6259 ( .B1(n6029), .B2(n6092), .A(n5047), .ZN(U2850) );
  NAND2_X1 U6260 ( .A1(n5049), .A2(n5048), .ZN(n5050) );
  NAND2_X1 U6261 ( .A1(n5051), .A2(n5050), .ZN(n5760) );
  INV_X1 U6262 ( .A(EBX_REG_14__SCAN_IN), .ZN(n6663) );
  OAI222_X1 U6263 ( .A1(n5760), .A2(n6091), .B1(n6096), .B2(n6663), .C1(n6092), 
        .C2(n5052), .ZN(U2845) );
  NOR2_X1 U6264 ( .A1(n5426), .A2(n5053), .ZN(n5054) );
  AND2_X1 U6265 ( .A1(n5428), .A2(n5054), .ZN(n5496) );
  AOI21_X1 U6266 ( .B1(n5056), .B2(n5055), .A(n5496), .ZN(n5300) );
  INV_X1 U6267 ( .A(n5300), .ZN(n5192) );
  AOI22_X1 U6268 ( .A1(n5499), .A2(DATAI_10_), .B1(n6103), .B2(
        EAX_REG_10__SCAN_IN), .ZN(n5057) );
  OAI21_X1 U6269 ( .B1(n5192), .B2(n5914), .A(n5057), .ZN(U2881) );
  OR2_X1 U6270 ( .A1(n5059), .A2(n5058), .ZN(n5060) );
  NAND2_X1 U6271 ( .A1(n5061), .A2(n5060), .ZN(n6228) );
  INV_X1 U6272 ( .A(EBX_REG_8__SCAN_IN), .ZN(n6671) );
  OAI222_X1 U6273 ( .A1(n6228), .A2(n6091), .B1(n6096), .B2(n6671), .C1(n6092), 
        .C2(n5228), .ZN(U2851) );
  OAI222_X1 U6274 ( .A1(n5914), .A2(n5081), .B1(n5203), .B2(n6632), .C1(n5472), 
        .C2(n3739), .ZN(U2884) );
  OR2_X1 U6275 ( .A1(n5064), .A2(n5063), .ZN(n5065) );
  NAND2_X1 U6276 ( .A1(n5942), .A2(n5065), .ZN(n6011) );
  INV_X1 U6277 ( .A(EBX_REG_16__SCAN_IN), .ZN(n5069) );
  OAI21_X1 U6278 ( .B1(n4963), .B2(n5068), .A(n5067), .ZN(n5590) );
  OAI222_X1 U6279 ( .A1(n6011), .A2(n6091), .B1(n6096), .B2(n5069), .C1(n6092), 
        .C2(n5590), .ZN(U2843) );
  INV_X1 U6280 ( .A(n5070), .ZN(n5077) );
  AOI22_X1 U6281 ( .A1(EBX_REG_7__SCAN_IN), .A2(n6695), .B1(n6697), .B2(n6239), 
        .ZN(n5072) );
  NAND2_X1 U6282 ( .A1(n5071), .A2(n6074), .ZN(n6691) );
  OAI211_X1 U6283 ( .C1(n6693), .C2(n5073), .A(n5072), .B(n6691), .ZN(n5076)
         );
  INV_X1 U6284 ( .A(REIP_REG_6__SCAN_IN), .ZN(n6480) );
  INV_X1 U6285 ( .A(n6042), .ZN(n5074) );
  NAND2_X1 U6286 ( .A1(n6069), .A2(n5074), .ZN(n6047) );
  NOR2_X1 U6287 ( .A1(n6047), .A2(n6477), .ZN(n5263) );
  NAND2_X1 U6288 ( .A1(REIP_REG_5__SCAN_IN), .A2(n5263), .ZN(n5217) );
  NOR3_X1 U6289 ( .A1(REIP_REG_7__SCAN_IN), .A2(n6480), .A3(n5217), .ZN(n5075)
         );
  AOI211_X1 U6290 ( .C1(n6077), .C2(n5077), .A(n5076), .B(n5075), .ZN(n5080)
         );
  NOR2_X1 U6291 ( .A1(REIP_REG_6__SCAN_IN), .A2(n5217), .ZN(n6039) );
  OAI21_X1 U6292 ( .B1(n6018), .B2(n5078), .A(n6074), .ZN(n6036) );
  OAI21_X1 U6293 ( .B1(n6039), .B2(n6036), .A(REIP_REG_7__SCAN_IN), .ZN(n5079)
         );
  OAI211_X1 U6294 ( .C1(n5081), .C2(n5995), .A(n5080), .B(n5079), .ZN(U2820)
         );
  OAI21_X1 U6295 ( .B1(n5084), .B2(n5083), .A(n5082), .ZN(n6232) );
  NAND2_X1 U6296 ( .A1(n3668), .A2(REIP_REG_8__SCAN_IN), .ZN(n6229) );
  NAND2_X1 U6297 ( .A1(n6186), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n5085)
         );
  OAI211_X1 U6298 ( .C1(n6195), .C2(n5221), .A(n6229), .B(n5085), .ZN(n5086)
         );
  AOI21_X1 U6299 ( .B1(n5087), .B2(n6165), .A(n5086), .ZN(n5088) );
  OAI21_X1 U6300 ( .B1(n6232), .B2(n6169), .A(n5088), .ZN(U2978) );
  INV_X1 U6301 ( .A(DATAI_9_), .ZN(n6731) );
  INV_X1 U6302 ( .A(EAX_REG_9__SCAN_IN), .ZN(n6121) );
  OAI222_X1 U6303 ( .A1(n6029), .A2(n5914), .B1(n5203), .B2(n6731), .C1(n5472), 
        .C2(n6121), .ZN(U2882) );
  NAND3_X1 U6304 ( .A1(n5127), .A2(n5089), .A3(n6391), .ZN(n5090) );
  AOI21_X1 U6305 ( .B1(n5090), .B2(n5800), .A(n5097), .ZN(n5095) );
  NOR2_X1 U6306 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5091), .ZN(n5098)
         );
  OAI211_X1 U6307 ( .C1(n6717), .C2(n5098), .A(n5093), .B(n5092), .ZN(n5094)
         );
  NAND2_X1 U6308 ( .A1(n5120), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n5101) );
  AOI22_X1 U6309 ( .A1(n5097), .A2(n5797), .B1(n5096), .B2(n5132), .ZN(n5122)
         );
  INV_X1 U6310 ( .A(n5098), .ZN(n5121) );
  OAI22_X1 U6311 ( .A1(n5828), .A2(n5122), .B1(n5155), .B2(n5121), .ZN(n5099)
         );
  AOI21_X1 U6312 ( .B1(n5158), .B2(n5124), .A(n5099), .ZN(n5100) );
  OAI211_X1 U6313 ( .C1(n5127), .C2(n5156), .A(n5101), .B(n5100), .ZN(U3025)
         );
  NAND2_X1 U6314 ( .A1(n5120), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n5104) );
  OAI22_X1 U6315 ( .A1(n5807), .A2(n5122), .B1(n5173), .B2(n5121), .ZN(n5102)
         );
  AOI21_X1 U6316 ( .B1(n6310), .B2(n5124), .A(n5102), .ZN(n5103) );
  OAI211_X1 U6317 ( .C1(n5127), .C2(n6379), .A(n5104), .B(n5103), .ZN(U3020)
         );
  NAND2_X1 U6318 ( .A1(n5120), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n5107) );
  OAI22_X1 U6319 ( .A1(n5839), .A2(n5122), .B1(n5167), .B2(n5121), .ZN(n5105)
         );
  AOI21_X1 U6320 ( .B1(n5170), .B2(n5124), .A(n5105), .ZN(n5106) );
  OAI211_X1 U6321 ( .C1(n5127), .C2(n5168), .A(n5107), .B(n5106), .ZN(U3027)
         );
  NAND2_X1 U6322 ( .A1(n5120), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n5110) );
  OAI22_X1 U6323 ( .A1(n5812), .A2(n5122), .B1(n5177), .B2(n5121), .ZN(n5108)
         );
  AOI21_X1 U6324 ( .B1(n6313), .B2(n5124), .A(n5108), .ZN(n5109) );
  OAI211_X1 U6325 ( .C1(n5127), .C2(n6390), .A(n5110), .B(n5109), .ZN(U3021)
         );
  NAND2_X1 U6326 ( .A1(n5120), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n5113) );
  OAI22_X1 U6327 ( .A1(n5824), .A2(n5122), .B1(n5143), .B2(n5121), .ZN(n5111)
         );
  AOI21_X1 U6328 ( .B1(n5146), .B2(n5124), .A(n5111), .ZN(n5112) );
  OAI211_X1 U6329 ( .C1(n5127), .C2(n5144), .A(n5113), .B(n5112), .ZN(U3024)
         );
  NAND2_X1 U6330 ( .A1(n5120), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n5116) );
  OAI22_X1 U6331 ( .A1(n5832), .A2(n5122), .B1(n5161), .B2(n5121), .ZN(n5114)
         );
  AOI21_X1 U6332 ( .B1(n5164), .B2(n5124), .A(n5114), .ZN(n5115) );
  OAI211_X1 U6333 ( .C1(n5127), .C2(n5162), .A(n5116), .B(n5115), .ZN(U3026)
         );
  NAND2_X1 U6334 ( .A1(n5120), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n5119) );
  OAI22_X1 U6335 ( .A1(n5820), .A2(n5122), .B1(n5149), .B2(n5121), .ZN(n5117)
         );
  AOI21_X1 U6336 ( .B1(n5152), .B2(n5124), .A(n5117), .ZN(n5118) );
  OAI211_X1 U6337 ( .C1(n5127), .C2(n5150), .A(n5119), .B(n5118), .ZN(U3023)
         );
  NAND2_X1 U6338 ( .A1(n5120), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n5126) );
  OAI22_X1 U6339 ( .A1(n5816), .A2(n5122), .B1(n5183), .B2(n5121), .ZN(n5123)
         );
  AOI21_X1 U6340 ( .B1(n6319), .B2(n5124), .A(n5123), .ZN(n5125) );
  OAI211_X1 U6341 ( .C1(n5127), .C2(n6323), .A(n5126), .B(n5125), .ZN(U3022)
         );
  OAI21_X1 U6342 ( .B1(n5185), .B2(n5129), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n5130) );
  NAND2_X1 U6343 ( .A1(n5130), .A2(n5797), .ZN(n5141) );
  INV_X1 U6344 ( .A(n5141), .ZN(n5134) );
  INV_X1 U6345 ( .A(n5131), .ZN(n5140) );
  INV_X1 U6346 ( .A(n5132), .ZN(n5794) );
  NOR2_X1 U6347 ( .A1(n5794), .A2(n6419), .ZN(n5133) );
  AOI22_X1 U6348 ( .A1(n5134), .A2(n5140), .B1(n5796), .B2(n5133), .ZN(n5188)
         );
  NOR2_X1 U6349 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5135), .ZN(n5142)
         );
  OAI22_X1 U6350 ( .A1(n6661), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B1(n6717), .B2(n5142), .ZN(n5136) );
  INV_X1 U6351 ( .A(n5136), .ZN(n5139) );
  NOR2_X1 U6352 ( .A1(n5138), .A2(n5137), .ZN(n5804) );
  OAI211_X1 U6353 ( .C1(n5141), .C2(n5140), .A(n5139), .B(n5804), .ZN(n5181)
         );
  NAND2_X1 U6354 ( .A1(n5181), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n5148)
         );
  INV_X1 U6355 ( .A(n5142), .ZN(n5182) );
  OAI22_X1 U6356 ( .A1(n6373), .A2(n5144), .B1(n5143), .B2(n5182), .ZN(n5145)
         );
  AOI21_X1 U6357 ( .B1(n5146), .B2(n5185), .A(n5145), .ZN(n5147) );
  OAI211_X1 U6358 ( .C1(n5188), .C2(n5824), .A(n5148), .B(n5147), .ZN(U3104)
         );
  NAND2_X1 U6359 ( .A1(n5181), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n5154)
         );
  OAI22_X1 U6360 ( .A1(n6373), .A2(n5150), .B1(n5149), .B2(n5182), .ZN(n5151)
         );
  AOI21_X1 U6361 ( .B1(n5152), .B2(n5185), .A(n5151), .ZN(n5153) );
  OAI211_X1 U6362 ( .C1(n5188), .C2(n5820), .A(n5154), .B(n5153), .ZN(U3103)
         );
  NAND2_X1 U6363 ( .A1(n5181), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n5160)
         );
  OAI22_X1 U6364 ( .A1(n6373), .A2(n5156), .B1(n5155), .B2(n5182), .ZN(n5157)
         );
  AOI21_X1 U6365 ( .B1(n5158), .B2(n5185), .A(n5157), .ZN(n5159) );
  OAI211_X1 U6366 ( .C1(n5188), .C2(n5828), .A(n5160), .B(n5159), .ZN(U3105)
         );
  NAND2_X1 U6367 ( .A1(n5181), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n5166)
         );
  OAI22_X1 U6368 ( .A1(n6373), .A2(n5162), .B1(n5161), .B2(n5182), .ZN(n5163)
         );
  AOI21_X1 U6369 ( .B1(n5164), .B2(n5185), .A(n5163), .ZN(n5165) );
  OAI211_X1 U6370 ( .C1(n5188), .C2(n5832), .A(n5166), .B(n5165), .ZN(U3106)
         );
  NAND2_X1 U6371 ( .A1(n5181), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n5172)
         );
  OAI22_X1 U6372 ( .A1(n6373), .A2(n5168), .B1(n5167), .B2(n5182), .ZN(n5169)
         );
  AOI21_X1 U6373 ( .B1(n5170), .B2(n5185), .A(n5169), .ZN(n5171) );
  OAI211_X1 U6374 ( .C1(n5188), .C2(n5839), .A(n5172), .B(n5171), .ZN(U3107)
         );
  NAND2_X1 U6375 ( .A1(n5181), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n5176)
         );
  OAI22_X1 U6376 ( .A1(n6373), .A2(n6379), .B1(n5173), .B2(n5182), .ZN(n5174)
         );
  AOI21_X1 U6377 ( .B1(n6310), .B2(n5185), .A(n5174), .ZN(n5175) );
  OAI211_X1 U6378 ( .C1(n5188), .C2(n5807), .A(n5176), .B(n5175), .ZN(U3100)
         );
  NAND2_X1 U6379 ( .A1(n5181), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n5180)
         );
  OAI22_X1 U6380 ( .A1(n6373), .A2(n6390), .B1(n5177), .B2(n5182), .ZN(n5178)
         );
  AOI21_X1 U6381 ( .B1(n6313), .B2(n5185), .A(n5178), .ZN(n5179) );
  OAI211_X1 U6382 ( .C1(n5188), .C2(n5812), .A(n5180), .B(n5179), .ZN(U3101)
         );
  NAND2_X1 U6383 ( .A1(n5181), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n5187)
         );
  OAI22_X1 U6384 ( .A1(n6373), .A2(n6323), .B1(n5183), .B2(n5182), .ZN(n5184)
         );
  AOI21_X1 U6385 ( .B1(n6319), .B2(n5185), .A(n5184), .ZN(n5186) );
  OAI211_X1 U6386 ( .C1(n5188), .C2(n5816), .A(n5187), .B(n5186), .ZN(U3102)
         );
  AND2_X1 U6387 ( .A1(n5190), .A2(n5189), .ZN(n5191) );
  OR2_X1 U6388 ( .A1(n5191), .A2(n6013), .ZN(n6211) );
  INV_X1 U6389 ( .A(EBX_REG_10__SCAN_IN), .ZN(n5276) );
  OAI222_X1 U6390 ( .A1(n6211), .A2(n6091), .B1(n6096), .B2(n5276), .C1(n6092), 
        .C2(n5192), .ZN(U2849) );
  INV_X1 U6391 ( .A(n5193), .ZN(n5194) );
  AOI21_X1 U6392 ( .B1(n4977), .B2(n5426), .A(n5194), .ZN(n6173) );
  INV_X1 U6393 ( .A(n5195), .ZN(n5199) );
  INV_X1 U6394 ( .A(n5196), .ZN(n5198) );
  OAI21_X1 U6395 ( .B1(n5199), .B2(n5198), .A(n5197), .ZN(n6250) );
  OAI22_X1 U6396 ( .A1(n6091), .A2(n6250), .B1(n5200), .B2(n6096), .ZN(n5201)
         );
  AOI21_X1 U6397 ( .B1(n6173), .B2(n6088), .A(n5201), .ZN(n5202) );
  INV_X1 U6398 ( .A(n5202), .ZN(U2853) );
  INV_X1 U6399 ( .A(n6173), .ZN(n5204) );
  INV_X1 U6400 ( .A(EAX_REG_6__SCAN_IN), .ZN(n6126) );
  OAI222_X1 U6401 ( .A1(n5204), .A2(n5914), .B1(n5203), .B2(n6733), .C1(n6126), 
        .C2(n5472), .ZN(U2885) );
  NAND2_X1 U6402 ( .A1(n5207), .A2(n3154), .ZN(n5205) );
  NAND2_X1 U6403 ( .A1(n5205), .A2(n5995), .ZN(n6073) );
  INV_X1 U6404 ( .A(n6073), .ZN(n6056) );
  OAI21_X1 U6405 ( .B1(n6018), .B2(REIP_REG_1__SCAN_IN), .A(n6074), .ZN(n6055)
         );
  NAND2_X1 U6406 ( .A1(n6695), .A2(EBX_REG_2__SCAN_IN), .ZN(n5213) );
  NAND2_X1 U6407 ( .A1(n5207), .A2(n5206), .ZN(n6048) );
  INV_X1 U6408 ( .A(n6048), .ZN(n6071) );
  AOI22_X1 U6409 ( .A1(n6071), .A2(n5208), .B1(n6697), .B2(n6279), .ZN(n5212)
         );
  INV_X1 U6410 ( .A(n6194), .ZN(n5209) );
  AOI22_X1 U6411 ( .A1(n6078), .A2(PHYADDRPOINTER_REG_2__SCAN_IN), .B1(n6077), 
        .B2(n5209), .ZN(n5211) );
  INV_X1 U6412 ( .A(REIP_REG_2__SCAN_IN), .ZN(n6054) );
  NAND3_X1 U6413 ( .A1(n6069), .A2(REIP_REG_1__SCAN_IN), .A3(n6054), .ZN(n5210) );
  NAND4_X1 U6414 ( .A1(n5213), .A2(n5212), .A3(n5211), .A4(n5210), .ZN(n5214)
         );
  AOI21_X1 U6415 ( .B1(REIP_REG_2__SCAN_IN), .B2(n6055), .A(n5214), .ZN(n5215)
         );
  OAI21_X1 U6416 ( .B1(n6056), .B2(n5216), .A(n5215), .ZN(U2825) );
  NAND2_X1 U6417 ( .A1(REIP_REG_7__SCAN_IN), .A2(REIP_REG_6__SCAN_IN), .ZN(
        n5218) );
  INV_X1 U6418 ( .A(REIP_REG_8__SCAN_IN), .ZN(n6483) );
  OAI21_X1 U6419 ( .B1(n5218), .B2(n5217), .A(n6483), .ZN(n5226) );
  INV_X1 U6420 ( .A(n5219), .ZN(n6027) );
  OAI21_X1 U6421 ( .B1(n6018), .B2(n6027), .A(n6074), .ZN(n6028) );
  INV_X1 U6422 ( .A(n6695), .ZN(n6043) );
  INV_X1 U6423 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n5220) );
  OAI22_X1 U6424 ( .A1(n6043), .A2(n6671), .B1(n5220), .B2(n6693), .ZN(n5225)
         );
  INV_X1 U6425 ( .A(n5221), .ZN(n5222) );
  INV_X1 U6426 ( .A(n6691), .ZN(n6045) );
  AOI21_X1 U6427 ( .B1(n6077), .B2(n5222), .A(n6045), .ZN(n5223) );
  OAI21_X1 U6428 ( .B1(n6085), .B2(n6228), .A(n5223), .ZN(n5224) );
  AOI211_X1 U6429 ( .C1(n5226), .C2(n6028), .A(n5225), .B(n5224), .ZN(n5227)
         );
  OAI21_X1 U6430 ( .B1(n5228), .B2(n5995), .A(n5227), .ZN(U2819) );
  AOI22_X1 U6431 ( .A1(EBX_REG_13__SCAN_IN), .A2(n6695), .B1(n6697), .B2(n5954), .ZN(n5229) );
  OAI211_X1 U6432 ( .C1(n6693), .C2(n5230), .A(n5229), .B(n6691), .ZN(n5237)
         );
  INV_X1 U6433 ( .A(REIP_REG_12__SCAN_IN), .ZN(n6635) );
  AND3_X1 U6434 ( .A1(n6069), .A2(n5231), .A3(n6635), .ZN(n5434) );
  OAI21_X1 U6435 ( .B1(n6018), .B2(n5231), .A(n6074), .ZN(n6016) );
  OAI21_X1 U6436 ( .B1(n5434), .B2(n6016), .A(REIP_REG_13__SCAN_IN), .ZN(n5234) );
  OR3_X1 U6437 ( .A1(n6018), .A2(REIP_REG_13__SCAN_IN), .A3(n5232), .ZN(n5233)
         );
  OAI211_X1 U6438 ( .C1(n5235), .C2(n6702), .A(n5234), .B(n5233), .ZN(n5236)
         );
  NOR2_X1 U6439 ( .A1(n5237), .A2(n5236), .ZN(n5238) );
  OAI21_X1 U6440 ( .B1(n5623), .B2(n5995), .A(n5238), .ZN(U2814) );
  NAND2_X1 U6441 ( .A1(n5240), .A2(n5239), .ZN(n5241) );
  XNOR2_X1 U6442 ( .A(n5242), .B(n5241), .ZN(n6222) );
  NAND2_X1 U6443 ( .A1(n6222), .A2(n6191), .ZN(n5245) );
  NAND2_X1 U6444 ( .A1(n3668), .A2(REIP_REG_9__SCAN_IN), .ZN(n6218) );
  OAI21_X1 U6445 ( .B1(n5618), .B2(n6567), .A(n6218), .ZN(n5243) );
  AOI21_X1 U6446 ( .B1(n6164), .B2(n6030), .A(n5243), .ZN(n5244) );
  OAI211_X1 U6447 ( .C1(n5634), .C2(n6029), .A(n5245), .B(n5244), .ZN(U2977)
         );
  NAND2_X1 U6448 ( .A1(n5937), .A2(n5247), .ZN(n5248) );
  NAND2_X1 U6449 ( .A1(n5304), .A2(n5248), .ZN(n5996) );
  NOR2_X2 U6450 ( .A1(n6103), .A2(n5249), .ZN(n6100) );
  AOI22_X1 U6451 ( .A1(n6100), .A2(DATAI_18_), .B1(EAX_REG_18__SCAN_IN), .B2(
        n6103), .ZN(n5252) );
  AND2_X1 U6452 ( .A1(n3133), .A2(n3146), .ZN(n5250) );
  NAND2_X1 U6453 ( .A1(n6104), .A2(DATAI_2_), .ZN(n5251) );
  OAI211_X1 U6454 ( .C1(n5996), .C2(n5914), .A(n5252), .B(n5251), .ZN(U2873)
         );
  NAND2_X1 U6455 ( .A1(n6693), .A2(n6702), .ZN(n5258) );
  OAI22_X1 U6456 ( .A1(n5253), .A2(n6549), .B1(n6043), .B2(n4398), .ZN(n5257)
         );
  OAI22_X1 U6457 ( .A1(n6085), .A2(n5255), .B1(n5254), .B2(n6048), .ZN(n5256)
         );
  AOI211_X1 U6458 ( .C1(PHYADDRPOINTER_REG_0__SCAN_IN), .C2(n5258), .A(n5257), 
        .B(n5256), .ZN(n5259) );
  OAI21_X1 U6459 ( .B1(n6056), .B2(n5260), .A(n5259), .ZN(U2827) );
  MUX2_X1 U6460 ( .A(n5318), .B(n5262), .S(n5261), .Z(n5308) );
  XNOR2_X1 U6461 ( .A(n5944), .B(n5308), .ZN(n6000) );
  OAI222_X1 U6462 ( .A1(n6092), .A2(n5996), .B1(n6096), .B2(n5991), .C1(n6000), 
        .C2(n6091), .ZN(U2841) );
  OAI21_X1 U6463 ( .B1(n5263), .B2(REIP_REG_5__SCAN_IN), .A(n6036), .ZN(n5264)
         );
  OAI21_X1 U6464 ( .B1(n6702), .B2(n5265), .A(n5264), .ZN(n5270) );
  INV_X1 U6465 ( .A(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n5268) );
  AOI22_X1 U6466 ( .A1(EBX_REG_5__SCAN_IN), .A2(n6695), .B1(n6697), .B2(n5266), 
        .ZN(n5267) );
  OAI211_X1 U6467 ( .C1(n6693), .C2(n5268), .A(n5267), .B(n6691), .ZN(n5269)
         );
  AOI211_X1 U6468 ( .C1(n5271), .C2(n6073), .A(n5270), .B(n5269), .ZN(n5272)
         );
  INV_X1 U6469 ( .A(n5272), .ZN(U2822) );
  INV_X1 U6470 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n5275) );
  INV_X1 U6471 ( .A(REIP_REG_10__SCAN_IN), .ZN(n6486) );
  NAND3_X1 U6472 ( .A1(n6069), .A2(n6486), .A3(n5273), .ZN(n5274) );
  OAI211_X1 U6473 ( .C1(n6693), .C2(n5275), .A(n6691), .B(n5274), .ZN(n5281)
         );
  NOR2_X1 U6474 ( .A1(n6018), .A2(REIP_REG_9__SCAN_IN), .ZN(n6026) );
  OAI21_X1 U6475 ( .B1(n6028), .B2(n6026), .A(REIP_REG_10__SCAN_IN), .ZN(n5279) );
  OAI22_X1 U6476 ( .A1(n6043), .A2(n5276), .B1(n6085), .B2(n6211), .ZN(n5277)
         );
  INV_X1 U6477 ( .A(n5277), .ZN(n5278) );
  OAI211_X1 U6478 ( .C1(n6702), .C2(n5298), .A(n5279), .B(n5278), .ZN(n5280)
         );
  AOI211_X1 U6479 ( .C1(n5300), .C2(n6698), .A(n5281), .B(n5280), .ZN(n5282)
         );
  INV_X1 U6480 ( .A(n5282), .ZN(U2817) );
  AOI22_X1 U6481 ( .A1(EBX_REG_14__SCAN_IN), .A2(n6695), .B1(
        PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n6078), .ZN(n5283) );
  OAI211_X1 U6482 ( .C1(n5760), .C2(n6085), .A(n5283), .B(n6691), .ZN(n5288)
         );
  INV_X1 U6483 ( .A(n6001), .ZN(n5286) );
  AOI21_X1 U6484 ( .B1(n6069), .B2(n5284), .A(REIP_REG_14__SCAN_IN), .ZN(n5285) );
  OAI22_X1 U6485 ( .A1(n5286), .A2(n5285), .B1(n5611), .B2(n6702), .ZN(n5287)
         );
  AOI211_X1 U6486 ( .C1(n5613), .C2(n6698), .A(n5288), .B(n5287), .ZN(n5289)
         );
  INV_X1 U6487 ( .A(n5289), .ZN(U2813) );
  INV_X1 U6488 ( .A(REIP_REG_15__SCAN_IN), .ZN(n6574) );
  INV_X1 U6489 ( .A(n5601), .ZN(n5290) );
  OAI22_X1 U6490 ( .A1(n6085), .A2(n5748), .B1(n6702), .B2(n5290), .ZN(n5294)
         );
  AOI22_X1 U6491 ( .A1(EBX_REG_15__SCAN_IN), .A2(n6695), .B1(
        REIP_REG_15__SCAN_IN), .B2(n6001), .ZN(n5291) );
  OAI211_X1 U6492 ( .C1(n6693), .C2(n5292), .A(n5291), .B(n6691), .ZN(n5293)
         );
  AOI211_X1 U6493 ( .C1(n6002), .C2(n6574), .A(n5294), .B(n5293), .ZN(n5295)
         );
  OAI21_X1 U6494 ( .B1(n5598), .B2(n5995), .A(n5295), .ZN(U2812) );
  NAND2_X1 U6495 ( .A1(n6158), .A2(n6156), .ZN(n5296) );
  XNOR2_X1 U6496 ( .A(n6157), .B(n5296), .ZN(n6213) );
  INV_X1 U6497 ( .A(n6213), .ZN(n5302) );
  AOI22_X1 U6498 ( .A1(n6186), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .B1(n3668), 
        .B2(REIP_REG_10__SCAN_IN), .ZN(n5297) );
  OAI21_X1 U6499 ( .B1(n6195), .B2(n5298), .A(n5297), .ZN(n5299) );
  AOI21_X1 U6500 ( .B1(n5300), .B2(n6165), .A(n5299), .ZN(n5301) );
  OAI21_X1 U6501 ( .B1(n5302), .B2(n6169), .A(n5301), .ZN(U2976) );
  AND2_X1 U6502 ( .A1(n5304), .A2(n5303), .ZN(n5305) );
  OR2_X1 U6503 ( .A1(n5305), .A2(n5314), .ZN(n5899) );
  INV_X1 U6504 ( .A(n5308), .ZN(n5306) );
  NAND2_X1 U6505 ( .A1(n5317), .A2(n5306), .ZN(n5310) );
  OAI21_X1 U6506 ( .B1(n5944), .B2(n5308), .A(n5307), .ZN(n5309) );
  NAND2_X1 U6507 ( .A1(n5310), .A2(n5309), .ZN(n5909) );
  OAI22_X1 U6508 ( .A1(n5909), .A2(n6091), .B1(n5901), .B2(n6096), .ZN(n5311)
         );
  INV_X1 U6509 ( .A(n5311), .ZN(n5312) );
  OAI21_X1 U6510 ( .B1(n5899), .B2(n6092), .A(n5312), .ZN(U2840) );
  OAI21_X1 U6511 ( .B1(n5314), .B2(n5313), .A(n5465), .ZN(n5892) );
  AOI22_X1 U6512 ( .A1(n6104), .A2(DATAI_4_), .B1(n6103), .B2(
        EAX_REG_20__SCAN_IN), .ZN(n5316) );
  NAND2_X1 U6513 ( .A1(n6100), .A2(DATAI_20_), .ZN(n5315) );
  OAI211_X1 U6514 ( .C1(n5892), .C2(n5914), .A(n5316), .B(n5315), .ZN(U2871)
         );
  INV_X1 U6515 ( .A(EBX_REG_20__SCAN_IN), .ZN(n5322) );
  MUX2_X1 U6516 ( .A(n5319), .B(n5318), .S(n5317), .Z(n5321) );
  XNOR2_X1 U6517 ( .A(n5321), .B(n5320), .ZN(n5706) );
  INV_X1 U6518 ( .A(n5706), .ZN(n5891) );
  OAI222_X1 U6519 ( .A1(n6092), .A2(n5892), .B1(n6096), .B2(n5322), .C1(n5891), 
        .C2(n6091), .ZN(U2839) );
  INV_X1 U6520 ( .A(EBX_REG_30__SCAN_IN), .ZN(n5323) );
  OAI222_X1 U6521 ( .A1(n6092), .A2(n5479), .B1(n6091), .B2(n5324), .C1(n5323), 
        .C2(n6096), .ZN(U2829) );
  OAI22_X1 U6522 ( .A1(n5383), .A2(n6091), .B1(n5325), .B2(n6096), .ZN(U2828)
         );
  INV_X1 U6523 ( .A(n5352), .ZN(n5330) );
  NOR2_X1 U6524 ( .A1(n5353), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5329)
         );
  XNOR2_X1 U6525 ( .A(n5392), .B(n5326), .ZN(n5377) );
  OAI21_X1 U6526 ( .B1(n5377), .B2(n6249), .A(n5327), .ZN(n5328) );
  AOI211_X1 U6527 ( .C1(INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n5330), .A(n5329), .B(n5328), .ZN(n5331) );
  OAI21_X1 U6528 ( .B1(n5332), .B2(n5780), .A(n5331), .ZN(U2989) );
  NOR2_X2 U6529 ( .A1(n5334), .A2(n5333), .ZN(n5338) );
  AOI22_X1 U6530 ( .A1(n5336), .A2(EAX_REG_31__SCAN_IN), .B1(n5335), .B2(
        PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n5337) );
  XNOR2_X1 U6531 ( .A(n5338), .B(n5337), .ZN(n5474) );
  AOI21_X1 U6532 ( .B1(n6186), .B2(PHYADDRPOINTER_REG_31__SCAN_IN), .A(n5339), 
        .ZN(n5340) );
  OAI21_X1 U6533 ( .B1(n6195), .B2(n5341), .A(n5340), .ZN(n5342) );
  AOI21_X1 U6534 ( .B1(n5474), .B2(n5593), .A(n5342), .ZN(n5343) );
  OAI21_X1 U6535 ( .B1(n5344), .B2(n6169), .A(n5343), .ZN(U2955) );
  NAND2_X1 U6536 ( .A1(n5345), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5350) );
  INV_X1 U6537 ( .A(n5520), .ZN(n5348) );
  XNOR2_X1 U6538 ( .A(n5351), .B(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5366)
         );
  OAI21_X1 U6539 ( .B1(INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n5735), .A(n5352), 
        .ZN(n5357) );
  NOR3_X1 U6540 ( .A1(n5353), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .A3(n6625), 
        .ZN(n5356) );
  NAND2_X1 U6541 ( .A1(n3668), .A2(REIP_REG_30__SCAN_IN), .ZN(n5360) );
  OAI21_X1 U6542 ( .B1(n5354), .B2(n6249), .A(n5360), .ZN(n5355) );
  AOI211_X1 U6543 ( .C1(INSTADDRPOINTER_REG_30__SCAN_IN), .C2(n5357), .A(n5356), .B(n5355), .ZN(n5358) );
  OAI21_X1 U6544 ( .B1(n5366), .B2(n5780), .A(n5358), .ZN(U2988) );
  NAND2_X1 U6545 ( .A1(n6164), .A2(n5359), .ZN(n5361) );
  OAI211_X1 U6546 ( .C1(n5362), .C2(n5618), .A(n5361), .B(n5360), .ZN(n5363)
         );
  AOI21_X1 U6547 ( .B1(n5364), .B2(n6165), .A(n5363), .ZN(n5365) );
  OAI21_X1 U6548 ( .B1(n5366), .B2(n6169), .A(n5365), .ZN(U2956) );
  AOI22_X1 U6549 ( .A1(n6100), .A2(DATAI_29_), .B1(EAX_REG_29__SCAN_IN), .B2(
        n6103), .ZN(n5369) );
  NAND2_X1 U6550 ( .A1(n6104), .A2(DATAI_13_), .ZN(n5368) );
  OAI211_X1 U6551 ( .C1(n5367), .C2(n5914), .A(n5369), .B(n5368), .ZN(U2862)
         );
  INV_X1 U6552 ( .A(n5377), .ZN(n5374) );
  AOI22_X1 U6553 ( .A1(PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n6078), .B1(n6077), 
        .B2(n5370), .ZN(n5372) );
  NAND2_X1 U6554 ( .A1(n6695), .A2(EBX_REG_29__SCAN_IN), .ZN(n5371) );
  OAI211_X1 U6555 ( .C1(n5397), .C2(n6520), .A(n5372), .B(n5371), .ZN(n5373)
         );
  AOI21_X1 U6556 ( .B1(n5374), .B2(n6697), .A(n5373), .ZN(n5376) );
  OAI211_X1 U6557 ( .C1(n5367), .C2(n5995), .A(n5376), .B(n5375), .ZN(U2798)
         );
  INV_X1 U6558 ( .A(EBX_REG_29__SCAN_IN), .ZN(n6571) );
  OAI222_X1 U6559 ( .A1(n6571), .A2(n6096), .B1(n6091), .B2(n5377), .C1(n5367), 
        .C2(n6092), .ZN(U2830) );
  INV_X1 U6560 ( .A(n5474), .ZN(n5387) );
  AOI22_X1 U6561 ( .A1(n5378), .A2(EBX_REG_31__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n6078), .ZN(n5382) );
  OAI21_X1 U6562 ( .B1(n6520), .B2(REIP_REG_31__SCAN_IN), .A(
        REIP_REG_30__SCAN_IN), .ZN(n5379) );
  OAI211_X1 U6563 ( .C1(REIP_REG_31__SCAN_IN), .C2(REIP_REG_30__SCAN_IN), .A(
        n5380), .B(n5379), .ZN(n5381) );
  OAI211_X1 U6564 ( .C1(n5383), .C2(n6085), .A(n5382), .B(n5381), .ZN(n5384)
         );
  AOI21_X1 U6565 ( .B1(REIP_REG_31__SCAN_IN), .B2(n5385), .A(n5384), .ZN(n5386) );
  OAI21_X1 U6566 ( .B1(n5387), .B2(n5995), .A(n5386), .ZN(U2796) );
  AOI21_X1 U6567 ( .B1(n5391), .B2(n5389), .A(n5390), .ZN(n5510) );
  INV_X1 U6568 ( .A(n5510), .ZN(n5482) );
  AOI21_X1 U6569 ( .B1(n5393), .B2(n5445), .A(n5392), .ZN(n5640) );
  INV_X1 U6570 ( .A(REIP_REG_28__SCAN_IN), .ZN(n6516) );
  OAI22_X1 U6571 ( .A1(n5394), .A2(n6693), .B1(n6702), .B2(n5508), .ZN(n5395)
         );
  AOI21_X1 U6572 ( .B1(EBX_REG_28__SCAN_IN), .B2(n6695), .A(n5395), .ZN(n5396)
         );
  OAI21_X1 U6573 ( .B1(n5397), .B2(n6516), .A(n5396), .ZN(n5399) );
  INV_X1 U6574 ( .A(REIP_REG_27__SCAN_IN), .ZN(n6513) );
  NOR3_X1 U6575 ( .A1(n5852), .A2(REIP_REG_28__SCAN_IN), .A3(n6513), .ZN(n5398) );
  AOI211_X1 U6576 ( .C1(n6697), .C2(n5640), .A(n5399), .B(n5398), .ZN(n5400)
         );
  OAI21_X1 U6577 ( .B1(n5482), .B2(n5995), .A(n5400), .ZN(U2799) );
  AOI21_X1 U6578 ( .B1(n5402), .B2(n5411), .A(n5443), .ZN(n5526) );
  INV_X1 U6579 ( .A(n5526), .ZN(n5488) );
  NAND2_X1 U6580 ( .A1(REIP_REG_24__SCAN_IN), .A2(n5418), .ZN(n5414) );
  OAI21_X1 U6581 ( .B1(n6508), .B2(n5414), .A(n6511), .ZN(n5409) );
  OR2_X1 U6582 ( .A1(n5417), .A2(n5404), .ZN(n5405) );
  NAND2_X1 U6583 ( .A1(n5447), .A2(n5405), .ZN(n5655) );
  OAI22_X1 U6584 ( .A1(n6043), .A2(n6732), .B1(n5524), .B2(n6693), .ZN(n5406)
         );
  AOI21_X1 U6585 ( .B1(n6077), .B2(n5522), .A(n5406), .ZN(n5407) );
  OAI21_X1 U6586 ( .B1(n5655), .B2(n6085), .A(n5407), .ZN(n5408) );
  AOI21_X1 U6587 ( .B1(n5409), .B2(n5847), .A(n5408), .ZN(n5410) );
  OAI21_X1 U6588 ( .B1(n5488), .B2(n5995), .A(n5410), .ZN(U2801) );
  INV_X1 U6589 ( .A(n5411), .ZN(n5412) );
  AOI21_X1 U6590 ( .B1(n5413), .B2(n5453), .A(n5412), .ZN(n5535) );
  OAI22_X1 U6591 ( .A1(REIP_REG_25__SCAN_IN), .A2(n5414), .B1(n5533), .B2(
        n6702), .ZN(n5423) );
  NOR2_X1 U6592 ( .A1(n5456), .A2(n5415), .ZN(n5416) );
  OR2_X1 U6593 ( .A1(n5417), .A2(n5416), .ZN(n5663) );
  AOI22_X1 U6594 ( .A1(n6695), .A2(EBX_REG_25__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n6078), .ZN(n5421) );
  INV_X1 U6595 ( .A(n5871), .ZN(n5419) );
  AND2_X1 U6596 ( .A1(n6506), .A2(n5418), .ZN(n5859) );
  OAI21_X1 U6597 ( .B1(n5419), .B2(n5859), .A(REIP_REG_25__SCAN_IN), .ZN(n5420) );
  OAI211_X1 U6598 ( .C1(n5663), .C2(n6085), .A(n5421), .B(n5420), .ZN(n5422)
         );
  AOI211_X1 U6599 ( .C1(n5535), .C2(n6698), .A(n5423), .B(n5422), .ZN(n5424)
         );
  INV_X1 U6600 ( .A(n5424), .ZN(U2802) );
  NOR2_X1 U6601 ( .A1(n5426), .A2(n5425), .ZN(n5427) );
  AND2_X1 U6602 ( .A1(n5428), .A2(n5427), .ZN(n5498) );
  OAI21_X1 U6603 ( .B1(n5498), .B2(n5429), .A(n4663), .ZN(n5633) );
  INV_X1 U6604 ( .A(n5629), .ZN(n5439) );
  INV_X1 U6605 ( .A(EBX_REG_12__SCAN_IN), .ZN(n5471) );
  OR2_X1 U6606 ( .A1(n6015), .A2(n5430), .ZN(n5431) );
  NAND2_X1 U6607 ( .A1(n5432), .A2(n5431), .ZN(n5774) );
  OAI22_X1 U6608 ( .A1(n5471), .A2(n6043), .B1(n6085), .B2(n5774), .ZN(n5433)
         );
  INV_X1 U6609 ( .A(n5433), .ZN(n5436) );
  AOI211_X1 U6610 ( .C1(REIP_REG_12__SCAN_IN), .C2(n6016), .A(n6045), .B(n5434), .ZN(n5435) );
  OAI211_X1 U6611 ( .C1(n5437), .C2(n6693), .A(n5436), .B(n5435), .ZN(n5438)
         );
  AOI21_X1 U6612 ( .B1(n6077), .B2(n5439), .A(n5438), .ZN(n5440) );
  OAI21_X1 U6613 ( .B1(n5633), .B2(n5995), .A(n5440), .ZN(U2815) );
  AOI22_X1 U6614 ( .A1(n5640), .A2(n6087), .B1(n5462), .B2(EBX_REG_28__SCAN_IN), .ZN(n5441) );
  OAI21_X1 U6615 ( .B1(n5482), .B2(n6092), .A(n5441), .ZN(U2831) );
  OR2_X1 U6616 ( .A1(n5443), .A2(n5442), .ZN(n5444) );
  AND2_X1 U6617 ( .A1(n5389), .A2(n5444), .ZN(n5849) );
  INV_X1 U6618 ( .A(n5849), .ZN(n5485) );
  INV_X1 U6619 ( .A(n5445), .ZN(n5446) );
  AOI21_X1 U6620 ( .B1(n5448), .B2(n5447), .A(n5446), .ZN(n5848) );
  AOI22_X1 U6621 ( .A1(n5848), .A2(n6087), .B1(EBX_REG_27__SCAN_IN), .B2(n5462), .ZN(n5449) );
  OAI21_X1 U6622 ( .B1(n5485), .B2(n6092), .A(n5449), .ZN(U2832) );
  OAI22_X1 U6623 ( .A1(n5655), .A2(n6091), .B1(n6732), .B2(n6096), .ZN(n5450)
         );
  INV_X1 U6624 ( .A(n5450), .ZN(n5451) );
  OAI21_X1 U6625 ( .B1(n5488), .B2(n6092), .A(n5451), .ZN(U2833) );
  INV_X1 U6626 ( .A(n5535), .ZN(n5491) );
  INV_X1 U6627 ( .A(EBX_REG_25__SCAN_IN), .ZN(n5452) );
  OAI222_X1 U6628 ( .A1(n6092), .A2(n5491), .B1(n6096), .B2(n5452), .C1(n5663), 
        .C2(n6091), .ZN(U2834) );
  OAI21_X1 U6629 ( .B1(n5553), .B2(n5454), .A(n5453), .ZN(n5543) );
  AND2_X1 U6630 ( .A1(n5680), .A2(n5455), .ZN(n5457) );
  OR2_X1 U6631 ( .A1(n5457), .A2(n5456), .ZN(n5862) );
  OAI22_X1 U6632 ( .A1(n5862), .A2(n6091), .B1(n5458), .B2(n6096), .ZN(n5459)
         );
  INV_X1 U6633 ( .A(n5459), .ZN(n5460) );
  OAI21_X1 U6634 ( .B1(n5543), .B2(n6092), .A(n5460), .ZN(U2835) );
  XNOR2_X1 U6635 ( .A(n5679), .B(n5675), .ZN(n5875) );
  AOI22_X1 U6636 ( .A1(n5875), .A2(n6087), .B1(EBX_REG_22__SCAN_IN), .B2(n5462), .ZN(n5463) );
  OAI21_X1 U6637 ( .B1(n5874), .B2(n6092), .A(n5463), .ZN(U2837) );
  AOI21_X1 U6638 ( .B1(n5466), .B2(n5465), .A(n3992), .ZN(n5921) );
  INV_X1 U6639 ( .A(n5921), .ZN(n5470) );
  INV_X1 U6640 ( .A(EBX_REG_21__SCAN_IN), .ZN(n5469) );
  OAI21_X1 U6641 ( .B1(n5468), .B2(n5467), .A(n5679), .ZN(n5883) );
  OAI222_X1 U6642 ( .A1(n6092), .A2(n5470), .B1(n6096), .B2(n5469), .C1(n5883), 
        .C2(n6091), .ZN(U2838) );
  OAI222_X1 U6643 ( .A1(n5774), .A2(n6091), .B1(n6096), .B2(n5471), .C1(n6092), 
        .C2(n5633), .ZN(U2847) );
  NAND3_X1 U6644 ( .A1(n5474), .A2(n5473), .A3(n5472), .ZN(n5476) );
  AOI22_X1 U6645 ( .A1(n6100), .A2(DATAI_31_), .B1(EAX_REG_31__SCAN_IN), .B2(
        n6103), .ZN(n5475) );
  NAND2_X1 U6646 ( .A1(n5476), .A2(n5475), .ZN(U2860) );
  AOI22_X1 U6647 ( .A1(n6100), .A2(DATAI_30_), .B1(EAX_REG_30__SCAN_IN), .B2(
        n6103), .ZN(n5478) );
  NAND2_X1 U6648 ( .A1(n6104), .A2(DATAI_14_), .ZN(n5477) );
  OAI211_X1 U6649 ( .C1(n5479), .C2(n5914), .A(n5478), .B(n5477), .ZN(U2861)
         );
  AOI22_X1 U6650 ( .A1(n6100), .A2(DATAI_28_), .B1(EAX_REG_28__SCAN_IN), .B2(
        n6103), .ZN(n5481) );
  NAND2_X1 U6651 ( .A1(n6104), .A2(DATAI_12_), .ZN(n5480) );
  OAI211_X1 U6652 ( .C1(n5482), .C2(n5914), .A(n5481), .B(n5480), .ZN(U2863)
         );
  AOI22_X1 U6653 ( .A1(n6104), .A2(DATAI_11_), .B1(n6103), .B2(
        EAX_REG_27__SCAN_IN), .ZN(n5484) );
  NAND2_X1 U6654 ( .A1(n6100), .A2(DATAI_27_), .ZN(n5483) );
  OAI211_X1 U6655 ( .C1(n5485), .C2(n5914), .A(n5484), .B(n5483), .ZN(U2864)
         );
  AOI22_X1 U6656 ( .A1(n6100), .A2(DATAI_26_), .B1(EAX_REG_26__SCAN_IN), .B2(
        n6103), .ZN(n5487) );
  NAND2_X1 U6657 ( .A1(n6104), .A2(DATAI_10_), .ZN(n5486) );
  OAI211_X1 U6658 ( .C1(n5488), .C2(n5914), .A(n5487), .B(n5486), .ZN(U2865)
         );
  AOI22_X1 U6659 ( .A1(n6100), .A2(DATAI_25_), .B1(EAX_REG_25__SCAN_IN), .B2(
        n6103), .ZN(n5490) );
  NAND2_X1 U6660 ( .A1(n6104), .A2(DATAI_9_), .ZN(n5489) );
  OAI211_X1 U6661 ( .C1(n5491), .C2(n5914), .A(n5490), .B(n5489), .ZN(U2866)
         );
  AOI22_X1 U6662 ( .A1(n6104), .A2(DATAI_8_), .B1(n6103), .B2(
        EAX_REG_24__SCAN_IN), .ZN(n5493) );
  NAND2_X1 U6663 ( .A1(n6100), .A2(DATAI_24_), .ZN(n5492) );
  OAI211_X1 U6664 ( .C1(n5543), .C2(n5914), .A(n5493), .B(n5492), .ZN(U2867)
         );
  AOI22_X1 U6665 ( .A1(n5499), .A2(DATAI_12_), .B1(n6103), .B2(
        EAX_REG_12__SCAN_IN), .ZN(n5494) );
  OAI21_X1 U6666 ( .B1(n5633), .B2(n5914), .A(n5494), .ZN(U2879) );
  NOR2_X1 U6667 ( .A1(n5496), .A2(n5495), .ZN(n5497) );
  OR2_X1 U6668 ( .A1(n5498), .A2(n5497), .ZN(n6093) );
  AOI22_X1 U6669 ( .A1(n5499), .A2(DATAI_11_), .B1(n6103), .B2(
        EAX_REG_11__SCAN_IN), .ZN(n5500) );
  OAI21_X1 U6670 ( .B1(n6093), .B2(n5914), .A(n5500), .ZN(U2880) );
  NAND2_X1 U6671 ( .A1(n5513), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5504) );
  INV_X1 U6672 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5502) );
  XNOR2_X1 U6673 ( .A(n5506), .B(n5505), .ZN(n5643) );
  NOR2_X1 U6674 ( .A1(n6248), .A2(n6516), .ZN(n5639) );
  AOI21_X1 U6675 ( .B1(n6186), .B2(PHYADDRPOINTER_REG_28__SCAN_IN), .A(n5639), 
        .ZN(n5507) );
  OAI21_X1 U6676 ( .B1(n6195), .B2(n5508), .A(n5507), .ZN(n5509) );
  AOI21_X1 U6677 ( .B1(n5510), .B2(n6165), .A(n5509), .ZN(n5511) );
  OAI21_X1 U6678 ( .B1(n5643), .B2(n6169), .A(n5511), .ZN(U2958) );
  NAND2_X1 U6679 ( .A1(n5513), .A2(n5512), .ZN(n5514) );
  XNOR2_X1 U6680 ( .A(n5514), .B(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5650)
         );
  NOR2_X1 U6681 ( .A1(n6248), .A2(n6513), .ZN(n5644) );
  AOI21_X1 U6682 ( .B1(n6186), .B2(PHYADDRPOINTER_REG_27__SCAN_IN), .A(n5644), 
        .ZN(n5515) );
  OAI21_X1 U6683 ( .B1(n6195), .B2(n5845), .A(n5515), .ZN(n5516) );
  AOI21_X1 U6684 ( .B1(n5849), .B2(n5593), .A(n5516), .ZN(n5517) );
  OAI21_X1 U6685 ( .B1(n5650), .B2(n6169), .A(n5517), .ZN(U2959) );
  NOR2_X1 U6686 ( .A1(n5519), .A2(n5518), .ZN(n5521) );
  XOR2_X1 U6687 ( .A(n5521), .B(n5520), .Z(n5658) );
  NAND2_X1 U6688 ( .A1(n6164), .A2(n5522), .ZN(n5523) );
  NAND2_X1 U6689 ( .A1(n3668), .A2(REIP_REG_26__SCAN_IN), .ZN(n5653) );
  OAI211_X1 U6690 ( .C1(n5618), .C2(n5524), .A(n5523), .B(n5653), .ZN(n5525)
         );
  AOI21_X1 U6691 ( .B1(n5526), .B2(n5593), .A(n5525), .ZN(n5527) );
  OAI21_X1 U6692 ( .B1(n5658), .B2(n6169), .A(n5527), .ZN(U2960) );
  AOI21_X1 U6693 ( .B1(n5530), .B2(n5529), .A(n5528), .ZN(n5666) );
  NAND2_X1 U6694 ( .A1(n3668), .A2(REIP_REG_25__SCAN_IN), .ZN(n5661) );
  INV_X1 U6695 ( .A(n5661), .ZN(n5531) );
  AOI21_X1 U6696 ( .B1(n6186), .B2(PHYADDRPOINTER_REG_25__SCAN_IN), .A(n5531), 
        .ZN(n5532) );
  OAI21_X1 U6697 ( .B1(n6195), .B2(n5533), .A(n5532), .ZN(n5534) );
  AOI21_X1 U6698 ( .B1(n5535), .B2(n6165), .A(n5534), .ZN(n5536) );
  OAI21_X1 U6699 ( .B1(n5666), .B2(n6169), .A(n5536), .ZN(U2961) );
  NAND2_X1 U6700 ( .A1(n5557), .A2(n5537), .ZN(n5547) );
  NAND3_X1 U6701 ( .A1(n2963), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5538) );
  OAI22_X1 U6702 ( .A1(n5547), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .B1(n5539), .B2(n5538), .ZN(n5540) );
  XNOR2_X1 U6703 ( .A(n5540), .B(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5674)
         );
  NOR2_X1 U6704 ( .A1(n6248), .A2(n6506), .ZN(n5667) );
  NOR2_X1 U6705 ( .A1(n5618), .A2(n5541), .ZN(n5542) );
  AOI211_X1 U6706 ( .C1(n6164), .C2(n5853), .A(n5667), .B(n5542), .ZN(n5545)
         );
  INV_X1 U6707 ( .A(n5543), .ZN(n5857) );
  NAND2_X1 U6708 ( .A1(n5857), .A2(n6165), .ZN(n5544) );
  OAI211_X1 U6709 ( .C1(n5674), .C2(n6169), .A(n5545), .B(n5544), .ZN(U2962)
         );
  INV_X1 U6710 ( .A(n5683), .ZN(n5546) );
  NAND3_X1 U6711 ( .A1(n2963), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .A3(n5546), .ZN(n5548) );
  OAI21_X1 U6712 ( .B1(n5549), .B2(n5548), .A(n5547), .ZN(n5550) );
  XNOR2_X1 U6713 ( .A(n5550), .B(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5688)
         );
  NOR2_X1 U6714 ( .A1(n4061), .A2(n5551), .ZN(n5552) );
  OR2_X1 U6715 ( .A1(n5553), .A2(n5552), .ZN(n5911) );
  INV_X1 U6716 ( .A(n5911), .ZN(n5915) );
  NAND2_X1 U6717 ( .A1(n3668), .A2(REIP_REG_23__SCAN_IN), .ZN(n5682) );
  NAND2_X1 U6718 ( .A1(n6186), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5554)
         );
  OAI211_X1 U6719 ( .C1(n6195), .C2(n5864), .A(n5682), .B(n5554), .ZN(n5555)
         );
  AOI21_X1 U6720 ( .B1(n5915), .B2(n5593), .A(n5555), .ZN(n5556) );
  OAI21_X1 U6721 ( .B1(n5688), .B2(n6169), .A(n5556), .ZN(U2963) );
  AOI21_X1 U6722 ( .B1(n5559), .B2(n5558), .A(n5557), .ZN(n5703) );
  NAND2_X1 U6723 ( .A1(n3668), .A2(REIP_REG_21__SCAN_IN), .ZN(n5697) );
  NAND2_X1 U6724 ( .A1(n6186), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n5560)
         );
  OAI211_X1 U6725 ( .C1(n6195), .C2(n5881), .A(n5697), .B(n5560), .ZN(n5561)
         );
  AOI21_X1 U6726 ( .B1(n5921), .B2(n5593), .A(n5561), .ZN(n5562) );
  OAI21_X1 U6727 ( .B1(n5703), .B2(n6169), .A(n5562), .ZN(U2965) );
  XNOR2_X1 U6728 ( .A(n6160), .B(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5563)
         );
  XNOR2_X1 U6729 ( .A(n5564), .B(n5563), .ZN(n5715) );
  AND2_X1 U6730 ( .A1(n3668), .A2(REIP_REG_20__SCAN_IN), .ZN(n5705) );
  NOR2_X1 U6731 ( .A1(n5618), .A2(n5898), .ZN(n5565) );
  AOI211_X1 U6732 ( .C1(n6164), .C2(n5890), .A(n5705), .B(n5565), .ZN(n5568)
         );
  INV_X1 U6733 ( .A(n5892), .ZN(n5566) );
  NAND2_X1 U6734 ( .A1(n5566), .A2(n6165), .ZN(n5567) );
  OAI211_X1 U6735 ( .C1(n5715), .C2(n6169), .A(n5568), .B(n5567), .ZN(U2966)
         );
  XNOR2_X1 U6736 ( .A(n6160), .B(n6641), .ZN(n5569) );
  XNOR2_X1 U6737 ( .A(n5570), .B(n5569), .ZN(n5716) );
  NAND2_X1 U6738 ( .A1(n5716), .A2(n6191), .ZN(n5573) );
  NOR2_X1 U6739 ( .A1(n6248), .A2(n6501), .ZN(n5717) );
  NOR2_X1 U6740 ( .A1(n6195), .A2(n5900), .ZN(n5571) );
  AOI211_X1 U6741 ( .C1(n6186), .C2(PHYADDRPOINTER_REG_19__SCAN_IN), .A(n5717), 
        .B(n5571), .ZN(n5572) );
  OAI211_X1 U6742 ( .C1(n5634), .C2(n5899), .A(n5573), .B(n5572), .ZN(U2967)
         );
  NAND3_X1 U6743 ( .A1(n5931), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .A3(n2963), .ZN(n5927) );
  OR2_X1 U6744 ( .A1(n5628), .A2(n5576), .ZN(n5578) );
  NOR2_X1 U6745 ( .A1(n2963), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5928)
         );
  NAND3_X1 U6746 ( .A1(n5595), .A2(n5928), .A3(n5579), .ZN(n5932) );
  NAND2_X1 U6747 ( .A1(n5927), .A2(n5932), .ZN(n5580) );
  XNOR2_X1 U6748 ( .A(n5580), .B(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5731)
         );
  NAND2_X1 U6749 ( .A1(n3668), .A2(REIP_REG_18__SCAN_IN), .ZN(n5725) );
  OAI21_X1 U6750 ( .B1(n5618), .B2(n5581), .A(n5725), .ZN(n5583) );
  NOR2_X1 U6751 ( .A1(n5996), .A2(n5634), .ZN(n5582) );
  AOI211_X1 U6752 ( .C1(n6164), .C2(n5998), .A(n5583), .B(n5582), .ZN(n5584)
         );
  OAI21_X1 U6753 ( .B1(n5731), .B2(n6169), .A(n5584), .ZN(U2968) );
  MUX2_X1 U6754 ( .A(n5579), .B(INSTADDRPOINTER_REG_16__SCAN_IN), .S(n2963), 
        .Z(n5589) );
  INV_X1 U6755 ( .A(n5589), .ZN(n5588) );
  NAND2_X1 U6756 ( .A1(n5586), .A2(n5585), .ZN(n5587) );
  MUX2_X1 U6757 ( .A(n5589), .B(n5588), .S(n5587), .Z(n5742) );
  INV_X1 U6758 ( .A(n5590), .ZN(n6102) );
  NAND2_X1 U6759 ( .A1(n3668), .A2(REIP_REG_16__SCAN_IN), .ZN(n5736) );
  NAND2_X1 U6760 ( .A1(n6186), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n5591)
         );
  OAI211_X1 U6761 ( .C1(n6195), .C2(n6007), .A(n5736), .B(n5591), .ZN(n5592)
         );
  AOI21_X1 U6762 ( .B1(n6102), .B2(n5593), .A(n5592), .ZN(n5594) );
  OAI21_X1 U6763 ( .B1(n5742), .B2(n6169), .A(n5594), .ZN(U2970) );
  AOI21_X1 U6764 ( .B1(n5597), .B2(n5596), .A(n5595), .ZN(n5752) );
  NAND2_X1 U6765 ( .A1(n3668), .A2(REIP_REG_15__SCAN_IN), .ZN(n5746) );
  OAI21_X1 U6766 ( .B1(n5618), .B2(n5292), .A(n5746), .ZN(n5600) );
  NOR2_X1 U6767 ( .A1(n5598), .A2(n5634), .ZN(n5599) );
  AOI211_X1 U6768 ( .C1(n6164), .C2(n5601), .A(n5600), .B(n5599), .ZN(n5602)
         );
  OAI21_X1 U6769 ( .B1(n5752), .B2(n6169), .A(n5602), .ZN(U2971) );
  OR2_X1 U6770 ( .A1(n5628), .A2(n5624), .ZN(n5615) );
  NAND2_X1 U6771 ( .A1(n5615), .A2(n5603), .ZN(n5605) );
  AND2_X1 U6772 ( .A1(n5605), .A2(n5604), .ZN(n5608) );
  XNOR2_X1 U6773 ( .A(n6160), .B(n5606), .ZN(n5607) );
  XNOR2_X1 U6774 ( .A(n5608), .B(n5607), .ZN(n5768) );
  INV_X1 U6775 ( .A(REIP_REG_14__SCAN_IN), .ZN(n5609) );
  NOR2_X1 U6776 ( .A1(n6248), .A2(n5609), .ZN(n5764) );
  AOI21_X1 U6777 ( .B1(n6186), .B2(PHYADDRPOINTER_REG_14__SCAN_IN), .A(n5764), 
        .ZN(n5610) );
  OAI21_X1 U6778 ( .B1(n6195), .B2(n5611), .A(n5610), .ZN(n5612) );
  AOI21_X1 U6779 ( .B1(n5613), .B2(n6165), .A(n5612), .ZN(n5614) );
  OAI21_X1 U6780 ( .B1(n5768), .B2(n6169), .A(n5614), .ZN(U2972) );
  NAND2_X1 U6781 ( .A1(n5615), .A2(n5625), .ZN(n5617) );
  XNOR2_X1 U6782 ( .A(n5617), .B(n5616), .ZN(n5956) );
  NAND2_X1 U6783 ( .A1(n5956), .A2(n6191), .ZN(n5622) );
  NAND2_X1 U6784 ( .A1(n3668), .A2(REIP_REG_13__SCAN_IN), .ZN(n5952) );
  OAI21_X1 U6785 ( .B1(n5618), .B2(n5230), .A(n5952), .ZN(n5619) );
  AOI21_X1 U6786 ( .B1(n6164), .B2(n5620), .A(n5619), .ZN(n5621) );
  OAI211_X1 U6787 ( .C1(n5634), .C2(n5623), .A(n5622), .B(n5621), .ZN(U2973)
         );
  INV_X1 U6788 ( .A(n5624), .ZN(n5626) );
  NAND2_X1 U6789 ( .A1(n5626), .A2(n5625), .ZN(n5627) );
  XNOR2_X1 U6790 ( .A(n5628), .B(n5627), .ZN(n5769) );
  NAND2_X1 U6791 ( .A1(n5769), .A2(n6191), .ZN(n5632) );
  NOR2_X1 U6792 ( .A1(n6248), .A2(n6635), .ZN(n5777) );
  NOR2_X1 U6793 ( .A1(n6195), .A2(n5629), .ZN(n5630) );
  AOI211_X1 U6794 ( .C1(n6186), .C2(PHYADDRPOINTER_REG_12__SCAN_IN), .A(n5777), 
        .B(n5630), .ZN(n5631) );
  OAI211_X1 U6795 ( .C1(n5634), .C2(n5633), .A(n5632), .B(n5631), .ZN(U2974)
         );
  INV_X1 U6796 ( .A(n5635), .ZN(n5636) );
  NOR3_X1 U6797 ( .A1(n5646), .A2(n5637), .A3(n5636), .ZN(n5638) );
  AOI211_X1 U6798 ( .C1(n5640), .C2(n6280), .A(n5639), .B(n5638), .ZN(n5642)
         );
  NAND2_X1 U6799 ( .A1(n5648), .A2(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5641) );
  OAI211_X1 U6800 ( .C1(n5643), .C2(n5780), .A(n5642), .B(n5641), .ZN(U2990)
         );
  AOI21_X1 U6801 ( .B1(n5848), .B2(n6280), .A(n5644), .ZN(n5645) );
  OAI21_X1 U6802 ( .B1(INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n5646), .A(n5645), 
        .ZN(n5647) );
  AOI21_X1 U6803 ( .B1(INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n5648), .A(n5647), 
        .ZN(n5649) );
  OAI21_X1 U6804 ( .B1(n5650), .B2(n5780), .A(n5649), .ZN(U2991) );
  INV_X1 U6805 ( .A(n5651), .ZN(n5670) );
  XNOR2_X1 U6806 ( .A(n5659), .B(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5652)
         );
  NAND2_X1 U6807 ( .A1(n5660), .A2(n5652), .ZN(n5654) );
  OAI211_X1 U6808 ( .C1(n6249), .C2(n5655), .A(n5654), .B(n5653), .ZN(n5656)
         );
  AOI21_X1 U6809 ( .B1(INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n5670), .A(n5656), 
        .ZN(n5657) );
  OAI21_X1 U6810 ( .B1(n5658), .B2(n5780), .A(n5657), .ZN(U2992) );
  NAND2_X1 U6811 ( .A1(n5660), .A2(n5659), .ZN(n5662) );
  OAI211_X1 U6812 ( .C1(n6249), .C2(n5663), .A(n5662), .B(n5661), .ZN(n5664)
         );
  AOI21_X1 U6813 ( .B1(INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n5670), .A(n5664), 
        .ZN(n5665) );
  OAI21_X1 U6814 ( .B1(n5666), .B2(n5780), .A(n5665), .ZN(U2993) );
  INV_X1 U6815 ( .A(n5862), .ZN(n5668) );
  AOI21_X1 U6816 ( .B1(n5668), .B2(n6280), .A(n5667), .ZN(n5673) );
  NOR3_X1 U6817 ( .A1(n5698), .A2(n5683), .A3(n5669), .ZN(n5671) );
  OAI21_X1 U6818 ( .B1(INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n5671), .A(n5670), 
        .ZN(n5672) );
  OAI211_X1 U6819 ( .C1(n5674), .C2(n5780), .A(n5673), .B(n5672), .ZN(U2994)
         );
  INV_X1 U6820 ( .A(n5675), .ZN(n5678) );
  INV_X1 U6821 ( .A(n5676), .ZN(n5677) );
  OAI21_X1 U6822 ( .B1(n5679), .B2(n5678), .A(n5677), .ZN(n5681) );
  NAND2_X1 U6823 ( .A1(n5681), .A2(n5680), .ZN(n5910) );
  OAI21_X1 U6824 ( .B1(n5910), .B2(n6249), .A(n5682), .ZN(n5685) );
  NOR3_X1 U6825 ( .A1(n5698), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .A3(n5683), 
        .ZN(n5684) );
  AOI211_X1 U6826 ( .C1(INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n5686), .A(n5685), .B(n5684), .ZN(n5687) );
  OAI21_X1 U6827 ( .B1(n5688), .B2(n5780), .A(n5687), .ZN(U2995) );
  INV_X1 U6828 ( .A(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5695) );
  XNOR2_X1 U6829 ( .A(INSTADDRPOINTER_REG_22__SCAN_IN), .B(
        INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5690) );
  NOR2_X1 U6830 ( .A1(n5698), .A2(n5690), .ZN(n5691) );
  AOI211_X1 U6831 ( .C1(n6280), .C2(n5875), .A(n5692), .B(n5691), .ZN(n5693)
         );
  OAI211_X1 U6832 ( .C1(n5696), .C2(n5695), .A(n5694), .B(n5693), .ZN(U2996)
         );
  INV_X1 U6833 ( .A(n5696), .ZN(n5701) );
  OAI21_X1 U6834 ( .B1(n5883), .B2(n6249), .A(n5697), .ZN(n5700) );
  NOR2_X1 U6835 ( .A1(n5698), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5699)
         );
  AOI211_X1 U6836 ( .C1(INSTADDRPOINTER_REG_21__SCAN_IN), .C2(n5701), .A(n5700), .B(n5699), .ZN(n5702) );
  OAI21_X1 U6837 ( .B1(n5703), .B2(n5780), .A(n5702), .ZN(U2997) );
  NOR3_X1 U6838 ( .A1(n5707), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .A3(n6641), 
        .ZN(n5704) );
  AOI211_X1 U6839 ( .C1(n6280), .C2(n5706), .A(n5705), .B(n5704), .ZN(n5714)
         );
  NOR2_X1 U6840 ( .A1(n5707), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5721)
         );
  OAI21_X1 U6841 ( .B1(n5708), .B2(n5948), .A(n6207), .ZN(n5710) );
  AND2_X1 U6842 ( .A1(n5710), .A2(n5709), .ZN(n5949) );
  OR2_X1 U6843 ( .A1(n6284), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5711)
         );
  NAND2_X1 U6844 ( .A1(n5949), .A2(n5711), .ZN(n5727) );
  INV_X1 U6845 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5728) );
  AND2_X1 U6846 ( .A1(n6210), .A2(n5728), .ZN(n5712) );
  OR2_X1 U6847 ( .A1(n5727), .A2(n5712), .ZN(n5720) );
  OAI21_X1 U6848 ( .B1(n5721), .B2(n5720), .A(INSTADDRPOINTER_REG_20__SCAN_IN), 
        .ZN(n5713) );
  OAI211_X1 U6849 ( .C1(n5715), .C2(n5780), .A(n5714), .B(n5713), .ZN(U2998)
         );
  INV_X1 U6850 ( .A(n5716), .ZN(n5724) );
  INV_X1 U6851 ( .A(n5717), .ZN(n5718) );
  OAI21_X1 U6852 ( .B1(n5909), .B2(n6249), .A(n5718), .ZN(n5719) );
  AOI21_X1 U6853 ( .B1(n5720), .B2(INSTADDRPOINTER_REG_19__SCAN_IN), .A(n5719), 
        .ZN(n5723) );
  INV_X1 U6854 ( .A(n5721), .ZN(n5722) );
  OAI211_X1 U6855 ( .C1(n5724), .C2(n5780), .A(n5723), .B(n5722), .ZN(U2999)
         );
  OAI21_X1 U6856 ( .B1(n6000), .B2(n6249), .A(n5725), .ZN(n5726) );
  AOI21_X1 U6857 ( .B1(n5727), .B2(INSTADDRPOINTER_REG_18__SCAN_IN), .A(n5726), 
        .ZN(n5730) );
  NAND3_X1 U6858 ( .A1(n5940), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .A3(n5728), .ZN(n5729) );
  OAI211_X1 U6859 ( .C1(n5731), .C2(n5780), .A(n5730), .B(n5729), .ZN(U3000)
         );
  AOI211_X1 U6860 ( .C1(n5579), .C2(n5744), .A(n6196), .B(n5743), .ZN(n5740)
         );
  INV_X1 U6861 ( .A(n5743), .ZN(n5734) );
  INV_X1 U6862 ( .A(n5732), .ZN(n5753) );
  AOI22_X1 U6863 ( .A1(n5753), .A2(n6207), .B1(n6206), .B2(n5733), .ZN(n6204)
         );
  OAI21_X1 U6864 ( .B1(n5735), .B2(n5734), .A(n6204), .ZN(n5750) );
  NAND2_X1 U6865 ( .A1(n5750), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5737) );
  OAI211_X1 U6866 ( .C1(n6249), .C2(n6011), .A(n5737), .B(n5736), .ZN(n5738)
         );
  AOI21_X1 U6867 ( .B1(n5740), .B2(n5739), .A(n5738), .ZN(n5741) );
  OAI21_X1 U6868 ( .B1(n5742), .B2(n5780), .A(n5741), .ZN(U3002) );
  NOR2_X1 U6869 ( .A1(n6196), .A2(n5743), .ZN(n5745) );
  NAND2_X1 U6870 ( .A1(n5745), .A2(n5744), .ZN(n5747) );
  OAI211_X1 U6871 ( .C1(n6249), .C2(n5748), .A(n5747), .B(n5746), .ZN(n5749)
         );
  AOI21_X1 U6872 ( .B1(n5750), .B2(INSTADDRPOINTER_REG_15__SCAN_IN), .A(n5749), 
        .ZN(n5751) );
  OAI21_X1 U6873 ( .B1(n5752), .B2(n5780), .A(n5751), .ZN(U3003) );
  AOI21_X1 U6874 ( .B1(n5754), .B2(n5753), .A(INSTADDRPOINTER_REG_13__SCAN_IN), 
        .ZN(n5759) );
  INV_X1 U6875 ( .A(n5755), .ZN(n5951) );
  OR2_X1 U6876 ( .A1(n5951), .A2(n5756), .ZN(n5757) );
  OAI211_X1 U6877 ( .C1(n5761), .C2(n5758), .A(n6204), .B(n5757), .ZN(n5955)
         );
  OAI21_X1 U6878 ( .B1(n5759), .B2(n5955), .A(INSTADDRPOINTER_REG_14__SCAN_IN), 
        .ZN(n5767) );
  INV_X1 U6879 ( .A(n5760), .ZN(n5765) );
  INV_X1 U6880 ( .A(n5761), .ZN(n5762) );
  NOR3_X1 U6881 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n6196), .A3(n5762), 
        .ZN(n5763) );
  AOI211_X1 U6882 ( .C1(n6280), .C2(n5765), .A(n5764), .B(n5763), .ZN(n5766)
         );
  OAI211_X1 U6883 ( .C1(n5768), .C2(n5780), .A(n5767), .B(n5766), .ZN(U3004)
         );
  INV_X1 U6884 ( .A(n5769), .ZN(n5781) );
  OAI21_X1 U6885 ( .B1(n5771), .B2(n5770), .A(n6202), .ZN(n5773) );
  AOI21_X1 U6886 ( .B1(n6204), .B2(n5773), .A(n5772), .ZN(n5778) );
  NOR2_X1 U6887 ( .A1(n6249), .A2(n5774), .ZN(n5776) );
  NOR3_X1 U6888 ( .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n6196), .A3(n6202), 
        .ZN(n5775) );
  NOR4_X1 U6889 ( .A1(n5778), .A2(n5777), .A3(n5776), .A4(n5775), .ZN(n5779)
         );
  OAI21_X1 U6890 ( .B1(n5781), .B2(n5780), .A(n5779), .ZN(U3006) );
  OAI21_X1 U6891 ( .B1(STATEBS16_REG_SCAN_IN), .B2(n5783), .A(n5782), .ZN(
        n5784) );
  OAI21_X1 U6892 ( .B1(n5789), .B2(n5785), .A(n5784), .ZN(n5786) );
  MUX2_X1 U6893 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n5786), .S(n6291), 
        .Z(U3464) );
  XNOR2_X1 U6894 ( .A(n5788), .B(n5787), .ZN(n5792) );
  OAI22_X1 U6895 ( .A1(n5792), .A2(n5791), .B1(n5790), .B2(n5789), .ZN(n5793)
         );
  MUX2_X1 U6896 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n5793), .S(n6291), 
        .Z(U3463) );
  NOR2_X1 U6897 ( .A1(n5794), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n5795)
         );
  AOI22_X1 U6898 ( .A1(n5799), .A2(n5797), .B1(n5796), .B2(n5795), .ZN(n5838)
         );
  NOR2_X1 U6899 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5798), .ZN(n5836)
         );
  INV_X1 U6900 ( .A(n5799), .ZN(n5803) );
  OAI21_X1 U6901 ( .B1(n5801), .B2(n5841), .A(n5800), .ZN(n5802) );
  NAND2_X1 U6902 ( .A1(n5803), .A2(n5802), .ZN(n5805) );
  OAI221_X1 U6903 ( .B1(n5836), .B2(n6717), .C1(n5836), .C2(n5805), .A(n5804), 
        .ZN(n5835) );
  AOI22_X1 U6904 ( .A1(n6375), .A2(n5836), .B1(INSTQUEUE_REG_2__0__SCAN_IN), 
        .B2(n5835), .ZN(n5806) );
  OAI21_X1 U6905 ( .B1(n5807), .B2(n5838), .A(n5806), .ZN(n5808) );
  AOI21_X1 U6906 ( .B1(n5809), .B2(n5841), .A(n5808), .ZN(n5810) );
  OAI21_X1 U6907 ( .B1(n6377), .B2(n5843), .A(n5810), .ZN(U3036) );
  AOI22_X1 U6908 ( .A1(n6383), .A2(n5836), .B1(INSTQUEUE_REG_2__1__SCAN_IN), 
        .B2(n5835), .ZN(n5811) );
  OAI21_X1 U6909 ( .B1(n5812), .B2(n5838), .A(n5811), .ZN(n5813) );
  AOI21_X1 U6910 ( .B1(n6343), .B2(n5841), .A(n5813), .ZN(n5814) );
  OAI21_X1 U6911 ( .B1(n6387), .B2(n5843), .A(n5814), .ZN(U3037) );
  AOI22_X1 U6912 ( .A1(n6325), .A2(n5836), .B1(INSTQUEUE_REG_2__2__SCAN_IN), 
        .B2(n5835), .ZN(n5815) );
  OAI21_X1 U6913 ( .B1(n5816), .B2(n5838), .A(n5815), .ZN(n5817) );
  AOI21_X1 U6914 ( .B1(n6326), .B2(n5841), .A(n5817), .ZN(n5818) );
  OAI21_X1 U6915 ( .B1(n6330), .B2(n5843), .A(n5818), .ZN(U3038) );
  AOI22_X1 U6916 ( .A1(n6346), .A2(n5836), .B1(INSTQUEUE_REG_2__3__SCAN_IN), 
        .B2(n5835), .ZN(n5819) );
  OAI21_X1 U6917 ( .B1(n5820), .B2(n5838), .A(n5819), .ZN(n5821) );
  AOI21_X1 U6918 ( .B1(n6347), .B2(n5841), .A(n5821), .ZN(n5822) );
  OAI21_X1 U6919 ( .B1(n6351), .B2(n5843), .A(n5822), .ZN(U3039) );
  AOI22_X1 U6920 ( .A1(n6296), .A2(n5836), .B1(INSTQUEUE_REG_2__4__SCAN_IN), 
        .B2(n5835), .ZN(n5823) );
  OAI21_X1 U6921 ( .B1(n5824), .B2(n5838), .A(n5823), .ZN(n5825) );
  AOI21_X1 U6922 ( .B1(n6297), .B2(n5841), .A(n5825), .ZN(n5826) );
  OAI21_X1 U6923 ( .B1(n6301), .B2(n5843), .A(n5826), .ZN(U3040) );
  AOI22_X1 U6924 ( .A1(n6352), .A2(n5836), .B1(INSTQUEUE_REG_2__5__SCAN_IN), 
        .B2(n5835), .ZN(n5827) );
  OAI21_X1 U6925 ( .B1(n5828), .B2(n5838), .A(n5827), .ZN(n5829) );
  AOI21_X1 U6926 ( .B1(n6353), .B2(n5841), .A(n5829), .ZN(n5830) );
  OAI21_X1 U6927 ( .B1(n6357), .B2(n5843), .A(n5830), .ZN(U3041) );
  AOI22_X1 U6928 ( .A1(n6358), .A2(n5836), .B1(INSTQUEUE_REG_2__6__SCAN_IN), 
        .B2(n5835), .ZN(n5831) );
  OAI21_X1 U6929 ( .B1(n5832), .B2(n5838), .A(n5831), .ZN(n5833) );
  AOI21_X1 U6930 ( .B1(n6359), .B2(n5841), .A(n5833), .ZN(n5834) );
  OAI21_X1 U6931 ( .B1(n6363), .B2(n5843), .A(n5834), .ZN(U3042) );
  AOI22_X1 U6932 ( .A1(n6365), .A2(n5836), .B1(INSTQUEUE_REG_2__7__SCAN_IN), 
        .B2(n5835), .ZN(n5837) );
  OAI21_X1 U6933 ( .B1(n5839), .B2(n5838), .A(n5837), .ZN(n5840) );
  AOI21_X1 U6934 ( .B1(n6366), .B2(n5841), .A(n5840), .ZN(n5842) );
  OAI21_X1 U6935 ( .B1(n6374), .B2(n5843), .A(n5842), .ZN(U3043) );
  AND2_X1 U6936 ( .A1(n6136), .A2(DATAO_REG_31__SCAN_IN), .ZN(U2892) );
  AOI22_X1 U6937 ( .A1(EBX_REG_27__SCAN_IN), .A2(n6695), .B1(
        PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n6078), .ZN(n5844) );
  OAI21_X1 U6938 ( .B1(n5845), .B2(n6702), .A(n5844), .ZN(n5846) );
  AOI21_X1 U6939 ( .B1(REIP_REG_27__SCAN_IN), .B2(n5847), .A(n5846), .ZN(n5851) );
  AOI22_X1 U6940 ( .A1(n5849), .A2(n6698), .B1(n5848), .B2(n6697), .ZN(n5850)
         );
  OAI211_X1 U6941 ( .C1(REIP_REG_27__SCAN_IN), .C2(n5852), .A(n5851), .B(n5850), .ZN(U2800) );
  AOI22_X1 U6942 ( .A1(PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n6078), .B1(n6077), 
        .B2(n5853), .ZN(n5855) );
  NAND2_X1 U6943 ( .A1(n6695), .A2(EBX_REG_24__SCAN_IN), .ZN(n5854) );
  OAI211_X1 U6944 ( .C1(n5871), .C2(n6506), .A(n5855), .B(n5854), .ZN(n5856)
         );
  AOI21_X1 U6945 ( .B1(n5857), .B2(n6698), .A(n5856), .ZN(n5858) );
  INV_X1 U6946 ( .A(n5858), .ZN(n5860) );
  NOR2_X1 U6947 ( .A1(n5860), .A2(n5859), .ZN(n5861) );
  OAI21_X1 U6948 ( .B1(n5862), .B2(n6085), .A(n5861), .ZN(U2803) );
  INV_X1 U6949 ( .A(REIP_REG_21__SCAN_IN), .ZN(n5863) );
  NOR2_X1 U6950 ( .A1(n5863), .A2(n5876), .ZN(n5872) );
  AOI21_X1 U6951 ( .B1(REIP_REG_22__SCAN_IN), .B2(n5872), .A(
        REIP_REG_23__SCAN_IN), .ZN(n5870) );
  INV_X1 U6952 ( .A(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5865) );
  OAI22_X1 U6953 ( .A1(n5865), .A2(n6693), .B1(n5864), .B2(n6702), .ZN(n5866)
         );
  AOI21_X1 U6954 ( .B1(EBX_REG_23__SCAN_IN), .B2(n6695), .A(n5866), .ZN(n5869)
         );
  OAI22_X1 U6955 ( .A1(n5911), .A2(n5995), .B1(n5910), .B2(n6085), .ZN(n5867)
         );
  INV_X1 U6956 ( .A(n5867), .ZN(n5868) );
  OAI211_X1 U6957 ( .C1(n5871), .C2(n5870), .A(n5869), .B(n5868), .ZN(U2804)
         );
  AOI22_X1 U6958 ( .A1(EBX_REG_22__SCAN_IN), .A2(n6695), .B1(
        PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n6078), .ZN(n5880) );
  AOI22_X1 U6959 ( .A1(n5873), .A2(n6077), .B1(n5872), .B2(n4018), .ZN(n5879)
         );
  INV_X1 U6960 ( .A(n5874), .ZN(n5918) );
  AOI22_X1 U6961 ( .A1(n5918), .A2(n6698), .B1(n6697), .B2(n5875), .ZN(n5878)
         );
  NOR2_X1 U6962 ( .A1(REIP_REG_21__SCAN_IN), .A2(n5876), .ZN(n5885) );
  OAI21_X1 U6963 ( .B1(n5885), .B2(n5895), .A(REIP_REG_22__SCAN_IN), .ZN(n5877) );
  NAND4_X1 U6964 ( .A1(n5880), .A2(n5879), .A3(n5878), .A4(n5877), .ZN(U2805)
         );
  AOI22_X1 U6965 ( .A1(EBX_REG_21__SCAN_IN), .A2(n6695), .B1(
        PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n6078), .ZN(n5889) );
  INV_X1 U6966 ( .A(n5881), .ZN(n5882) );
  AOI22_X1 U6967 ( .A1(n5882), .A2(n6077), .B1(REIP_REG_21__SCAN_IN), .B2(
        n5895), .ZN(n5888) );
  INV_X1 U6968 ( .A(n5883), .ZN(n5884) );
  AOI22_X1 U6969 ( .A1(n5921), .A2(n6698), .B1(n5884), .B2(n6697), .ZN(n5887)
         );
  INV_X1 U6970 ( .A(n5885), .ZN(n5886) );
  NAND4_X1 U6971 ( .A1(n5889), .A2(n5888), .A3(n5887), .A4(n5886), .ZN(U2806)
         );
  AOI22_X1 U6972 ( .A1(EBX_REG_20__SCAN_IN), .A2(n6695), .B1(n5890), .B2(n6077), .ZN(n5897) );
  OAI22_X1 U6973 ( .A1(n5892), .A2(n5995), .B1(n5891), .B2(n6085), .ZN(n5893)
         );
  AOI221_X1 U6974 ( .B1(REIP_REG_20__SCAN_IN), .B2(n5895), .C1(n5894), .C2(
        n5895), .A(n5893), .ZN(n5896) );
  OAI211_X1 U6975 ( .C1(n5898), .C2(n6693), .A(n5897), .B(n5896), .ZN(U2807)
         );
  INV_X1 U6976 ( .A(n5899), .ZN(n5924) );
  NOR3_X1 U6977 ( .A1(REIP_REG_19__SCAN_IN), .A2(n6499), .A3(n5906), .ZN(n5905) );
  OAI22_X1 U6978 ( .A1(n5901), .A2(n6043), .B1(n5900), .B2(n6702), .ZN(n5902)
         );
  AOI211_X1 U6979 ( .C1(n6078), .C2(PHYADDRPOINTER_REG_19__SCAN_IN), .A(n5902), 
        .B(n6045), .ZN(n5903) );
  INV_X1 U6980 ( .A(n5903), .ZN(n5904) );
  AOI211_X1 U6981 ( .C1(n5924), .C2(n6698), .A(n5905), .B(n5904), .ZN(n5908)
         );
  NOR2_X1 U6982 ( .A1(REIP_REG_18__SCAN_IN), .A2(n5906), .ZN(n5992) );
  OAI21_X1 U6983 ( .B1(n5992), .B2(n6688), .A(REIP_REG_19__SCAN_IN), .ZN(n5907) );
  OAI211_X1 U6984 ( .C1(n5909), .C2(n6085), .A(n5908), .B(n5907), .ZN(U2808)
         );
  OAI22_X1 U6985 ( .A1(n5911), .A2(n6092), .B1(n5910), .B2(n6091), .ZN(n5912)
         );
  INV_X1 U6986 ( .A(n5912), .ZN(n5913) );
  OAI21_X1 U6987 ( .B1(n6657), .B2(n6096), .A(n5913), .ZN(U2836) );
  INV_X1 U6988 ( .A(n5914), .ZN(n6101) );
  AOI22_X1 U6989 ( .A1(n5915), .A2(n6101), .B1(n6100), .B2(DATAI_23_), .ZN(
        n5917) );
  AOI22_X1 U6990 ( .A1(n6104), .A2(DATAI_7_), .B1(n6103), .B2(
        EAX_REG_23__SCAN_IN), .ZN(n5916) );
  NAND2_X1 U6991 ( .A1(n5917), .A2(n5916), .ZN(U2868) );
  AOI22_X1 U6992 ( .A1(n5918), .A2(n6101), .B1(n6100), .B2(DATAI_22_), .ZN(
        n5920) );
  AOI22_X1 U6993 ( .A1(n6104), .A2(DATAI_6_), .B1(n6103), .B2(
        EAX_REG_22__SCAN_IN), .ZN(n5919) );
  NAND2_X1 U6994 ( .A1(n5920), .A2(n5919), .ZN(U2869) );
  AOI22_X1 U6995 ( .A1(n5921), .A2(n6101), .B1(n6100), .B2(DATAI_21_), .ZN(
        n5923) );
  AOI22_X1 U6996 ( .A1(n6104), .A2(DATAI_5_), .B1(n6103), .B2(
        EAX_REG_21__SCAN_IN), .ZN(n5922) );
  NAND2_X1 U6997 ( .A1(n5923), .A2(n5922), .ZN(U2870) );
  AOI22_X1 U6998 ( .A1(n5924), .A2(n6101), .B1(n6100), .B2(DATAI_19_), .ZN(
        n5926) );
  AOI22_X1 U6999 ( .A1(n6104), .A2(DATAI_3_), .B1(n6103), .B2(
        EAX_REG_19__SCAN_IN), .ZN(n5925) );
  NAND2_X1 U7000 ( .A1(n5926), .A2(n5925), .ZN(U2872) );
  AOI22_X1 U7001 ( .A1(n3668), .A2(REIP_REG_17__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n6186), .ZN(n5939) );
  INV_X1 U7002 ( .A(n5927), .ZN(n5934) );
  INV_X1 U7003 ( .A(n5928), .ZN(n5930) );
  NAND2_X1 U7004 ( .A1(n2967), .A2(n5579), .ZN(n5929) );
  AOI22_X1 U7005 ( .A1(n5931), .A2(n5930), .B1(INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n5929), .ZN(n5933) );
  OAI21_X1 U7006 ( .B1(n5934), .B2(n5933), .A(n5932), .ZN(n5945) );
  NAND2_X1 U7007 ( .A1(n5067), .A2(n5935), .ZN(n5936) );
  AND2_X1 U7008 ( .A1(n5937), .A2(n5936), .ZN(n6699) );
  AOI22_X1 U7009 ( .A1(n5945), .A2(n6191), .B1(n6165), .B2(n6699), .ZN(n5938)
         );
  OAI211_X1 U7010 ( .C1(n6195), .C2(n6703), .A(n5939), .B(n5938), .ZN(U2969)
         );
  AOI22_X1 U7011 ( .A1(REIP_REG_17__SCAN_IN), .A2(n3668), .B1(n5940), .B2(
        n5948), .ZN(n5947) );
  NAND2_X1 U7012 ( .A1(n5942), .A2(n5941), .ZN(n5943) );
  AND2_X1 U7013 ( .A1(n5944), .A2(n5943), .ZN(n6696) );
  AOI22_X1 U7014 ( .A1(n5945), .A2(n6282), .B1(n6280), .B2(n6696), .ZN(n5946)
         );
  OAI211_X1 U7015 ( .C1(n5949), .C2(n5948), .A(n5947), .B(n5946), .ZN(U3001)
         );
  NAND2_X1 U7016 ( .A1(n5951), .A2(n5950), .ZN(n5959) );
  INV_X1 U7017 ( .A(n5952), .ZN(n5953) );
  AOI21_X1 U7018 ( .B1(n5954), .B2(n6280), .A(n5953), .ZN(n5958) );
  AOI22_X1 U7019 ( .A1(n5956), .A2(n6282), .B1(INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n5955), .ZN(n5957) );
  OAI211_X1 U7020 ( .C1(n6196), .C2(n5959), .A(n5958), .B(n5957), .ZN(U3005)
         );
  INV_X1 U7021 ( .A(n6542), .ZN(n5961) );
  NAND3_X1 U7022 ( .A1(n5962), .A2(n5961), .A3(n5960), .ZN(n5964) );
  OAI22_X1 U7023 ( .A1(n5965), .A2(n5964), .B1(n5963), .B2(n6540), .ZN(U3455)
         );
  INV_X1 U7024 ( .A(STATE_REG_2__SCAN_IN), .ZN(n6716) );
  AOI21_X1 U7025 ( .B1(STATE_REG_1__SCAN_IN), .B2(n6716), .A(n6466), .ZN(n5971) );
  INV_X1 U7026 ( .A(ADS_N_REG_SCAN_IN), .ZN(n5966) );
  NAND2_X1 U7027 ( .A1(n6466), .A2(STATE_REG_1__SCAN_IN), .ZN(n6509) );
  INV_X1 U7028 ( .A(n6509), .ZN(n6485) );
  AOI21_X1 U7029 ( .B1(n5971), .B2(n5966), .A(n6485), .ZN(U2789) );
  NAND2_X1 U7030 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n6560), .ZN(n5969) );
  OAI21_X1 U7031 ( .B1(n5967), .B2(n6447), .A(CODEFETCH_REG_SCAN_IN), .ZN(
        n5968) );
  OAI21_X1 U7032 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n5969), .A(n5968), .ZN(
        U2790) );
  INV_X1 U7033 ( .A(n6485), .ZN(n6565) );
  NOR2_X1 U7034 ( .A1(STATE_REG_0__SCAN_IN), .A2(STATE_REG_2__SCAN_IN), .ZN(
        n5972) );
  OAI21_X1 U7035 ( .B1(D_C_N_REG_SCAN_IN), .B2(n5972), .A(n6565), .ZN(n5970)
         );
  OAI21_X1 U7036 ( .B1(CODEFETCH_REG_SCAN_IN), .B2(n6565), .A(n5970), .ZN(
        U2791) );
  NOR2_X1 U7037 ( .A1(n6485), .A2(n5971), .ZN(n6528) );
  OAI21_X1 U7038 ( .B1(n5972), .B2(BS16_N), .A(n6528), .ZN(n6526) );
  OAI21_X1 U7039 ( .B1(n6528), .B2(n5973), .A(n6526), .ZN(U2792) );
  OAI21_X1 U7040 ( .B1(n5974), .B2(n6647), .A(n6169), .ZN(U2793) );
  NOR4_X1 U7041 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(
        DATAWIDTH_REG_21__SCAN_IN), .A3(DATAWIDTH_REG_22__SCAN_IN), .A4(
        DATAWIDTH_REG_23__SCAN_IN), .ZN(n5978) );
  NOR4_X1 U7042 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(
        DATAWIDTH_REG_17__SCAN_IN), .A3(DATAWIDTH_REG_18__SCAN_IN), .A4(
        DATAWIDTH_REG_19__SCAN_IN), .ZN(n5977) );
  NOR4_X1 U7043 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(
        DATAWIDTH_REG_29__SCAN_IN), .A3(DATAWIDTH_REG_30__SCAN_IN), .A4(
        DATAWIDTH_REG_31__SCAN_IN), .ZN(n5976) );
  NOR4_X1 U7044 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(
        DATAWIDTH_REG_25__SCAN_IN), .A3(DATAWIDTH_REG_26__SCAN_IN), .A4(
        DATAWIDTH_REG_27__SCAN_IN), .ZN(n5975) );
  NAND4_X1 U7045 ( .A1(n5978), .A2(n5977), .A3(n5976), .A4(n5975), .ZN(n5984)
         );
  NOR4_X1 U7046 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(DATAWIDTH_REG_3__SCAN_IN), 
        .A3(DATAWIDTH_REG_4__SCAN_IN), .A4(DATAWIDTH_REG_6__SCAN_IN), .ZN(
        n5982) );
  AOI211_X1 U7047 ( .C1(DATAWIDTH_REG_1__SCAN_IN), .C2(
        DATAWIDTH_REG_0__SCAN_IN), .A(DATAWIDTH_REG_5__SCAN_IN), .B(
        DATAWIDTH_REG_15__SCAN_IN), .ZN(n5981) );
  NOR4_X1 U7048 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(
        DATAWIDTH_REG_12__SCAN_IN), .A3(DATAWIDTH_REG_13__SCAN_IN), .A4(
        DATAWIDTH_REG_14__SCAN_IN), .ZN(n5980) );
  NOR4_X1 U7049 ( .A1(DATAWIDTH_REG_7__SCAN_IN), .A2(DATAWIDTH_REG_8__SCAN_IN), 
        .A3(DATAWIDTH_REG_9__SCAN_IN), .A4(DATAWIDTH_REG_10__SCAN_IN), .ZN(
        n5979) );
  NAND4_X1 U7050 ( .A1(n5982), .A2(n5981), .A3(n5980), .A4(n5979), .ZN(n5983)
         );
  NOR2_X1 U7051 ( .A1(n5984), .A2(n5983), .ZN(n6547) );
  INV_X1 U7052 ( .A(BYTEENABLE_REG_1__SCAN_IN), .ZN(n5986) );
  NOR3_X1 U7053 ( .A1(REIP_REG_0__SCAN_IN), .A2(DATAWIDTH_REG_1__SCAN_IN), 
        .A3(DATAWIDTH_REG_0__SCAN_IN), .ZN(n5987) );
  OAI21_X1 U7054 ( .B1(REIP_REG_1__SCAN_IN), .B2(n5987), .A(n6547), .ZN(n5985)
         );
  OAI21_X1 U7055 ( .B1(n6547), .B2(n5986), .A(n5985), .ZN(U2794) );
  INV_X1 U7056 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6527) );
  AOI21_X1 U7057 ( .B1(n6573), .B2(n6527), .A(n5987), .ZN(n5989) );
  INV_X1 U7058 ( .A(BYTEENABLE_REG_3__SCAN_IN), .ZN(n5988) );
  INV_X1 U7059 ( .A(n6547), .ZN(n6550) );
  AOI22_X1 U7060 ( .A1(n6547), .A2(n5989), .B1(n5988), .B2(n6550), .ZN(U2795)
         );
  AOI21_X1 U7061 ( .B1(n6078), .B2(PHYADDRPOINTER_REG_18__SCAN_IN), .A(n6045), 
        .ZN(n5990) );
  OAI21_X1 U7062 ( .B1(n6043), .B2(n5991), .A(n5990), .ZN(n5993) );
  AOI211_X1 U7063 ( .C1(REIP_REG_18__SCAN_IN), .C2(n6688), .A(n5993), .B(n5992), .ZN(n5994) );
  OAI21_X1 U7064 ( .B1(n5996), .B2(n5995), .A(n5994), .ZN(n5997) );
  AOI21_X1 U7065 ( .B1(n5998), .B2(n6077), .A(n5997), .ZN(n5999) );
  OAI21_X1 U7066 ( .B1(n6085), .B2(n6000), .A(n5999), .ZN(U2809) );
  AOI21_X1 U7067 ( .B1(n6002), .B2(n6574), .A(n6001), .ZN(n6004) );
  AOI21_X1 U7068 ( .B1(n6078), .B2(PHYADDRPOINTER_REG_16__SCAN_IN), .A(n6045), 
        .ZN(n6003) );
  OAI221_X1 U7069 ( .B1(REIP_REG_16__SCAN_IN), .B2(n6005), .C1(n6496), .C2(
        n6004), .A(n6003), .ZN(n6006) );
  AOI21_X1 U7070 ( .B1(EBX_REG_16__SCAN_IN), .B2(n6695), .A(n6006), .ZN(n6010)
         );
  INV_X1 U7071 ( .A(n6007), .ZN(n6008) );
  AOI22_X1 U7072 ( .A1(n6102), .A2(n6698), .B1(n6008), .B2(n6077), .ZN(n6009)
         );
  OAI211_X1 U7073 ( .C1(n6085), .C2(n6011), .A(n6010), .B(n6009), .ZN(U2811)
         );
  AOI22_X1 U7074 ( .A1(EBX_REG_11__SCAN_IN), .A2(n6695), .B1(
        PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n6078), .ZN(n6025) );
  NOR2_X1 U7075 ( .A1(n6013), .A2(n6012), .ZN(n6014) );
  OR2_X1 U7076 ( .A1(n6015), .A2(n6014), .ZN(n6197) );
  INV_X1 U7077 ( .A(n6197), .ZN(n6022) );
  INV_X1 U7078 ( .A(n6016), .ZN(n6020) );
  OR3_X1 U7079 ( .A1(n6018), .A2(REIP_REG_11__SCAN_IN), .A3(n6017), .ZN(n6019)
         );
  OAI21_X1 U7080 ( .B1(n6020), .B2(n6488), .A(n6019), .ZN(n6021) );
  AOI21_X1 U7081 ( .B1(n6697), .B2(n6022), .A(n6021), .ZN(n6024) );
  INV_X1 U7082 ( .A(n6093), .ZN(n6166) );
  AOI22_X1 U7083 ( .A1(n6166), .A2(n6698), .B1(n6077), .B2(n6163), .ZN(n6023)
         );
  NAND4_X1 U7084 ( .A1(n6025), .A2(n6024), .A3(n6023), .A4(n6691), .ZN(U2816)
         );
  AOI22_X1 U7085 ( .A1(EBX_REG_9__SCAN_IN), .A2(n6695), .B1(n6027), .B2(n6026), 
        .ZN(n6035) );
  AOI22_X1 U7086 ( .A1(PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n6078), .B1(
        REIP_REG_9__SCAN_IN), .B2(n6028), .ZN(n6034) );
  AOI21_X1 U7087 ( .B1(n6697), .B2(n6220), .A(n6045), .ZN(n6033) );
  INV_X1 U7088 ( .A(n6029), .ZN(n6031) );
  AOI22_X1 U7089 ( .A1(n6031), .A2(n6698), .B1(n6077), .B2(n6030), .ZN(n6032)
         );
  NAND4_X1 U7090 ( .A1(n6035), .A2(n6034), .A3(n6033), .A4(n6032), .ZN(U2818)
         );
  AOI22_X1 U7091 ( .A1(EBX_REG_6__SCAN_IN), .A2(n6695), .B1(
        REIP_REG_6__SCAN_IN), .B2(n6036), .ZN(n6038) );
  AOI21_X1 U7092 ( .B1(n6078), .B2(PHYADDRPOINTER_REG_6__SCAN_IN), .A(n6045), 
        .ZN(n6037) );
  OAI211_X1 U7093 ( .C1(n6085), .C2(n6250), .A(n6038), .B(n6037), .ZN(n6040)
         );
  AOI211_X1 U7094 ( .C1(n6173), .C2(n6698), .A(n6040), .B(n6039), .ZN(n6041)
         );
  OAI21_X1 U7095 ( .B1(n6177), .B2(n6702), .A(n6041), .ZN(U2821) );
  NAND2_X1 U7096 ( .A1(n6069), .A2(n6042), .ZN(n6068) );
  AND2_X1 U7097 ( .A1(n6068), .A2(n6074), .ZN(n6062) );
  OAI22_X1 U7098 ( .A1(n6043), .A2(n6581), .B1(n6062), .B2(n6477), .ZN(n6044)
         );
  AOI211_X1 U7099 ( .C1(n6078), .C2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n6045), 
        .B(n6044), .ZN(n6053) );
  INV_X1 U7100 ( .A(n6046), .ZN(n6182) );
  NOR2_X1 U7101 ( .A1(n6047), .A2(REIP_REG_4__SCAN_IN), .ZN(n6051) );
  OAI22_X1 U7102 ( .A1(n6085), .A2(n6256), .B1(n6049), .B2(n6048), .ZN(n6050)
         );
  AOI211_X1 U7103 ( .C1(n6182), .C2(n6073), .A(n6051), .B(n6050), .ZN(n6052)
         );
  OAI211_X1 U7104 ( .C1(n6185), .C2(n6702), .A(n6053), .B(n6052), .ZN(U2823)
         );
  OR2_X1 U7105 ( .A1(n6055), .A2(n6054), .ZN(n6067) );
  AOI22_X1 U7106 ( .A1(PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n6078), .B1(n6697), 
        .B2(n6266), .ZN(n6066) );
  NOR2_X1 U7107 ( .A1(n6057), .A2(n6056), .ZN(n6064) );
  INV_X1 U7108 ( .A(REIP_REG_3__SCAN_IN), .ZN(n6474) );
  AOI22_X1 U7109 ( .A1(n6071), .A2(n6059), .B1(n6077), .B2(n6058), .ZN(n6061)
         );
  NAND2_X1 U7110 ( .A1(n6695), .A2(EBX_REG_3__SCAN_IN), .ZN(n6060) );
  OAI211_X1 U7111 ( .C1(n6062), .C2(n6474), .A(n6061), .B(n6060), .ZN(n6063)
         );
  NOR2_X1 U7112 ( .A1(n6064), .A2(n6063), .ZN(n6065) );
  OAI211_X1 U7113 ( .C1(n6068), .C2(n6067), .A(n6066), .B(n6065), .ZN(U2824)
         );
  AOI22_X1 U7114 ( .A1(n6695), .A2(EBX_REG_1__SCAN_IN), .B1(n6069), .B2(n6573), 
        .ZN(n6084) );
  NAND2_X1 U7115 ( .A1(n6071), .A2(n6070), .ZN(n6082) );
  NAND2_X1 U7116 ( .A1(n6073), .A2(n6072), .ZN(n6081) );
  INV_X1 U7117 ( .A(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n6076) );
  INV_X1 U7118 ( .A(n6074), .ZN(n6075) );
  AOI22_X1 U7119 ( .A1(n6077), .A2(n6076), .B1(n6075), .B2(REIP_REG_1__SCAN_IN), .ZN(n6080) );
  NAND2_X1 U7120 ( .A1(n6078), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n6079)
         );
  AND4_X1 U7121 ( .A1(n6082), .A2(n6081), .A3(n6080), .A4(n6079), .ZN(n6083)
         );
  OAI211_X1 U7122 ( .C1(n6086), .C2(n6085), .A(n6084), .B(n6083), .ZN(U2826)
         );
  AOI22_X1 U7123 ( .A1(n6699), .A2(n6088), .B1(n6087), .B2(n6696), .ZN(n6089)
         );
  OAI21_X1 U7124 ( .B1(n6090), .B2(n6096), .A(n6089), .ZN(U2842) );
  OAI22_X1 U7125 ( .A1(n6093), .A2(n6092), .B1(n6091), .B2(n6197), .ZN(n6094)
         );
  INV_X1 U7126 ( .A(n6094), .ZN(n6095) );
  OAI21_X1 U7127 ( .B1(n6097), .B2(n6096), .A(n6095), .ZN(U2848) );
  AOI22_X1 U7128 ( .A1(n6699), .A2(n6101), .B1(n6100), .B2(DATAI_17_), .ZN(
        n6099) );
  AOI22_X1 U7129 ( .A1(n6104), .A2(DATAI_1_), .B1(n6103), .B2(
        EAX_REG_17__SCAN_IN), .ZN(n6098) );
  NAND2_X1 U7130 ( .A1(n6099), .A2(n6098), .ZN(U2874) );
  AOI22_X1 U7131 ( .A1(n6102), .A2(n6101), .B1(n6100), .B2(DATAI_16_), .ZN(
        n6106) );
  AOI22_X1 U7132 ( .A1(n6104), .A2(DATAI_0_), .B1(n6103), .B2(
        EAX_REG_16__SCAN_IN), .ZN(n6105) );
  NAND2_X1 U7133 ( .A1(n6106), .A2(n6105), .ZN(U2875) );
  INV_X1 U7134 ( .A(UWORD_REG_11__SCAN_IN), .ZN(n6627) );
  AOI22_X1 U7135 ( .A1(n6136), .A2(DATAO_REG_27__SCAN_IN), .B1(n6108), .B2(
        EAX_REG_27__SCAN_IN), .ZN(n6107) );
  OAI21_X1 U7136 ( .B1(n6627), .B2(n6110), .A(n6107), .ZN(U2896) );
  INV_X1 U7137 ( .A(DATAO_REG_23__SCAN_IN), .ZN(n6674) );
  AOI22_X1 U7138 ( .A1(n6108), .A2(EAX_REG_23__SCAN_IN), .B1(n6553), .B2(
        UWORD_REG_7__SCAN_IN), .ZN(n6109) );
  OAI21_X1 U7139 ( .B1(n6674), .B2(n6119), .A(n6109), .ZN(U2900) );
  INV_X1 U7140 ( .A(EAX_REG_15__SCAN_IN), .ZN(n6726) );
  INV_X1 U7141 ( .A(DATAO_REG_15__SCAN_IN), .ZN(n6650) );
  OAI222_X1 U7142 ( .A1(n6110), .A2(n4432), .B1(n6138), .B2(n6726), .C1(n6650), 
        .C2(n6119), .ZN(U2908) );
  AOI22_X1 U7143 ( .A1(LWORD_REG_14__SCAN_IN), .A2(n6553), .B1(n6136), .B2(
        DATAO_REG_14__SCAN_IN), .ZN(n6111) );
  OAI21_X1 U7144 ( .B1(n6610), .B2(n6138), .A(n6111), .ZN(U2909) );
  AOI22_X1 U7145 ( .A1(LWORD_REG_13__SCAN_IN), .A2(n6553), .B1(n6136), .B2(
        DATAO_REG_13__SCAN_IN), .ZN(n6112) );
  OAI21_X1 U7146 ( .B1(n6725), .B2(n6138), .A(n6112), .ZN(U2910) );
  INV_X1 U7147 ( .A(EAX_REG_12__SCAN_IN), .ZN(n6114) );
  AOI22_X1 U7148 ( .A1(LWORD_REG_12__SCAN_IN), .A2(n6553), .B1(n6136), .B2(
        DATAO_REG_12__SCAN_IN), .ZN(n6113) );
  OAI21_X1 U7149 ( .B1(n6114), .B2(n6138), .A(n6113), .ZN(U2911) );
  INV_X1 U7150 ( .A(EAX_REG_11__SCAN_IN), .ZN(n6116) );
  AOI22_X1 U7151 ( .A1(LWORD_REG_11__SCAN_IN), .A2(n6553), .B1(n6136), .B2(
        DATAO_REG_11__SCAN_IN), .ZN(n6115) );
  OAI21_X1 U7152 ( .B1(n6116), .B2(n6138), .A(n6115), .ZN(U2912) );
  INV_X1 U7153 ( .A(DATAO_REG_10__SCAN_IN), .ZN(n6593) );
  AOI22_X1 U7154 ( .A1(EAX_REG_10__SCAN_IN), .A2(n6132), .B1(
        LWORD_REG_10__SCAN_IN), .B2(n6117), .ZN(n6118) );
  OAI21_X1 U7155 ( .B1(n6593), .B2(n6119), .A(n6118), .ZN(U2913) );
  AOI22_X1 U7156 ( .A1(LWORD_REG_9__SCAN_IN), .A2(n6553), .B1(n6136), .B2(
        DATAO_REG_9__SCAN_IN), .ZN(n6120) );
  OAI21_X1 U7157 ( .B1(n6121), .B2(n6138), .A(n6120), .ZN(U2914) );
  INV_X1 U7158 ( .A(EAX_REG_8__SCAN_IN), .ZN(n6123) );
  AOI22_X1 U7159 ( .A1(LWORD_REG_8__SCAN_IN), .A2(n6553), .B1(n6136), .B2(
        DATAO_REG_8__SCAN_IN), .ZN(n6122) );
  OAI21_X1 U7160 ( .B1(n6123), .B2(n6138), .A(n6122), .ZN(U2915) );
  AOI22_X1 U7161 ( .A1(LWORD_REG_7__SCAN_IN), .A2(n6553), .B1(n6136), .B2(
        DATAO_REG_7__SCAN_IN), .ZN(n6124) );
  OAI21_X1 U7162 ( .B1(n3739), .B2(n6138), .A(n6124), .ZN(U2916) );
  AOI22_X1 U7163 ( .A1(LWORD_REG_6__SCAN_IN), .A2(n6553), .B1(n6136), .B2(
        DATAO_REG_6__SCAN_IN), .ZN(n6125) );
  OAI21_X1 U7164 ( .B1(n6126), .B2(n6138), .A(n6125), .ZN(U2917) );
  AOI22_X1 U7165 ( .A1(LWORD_REG_5__SCAN_IN), .A2(n6553), .B1(n6136), .B2(
        DATAO_REG_5__SCAN_IN), .ZN(n6127) );
  OAI21_X1 U7166 ( .B1(n3771), .B2(n6138), .A(n6127), .ZN(U2918) );
  AOI22_X1 U7167 ( .A1(LWORD_REG_4__SCAN_IN), .A2(n6553), .B1(n6136), .B2(
        DATAO_REG_4__SCAN_IN), .ZN(n6128) );
  OAI21_X1 U7168 ( .B1(n6129), .B2(n6138), .A(n6128), .ZN(U2919) );
  AOI22_X1 U7169 ( .A1(LWORD_REG_3__SCAN_IN), .A2(n6553), .B1(n6136), .B2(
        DATAO_REG_3__SCAN_IN), .ZN(n6130) );
  OAI21_X1 U7170 ( .B1(n6131), .B2(n6138), .A(n6130), .ZN(U2920) );
  AOI222_X1 U7171 ( .A1(n6553), .A2(LWORD_REG_2__SCAN_IN), .B1(n6132), .B2(
        EAX_REG_2__SCAN_IN), .C1(DATAO_REG_2__SCAN_IN), .C2(n6136), .ZN(n6133)
         );
  INV_X1 U7172 ( .A(n6133), .ZN(U2921) );
  AOI22_X1 U7173 ( .A1(LWORD_REG_1__SCAN_IN), .A2(n6553), .B1(n6136), .B2(
        DATAO_REG_1__SCAN_IN), .ZN(n6134) );
  OAI21_X1 U7174 ( .B1(n6135), .B2(n6138), .A(n6134), .ZN(U2922) );
  AOI22_X1 U7175 ( .A1(LWORD_REG_0__SCAN_IN), .A2(n6553), .B1(n6136), .B2(
        DATAO_REG_0__SCAN_IN), .ZN(n6137) );
  OAI21_X1 U7176 ( .B1(n6673), .B2(n6138), .A(n6137), .ZN(U2923) );
  AOI22_X1 U7177 ( .A1(EAX_REG_24__SCAN_IN), .A2(n4572), .B1(n6153), .B2(
        UWORD_REG_8__SCAN_IN), .ZN(n6139) );
  NAND2_X1 U7178 ( .A1(n6143), .A2(DATAI_8_), .ZN(n6147) );
  NAND2_X1 U7179 ( .A1(n6139), .A2(n6147), .ZN(U2932) );
  AOI22_X1 U7180 ( .A1(EAX_REG_26__SCAN_IN), .A2(n4572), .B1(n6153), .B2(
        UWORD_REG_10__SCAN_IN), .ZN(n6140) );
  NAND2_X1 U7181 ( .A1(n6143), .A2(DATAI_10_), .ZN(n6149) );
  NAND2_X1 U7182 ( .A1(n6140), .A2(n6149), .ZN(U2934) );
  NAND2_X1 U7183 ( .A1(n6143), .A2(DATAI_11_), .ZN(n6151) );
  INV_X1 U7184 ( .A(n6151), .ZN(n6141) );
  AOI21_X1 U7185 ( .B1(n4572), .B2(EAX_REG_27__SCAN_IN), .A(n6141), .ZN(n6142)
         );
  OAI21_X1 U7186 ( .B1(n6627), .B2(n6146), .A(n6142), .ZN(U2935) );
  INV_X1 U7187 ( .A(UWORD_REG_12__SCAN_IN), .ZN(n6608) );
  NAND2_X1 U7188 ( .A1(n6143), .A2(DATAI_12_), .ZN(n6154) );
  INV_X1 U7189 ( .A(n6154), .ZN(n6144) );
  AOI21_X1 U7190 ( .B1(n4572), .B2(EAX_REG_28__SCAN_IN), .A(n6144), .ZN(n6145)
         );
  OAI21_X1 U7191 ( .B1(n6608), .B2(n6146), .A(n6145), .ZN(U2936) );
  AOI22_X1 U7192 ( .A1(EAX_REG_8__SCAN_IN), .A2(n4572), .B1(n6153), .B2(
        LWORD_REG_8__SCAN_IN), .ZN(n6148) );
  NAND2_X1 U7193 ( .A1(n6148), .A2(n6147), .ZN(U2947) );
  AOI22_X1 U7194 ( .A1(EAX_REG_10__SCAN_IN), .A2(n4572), .B1(n6153), .B2(
        LWORD_REG_10__SCAN_IN), .ZN(n6150) );
  NAND2_X1 U7195 ( .A1(n6150), .A2(n6149), .ZN(U2949) );
  AOI22_X1 U7196 ( .A1(EAX_REG_11__SCAN_IN), .A2(n4572), .B1(n6153), .B2(
        LWORD_REG_11__SCAN_IN), .ZN(n6152) );
  NAND2_X1 U7197 ( .A1(n6152), .A2(n6151), .ZN(U2950) );
  AOI22_X1 U7198 ( .A1(EAX_REG_12__SCAN_IN), .A2(n4572), .B1(n6153), .B2(
        LWORD_REG_12__SCAN_IN), .ZN(n6155) );
  NAND2_X1 U7199 ( .A1(n6155), .A2(n6154), .ZN(U2951) );
  NAND2_X1 U7200 ( .A1(n6157), .A2(n6156), .ZN(n6159) );
  NAND2_X1 U7201 ( .A1(n6159), .A2(n6158), .ZN(n6162) );
  XNOR2_X1 U7202 ( .A(n6160), .B(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n6161)
         );
  XNOR2_X1 U7203 ( .A(n6162), .B(n6161), .ZN(n6198) );
  AOI22_X1 U7204 ( .A1(n3668), .A2(REIP_REG_11__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n6186), .ZN(n6168) );
  AOI22_X1 U7205 ( .A1(n6166), .A2(n6165), .B1(n6164), .B2(n6163), .ZN(n6167)
         );
  OAI211_X1 U7206 ( .C1(n6198), .C2(n6169), .A(n6168), .B(n6167), .ZN(U2975)
         );
  AOI22_X1 U7207 ( .A1(n3668), .A2(REIP_REG_6__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n6186), .ZN(n6176) );
  OAI21_X1 U7208 ( .B1(n6172), .B2(n6171), .A(n6170), .ZN(n6247) );
  INV_X1 U7209 ( .A(n6247), .ZN(n6174) );
  AOI22_X1 U7210 ( .A1(n6174), .A2(n6191), .B1(n6165), .B2(n6173), .ZN(n6175)
         );
  OAI211_X1 U7211 ( .C1(n6195), .C2(n6177), .A(n6176), .B(n6175), .ZN(U2980)
         );
  AOI22_X1 U7212 ( .A1(n3668), .A2(REIP_REG_4__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n6186), .ZN(n6184) );
  OAI21_X1 U7213 ( .B1(n6180), .B2(n6179), .A(n6178), .ZN(n6181) );
  INV_X1 U7214 ( .A(n6181), .ZN(n6257) );
  AOI22_X1 U7215 ( .A1(n6257), .A2(n6191), .B1(n6165), .B2(n6182), .ZN(n6183)
         );
  OAI211_X1 U7216 ( .C1(n6195), .C2(n6185), .A(n6184), .B(n6183), .ZN(U2982)
         );
  AOI22_X1 U7217 ( .A1(n3668), .A2(REIP_REG_2__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n6186), .ZN(n6193) );
  XOR2_X1 U7218 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .B(n6187), .Z(n6189) );
  XNOR2_X1 U7219 ( .A(n6189), .B(n6188), .ZN(n6283) );
  AOI22_X1 U7220 ( .A1(n6283), .A2(n6191), .B1(n6165), .B2(n6190), .ZN(n6192)
         );
  OAI211_X1 U7221 ( .C1(n6195), .C2(n6194), .A(n6193), .B(n6192), .ZN(U2984)
         );
  INV_X1 U7222 ( .A(n6196), .ZN(n6201) );
  OAI22_X1 U7223 ( .A1(n6249), .A2(n6197), .B1(n6488), .B2(n6248), .ZN(n6200)
         );
  NOR2_X1 U7224 ( .A1(n6198), .A2(n5780), .ZN(n6199) );
  AOI211_X1 U7225 ( .C1(n6202), .C2(n6201), .A(n6200), .B(n6199), .ZN(n6203)
         );
  OAI21_X1 U7226 ( .B1(n6204), .B2(n6202), .A(n6203), .ZN(U3007) );
  AOI22_X1 U7227 ( .A1(n6208), .A2(n6207), .B1(n6206), .B2(n6205), .ZN(n6209)
         );
  INV_X1 U7228 ( .A(n6209), .ZN(n6241) );
  AOI21_X1 U7229 ( .B1(n6227), .B2(n6210), .A(n6241), .ZN(n6226) );
  OAI22_X1 U7230 ( .A1(n6249), .A2(n6211), .B1(n6486), .B2(n6248), .ZN(n6212)
         );
  AOI21_X1 U7231 ( .B1(n6213), .B2(n6282), .A(n6212), .ZN(n6217) );
  OAI21_X1 U7232 ( .B1(n6284), .B2(n6274), .A(n6276), .ZN(n6260) );
  NAND2_X1 U7233 ( .A1(n6214), .A2(n6260), .ZN(n6245) );
  NOR2_X1 U7234 ( .A1(n6227), .A2(n6245), .ZN(n6221) );
  OAI211_X1 U7235 ( .C1(INSTADDRPOINTER_REG_10__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_9__SCAN_IN), .A(n6221), .B(n6215), .ZN(n6216) );
  OAI211_X1 U7236 ( .C1(n6226), .C2(n3418), .A(n6217), .B(n6216), .ZN(U3008)
         );
  INV_X1 U7237 ( .A(n6218), .ZN(n6219) );
  AOI21_X1 U7238 ( .B1(n6280), .B2(n6220), .A(n6219), .ZN(n6224) );
  AOI22_X1 U7239 ( .A1(n6222), .A2(n6282), .B1(n6221), .B2(n6225), .ZN(n6223)
         );
  OAI211_X1 U7240 ( .C1(n6226), .C2(n6225), .A(n6224), .B(n6223), .ZN(U3009)
         );
  OAI21_X1 U7241 ( .B1(INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_7__SCAN_IN), .A(n6227), .ZN(n6236) );
  INV_X1 U7242 ( .A(n6228), .ZN(n6231) );
  INV_X1 U7243 ( .A(n6229), .ZN(n6230) );
  AOI21_X1 U7244 ( .B1(n6280), .B2(n6231), .A(n6230), .ZN(n6235) );
  INV_X1 U7245 ( .A(n6232), .ZN(n6233) );
  AOI22_X1 U7246 ( .A1(n6233), .A2(n6282), .B1(INSTADDRPOINTER_REG_8__SCAN_IN), 
        .B2(n6241), .ZN(n6234) );
  OAI211_X1 U7247 ( .C1(n6245), .C2(n6236), .A(n6235), .B(n6234), .ZN(U3010)
         );
  INV_X1 U7248 ( .A(n6237), .ZN(n6238) );
  AOI21_X1 U7249 ( .B1(n6280), .B2(n6239), .A(n6238), .ZN(n6244) );
  INV_X1 U7250 ( .A(n6240), .ZN(n6242) );
  AOI22_X1 U7251 ( .A1(n6242), .A2(n6282), .B1(INSTADDRPOINTER_REG_7__SCAN_IN), 
        .B2(n6241), .ZN(n6243) );
  OAI211_X1 U7252 ( .C1(INSTADDRPOINTER_REG_7__SCAN_IN), .C2(n6245), .A(n6244), 
        .B(n6243), .ZN(U3011) );
  NAND2_X1 U7253 ( .A1(n6246), .A2(n6260), .ZN(n6255) );
  OAI222_X1 U7254 ( .A1(n6250), .A2(n6249), .B1(n6248), .B2(n6480), .C1(n5780), 
        .C2(n6247), .ZN(n6251) );
  INV_X1 U7255 ( .A(n6251), .ZN(n6252) );
  OAI221_X1 U7256 ( .B1(INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n6255), .C1(n6254), .C2(n6253), .A(n6252), .ZN(U3012) );
  NOR2_X1 U7257 ( .A1(n6276), .A2(n6259), .ZN(n6277) );
  NOR2_X1 U7258 ( .A1(n6277), .A2(n6281), .ZN(n6273) );
  INV_X1 U7259 ( .A(n6256), .ZN(n6258) );
  AOI222_X1 U7260 ( .A1(REIP_REG_4__SCAN_IN), .A2(n3668), .B1(n6280), .B2(
        n6258), .C1(n6282), .C2(n6257), .ZN(n6263) );
  AND2_X1 U7261 ( .A1(n6260), .A2(n6259), .ZN(n6269) );
  OAI211_X1 U7262 ( .C1(INSTADDRPOINTER_REG_4__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_3__SCAN_IN), .A(n6269), .B(n6261), .ZN(n6262) );
  OAI211_X1 U7263 ( .C1(n6273), .C2(n6646), .A(n6263), .B(n6262), .ZN(U3014)
         );
  INV_X1 U7264 ( .A(n6264), .ZN(n6265) );
  AOI21_X1 U7265 ( .B1(n6280), .B2(n6266), .A(n6265), .ZN(n6271) );
  INV_X1 U7266 ( .A(n6267), .ZN(n6268) );
  AOI22_X1 U7267 ( .A1(n6269), .A2(n6272), .B1(n6268), .B2(n6282), .ZN(n6270)
         );
  OAI211_X1 U7268 ( .C1(n6273), .C2(n6272), .A(n6271), .B(n6270), .ZN(U3015)
         );
  NOR3_X1 U7269 ( .A1(n6276), .A2(n6275), .A3(n6274), .ZN(n6278) );
  AOI211_X1 U7270 ( .C1(n6280), .C2(n6279), .A(n6278), .B(n6277), .ZN(n6290)
         );
  AOI22_X1 U7271 ( .A1(n6283), .A2(n6282), .B1(INSTADDRPOINTER_REG_2__SCAN_IN), 
        .B2(n6281), .ZN(n6289) );
  NAND2_X1 U7272 ( .A1(n3668), .A2(REIP_REG_2__SCAN_IN), .ZN(n6288) );
  INV_X1 U7273 ( .A(n6284), .ZN(n6286) );
  NAND3_X1 U7274 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n6286), .A3(n6285), 
        .ZN(n6287) );
  NAND4_X1 U7275 ( .A1(n6290), .A2(n6289), .A3(n6288), .A4(n6287), .ZN(U3016)
         );
  NOR2_X1 U7276 ( .A1(n6417), .A2(n6291), .ZN(U3019) );
  AOI22_X1 U7277 ( .A1(n6303), .A2(n6326), .B1(n6325), .B2(n6302), .ZN(n6293)
         );
  AOI22_X1 U7278 ( .A1(INSTQUEUE_REG_3__2__SCAN_IN), .A2(n6305), .B1(n6327), 
        .B2(n6304), .ZN(n6292) );
  OAI211_X1 U7279 ( .C1(n6308), .C2(n6330), .A(n6293), .B(n6292), .ZN(U3046)
         );
  AOI22_X1 U7280 ( .A1(n6303), .A2(n6347), .B1(n6346), .B2(n6302), .ZN(n6295)
         );
  AOI22_X1 U7281 ( .A1(INSTQUEUE_REG_3__3__SCAN_IN), .A2(n6305), .B1(n6348), 
        .B2(n6304), .ZN(n6294) );
  OAI211_X1 U7282 ( .C1(n6308), .C2(n6351), .A(n6295), .B(n6294), .ZN(U3047)
         );
  AOI22_X1 U7283 ( .A1(n6303), .A2(n6297), .B1(n6296), .B2(n6302), .ZN(n6300)
         );
  AOI22_X1 U7284 ( .A1(INSTQUEUE_REG_3__4__SCAN_IN), .A2(n6305), .B1(n6298), 
        .B2(n6304), .ZN(n6299) );
  OAI211_X1 U7285 ( .C1(n6308), .C2(n6301), .A(n6300), .B(n6299), .ZN(U3048)
         );
  AOI22_X1 U7286 ( .A1(n6303), .A2(n6366), .B1(n6365), .B2(n6302), .ZN(n6307)
         );
  AOI22_X1 U7287 ( .A1(INSTQUEUE_REG_3__7__SCAN_IN), .A2(n6305), .B1(n6369), 
        .B2(n6304), .ZN(n6306) );
  OAI211_X1 U7288 ( .C1(n6308), .C2(n6374), .A(n6307), .B(n6306), .ZN(U3051)
         );
  INV_X1 U7289 ( .A(n6309), .ZN(n6317) );
  AOI22_X1 U7290 ( .A1(n6376), .A2(n6317), .B1(n6375), .B2(n6316), .ZN(n6312)
         );
  AOI22_X1 U7291 ( .A1(n6320), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n6310), 
        .B2(n6318), .ZN(n6311) );
  OAI211_X1 U7292 ( .C1(n6379), .C2(n6341), .A(n6312), .B(n6311), .ZN(U3068)
         );
  AOI22_X1 U7293 ( .A1(n6386), .A2(n6317), .B1(n6383), .B2(n6316), .ZN(n6315)
         );
  AOI22_X1 U7294 ( .A1(n6320), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n6313), 
        .B2(n6318), .ZN(n6314) );
  OAI211_X1 U7295 ( .C1(n6390), .C2(n6341), .A(n6315), .B(n6314), .ZN(U3069)
         );
  AOI22_X1 U7296 ( .A1(n6327), .A2(n6317), .B1(n6325), .B2(n6316), .ZN(n6322)
         );
  AOI22_X1 U7297 ( .A1(n6320), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n6319), 
        .B2(n6318), .ZN(n6321) );
  OAI211_X1 U7298 ( .C1(n6323), .C2(n6341), .A(n6322), .B(n6321), .ZN(U3070)
         );
  INV_X1 U7299 ( .A(n6324), .ZN(n6335) );
  AOI22_X1 U7300 ( .A1(n6336), .A2(n6326), .B1(n6325), .B2(n6335), .ZN(n6329)
         );
  AOI22_X1 U7301 ( .A1(INSTQUEUE_REG_7__2__SCAN_IN), .A2(n6338), .B1(n6327), 
        .B2(n6337), .ZN(n6328) );
  OAI211_X1 U7302 ( .C1(n6330), .C2(n6341), .A(n6329), .B(n6328), .ZN(U3078)
         );
  AOI22_X1 U7303 ( .A1(n6336), .A2(n6347), .B1(n6346), .B2(n6335), .ZN(n6332)
         );
  AOI22_X1 U7304 ( .A1(INSTQUEUE_REG_7__3__SCAN_IN), .A2(n6338), .B1(n6348), 
        .B2(n6337), .ZN(n6331) );
  OAI211_X1 U7305 ( .C1(n6351), .C2(n6341), .A(n6332), .B(n6331), .ZN(U3079)
         );
  AOI22_X1 U7306 ( .A1(n6336), .A2(n6353), .B1(n6352), .B2(n6335), .ZN(n6334)
         );
  AOI22_X1 U7307 ( .A1(INSTQUEUE_REG_7__5__SCAN_IN), .A2(n6338), .B1(n6354), 
        .B2(n6337), .ZN(n6333) );
  OAI211_X1 U7308 ( .C1(n6357), .C2(n6341), .A(n6334), .B(n6333), .ZN(U3081)
         );
  AOI22_X1 U7309 ( .A1(n6336), .A2(n6359), .B1(n6358), .B2(n6335), .ZN(n6340)
         );
  AOI22_X1 U7310 ( .A1(INSTQUEUE_REG_7__6__SCAN_IN), .A2(n6338), .B1(n6360), 
        .B2(n6337), .ZN(n6339) );
  OAI211_X1 U7311 ( .C1(n6363), .C2(n6341), .A(n6340), .B(n6339), .ZN(U3082)
         );
  INV_X1 U7312 ( .A(n6342), .ZN(n6364) );
  AOI22_X1 U7313 ( .A1(n6367), .A2(n6343), .B1(n6383), .B2(n6364), .ZN(n6345)
         );
  AOI22_X1 U7314 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(n6370), .B1(n6386), 
        .B2(n6368), .ZN(n6344) );
  OAI211_X1 U7315 ( .C1(n6387), .C2(n6373), .A(n6345), .B(n6344), .ZN(U3109)
         );
  AOI22_X1 U7316 ( .A1(n6367), .A2(n6347), .B1(n6346), .B2(n6364), .ZN(n6350)
         );
  AOI22_X1 U7317 ( .A1(INSTQUEUE_REG_11__3__SCAN_IN), .A2(n6370), .B1(n6348), 
        .B2(n6368), .ZN(n6349) );
  OAI211_X1 U7318 ( .C1(n6351), .C2(n6373), .A(n6350), .B(n6349), .ZN(U3111)
         );
  AOI22_X1 U7319 ( .A1(n6367), .A2(n6353), .B1(n6352), .B2(n6364), .ZN(n6356)
         );
  AOI22_X1 U7320 ( .A1(INSTQUEUE_REG_11__5__SCAN_IN), .A2(n6370), .B1(n6354), 
        .B2(n6368), .ZN(n6355) );
  OAI211_X1 U7321 ( .C1(n6357), .C2(n6373), .A(n6356), .B(n6355), .ZN(U3113)
         );
  AOI22_X1 U7322 ( .A1(n6367), .A2(n6359), .B1(n6358), .B2(n6364), .ZN(n6362)
         );
  AOI22_X1 U7323 ( .A1(INSTQUEUE_REG_11__6__SCAN_IN), .A2(n6370), .B1(n6360), 
        .B2(n6368), .ZN(n6361) );
  OAI211_X1 U7324 ( .C1(n6363), .C2(n6373), .A(n6362), .B(n6361), .ZN(U3114)
         );
  AOI22_X1 U7325 ( .A1(n6367), .A2(n6366), .B1(n6365), .B2(n6364), .ZN(n6372)
         );
  AOI22_X1 U7326 ( .A1(INSTQUEUE_REG_11__7__SCAN_IN), .A2(n6370), .B1(n6369), 
        .B2(n6368), .ZN(n6371) );
  OAI211_X1 U7327 ( .C1(n6374), .C2(n6373), .A(n6372), .B(n6371), .ZN(U3115)
         );
  AOI22_X1 U7328 ( .A1(n6376), .A2(n6385), .B1(n6384), .B2(n6375), .ZN(n6382)
         );
  OR2_X1 U7329 ( .A1(n6388), .A2(n6377), .ZN(n6378) );
  OAI21_X1 U7330 ( .B1(n6391), .B2(n6379), .A(n6378), .ZN(n6380) );
  INV_X1 U7331 ( .A(n6380), .ZN(n6381) );
  OAI211_X1 U7332 ( .C1(n6395), .C2(n6710), .A(n6382), .B(n6381), .ZN(U3140)
         );
  INV_X1 U7333 ( .A(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n6583) );
  AOI22_X1 U7334 ( .A1(n6386), .A2(n6385), .B1(n6384), .B2(n6383), .ZN(n6394)
         );
  OR2_X1 U7335 ( .A1(n6388), .A2(n6387), .ZN(n6389) );
  OAI21_X1 U7336 ( .B1(n6391), .B2(n6390), .A(n6389), .ZN(n6392) );
  INV_X1 U7337 ( .A(n6392), .ZN(n6393) );
  OAI211_X1 U7338 ( .C1(n6395), .C2(n6583), .A(n6394), .B(n6393), .ZN(U3141)
         );
  INV_X1 U7339 ( .A(n6396), .ZN(n6398) );
  NOR3_X1 U7340 ( .A1(n6399), .A2(n6398), .A3(n6397), .ZN(n6422) );
  INV_X1 U7341 ( .A(n6416), .ZN(n6420) );
  INV_X1 U7342 ( .A(n6411), .ZN(n6414) );
  AOI22_X1 U7343 ( .A1(n6403), .A2(n6402), .B1(n6401), .B2(n6400), .ZN(n6537)
         );
  NAND2_X1 U7344 ( .A1(n6404), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n6543) );
  AND3_X1 U7345 ( .A1(n6537), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A3(n6543), 
        .ZN(n6405) );
  INV_X1 U7346 ( .A(n6405), .ZN(n6409) );
  OAI22_X1 U7347 ( .A1(n6407), .A2(n6406), .B1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n6405), .ZN(n6408) );
  OAI21_X1 U7348 ( .B1(n6409), .B2(n6612), .A(n6408), .ZN(n6410) );
  INV_X1 U7349 ( .A(n6410), .ZN(n6413) );
  OAI21_X1 U7350 ( .B1(n6411), .B2(n6410), .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), 
        .ZN(n6412) );
  OAI21_X1 U7351 ( .B1(n6414), .B2(n6413), .A(n6412), .ZN(n6415) );
  OAI21_X1 U7352 ( .B1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n6416), .A(n6415), 
        .ZN(n6418) );
  OAI211_X1 U7353 ( .C1(n6420), .C2(n6419), .A(n6418), .B(n6417), .ZN(n6421)
         );
  NAND3_X1 U7354 ( .A1(n6423), .A2(n6422), .A3(n6421), .ZN(n6424) );
  AOI221_X1 U7355 ( .B1(FLUSH_REG_SCAN_IN), .B2(n6425), .C1(MORE_REG_SCAN_IN), 
        .C2(n6425), .A(n6424), .ZN(n6433) );
  NOR2_X1 U7356 ( .A1(n6433), .A2(STATE2_REG_1__SCAN_IN), .ZN(n6432) );
  OR2_X1 U7357 ( .A1(n6427), .A2(n6426), .ZN(n6431) );
  NAND3_X1 U7358 ( .A1(STATE2_REG_2__SCAN_IN), .A2(READY_N), .A3(n6443), .ZN(
        n6428) );
  NAND2_X1 U7359 ( .A1(n6429), .A2(n6428), .ZN(n6430) );
  NAND2_X1 U7360 ( .A1(n6431), .A2(n6430), .ZN(n6434) );
  OR2_X1 U7361 ( .A1(n6432), .A2(n6434), .ZN(n6531) );
  INV_X1 U7362 ( .A(n6531), .ZN(n6445) );
  AOI21_X1 U7363 ( .B1(READY_N), .B2(n6661), .A(n6445), .ZN(n6444) );
  INV_X1 U7364 ( .A(n6433), .ZN(n6439) );
  INV_X1 U7365 ( .A(n6434), .ZN(n6436) );
  NOR2_X1 U7366 ( .A1(n6451), .A2(n6533), .ZN(n6435) );
  AOI211_X1 U7367 ( .C1(STATE2_REG_1__SCAN_IN), .C2(n6436), .A(
        STATE2_REG_0__SCAN_IN), .B(n6435), .ZN(n6437) );
  AOI211_X1 U7368 ( .C1(n6440), .C2(n6439), .A(n6438), .B(n6437), .ZN(n6441)
         );
  OAI221_X1 U7369 ( .B1(n6443), .B2(n6444), .C1(n6443), .C2(n6442), .A(n6441), 
        .ZN(U3148) );
  NOR3_X1 U7370 ( .A1(n6454), .A2(n6444), .A3(n6536), .ZN(n6449) );
  AOI221_X1 U7371 ( .B1(READY_N), .B2(n6447), .C1(n6446), .C2(n6447), .A(n6445), .ZN(n6448) );
  OR3_X1 U7372 ( .A1(n6450), .A2(n6449), .A3(n6448), .ZN(U3149) );
  OAI211_X1 U7373 ( .C1(STATE2_REG_2__SCAN_IN), .C2(n6554), .A(n6529), .B(
        n6451), .ZN(n6453) );
  OAI21_X1 U7374 ( .B1(n6454), .B2(n6453), .A(n6452), .ZN(U3150) );
  INV_X1 U7375 ( .A(n6528), .ZN(n6455) );
  AND2_X1 U7376 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(n6455), .ZN(U3151) );
  AND2_X1 U7377 ( .A1(DATAWIDTH_REG_30__SCAN_IN), .A2(n6455), .ZN(U3152) );
  AND2_X1 U7378 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(n6455), .ZN(U3153) );
  AND2_X1 U7379 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(n6455), .ZN(U3154) );
  AND2_X1 U7380 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(n6455), .ZN(U3155) );
  AND2_X1 U7381 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(n6455), .ZN(U3156) );
  AND2_X1 U7382 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(n6455), .ZN(U3157) );
  AND2_X1 U7383 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(n6455), .ZN(U3158) );
  AND2_X1 U7384 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(n6455), .ZN(U3159) );
  AND2_X1 U7385 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(n6455), .ZN(U3160) );
  AND2_X1 U7386 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(n6455), .ZN(U3161) );
  AND2_X1 U7387 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(n6455), .ZN(U3162) );
  AND2_X1 U7388 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(n6455), .ZN(U3163) );
  AND2_X1 U7389 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(n6455), .ZN(U3164) );
  AND2_X1 U7390 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(n6455), .ZN(U3165) );
  AND2_X1 U7391 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(n6455), .ZN(U3166) );
  INV_X1 U7392 ( .A(DATAWIDTH_REG_15__SCAN_IN), .ZN(n6626) );
  NOR2_X1 U7393 ( .A1(n6528), .A2(n6626), .ZN(U3167) );
  AND2_X1 U7394 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(n6455), .ZN(U3168) );
  AND2_X1 U7395 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(n6455), .ZN(U3169) );
  AND2_X1 U7396 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(n6455), .ZN(U3170) );
  AND2_X1 U7397 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(n6455), .ZN(U3171) );
  AND2_X1 U7398 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(n6455), .ZN(U3172) );
  AND2_X1 U7399 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(n6455), .ZN(U3173) );
  AND2_X1 U7400 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(n6455), .ZN(U3174) );
  AND2_X1 U7401 ( .A1(DATAWIDTH_REG_7__SCAN_IN), .A2(n6455), .ZN(U3175) );
  AND2_X1 U7402 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(n6455), .ZN(U3176) );
  INV_X1 U7403 ( .A(DATAWIDTH_REG_5__SCAN_IN), .ZN(n6644) );
  NOR2_X1 U7404 ( .A1(n6528), .A2(n6644), .ZN(U3177) );
  AND2_X1 U7405 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(n6455), .ZN(U3178) );
  AND2_X1 U7406 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(n6455), .ZN(U3179) );
  AND2_X1 U7407 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(n6455), .ZN(U3180) );
  NOR2_X1 U7408 ( .A1(n6716), .A2(n6462), .ZN(n6463) );
  AOI22_X1 U7409 ( .A1(READY_N), .A2(STATE_REG_1__SCAN_IN), .B1(
        STATE_REG_2__SCAN_IN), .B2(HOLD), .ZN(n6471) );
  AND2_X1 U7410 ( .A1(STATE_REG_1__SCAN_IN), .A2(HOLD), .ZN(n6459) );
  INV_X1 U7411 ( .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6457) );
  INV_X1 U7412 ( .A(NA_N), .ZN(n6464) );
  AOI221_X1 U7413 ( .B1(STATE_REG_1__SCAN_IN), .B2(STATE_REG_2__SCAN_IN), .C1(
        n6464), .C2(STATE_REG_2__SCAN_IN), .A(STATE_REG_0__SCAN_IN), .ZN(n6468) );
  AOI221_X1 U7414 ( .B1(n6459), .B2(n6565), .C1(n6457), .C2(n6565), .A(n6468), 
        .ZN(n6456) );
  OAI21_X1 U7415 ( .B1(n6463), .B2(n6471), .A(n6456), .ZN(U3181) );
  NOR2_X1 U7416 ( .A1(n6466), .A2(n6457), .ZN(n6465) );
  NAND2_X1 U7417 ( .A1(STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n6458) );
  OAI21_X1 U7418 ( .B1(n6465), .B2(n6459), .A(n6458), .ZN(n6460) );
  OAI211_X1 U7419 ( .C1(n6462), .C2(n6554), .A(n6461), .B(n6460), .ZN(U3182)
         );
  AOI21_X1 U7420 ( .B1(n6465), .B2(n6464), .A(n6463), .ZN(n6470) );
  AOI221_X1 U7421 ( .B1(NA_N), .B2(STATE_REG_1__SCAN_IN), .C1(n6554), .C2(
        STATE_REG_1__SCAN_IN), .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6467) );
  AOI221_X1 U7422 ( .B1(STATE_REG_2__SCAN_IN), .B2(HOLD), .C1(n6467), .C2(HOLD), .A(n6466), .ZN(n6469) );
  OAI22_X1 U7423 ( .A1(n6471), .A2(n6470), .B1(n6469), .B2(n6468), .ZN(U3183)
         );
  NOR2_X2 U7424 ( .A1(n6716), .A2(n6565), .ZN(n6521) );
  INV_X1 U7425 ( .A(n6521), .ZN(n6519) );
  NAND2_X1 U7426 ( .A1(n6716), .A2(n6485), .ZN(n6523) );
  INV_X1 U7427 ( .A(n6523), .ZN(n6517) );
  AOI22_X1 U7428 ( .A1(REIP_REG_2__SCAN_IN), .A2(n6517), .B1(
        ADDRESS_REG_0__SCAN_IN), .B2(n6509), .ZN(n6472) );
  OAI21_X1 U7429 ( .B1(n6573), .B2(n6519), .A(n6472), .ZN(U3184) );
  AOI22_X1 U7430 ( .A1(REIP_REG_2__SCAN_IN), .A2(n6521), .B1(
        ADDRESS_REG_1__SCAN_IN), .B2(n6509), .ZN(n6473) );
  OAI21_X1 U7431 ( .B1(n6474), .B2(n6523), .A(n6473), .ZN(U3185) );
  AOI22_X1 U7432 ( .A1(REIP_REG_3__SCAN_IN), .A2(n6521), .B1(
        ADDRESS_REG_2__SCAN_IN), .B2(n6509), .ZN(n6475) );
  OAI21_X1 U7433 ( .B1(n6477), .B2(n6523), .A(n6475), .ZN(U3186) );
  AOI22_X1 U7434 ( .A1(REIP_REG_5__SCAN_IN), .A2(n6517), .B1(
        ADDRESS_REG_3__SCAN_IN), .B2(n6509), .ZN(n6476) );
  OAI21_X1 U7435 ( .B1(n6477), .B2(n6519), .A(n6476), .ZN(U3187) );
  AOI22_X1 U7436 ( .A1(REIP_REG_5__SCAN_IN), .A2(n6521), .B1(
        ADDRESS_REG_4__SCAN_IN), .B2(n6509), .ZN(n6478) );
  OAI21_X1 U7437 ( .B1(n6480), .B2(n6523), .A(n6478), .ZN(U3188) );
  AOI22_X1 U7438 ( .A1(REIP_REG_7__SCAN_IN), .A2(n6517), .B1(
        ADDRESS_REG_5__SCAN_IN), .B2(n6509), .ZN(n6479) );
  OAI21_X1 U7439 ( .B1(n6480), .B2(n6519), .A(n6479), .ZN(U3189) );
  AOI22_X1 U7440 ( .A1(REIP_REG_7__SCAN_IN), .A2(n6521), .B1(
        ADDRESS_REG_6__SCAN_IN), .B2(n6509), .ZN(n6481) );
  OAI21_X1 U7441 ( .B1(n6483), .B2(n6523), .A(n6481), .ZN(U3190) );
  AOI22_X1 U7442 ( .A1(REIP_REG_9__SCAN_IN), .A2(n6517), .B1(
        ADDRESS_REG_7__SCAN_IN), .B2(n6509), .ZN(n6482) );
  OAI21_X1 U7443 ( .B1(n6483), .B2(n6519), .A(n6482), .ZN(U3191) );
  INV_X1 U7444 ( .A(ADDRESS_REG_8__SCAN_IN), .ZN(n6643) );
  OAI222_X1 U7445 ( .A1(n6523), .A2(n6486), .B1(n6643), .B2(n6485), .C1(n6484), 
        .C2(n6519), .ZN(U3192) );
  AOI22_X1 U7446 ( .A1(REIP_REG_10__SCAN_IN), .A2(n6521), .B1(
        ADDRESS_REG_9__SCAN_IN), .B2(n6509), .ZN(n6487) );
  OAI21_X1 U7447 ( .B1(n6488), .B2(n6523), .A(n6487), .ZN(U3193) );
  AOI22_X1 U7448 ( .A1(REIP_REG_11__SCAN_IN), .A2(n6521), .B1(
        ADDRESS_REG_10__SCAN_IN), .B2(n6509), .ZN(n6489) );
  OAI21_X1 U7449 ( .B1(n6635), .B2(n6523), .A(n6489), .ZN(U3194) );
  AOI22_X1 U7450 ( .A1(REIP_REG_13__SCAN_IN), .A2(n6517), .B1(
        ADDRESS_REG_11__SCAN_IN), .B2(n6509), .ZN(n6490) );
  OAI21_X1 U7451 ( .B1(n6635), .B2(n6519), .A(n6490), .ZN(U3195) );
  AOI22_X1 U7452 ( .A1(REIP_REG_14__SCAN_IN), .A2(n6517), .B1(
        ADDRESS_REG_12__SCAN_IN), .B2(n6509), .ZN(n6491) );
  OAI21_X1 U7453 ( .B1(n6492), .B2(n6519), .A(n6491), .ZN(U3196) );
  AOI22_X1 U7454 ( .A1(REIP_REG_14__SCAN_IN), .A2(n6521), .B1(
        ADDRESS_REG_13__SCAN_IN), .B2(n6509), .ZN(n6493) );
  OAI21_X1 U7455 ( .B1(n6574), .B2(n6523), .A(n6493), .ZN(U3197) );
  AOI22_X1 U7456 ( .A1(REIP_REG_15__SCAN_IN), .A2(n6521), .B1(
        ADDRESS_REG_14__SCAN_IN), .B2(n6509), .ZN(n6494) );
  OAI21_X1 U7457 ( .B1(n6496), .B2(n6523), .A(n6494), .ZN(U3198) );
  AOI22_X1 U7458 ( .A1(REIP_REG_17__SCAN_IN), .A2(n6517), .B1(
        ADDRESS_REG_15__SCAN_IN), .B2(n6509), .ZN(n6495) );
  OAI21_X1 U7459 ( .B1(n6496), .B2(n6519), .A(n6495), .ZN(U3199) );
  AOI22_X1 U7460 ( .A1(REIP_REG_17__SCAN_IN), .A2(n6521), .B1(
        ADDRESS_REG_16__SCAN_IN), .B2(n6509), .ZN(n6497) );
  OAI21_X1 U7461 ( .B1(n6499), .B2(n6523), .A(n6497), .ZN(U3200) );
  AOI22_X1 U7462 ( .A1(REIP_REG_19__SCAN_IN), .A2(n6517), .B1(
        ADDRESS_REG_17__SCAN_IN), .B2(n6509), .ZN(n6498) );
  OAI21_X1 U7463 ( .B1(n6499), .B2(n6519), .A(n6498), .ZN(U3201) );
  AOI22_X1 U7464 ( .A1(REIP_REG_20__SCAN_IN), .A2(n6517), .B1(
        ADDRESS_REG_18__SCAN_IN), .B2(n6509), .ZN(n6500) );
  OAI21_X1 U7465 ( .B1(n6501), .B2(n6519), .A(n6500), .ZN(U3202) );
  AOI222_X1 U7466 ( .A1(n6521), .A2(REIP_REG_20__SCAN_IN), .B1(
        ADDRESS_REG_19__SCAN_IN), .B2(n6565), .C1(REIP_REG_21__SCAN_IN), .C2(
        n6517), .ZN(n6502) );
  INV_X1 U7467 ( .A(n6502), .ZN(U3203) );
  AOI22_X1 U7468 ( .A1(REIP_REG_21__SCAN_IN), .A2(n6521), .B1(
        ADDRESS_REG_20__SCAN_IN), .B2(n6509), .ZN(n6503) );
  OAI21_X1 U7469 ( .B1(n4018), .B2(n6523), .A(n6503), .ZN(U3204) );
  AOI22_X1 U7470 ( .A1(REIP_REG_23__SCAN_IN), .A2(n6517), .B1(
        ADDRESS_REG_21__SCAN_IN), .B2(n6509), .ZN(n6504) );
  OAI21_X1 U7471 ( .B1(n4018), .B2(n6519), .A(n6504), .ZN(U3205) );
  AOI22_X1 U7472 ( .A1(REIP_REG_23__SCAN_IN), .A2(n6521), .B1(
        ADDRESS_REG_22__SCAN_IN), .B2(n6509), .ZN(n6505) );
  OAI21_X1 U7473 ( .B1(n6506), .B2(n6523), .A(n6505), .ZN(U3206) );
  AOI22_X1 U7474 ( .A1(REIP_REG_24__SCAN_IN), .A2(n6521), .B1(
        ADDRESS_REG_23__SCAN_IN), .B2(n6509), .ZN(n6507) );
  OAI21_X1 U7475 ( .B1(n6508), .B2(n6523), .A(n6507), .ZN(U3207) );
  AOI22_X1 U7476 ( .A1(REIP_REG_25__SCAN_IN), .A2(n6521), .B1(
        ADDRESS_REG_24__SCAN_IN), .B2(n6509), .ZN(n6510) );
  OAI21_X1 U7477 ( .B1(n6511), .B2(n6523), .A(n6510), .ZN(U3208) );
  AOI22_X1 U7478 ( .A1(REIP_REG_26__SCAN_IN), .A2(n6521), .B1(
        ADDRESS_REG_25__SCAN_IN), .B2(n6565), .ZN(n6512) );
  OAI21_X1 U7479 ( .B1(n6513), .B2(n6523), .A(n6512), .ZN(U3209) );
  AOI22_X1 U7480 ( .A1(REIP_REG_27__SCAN_IN), .A2(n6521), .B1(
        ADDRESS_REG_26__SCAN_IN), .B2(n6565), .ZN(n6514) );
  OAI21_X1 U7481 ( .B1(n6516), .B2(n6523), .A(n6514), .ZN(U3210) );
  AOI22_X1 U7482 ( .A1(REIP_REG_29__SCAN_IN), .A2(n6517), .B1(
        ADDRESS_REG_27__SCAN_IN), .B2(n6565), .ZN(n6515) );
  OAI21_X1 U7483 ( .B1(n6516), .B2(n6519), .A(n6515), .ZN(U3211) );
  AOI22_X1 U7484 ( .A1(REIP_REG_30__SCAN_IN), .A2(n6517), .B1(
        ADDRESS_REG_28__SCAN_IN), .B2(n6565), .ZN(n6518) );
  OAI21_X1 U7485 ( .B1(n6520), .B2(n6519), .A(n6518), .ZN(U3212) );
  AOI22_X1 U7486 ( .A1(REIP_REG_30__SCAN_IN), .A2(n6521), .B1(
        ADDRESS_REG_29__SCAN_IN), .B2(n6565), .ZN(n6522) );
  OAI21_X1 U7487 ( .B1(n6524), .B2(n6523), .A(n6522), .ZN(U3213) );
  MUX2_X1 U7488 ( .A(BYTEENABLE_REG_3__SCAN_IN), .B(BE_N_REG_3__SCAN_IN), .S(
        n6565), .Z(U3445) );
  MUX2_X1 U7489 ( .A(BYTEENABLE_REG_2__SCAN_IN), .B(BE_N_REG_2__SCAN_IN), .S(
        n6565), .Z(U3446) );
  MUX2_X1 U7490 ( .A(BYTEENABLE_REG_1__SCAN_IN), .B(BE_N_REG_1__SCAN_IN), .S(
        n6565), .Z(U3447) );
  MUX2_X1 U7491 ( .A(BYTEENABLE_REG_0__SCAN_IN), .B(BE_N_REG_0__SCAN_IN), .S(
        n6565), .Z(U3448) );
  OAI21_X1 U7492 ( .B1(DATAWIDTH_REG_0__SCAN_IN), .B2(n6528), .A(n6526), .ZN(
        n6525) );
  INV_X1 U7493 ( .A(n6525), .ZN(U3451) );
  OAI21_X1 U7494 ( .B1(n6528), .B2(n6527), .A(n6526), .ZN(U3452) );
  OAI211_X1 U7495 ( .C1(n6717), .C2(n6531), .A(n6530), .B(n6529), .ZN(U3453)
         );
  OAI22_X1 U7496 ( .A1(n6534), .A2(n6542), .B1(n6533), .B2(n6532), .ZN(n6535)
         );
  MUX2_X1 U7497 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n6535), .S(n6540), 
        .Z(U3456) );
  OAI22_X1 U7498 ( .A1(n6537), .A2(n6542), .B1(INSTADDRPOINTER_REG_0__SCAN_IN), 
        .B2(n6536), .ZN(n6539) );
  OAI22_X1 U7499 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n6540), .B1(n6539), .B2(n6538), .ZN(n6541) );
  OAI21_X1 U7500 ( .B1(n6543), .B2(n6542), .A(n6541), .ZN(U3461) );
  AOI21_X1 U7501 ( .B1(REIP_REG_0__SCAN_IN), .B2(DATAWIDTH_REG_0__SCAN_IN), 
        .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6544) );
  AOI22_X1 U7502 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_0__SCAN_IN), .B1(
        n6544), .B2(n6573), .ZN(n6546) );
  INV_X1 U7503 ( .A(BYTEENABLE_REG_2__SCAN_IN), .ZN(n6545) );
  AOI22_X1 U7504 ( .A1(n6547), .A2(n6546), .B1(n6545), .B2(n6550), .ZN(U3468)
         );
  INV_X1 U7505 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n6551) );
  NOR2_X1 U7506 ( .A1(n6550), .A2(REIP_REG_1__SCAN_IN), .ZN(n6548) );
  AOI22_X1 U7507 ( .A1(n6551), .A2(n6550), .B1(n6549), .B2(n6548), .ZN(U3469)
         );
  NAND2_X1 U7508 ( .A1(n6565), .A2(W_R_N_REG_SCAN_IN), .ZN(n6552) );
  OAI21_X1 U7509 ( .B1(n6565), .B2(READREQUEST_REG_SCAN_IN), .A(n6552), .ZN(
        U3470) );
  AND2_X1 U7510 ( .A1(n6554), .A2(n6553), .ZN(n6555) );
  NOR4_X1 U7511 ( .A1(n6557), .A2(n6556), .A3(n5797), .A4(n6555), .ZN(n6564)
         );
  OAI211_X1 U7512 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n6559), .A(n6558), .B(
        STATE2_REG_2__SCAN_IN), .ZN(n6561) );
  AOI21_X1 U7513 ( .B1(n6561), .B2(STATE2_REG_0__SCAN_IN), .A(n6560), .ZN(
        n6563) );
  NAND2_X1 U7514 ( .A1(n6564), .A2(REQUESTPENDING_REG_SCAN_IN), .ZN(n6562) );
  OAI21_X1 U7515 ( .B1(n6564), .B2(n6563), .A(n6562), .ZN(U3472) );
  MUX2_X1 U7516 ( .A(MEMORYFETCH_REG_SCAN_IN), .B(M_IO_N_REG_SCAN_IN), .S(
        n6565), .Z(U3473) );
  AOI22_X1 U7517 ( .A1(n6567), .A2(keyinput50), .B1(keyinput51), .B2(n6731), 
        .ZN(n6566) );
  OAI221_X1 U7518 ( .B1(n6567), .B2(keyinput50), .C1(n6731), .C2(keyinput51), 
        .A(n6566), .ZN(n6578) );
  INV_X1 U7519 ( .A(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n6569) );
  AOI22_X1 U7520 ( .A1(n6569), .A2(keyinput46), .B1(keyinput30), .B2(n6732), 
        .ZN(n6568) );
  OAI221_X1 U7521 ( .B1(n6569), .B2(keyinput46), .C1(n6732), .C2(keyinput30), 
        .A(n6568), .ZN(n6577) );
  AOI22_X1 U7522 ( .A1(n6733), .A2(keyinput58), .B1(n6571), .B2(keyinput48), 
        .ZN(n6570) );
  OAI221_X1 U7523 ( .B1(n6733), .B2(keyinput58), .C1(n6571), .C2(keyinput48), 
        .A(n6570), .ZN(n6576) );
  AOI22_X1 U7524 ( .A1(n6574), .A2(keyinput13), .B1(keyinput11), .B2(n6573), 
        .ZN(n6572) );
  OAI221_X1 U7525 ( .B1(n6574), .B2(keyinput13), .C1(n6573), .C2(keyinput11), 
        .A(n6572), .ZN(n6575) );
  NOR4_X1 U7526 ( .A1(n6578), .A2(n6577), .A3(n6576), .A4(n6575), .ZN(n6623)
         );
  AOI22_X1 U7527 ( .A1(n6581), .A2(keyinput49), .B1(keyinput29), .B2(n6580), 
        .ZN(n6579) );
  OAI221_X1 U7528 ( .B1(n6581), .B2(keyinput49), .C1(n6580), .C2(keyinput29), 
        .A(n6579), .ZN(n6591) );
  AOI22_X1 U7529 ( .A1(n6716), .A2(keyinput9), .B1(n6583), .B2(keyinput44), 
        .ZN(n6582) );
  OAI221_X1 U7530 ( .B1(n6716), .B2(keyinput9), .C1(n6583), .C2(keyinput44), 
        .A(n6582), .ZN(n6590) );
  AOI22_X1 U7531 ( .A1(n4312), .A2(keyinput45), .B1(n6723), .B2(keyinput57), 
        .ZN(n6584) );
  OAI221_X1 U7532 ( .B1(n4312), .B2(keyinput45), .C1(n6723), .C2(keyinput57), 
        .A(n6584), .ZN(n6589) );
  INV_X1 U7533 ( .A(DATAI_21_), .ZN(n6585) );
  XOR2_X1 U7534 ( .A(n6585), .B(keyinput5), .Z(n6587) );
  XNOR2_X1 U7535 ( .A(INSTQUEUE_REG_7__3__SCAN_IN), .B(keyinput19), .ZN(n6586)
         );
  NAND2_X1 U7536 ( .A1(n6587), .A2(n6586), .ZN(n6588) );
  NOR4_X1 U7537 ( .A1(n6591), .A2(n6590), .A3(n6589), .A4(n6588), .ZN(n6622)
         );
  INV_X1 U7538 ( .A(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n6709) );
  AOI22_X1 U7539 ( .A1(n6709), .A2(keyinput22), .B1(keyinput55), .B2(n6593), 
        .ZN(n6592) );
  OAI221_X1 U7540 ( .B1(n6709), .B2(keyinput22), .C1(n6593), .C2(keyinput55), 
        .A(n6592), .ZN(n6605) );
  INV_X1 U7541 ( .A(LWORD_REG_6__SCAN_IN), .ZN(n6595) );
  AOI22_X1 U7542 ( .A1(n6596), .A2(keyinput24), .B1(keyinput6), .B2(n6595), 
        .ZN(n6594) );
  OAI221_X1 U7543 ( .B1(n6596), .B2(keyinput24), .C1(n6595), .C2(keyinput6), 
        .A(n6594), .ZN(n6604) );
  AOI22_X1 U7544 ( .A1(n6599), .A2(keyinput54), .B1(n6598), .B2(keyinput40), 
        .ZN(n6597) );
  OAI221_X1 U7545 ( .B1(n6599), .B2(keyinput54), .C1(n6598), .C2(keyinput40), 
        .A(n6597), .ZN(n6603) );
  XOR2_X1 U7546 ( .A(n4432), .B(keyinput37), .Z(n6601) );
  XNOR2_X1 U7547 ( .A(INSTQUEUE_REG_1__1__SCAN_IN), .B(keyinput21), .ZN(n6600)
         );
  NAND2_X1 U7548 ( .A1(n6601), .A2(n6600), .ZN(n6602) );
  NOR4_X1 U7549 ( .A1(n6605), .A2(n6604), .A3(n6603), .A4(n6602), .ZN(n6621)
         );
  INV_X1 U7550 ( .A(DATAO_REG_2__SCAN_IN), .ZN(n6607) );
  AOI22_X1 U7551 ( .A1(n6608), .A2(keyinput62), .B1(keyinput43), .B2(n6607), 
        .ZN(n6606) );
  OAI221_X1 U7552 ( .B1(n6608), .B2(keyinput62), .C1(n6607), .C2(keyinput43), 
        .A(n6606), .ZN(n6619) );
  INV_X1 U7553 ( .A(DATAI_19_), .ZN(n6704) );
  AOI22_X1 U7554 ( .A1(n6610), .A2(keyinput10), .B1(keyinput27), .B2(n6704), 
        .ZN(n6609) );
  OAI221_X1 U7555 ( .B1(n6610), .B2(keyinput10), .C1(n6704), .C2(keyinput27), 
        .A(n6609), .ZN(n6618) );
  INV_X1 U7556 ( .A(UWORD_REG_3__SCAN_IN), .ZN(n6613) );
  AOI22_X1 U7557 ( .A1(n6613), .A2(keyinput17), .B1(n6612), .B2(keyinput25), 
        .ZN(n6611) );
  OAI221_X1 U7558 ( .B1(n6613), .B2(keyinput17), .C1(n6612), .C2(keyinput25), 
        .A(n6611), .ZN(n6617) );
  XNOR2_X1 U7559 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(keyinput59), .ZN(
        n6615) );
  XNOR2_X1 U7560 ( .A(INSTQUEUE_REG_5__5__SCAN_IN), .B(keyinput38), .ZN(n6614)
         );
  NAND2_X1 U7561 ( .A1(n6615), .A2(n6614), .ZN(n6616) );
  NOR4_X1 U7562 ( .A1(n6619), .A2(n6618), .A3(n6617), .A4(n6616), .ZN(n6620)
         );
  NAND4_X1 U7563 ( .A1(n6623), .A2(n6622), .A3(n6621), .A4(n6620), .ZN(n6687)
         );
  AOI22_X1 U7564 ( .A1(n6626), .A2(keyinput15), .B1(n6625), .B2(keyinput3), 
        .ZN(n6624) );
  OAI221_X1 U7565 ( .B1(n6626), .B2(keyinput15), .C1(n6625), .C2(keyinput3), 
        .A(n6624), .ZN(n6630) );
  XNOR2_X1 U7566 ( .A(n6627), .B(keyinput8), .ZN(n6629) );
  XOR2_X1 U7567 ( .A(INSTQUEUE_REG_5__6__SCAN_IN), .B(keyinput63), .Z(n6628)
         );
  OR3_X1 U7568 ( .A1(n6630), .A2(n6629), .A3(n6628), .ZN(n6638) );
  AOI22_X1 U7569 ( .A1(n6725), .A2(keyinput20), .B1(keyinput61), .B2(n6632), 
        .ZN(n6631) );
  OAI221_X1 U7570 ( .B1(n6725), .B2(keyinput20), .C1(n6632), .C2(keyinput61), 
        .A(n6631), .ZN(n6637) );
  INV_X1 U7571 ( .A(DATAI_31_), .ZN(n6634) );
  AOI22_X1 U7572 ( .A1(n6635), .A2(keyinput28), .B1(n6634), .B2(keyinput16), 
        .ZN(n6633) );
  OAI221_X1 U7573 ( .B1(n6635), .B2(keyinput28), .C1(n6634), .C2(keyinput16), 
        .A(n6633), .ZN(n6636) );
  NOR3_X1 U7574 ( .A1(n6638), .A2(n6637), .A3(n6636), .ZN(n6685) );
  INV_X1 U7575 ( .A(ADDRESS_REG_19__SCAN_IN), .ZN(n6640) );
  AOI22_X1 U7576 ( .A1(n6641), .A2(keyinput14), .B1(keyinput53), .B2(n6640), 
        .ZN(n6639) );
  OAI221_X1 U7577 ( .B1(n6641), .B2(keyinput14), .C1(n6640), .C2(keyinput53), 
        .A(n6639), .ZN(n6654) );
  AOI22_X1 U7578 ( .A1(n6644), .A2(keyinput60), .B1(keyinput47), .B2(n6643), 
        .ZN(n6642) );
  OAI221_X1 U7579 ( .B1(n6644), .B2(keyinput60), .C1(n6643), .C2(keyinput47), 
        .A(n6642), .ZN(n6653) );
  AOI22_X1 U7580 ( .A1(n6647), .A2(keyinput12), .B1(n6646), .B2(keyinput52), 
        .ZN(n6645) );
  OAI221_X1 U7581 ( .B1(n6647), .B2(keyinput12), .C1(n6646), .C2(keyinput52), 
        .A(n6645), .ZN(n6652) );
  AOI22_X1 U7582 ( .A1(n6650), .A2(keyinput41), .B1(keyinput35), .B2(n6649), 
        .ZN(n6648) );
  OAI221_X1 U7583 ( .B1(n6650), .B2(keyinput41), .C1(n6649), .C2(keyinput35), 
        .A(n6648), .ZN(n6651) );
  NOR4_X1 U7584 ( .A1(n6654), .A2(n6653), .A3(n6652), .A4(n6651), .ZN(n6684)
         );
  AOI22_X1 U7585 ( .A1(n6657), .A2(keyinput26), .B1(keyinput18), .B2(n6656), 
        .ZN(n6655) );
  OAI221_X1 U7586 ( .B1(n6657), .B2(keyinput26), .C1(n6656), .C2(keyinput18), 
        .A(n6655), .ZN(n6669) );
  INV_X1 U7587 ( .A(UWORD_REG_1__SCAN_IN), .ZN(n6659) );
  AOI22_X1 U7588 ( .A1(n6659), .A2(keyinput42), .B1(n6724), .B2(keyinput56), 
        .ZN(n6658) );
  OAI221_X1 U7589 ( .B1(n6659), .B2(keyinput42), .C1(n6724), .C2(keyinput56), 
        .A(n6658), .ZN(n6668) );
  INV_X1 U7590 ( .A(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n6662) );
  AOI22_X1 U7591 ( .A1(n6662), .A2(keyinput36), .B1(n6661), .B2(keyinput31), 
        .ZN(n6660) );
  OAI221_X1 U7592 ( .B1(n6662), .B2(keyinput36), .C1(n6661), .C2(keyinput31), 
        .A(n6660), .ZN(n6667) );
  XOR2_X1 U7593 ( .A(n6663), .B(keyinput4), .Z(n6665) );
  XNOR2_X1 U7594 ( .A(INSTQUEUE_REG_9__4__SCAN_IN), .B(keyinput1), .ZN(n6664)
         );
  NAND2_X1 U7595 ( .A1(n6665), .A2(n6664), .ZN(n6666) );
  NOR4_X1 U7596 ( .A1(n6669), .A2(n6668), .A3(n6667), .A4(n6666), .ZN(n6683)
         );
  AOI22_X1 U7597 ( .A1(n3899), .A2(keyinput0), .B1(n6671), .B2(keyinput34), 
        .ZN(n6670) );
  OAI221_X1 U7598 ( .B1(n3899), .B2(keyinput0), .C1(n6671), .C2(keyinput34), 
        .A(n6670), .ZN(n6681) );
  AOI22_X1 U7599 ( .A1(n6674), .A2(keyinput39), .B1(n6673), .B2(keyinput2), 
        .ZN(n6672) );
  OAI221_X1 U7600 ( .B1(n6674), .B2(keyinput39), .C1(n6673), .C2(keyinput2), 
        .A(n6672), .ZN(n6680) );
  AOI22_X1 U7601 ( .A1(n6726), .A2(keyinput33), .B1(n6710), .B2(keyinput7), 
        .ZN(n6675) );
  OAI221_X1 U7602 ( .B1(n6726), .B2(keyinput33), .C1(n6710), .C2(keyinput7), 
        .A(n6675), .ZN(n6679) );
  AOI22_X1 U7603 ( .A1(n6677), .A2(keyinput23), .B1(keyinput32), .B2(n6717), 
        .ZN(n6676) );
  OAI221_X1 U7604 ( .B1(n6677), .B2(keyinput23), .C1(n6717), .C2(keyinput32), 
        .A(n6676), .ZN(n6678) );
  NOR4_X1 U7605 ( .A1(n6681), .A2(n6680), .A3(n6679), .A4(n6678), .ZN(n6682)
         );
  NAND4_X1 U7606 ( .A1(n6685), .A2(n6684), .A3(n6683), .A4(n6682), .ZN(n6686)
         );
  NOR2_X1 U7607 ( .A1(n6687), .A2(n6686), .ZN(n6744) );
  INV_X1 U7608 ( .A(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n6692) );
  OAI21_X1 U7609 ( .B1(REIP_REG_17__SCAN_IN), .B2(n6689), .A(n6688), .ZN(n6690) );
  OAI211_X1 U7610 ( .C1(n6693), .C2(n6692), .A(n6691), .B(n6690), .ZN(n6694)
         );
  AOI21_X1 U7611 ( .B1(EBX_REG_17__SCAN_IN), .B2(n6695), .A(n6694), .ZN(n6701)
         );
  AOI22_X1 U7612 ( .A1(n6699), .A2(n6698), .B1(n6697), .B2(n6696), .ZN(n6700)
         );
  OAI211_X1 U7613 ( .C1(n6703), .C2(n6702), .A(n6701), .B(n6700), .ZN(n6742)
         );
  NAND4_X1 U7614 ( .A1(EBX_REG_29__SCAN_IN), .A2(UWORD_REG_12__SCAN_IN), .A3(
        DATAO_REG_2__SCAN_IN), .A4(n6704), .ZN(n6708) );
  NAND4_X1 U7615 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        LWORD_REG_15__SCAN_IN), .A3(DATAO_REG_10__SCAN_IN), .A4(
        ADDRESS_REG_8__SCAN_IN), .ZN(n6707) );
  NAND4_X1 U7616 ( .A1(DATAI_31_), .A2(ADDRESS_REG_19__SCAN_IN), .A3(
        UWORD_REG_0__SCAN_IN), .A4(DATAWIDTH_REG_15__SCAN_IN), .ZN(n6706) );
  NAND4_X1 U7617 ( .A1(INSTADDRPOINTER_REG_29__SCAN_IN), .A2(DATAI_7_), .A3(
        UWORD_REG_1__SCAN_IN), .A4(DATAO_REG_23__SCAN_IN), .ZN(n6705) );
  NOR4_X1 U7618 ( .A1(n6708), .A2(n6707), .A3(n6706), .A4(n6705), .ZN(n6722)
         );
  NOR4_X1 U7619 ( .A1(INSTQUEUE_REG_6__0__SCAN_IN), .A2(
        INSTQUEUE_REG_5__6__SCAN_IN), .A3(n6710), .A4(n6709), .ZN(n6721) );
  NOR3_X1 U7620 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n6711), .A3(
        INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n6712) );
  NAND3_X1 U7621 ( .A1(n6712), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .A3(n6662), 
        .ZN(n6719) );
  INV_X1 U7622 ( .A(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n6715) );
  INV_X1 U7623 ( .A(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n6714) );
  INV_X1 U7624 ( .A(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n6713) );
  NAND4_X1 U7625 ( .A1(n6715), .A2(n6714), .A3(n6583), .A4(n6713), .ZN(n6718)
         );
  NOR4_X1 U7626 ( .A1(n6719), .A2(n6718), .A3(n6717), .A4(n6716), .ZN(n6720)
         );
  NAND3_X1 U7627 ( .A1(n6722), .A2(n6721), .A3(n6720), .ZN(n6740) );
  NOR4_X1 U7628 ( .A1(EBX_REG_14__SCAN_IN), .A2(EBX_REG_8__SCAN_IN), .A3(
        PHYADDRPOINTER_REG_9__SCAN_IN), .A4(n6723), .ZN(n6730) );
  NOR4_X1 U7629 ( .A1(INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .A3(EBX_REG_4__SCAN_IN), .A4(
        REIP_REG_1__SCAN_IN), .ZN(n6729) );
  NOR4_X1 U7630 ( .A1(EAX_REG_16__SCAN_IN), .A2(REIP_REG_15__SCAN_IN), .A3(
        REIP_REG_12__SCAN_IN), .A4(n6724), .ZN(n6728) );
  NOR4_X1 U7631 ( .A1(EAX_REG_14__SCAN_IN), .A2(EAX_REG_0__SCAN_IN), .A3(n6726), .A4(n6725), .ZN(n6727) );
  NAND4_X1 U7632 ( .A1(n6730), .A2(n6729), .A3(n6728), .A4(n6727), .ZN(n6739)
         );
  NOR4_X1 U7633 ( .A1(EAX_REG_22__SCAN_IN), .A2(DATAI_21_), .A3(n6732), .A4(
        n6731), .ZN(n6737) );
  NOR4_X1 U7634 ( .A1(DATAO_REG_16__SCAN_IN), .A2(DATAO_REG_15__SCAN_IN), .A3(
        UWORD_REG_11__SCAN_IN), .A4(n6733), .ZN(n6736) );
  NOR4_X1 U7635 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(FLUSH_REG_SCAN_IN), .A3(
        LWORD_REG_6__SCAN_IN), .A4(UWORD_REG_3__SCAN_IN), .ZN(n6735) );
  NOR4_X1 U7636 ( .A1(EBX_REG_23__SCAN_IN), .A2(EAX_REG_18__SCAN_IN), .A3(
        DATAO_REG_28__SCAN_IN), .A4(DATAI_0_), .ZN(n6734) );
  NAND4_X1 U7637 ( .A1(n6737), .A2(n6736), .A3(n6735), .A4(n6734), .ZN(n6738)
         );
  NOR3_X1 U7638 ( .A1(n6740), .A2(n6739), .A3(n6738), .ZN(n6741) );
  XNOR2_X1 U7639 ( .A(n6742), .B(n6741), .ZN(n6743) );
  XNOR2_X1 U7640 ( .A(n6744), .B(n6743), .ZN(U2810) );
  AND4_X1 U3857 ( .A1(n3001), .A2(n3000), .A3(n2999), .A4(n2998), .ZN(n3012)
         );
  AND4_X1 U3942 ( .A1(n3093), .A2(n3092), .A3(n3091), .A4(n3090), .ZN(n3100)
         );
  INV_X1 U3414 ( .A(n3261), .ZN(n4223) );
  AOI21_X1 U4655 ( .B1(n4837), .B2(n3166), .A(n6661), .ZN(n4397) );
  BUF_X1 U3492 ( .A(n4174), .Z(n4156) );
  OAI21_X1 U4027 ( .B1(n3293), .B2(n6400), .A(n3175), .ZN(n3217) );
  AND4_X1 U3419 ( .A1(n3005), .A2(n3004), .A3(n3003), .A4(n3002), .ZN(n3011)
         );
  CLKBUF_X1 U3425 ( .A(n3365), .Z(n4457) );
  OR2_X2 U3432 ( .A1(n3059), .A2(n3058), .ZN(n4473) );
  CLKBUF_X1 U3436 ( .A(n3694), .Z(n6403) );
  CLKBUF_X1 U3442 ( .A(n5403), .Z(n5447) );
  INV_X1 U34740 ( .A(n3655), .ZN(n3166) );
  CLKBUF_X1 U3533 ( .A(n4199), .Z(n5390) );
  CLKBUF_X1 U3582 ( .A(n3201), .Z(n3203) );
  CLKBUF_X1 U3611 ( .A(n3517), .Z(n4494) );
  CLKBUF_X1 U3618 ( .A(n3715), .Z(n4743) );
  CLKBUF_X1 U3862 ( .A(n5062), .Z(n5942) );
  XNOR2_X1 U3910 ( .A(n3203), .B(n3202), .ZN(n5785) );
endmodule

