

module b14_C_2inp_gates_syn ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, 
        REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, 
        REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, 
        REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, 
        REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, 
        REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, 
        REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, 
        REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, 
        IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, 
        IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, 
        IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, 
        IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, 
        IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, 
        IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, 
        IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, 
        IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, 
        IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, 
        IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, 
        IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, 
        D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, 
        D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, 
        D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, 
        D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, 
        D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, 
        D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, 
        D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, 
        D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, 
        D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, 
        D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, 
        REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, 
        REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, 
        REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, 
        REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, 
        REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, 
        REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, 
        REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, 
        REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, 
        REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, 
        REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, 
        REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, 
        REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, 
        REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, 
        REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, 
        REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, 
        REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, 
        REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, 
        REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, 
        REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, 
        REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, 
        REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, 
        REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, 
        REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, 
        REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, 
        REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, 
        REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, 
        REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, 
        REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, 
        REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, 
        REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, 
        REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, 
        REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, 
        ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, 
        ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, 
        ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, 
        ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, 
        ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, 
        ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, 
        ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, 
        REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, 
        REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, U3352, U3351, U3350, U3349, 
        U3348, U3347, U3346, U3345, U3344, U3343, U3342, U3341, U3340, U3339, 
        U3338, U3337, U3336, U3335, U3334, U3333, U3332, U3331, U3330, U3329, 
        U3328, U3327, U3326, U3325, U3324, U3323, U3322, U3321, U3458, U3459, 
        U3320, U3319, U3318, U3317, U3316, U3315, U3314, U3313, U3312, U3311, 
        U3310, U3309, U3308, U3307, U3306, U3305, U3304, U3303, U3302, U3301, 
        U3300, U3299, U3298, U3297, U3296, U3295, U3294, U3293, U3292, U3291, 
        U3467, U3469, U3471, U3473, U3475, U3477, U3479, U3481, U3483, U3485, 
        U3487, U3489, U3491, U3493, U3495, U3497, U3499, U3501, U3503, U3505, 
        U3506, U3507, U3508, U3509, U3510, U3511, U3512, U3513, U3514, U3515, 
        U3516, U3517, U3518, U3519, U3520, U3521, U3522, U3523, U3524, U3525, 
        U3526, U3527, U3528, U3529, U3530, U3531, U3532, U3533, U3534, U3535, 
        U3536, U3537, U3538, U3539, U3540, U3541, U3542, U3543, U3544, U3545, 
        U3546, U3547, U3548, U3549, U3290, U3289, U3288, U3287, U3286, U3285, 
        U3284, U3283, U3282, U3281, U3280, U3279, U3278, U3277, U3276, U3275, 
        U3274, U3273, U3272, U3271, U3270, U3269, U3268, U3267, U3266, U3265, 
        U3264, U3263, U3262, U3354, U3261, U3260, U3259, U3258, U3257, U3256, 
        U3255, U3254, U3253, U3252, U3251, U3250, U3249, U3248, U3247, U3246, 
        U3245, U3244, U3243, U3242, U3241, U3240, U3550, U3551, U3552, U3553, 
        U3554, U3555, U3556, U3557, U3558, U3559, U3560, U3561, U3562, U3563, 
        U3564, U3565, U3566, U3567, U3568, U3569, U3570, U3571, U3572, U3573, 
        U3574, U3575, U3576, U3577, U3578, U3579, U3580, U3581, U3239, U3238, 
        U3237, U3236, U3235, U3234, U3233, U3232, U3231, U3230, U3229, U3228, 
        U3227, U3226, U3225, U3224, U3223, U3222, U3221, U3220, U3219, U3218, 
        U3217, U3216, U3215, U3214, U3213, U3212, U3211, U3210, U3149, U3148, 
        U4043, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, 
        keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, 
        keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, 
        keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, 
        keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, 
        keyinput29, keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, 
        keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, 
        keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, 
        keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, 
        keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, 
        keyinput59, keyinput60, keyinput61, keyinput62, keyinput63, keyinput64, 
        keyinput65, keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, 
        keyinput71, keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, 
        keyinput77, keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, 
        keyinput83, keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, 
        keyinput89, keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, 
        keyinput95, keyinput96, keyinput97, keyinput98, keyinput99, 
        keyinput100, keyinput101, keyinput102, keyinput103, keyinput104, 
        keyinput105, keyinput106, keyinput107, keyinput108, keyinput109, 
        keyinput110, keyinput111, keyinput112, keyinput113, keyinput114, 
        keyinput115, keyinput116, keyinput117, keyinput118, keyinput119, 
        keyinput120, keyinput121, keyinput122, keyinput123, keyinput124, 
        keyinput125, keyinput126, keyinput127 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
         REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
         REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
         REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
         REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
         REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
         REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
         REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
         IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
         IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
         IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
         IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
         IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
         IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
         IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
         IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
         IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
         IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
         IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
         D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
         D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN,
         D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
         D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
         D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
         D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
         D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
         D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
         D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
         D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
         D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
         REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
         REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
         REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
         REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
         REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
         REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
         REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
         REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
         REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
         REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
         REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
         REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
         REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
         REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
         REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
         REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
         REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
         REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
         REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
         REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
         REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
         REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
         REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
         REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
         REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
         REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
         REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
         REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
         REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
         REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
         REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
         REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
         ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
         ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
         ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
         ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
         ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
         ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
         DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
         DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
         DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
         DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
         DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
         DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
         DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
         DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
         DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
         DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
         DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
         REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
         REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
         REG3_REG_22__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141,
         n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151,
         n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161,
         n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171,
         n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181,
         n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191,
         n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201,
         n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211,
         n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221,
         n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231,
         n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241,
         n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251,
         n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261,
         n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271,
         n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281,
         n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291,
         n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301,
         n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311,
         n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321,
         n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331,
         n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341,
         n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351,
         n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361,
         n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371,
         n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381,
         n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391,
         n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401,
         n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411,
         n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421,
         n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431,
         n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441,
         n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451,
         n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461,
         n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471,
         n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481,
         n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491,
         n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501,
         n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511,
         n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521,
         n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531,
         n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541,
         n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551,
         n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561,
         n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571,
         n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581,
         n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591,
         n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601,
         n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611,
         n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621,
         n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631,
         n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641,
         n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651,
         n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661,
         n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671,
         n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681,
         n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691,
         n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701,
         n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711,
         n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721,
         n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731,
         n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741,
         n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751,
         n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761,
         n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771,
         n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781,
         n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791,
         n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801,
         n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811,
         n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821,
         n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831,
         n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841,
         n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851,
         n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861,
         n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871,
         n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881,
         n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891,
         n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901,
         n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911,
         n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921,
         n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931,
         n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941,
         n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951,
         n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961,
         n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971,
         n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981,
         n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991,
         n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001,
         n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011,
         n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021,
         n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031,
         n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041,
         n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051,
         n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061,
         n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071,
         n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081,
         n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091,
         n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101,
         n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111,
         n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121,
         n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131,
         n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141,
         n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151,
         n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161,
         n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171,
         n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181,
         n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191,
         n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201,
         n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211,
         n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221,
         n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231,
         n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241,
         n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251,
         n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261,
         n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271,
         n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281,
         n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291,
         n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301,
         n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311,
         n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321,
         n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331,
         n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341,
         n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351,
         n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361,
         n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371,
         n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381,
         n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391,
         n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401,
         n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411,
         n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421,
         n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431,
         n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441,
         n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451,
         n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461,
         n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471,
         n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481,
         n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491,
         n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501,
         n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511,
         n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521,
         n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531,
         n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541,
         n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551,
         n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561,
         n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571,
         n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581,
         n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591,
         n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601,
         n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611,
         n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621,
         n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631,
         n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641,
         n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651,
         n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661,
         n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671,
         n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681,
         n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691,
         n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701,
         n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711,
         n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721,
         n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731,
         n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741,
         n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751,
         n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761,
         n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771,
         n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781,
         n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791,
         n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801,
         n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811,
         n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821,
         n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831,
         n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841,
         n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851,
         n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861,
         n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871,
         n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881,
         n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891,
         n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901,
         n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911,
         n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921,
         n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931,
         n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941,
         n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951,
         n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961,
         n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971,
         n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981,
         n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991,
         n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001,
         n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011,
         n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021,
         n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031,
         n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041,
         n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051,
         n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061,
         n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071,
         n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081,
         n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091,
         n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101,
         n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111,
         n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121,
         n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131,
         n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141,
         n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151,
         n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161,
         n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171,
         n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181,
         n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191,
         n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201,
         n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211,
         n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221,
         n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231,
         n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241,
         n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251,
         n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261,
         n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271,
         n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281,
         n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291,
         n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301,
         n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311,
         n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321,
         n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331,
         n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341,
         n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351,
         n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361,
         n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371,
         n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381,
         n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391,
         n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401,
         n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411,
         n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421,
         n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431,
         n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441,
         n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451,
         n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461,
         n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471,
         n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481,
         n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491,
         n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501,
         n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511,
         n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521,
         n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531,
         n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541,
         n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551,
         n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561,
         n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571,
         n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581,
         n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591,
         n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601,
         n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611,
         n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621,
         n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631,
         n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641,
         n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651,
         n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661,
         n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671,
         n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681,
         n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691,
         n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701,
         n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711,
         n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721,
         n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731,
         n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741,
         n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751,
         n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761,
         n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771,
         n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781,
         n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791,
         n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801,
         n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811,
         n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821,
         n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831,
         n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841,
         n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851,
         n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861,
         n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871,
         n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881,
         n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891,
         n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901,
         n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911,
         n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921,
         n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931,
         n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941,
         n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951,
         n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961,
         n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971,
         n4972, n4973, n4974, n4975, n4976, n4977, n4978;

  CLKBUF_X1 U2374 ( .A(n2535), .Z(n2135) );
  INV_X1 U2375 ( .A(n4288), .ZN(n3918) );
  INV_X1 U2376 ( .A(n2414), .ZN(n2916) );
  INV_X1 U2377 ( .A(n2991), .ZN(n3629) );
  CLKBUF_X2 U2378 ( .A(n2535), .Z(n2136) );
  CLKBUF_X1 U2379 ( .A(n2493), .Z(n2132) );
  CLKBUF_X1 U2380 ( .A(n2470), .Z(n2137) );
  NAND4_X2 U2381 ( .A1(n2460), .A2(n2459), .A3(n2458), .A4(n2457), .ZN(n2990)
         );
  NAND2_X1 U2382 ( .A1(n2469), .A2(n2470), .ZN(n3033) );
  INV_X1 U2383 ( .A(n2535), .ZN(n2138) );
  OR2_X1 U2384 ( .A1(n3007), .A2(n3843), .ZN(n3925) );
  INV_X1 U2385 ( .A(n3033), .ZN(n3500) );
  INV_X2 U2386 ( .A(IR_REG_15__SCAN_IN), .ZN(n3154) );
  XNOR2_X1 U2388 ( .A(n4353), .B(n4344), .ZN(n4874) );
  XNOR2_X1 U2389 ( .A(n2244), .B(n3413), .ZN(n3424) );
  INV_X1 U2390 ( .A(n4908), .ZN(n4485) );
  OR3_X1 U2391 ( .A1(n3531), .A2(n2469), .A3(n4937), .ZN(n4647) );
  NAND4_X1 U2392 ( .A1(n2664), .A2(n2663), .A3(n2662), .A4(n2661), .ZN(n4288)
         );
  INV_X2 U2393 ( .A(n3499), .ZN(n4908) );
  NAND2_X2 U2394 ( .A1(n4827), .A2(n2243), .ZN(n2239) );
  NAND4_X2 U2395 ( .A1(n2415), .A2(n2445), .A3(n2515), .A4(n2530), .ZN(n2550)
         );
  NAND2_X2 U2396 ( .A1(n2157), .A2(IR_REG_31__SCAN_IN), .ZN(n2464) );
  XNOR2_X2 U2397 ( .A(n3400), .B(n3394), .ZN(n3399) );
  OR2_X4 U2398 ( .A1(n3118), .A2(n2456), .ZN(n2509) );
  XNOR2_X2 U2399 ( .A(n2451), .B(n2452), .ZN(n2456) );
  NAND2_X2 U2400 ( .A1(n4016), .A2(IR_REG_31__SCAN_IN), .ZN(n2454) );
  XNOR2_X2 U2401 ( .A(n3771), .B(n3773), .ZN(n3775) );
  AND2_X1 U2402 ( .A1(n4180), .A2(n3842), .ZN(n3843) );
  NAND4_X1 U2403 ( .A1(n2639), .A2(n2638), .A3(n2637), .A4(n2636), .ZN(n4289)
         );
  NAND4_X2 U2404 ( .A1(n2548), .A2(n2547), .A3(n2546), .A4(n2545), .ZN(n3830)
         );
  INV_X4 U2405 ( .A(n2849), .ZN(n2914) );
  NAND4_X2 U2406 ( .A1(n2405), .A2(n2497), .A3(n2496), .A4(n2495), .ZN(n3643)
         );
  INV_X1 U2407 ( .A(n2133), .ZN(n2898) );
  INV_X2 U2408 ( .A(n2494), .ZN(n3465) );
  XNOR2_X1 U2409 ( .A(n2435), .B(IR_REG_20__SCAN_IN), .ZN(n2470) );
  INV_X2 U2410 ( .A(IR_REG_7__SCAN_IN), .ZN(n2609) );
  OR2_X1 U2411 ( .A1(n4021), .A2(n4020), .ZN(n2286) );
  OAI21_X1 U2412 ( .B1(n4100), .B2(n4102), .A(n4101), .ZN(n4021) );
  NAND2_X1 U2413 ( .A1(n2342), .A2(n2340), .ZN(n2343) );
  NAND2_X1 U2414 ( .A1(n2151), .A2(n2289), .ZN(n3573) );
  AND2_X1 U2415 ( .A1(n3989), .A2(n4645), .ZN(n2406) );
  OR2_X1 U2416 ( .A1(n3546), .A2(n2249), .ZN(n2246) );
  AOI21_X1 U2417 ( .B1(n2326), .B2(n2142), .A(n2325), .ZN(n2324) );
  AOI21_X1 U2418 ( .B1(n2160), .B2(n2378), .A(n3015), .ZN(n2374) );
  AND2_X1 U2419 ( .A1(n3710), .A2(n3002), .ZN(n3001) );
  AND2_X1 U2420 ( .A1(n3724), .A2(n3000), .ZN(n3002) );
  AOI21_X1 U2421 ( .B1(n2328), .B2(n2142), .A(n2171), .ZN(n2327) );
  NAND2_X1 U2422 ( .A1(n4243), .A2(n4239), .ZN(n4180) );
  NAND2_X1 U2423 ( .A1(n3035), .A2(n4206), .ZN(n3639) );
  NAND2_X1 U2424 ( .A1(n4214), .A2(n4211), .ZN(n4171) );
  NAND3_X1 U2425 ( .A1(n2240), .A2(n2172), .A3(n2239), .ZN(n2244) );
  NAND2_X1 U2426 ( .A1(n3039), .A2(n4225), .ZN(n3716) );
  NAND4_X1 U2427 ( .A1(n2623), .A2(n2622), .A3(n2621), .A4(n2620), .ZN(n3811)
         );
  NAND2_X2 U2428 ( .A1(n2471), .A2(n2137), .ZN(n3076) );
  NAND2_X1 U2429 ( .A1(n2569), .A2(n2568), .ZN(n4291) );
  NAND2_X1 U2430 ( .A1(n4290), .A2(n3700), .ZN(n4225) );
  OR2_X1 U2431 ( .A1(n4290), .A2(n3700), .ZN(n3039) );
  NAND4_X1 U2432 ( .A1(n2608), .A2(n2607), .A3(n2606), .A4(n2605), .ZN(n3796)
         );
  NAND4_X1 U2433 ( .A1(n2689), .A2(n2688), .A3(n2687), .A4(n2686), .ZN(n4287)
         );
  INV_X1 U2434 ( .A(n3537), .ZN(n3636) );
  AND3_X1 U2435 ( .A1(n2567), .A2(n2566), .A3(n2565), .ZN(n2568) );
  NAND4_X2 U2436 ( .A1(n2591), .A2(n2590), .A3(n2589), .A4(n2588), .ZN(n4290)
         );
  AND2_X2 U2437 ( .A1(n2962), .A2(n3033), .ZN(n2414) );
  AND2_X2 U2438 ( .A1(n2964), .A2(n3033), .ZN(n2849) );
  NAND2_X1 U2439 ( .A1(n2972), .A2(REG1_REG_3__SCAN_IN), .ZN(n2514) );
  INV_X2 U2440 ( .A(n2518), .ZN(n3085) );
  NAND2_X1 U2441 ( .A1(n2430), .A2(n4805), .ZN(n2962) );
  XNOR2_X1 U2442 ( .A(n2440), .B(IR_REG_26__SCAN_IN), .ZN(n4805) );
  NOR2_X1 U2443 ( .A1(n2927), .A2(n2428), .ZN(n2430) );
  OR2_X1 U2444 ( .A1(n2440), .A2(IR_REG_27__SCAN_IN), .ZN(n2441) );
  XNOR2_X1 U2445 ( .A(n2465), .B(n2466), .ZN(n4376) );
  NAND2_X1 U2446 ( .A1(n2196), .A2(IR_REG_31__SCAN_IN), .ZN(n2498) );
  NAND2_X1 U2447 ( .A1(n2443), .A2(n2445), .ZN(n2196) );
  NAND3_X1 U2448 ( .A1(n3207), .A2(n2609), .A3(n2592), .ZN(n3128) );
  INV_X1 U2449 ( .A(IR_REG_3__SCAN_IN), .ZN(n2530) );
  INV_X1 U2450 ( .A(IR_REG_25__SCAN_IN), .ZN(n2447) );
  INV_X1 U2451 ( .A(IR_REG_28__SCAN_IN), .ZN(n2969) );
  INV_X1 U2452 ( .A(IR_REG_11__SCAN_IN), .ZN(n2690) );
  INV_X1 U2453 ( .A(IR_REG_26__SCAN_IN), .ZN(n2448) );
  INV_X1 U2454 ( .A(IR_REG_6__SCAN_IN), .ZN(n2592) );
  NOR2_X1 U2455 ( .A1(IR_REG_20__SCAN_IN), .A2(IR_REG_19__SCAN_IN), .ZN(n2431)
         );
  INV_X1 U2456 ( .A(IR_REG_13__SCAN_IN), .ZN(n2714) );
  INV_X1 U2457 ( .A(IR_REG_14__SCAN_IN), .ZN(n2730) );
  INV_X1 U2458 ( .A(IR_REG_27__SCAN_IN), .ZN(n3087) );
  NOR2_X1 U2459 ( .A1(IR_REG_16__SCAN_IN), .A2(IR_REG_9__SCAN_IN), .ZN(n2417)
         );
  OR2_X1 U2460 ( .A1(n2433), .A2(n2763), .ZN(n2465) );
  OAI21_X1 U2461 ( .B1(n4419), .B2(n3031), .A(n2345), .ZN(n4390) );
  NAND2_X2 U2462 ( .A1(n3573), .A2(n2600), .ZN(n3522) );
  NAND2_X1 U2464 ( .A1(n4804), .A2(n3118), .ZN(n2493) );
  NAND3_X2 U2465 ( .A1(n2422), .A2(n2421), .A3(n2423), .ZN(n2764) );
  INV_X1 U2466 ( .A(n2525), .ZN(n2134) );
  AND2_X4 U2467 ( .A1(n2455), .A2(n2456), .ZN(n2525) );
  OAI211_X2 U2468 ( .C1(n4612), .C2(n2350), .A(n2348), .B(n2346), .ZN(n4543)
         );
  OAI22_X2 U2469 ( .A1(n4543), .A2(n3021), .B1(n4032), .B2(n4558), .ZN(n4526)
         );
  AOI21_X2 U2470 ( .B1(n4036), .B2(n2832), .A(n2401), .ZN(n4078) );
  AOI21_X2 U2471 ( .B1(n2291), .B2(n2140), .A(n2290), .ZN(n4036) );
  AOI21_X1 U2472 ( .B1(n3627), .B2(n3628), .A(n2492), .ZN(n3558) );
  OAI21_X2 U2473 ( .B1(n3787), .B2(n2705), .A(n2704), .ZN(n3903) );
  NAND2_X2 U2474 ( .A1(n2670), .A2(n3753), .ZN(n3787) );
  NAND2_X1 U2475 ( .A1(n2962), .A2(n3500), .ZN(n2535) );
  OAI22_X2 U2476 ( .A1(n4453), .A2(n3028), .B1(n4441), .B2(n4463), .ZN(n4435)
         );
  AND2_X4 U2477 ( .A1(n3118), .A2(n2456), .ZN(n2494) );
  XNOR2_X2 U2478 ( .A(n2454), .B(IR_REG_30__SCAN_IN), .ZN(n3118) );
  INV_X4 U2479 ( .A(n2645), .ZN(n2504) );
  AND2_X4 U2480 ( .A1(n2962), .A2(n3500), .ZN(n2549) );
  XNOR2_X2 U2481 ( .A(n2464), .B(IR_REG_22__SCAN_IN), .ZN(n2468) );
  NAND2_X1 U2482 ( .A1(n4340), .A2(n4339), .ZN(n4852) );
  NAND2_X1 U2483 ( .A1(n4346), .A2(n4347), .ZN(n4363) );
  NAND2_X1 U2484 ( .A1(n3402), .A2(n3401), .ZN(n3403) );
  INV_X1 U2485 ( .A(n3542), .ZN(n2277) );
  AOI21_X1 U2486 ( .B1(n4848), .B2(n4327), .A(n2407), .ZN(n4349) );
  NAND2_X1 U2487 ( .A1(n2362), .A2(n4677), .ZN(n2361) );
  NAND2_X1 U2488 ( .A1(n2381), .A2(n2379), .ZN(n4437) );
  NOR2_X1 U2489 ( .A1(n2380), .A2(n4160), .ZN(n2379) );
  INV_X1 U2490 ( .A(n2382), .ZN(n2380) );
  AND2_X1 U2491 ( .A1(n4285), .A2(n4440), .ZN(n4157) );
  INV_X1 U2492 ( .A(n2855), .ZN(n2854) );
  INV_X1 U2493 ( .A(n2793), .ZN(n2792) );
  AND2_X1 U2494 ( .A1(n4601), .A2(n2162), .ZN(n2351) );
  AOI21_X1 U2495 ( .B1(n3038), .B2(n4219), .A(n2390), .ZN(n2389) );
  INV_X1 U2496 ( .A(n4232), .ZN(n2390) );
  OR2_X1 U2497 ( .A1(n3504), .A2(n3617), .ZN(n4214) );
  AND2_X1 U2498 ( .A1(n2345), .A2(n2341), .ZN(n2340) );
  NAND2_X1 U2499 ( .A1(n4435), .A2(n3029), .ZN(n2342) );
  NAND2_X1 U2500 ( .A1(n3030), .A2(n3029), .ZN(n2341) );
  INV_X1 U2501 ( .A(IR_REG_5__SCAN_IN), .ZN(n2416) );
  AND2_X1 U2502 ( .A1(n4000), .A2(n2306), .ZN(n2305) );
  NAND2_X1 U2503 ( .A1(n2748), .A2(n2307), .ZN(n2306) );
  INV_X1 U2504 ( .A(n4113), .ZN(n2307) );
  OR2_X1 U2505 ( .A1(n2298), .A2(n2402), .ZN(n2296) );
  AND2_X1 U2506 ( .A1(n4028), .A2(n2299), .ZN(n2298) );
  NAND2_X1 U2507 ( .A1(n4089), .A2(n4090), .ZN(n2299) );
  INV_X1 U2508 ( .A(n3436), .ZN(n2206) );
  NOR2_X1 U2509 ( .A1(n3435), .A2(n3412), .ZN(n3419) );
  AND2_X1 U2510 ( .A1(n4816), .A2(REG1_REG_5__SCAN_IN), .ZN(n3412) );
  XNOR2_X1 U2511 ( .A(n4349), .B(n4809), .ZN(n4328) );
  NAND2_X1 U2512 ( .A1(n4345), .A2(n4869), .ZN(n4346) );
  INV_X1 U2513 ( .A(n4343), .ZN(n2210) );
  NAND2_X1 U2514 ( .A1(n2905), .A2(REG3_REG_28__SCAN_IN), .ZN(n4405) );
  OR2_X1 U2515 ( .A1(n2896), .A2(n2895), .ZN(n2907) );
  NAND2_X1 U2516 ( .A1(n2854), .A2(n2213), .ZN(n2883) );
  AOI21_X1 U2517 ( .B1(n4526), .B2(n2334), .A(n2331), .ZN(n2330) );
  INV_X1 U2518 ( .A(n2332), .ZN(n2331) );
  AOI21_X1 U2519 ( .B1(n2334), .B2(n2333), .A(n2187), .ZN(n2332) );
  AOI21_X1 U2520 ( .B1(n2999), .B2(n3716), .A(n2411), .ZN(n3724) );
  AND2_X1 U2521 ( .A1(n4291), .A2(n3831), .ZN(n2999) );
  NAND2_X1 U2522 ( .A1(n4393), .A2(n4385), .ZN(n4383) );
  NAND2_X1 U2523 ( .A1(n4334), .A2(REG1_REG_14__SCAN_IN), .ZN(n4340) );
  NAND2_X1 U2524 ( .A1(n3052), .A2(n2396), .ZN(n2395) );
  INV_X1 U2525 ( .A(n2398), .ZN(n2396) );
  INV_X1 U2526 ( .A(n3003), .ZN(n2328) );
  XNOR2_X1 U2527 ( .A(n2554), .B(n2849), .ZN(n2577) );
  AND2_X1 U2528 ( .A1(n2301), .A2(n4090), .ZN(n2297) );
  AND2_X1 U2529 ( .A1(n3097), .A2(n3098), .ZN(n2853) );
  INV_X1 U2530 ( .A(n2361), .ZN(n2360) );
  NOR2_X1 U2531 ( .A1(n4073), .A2(n2222), .ZN(n2221) );
  AND2_X1 U2532 ( .A1(n2399), .A2(n4632), .ZN(n2398) );
  NAND2_X1 U2533 ( .A1(n4656), .A2(n4229), .ZN(n2399) );
  AND2_X1 U2534 ( .A1(n3848), .A2(n3930), .ZN(n3009) );
  INV_X1 U2535 ( .A(n4227), .ZN(n2372) );
  OAI21_X1 U2536 ( .B1(n2144), .B2(n2372), .A(n4238), .ZN(n2371) );
  OR2_X1 U2537 ( .A1(n3811), .A2(n3801), .ZN(n4227) );
  OR2_X1 U2538 ( .A1(n3796), .A2(n3070), .ZN(n4226) );
  AND2_X1 U2539 ( .A1(n2560), .A2(REG3_REG_6__SCAN_IN), .ZN(n2583) );
  INV_X1 U2540 ( .A(n2562), .ZN(n2560) );
  AND2_X1 U2541 ( .A1(n2468), .A2(n2469), .ZN(n3382) );
  NOR2_X1 U2542 ( .A1(n4446), .A2(n4456), .ZN(n2234) );
  AND2_X1 U2543 ( .A1(n3629), .A2(n3537), .ZN(n4208) );
  NOR2_X1 U2544 ( .A1(n2764), .A2(n2450), .ZN(n2429) );
  NAND2_X1 U2545 ( .A1(n2923), .A2(IR_REG_31__SCAN_IN), .ZN(n2946) );
  OR2_X1 U2546 ( .A1(n2655), .A2(IR_REG_10__SCAN_IN), .ZN(n2717) );
  NAND2_X1 U2547 ( .A1(n2582), .A2(n2412), .ZN(n2287) );
  NAND2_X1 U2548 ( .A1(n3563), .A2(n2575), .ZN(n2289) );
  AND2_X1 U2549 ( .A1(n2571), .A2(DATAI_21_), .ZN(n4040) );
  INV_X1 U2550 ( .A(n2297), .ZN(n2293) );
  NAND2_X1 U2551 ( .A1(n2792), .A2(n2221), .ZN(n2819) );
  OR2_X1 U2552 ( .A1(n4059), .A2(n2322), .ZN(n2321) );
  NAND2_X1 U2553 ( .A1(n2218), .A2(REG3_REG_16__SCAN_IN), .ZN(n2754) );
  AOI21_X1 U2554 ( .B1(n3095), .B2(n2868), .A(n2867), .ZN(n4056) );
  OAI22_X1 U2555 ( .A1(n2645), .A2(n3597), .B1(n3609), .B2(n2135), .ZN(n2558)
         );
  INV_X1 U2556 ( .A(n4070), .ZN(n2294) );
  NOR2_X1 U2557 ( .A1(n2317), .A2(n2311), .ZN(n2310) );
  INV_X1 U2558 ( .A(n2853), .ZN(n2311) );
  INV_X1 U2559 ( .A(n4059), .ZN(n2320) );
  INV_X1 U2560 ( .A(n2509), .ZN(n2972) );
  NAND2_X1 U2561 ( .A1(n2494), .A2(REG2_REG_0__SCAN_IN), .ZN(n2475) );
  OR2_X1 U2562 ( .A1(n2509), .A2(n4968), .ZN(n2474) );
  NOR2_X1 U2563 ( .A1(n3433), .A2(n4828), .ZN(n2243) );
  OAI21_X1 U2564 ( .B1(n3449), .B2(n3448), .A(n2408), .ZN(n3540) );
  OR2_X1 U2565 ( .A1(n3446), .A2(n2587), .ZN(n3442) );
  OAI21_X1 U2566 ( .B1(n3543), .B2(n2276), .A(n2275), .ZN(n2201) );
  NAND2_X1 U2567 ( .A1(n3544), .A2(n2179), .ZN(n2275) );
  NAND2_X1 U2568 ( .A1(n2277), .A2(n2179), .ZN(n2276) );
  NAND2_X1 U2569 ( .A1(n3881), .A2(n3880), .ZN(n4330) );
  OR2_X1 U2570 ( .A1(n4811), .A2(n3954), .ZN(n3880) );
  INV_X1 U2571 ( .A(n4932), .ZN(n4846) );
  NAND2_X1 U2572 ( .A1(n2198), .A2(n2197), .ZN(n4333) );
  AOI21_X1 U2573 ( .B1(n4331), .B2(n4745), .A(n4842), .ZN(n2197) );
  OR2_X1 U2574 ( .A1(n3882), .A2(n2199), .ZN(n2198) );
  INV_X1 U2575 ( .A(n4331), .ZN(n2199) );
  NAND2_X1 U2576 ( .A1(n4852), .A2(n4342), .ZN(n2211) );
  NAND2_X1 U2577 ( .A1(n4874), .A2(n4873), .ZN(n4872) );
  INV_X1 U2578 ( .A(IR_REG_19__SCAN_IN), .ZN(n2466) );
  AOI21_X1 U2579 ( .B1(n2256), .B2(n2257), .A(n2255), .ZN(n2254) );
  INV_X1 U2580 ( .A(n4371), .ZN(n2255) );
  INV_X1 U2581 ( .A(n4356), .ZN(n2256) );
  INV_X1 U2582 ( .A(n4891), .ZN(n2259) );
  INV_X1 U2583 ( .A(n4881), .ZN(n2283) );
  NAND2_X1 U2584 ( .A1(n2343), .A2(n2155), .ZN(n4679) );
  OR2_X1 U2585 ( .A1(n4284), .A2(n4145), .ZN(n4200) );
  OR2_X1 U2586 ( .A1(n4268), .A2(n4428), .ZN(n2345) );
  AND2_X1 U2587 ( .A1(n4396), .A2(n4395), .ZN(n4202) );
  INV_X1 U2588 ( .A(n4420), .ZN(n4428) );
  NAND2_X1 U2589 ( .A1(n2840), .A2(n2839), .ZN(n2855) );
  INV_X1 U2590 ( .A(n2842), .ZN(n2840) );
  INV_X1 U2591 ( .A(n4457), .ZN(n4497) );
  NAND2_X1 U2592 ( .A1(n2792), .A2(n2219), .ZN(n2842) );
  NOR2_X1 U2593 ( .A1(n2220), .A2(n3255), .ZN(n2219) );
  INV_X1 U2594 ( .A(n2221), .ZN(n2220) );
  NAND2_X1 U2595 ( .A1(n4553), .A2(n4040), .ZN(n3022) );
  NAND2_X1 U2596 ( .A1(n2349), .A2(n2347), .ZN(n2346) );
  AOI21_X1 U2597 ( .B1(n2349), .B2(n2143), .A(n2141), .ZN(n2348) );
  INV_X1 U2598 ( .A(n3020), .ZN(n2347) );
  NAND2_X1 U2599 ( .A1(n2775), .A2(REG3_REG_18__SCAN_IN), .ZN(n2793) );
  INV_X1 U2600 ( .A(n2777), .ZN(n2775) );
  NAND2_X1 U2601 ( .A1(n2217), .A2(REG3_REG_17__SCAN_IN), .ZN(n2777) );
  INV_X1 U2602 ( .A(n2754), .ZN(n2217) );
  AND2_X1 U2603 ( .A1(n2352), .A2(n2351), .ZN(n4603) );
  NAND2_X1 U2604 ( .A1(n4544), .A2(n4545), .ZN(n4606) );
  NAND2_X1 U2605 ( .A1(n4644), .A2(n3017), .ZN(n2339) );
  NAND2_X1 U2606 ( .A1(n2164), .A2(n2385), .ZN(n2384) );
  NAND2_X1 U2607 ( .A1(n2343), .A2(n2186), .ZN(n4676) );
  NAND2_X1 U2608 ( .A1(n4680), .A2(n4943), .ZN(n2227) );
  INV_X1 U2609 ( .A(n4040), .ZN(n4536) );
  NOR2_X1 U2610 ( .A1(n4011), .A2(n4589), .ZN(n2238) );
  NAND2_X1 U2611 ( .A1(n4635), .A2(n2146), .ZN(n4556) );
  AND2_X1 U2612 ( .A1(n3069), .A2(n2230), .ZN(n2229) );
  NOR2_X1 U2613 ( .A1(n2998), .A2(n3706), .ZN(n2230) );
  AND3_X1 U2614 ( .A1(n3067), .A2(n3066), .A3(n3065), .ZN(n3080) );
  NAND2_X1 U2615 ( .A1(n3646), .A2(n3636), .ZN(n3664) );
  OR2_X1 U2616 ( .A1(n2468), .A2(n4902), .ZN(n4937) );
  INV_X1 U2617 ( .A(IR_REG_29__SCAN_IN), .ZN(n2452) );
  NOR2_X1 U2618 ( .A1(n2764), .A2(n2161), .ZN(n2453) );
  NAND2_X1 U2619 ( .A1(n2717), .A2(IR_REG_31__SCAN_IN), .ZN(n2691) );
  NOR2_X1 U2620 ( .A1(n2550), .A2(IR_REG_5__SCAN_IN), .ZN(n2625) );
  NAND2_X1 U2621 ( .A1(n2517), .A2(IR_REG_31__SCAN_IN), .ZN(n2531) );
  INV_X1 U2622 ( .A(n2196), .ZN(n2516) );
  AND2_X1 U2623 ( .A1(n2883), .A2(n2870), .ZN(n4465) );
  AOI21_X1 U2624 ( .B1(n2305), .B2(n2183), .A(n2150), .ZN(n2302) );
  INV_X1 U2625 ( .A(n4479), .ZN(n4441) );
  INV_X1 U2626 ( .A(n4553), .ZN(n4083) );
  OAI21_X1 U2627 ( .B1(n4413), .B2(n2132), .A(n2912), .ZN(n4430) );
  NAND2_X1 U2628 ( .A1(n2903), .A2(n2902), .ZN(n4443) );
  OR2_X1 U2629 ( .A1(n2509), .A2(n4977), .ZN(n2590) );
  NAND2_X1 U2630 ( .A1(n2525), .A2(REG0_REG_2__SCAN_IN), .ZN(n2495) );
  OR2_X1 U2631 ( .A1(n2509), .A2(n3387), .ZN(n2496) );
  NAND2_X1 U2632 ( .A1(n2494), .A2(REG2_REG_1__SCAN_IN), .ZN(n2459) );
  NAND2_X1 U2633 ( .A1(n2525), .A2(REG0_REG_1__SCAN_IN), .ZN(n2458) );
  AND2_X1 U2634 ( .A1(n3392), .A2(n3390), .ZN(n4823) );
  NAND2_X1 U2635 ( .A1(n2203), .A2(n2202), .ZN(n3435) );
  NAND2_X1 U2636 ( .A1(n3411), .A2(n2206), .ZN(n2202) );
  XNOR2_X1 U2637 ( .A(n3546), .B(n3444), .ZN(n3547) );
  NAND2_X1 U2638 ( .A1(n3882), .A2(REG1_REG_12__SCAN_IN), .ZN(n4332) );
  XNOR2_X1 U2639 ( .A(n2262), .B(n2261), .ZN(n4334) );
  INV_X1 U2640 ( .A(n4809), .ZN(n2261) );
  OAI21_X1 U2641 ( .B1(n4351), .B2(n4858), .A(n2253), .ZN(n4857) );
  OAI211_X1 U2642 ( .C1(n4852), .C2(n2269), .A(n4870), .B(n2267), .ZN(n4869)
         );
  NAND2_X1 U2643 ( .A1(n2271), .A2(n2274), .ZN(n2269) );
  NAND2_X1 U2644 ( .A1(n4852), .A2(n2185), .ZN(n2267) );
  INV_X1 U2645 ( .A(n4863), .ZN(n4896) );
  NAND2_X1 U2646 ( .A1(n4370), .A2(n4369), .ZN(n4890) );
  AND2_X1 U2647 ( .A1(n4370), .A2(n2257), .ZN(n4889) );
  NAND2_X1 U2648 ( .A1(n4363), .A2(n4362), .ZN(n4882) );
  NAND2_X1 U2649 ( .A1(n2358), .A2(n4898), .ZN(n2357) );
  XNOR2_X1 U2650 ( .A(n4383), .B(n3086), .ZN(n4671) );
  NAND2_X1 U2651 ( .A1(n4967), .A2(n4943), .ZN(n4802) );
  INV_X1 U2652 ( .A(n4965), .ZN(n4967) );
  XNOR2_X1 U2653 ( .A(IR_REG_27__SCAN_IN), .B(IR_REG_28__SCAN_IN), .ZN(n2437)
         );
  NAND2_X1 U2654 ( .A1(n2792), .A2(REG3_REG_19__SCAN_IN), .ZN(n2806) );
  NOR2_X1 U2655 ( .A1(n3444), .A2(n3736), .ZN(n2249) );
  OR2_X1 U2656 ( .A1(n4814), .A2(REG2_REG_8__SCAN_IN), .ZN(n2248) );
  INV_X1 U2657 ( .A(n3548), .ZN(n2251) );
  AND2_X1 U2658 ( .A1(n4862), .A2(REG1_REG_15__SCAN_IN), .ZN(n4343) );
  NOR2_X1 U2659 ( .A1(n4050), .A2(n4062), .ZN(n2213) );
  AOI21_X1 U2660 ( .B1(n4136), .B2(n4472), .A(n2383), .ZN(n2382) );
  NAND2_X1 U2661 ( .A1(n4163), .A2(n3054), .ZN(n4472) );
  INV_X1 U2662 ( .A(n3022), .ZN(n2333) );
  AND2_X1 U2663 ( .A1(n3052), .A2(n4229), .ZN(n2397) );
  NAND2_X1 U2664 ( .A1(n2395), .A2(n2394), .ZN(n2393) );
  INV_X1 U2665 ( .A(n2404), .ZN(n2394) );
  NOR2_X1 U2666 ( .A1(n2726), .A2(n2725), .ZN(n2218) );
  NAND2_X1 U2667 ( .A1(n4245), .A2(n2377), .ZN(n2376) );
  INV_X1 U2668 ( .A(n4245), .ZN(n2378) );
  NOR2_X1 U2669 ( .A1(n3244), .A2(n2658), .ZN(n2216) );
  INV_X1 U2670 ( .A(n2659), .ZN(n2657) );
  INV_X1 U2671 ( .A(n2327), .ZN(n2325) );
  INV_X1 U2672 ( .A(n4217), .ZN(n2387) );
  INV_X1 U2673 ( .A(n2389), .ZN(n2385) );
  CLKBUF_X1 U2674 ( .A(n3035), .Z(n4209) );
  NAND2_X1 U2675 ( .A1(n2989), .A2(n2472), .ZN(n3035) );
  NAND2_X1 U2676 ( .A1(n2990), .A2(n3646), .ZN(n4206) );
  NAND2_X1 U2677 ( .A1(n2345), .A2(n3031), .ZN(n2344) );
  NAND2_X1 U2678 ( .A1(n4428), .A2(n2234), .ZN(n2233) );
  AND2_X1 U2679 ( .A1(n3801), .A2(n2237), .ZN(n2236) );
  INV_X1 U2680 ( .A(n3639), .ZN(n3640) );
  XNOR2_X1 U2681 ( .A(IR_REG_1__SCAN_IN), .B(keyinput62), .ZN(n3295) );
  OR2_X1 U2682 ( .A1(n2640), .A2(IR_REG_9__SCAN_IN), .ZN(n2655) );
  NAND2_X1 U2683 ( .A1(n2583), .A2(n2170), .ZN(n2634) );
  INV_X1 U2684 ( .A(n4430), .ZN(n3032) );
  NAND2_X1 U2685 ( .A1(n2583), .A2(n2148), .ZN(n2618) );
  XNOR2_X1 U2686 ( .A(n2521), .B(n2849), .ZN(n2522) );
  NAND2_X1 U2687 ( .A1(n4093), .A2(n2297), .ZN(n2295) );
  OR2_X1 U2688 ( .A1(n2634), .A2(n3659), .ZN(n2659) );
  OAI22_X1 U2689 ( .A1(n2645), .A2(n2989), .B1(n3646), .B2(n2535), .ZN(n2489)
         );
  XNOR2_X1 U2690 ( .A(n2467), .B(n2849), .ZN(n2491) );
  NAND3_X1 U2691 ( .A1(REG3_REG_3__SCAN_IN), .A2(REG3_REG_4__SCAN_IN), .A3(
        REG3_REG_5__SCAN_IN), .ZN(n2562) );
  INV_X1 U2692 ( .A(n2982), .ZN(n2980) );
  NAND2_X1 U2693 ( .A1(n2304), .A2(n2748), .ZN(n4111) );
  NAND2_X1 U2694 ( .A1(n2724), .A2(n2723), .ZN(n2304) );
  NAND2_X1 U2695 ( .A1(n4317), .A2(n3380), .ZN(n3400) );
  NAND2_X1 U2696 ( .A1(n3389), .A2(n3388), .ZN(n3406) );
  INV_X1 U2697 ( .A(n4817), .ZN(n3394) );
  NAND2_X1 U2698 ( .A1(n3404), .A2(n2241), .ZN(n2240) );
  INV_X1 U2699 ( .A(n3433), .ZN(n2241) );
  AND2_X1 U2700 ( .A1(n3541), .A2(n4814), .ZN(n3542) );
  AND2_X1 U2701 ( .A1(n3451), .A2(REG1_REG_8__SCAN_IN), .ZN(n3543) );
  NAND2_X1 U2702 ( .A1(n4846), .A2(REG1_REG_13__SCAN_IN), .ZN(n2263) );
  NAND2_X1 U2703 ( .A1(n4328), .A2(REG2_REG_14__SCAN_IN), .ZN(n4352) );
  INV_X1 U2704 ( .A(n2270), .ZN(n2268) );
  NOR2_X1 U2705 ( .A1(n4344), .A2(n4854), .ZN(n2270) );
  INV_X1 U2706 ( .A(n2272), .ZN(n2271) );
  OAI21_X1 U2707 ( .B1(n2274), .B2(n4342), .A(n2273), .ZN(n2272) );
  NAND2_X1 U2708 ( .A1(n4928), .A2(n4343), .ZN(n2273) );
  OR2_X1 U2709 ( .A1(n4928), .A2(n4343), .ZN(n2274) );
  AND2_X1 U2710 ( .A1(n4403), .A2(n4402), .ZN(n4404) );
  NOR2_X1 U2711 ( .A1(n4397), .A2(n2365), .ZN(n2364) );
  INV_X1 U2712 ( .A(n4426), .ZN(n2365) );
  OAI21_X1 U2713 ( .B1(n2364), .B2(n2361), .A(n2223), .ZN(n2358) );
  NAND2_X1 U2714 ( .A1(n2363), .A2(n4674), .ZN(n2223) );
  INV_X1 U2715 ( .A(n4202), .ZN(n4389) );
  AND2_X1 U2716 ( .A1(n2907), .A2(n2897), .ZN(n4421) );
  AND2_X1 U2717 ( .A1(n2848), .A2(n2847), .ZN(n4517) );
  OR2_X1 U2718 ( .A1(n4606), .A2(n4565), .ZN(n4567) );
  NOR2_X1 U2719 ( .A1(n4632), .A2(n2338), .ZN(n2337) );
  INV_X1 U2720 ( .A(n3018), .ZN(n2338) );
  NAND2_X1 U2721 ( .A1(n4657), .A2(n4229), .ZN(n2392) );
  NAND2_X1 U2722 ( .A1(n4653), .A2(n4229), .ZN(n4620) );
  AND3_X1 U2723 ( .A1(n2713), .A2(n2712), .A3(n2711), .ZN(n4651) );
  OR2_X1 U2724 ( .A1(n4657), .A2(n4656), .ZN(n4653) );
  INV_X1 U2725 ( .A(REG3_REG_15__SCAN_IN), .ZN(n2725) );
  INV_X1 U2726 ( .A(n2218), .ZN(n2738) );
  NAND2_X1 U2727 ( .A1(n2706), .A2(REG3_REG_14__SCAN_IN), .ZN(n2726) );
  INV_X1 U2728 ( .A(n2707), .ZN(n2706) );
  NAND2_X1 U2729 ( .A1(n2657), .A2(n2215), .ZN(n2707) );
  AND2_X1 U2730 ( .A1(n2216), .A2(REG3_REG_13__SCAN_IN), .ZN(n2215) );
  NAND2_X1 U2731 ( .A1(n3011), .A2(n3010), .ZN(n3965) );
  INV_X1 U2732 ( .A(n3009), .ZN(n3010) );
  NAND2_X1 U2733 ( .A1(n2657), .A2(REG3_REG_11__SCAN_IN), .ZN(n2683) );
  NAND2_X1 U2734 ( .A1(n2657), .A2(n2216), .ZN(n2685) );
  NAND2_X1 U2735 ( .A1(n3042), .A2(n4243), .ZN(n3962) );
  AOI21_X1 U2736 ( .B1(n2370), .B2(n2372), .A(n2368), .ZN(n2367) );
  INV_X1 U2737 ( .A(n2371), .ZN(n2370) );
  NAND2_X1 U2738 ( .A1(n3041), .A2(n2144), .ZN(n2369) );
  CLKBUF_X1 U2739 ( .A(n3808), .Z(n3809) );
  NAND2_X1 U2740 ( .A1(n2583), .A2(REG3_REG_7__SCAN_IN), .ZN(n2603) );
  NAND2_X1 U2741 ( .A1(n2391), .A2(n2389), .ZN(n2388) );
  NAND2_X1 U2742 ( .A1(n3502), .A2(n4219), .ZN(n2391) );
  INV_X1 U2743 ( .A(n4622), .ZN(n4650) );
  AND2_X1 U2744 ( .A1(n3382), .A2(n4819), .ZN(n4623) );
  AND2_X1 U2745 ( .A1(n3382), .A2(n4307), .ZN(n4622) );
  NOR2_X1 U2746 ( .A1(n4462), .A2(n2233), .ZN(n3074) );
  INV_X1 U2747 ( .A(n2234), .ZN(n2232) );
  CLKBUF_X1 U2748 ( .A(n4462), .Z(n4483) );
  INV_X1 U2749 ( .A(n4065), .ZN(n4484) );
  INV_X1 U2750 ( .A(n3043), .ZN(n3973) );
  NAND2_X1 U2751 ( .A1(n3802), .A2(n2147), .ZN(n3928) );
  INV_X1 U2752 ( .A(n3005), .ZN(n3801) );
  NAND2_X1 U2753 ( .A1(n3802), .A2(n3801), .ZN(n3816) );
  AND2_X1 U2754 ( .A1(n3069), .A2(n3602), .ZN(n2228) );
  NAND2_X1 U2755 ( .A1(n4924), .A2(n2962), .ZN(n3531) );
  NAND2_X1 U2756 ( .A1(n2465), .A2(n2434), .ZN(n2435) );
  INV_X1 U2757 ( .A(IR_REG_17__SCAN_IN), .ZN(n2423) );
  NAND2_X1 U2758 ( .A1(n2444), .A2(n2445), .ZN(n2264) );
  INV_X1 U2759 ( .A(IR_REG_31__SCAN_IN), .ZN(n2444) );
  NAND3_X1 U2760 ( .A1(IR_REG_0__SCAN_IN), .A2(IR_REG_31__SCAN_IN), .A3(
        IR_REG_1__SCAN_IN), .ZN(n2265) );
  NAND2_X1 U2761 ( .A1(n2288), .A2(n2289), .ZN(n3572) );
  AND2_X1 U2762 ( .A1(n3826), .A2(n2287), .ZN(n2288) );
  XNOR2_X1 U2763 ( .A(n2919), .B(n2920), .ZN(n4020) );
  XNOR2_X1 U2764 ( .A(n2491), .B(n2489), .ZN(n3627) );
  AND2_X1 U2765 ( .A1(n2837), .A2(n2836), .ZN(n4043) );
  INV_X1 U2766 ( .A(n2292), .ZN(n2290) );
  AOI21_X1 U2767 ( .B1(n2140), .B2(n2293), .A(n4069), .ZN(n2292) );
  AND2_X1 U2768 ( .A1(n2842), .A2(n2820), .ZN(n4538) );
  AND2_X1 U2769 ( .A1(n2889), .A2(n2888), .ZN(n4459) );
  OR2_X1 U2770 ( .A1(n4448), .A2(n2133), .ZN(n2889) );
  INV_X1 U2771 ( .A(n2314), .ZN(n4047) );
  OAI21_X1 U2772 ( .B1(n3095), .B2(n2315), .A(n2318), .ZN(n2314) );
  INV_X1 U2773 ( .A(n2321), .ZN(n2315) );
  XOR2_X1 U2774 ( .A(n2750), .B(n2749), .Z(n4000) );
  AND3_X1 U2775 ( .A1(n2742), .A2(n2741), .A3(n2740), .ZN(n4652) );
  NAND2_X1 U2776 ( .A1(n3095), .A2(n2145), .ZN(n4057) );
  OR2_X1 U2777 ( .A1(n2518), .A2(n2479), .ZN(n2480) );
  INV_X1 U2778 ( .A(n4118), .ZN(n4082) );
  INV_X1 U2779 ( .A(n4117), .ZN(n4095) );
  INV_X1 U2780 ( .A(n4119), .ZN(n4096) );
  AOI21_X1 U2781 ( .B1(n2316), .B2(n2319), .A(n2313), .ZN(n2312) );
  INV_X1 U2782 ( .A(n4048), .ZN(n2313) );
  AOI21_X1 U2783 ( .B1(n4621), .B2(n2504), .A(n2736), .ZN(n4113) );
  NAND2_X1 U2784 ( .A1(n2978), .A2(n2977), .ZN(n4284) );
  OR2_X1 U2785 ( .A1(n4405), .A2(n2132), .ZN(n2978) );
  NAND2_X1 U2786 ( .A1(n2875), .A2(n2874), .ZN(n4479) );
  NAND2_X1 U2787 ( .A1(n2861), .A2(n2860), .ZN(n4457) );
  OR2_X1 U2788 ( .A1(n4487), .A2(n2133), .ZN(n2861) );
  INV_X1 U2789 ( .A(n4043), .ZN(n4532) );
  OR2_X1 U2790 ( .A1(n4072), .A2(n2132), .ZN(n2812) );
  NAND2_X1 U2791 ( .A1(n2783), .A2(n2782), .ZN(n4608) );
  OR2_X1 U2792 ( .A1(n4597), .A2(n2132), .ZN(n2783) );
  NAND2_X1 U2793 ( .A1(n2760), .A2(n2759), .ZN(n4624) );
  INV_X1 U2794 ( .A(n4652), .ZN(n4116) );
  OR2_X1 U2795 ( .A1(n3462), .A2(n3420), .ZN(n2569) );
  AND2_X1 U2796 ( .A1(n4924), .A2(n3094), .ZN(n3521) );
  NAND2_X1 U2797 ( .A1(n2898), .A2(REG3_REG_0__SCAN_IN), .ZN(n2478) );
  XNOR2_X1 U2798 ( .A(n3406), .B(n3394), .ZN(n3405) );
  NAND2_X1 U2799 ( .A1(n2240), .A2(n2239), .ZN(n3432) );
  AND2_X1 U2800 ( .A1(n2242), .A2(n2245), .ZN(n3434) );
  NAND2_X1 U2801 ( .A1(n4827), .A2(REG2_REG_4__SCAN_IN), .ZN(n2242) );
  NAND2_X1 U2802 ( .A1(n2204), .A2(n2208), .ZN(n2207) );
  NAND2_X1 U2803 ( .A1(n4831), .A2(REG1_REG_4__SCAN_IN), .ZN(n2204) );
  XNOR2_X1 U2804 ( .A(n3419), .B(n3413), .ZN(n2209) );
  AOI22_X1 U2805 ( .A1(n3419), .A2(n2167), .B1(n3413), .B2(n3420), .ZN(n3449)
         );
  AND2_X1 U2806 ( .A1(n2195), .A2(n2250), .ZN(n3549) );
  NAND2_X1 U2807 ( .A1(n3547), .A2(REG2_REG_8__SCAN_IN), .ZN(n2250) );
  NOR2_X1 U2808 ( .A1(n3543), .A2(n3542), .ZN(n3545) );
  XNOR2_X1 U2809 ( .A(n2201), .B(n3773), .ZN(n3658) );
  CLKBUF_X1 U2810 ( .A(n3771), .Z(n3772) );
  NAND2_X1 U2811 ( .A1(n3776), .A2(n2200), .ZN(n3779) );
  OR2_X1 U2812 ( .A1(n2201), .A2(n3777), .ZN(n2200) );
  INV_X1 U2813 ( .A(n4333), .ZN(n4841) );
  AND2_X1 U2814 ( .A1(n4352), .A2(n4351), .ZN(n4859) );
  INV_X1 U2815 ( .A(n2211), .ZN(n4853) );
  AND2_X1 U2816 ( .A1(n4823), .A2(n4305), .ZN(n4877) );
  AND2_X1 U2817 ( .A1(n4823), .A2(n4819), .ZN(n4863) );
  OAI21_X1 U2818 ( .B1(n4355), .B2(n2258), .A(n2254), .ZN(n2260) );
  NAND2_X1 U2819 ( .A1(n2279), .A2(n2278), .ZN(n4366) );
  NAND2_X1 U2820 ( .A1(n2282), .A2(n2156), .ZN(n2278) );
  AND2_X1 U2821 ( .A1(n4347), .A2(n2156), .ZN(n2280) );
  NAND2_X1 U2822 ( .A1(n4405), .A2(n2908), .ZN(n4413) );
  XNOR2_X1 U2823 ( .A(n4390), .B(n4202), .ZN(n4410) );
  NAND2_X1 U2824 ( .A1(n2336), .A2(n3022), .ZN(n2335) );
  NOR2_X1 U2825 ( .A1(n4603), .A2(n2143), .ZN(n4578) );
  NAND2_X1 U2826 ( .A1(n3711), .A2(n3001), .ZN(n2329) );
  AND2_X1 U2827 ( .A1(n3499), .A2(n3501), .ZN(n4904) );
  NAND2_X1 U2828 ( .A1(n2212), .A2(n2149), .ZN(n4752) );
  INV_X1 U2829 ( .A(n4675), .ZN(n2212) );
  AND2_X1 U2830 ( .A1(n4635), .A2(n2238), .ZN(n4580) );
  XNOR2_X1 U2831 ( .A(n2925), .B(n2924), .ZN(n3373) );
  INV_X1 U2832 ( .A(n2456), .ZN(n4804) );
  NAND2_X1 U2833 ( .A1(n2463), .A2(IR_REG_31__SCAN_IN), .ZN(n2432) );
  XNOR2_X1 U2834 ( .A(n2718), .B(IR_REG_14__SCAN_IN), .ZN(n4809) );
  XNOR2_X1 U2835 ( .A(n2678), .B(IR_REG_13__SCAN_IN), .ZN(n4932) );
  XNOR2_X1 U2836 ( .A(n2691), .B(n2690), .ZN(n4811) );
  XNOR2_X1 U2837 ( .A(n2626), .B(IR_REG_9__SCAN_IN), .ZN(n4813) );
  XNOR2_X1 U2838 ( .A(n2551), .B(IR_REG_5__SCAN_IN), .ZN(n4816) );
  XNOR2_X1 U2839 ( .A(n2534), .B(n2533), .ZN(n3409) );
  XNOR2_X1 U2840 ( .A(n2531), .B(IR_REG_3__SCAN_IN), .ZN(n4817) );
  AOI21_X1 U2841 ( .B1(n4888), .B2(n2169), .A(n4887), .ZN(n4895) );
  NAND2_X1 U2842 ( .A1(n2226), .A2(n2224), .ZN(U3547) );
  OR2_X1 U2843 ( .A1(n4975), .A2(n2225), .ZN(n2224) );
  NAND2_X1 U2844 ( .A1(n4752), .A2(n4975), .ZN(n2226) );
  INV_X1 U2845 ( .A(REG1_REG_29__SCAN_IN), .ZN(n2225) );
  AND2_X1 U2846 ( .A1(n3092), .A2(n3091), .ZN(n3093) );
  NOR2_X1 U2847 ( .A1(n3964), .A2(n3012), .ZN(n2139) );
  AND2_X1 U2848 ( .A1(n2296), .A2(n2294), .ZN(n2140) );
  AND2_X1 U2849 ( .A1(n4591), .A2(n4579), .ZN(n2141) );
  NAND2_X1 U2850 ( .A1(n3811), .A2(n3005), .ZN(n2142) );
  AND2_X1 U2851 ( .A1(n4572), .A2(n4595), .ZN(n2143) );
  AND2_X1 U2852 ( .A1(n2373), .A2(n4224), .ZN(n2144) );
  NAND2_X1 U2853 ( .A1(n4612), .A2(n3020), .ZN(n2352) );
  AND2_X1 U2854 ( .A1(n2868), .A2(n2867), .ZN(n2145) );
  AND2_X1 U2855 ( .A1(n2238), .A2(n4579), .ZN(n2146) );
  AND2_X1 U2856 ( .A1(n2236), .A2(n3757), .ZN(n2147) );
  INV_X1 U2857 ( .A(n3817), .ZN(n2237) );
  AND2_X1 U2858 ( .A1(REG3_REG_7__SCAN_IN), .A2(REG3_REG_8__SCAN_IN), .ZN(
        n2148) );
  AND4_X2 U2859 ( .A1(n4676), .A2(n4681), .A3(n2227), .A4(n2180), .ZN(n2149)
         );
  NAND2_X1 U2860 ( .A1(n2339), .A2(n3018), .ZN(n4629) );
  NAND2_X1 U2861 ( .A1(n2335), .A2(n2334), .ZN(n4510) );
  NAND2_X1 U2862 ( .A1(n2295), .A2(n2296), .ZN(n4068) );
  AND2_X1 U2863 ( .A1(n4126), .A2(n4230), .ZN(n4176) );
  INV_X1 U2864 ( .A(n4176), .ZN(n3015) );
  AND2_X1 U2865 ( .A1(n2752), .A2(n2751), .ZN(n2150) );
  INV_X1 U2866 ( .A(n4591), .ZN(n3482) );
  AND2_X1 U2867 ( .A1(n2799), .A2(n2798), .ZN(n4591) );
  AND3_X1 U2868 ( .A1(n2287), .A2(n2597), .A3(n3826), .ZN(n2151) );
  OR2_X1 U2869 ( .A1(n3013), .A2(n2158), .ZN(n2152) );
  NOR2_X1 U2870 ( .A1(n3444), .A2(n4814), .ZN(n2153) );
  AND2_X1 U2871 ( .A1(n2329), .A2(n2193), .ZN(n2154) );
  AND2_X1 U2872 ( .A1(n4389), .A2(n2344), .ZN(n2155) );
  NAND2_X1 U2873 ( .A1(n3802), .A2(n2236), .ZN(n2235) );
  OR2_X1 U2874 ( .A1(n4926), .A2(n4364), .ZN(n2156) );
  NAND2_X1 U2875 ( .A1(n2392), .A2(n2398), .ZN(n4544) );
  OR2_X1 U2876 ( .A1(n2463), .A2(IR_REG_21__SCAN_IN), .ZN(n2157) );
  NOR2_X1 U2877 ( .A1(n4501), .A2(n3073), .ZN(n4482) );
  AND3_X1 U2878 ( .A1(n2724), .A2(n2308), .A3(n2723), .ZN(n3998) );
  AND2_X1 U2879 ( .A1(n3983), .A2(n3043), .ZN(n2158) );
  OR2_X1 U2880 ( .A1(n4462), .A2(n2232), .ZN(n2159) );
  AND2_X1 U2881 ( .A1(n4248), .A2(n2376), .ZN(n2160) );
  INV_X1 U2882 ( .A(n2998), .ZN(n3602) );
  OR2_X1 U2883 ( .A1(n2450), .A2(n2449), .ZN(n2161) );
  NAND2_X1 U2884 ( .A1(n4624), .A2(n4011), .ZN(n2162) );
  NAND2_X1 U2885 ( .A1(n4083), .A2(n4536), .ZN(n2163) );
  NOR2_X1 U2886 ( .A1(n4394), .A2(n4399), .ZN(n4393) );
  NAND2_X1 U2887 ( .A1(n2309), .A2(n2312), .ZN(n4100) );
  OAI21_X1 U2888 ( .B1(n4093), .B2(n4089), .A(n4090), .ZN(n4027) );
  NAND2_X1 U2889 ( .A1(n2381), .A2(n2382), .ZN(n4454) );
  NOR2_X1 U2890 ( .A1(n4233), .A2(n2387), .ZN(n2164) );
  INV_X1 U2891 ( .A(n3921), .ZN(n3930) );
  OR2_X1 U2892 ( .A1(n4591), .A2(n4579), .ZN(n2165) );
  OR2_X1 U2893 ( .A1(n4462), .A2(n4456), .ZN(n2166) );
  NAND2_X2 U2894 ( .A1(n3076), .A2(n2414), .ZN(n2645) );
  OR2_X1 U2895 ( .A1(n3413), .A2(n3420), .ZN(n2167) );
  INV_X1 U2896 ( .A(n2472), .ZN(n3646) );
  OAI21_X1 U2897 ( .B1(n2518), .B2(n3107), .A(n2446), .ZN(n2472) );
  AND2_X1 U2898 ( .A1(n2295), .A2(n2140), .ZN(n2168) );
  NAND2_X1 U2899 ( .A1(n4363), .A2(n2281), .ZN(n2169) );
  AND2_X1 U2900 ( .A1(n4511), .A2(n2163), .ZN(n2334) );
  AND2_X1 U2901 ( .A1(n2148), .A2(REG3_REG_9__SCAN_IN), .ZN(n2170) );
  AND2_X1 U2902 ( .A1(n4253), .A2(n4545), .ZN(n4632) );
  AND2_X1 U2903 ( .A1(n3006), .A2(n3801), .ZN(n2171) );
  NAND2_X1 U2904 ( .A1(n4333), .A2(n2263), .ZN(n2262) );
  NAND2_X1 U2905 ( .A1(n4816), .A2(REG2_REG_5__SCAN_IN), .ZN(n2172) );
  INV_X1 U2906 ( .A(n2350), .ZN(n2349) );
  OAI21_X1 U2907 ( .B1(n2351), .B2(n2143), .A(n2165), .ZN(n2350) );
  INV_X1 U2908 ( .A(n3404), .ZN(n2245) );
  AND2_X1 U2909 ( .A1(n3403), .A2(n4833), .ZN(n3404) );
  AND2_X1 U2910 ( .A1(n2352), .A2(n2162), .ZN(n2173) );
  AND2_X1 U2911 ( .A1(n2147), .A2(n3930), .ZN(n2174) );
  AND2_X1 U2912 ( .A1(n2335), .A2(n2163), .ZN(n2175) );
  AND2_X1 U2913 ( .A1(n2206), .A2(REG1_REG_4__SCAN_IN), .ZN(n2176) );
  AND2_X1 U2914 ( .A1(n2211), .A2(n2210), .ZN(n2177) );
  NAND2_X1 U2915 ( .A1(n2251), .A2(n2248), .ZN(n2178) );
  INV_X1 U2916 ( .A(n2402), .ZN(n2301) );
  INV_X1 U2917 ( .A(n4975), .ZN(n4976) );
  AND2_X2 U2918 ( .A1(n3080), .A2(n3079), .ZN(n4975) );
  NAND2_X1 U2919 ( .A1(n4813), .A2(REG1_REG_9__SCAN_IN), .ZN(n2179) );
  INV_X1 U2920 ( .A(n2867), .ZN(n2322) );
  NAND2_X1 U2921 ( .A1(n2303), .A2(n2302), .ZN(n4007) );
  NAND2_X1 U2922 ( .A1(n2388), .A2(n4217), .ZN(n3742) );
  NAND2_X1 U2923 ( .A1(n2369), .A2(n4227), .ZN(n3810) );
  OR3_X1 U2924 ( .A1(n4678), .A2(n4959), .A3(n4677), .ZN(n2180) );
  AND2_X1 U2925 ( .A1(n4674), .A2(n4744), .ZN(n2181) );
  OR2_X1 U2926 ( .A1(n2882), .A2(n2881), .ZN(n2182) );
  INV_X1 U2927 ( .A(n4161), .ZN(n2383) );
  INV_X1 U2928 ( .A(n2319), .ZN(n2318) );
  OAI22_X1 U2929 ( .A1(n2145), .A2(n2320), .B1(n2868), .B2(n2867), .ZN(n2319)
         );
  NAND2_X1 U2930 ( .A1(n3918), .A2(n3852), .ZN(n4243) );
  INV_X1 U2931 ( .A(n4243), .ZN(n2377) );
  AND2_X1 U2932 ( .A1(n2308), .A2(n4113), .ZN(n2183) );
  INV_X1 U2933 ( .A(n4011), .ZN(n4613) );
  INV_X1 U2934 ( .A(n3071), .ZN(n4558) );
  AND2_X1 U2935 ( .A1(n4332), .A2(n4331), .ZN(n2184) );
  NAND2_X1 U2936 ( .A1(n4200), .A2(n4199), .ZN(n4677) );
  AND2_X1 U2937 ( .A1(n2268), .A2(n2271), .ZN(n2185) );
  NAND2_X1 U2938 ( .A1(n4635), .A2(n4613), .ZN(n4594) );
  OR2_X1 U2939 ( .A1(n4289), .A2(n2237), .ZN(n4236) );
  INV_X1 U2940 ( .A(n4236), .ZN(n2368) );
  INV_X1 U2941 ( .A(n2317), .ZN(n2316) );
  OAI21_X1 U2942 ( .B1(n2319), .B2(n2321), .A(n2182), .ZN(n2317) );
  AND2_X1 U2943 ( .A1(n2155), .A2(n2181), .ZN(n2186) );
  NOR2_X1 U2944 ( .A1(n4043), .A2(n4514), .ZN(n2187) );
  INV_X1 U2945 ( .A(n2363), .ZN(n2362) );
  OAI21_X1 U2946 ( .B1(n4397), .B2(n4140), .A(n4396), .ZN(n2363) );
  NAND2_X1 U2947 ( .A1(n3563), .A2(n3824), .ZN(n2188) );
  NOR2_X1 U2948 ( .A1(n4858), .A2(n3993), .ZN(n2189) );
  NAND2_X1 U2949 ( .A1(n4813), .A2(REG2_REG_9__SCAN_IN), .ZN(n2190) );
  AND2_X1 U2950 ( .A1(n2146), .A2(n4558), .ZN(n2191) );
  INV_X1 U2951 ( .A(n3076), .ZN(n4943) );
  AND2_X1 U2952 ( .A1(n3512), .A2(n2229), .ZN(n3704) );
  NOR2_X1 U2953 ( .A1(n3666), .A2(n3590), .ZN(n3511) );
  NAND2_X1 U2954 ( .A1(n3512), .A2(n3602), .ZN(n3601) );
  NAND2_X1 U2955 ( .A1(n3512), .A2(n2228), .ZN(n3705) );
  AND2_X1 U2956 ( .A1(n3057), .A2(n4276), .ZN(n4655) );
  AND2_X1 U2957 ( .A1(n3511), .A2(n3609), .ZN(n3512) );
  INV_X1 U2958 ( .A(n4069), .ZN(n2300) );
  NOR2_X1 U2959 ( .A1(n3545), .A2(n3544), .ZN(n2192) );
  AND2_X1 U2960 ( .A1(n3004), .A2(n3003), .ZN(n2193) );
  INV_X1 U2961 ( .A(REG3_REG_19__SCAN_IN), .ZN(n2222) );
  INV_X1 U2962 ( .A(n2235), .ZN(n3815) );
  INV_X1 U2963 ( .A(n2258), .ZN(n2257) );
  NAND2_X1 U2964 ( .A1(n4369), .A2(n2259), .ZN(n2258) );
  AND2_X1 U2965 ( .A1(n2213), .A2(REG3_REG_26__SCAN_IN), .ZN(n2194) );
  NAND2_X1 U2966 ( .A1(n3546), .A2(n4814), .ZN(n2195) );
  INV_X1 U2967 ( .A(IR_REG_30__SCAN_IN), .ZN(n4017) );
  INV_X1 U2968 ( .A(REG3_REG_26__SCAN_IN), .ZN(n2214) );
  INV_X1 U2969 ( .A(n2282), .ZN(n2281) );
  NAND2_X1 U2970 ( .A1(n4362), .A2(n2283), .ZN(n2282) );
  INV_X2 U2971 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  NAND3_X1 U2972 ( .A1(n2196), .A2(n2264), .A3(n2265), .ZN(n3383) );
  NAND4_X1 U2973 ( .A1(n2196), .A2(REG1_REG_1__SCAN_IN), .A3(n2265), .A4(n2264), .ZN(n3385) );
  NAND2_X1 U2974 ( .A1(n4831), .A2(n2176), .ZN(n2203) );
  INV_X1 U2975 ( .A(n3411), .ZN(n2208) );
  NOR3_X1 U2976 ( .A1(n4880), .A2(n3435), .A3(n2205), .ZN(n3440) );
  NOR2_X1 U2977 ( .A1(n2207), .A2(n2206), .ZN(n2205) );
  XNOR2_X1 U2978 ( .A(n2209), .B(REG1_REG_6__SCAN_IN), .ZN(n3416) );
  NAND3_X1 U2979 ( .A1(n2357), .A2(n2355), .A3(n2353), .ZN(n4675) );
  NAND2_X1 U2980 ( .A1(n2854), .A2(n2194), .ZN(n2896) );
  NAND2_X1 U2981 ( .A1(n2854), .A2(REG3_REG_24__SCAN_IN), .ZN(n2869) );
  INV_X1 U2982 ( .A(n2231), .ZN(n4394) );
  NOR3_X2 U2983 ( .A1(n4462), .A2(n2233), .A3(n4391), .ZN(n2231) );
  AND2_X2 U2984 ( .A1(n3802), .A2(n2174), .ZN(n3974) );
  NAND2_X1 U2985 ( .A1(n4635), .A2(n2191), .ZN(n4557) );
  INV_X1 U2986 ( .A(n2244), .ZN(n3422) );
  AND2_X2 U2987 ( .A1(n2252), .A2(n2190), .ZN(n3771) );
  NAND2_X1 U2988 ( .A1(n2247), .A2(n2246), .ZN(n2252) );
  AOI21_X1 U2989 ( .B1(n3546), .B2(n2153), .A(n2178), .ZN(n2247) );
  INV_X1 U2990 ( .A(n2252), .ZN(n3657) );
  NAND2_X1 U2991 ( .A1(n4328), .A2(n2189), .ZN(n2253) );
  NAND2_X1 U2992 ( .A1(n4355), .A2(n4356), .ZN(n4370) );
  INV_X1 U2993 ( .A(n2260), .ZN(n4373) );
  INV_X2 U2994 ( .A(IR_REG_1__SCAN_IN), .ZN(n2445) );
  INV_X1 U2995 ( .A(n3383), .ZN(n4299) );
  OAI211_X1 U2996 ( .C1(n4852), .C2(n2274), .A(n2271), .B(n2266), .ZN(n4871)
         );
  NAND2_X1 U2997 ( .A1(n4852), .A2(n2270), .ZN(n2266) );
  NAND2_X1 U2998 ( .A1(n4346), .A2(n2280), .ZN(n2279) );
  NAND2_X1 U2999 ( .A1(n2992), .A2(n3068), .ZN(n3666) );
  AOI21_X1 U3000 ( .B1(n4378), .B2(n4893), .A(n4377), .ZN(n4379) );
  XNOR2_X2 U3001 ( .A(n4323), .B(n4810), .ZN(n4326) );
  OAI211_X1 U3002 ( .C1(n2286), .C2(n2285), .A(n2284), .B(n2987), .ZN(U3217)
         );
  NAND2_X1 U3003 ( .A1(n2286), .A2(n2400), .ZN(n2284) );
  NAND2_X1 U3004 ( .A1(n2955), .A2(n2953), .ZN(n2285) );
  INV_X1 U3005 ( .A(n4093), .ZN(n2291) );
  NAND3_X1 U3006 ( .A1(n2724), .A2(n2723), .A3(n2305), .ZN(n2303) );
  INV_X1 U3007 ( .A(n2748), .ZN(n2308) );
  NAND2_X1 U3008 ( .A1(n3096), .A2(n2853), .ZN(n3095) );
  NAND2_X1 U3009 ( .A1(n3096), .A2(n2310), .ZN(n2309) );
  NOR2_X1 U3010 ( .A1(n2764), .A2(IR_REG_18__SCAN_IN), .ZN(n2433) );
  NOR2_X2 U3011 ( .A1(n2420), .A2(n3128), .ZN(n2421) );
  NOR2_X2 U3012 ( .A1(n2550), .A2(n2418), .ZN(n2422) );
  INV_X1 U3013 ( .A(n3004), .ZN(n2326) );
  NAND2_X1 U3014 ( .A1(n2324), .A2(n2323), .ZN(n3808) );
  NAND3_X1 U3015 ( .A1(n3711), .A2(n2142), .A3(n3001), .ZN(n2323) );
  INV_X1 U3016 ( .A(n4526), .ZN(n2336) );
  INV_X1 U3017 ( .A(n2330), .ZN(n4492) );
  NAND2_X1 U3018 ( .A1(n2339), .A2(n2337), .ZN(n4630) );
  OAI21_X2 U3019 ( .B1(n4435), .B2(n3030), .A(n3029), .ZN(n4419) );
  AND2_X1 U3020 ( .A1(n2422), .A2(n2421), .ZN(n2761) );
  AOI21_X1 U3021 ( .B1(n4425), .B2(n4426), .A(n4139), .ZN(n4398) );
  INV_X1 U3022 ( .A(n2354), .ZN(n2353) );
  OAI21_X1 U3023 ( .B1(n2359), .B2(n4425), .A(n4404), .ZN(n2354) );
  NAND3_X1 U3024 ( .A1(n4425), .A2(n2364), .A3(n2356), .ZN(n2355) );
  AND2_X1 U3025 ( .A1(n4674), .A2(n4898), .ZN(n2356) );
  NAND2_X1 U3026 ( .A1(n2360), .A2(n4898), .ZN(n2359) );
  NAND2_X1 U3027 ( .A1(n3041), .A2(n2370), .ZN(n2366) );
  NAND2_X1 U3028 ( .A1(n2366), .A2(n2367), .ZN(n3840) );
  NAND2_X1 U3029 ( .A1(n3041), .A2(n4224), .ZN(n3793) );
  INV_X1 U3030 ( .A(n4235), .ZN(n2373) );
  OAI21_X1 U3031 ( .B1(n3042), .B2(n2378), .A(n2160), .ZN(n3981) );
  NAND2_X1 U3032 ( .A1(n2375), .A2(n2374), .ZN(n3046) );
  NAND2_X1 U3033 ( .A1(n3042), .A2(n2160), .ZN(n2375) );
  NAND2_X1 U3034 ( .A1(n4471), .A2(n4136), .ZN(n2381) );
  NAND3_X1 U3035 ( .A1(n2386), .A2(n2384), .A3(n4221), .ZN(n3699) );
  NAND3_X1 U3036 ( .A1(n2164), .A2(n4219), .A3(n3502), .ZN(n2386) );
  OAI21_X1 U3037 ( .B1(n3502), .B2(n3038), .A(n4219), .ZN(n3596) );
  NAND3_X2 U3038 ( .A1(n2478), .A2(n2476), .A3(n2477), .ZN(n2991) );
  NAND4_X1 U3039 ( .A1(n3035), .A2(n3629), .A3(n4206), .A4(n3537), .ZN(n3641)
         );
  AOI21_X1 U3040 ( .B1(n4657), .B2(n2397), .A(n2393), .ZN(n4527) );
  OAI21_X1 U3041 ( .B1(n4411), .B2(n4747), .A(n3081), .ZN(n3082) );
  INV_X1 U3042 ( .A(n4852), .ZN(n4855) );
  NAND2_X1 U3043 ( .A1(n3779), .A2(n3778), .ZN(n3881) );
  AOI21_X1 U3044 ( .B1(n4882), .B2(n4881), .A(n4880), .ZN(n4888) );
  NAND2_X1 U3045 ( .A1(n2518), .A2(n4299), .ZN(n2446) );
  AND2_X1 U3046 ( .A1(n3410), .A2(n4833), .ZN(n3411) );
  XNOR2_X1 U3047 ( .A(n3410), .B(n3409), .ZN(n4831) );
  XNOR2_X1 U3048 ( .A(n3540), .B(n4814), .ZN(n3451) );
  NAND4_X4 U3049 ( .A1(n2514), .A2(n2513), .A3(n2512), .A4(n2511), .ZN(n3504)
         );
  OR2_X1 U3050 ( .A1(n2509), .A2(n4293), .ZN(n2457) );
  INV_X1 U3051 ( .A(n3989), .ZN(n4646) );
  INV_X1 U3052 ( .A(n2967), .ZN(n2926) );
  NAND2_X1 U3053 ( .A1(n2967), .A2(IR_REG_31__SCAN_IN), .ZN(n2440) );
  NAND2_X1 U3054 ( .A1(n2429), .A2(n2447), .ZN(n2967) );
  NAND2_X1 U3055 ( .A1(n2414), .A2(n2499), .ZN(n2500) );
  OR2_X1 U3056 ( .A1(n2453), .A2(n2763), .ZN(n2451) );
  AND2_X1 U3057 ( .A1(n2991), .A2(n3537), .ZN(n3638) );
  INV_X1 U3058 ( .A(n2990), .ZN(n2989) );
  OAI21_X2 U3059 ( .B1(n2571), .B2(n2443), .A(n2480), .ZN(n3537) );
  INV_X2 U3060 ( .A(n2518), .ZN(n2571) );
  OAI21_X1 U3061 ( .B1(n3699), .B2(n3040), .A(n4225), .ZN(n3727) );
  NAND2_X1 U3062 ( .A1(n2982), .A2(n2952), .ZN(n4109) );
  INV_X1 U3063 ( .A(n4109), .ZN(n2953) );
  AND3_X1 U3064 ( .A1(n2954), .A2(n2403), .A3(n2953), .ZN(n2400) );
  AND2_X1 U3065 ( .A1(n2831), .A2(n4037), .ZN(n2401) );
  AND2_X1 U3066 ( .A1(n2805), .A2(n2804), .ZN(n2402) );
  OR2_X1 U3067 ( .A1(n2922), .A2(n2921), .ZN(n2403) );
  AND2_X1 U3068 ( .A1(n4132), .A2(n4131), .ZN(n2404) );
  OR2_X1 U3069 ( .A1(n2133), .A2(n3680), .ZN(n2405) );
  AND2_X1 U3070 ( .A1(n4846), .A2(REG2_REG_13__SCAN_IN), .ZN(n2407) );
  INV_X1 U3071 ( .A(n4815), .ZN(n3413) );
  INV_X1 U3072 ( .A(n3811), .ZN(n3006) );
  OR2_X1 U3073 ( .A1(n3447), .A2(REG1_REG_7__SCAN_IN), .ZN(n2408) );
  INV_X1 U3074 ( .A(n4160), .ZN(n3056) );
  AND3_X1 U3075 ( .A1(n4678), .A2(n4677), .A3(n4744), .ZN(n2409) );
  XNOR2_X1 U3076 ( .A(n2612), .B(IR_REG_8__SCAN_IN), .ZN(n4814) );
  AND2_X1 U3077 ( .A1(n3078), .A2(n3077), .ZN(n2410) );
  INV_X1 U3078 ( .A(n2955), .ZN(n2954) );
  INV_X1 U3079 ( .A(REG3_REG_9__SCAN_IN), .ZN(n2617) );
  INV_X1 U3080 ( .A(REG3_REG_13__SCAN_IN), .ZN(n2671) );
  AND2_X1 U3081 ( .A1(n4290), .A2(n3706), .ZN(n2411) );
  NAND2_X1 U3082 ( .A1(n2581), .A2(n2580), .ZN(n2412) );
  INV_X1 U3083 ( .A(n3831), .ZN(n3069) );
  INV_X1 U3084 ( .A(n4928), .ZN(n4344) );
  AND2_X1 U3085 ( .A1(n4862), .A2(REG2_REG_15__SCAN_IN), .ZN(n2413) );
  INV_X1 U3086 ( .A(IR_REG_10__SCAN_IN), .ZN(n2419) );
  AND2_X1 U3087 ( .A1(n3960), .A2(n3044), .ZN(n4245) );
  INV_X1 U3088 ( .A(n3571), .ZN(n2597) );
  AND2_X1 U3089 ( .A1(n4158), .A2(n4436), .ZN(n4263) );
  AND2_X1 U3090 ( .A1(n2703), .A2(n3865), .ZN(n2704) );
  INV_X1 U3091 ( .A(n2750), .ZN(n2751) );
  INV_X1 U3092 ( .A(n2749), .ZN(n2752) );
  OR2_X1 U3093 ( .A1(n3050), .A2(n4565), .ZN(n4546) );
  AND2_X1 U3094 ( .A1(n2448), .A2(IR_REG_27__SCAN_IN), .ZN(n2439) );
  INV_X1 U3095 ( .A(IR_REG_12__SCAN_IN), .ZN(n3133) );
  NAND2_X1 U3096 ( .A1(n2556), .A2(n2576), .ZN(n2578) );
  INV_X1 U3097 ( .A(n3118), .ZN(n2455) );
  NAND2_X1 U3098 ( .A1(n2262), .A2(n4809), .ZN(n4339) );
  INV_X1 U3099 ( .A(n3700), .ZN(n3706) );
  OAI22_X1 U3100 ( .A1(n4651), .A2(n2913), .B1(n3986), .B2(n2135), .ZN(n3904)
         );
  OR2_X1 U3101 ( .A1(n4504), .A2(n2133), .ZN(n2848) );
  INV_X1 U3102 ( .A(REG1_REG_18__SCAN_IN), .ZN(n4364) );
  OR2_X1 U3103 ( .A1(n4029), .A2(n2133), .ZN(n2799) );
  INV_X1 U3104 ( .A(n4443), .ZN(n4268) );
  OR2_X1 U3105 ( .A1(n3531), .A2(n3062), .ZN(n3494) );
  INV_X1 U3106 ( .A(n3734), .ZN(n3070) );
  OR2_X1 U3107 ( .A1(n2157), .A2(IR_REG_22__SCAN_IN), .ZN(n2923) );
  INV_X2 U3108 ( .A(IR_REG_2__SCAN_IN), .ZN(n2515) );
  OR2_X1 U3109 ( .A1(n2631), .A2(n2630), .ZN(n2650) );
  INV_X1 U3110 ( .A(n4521), .ZN(n4514) );
  INV_X1 U3111 ( .A(n3409), .ZN(n4833) );
  INV_X1 U3112 ( .A(REG3_REG_10__SCAN_IN), .ZN(n3659) );
  INV_X1 U3113 ( .A(n3990), .ZN(n3986) );
  AOI21_X1 U3114 ( .B1(n3579), .B2(n2995), .A(n2994), .ZN(n3491) );
  INV_X1 U3115 ( .A(n3664), .ZN(n3068) );
  OR2_X1 U3116 ( .A1(n2948), .A2(n2137), .ZN(n4627) );
  INV_X1 U3117 ( .A(n4627), .ZN(n4661) );
  INV_X1 U3118 ( .A(n3757), .ZN(n3852) );
  INV_X1 U3119 ( .A(n4623), .ZN(n4901) );
  NAND2_X1 U3120 ( .A1(n2946), .A2(n2945), .ZN(n2944) );
  INV_X1 U3121 ( .A(n2764), .ZN(n2765) );
  INV_X1 U3122 ( .A(n4122), .ZN(n4086) );
  AND2_X1 U3123 ( .A1(n3079), .A2(n2943), .ZN(n2982) );
  NAND2_X1 U3124 ( .A1(n2812), .A2(n2811), .ZN(n4574) );
  NAND2_X1 U3125 ( .A1(n2494), .A2(REG2_REG_11__SCAN_IN), .ZN(n2662) );
  NAND2_X1 U3126 ( .A1(n4297), .A2(n3379), .ZN(n4318) );
  NAND2_X1 U3127 ( .A1(n4886), .A2(n4885), .ZN(n4887) );
  AND2_X1 U3128 ( .A1(n4823), .A2(n4309), .ZN(n4893) );
  INV_X1 U3129 ( .A(n4655), .ZN(n4898) );
  AND2_X1 U3130 ( .A1(n3499), .A2(n4376), .ZN(n4600) );
  AND2_X1 U3131 ( .A1(n4600), .A2(n4943), .ZN(n4664) );
  AND2_X1 U3132 ( .A1(n2931), .A2(n2930), .ZN(n3079) );
  INV_X1 U3133 ( .A(n4164), .ZN(n3086) );
  INV_X1 U3134 ( .A(n3079), .ZN(n3497) );
  INV_X1 U3135 ( .A(IR_REG_24__SCAN_IN), .ZN(n2924) );
  OAI21_X1 U3136 ( .B1(n2946), .B2(n2945), .A(n2944), .ZN(n3381) );
  XNOR2_X1 U3137 ( .A(n2610), .B(n2609), .ZN(n3446) );
  AND2_X1 U3138 ( .A1(n3392), .A2(n3391), .ZN(n4883) );
  NOR2_X1 U3139 ( .A1(n2956), .A2(n2986), .ZN(n2987) );
  AND2_X1 U3140 ( .A1(n2966), .A2(n3530), .ZN(n4122) );
  NAND2_X1 U3141 ( .A1(n2825), .A2(n2824), .ZN(n4553) );
  INV_X1 U3142 ( .A(n4893), .ZN(n4856) );
  NAND2_X1 U3143 ( .A1(n4485), .A2(n3594), .ZN(n4666) );
  INV_X1 U3144 ( .A(n4664), .ZN(n4639) );
  NAND2_X1 U3145 ( .A1(n4975), .A2(n4943), .ZN(n4747) );
  AND2_X1 U3146 ( .A1(n3080), .A2(n3497), .ZN(n4798) );
  INV_X1 U3147 ( .A(n4798), .ZN(n4965) );
  INV_X1 U31480 ( .A(n4921), .ZN(n4923) );
  AND2_X1 U31490 ( .A1(n3381), .A2(STATE_REG_SCAN_IN), .ZN(n4924) );
  XNOR2_X1 U3150 ( .A(n2746), .B(n2745), .ZN(n4928) );
  CLKBUF_X2 U3151 ( .A(n3521), .Z(U4043) );
  OAI21_X1 U3152 ( .B1(n4671), .B2(n4802), .A(n3093), .ZN(U3517) );
  NOR2_X2 U3153 ( .A1(IR_REG_0__SCAN_IN), .A2(IR_REG_4__SCAN_IN), .ZN(n2415)
         );
  NAND4_X1 U3154 ( .A1(n2417), .A2(n2730), .A3(n2416), .A4(n3133), .ZN(n2418)
         );
  NAND4_X1 U3155 ( .A1(n2690), .A2(n3154), .A3(n2419), .A4(n2714), .ZN(n2420)
         );
  NOR2_X1 U3156 ( .A1(IR_REG_21__SCAN_IN), .A2(IR_REG_18__SCAN_IN), .ZN(n2425)
         );
  NOR2_X1 U3157 ( .A1(IR_REG_22__SCAN_IN), .A2(IR_REG_23__SCAN_IN), .ZN(n2424)
         );
  NAND4_X1 U3158 ( .A1(n2431), .A2(n2425), .A3(n2424), .A4(n2924), .ZN(n2450)
         );
  NOR2_X1 U3159 ( .A1(n2429), .A2(n2763), .ZN(n2426) );
  MUX2_X1 U3160 ( .A(n2763), .B(n2426), .S(IR_REG_25__SCAN_IN), .Z(n2927) );
  NAND2_X1 U3161 ( .A1(IR_REG_24__SCAN_IN), .A2(IR_REG_23__SCAN_IN), .ZN(n2427) );
  OAI21_X1 U3162 ( .B1(IR_REG_24__SCAN_IN), .B2(IR_REG_23__SCAN_IN), .A(n2427), 
        .ZN(n2428) );
  NAND2_X1 U3163 ( .A1(n2433), .A2(n2431), .ZN(n2463) );
  XNOR2_X2 U3164 ( .A(n2432), .B(IR_REG_21__SCAN_IN), .ZN(n2469) );
  OR2_X1 U3165 ( .A1(n2763), .A2(n2466), .ZN(n2434) );
  NAND3_X1 U3166 ( .A1(n3087), .A2(IR_REG_31__SCAN_IN), .A3(IR_REG_26__SCAN_IN), .ZN(n2436) );
  OAI211_X1 U3167 ( .C1(IR_REG_31__SCAN_IN), .C2(n3087), .A(n2437), .B(n2436), 
        .ZN(n2438) );
  AOI21_X1 U3168 ( .B1(n2926), .B2(n2439), .A(n2438), .ZN(n2442) );
  AND2_X4 U3169 ( .A1(n2442), .A2(n2441), .ZN(n2518) );
  INV_X2 U3170 ( .A(IR_REG_0__SCAN_IN), .ZN(n2443) );
  NAND2_X1 U3171 ( .A1(n2414), .A2(n2472), .ZN(n2462) );
  NAND4_X1 U3172 ( .A1(n3087), .A2(n2448), .A3(n2969), .A4(n2447), .ZN(n2449)
         );
  NAND2_X1 U3173 ( .A1(n2453), .A2(n2452), .ZN(n4016) );
  INV_X1 U3174 ( .A(REG3_REG_1__SCAN_IN), .ZN(n3630) );
  OR2_X1 U3175 ( .A1(n2493), .A2(n3630), .ZN(n2460) );
  INV_X1 U3176 ( .A(REG2_REG_1__SCAN_IN), .ZN(n3653) );
  INV_X1 U3177 ( .A(REG1_REG_1__SCAN_IN), .ZN(n4293) );
  NAND2_X1 U3178 ( .A1(n2990), .A2(n2549), .ZN(n2461) );
  NAND2_X1 U3179 ( .A1(n2462), .A2(n2461), .ZN(n2467) );
  NAND2_X1 U3180 ( .A1(n2468), .A2(n4376), .ZN(n2964) );
  INV_X1 U3181 ( .A(n2468), .ZN(n2947) );
  INV_X1 U3182 ( .A(n2469), .ZN(n4203) );
  NAND2_X1 U3183 ( .A1(n2947), .A2(n4203), .ZN(n2948) );
  INV_X1 U3184 ( .A(n2948), .ZN(n2471) );
  INV_X1 U3185 ( .A(n2137), .ZN(n4807) );
  INV_X1 U3186 ( .A(n2525), .ZN(n2601) );
  INV_X1 U3187 ( .A(REG0_REG_0__SCAN_IN), .ZN(n2473) );
  OR2_X1 U3188 ( .A1(n2134), .A2(n2473), .ZN(n2477) );
  INV_X1 U3189 ( .A(REG1_REG_0__SCAN_IN), .ZN(n4968) );
  AND2_X1 U3190 ( .A1(n2475), .A2(n2474), .ZN(n2476) );
  INV_X1 U3191 ( .A(DATAI_0_), .ZN(n2479) );
  INV_X1 U3192 ( .A(n2962), .ZN(n3094) );
  AOI22_X1 U3193 ( .A1(n2549), .A2(n3537), .B1(n3094), .B2(IR_REG_0__SCAN_IN), 
        .ZN(n2481) );
  OAI21_X1 U3194 ( .B1(n2645), .B2(n3629), .A(n2481), .ZN(n3534) );
  NAND2_X1 U3195 ( .A1(n2991), .A2(n2549), .ZN(n2484) );
  NAND2_X1 U3196 ( .A1(n2414), .A2(n3537), .ZN(n2485) );
  OR2_X1 U3197 ( .A1(n2962), .A2(n4968), .ZN(n2482) );
  AND2_X1 U3198 ( .A1(n2485), .A2(n2482), .ZN(n2483) );
  NAND2_X1 U3199 ( .A1(n2484), .A2(n2483), .ZN(n3535) );
  NAND2_X1 U3200 ( .A1(n3534), .A2(n3535), .ZN(n2488) );
  INV_X1 U3201 ( .A(n2485), .ZN(n2486) );
  OR2_X1 U3202 ( .A1(n2914), .A2(n2486), .ZN(n2487) );
  NAND2_X1 U3203 ( .A1(n2488), .A2(n2487), .ZN(n3628) );
  INV_X1 U3204 ( .A(n2489), .ZN(n2490) );
  NOR2_X1 U3205 ( .A1(n2491), .A2(n2490), .ZN(n2492) );
  INV_X1 U3206 ( .A(REG3_REG_2__SCAN_IN), .ZN(n3680) );
  NAND2_X1 U3207 ( .A1(n2494), .A2(REG2_REG_2__SCAN_IN), .ZN(n2497) );
  INV_X1 U3208 ( .A(REG1_REG_2__SCAN_IN), .ZN(n3387) );
  NAND2_X1 U3209 ( .A1(n3643), .A2(n2549), .ZN(n2501) );
  XNOR2_X2 U32100 ( .A(n2498), .B(n2515), .ZN(n3386) );
  MUX2_X1 U32110 ( .A(n3386), .B(n3113), .S(n2571), .Z(n2992) );
  INV_X1 U32120 ( .A(n2992), .ZN(n2499) );
  NAND2_X1 U32130 ( .A1(n2501), .A2(n2500), .ZN(n2502) );
  XNOR2_X1 U32140 ( .A(n2502), .B(n2849), .ZN(n2505) );
  NOR2_X1 U32150 ( .A1(n2136), .A2(n2992), .ZN(n2503) );
  AOI21_X1 U32160 ( .B1(n2504), .B2(n3643), .A(n2503), .ZN(n2506) );
  OR2_X1 U32170 ( .A1(n2505), .A2(n2506), .ZN(n2507) );
  NAND2_X1 U32180 ( .A1(n2506), .A2(n2505), .ZN(n2508) );
  AND2_X1 U32190 ( .A1(n2507), .A2(n2508), .ZN(n3557) );
  NAND2_X1 U32200 ( .A1(n3558), .A2(n3557), .ZN(n3556) );
  NAND2_X1 U32210 ( .A1(n3556), .A2(n2508), .ZN(n3622) );
  OR2_X1 U32220 ( .A1(n2132), .A2(REG3_REG_3__SCAN_IN), .ZN(n2513) );
  INV_X1 U32230 ( .A(REG2_REG_3__SCAN_IN), .ZN(n3588) );
  OR2_X1 U32240 ( .A1(n3465), .A2(n3588), .ZN(n2512) );
  INV_X1 U32250 ( .A(REG0_REG_3__SCAN_IN), .ZN(n2510) );
  OR2_X1 U32260 ( .A1(n2601), .A2(n2510), .ZN(n2511) );
  NAND2_X1 U32270 ( .A1(n3504), .A2(n2138), .ZN(n2520) );
  NAND2_X1 U32280 ( .A1(n2516), .A2(n2515), .ZN(n2517) );
  MUX2_X1 U32290 ( .A(n4817), .B(DATAI_3_), .S(n3085), .Z(n3590) );
  NAND2_X1 U32300 ( .A1(n2414), .A2(n3590), .ZN(n2519) );
  NAND2_X1 U32310 ( .A1(n2520), .A2(n2519), .ZN(n2521) );
  INV_X1 U32320 ( .A(n3504), .ZN(n3677) );
  INV_X1 U32330 ( .A(n3590), .ZN(n3617) );
  OAI22_X1 U32340 ( .A1(n2645), .A2(n3677), .B1(n3617), .B2(n2136), .ZN(n2523)
         );
  XNOR2_X1 U32350 ( .A(n2522), .B(n2523), .ZN(n3623) );
  NAND2_X1 U32360 ( .A1(n3622), .A2(n3623), .ZN(n3621) );
  INV_X1 U32370 ( .A(n2522), .ZN(n2524) );
  OR2_X1 U32380 ( .A1(n2524), .A2(n2523), .ZN(n3611) );
  NAND2_X1 U32390 ( .A1(n2525), .A2(REG0_REG_4__SCAN_IN), .ZN(n2529) );
  INV_X1 U32400 ( .A(REG1_REG_4__SCAN_IN), .ZN(n4830) );
  OR2_X1 U32410 ( .A1(n2509), .A2(n4830), .ZN(n2528) );
  XNOR2_X1 U32420 ( .A(REG3_REG_4__SCAN_IN), .B(REG3_REG_3__SCAN_IN), .ZN(
        n3616) );
  OR2_X1 U32430 ( .A1(n2132), .A2(n3616), .ZN(n2527) );
  INV_X1 U32440 ( .A(REG2_REG_4__SCAN_IN), .ZN(n4828) );
  OR2_X1 U32450 ( .A1(n3465), .A2(n4828), .ZN(n2526) );
  NAND4_X1 U32460 ( .A1(n2529), .A2(n2528), .A3(n2527), .A4(n2526), .ZN(n3620)
         );
  INV_X1 U32470 ( .A(n3620), .ZN(n3597) );
  NAND2_X1 U32480 ( .A1(n2531), .A2(n2530), .ZN(n2532) );
  NAND2_X1 U32490 ( .A1(n2532), .A2(IR_REG_31__SCAN_IN), .ZN(n2534) );
  INV_X1 U32500 ( .A(IR_REG_4__SCAN_IN), .ZN(n2533) );
  INV_X1 U32510 ( .A(DATAI_4_), .ZN(n3109) );
  MUX2_X1 U32520 ( .A(n3409), .B(n3109), .S(n2571), .Z(n3609) );
  NAND2_X1 U32530 ( .A1(n3620), .A2(n2138), .ZN(n2537) );
  OR2_X1 U32540 ( .A1(n2916), .A2(n3609), .ZN(n2536) );
  NAND2_X1 U32550 ( .A1(n2537), .A2(n2536), .ZN(n2538) );
  XNOR2_X1 U32560 ( .A(n2538), .B(n2849), .ZN(n2557) );
  XNOR2_X1 U32570 ( .A(n2558), .B(n2557), .ZN(n3612) );
  AND2_X1 U32580 ( .A1(n3611), .A2(n3612), .ZN(n2539) );
  NAND2_X1 U32590 ( .A1(n3621), .A2(n2539), .ZN(n3563) );
  INV_X1 U32600 ( .A(REG3_REG_5__SCAN_IN), .ZN(n2541) );
  NAND2_X1 U32610 ( .A1(REG3_REG_4__SCAN_IN), .A2(REG3_REG_3__SCAN_IN), .ZN(
        n2540) );
  NAND2_X1 U32620 ( .A1(n2541), .A2(n2540), .ZN(n2542) );
  NAND2_X1 U32630 ( .A1(n2562), .A2(n2542), .ZN(n3604) );
  OR2_X1 U32640 ( .A1(n2132), .A2(n3604), .ZN(n2548) );
  NAND2_X1 U32650 ( .A1(n2525), .A2(REG0_REG_5__SCAN_IN), .ZN(n2547) );
  INV_X1 U32660 ( .A(REG1_REG_5__SCAN_IN), .ZN(n2543) );
  OR2_X1 U32670 ( .A1(n2509), .A2(n2543), .ZN(n2546) );
  INV_X1 U32680 ( .A(REG2_REG_5__SCAN_IN), .ZN(n2544) );
  OR2_X1 U32690 ( .A1(n3465), .A2(n2544), .ZN(n2545) );
  NAND2_X1 U32700 ( .A1(n3830), .A2(n2549), .ZN(n2553) );
  NAND2_X1 U32710 ( .A1(n2550), .A2(IR_REG_31__SCAN_IN), .ZN(n2551) );
  MUX2_X1 U32720 ( .A(n4816), .B(DATAI_5_), .S(n3085), .Z(n2998) );
  NAND2_X1 U32730 ( .A1(n2414), .A2(n2998), .ZN(n2552) );
  NAND2_X1 U32740 ( .A1(n2553), .A2(n2552), .ZN(n2554) );
  INV_X1 U32750 ( .A(n2577), .ZN(n2556) );
  INV_X1 U32760 ( .A(n3830), .ZN(n2555) );
  OAI22_X1 U32770 ( .A1(n2645), .A2(n2555), .B1(n3602), .B2(n2135), .ZN(n2576)
         );
  INV_X1 U32780 ( .A(n2557), .ZN(n2559) );
  NAND2_X1 U32790 ( .A1(n2559), .A2(n2558), .ZN(n3564) );
  AND2_X1 U32800 ( .A1(n2578), .A2(n3564), .ZN(n3824) );
  INV_X1 U32810 ( .A(REG1_REG_6__SCAN_IN), .ZN(n3420) );
  INV_X1 U32820 ( .A(n2583), .ZN(n2585) );
  INV_X1 U32830 ( .A(REG3_REG_6__SCAN_IN), .ZN(n2561) );
  NAND2_X1 U32840 ( .A1(n2562), .A2(n2561), .ZN(n2563) );
  NAND2_X1 U32850 ( .A1(n2585), .A2(n2563), .ZN(n3834) );
  OR2_X1 U32860 ( .A1(n2133), .A2(n3834), .ZN(n2567) );
  NAND2_X1 U32870 ( .A1(n2525), .A2(REG0_REG_6__SCAN_IN), .ZN(n2566) );
  INV_X1 U32880 ( .A(REG2_REG_6__SCAN_IN), .ZN(n2564) );
  OR2_X1 U32890 ( .A1(n3465), .A2(n2564), .ZN(n2565) );
  NAND2_X1 U32900 ( .A1(n4291), .A2(n2138), .ZN(n2573) );
  INV_X1 U32910 ( .A(IR_REG_31__SCAN_IN), .ZN(n2763) );
  OR2_X1 U32920 ( .A1(n2625), .A2(n2763), .ZN(n2570) );
  XNOR2_X1 U32930 ( .A(n2570), .B(IR_REG_6__SCAN_IN), .ZN(n4815) );
  MUX2_X1 U32940 ( .A(n4815), .B(DATAI_6_), .S(n3085), .Z(n3831) );
  NAND2_X1 U32950 ( .A1(n2414), .A2(n3831), .ZN(n2572) );
  NAND2_X1 U32960 ( .A1(n2573), .A2(n2572), .ZN(n2574) );
  XNOR2_X1 U32970 ( .A(n2574), .B(n2914), .ZN(n2581) );
  INV_X1 U32980 ( .A(n4291), .ZN(n3714) );
  OAI22_X1 U32990 ( .A1(n2913), .A2(n3714), .B1(n3069), .B2(n2135), .ZN(n2580)
         );
  AND2_X1 U33000 ( .A1(n3824), .A2(n2412), .ZN(n2575) );
  XNOR2_X1 U33010 ( .A(n2577), .B(n2576), .ZN(n3562) );
  INV_X1 U33020 ( .A(n3562), .ZN(n2579) );
  NAND2_X1 U33030 ( .A1(n2579), .A2(n2578), .ZN(n3825) );
  INV_X1 U33040 ( .A(n3825), .ZN(n2582) );
  OR2_X1 U33050 ( .A1(n2581), .A2(n2580), .ZN(n3826) );
  INV_X1 U33060 ( .A(REG3_REG_7__SCAN_IN), .ZN(n2584) );
  NAND2_X1 U33070 ( .A1(n2585), .A2(n2584), .ZN(n2586) );
  NAND2_X1 U33080 ( .A1(n2603), .A2(n2586), .ZN(n3709) );
  OR2_X1 U33090 ( .A1(n2132), .A2(n3709), .ZN(n2591) );
  NAND2_X1 U33100 ( .A1(n2525), .A2(REG0_REG_7__SCAN_IN), .ZN(n2589) );
  INV_X1 U33110 ( .A(REG2_REG_7__SCAN_IN), .ZN(n2587) );
  OR2_X1 U33120 ( .A1(n3465), .A2(n2587), .ZN(n2588) );
  NAND2_X1 U33130 ( .A1(n4290), .A2(n2549), .ZN(n2595) );
  NAND2_X1 U33140 ( .A1(n2625), .A2(n2592), .ZN(n2593) );
  NAND2_X1 U33150 ( .A1(n2593), .A2(IR_REG_31__SCAN_IN), .ZN(n2610) );
  INV_X1 U33160 ( .A(DATAI_7_), .ZN(n3111) );
  MUX2_X1 U33170 ( .A(n3446), .B(n3111), .S(n3085), .Z(n3700) );
  OR2_X1 U33180 ( .A1(n2916), .A2(n3700), .ZN(n2594) );
  NAND2_X1 U33190 ( .A1(n2595), .A2(n2594), .ZN(n2596) );
  XNOR2_X1 U33200 ( .A(n2596), .B(n2914), .ZN(n2599) );
  INV_X1 U33210 ( .A(n4290), .ZN(n3732) );
  OAI22_X1 U33220 ( .A1(n2913), .A2(n3732), .B1(n3700), .B2(n2136), .ZN(n2598)
         );
  XNOR2_X1 U33230 ( .A(n2599), .B(n2598), .ZN(n3571) );
  NAND2_X1 U33240 ( .A1(n2599), .A2(n2598), .ZN(n2600) );
  NAND2_X1 U33250 ( .A1(n2972), .A2(REG1_REG_8__SCAN_IN), .ZN(n2608) );
  INV_X1 U33260 ( .A(REG0_REG_8__SCAN_IN), .ZN(n3267) );
  OR2_X1 U33270 ( .A1(n2601), .A2(n3267), .ZN(n2607) );
  INV_X1 U33280 ( .A(REG3_REG_8__SCAN_IN), .ZN(n2602) );
  NAND2_X1 U33290 ( .A1(n2603), .A2(n2602), .ZN(n2604) );
  NAND2_X1 U33300 ( .A1(n2618), .A2(n2604), .ZN(n3735) );
  OR2_X1 U33310 ( .A1(n2132), .A2(n3735), .ZN(n2606) );
  INV_X1 U33320 ( .A(REG2_REG_8__SCAN_IN), .ZN(n3736) );
  OR2_X1 U33330 ( .A1(n3465), .A2(n3736), .ZN(n2605) );
  NAND2_X1 U33340 ( .A1(n3796), .A2(n2549), .ZN(n2614) );
  NAND2_X1 U33350 ( .A1(n2610), .A2(n2609), .ZN(n2611) );
  NAND2_X1 U33360 ( .A1(n2611), .A2(IR_REG_31__SCAN_IN), .ZN(n2612) );
  MUX2_X1 U33370 ( .A(n4814), .B(DATAI_8_), .S(n3085), .Z(n3734) );
  NAND2_X1 U33380 ( .A1(n2414), .A2(n3734), .ZN(n2613) );
  NAND2_X1 U33390 ( .A1(n2614), .A2(n2613), .ZN(n2615) );
  XNOR2_X1 U33400 ( .A(n2615), .B(n2914), .ZN(n3686) );
  INV_X1 U33410 ( .A(n3796), .ZN(n2616) );
  OAI22_X1 U33420 ( .A1(n2913), .A2(n2616), .B1(n3070), .B2(n2136), .ZN(n3687)
         );
  AND2_X1 U33430 ( .A1(n3686), .A2(n3687), .ZN(n2631) );
  NAND2_X1 U33440 ( .A1(n2972), .A2(REG1_REG_9__SCAN_IN), .ZN(n2623) );
  INV_X1 U33450 ( .A(REG0_REG_9__SCAN_IN), .ZN(n3271) );
  OR2_X1 U33460 ( .A1(n2601), .A2(n3271), .ZN(n2622) );
  NAND2_X1 U33470 ( .A1(n2618), .A2(n2617), .ZN(n2619) );
  NAND2_X1 U33480 ( .A1(n2634), .A2(n2619), .ZN(n3695) );
  OR2_X1 U33490 ( .A1(n2133), .A2(n3695), .ZN(n2621) );
  INV_X1 U33500 ( .A(REG2_REG_9__SCAN_IN), .ZN(n3800) );
  OR2_X1 U33510 ( .A1(n3465), .A2(n3800), .ZN(n2620) );
  NAND2_X1 U33520 ( .A1(n3811), .A2(n2549), .ZN(n2628) );
  INV_X1 U3353 ( .A(n3128), .ZN(n2624) );
  NAND2_X1 U33540 ( .A1(n2625), .A2(n2624), .ZN(n2640) );
  NAND2_X1 U3355 ( .A1(n2640), .A2(IR_REG_31__SCAN_IN), .ZN(n2626) );
  MUX2_X1 U3356 ( .A(n4813), .B(DATAI_9_), .S(n3085), .Z(n3005) );
  NAND2_X1 U3357 ( .A1(n2414), .A2(n3005), .ZN(n2627) );
  NAND2_X1 U3358 ( .A1(n2628), .A2(n2627), .ZN(n2629) );
  XNOR2_X1 U3359 ( .A(n2629), .B(n2914), .ZN(n3685) );
  OAI22_X1 U3360 ( .A1(n2913), .A2(n3006), .B1(n3801), .B2(n2135), .ZN(n3684)
         );
  AND2_X1 U3361 ( .A1(n3685), .A2(n3684), .ZN(n2630) );
  OAI21_X1 U3362 ( .B1(n3686), .B2(n3687), .A(n3684), .ZN(n2632) );
  INV_X1 U3363 ( .A(n3685), .ZN(n3763) );
  NAND2_X1 U3364 ( .A1(n2632), .A2(n3763), .ZN(n2648) );
  NAND2_X1 U3365 ( .A1(n2525), .A2(REG0_REG_10__SCAN_IN), .ZN(n2639) );
  INV_X1 U3366 ( .A(REG1_REG_10__SCAN_IN), .ZN(n2633) );
  OR2_X1 U3367 ( .A1(n3462), .A2(n2633), .ZN(n2638) );
  NAND2_X1 U3368 ( .A1(n2634), .A2(n3659), .ZN(n2635) );
  NAND2_X1 U3369 ( .A1(n2659), .A2(n2635), .ZN(n3818) );
  OR2_X1 U3370 ( .A1(n2132), .A2(n3818), .ZN(n2637) );
  INV_X1 U3371 ( .A(REG2_REG_10__SCAN_IN), .ZN(n3819) );
  OR2_X1 U3372 ( .A1(n3465), .A2(n3819), .ZN(n2636) );
  NAND2_X1 U3373 ( .A1(n4289), .A2(n2138), .ZN(n2643) );
  NAND2_X1 U3374 ( .A1(n2655), .A2(IR_REG_31__SCAN_IN), .ZN(n2641) );
  XNOR2_X1 U3375 ( .A(n2641), .B(IR_REG_10__SCAN_IN), .ZN(n3773) );
  MUX2_X1 U3376 ( .A(n3773), .B(DATAI_10_), .S(n3085), .Z(n3817) );
  NAND2_X1 U3377 ( .A1(n2414), .A2(n3817), .ZN(n2642) );
  NAND2_X1 U3378 ( .A1(n2643), .A2(n2642), .ZN(n2644) );
  XNOR2_X1 U3379 ( .A(n2644), .B(n2849), .ZN(n2651) );
  INV_X2 U3380 ( .A(n2504), .ZN(n2913) );
  INV_X1 U3381 ( .A(n4289), .ZN(n3794) );
  OAI22_X1 U3382 ( .A1(n2913), .A2(n3794), .B1(n2237), .B2(n2136), .ZN(n2652)
         );
  XNOR2_X1 U3383 ( .A(n2651), .B(n2652), .ZN(n3765) );
  INV_X1 U3384 ( .A(n3687), .ZN(n3689) );
  INV_X1 U3385 ( .A(n3684), .ZN(n3762) );
  INV_X1 U3386 ( .A(n3686), .ZN(n2646) );
  NAND3_X1 U3387 ( .A1(n3689), .A2(n3762), .A3(n2646), .ZN(n2647) );
  AND3_X1 U3388 ( .A1(n2648), .A2(n3765), .A3(n2647), .ZN(n2649) );
  OAI21_X2 U3389 ( .B1(n3522), .B2(n2650), .A(n2649), .ZN(n3764) );
  INV_X1 U3390 ( .A(n2651), .ZN(n2653) );
  NAND2_X1 U3391 ( .A1(n2653), .A2(n2652), .ZN(n2654) );
  NAND2_X1 U3392 ( .A1(n3764), .A2(n2654), .ZN(n3752) );
  INV_X1 U3393 ( .A(DATAI_11_), .ZN(n2656) );
  MUX2_X1 U3394 ( .A(n4811), .B(n2656), .S(n3085), .Z(n3757) );
  NAND2_X1 U3395 ( .A1(n3852), .A2(n2414), .ZN(n2666) );
  INV_X1 U3396 ( .A(REG3_REG_11__SCAN_IN), .ZN(n2658) );
  NAND2_X1 U3397 ( .A1(n2659), .A2(n2658), .ZN(n2660) );
  NAND2_X1 U3398 ( .A1(n2683), .A2(n2660), .ZN(n3854) );
  OR2_X1 U3399 ( .A1(n2133), .A2(n3854), .ZN(n2664) );
  INV_X1 U3400 ( .A(REG1_REG_11__SCAN_IN), .ZN(n3954) );
  OR2_X1 U3401 ( .A1(n2509), .A2(n3954), .ZN(n2663) );
  NAND2_X1 U3402 ( .A1(n2525), .A2(REG0_REG_11__SCAN_IN), .ZN(n2661) );
  NAND2_X1 U3403 ( .A1(n4288), .A2(n2549), .ZN(n2665) );
  NAND2_X1 U3404 ( .A1(n2666), .A2(n2665), .ZN(n2667) );
  XNOR2_X1 U3405 ( .A(n2667), .B(n2914), .ZN(n2669) );
  OAI22_X1 U3406 ( .A1(n2913), .A2(n3918), .B1(n3757), .B2(n2136), .ZN(n2668)
         );
  OR2_X1 U3407 ( .A1(n2669), .A2(n2668), .ZN(n3754) );
  NAND2_X1 U3408 ( .A1(n3752), .A2(n3754), .ZN(n2670) );
  NAND2_X1 U3409 ( .A1(n2669), .A2(n2668), .ZN(n3753) );
  NAND2_X1 U3410 ( .A1(n2685), .A2(n2671), .ZN(n2672) );
  AND2_X1 U3411 ( .A1(n2707), .A2(n2672), .ZN(n3976) );
  NAND2_X1 U3412 ( .A1(n3976), .A2(n2898), .ZN(n2676) );
  NAND2_X1 U3413 ( .A1(n2494), .A2(REG2_REG_13__SCAN_IN), .ZN(n2675) );
  INV_X1 U3414 ( .A(REG0_REG_13__SCAN_IN), .ZN(n4795) );
  OR2_X1 U3415 ( .A1(n2601), .A2(n4795), .ZN(n2674) );
  INV_X1 U3416 ( .A(REG1_REG_13__SCAN_IN), .ZN(n4740) );
  OR2_X1 U3417 ( .A1(n3462), .A2(n4740), .ZN(n2673) );
  NAND4_X1 U3418 ( .A1(n2676), .A2(n2675), .A3(n2674), .A4(n2673), .ZN(n3983)
         );
  NAND2_X1 U3419 ( .A1(n3983), .A2(n2138), .ZN(n2680) );
  NOR2_X1 U3420 ( .A1(IR_REG_11__SCAN_IN), .A2(IR_REG_12__SCAN_IN), .ZN(n2715)
         );
  OR2_X1 U3421 ( .A1(n2715), .A2(n2763), .ZN(n2677) );
  NAND2_X1 U3422 ( .A1(n2691), .A2(n2677), .ZN(n2678) );
  MUX2_X1 U3423 ( .A(n4846), .B(DATAI_13_), .S(n3085), .Z(n3043) );
  NAND2_X1 U3424 ( .A1(n2414), .A2(n3043), .ZN(n2679) );
  NAND2_X1 U3425 ( .A1(n2680), .A2(n2679), .ZN(n2681) );
  XNOR2_X1 U3426 ( .A(n2681), .B(n2914), .ZN(n2700) );
  INV_X1 U3427 ( .A(n3983), .ZN(n3919) );
  NAND2_X1 U3428 ( .A1(n2549), .A2(n3043), .ZN(n2682) );
  OAI21_X1 U3429 ( .B1(n2913), .B2(n3919), .A(n2682), .ZN(n2699) );
  NAND2_X1 U3430 ( .A1(n2700), .A2(n2699), .ZN(n3864) );
  NAND2_X1 U3431 ( .A1(n2525), .A2(REG0_REG_12__SCAN_IN), .ZN(n2689) );
  INV_X1 U3432 ( .A(REG1_REG_12__SCAN_IN), .ZN(n4745) );
  OR2_X1 U3433 ( .A1(n3462), .A2(n4745), .ZN(n2688) );
  INV_X1 U3434 ( .A(REG3_REG_12__SCAN_IN), .ZN(n3244) );
  NAND2_X1 U3435 ( .A1(n2683), .A2(n3244), .ZN(n2684) );
  NAND2_X1 U3436 ( .A1(n2685), .A2(n2684), .ZN(n3932) );
  OR2_X1 U3437 ( .A1(n2132), .A2(n3932), .ZN(n2687) );
  OR2_X1 U3438 ( .A1(n3465), .A2(n3332), .ZN(n2686) );
  NAND2_X1 U3439 ( .A1(n4287), .A2(n2138), .ZN(n2695) );
  NAND2_X1 U3440 ( .A1(n2691), .A2(n2690), .ZN(n2692) );
  NAND2_X1 U3441 ( .A1(n2692), .A2(IR_REG_31__SCAN_IN), .ZN(n2693) );
  XNOR2_X1 U3442 ( .A(n2693), .B(IR_REG_12__SCAN_IN), .ZN(n4810) );
  MUX2_X1 U3443 ( .A(n4810), .B(DATAI_12_), .S(n3085), .Z(n3921) );
  NAND2_X1 U3444 ( .A1(n2414), .A2(n3921), .ZN(n2694) );
  NAND2_X1 U3445 ( .A1(n2695), .A2(n2694), .ZN(n2696) );
  XNOR2_X1 U3446 ( .A(n2696), .B(n2914), .ZN(n3867) );
  INV_X1 U3447 ( .A(n4287), .ZN(n3848) );
  OAI22_X1 U3448 ( .A1(n2913), .A2(n3848), .B1(n3930), .B2(n2136), .ZN(n3866)
         );
  NAND2_X1 U3449 ( .A1(n3867), .A2(n3866), .ZN(n2697) );
  NAND2_X1 U3450 ( .A1(n3864), .A2(n2697), .ZN(n2705) );
  INV_X1 U3451 ( .A(n3866), .ZN(n2698) );
  INV_X1 U3452 ( .A(n3867), .ZN(n3869) );
  NAND3_X1 U3453 ( .A1(n3864), .A2(n2698), .A3(n3869), .ZN(n2703) );
  INV_X1 U3454 ( .A(n2699), .ZN(n2702) );
  INV_X1 U3455 ( .A(n2700), .ZN(n2701) );
  NAND2_X1 U3456 ( .A1(n2702), .A2(n2701), .ZN(n3865) );
  INV_X1 U3457 ( .A(REG3_REG_14__SCAN_IN), .ZN(n3338) );
  NAND2_X1 U34580 ( .A1(n2707), .A2(n3338), .ZN(n2708) );
  NAND2_X1 U34590 ( .A1(n2726), .A2(n2708), .ZN(n3992) );
  OR2_X1 U3460 ( .A1(n3992), .A2(n2133), .ZN(n2713) );
  INV_X1 U3461 ( .A(REG0_REG_14__SCAN_IN), .ZN(n4791) );
  OR2_X1 U3462 ( .A1(n2601), .A2(n4791), .ZN(n2710) );
  INV_X1 U3463 ( .A(REG1_REG_14__SCAN_IN), .ZN(n4736) );
  OR2_X1 U3464 ( .A1(n3462), .A2(n4736), .ZN(n2709) );
  AND2_X1 U3465 ( .A1(n2710), .A2(n2709), .ZN(n2712) );
  INV_X1 U3466 ( .A(REG2_REG_14__SCAN_IN), .ZN(n3993) );
  OR2_X1 U34670 ( .A1(n3465), .A2(n3993), .ZN(n2711) );
  NAND2_X1 U3468 ( .A1(n2715), .A2(n2714), .ZN(n2716) );
  NOR2_X1 U34690 ( .A1(n2717), .A2(n2716), .ZN(n2731) );
  OR2_X1 U3470 ( .A1(n2731), .A2(n2763), .ZN(n2718) );
  MUX2_X1 U34710 ( .A(n4809), .B(DATAI_14_), .S(n3085), .Z(n3990) );
  OAI22_X1 U3472 ( .A1(n4651), .A2(n2136), .B1(n3986), .B2(n2916), .ZN(n2719)
         );
  XNOR2_X1 U34730 ( .A(n2719), .B(n2849), .ZN(n3905) );
  NAND2_X1 U3474 ( .A1(n3903), .A2(n3905), .ZN(n2720) );
  NAND2_X1 U34750 ( .A1(n2720), .A2(n3904), .ZN(n2724) );
  INV_X1 U3476 ( .A(n3903), .ZN(n2722) );
  INV_X1 U34770 ( .A(n3905), .ZN(n2721) );
  NAND2_X1 U3478 ( .A1(n2722), .A2(n2721), .ZN(n2723) );
  NAND2_X1 U34790 ( .A1(n2726), .A2(n2725), .ZN(n2727) );
  NAND2_X1 U3480 ( .A1(n2738), .A2(n2727), .ZN(n4648) );
  AOI22_X1 U34810 ( .A1(n2972), .A2(REG1_REG_15__SCAN_IN), .B1(n2525), .B2(
        REG0_REG_15__SCAN_IN), .ZN(n2729) );
  INV_X1 U3482 ( .A(REG2_REG_15__SCAN_IN), .ZN(n4649) );
  OR2_X1 U34830 ( .A1(n3465), .A2(n4649), .ZN(n2728) );
  OAI211_X1 U3484 ( .C1(n4648), .C2(n2133), .A(n2729), .B(n2728), .ZN(n4621)
         );
  NAND2_X1 U34850 ( .A1(n4621), .A2(n2138), .ZN(n2734) );
  NAND2_X1 U3486 ( .A1(n2731), .A2(n2730), .ZN(n2732) );
  NAND2_X1 U34870 ( .A1(n2732), .A2(IR_REG_31__SCAN_IN), .ZN(n2743) );
  XNOR2_X1 U3488 ( .A(n2743), .B(IR_REG_15__SCAN_IN), .ZN(n4862) );
  MUX2_X1 U34890 ( .A(DATAI_15_), .B(n4862), .S(n2518), .Z(n4660) );
  NAND2_X1 U3490 ( .A1(n4660), .A2(n2414), .ZN(n2733) );
  NAND2_X1 U34910 ( .A1(n2734), .A2(n2733), .ZN(n2735) );
  XNOR2_X1 U3492 ( .A(n2735), .B(n2914), .ZN(n2748) );
  AND2_X1 U34930 ( .A1(n4660), .A2(n2549), .ZN(n2736) );
  INV_X1 U3494 ( .A(REG3_REG_16__SCAN_IN), .ZN(n2737) );
  NAND2_X1 U34950 ( .A1(n2738), .A2(n2737), .ZN(n2739) );
  NAND2_X1 U3496 ( .A1(n2754), .A2(n2739), .ZN(n4636) );
  OR2_X1 U34970 ( .A1(n4636), .A2(n2132), .ZN(n2742) );
  AOI22_X1 U3498 ( .A1(n2972), .A2(REG1_REG_16__SCAN_IN), .B1(n2525), .B2(
        REG0_REG_16__SCAN_IN), .ZN(n2741) );
  NAND2_X1 U34990 ( .A1(n2494), .A2(REG2_REG_16__SCAN_IN), .ZN(n2740) );
  INV_X1 U3500 ( .A(DATAI_16_), .ZN(n4927) );
  NAND2_X1 U35010 ( .A1(n2743), .A2(n3154), .ZN(n2744) );
  NAND2_X1 U3502 ( .A1(n2744), .A2(IR_REG_31__SCAN_IN), .ZN(n2746) );
  INV_X1 U35030 ( .A(IR_REG_16__SCAN_IN), .ZN(n2745) );
  MUX2_X1 U3504 ( .A(n4927), .B(n4928), .S(n2518), .Z(n4633) );
  OAI22_X1 U35050 ( .A1(n4652), .A2(n2913), .B1(n4633), .B2(n2135), .ZN(n2750)
         );
  OAI22_X1 U35060 ( .A1(n4652), .A2(n2135), .B1(n4633), .B2(n2916), .ZN(n2747)
         );
  XNOR2_X1 U35070 ( .A(n2747), .B(n2914), .ZN(n2749) );
  INV_X1 U35080 ( .A(REG3_REG_17__SCAN_IN), .ZN(n2753) );
  NAND2_X1 U35090 ( .A1(n2754), .A2(n2753), .ZN(n2755) );
  AND2_X1 U35100 ( .A1(n2777), .A2(n2755), .ZN(n4615) );
  NAND2_X1 U35110 ( .A1(n4615), .A2(n2898), .ZN(n2760) );
  INV_X1 U35120 ( .A(REG2_REG_17__SCAN_IN), .ZN(n3322) );
  NAND2_X1 U35130 ( .A1(n2525), .A2(REG0_REG_17__SCAN_IN), .ZN(n2757) );
  INV_X1 U35140 ( .A(REG1_REG_17__SCAN_IN), .ZN(n4724) );
  OR2_X1 U35150 ( .A1(n2509), .A2(n4724), .ZN(n2756) );
  OAI211_X1 U35160 ( .C1(n3322), .C2(n3465), .A(n2757), .B(n2756), .ZN(n2758)
         );
  INV_X1 U35170 ( .A(n2758), .ZN(n2759) );
  NAND2_X1 U35180 ( .A1(n4624), .A2(n2549), .ZN(n2768) );
  NOR2_X1 U35190 ( .A1(n2761), .A2(n2763), .ZN(n2762) );
  MUX2_X1 U35200 ( .A(n2763), .B(n2762), .S(IR_REG_17__SCAN_IN), .Z(n2766) );
  NOR2_X1 U35210 ( .A1(n2766), .A2(n2765), .ZN(n4368) );
  MUX2_X1 U35220 ( .A(n4368), .B(DATAI_17_), .S(n3085), .Z(n4011) );
  NAND2_X1 U35230 ( .A1(n2414), .A2(n4011), .ZN(n2767) );
  NAND2_X1 U35240 ( .A1(n2768), .A2(n2767), .ZN(n2769) );
  XNOR2_X1 U35250 ( .A(n2769), .B(n2914), .ZN(n4009) );
  NAND2_X1 U35260 ( .A1(n4624), .A2(n2504), .ZN(n2771) );
  NAND2_X1 U35270 ( .A1(n2138), .A2(n4011), .ZN(n2770) );
  NAND2_X1 U35280 ( .A1(n2771), .A2(n2770), .ZN(n4008) );
  NOR2_X1 U35290 ( .A1(n4009), .A2(n4008), .ZN(n2774) );
  INV_X1 U35300 ( .A(n4009), .ZN(n2773) );
  INV_X1 U35310 ( .A(n4008), .ZN(n2772) );
  OAI22_X2 U35320 ( .A1(n4007), .A2(n2774), .B1(n2773), .B2(n2772), .ZN(n4093)
         );
  INV_X1 U35330 ( .A(REG3_REG_18__SCAN_IN), .ZN(n2776) );
  NAND2_X1 U35340 ( .A1(n2777), .A2(n2776), .ZN(n2778) );
  NAND2_X1 U35350 ( .A1(n2793), .A2(n2778), .ZN(n4597) );
  NAND2_X1 U35360 ( .A1(n2494), .A2(REG2_REG_18__SCAN_IN), .ZN(n2780) );
  INV_X1 U35370 ( .A(REG0_REG_18__SCAN_IN), .ZN(n3172) );
  OR2_X1 U35380 ( .A1(n2601), .A2(n3172), .ZN(n2779) );
  OAI211_X1 U35390 ( .C1(n2509), .C2(n4364), .A(n2780), .B(n2779), .ZN(n2781)
         );
  INV_X1 U35400 ( .A(n2781), .ZN(n2782) );
  NAND2_X1 U35410 ( .A1(n4608), .A2(n2549), .ZN(n2787) );
  NAND2_X1 U35420 ( .A1(n2764), .A2(IR_REG_31__SCAN_IN), .ZN(n2784) );
  XNOR2_X1 U35430 ( .A(n2784), .B(IR_REG_18__SCAN_IN), .ZN(n4367) );
  INV_X1 U35440 ( .A(n4367), .ZN(n4926) );
  INV_X1 U35450 ( .A(DATAI_18_), .ZN(n2785) );
  MUX2_X1 U35460 ( .A(n4926), .B(n2785), .S(n3085), .Z(n4595) );
  OR2_X1 U35470 ( .A1(n2916), .A2(n4595), .ZN(n2786) );
  NAND2_X1 U35480 ( .A1(n2787), .A2(n2786), .ZN(n2788) );
  XNOR2_X1 U35490 ( .A(n2788), .B(n2849), .ZN(n2791) );
  NOR2_X1 U35500 ( .A1(n2135), .A2(n4595), .ZN(n2789) );
  AOI21_X1 U35510 ( .B1(n4608), .B2(n2504), .A(n2789), .ZN(n2790) );
  NOR2_X1 U35520 ( .A1(n2791), .A2(n2790), .ZN(n4089) );
  NAND2_X1 U35530 ( .A1(n2791), .A2(n2790), .ZN(n4090) );
  NAND2_X1 U35540 ( .A1(n2793), .A2(n2222), .ZN(n2794) );
  NAND2_X1 U35550 ( .A1(n2806), .A2(n2794), .ZN(n4029) );
  INV_X1 U35560 ( .A(REG1_REG_19__SCAN_IN), .ZN(n4716) );
  NAND2_X1 U35570 ( .A1(n2525), .A2(REG0_REG_19__SCAN_IN), .ZN(n2796) );
  NAND2_X1 U35580 ( .A1(n2494), .A2(REG2_REG_19__SCAN_IN), .ZN(n2795) );
  OAI211_X1 U35590 ( .C1(n3462), .C2(n4716), .A(n2796), .B(n2795), .ZN(n2797)
         );
  INV_X1 U35600 ( .A(n2797), .ZN(n2798) );
  INV_X1 U35610 ( .A(DATAI_19_), .ZN(n2800) );
  MUX2_X1 U35620 ( .A(n4376), .B(n2800), .S(n3085), .Z(n4579) );
  OAI22_X1 U35630 ( .A1(n4591), .A2(n2913), .B1(n4579), .B2(n2135), .ZN(n2803)
         );
  OAI22_X1 U35640 ( .A1(n4591), .A2(n2136), .B1(n4579), .B2(n2916), .ZN(n2801)
         );
  XNOR2_X1 U35650 ( .A(n2801), .B(n2914), .ZN(n2802) );
  XOR2_X1 U35660 ( .A(n2803), .B(n2802), .Z(n4028) );
  INV_X1 U35670 ( .A(n2802), .ZN(n2805) );
  INV_X1 U35680 ( .A(n2803), .ZN(n2804) );
  INV_X1 U35690 ( .A(REG3_REG_20__SCAN_IN), .ZN(n4073) );
  NAND2_X1 U35700 ( .A1(n2806), .A2(n4073), .ZN(n2807) );
  NAND2_X1 U35710 ( .A1(n2819), .A2(n2807), .ZN(n4072) );
  INV_X1 U35720 ( .A(REG0_REG_20__SCAN_IN), .ZN(n4776) );
  NAND2_X1 U35730 ( .A1(n2494), .A2(REG2_REG_20__SCAN_IN), .ZN(n2809) );
  NAND2_X1 U35740 ( .A1(n2972), .A2(REG1_REG_20__SCAN_IN), .ZN(n2808) );
  OAI211_X1 U35750 ( .C1(n2601), .C2(n4776), .A(n2809), .B(n2808), .ZN(n2810)
         );
  INV_X1 U35760 ( .A(n2810), .ZN(n2811) );
  NAND2_X1 U35770 ( .A1(n4574), .A2(n2138), .ZN(n2814) );
  AND2_X1 U35780 ( .A1(n3085), .A2(DATAI_20_), .ZN(n3071) );
  OR2_X1 U35790 ( .A1(n2916), .A2(n4558), .ZN(n2813) );
  NAND2_X1 U35800 ( .A1(n2814), .A2(n2813), .ZN(n2815) );
  XNOR2_X1 U35810 ( .A(n2815), .B(n2849), .ZN(n2818) );
  NOR2_X1 U3582 ( .A1(n2136), .A2(n4558), .ZN(n2816) );
  AOI21_X1 U3583 ( .B1(n4574), .B2(n2504), .A(n2816), .ZN(n2817) );
  NOR2_X1 U3584 ( .A1(n2818), .A2(n2817), .ZN(n4070) );
  AND2_X1 U3585 ( .A1(n2818), .A2(n2817), .ZN(n4069) );
  INV_X1 U3586 ( .A(REG3_REG_21__SCAN_IN), .ZN(n3255) );
  NAND2_X1 U3587 ( .A1(n2819), .A2(n3255), .ZN(n2820) );
  NAND2_X1 U3588 ( .A1(n4538), .A2(n2898), .ZN(n2825) );
  INV_X1 U3589 ( .A(REG1_REG_21__SCAN_IN), .ZN(n4708) );
  NAND2_X1 U3590 ( .A1(n2525), .A2(REG0_REG_21__SCAN_IN), .ZN(n2822) );
  NAND2_X1 U3591 ( .A1(n2494), .A2(REG2_REG_21__SCAN_IN), .ZN(n2821) );
  OAI211_X1 U3592 ( .C1(n2509), .C2(n4708), .A(n2822), .B(n2821), .ZN(n2823)
         );
  INV_X1 U3593 ( .A(n2823), .ZN(n2824) );
  NAND2_X1 U3594 ( .A1(n4553), .A2(n2138), .ZN(n2827) );
  OR2_X1 U3595 ( .A1(n2916), .A2(n4536), .ZN(n2826) );
  NAND2_X1 U3596 ( .A1(n2827), .A2(n2826), .ZN(n2828) );
  XNOR2_X1 U3597 ( .A(n2828), .B(n2849), .ZN(n4038) );
  NOR2_X1 U3598 ( .A1(n2135), .A2(n4536), .ZN(n2829) );
  AOI21_X1 U3599 ( .B1(n4553), .B2(n2504), .A(n2829), .ZN(n2830) );
  NAND2_X1 U3600 ( .A1(n4038), .A2(n2830), .ZN(n2832) );
  INV_X1 U3601 ( .A(n4038), .ZN(n2831) );
  INV_X1 U3602 ( .A(n2830), .ZN(n4037) );
  XNOR2_X1 U3603 ( .A(n2842), .B(REG3_REG_22__SCAN_IN), .ZN(n4520) );
  NAND2_X1 U3604 ( .A1(n4520), .A2(n2898), .ZN(n2837) );
  INV_X1 U3605 ( .A(REG1_REG_22__SCAN_IN), .ZN(n3176) );
  NAND2_X1 U3606 ( .A1(n2494), .A2(REG2_REG_22__SCAN_IN), .ZN(n2834) );
  INV_X1 U3607 ( .A(REG0_REG_22__SCAN_IN), .ZN(n3174) );
  OR2_X1 U3608 ( .A1(n2601), .A2(n3174), .ZN(n2833) );
  OAI211_X1 U3609 ( .C1(n2509), .C2(n3176), .A(n2834), .B(n2833), .ZN(n2835)
         );
  INV_X1 U3610 ( .A(n2835), .ZN(n2836) );
  AND2_X1 U3611 ( .A1(n3085), .A2(DATAI_22_), .ZN(n4521) );
  OAI22_X1 U3612 ( .A1(n4043), .A2(n2913), .B1(n4514), .B2(n2135), .ZN(n2851)
         );
  OAI22_X1 U3613 ( .A1(n4043), .A2(n2136), .B1(n4514), .B2(n2916), .ZN(n2838)
         );
  XNOR2_X1 U3614 ( .A(n2838), .B(n2914), .ZN(n2852) );
  XOR2_X1 U3615 ( .A(n2851), .B(n2852), .Z(n4079) );
  NAND2_X1 U3616 ( .A1(n4078), .A2(n4079), .ZN(n3096) );
  AND2_X1 U3617 ( .A1(REG3_REG_23__SCAN_IN), .A2(REG3_REG_22__SCAN_IN), .ZN(
        n2839) );
  INV_X1 U3618 ( .A(REG3_REG_22__SCAN_IN), .ZN(n4081) );
  INV_X1 U3619 ( .A(REG3_REG_23__SCAN_IN), .ZN(n2841) );
  OAI21_X1 U3620 ( .B1(n2842), .B2(n4081), .A(n2841), .ZN(n2843) );
  NAND2_X1 U3621 ( .A1(n2855), .A2(n2843), .ZN(n4504) );
  INV_X1 U3622 ( .A(REG1_REG_23__SCAN_IN), .ZN(n4700) );
  NAND2_X1 U3623 ( .A1(n2494), .A2(REG2_REG_23__SCAN_IN), .ZN(n2845) );
  NAND2_X1 U3624 ( .A1(n2525), .A2(REG0_REG_23__SCAN_IN), .ZN(n2844) );
  OAI211_X1 U3625 ( .C1(n3462), .C2(n4700), .A(n2845), .B(n2844), .ZN(n2846)
         );
  INV_X1 U3626 ( .A(n2846), .ZN(n2847) );
  NAND2_X1 U3627 ( .A1(n2571), .A2(DATAI_23_), .ZN(n4503) );
  OAI22_X1 U3628 ( .A1(n4517), .A2(n2135), .B1(n4503), .B2(n2916), .ZN(n2850)
         );
  XNOR2_X1 U3629 ( .A(n2850), .B(n2849), .ZN(n2863) );
  OAI22_X1 U3630 ( .A1(n4517), .A2(n2913), .B1(n4503), .B2(n2136), .ZN(n2864)
         );
  XNOR2_X1 U3631 ( .A(n2863), .B(n2864), .ZN(n3097) );
  OR2_X1 U3632 ( .A1(n2852), .A2(n2851), .ZN(n3098) );
  INV_X1 U3633 ( .A(REG3_REG_24__SCAN_IN), .ZN(n4062) );
  NAND2_X1 U3634 ( .A1(n2855), .A2(n4062), .ZN(n2856) );
  NAND2_X1 U3635 ( .A1(n2869), .A2(n2856), .ZN(n4487) );
  INV_X1 U3636 ( .A(REG1_REG_24__SCAN_IN), .ZN(n4696) );
  NAND2_X1 U3637 ( .A1(n2525), .A2(REG0_REG_24__SCAN_IN), .ZN(n2858) );
  NAND2_X1 U3638 ( .A1(n2494), .A2(REG2_REG_24__SCAN_IN), .ZN(n2857) );
  OAI211_X1 U3639 ( .C1(n3462), .C2(n4696), .A(n2858), .B(n2857), .ZN(n2859)
         );
  INV_X1 U3640 ( .A(n2859), .ZN(n2860) );
  AND2_X1 U3641 ( .A1(n3085), .A2(DATAI_24_), .ZN(n4065) );
  NOR2_X1 U3642 ( .A1(n2135), .A2(n4484), .ZN(n2862) );
  AOI21_X1 U3643 ( .B1(n4457), .B2(n2504), .A(n2862), .ZN(n2867) );
  INV_X1 U3644 ( .A(n2863), .ZN(n2865) );
  NAND2_X1 U3645 ( .A1(n2865), .A2(n2864), .ZN(n2868) );
  OAI22_X1 U3646 ( .A1(n4497), .A2(n2136), .B1(n4484), .B2(n2916), .ZN(n2866)
         );
  XNOR2_X1 U3647 ( .A(n2866), .B(n2914), .ZN(n4059) );
  INV_X1 U3648 ( .A(REG3_REG_25__SCAN_IN), .ZN(n4050) );
  NAND2_X1 U3649 ( .A1(n2869), .A2(n4050), .ZN(n2870) );
  NAND2_X1 U3650 ( .A1(n4465), .A2(n2898), .ZN(n2875) );
  INV_X1 U3651 ( .A(REG1_REG_25__SCAN_IN), .ZN(n3183) );
  NAND2_X1 U3652 ( .A1(n2494), .A2(REG2_REG_25__SCAN_IN), .ZN(n2872) );
  NAND2_X1 U3653 ( .A1(n2525), .A2(REG0_REG_25__SCAN_IN), .ZN(n2871) );
  OAI211_X1 U3654 ( .C1(n3462), .C2(n3183), .A(n2872), .B(n2871), .ZN(n2873)
         );
  INV_X1 U3655 ( .A(n2873), .ZN(n2874) );
  NAND2_X1 U3656 ( .A1(n4479), .A2(n2549), .ZN(n2877) );
  AND2_X1 U3657 ( .A1(n3085), .A2(DATAI_25_), .ZN(n4456) );
  INV_X1 U3658 ( .A(n4456), .ZN(n4463) );
  OR2_X1 U3659 ( .A1(n2916), .A2(n4463), .ZN(n2876) );
  NAND2_X1 U3660 ( .A1(n2877), .A2(n2876), .ZN(n2878) );
  XNOR2_X1 U3661 ( .A(n2878), .B(n2914), .ZN(n2882) );
  NAND2_X1 U3662 ( .A1(n4479), .A2(n2504), .ZN(n2880) );
  NAND2_X1 U3663 ( .A1(n2138), .A2(n4456), .ZN(n2879) );
  NAND2_X1 U3664 ( .A1(n2880), .A2(n2879), .ZN(n2881) );
  NAND2_X1 U3665 ( .A1(n2882), .A2(n2881), .ZN(n4048) );
  NAND2_X1 U3666 ( .A1(n2883), .A2(n2214), .ZN(n2884) );
  NAND2_X1 U3667 ( .A1(n2896), .A2(n2884), .ZN(n4448) );
  INV_X1 U3668 ( .A(REG1_REG_26__SCAN_IN), .ZN(n4688) );
  NAND2_X1 U3669 ( .A1(n2525), .A2(REG0_REG_26__SCAN_IN), .ZN(n2886) );
  NAND2_X1 U3670 ( .A1(n2494), .A2(REG2_REG_26__SCAN_IN), .ZN(n2885) );
  OAI211_X1 U3671 ( .C1(n3462), .C2(n4688), .A(n2886), .B(n2885), .ZN(n2887)
         );
  INV_X1 U3672 ( .A(n2887), .ZN(n2888) );
  NAND2_X1 U3673 ( .A1(n3085), .A2(DATAI_26_), .ZN(n4440) );
  OAI22_X1 U3674 ( .A1(n4459), .A2(n2136), .B1(n4440), .B2(n2916), .ZN(n2890)
         );
  XNOR2_X1 U3675 ( .A(n2890), .B(n2914), .ZN(n2891) );
  OAI22_X1 U3676 ( .A1(n4459), .A2(n2913), .B1(n4440), .B2(n2136), .ZN(n2892)
         );
  AND2_X1 U3677 ( .A1(n2891), .A2(n2892), .ZN(n4102) );
  INV_X1 U3678 ( .A(n2891), .ZN(n2894) );
  INV_X1 U3679 ( .A(n2892), .ZN(n2893) );
  NAND2_X1 U3680 ( .A1(n2894), .A2(n2893), .ZN(n4101) );
  INV_X1 U3681 ( .A(REG3_REG_27__SCAN_IN), .ZN(n2895) );
  NAND2_X1 U3682 ( .A1(n2896), .A2(n2895), .ZN(n2897) );
  NAND2_X1 U3683 ( .A1(n4421), .A2(n2898), .ZN(n2903) );
  INV_X1 U3684 ( .A(REG2_REG_27__SCAN_IN), .ZN(n4422) );
  NAND2_X1 U3685 ( .A1(n2525), .A2(REG0_REG_27__SCAN_IN), .ZN(n2900) );
  INV_X1 U3686 ( .A(REG1_REG_27__SCAN_IN), .ZN(n3185) );
  OR2_X1 U3687 ( .A1(n2509), .A2(n3185), .ZN(n2899) );
  OAI211_X1 U3688 ( .C1(n4422), .C2(n3465), .A(n2900), .B(n2899), .ZN(n2901)
         );
  INV_X1 U3689 ( .A(n2901), .ZN(n2902) );
  AND2_X1 U3690 ( .A1(n2571), .A2(DATAI_27_), .ZN(n4420) );
  OAI22_X1 U3691 ( .A1(n4268), .A2(n2136), .B1(n4428), .B2(n2916), .ZN(n2904)
         );
  XNOR2_X1 U3692 ( .A(n2904), .B(n2914), .ZN(n2919) );
  OAI22_X1 U3693 ( .A1(n4268), .A2(n2913), .B1(n4428), .B2(n2135), .ZN(n2920)
         );
  INV_X1 U3694 ( .A(n2907), .ZN(n2905) );
  INV_X1 U3695 ( .A(REG3_REG_28__SCAN_IN), .ZN(n2906) );
  NAND2_X1 U3696 ( .A1(n2907), .A2(n2906), .ZN(n2908) );
  INV_X1 U3697 ( .A(REG1_REG_28__SCAN_IN), .ZN(n3189) );
  NAND2_X1 U3698 ( .A1(n2494), .A2(REG2_REG_28__SCAN_IN), .ZN(n2910) );
  INV_X1 U3699 ( .A(REG0_REG_28__SCAN_IN), .ZN(n3188) );
  OR2_X1 U3700 ( .A1(n2601), .A2(n3188), .ZN(n2909) );
  OAI211_X1 U3701 ( .C1(n2509), .C2(n3189), .A(n2910), .B(n2909), .ZN(n2911)
         );
  INV_X1 U3702 ( .A(n2911), .ZN(n2912) );
  AND2_X1 U3703 ( .A1(n3085), .A2(DATAI_28_), .ZN(n4391) );
  INV_X1 U3704 ( .A(n4391), .ZN(n3075) );
  OAI22_X1 U3705 ( .A1(n3032), .A2(n2913), .B1(n3075), .B2(n2135), .ZN(n2915)
         );
  XNOR2_X1 U3706 ( .A(n2915), .B(n2914), .ZN(n2918) );
  OAI22_X1 U3707 ( .A1(n3032), .A2(n2135), .B1(n3075), .B2(n2916), .ZN(n2917)
         );
  XNOR2_X1 U3708 ( .A(n2918), .B(n2917), .ZN(n2955) );
  INV_X1 U3709 ( .A(n2919), .ZN(n2922) );
  INV_X1 U3710 ( .A(n2920), .ZN(n2921) );
  INV_X1 U3711 ( .A(IR_REG_23__SCAN_IN), .ZN(n2945) );
  NAND2_X1 U3712 ( .A1(n2944), .A2(IR_REG_31__SCAN_IN), .ZN(n2925) );
  INV_X1 U3713 ( .A(n3373), .ZN(n4806) );
  INV_X1 U3714 ( .A(B_REG_SCAN_IN), .ZN(n3312) );
  NAND2_X1 U3715 ( .A1(n4806), .A2(n3312), .ZN(n2929) );
  OR2_X1 U3716 ( .A1(n2927), .A2(n2926), .ZN(n3367) );
  NAND3_X1 U3717 ( .A1(n3373), .A2(B_REG_SCAN_IN), .A3(n3367), .ZN(n2928) );
  NAND3_X1 U3718 ( .A1(n2929), .A2(n2928), .A3(n4805), .ZN(n3371) );
  OR2_X1 U3719 ( .A1(n3371), .A2(D_REG_0__SCAN_IN), .ZN(n2931) );
  INV_X1 U3720 ( .A(n4805), .ZN(n3372) );
  NAND2_X1 U3721 ( .A1(n3373), .A2(n3372), .ZN(n2930) );
  NOR4_X1 U3722 ( .A1(D_REG_8__SCAN_IN), .A2(D_REG_26__SCAN_IN), .A3(
        D_REG_16__SCAN_IN), .A4(D_REG_23__SCAN_IN), .ZN(n3121) );
  NOR2_X1 U3723 ( .A1(D_REG_30__SCAN_IN), .A2(D_REG_31__SCAN_IN), .ZN(n2934)
         );
  NOR4_X1 U3724 ( .A1(D_REG_5__SCAN_IN), .A2(D_REG_18__SCAN_IN), .A3(
        D_REG_6__SCAN_IN), .A4(D_REG_24__SCAN_IN), .ZN(n2933) );
  NOR4_X1 U3725 ( .A1(D_REG_11__SCAN_IN), .A2(D_REG_12__SCAN_IN), .A3(
        D_REG_2__SCAN_IN), .A4(D_REG_21__SCAN_IN), .ZN(n2932) );
  NAND4_X1 U3726 ( .A1(n3121), .A2(n2934), .A3(n2933), .A4(n2932), .ZN(n2940)
         );
  NOR4_X1 U3727 ( .A1(D_REG_7__SCAN_IN), .A2(D_REG_9__SCAN_IN), .A3(
        D_REG_13__SCAN_IN), .A4(D_REG_14__SCAN_IN), .ZN(n2938) );
  NOR4_X1 U3728 ( .A1(D_REG_29__SCAN_IN), .A2(D_REG_3__SCAN_IN), .A3(
        D_REG_4__SCAN_IN), .A4(D_REG_10__SCAN_IN), .ZN(n2937) );
  NOR4_X1 U3729 ( .A1(D_REG_20__SCAN_IN), .A2(D_REG_28__SCAN_IN), .A3(
        D_REG_25__SCAN_IN), .A4(D_REG_27__SCAN_IN), .ZN(n2936) );
  NOR4_X1 U3730 ( .A1(D_REG_15__SCAN_IN), .A2(D_REG_17__SCAN_IN), .A3(
        D_REG_22__SCAN_IN), .A4(D_REG_19__SCAN_IN), .ZN(n2935) );
  NAND4_X1 U3731 ( .A1(n2938), .A2(n2937), .A3(n2936), .A4(n2935), .ZN(n2939)
         );
  NOR2_X1 U3732 ( .A1(n2940), .A2(n2939), .ZN(n3064) );
  AND2_X1 U3733 ( .A1(n3064), .A2(D_REG_1__SCAN_IN), .ZN(n2941) );
  OR2_X1 U3734 ( .A1(n3371), .A2(n2941), .ZN(n2942) );
  NAND2_X1 U3735 ( .A1(n3372), .A2(n3367), .ZN(n3376) );
  NAND2_X1 U3736 ( .A1(n2942), .A2(n3376), .ZN(n3495) );
  INV_X1 U3737 ( .A(n3495), .ZN(n2943) );
  INV_X1 U3738 ( .A(n3382), .ZN(n2951) );
  NAND2_X1 U3739 ( .A1(n2137), .A2(n4376), .ZN(n2959) );
  INV_X1 U3740 ( .A(n2959), .ZN(n2949) );
  OR2_X1 U3741 ( .A1(n2948), .A2(n2949), .ZN(n2950) );
  NAND2_X1 U3742 ( .A1(n2951), .A2(n2950), .ZN(n2957) );
  NOR2_X1 U3743 ( .A1(n3531), .A2(n2957), .ZN(n2952) );
  NOR3_X1 U3744 ( .A1(n2954), .A2(n4109), .A3(n2403), .ZN(n2956) );
  NAND2_X1 U3745 ( .A1(n2957), .A2(n4627), .ZN(n2958) );
  NAND2_X1 U3746 ( .A1(n2980), .A2(n2958), .ZN(n2961) );
  AND2_X1 U3747 ( .A1(n3382), .A2(n2959), .ZN(n3062) );
  INV_X1 U3748 ( .A(n3062), .ZN(n2960) );
  NAND2_X1 U3749 ( .A1(n2961), .A2(n2960), .ZN(n3532) );
  NAND2_X1 U3750 ( .A1(n2962), .A2(n3381), .ZN(n2963) );
  OAI21_X1 U3751 ( .B1(n3532), .B2(n2963), .A(STATE_REG_SCAN_IN), .ZN(n2966)
         );
  INV_X1 U3752 ( .A(n2964), .ZN(n2965) );
  AND3_X1 U3753 ( .A1(n2138), .A2(n4924), .A3(n2965), .ZN(n4279) );
  NAND2_X1 U3754 ( .A1(n2980), .A2(n4279), .ZN(n3530) );
  OR3_X1 U3755 ( .A1(n2967), .A2(IR_REG_27__SCAN_IN), .A3(IR_REG_26__SCAN_IN), 
        .ZN(n2968) );
  NAND2_X1 U3756 ( .A1(n2968), .A2(IR_REG_31__SCAN_IN), .ZN(n2970) );
  XNOR2_X1 U3757 ( .A(n2970), .B(n2969), .ZN(n4819) );
  NAND2_X1 U3758 ( .A1(n4279), .A2(n4819), .ZN(n2971) );
  NOR2_X2 U3759 ( .A1(n2980), .A2(n2971), .ZN(n4117) );
  INV_X1 U3760 ( .A(REG2_REG_29__SCAN_IN), .ZN(n2975) );
  NAND2_X1 U3761 ( .A1(n2525), .A2(REG0_REG_29__SCAN_IN), .ZN(n2974) );
  NAND2_X1 U3762 ( .A1(n2972), .A2(REG1_REG_29__SCAN_IN), .ZN(n2973) );
  OAI211_X1 U3763 ( .C1(n2975), .C2(n3465), .A(n2974), .B(n2973), .ZN(n2976)
         );
  INV_X1 U3764 ( .A(n2976), .ZN(n2977) );
  INV_X1 U3765 ( .A(n4819), .ZN(n4307) );
  NAND2_X1 U3766 ( .A1(n4279), .A2(n4307), .ZN(n2979) );
  NOR2_X2 U3767 ( .A1(n2980), .A2(n2979), .ZN(n4118) );
  AOI22_X1 U3768 ( .A1(n4117), .A2(n4284), .B1(n4443), .B2(n4118), .ZN(n2985)
         );
  NOR2_X1 U3769 ( .A1(n3531), .A2(n4627), .ZN(n2981) );
  NAND2_X1 U3770 ( .A1(n2982), .A2(n2981), .ZN(n2983) );
  INV_X1 U3771 ( .A(n4376), .ZN(n4808) );
  NAND2_X1 U3772 ( .A1(n2137), .A2(n4808), .ZN(n4902) );
  NAND2_X1 U3773 ( .A1(n2983), .A2(n4647), .ZN(n4119) );
  AOI22_X1 U3774 ( .A1(n4119), .A2(n4391), .B1(REG3_REG_28__SCAN_IN), .B2(
        U3149), .ZN(n2984) );
  OAI211_X1 U3775 ( .C1(n4122), .C2(n4413), .A(n2985), .B(n2984), .ZN(n2986)
         );
  INV_X1 U3776 ( .A(n3643), .ZN(n2988) );
  NAND2_X1 U3777 ( .A1(n2988), .A2(n2499), .ZN(n3037) );
  NAND2_X1 U3778 ( .A1(n3643), .A2(n2992), .ZN(n4212) );
  NAND2_X1 U3779 ( .A1(n3037), .A2(n4212), .ZN(n4172) );
  NAND2_X1 U3780 ( .A1(n3639), .A2(n3638), .ZN(n3637) );
  NAND2_X1 U3781 ( .A1(n2990), .A2(n2472), .ZN(n3667) );
  NAND3_X1 U3782 ( .A1(n4172), .A2(n3637), .A3(n3667), .ZN(n3670) );
  OR2_X1 U3783 ( .A1(n3643), .A2(n2499), .ZN(n2993) );
  NAND2_X1 U3784 ( .A1(n3670), .A2(n2993), .ZN(n3579) );
  NAND2_X1 U3785 ( .A1(n3504), .A2(n3590), .ZN(n2995) );
  NOR2_X1 U3786 ( .A1(n3504), .A2(n3590), .ZN(n2994) );
  OR2_X1 U3787 ( .A1(n3620), .A2(n3609), .ZN(n4215) );
  NAND2_X1 U3788 ( .A1(n3620), .A2(n3609), .ZN(n4219) );
  NAND2_X1 U3789 ( .A1(n4215), .A2(n4219), .ZN(n3503) );
  NAND2_X1 U3790 ( .A1(n3491), .A2(n3503), .ZN(n3493) );
  INV_X1 U3791 ( .A(n3609), .ZN(n3505) );
  NAND2_X1 U3792 ( .A1(n3620), .A2(n3505), .ZN(n2996) );
  NAND2_X1 U3793 ( .A1(n3493), .A2(n2996), .ZN(n3595) );
  OR2_X1 U3794 ( .A1(n3830), .A2(n2998), .ZN(n2997) );
  NAND2_X1 U3795 ( .A1(n3595), .A2(n2997), .ZN(n3711) );
  NAND2_X1 U3796 ( .A1(n3830), .A2(n2998), .ZN(n3710) );
  NAND2_X1 U3797 ( .A1(n3796), .A2(n3734), .ZN(n3000) );
  OAI21_X1 U3798 ( .B1(n3831), .B2(n4291), .A(n3716), .ZN(n3722) );
  NAND2_X1 U3799 ( .A1(n3002), .A2(n3722), .ZN(n3004) );
  OR2_X1 U3800 ( .A1(n3796), .A2(n3734), .ZN(n3003) );
  INV_X1 U3801 ( .A(n3808), .ZN(n3014) );
  NOR2_X1 U3802 ( .A1(n4289), .A2(n3817), .ZN(n3841) );
  AND2_X1 U3803 ( .A1(n3918), .A2(n3757), .ZN(n3007) );
  OR2_X1 U3804 ( .A1(n3841), .A2(n3007), .ZN(n3924) );
  OR2_X1 U3805 ( .A1(n3924), .A2(n3009), .ZN(n3964) );
  NOR2_X1 U3806 ( .A1(n3983), .A2(n3043), .ZN(n3012) );
  NAND2_X1 U3807 ( .A1(n4288), .A2(n3757), .ZN(n4239) );
  NAND2_X1 U3808 ( .A1(n4289), .A2(n3817), .ZN(n3842) );
  NAND2_X1 U3809 ( .A1(n4287), .A2(n3921), .ZN(n3008) );
  NAND2_X1 U3810 ( .A1(n3925), .A2(n3008), .ZN(n3011) );
  NOR2_X1 U3811 ( .A1(n3965), .A2(n3012), .ZN(n3013) );
  AOI21_X1 U3812 ( .B1(n3014), .B2(n2139), .A(n2152), .ZN(n3987) );
  NAND2_X1 U3813 ( .A1(n4651), .A2(n3990), .ZN(n4126) );
  INV_X1 U3814 ( .A(n4651), .ZN(n4286) );
  NAND2_X1 U3815 ( .A1(n4286), .A2(n3986), .ZN(n4230) );
  NAND2_X1 U3816 ( .A1(n3987), .A2(n3015), .ZN(n3988) );
  NAND2_X1 U3817 ( .A1(n4651), .A2(n3986), .ZN(n3016) );
  NAND2_X1 U3818 ( .A1(n3988), .A2(n3016), .ZN(n4644) );
  NAND2_X1 U3819 ( .A1(n4621), .A2(n4660), .ZN(n3017) );
  OR2_X1 U3820 ( .A1(n4621), .A2(n4660), .ZN(n3018) );
  INV_X1 U3821 ( .A(n4633), .ZN(n4001) );
  NAND2_X1 U3822 ( .A1(n4652), .A2(n4001), .ZN(n4253) );
  NAND2_X1 U3823 ( .A1(n4116), .A2(n4633), .ZN(n4545) );
  NAND2_X1 U3824 ( .A1(n4116), .A2(n4001), .ZN(n3019) );
  NAND2_X2 U3825 ( .A1(n4630), .A2(n3019), .ZN(n4612) );
  OR2_X1 U3826 ( .A1(n4624), .A2(n4011), .ZN(n3020) );
  OR2_X1 U3827 ( .A1(n4608), .A2(n4595), .ZN(n4568) );
  NAND2_X1 U3828 ( .A1(n4608), .A2(n4595), .ZN(n4569) );
  NAND2_X1 U3829 ( .A1(n4568), .A2(n4569), .ZN(n4601) );
  INV_X1 U3830 ( .A(n4608), .ZN(n4572) );
  INV_X1 U3831 ( .A(n4579), .ZN(n4030) );
  NOR2_X1 U3832 ( .A1(n4574), .A2(n3071), .ZN(n3021) );
  INV_X1 U3833 ( .A(n4574), .ZN(n4032) );
  NAND2_X1 U3834 ( .A1(n4043), .A2(n4521), .ZN(n4493) );
  NAND2_X1 U3835 ( .A1(n4532), .A2(n4514), .ZN(n3054) );
  NAND2_X1 U3836 ( .A1(n4493), .A2(n3054), .ZN(n4511) );
  NAND2_X1 U3837 ( .A1(n4517), .A2(n4503), .ZN(n3024) );
  NOR2_X1 U3838 ( .A1(n4517), .A2(n4503), .ZN(n3023) );
  AOI21_X1 U3839 ( .B1(n4492), .B2(n3024), .A(n3023), .ZN(n4470) );
  NAND2_X1 U3840 ( .A1(n4457), .A2(n4065), .ZN(n3025) );
  NAND2_X1 U3841 ( .A1(n4470), .A2(n3025), .ZN(n3027) );
  NAND2_X1 U3842 ( .A1(n4497), .A2(n4484), .ZN(n3026) );
  NAND2_X1 U3843 ( .A1(n3027), .A2(n3026), .ZN(n4453) );
  NOR2_X1 U3844 ( .A1(n4479), .A2(n4456), .ZN(n3028) );
  NOR2_X1 U3845 ( .A1(n4459), .A2(n4440), .ZN(n3030) );
  NAND2_X1 U3846 ( .A1(n4459), .A2(n4440), .ZN(n3029) );
  NOR2_X1 U3847 ( .A1(n4443), .A2(n4420), .ZN(n3031) );
  NAND2_X1 U3848 ( .A1(n3032), .A2(n4391), .ZN(n4396) );
  NAND2_X1 U3849 ( .A1(n4430), .A2(n3075), .ZN(n4395) );
  XNOR2_X1 U3850 ( .A(n2468), .B(n3033), .ZN(n3034) );
  NAND2_X1 U3851 ( .A1(n3034), .A2(n4376), .ZN(n3650) );
  NAND2_X1 U3852 ( .A1(n3650), .A2(n4937), .ZN(n4744) );
  NAND2_X1 U3853 ( .A1(n3641), .A2(n4209), .ZN(n3036) );
  INV_X1 U3854 ( .A(n4172), .ZN(n3668) );
  NAND2_X1 U3855 ( .A1(n3036), .A2(n3668), .ZN(n3672) );
  NAND2_X1 U3856 ( .A1(n3672), .A2(n3037), .ZN(n3581) );
  NAND2_X1 U3857 ( .A1(n3504), .A2(n3617), .ZN(n4211) );
  INV_X1 U3858 ( .A(n4171), .ZN(n3582) );
  NAND2_X1 U3859 ( .A1(n3581), .A2(n3582), .ZN(n3580) );
  NAND2_X1 U3860 ( .A1(n3580), .A2(n4214), .ZN(n3502) );
  INV_X1 U3861 ( .A(n4215), .ZN(n3038) );
  OR2_X1 U3862 ( .A1(n3830), .A2(n3602), .ZN(n4232) );
  NAND2_X1 U3863 ( .A1(n3830), .A2(n3602), .ZN(n4217) );
  AND2_X1 U3864 ( .A1(n4291), .A2(n3069), .ZN(n4233) );
  OR2_X1 U3865 ( .A1(n4291), .A2(n3069), .ZN(n4221) );
  INV_X1 U3866 ( .A(n3039), .ZN(n3040) );
  NAND2_X1 U3867 ( .A1(n3727), .A2(n4226), .ZN(n3041) );
  NAND2_X1 U3868 ( .A1(n3796), .A2(n3070), .ZN(n4224) );
  AND2_X1 U3869 ( .A1(n3811), .A2(n3801), .ZN(n4235) );
  NAND2_X1 U3870 ( .A1(n4289), .A2(n2237), .ZN(n4238) );
  NAND2_X1 U3871 ( .A1(n3840), .A2(n4239), .ZN(n3042) );
  NAND2_X1 U3872 ( .A1(n4287), .A2(n3930), .ZN(n3960) );
  NAND2_X1 U3873 ( .A1(n3983), .A2(n3973), .ZN(n3044) );
  NOR2_X1 U3874 ( .A1(n4287), .A2(n3930), .ZN(n3961) );
  NOR2_X1 U3875 ( .A1(n3983), .A2(n3973), .ZN(n3045) );
  AOI21_X1 U3876 ( .B1(n4245), .B2(n3961), .A(n3045), .ZN(n4248) );
  NAND2_X1 U3877 ( .A1(n3046), .A2(n4126), .ZN(n4657) );
  INV_X1 U3878 ( .A(n4660), .ZN(n4645) );
  NAND2_X1 U3879 ( .A1(n4621), .A2(n4645), .ZN(n4229) );
  OR2_X1 U3880 ( .A1(n4621), .A2(n4645), .ZN(n4127) );
  NAND2_X1 U3881 ( .A1(n4229), .A2(n4127), .ZN(n4656) );
  AND2_X1 U3882 ( .A1(n4574), .A2(n4558), .ZN(n4252) );
  NAND2_X1 U3883 ( .A1(n3482), .A2(n4579), .ZN(n3047) );
  NAND2_X1 U3884 ( .A1(n3047), .A2(n4569), .ZN(n3050) );
  AND2_X1 U3885 ( .A1(n4624), .A2(n4613), .ZN(n4565) );
  NOR2_X1 U3886 ( .A1(n4252), .A2(n4546), .ZN(n3048) );
  AND2_X1 U3887 ( .A1(n3048), .A2(n4545), .ZN(n3052) );
  OR2_X1 U3888 ( .A1(n4624), .A2(n4613), .ZN(n4566) );
  AND2_X1 U3889 ( .A1(n4568), .A2(n4566), .ZN(n3049) );
  OAI22_X1 U3890 ( .A1(n3050), .A2(n3049), .B1(n4579), .B2(n3482), .ZN(n4547)
         );
  NOR2_X1 U3891 ( .A1(n4574), .A2(n4558), .ZN(n3051) );
  OR2_X1 U3892 ( .A1(n4547), .A2(n3051), .ZN(n4132) );
  INV_X1 U3893 ( .A(n4252), .ZN(n4131) );
  NAND2_X1 U3894 ( .A1(n4083), .A2(n4040), .ZN(n4257) );
  NAND2_X1 U3895 ( .A1(n4527), .A2(n4257), .ZN(n3053) );
  NAND2_X1 U3896 ( .A1(n4553), .A2(n4536), .ZN(n4255) );
  NAND2_X1 U3897 ( .A1(n3053), .A2(n4255), .ZN(n4471) );
  INV_X1 U3898 ( .A(n4517), .ZN(n3518) );
  NAND2_X1 U3899 ( .A1(n3518), .A2(n4503), .ZN(n4163) );
  NAND2_X1 U3900 ( .A1(n4497), .A2(n4065), .ZN(n4162) );
  INV_X1 U3901 ( .A(n4503), .ZN(n3073) );
  NAND2_X1 U3902 ( .A1(n4517), .A2(n3073), .ZN(n4473) );
  NAND2_X1 U3903 ( .A1(n4162), .A2(n4473), .ZN(n4259) );
  NOR2_X1 U3904 ( .A1(n4472), .A2(n4493), .ZN(n3055) );
  NOR2_X1 U3905 ( .A1(n4259), .A2(n3055), .ZN(n4136) );
  NAND2_X1 U3906 ( .A1(n4457), .A2(n4484), .ZN(n4161) );
  AND2_X1 U3907 ( .A1(n4479), .A2(n4463), .ZN(n4160) );
  INV_X1 U3908 ( .A(n4440), .ZN(n4446) );
  NAND2_X1 U3909 ( .A1(n4459), .A2(n4446), .ZN(n4158) );
  NAND2_X1 U3910 ( .A1(n4441), .A2(n4456), .ZN(n4436) );
  INV_X1 U3911 ( .A(n4459), .ZN(n4285) );
  AOI21_X1 U3912 ( .B1(n4437), .B2(n4263), .A(n4157), .ZN(n4425) );
  XNOR2_X1 U3913 ( .A(n4443), .B(n4420), .ZN(n4426) );
  NOR2_X1 U3914 ( .A1(n4443), .A2(n4428), .ZN(n4139) );
  XOR2_X1 U3915 ( .A(n4389), .B(n4398), .Z(n3061) );
  NAND2_X1 U3916 ( .A1(n2468), .A2(n4808), .ZN(n3057) );
  NAND2_X1 U3917 ( .A1(n4807), .A2(n2469), .ZN(n4276) );
  NOR2_X1 U3918 ( .A1(n4627), .A2(n3075), .ZN(n3058) );
  AOI21_X1 U3919 ( .B1(n4443), .B2(n4622), .A(n3058), .ZN(n3060) );
  NAND2_X1 U3920 ( .A1(n4284), .A2(n4623), .ZN(n3059) );
  OAI211_X1 U3921 ( .C1(n3061), .C2(n4655), .A(n3060), .B(n3059), .ZN(n4416)
         );
  AOI21_X1 U3922 ( .B1(n4410), .B2(n4744), .A(n4416), .ZN(n3084) );
  OAI21_X1 U3923 ( .B1(n3371), .B2(D_REG_1__SCAN_IN), .A(n3376), .ZN(n3067) );
  NOR2_X1 U3924 ( .A1(n4937), .A2(n2469), .ZN(n3063) );
  NOR2_X1 U3925 ( .A1(n3494), .A2(n3063), .ZN(n3066) );
  OR2_X1 U3926 ( .A1(n3371), .A2(n3064), .ZN(n3065) );
  AND2_X2 U3927 ( .A1(n3704), .A2(n3070), .ZN(n3802) );
  NAND2_X1 U3928 ( .A1(n3974), .A2(n3973), .ZN(n3972) );
  NOR2_X2 U3929 ( .A1(n3972), .A2(n3990), .ZN(n3989) );
  AND2_X2 U3930 ( .A1(n2406), .A2(n4633), .ZN(n4635) );
  INV_X1 U3931 ( .A(n4595), .ZN(n4589) );
  OR2_X2 U3932 ( .A1(n4557), .A2(n4040), .ZN(n4535) );
  NOR2_X2 U3933 ( .A1(n4535), .A2(n4521), .ZN(n3072) );
  INV_X1 U3934 ( .A(n3072), .ZN(n4501) );
  NAND2_X1 U3935 ( .A1(n4482), .A2(n4484), .ZN(n4462) );
  OAI21_X1 U3936 ( .B1(n3074), .B2(n3075), .A(n4394), .ZN(n4411) );
  OR2_X1 U3937 ( .A1(n4411), .A2(n4802), .ZN(n3078) );
  NAND2_X1 U3938 ( .A1(n4965), .A2(REG0_REG_28__SCAN_IN), .ZN(n3077) );
  OAI21_X1 U3939 ( .B1(n3084), .B2(n4965), .A(n2410), .ZN(U3514) );
  NAND2_X1 U3940 ( .A1(n4976), .A2(REG1_REG_28__SCAN_IN), .ZN(n3081) );
  INV_X1 U3941 ( .A(n3082), .ZN(n3083) );
  OAI21_X1 U3942 ( .B1(n3084), .B2(n4976), .A(n3083), .ZN(U3546) );
  NAND2_X1 U3943 ( .A1(n2571), .A2(DATAI_29_), .ZN(n4145) );
  INV_X1 U3944 ( .A(n4145), .ZN(n4399) );
  NAND2_X1 U3945 ( .A1(n2571), .A2(DATAI_30_), .ZN(n4385) );
  NAND2_X1 U3946 ( .A1(n3085), .A2(DATAI_31_), .ZN(n4164) );
  NAND2_X1 U3947 ( .A1(n4965), .A2(REG0_REG_31__SCAN_IN), .ZN(n3092) );
  OAI21_X1 U3948 ( .B1(n2967), .B2(IR_REG_26__SCAN_IN), .A(IR_REG_31__SCAN_IN), 
        .ZN(n3088) );
  XNOR2_X1 U3949 ( .A(n3088), .B(n3087), .ZN(n4305) );
  INV_X1 U3950 ( .A(n4305), .ZN(n4821) );
  AOI21_X1 U3951 ( .B1(B_REG_SCAN_IN), .B2(n4821), .A(n4901), .ZN(n4401) );
  INV_X1 U3952 ( .A(REG2_REG_31__SCAN_IN), .ZN(n3311) );
  NAND2_X1 U3953 ( .A1(n2525), .A2(REG0_REG_31__SCAN_IN), .ZN(n3090) );
  INV_X1 U3954 ( .A(REG1_REG_31__SCAN_IN), .ZN(n4667) );
  OR2_X1 U3955 ( .A1(n2509), .A2(n4667), .ZN(n3089) );
  OAI211_X1 U3956 ( .C1(n3465), .C2(n3311), .A(n3090), .B(n3089), .ZN(n4165)
         );
  NAND2_X1 U3957 ( .A1(n4401), .A2(n4165), .ZN(n4384) );
  OAI21_X1 U3958 ( .B1(n4164), .B2(n4627), .A(n4384), .ZN(n4669) );
  NAND2_X1 U3959 ( .A1(n4798), .A2(n4669), .ZN(n3091) );
  INV_X1 U3960 ( .A(n3095), .ZN(n3100) );
  AOI21_X1 U3961 ( .B1(n3096), .B2(n3098), .A(n3097), .ZN(n3099) );
  NOR3_X1 U3962 ( .A1(n3100), .A2(n3099), .A3(n4109), .ZN(n3106) );
  NOR2_X1 U3963 ( .A1(n4122), .A2(n4504), .ZN(n3105) );
  NOR2_X1 U3964 ( .A1(n4043), .A2(n4082), .ZN(n3104) );
  NAND2_X1 U3965 ( .A1(n4457), .A2(n4117), .ZN(n3102) );
  NAND2_X1 U3966 ( .A1(U3149), .A2(REG3_REG_23__SCAN_IN), .ZN(n3101) );
  OAI211_X1 U3967 ( .C1(n4096), .C2(n4503), .A(n3102), .B(n3101), .ZN(n3103)
         );
  OR4_X1 U3968 ( .A1(n3106), .A2(n3105), .A3(n3104), .A4(n3103), .ZN(U3213) );
  INV_X1 U3969 ( .A(DATAI_1_), .ZN(n3107) );
  MUX2_X1 U3970 ( .A(n3383), .B(n3107), .S(U3149), .Z(n3108) );
  INV_X1 U3971 ( .A(n3108), .ZN(U3351) );
  MUX2_X1 U3972 ( .A(n3109), .B(n3409), .S(STATE_REG_SCAN_IN), .Z(n3110) );
  INV_X1 U3973 ( .A(n3110), .ZN(U3348) );
  MUX2_X1 U3974 ( .A(n3111), .B(n3446), .S(STATE_REG_SCAN_IN), .Z(n3112) );
  INV_X1 U3975 ( .A(n3112), .ZN(U3345) );
  INV_X1 U3976 ( .A(DATAI_2_), .ZN(n3113) );
  MUX2_X1 U3977 ( .A(n3386), .B(n3113), .S(U3149), .Z(n3114) );
  INV_X1 U3978 ( .A(n3114), .ZN(U3350) );
  INV_X1 U3979 ( .A(DATAI_17_), .ZN(n3345) );
  NAND2_X1 U3980 ( .A1(n4368), .A2(STATE_REG_SCAN_IN), .ZN(n3115) );
  OAI21_X1 U3981 ( .B1(STATE_REG_SCAN_IN), .B2(n3345), .A(n3115), .ZN(U3335)
         );
  INV_X1 U3982 ( .A(DATAI_10_), .ZN(n3116) );
  INV_X1 U3983 ( .A(n3773), .ZN(n3777) );
  MUX2_X1 U3984 ( .A(n3116), .B(n3777), .S(STATE_REG_SCAN_IN), .Z(n3117) );
  INV_X1 U3985 ( .A(n3117), .ZN(U3342) );
  INV_X1 U3986 ( .A(DATAI_30_), .ZN(n3308) );
  NAND2_X1 U3987 ( .A1(n3118), .A2(STATE_REG_SCAN_IN), .ZN(n3119) );
  OAI21_X1 U3988 ( .B1(STATE_REG_SCAN_IN), .B2(n3308), .A(n3119), .ZN(U3322)
         );
  INV_X1 U3989 ( .A(DATAI_27_), .ZN(n3222) );
  NAND2_X1 U3990 ( .A1(n4821), .A2(STATE_REG_SCAN_IN), .ZN(n3120) );
  OAI21_X1 U3991 ( .B1(STATE_REG_SCAN_IN), .B2(n3222), .A(n3120), .ZN(U3325)
         );
  INV_X1 U3992 ( .A(DATAO_REG_3__SCAN_IN), .ZN(n3469) );
  INV_X1 U3993 ( .A(n3121), .ZN(n3132) );
  INV_X1 U3994 ( .A(REG2_REG_25__SCAN_IN), .ZN(n3320) );
  NAND4_X1 U3995 ( .A1(REG2_REG_17__SCAN_IN), .A2(ADDR_REG_19__SCAN_IN), .A3(
        n3320), .A4(n4828), .ZN(n3131) );
  INV_X1 U3996 ( .A(ADDR_REG_7__SCAN_IN), .ZN(n3335) );
  NAND4_X1 U3997 ( .A1(ADDR_REG_0__SCAN_IN), .A2(ADDR_REG_6__SCAN_IN), .A3(
        n3680), .A4(n3335), .ZN(n3122) );
  NOR3_X1 U3998 ( .A1(ADDR_REG_5__SCAN_IN), .A2(n4830), .A3(n3122), .ZN(n3123)
         );
  INV_X1 U3999 ( .A(REG3_REG_3__SCAN_IN), .ZN(n3587) );
  NAND3_X1 U4000 ( .A1(DATAI_17_), .A2(n3123), .A3(n3587), .ZN(n3130) );
  INV_X1 U4001 ( .A(DATAI_20_), .ZN(n3346) );
  NOR4_X1 U4002 ( .A1(REG2_REG_27__SCAN_IN), .A2(REG2_REG_31__SCAN_IN), .A3(
        n3346), .A4(n3308), .ZN(n3125) );
  NOR4_X1 U4003 ( .A1(B_REG_SCAN_IN), .A2(REG3_REG_28__SCAN_IN), .A3(n4062), 
        .A4(n4073), .ZN(n3124) );
  NAND4_X1 U4004 ( .A1(n4364), .A2(ADDR_REG_3__SCAN_IN), .A3(n3125), .A4(n3124), .ZN(n3127) );
  INV_X1 U4005 ( .A(REG2_REG_19__SCAN_IN), .ZN(n3126) );
  OR4_X1 U4006 ( .A1(n3128), .A2(n3127), .A3(REG3_REG_0__SCAN_IN), .A4(n3126), 
        .ZN(n3129) );
  NOR4_X1 U4007 ( .A1(n3132), .A2(n3131), .A3(n3130), .A4(n3129), .ZN(n3169)
         );
  INV_X1 U4008 ( .A(DATAI_5_), .ZN(n3243) );
  AND4_X1 U4009 ( .A1(n3244), .A2(n2656), .A3(n3243), .A4(
        DATAO_REG_18__SCAN_IN), .ZN(n3138) );
  INV_X1 U4010 ( .A(ADDR_REG_15__SCAN_IN), .ZN(n4866) );
  INV_X1 U4011 ( .A(DATAI_26_), .ZN(n3241) );
  INV_X1 U4012 ( .A(DATAO_REG_15__SCAN_IN), .ZN(n3486) );
  AND4_X1 U4013 ( .A1(IR_REG_10__SCAN_IN), .A2(n4866), .A3(n3241), .A4(n3486), 
        .ZN(n3137) );
  INV_X1 U4014 ( .A(DATAI_28_), .ZN(n4818) );
  NAND4_X1 U4015 ( .A1(ADDR_REG_13__SCAN_IN), .A2(DATAO_REG_23__SCAN_IN), .A3(
        n3255), .A4(n4818), .ZN(n3135) );
  NAND3_X1 U4016 ( .A1(n3133), .A2(IR_REG_21__SCAN_IN), .A3(DATAI_24_), .ZN(
        n3134) );
  NOR2_X1 U4017 ( .A1(n3135), .A2(n3134), .ZN(n3136) );
  INV_X1 U4018 ( .A(DATAO_REG_13__SCAN_IN), .ZN(n3460) );
  AND4_X1 U4019 ( .A1(n3138), .A2(n3137), .A3(n3136), .A4(n3460), .ZN(n3168)
         );
  INV_X1 U4020 ( .A(DATAI_14_), .ZN(n3220) );
  INV_X1 U4021 ( .A(DATAO_REG_8__SCAN_IN), .ZN(n3473) );
  NAND4_X1 U4022 ( .A1(REG3_REG_8__SCAN_IN), .A2(DATAI_8_), .A3(n3220), .A4(
        n3473), .ZN(n3143) );
  INV_X1 U4023 ( .A(DATAO_REG_4__SCAN_IN), .ZN(n3456) );
  NAND4_X1 U4024 ( .A1(DATAO_REG_16__SCAN_IN), .A2(DATAO_REG_31__SCAN_IN), 
        .A3(n3222), .A4(n3456), .ZN(n3142) );
  INV_X1 U4025 ( .A(DATAI_21_), .ZN(n3139) );
  INV_X1 U4026 ( .A(DATAI_25_), .ZN(n3230) );
  INV_X1 U4027 ( .A(DATAO_REG_30__SCAN_IN), .ZN(n3467) );
  NAND4_X1 U4028 ( .A1(IR_REG_22__SCAN_IN), .A2(n3139), .A3(n3230), .A4(n3467), 
        .ZN(n3141) );
  INV_X1 U4029 ( .A(DATAO_REG_28__SCAN_IN), .ZN(n3839) );
  INV_X1 U4030 ( .A(DATAO_REG_5__SCAN_IN), .ZN(n3475) );
  INV_X1 U4031 ( .A(DATAO_REG_22__SCAN_IN), .ZN(n3490) );
  INV_X1 U4032 ( .A(DATAO_REG_27__SCAN_IN), .ZN(n3786) );
  NAND4_X1 U4033 ( .A1(n3839), .A2(n3475), .A3(n3490), .A4(n3786), .ZN(n3140)
         );
  NOR4_X1 U4034 ( .A1(n3143), .A2(n3142), .A3(n3141), .A4(n3140), .ZN(n3167)
         );
  NOR4_X1 U4035 ( .A1(REG0_REG_3__SCAN_IN), .A2(REG0_REG_8__SCAN_IN), .A3(
        n3271), .A4(n2473), .ZN(n3147) );
  INV_X1 U4036 ( .A(D_REG_2__SCAN_IN), .ZN(n4922) );
  NOR4_X1 U4037 ( .A1(IR_REG_1__SCAN_IN), .A2(REG3_REG_9__SCAN_IN), .A3(
        REG0_REG_14__SCAN_IN), .A4(REG0_REG_13__SCAN_IN), .ZN(n3144) );
  NAND4_X1 U4038 ( .A1(IR_REG_11__SCAN_IN), .A2(IR_REG_3__SCAN_IN), .A3(
        IR_REG_19__SCAN_IN), .A4(n3144), .ZN(n3145) );
  INV_X1 U4039 ( .A(DATAI_13_), .ZN(n4931) );
  NOR4_X1 U4040 ( .A1(n4922), .A2(n3145), .A3(n4931), .A4(DATAI_9_), .ZN(n3146) );
  NAND4_X1 U4041 ( .A1(n3147), .A2(n3146), .A3(D_REG_11__SCAN_IN), .A4(
        D_REG_12__SCAN_IN), .ZN(n3165) );
  INV_X1 U4042 ( .A(REG2_REG_12__SCAN_IN), .ZN(n3332) );
  INV_X1 U40430 ( .A(ADDR_REG_10__SCAN_IN), .ZN(n3333) );
  NOR4_X1 U4044 ( .A1(REG2_REG_10__SCAN_IN), .A2(n3332), .A3(n2671), .A4(n3333), .ZN(n3152) );
  NOR4_X1 U4045 ( .A1(REG3_REG_14__SCAN_IN), .A2(REG1_REG_11__SCAN_IN), .A3(
        REG1_REG_9__SCAN_IN), .A4(n4740), .ZN(n3149) );
  INV_X1 U4046 ( .A(DATAI_15_), .ZN(n4929) );
  INV_X1 U4047 ( .A(REG2_REG_11__SCAN_IN), .ZN(n3877) );
  NOR4_X1 U4048 ( .A1(IR_REG_30__SCAN_IN), .A2(REG2_REG_14__SCAN_IN), .A3(
        n4929), .A4(n3877), .ZN(n3148) );
  NAND2_X1 U4049 ( .A1(n3149), .A2(n3148), .ZN(n3150) );
  NOR4_X1 U4050 ( .A1(n3387), .A2(n2544), .A3(n3800), .A4(n3150), .ZN(n3151)
         );
  NAND3_X1 U4051 ( .A1(n3152), .A2(REG2_REG_1__SCAN_IN), .A3(n3151), .ZN(n3164) );
  INV_X1 U4052 ( .A(REG2_REG_26__SCAN_IN), .ZN(n3186) );
  NOR4_X1 U4053 ( .A1(REG1_REG_26__SCAN_IN), .A2(n3185), .A3(n3189), .A4(n3186), .ZN(n3157) );
  NOR4_X1 U4054 ( .A1(REG1_REG_30__SCAN_IN), .A2(REG0_REG_30__SCAN_IN), .A3(
        REG0_REG_31__SCAN_IN), .A4(n3188), .ZN(n3153) );
  AND4_X1 U4055 ( .A1(n3154), .A2(IR_REG_20__SCAN_IN), .A3(IR_REG_28__SCAN_IN), 
        .A4(n3153), .ZN(n3156) );
  NOR4_X1 U4056 ( .A1(DATAI_0_), .A2(DATAO_REG_2__SCAN_IN), .A3(
        DATAO_REG_19__SCAN_IN), .A4(DATAO_REG_20__SCAN_IN), .ZN(n3155) );
  NAND4_X1 U4057 ( .A1(n3157), .A2(n3156), .A3(n3155), .A4(
        DATAO_REG_9__SCAN_IN), .ZN(n3163) );
  INV_X1 U4058 ( .A(D_REG_29__SCAN_IN), .ZN(n4909) );
  INV_X1 U4059 ( .A(D_REG_24__SCAN_IN), .ZN(n4911) );
  NOR4_X1 U4060 ( .A1(REG1_REG_16__SCAN_IN), .A2(n4909), .A3(n4911), .A4(n3172), .ZN(n3161) );
  INV_X1 U4061 ( .A(D_REG_21__SCAN_IN), .ZN(n4913) );
  INV_X1 U4062 ( .A(D_REG_5__SCAN_IN), .ZN(n4920) );
  INV_X1 U4063 ( .A(D_REG_18__SCAN_IN), .ZN(n4914) );
  INV_X1 U4064 ( .A(D_REG_6__SCAN_IN), .ZN(n4919) );
  NOR4_X1 U4065 ( .A1(n4913), .A2(n4920), .A3(n4914), .A4(n4919), .ZN(n3160)
         );
  NOR4_X1 U4066 ( .A1(REG1_REG_24__SCAN_IN), .A2(n3183), .A3(n2841), .A4(n4700), .ZN(n3159) );
  NOR4_X1 U4067 ( .A1(REG1_REG_21__SCAN_IN), .A2(n3174), .A3(n3176), .A4(n4776), .ZN(n3158) );
  NAND4_X1 U4068 ( .A1(n3161), .A2(n3160), .A3(n3159), .A4(n3158), .ZN(n3162)
         );
  NOR4_X1 U4069 ( .A1(n3165), .A2(n3164), .A3(n3163), .A4(n3162), .ZN(n3166)
         );
  NAND4_X1 U4070 ( .A1(n3169), .A2(n3168), .A3(n3167), .A4(n3166), .ZN(n3365)
         );
  INV_X1 U4071 ( .A(REG1_REG_16__SCAN_IN), .ZN(n4870) );
  AOI22_X1 U4072 ( .A1(n4909), .A2(keyinput49), .B1(keyinput48), .B2(n4870), 
        .ZN(n3170) );
  OAI221_X1 U4073 ( .B1(n4909), .B2(keyinput49), .C1(n4870), .C2(keyinput48), 
        .A(n3170), .ZN(n3180) );
  AOI22_X1 U4074 ( .A1(n3172), .A2(keyinput79), .B1(n4776), .B2(keyinput60), 
        .ZN(n3171) );
  OAI221_X1 U4075 ( .B1(n3172), .B2(keyinput79), .C1(n4776), .C2(keyinput60), 
        .A(n3171), .ZN(n3179) );
  AOI22_X1 U4076 ( .A1(n4708), .A2(keyinput63), .B1(n3174), .B2(keyinput6), 
        .ZN(n3173) );
  OAI221_X1 U4077 ( .B1(n4708), .B2(keyinput63), .C1(n3174), .C2(keyinput6), 
        .A(n3173), .ZN(n3178) );
  AOI22_X1 U4078 ( .A1(n3176), .A2(keyinput13), .B1(n4700), .B2(keyinput2), 
        .ZN(n3175) );
  OAI221_X1 U4079 ( .B1(n3176), .B2(keyinput13), .C1(n4700), .C2(keyinput2), 
        .A(n3175), .ZN(n3177) );
  NOR4_X1 U4080 ( .A1(n3180), .A2(n3179), .A3(n3178), .A4(n3177), .ZN(n3217)
         );
  AOI22_X1 U4081 ( .A1(n2841), .A2(keyinput15), .B1(keyinput108), .B2(n4696), 
        .ZN(n3181) );
  OAI221_X1 U4082 ( .B1(n2841), .B2(keyinput15), .C1(n4696), .C2(keyinput108), 
        .A(n3181), .ZN(n3193) );
  AOI22_X1 U4083 ( .A1(n3183), .A2(keyinput125), .B1(n4688), .B2(keyinput45), 
        .ZN(n3182) );
  OAI221_X1 U4084 ( .B1(n3183), .B2(keyinput125), .C1(n4688), .C2(keyinput45), 
        .A(n3182), .ZN(n3192) );
  AOI22_X1 U4085 ( .A1(n3186), .A2(keyinput31), .B1(n3185), .B2(keyinput35), 
        .ZN(n3184) );
  OAI221_X1 U4086 ( .B1(n3186), .B2(keyinput31), .C1(n3185), .C2(keyinput35), 
        .A(n3184), .ZN(n3191) );
  AOI22_X1 U4087 ( .A1(n3189), .A2(keyinput76), .B1(n3188), .B2(keyinput42), 
        .ZN(n3187) );
  OAI221_X1 U4088 ( .B1(n3189), .B2(keyinput76), .C1(n3188), .C2(keyinput42), 
        .A(n3187), .ZN(n3190) );
  NOR4_X1 U4089 ( .A1(n3193), .A2(n3192), .A3(n3191), .A4(n3190), .ZN(n3216)
         );
  INV_X1 U4090 ( .A(D_REG_26__SCAN_IN), .ZN(n4910) );
  INV_X1 U4091 ( .A(DATAO_REG_20__SCAN_IN), .ZN(n3488) );
  AOI22_X1 U4092 ( .A1(n4910), .A2(keyinput119), .B1(keyinput111), .B2(n3488), 
        .ZN(n3194) );
  OAI221_X1 U4093 ( .B1(n4910), .B2(keyinput119), .C1(n3488), .C2(keyinput111), 
        .A(n3194), .ZN(n3203) );
  INV_X1 U4094 ( .A(DATAO_REG_9__SCAN_IN), .ZN(n3458) );
  INV_X1 U4095 ( .A(D_REG_8__SCAN_IN), .ZN(n4918) );
  AOI22_X1 U4096 ( .A1(n3458), .A2(keyinput23), .B1(n4918), .B2(keyinput27), 
        .ZN(n3195) );
  OAI221_X1 U4097 ( .B1(n3458), .B2(keyinput23), .C1(n4918), .C2(keyinput27), 
        .A(n3195), .ZN(n3202) );
  INV_X1 U4098 ( .A(REG1_REG_30__SCAN_IN), .ZN(n3461) );
  INV_X1 U4099 ( .A(REG0_REG_30__SCAN_IN), .ZN(n3197) );
  AOI22_X1 U4100 ( .A1(n3461), .A2(keyinput57), .B1(n3197), .B2(keyinput124), 
        .ZN(n3196) );
  OAI221_X1 U4101 ( .B1(n3461), .B2(keyinput57), .C1(n3197), .C2(keyinput124), 
        .A(n3196), .ZN(n3201) );
  XNOR2_X1 U4102 ( .A(REG0_REG_31__SCAN_IN), .B(keyinput99), .ZN(n3199) );
  XNOR2_X1 U4103 ( .A(IR_REG_28__SCAN_IN), .B(keyinput1), .ZN(n3198) );
  NAND2_X1 U4104 ( .A1(n3199), .A2(n3198), .ZN(n3200) );
  NOR4_X1 U4105 ( .A1(n3203), .A2(n3202), .A3(n3201), .A4(n3200), .ZN(n3215)
         );
  INV_X1 U4106 ( .A(DATAO_REG_31__SCAN_IN), .ZN(n3471) );
  AOI22_X1 U4107 ( .A1(n3471), .A2(keyinput25), .B1(n3456), .B2(keyinput38), 
        .ZN(n3204) );
  OAI221_X1 U4108 ( .B1(n3471), .B2(keyinput25), .C1(n3456), .C2(keyinput38), 
        .A(n3204), .ZN(n3213) );
  INV_X1 U4109 ( .A(DATAO_REG_19__SCAN_IN), .ZN(n3484) );
  AOI22_X1 U4110 ( .A1(n3154), .A2(keyinput115), .B1(keyinput51), .B2(n3484), 
        .ZN(n3205) );
  OAI221_X1 U4111 ( .B1(n3154), .B2(keyinput115), .C1(n3484), .C2(keyinput51), 
        .A(n3205), .ZN(n3212) );
  INV_X1 U4112 ( .A(DATAO_REG_2__SCAN_IN), .ZN(n3477) );
  AOI22_X1 U4113 ( .A1(n3477), .A2(keyinput91), .B1(n2479), .B2(keyinput103), 
        .ZN(n3206) );
  OAI221_X1 U4114 ( .B1(n3477), .B2(keyinput91), .C1(n2479), .C2(keyinput103), 
        .A(n3206), .ZN(n3211) );
  INV_X1 U4115 ( .A(IR_REG_8__SCAN_IN), .ZN(n3207) );
  XOR2_X1 U4116 ( .A(n3207), .B(keyinput59), .Z(n3209) );
  XNOR2_X1 U4117 ( .A(IR_REG_20__SCAN_IN), .B(keyinput71), .ZN(n3208) );
  NAND2_X1 U4118 ( .A1(n3209), .A2(n3208), .ZN(n3210) );
  NOR4_X1 U4119 ( .A1(n3213), .A2(n3212), .A3(n3211), .A4(n3210), .ZN(n3214)
         );
  NAND4_X1 U4120 ( .A1(n3217), .A2(n3216), .A3(n3215), .A4(n3214), .ZN(n3363)
         );
  AOI22_X1 U4121 ( .A1(n3490), .A2(keyinput5), .B1(keyinput16), .B2(n3786), 
        .ZN(n3218) );
  OAI221_X1 U4122 ( .B1(n3490), .B2(keyinput5), .C1(n3786), .C2(keyinput16), 
        .A(n3218), .ZN(n3228) );
  AOI22_X1 U4123 ( .A1(n3220), .A2(keyinput33), .B1(keyinput32), .B2(n3473), 
        .ZN(n3219) );
  OAI221_X1 U4124 ( .B1(n3220), .B2(keyinput33), .C1(n3473), .C2(keyinput32), 
        .A(n3219), .ZN(n3227) );
  INV_X1 U4125 ( .A(DATAO_REG_16__SCAN_IN), .ZN(n3479) );
  AOI22_X1 U4126 ( .A1(n3479), .A2(keyinput41), .B1(n3222), .B2(keyinput40), 
        .ZN(n3221) );
  OAI221_X1 U4127 ( .B1(n3479), .B2(keyinput41), .C1(n3222), .C2(keyinput40), 
        .A(n3221), .ZN(n3226) );
  XNOR2_X1 U4128 ( .A(REG3_REG_8__SCAN_IN), .B(keyinput34), .ZN(n3224) );
  XNOR2_X1 U4129 ( .A(keyinput0), .B(DATAI_8_), .ZN(n3223) );
  NAND2_X1 U4130 ( .A1(n3224), .A2(n3223), .ZN(n3225) );
  NOR4_X1 U4131 ( .A1(n3228), .A2(n3227), .A3(n3226), .A4(n3225), .ZN(n3265)
         );
  AOI22_X1 U4132 ( .A1(n3230), .A2(keyinput120), .B1(keyinput114), .B2(n3467), 
        .ZN(n3229) );
  OAI221_X1 U4133 ( .B1(n3230), .B2(keyinput120), .C1(n3467), .C2(keyinput114), 
        .A(n3229), .ZN(n3238) );
  AOI22_X1 U4134 ( .A1(n3475), .A2(keyinput10), .B1(n3839), .B2(keyinput14), 
        .ZN(n3231) );
  OAI221_X1 U4135 ( .B1(n3475), .B2(keyinput10), .C1(n3839), .C2(keyinput14), 
        .A(n3231), .ZN(n3237) );
  XNOR2_X1 U4136 ( .A(IR_REG_10__SCAN_IN), .B(keyinput112), .ZN(n3234) );
  XNOR2_X1 U4137 ( .A(DATAI_21_), .B(keyinput122), .ZN(n3233) );
  XNOR2_X1 U4138 ( .A(IR_REG_22__SCAN_IN), .B(keyinput121), .ZN(n3232) );
  NAND3_X1 U4139 ( .A1(n3234), .A2(n3233), .A3(n3232), .ZN(n3236) );
  XNOR2_X1 U4140 ( .A(n3486), .B(keyinput110), .ZN(n3235) );
  NOR4_X1 U4141 ( .A1(n3238), .A2(n3237), .A3(n3236), .A4(n3235), .ZN(n3264)
         );
  INV_X1 U4142 ( .A(D_REG_16__SCAN_IN), .ZN(n4915) );
  INV_X1 U4143 ( .A(D_REG_23__SCAN_IN), .ZN(n4912) );
  AOI22_X1 U4144 ( .A1(n4915), .A2(keyinput106), .B1(keyinput105), .B2(n4912), 
        .ZN(n3239) );
  OAI221_X1 U4145 ( .B1(n4915), .B2(keyinput106), .C1(n4912), .C2(keyinput105), 
        .A(n3239), .ZN(n3249) );
  AOI22_X1 U4146 ( .A1(n3241), .A2(keyinput104), .B1(keyinput92), .B2(n4866), 
        .ZN(n3240) );
  OAI221_X1 U4147 ( .B1(n3241), .B2(keyinput104), .C1(n4866), .C2(keyinput92), 
        .A(n3240), .ZN(n3248) );
  AOI22_X1 U4148 ( .A1(n3244), .A2(keyinput93), .B1(keyinput88), .B2(n3243), 
        .ZN(n3242) );
  OAI221_X1 U4149 ( .B1(n3244), .B2(keyinput93), .C1(n3243), .C2(keyinput88), 
        .A(n3242), .ZN(n3247) );
  INV_X1 U4150 ( .A(DATAO_REG_18__SCAN_IN), .ZN(n3481) );
  AOI22_X1 U4151 ( .A1(n3481), .A2(keyinput84), .B1(n2656), .B2(keyinput86), 
        .ZN(n3245) );
  OAI221_X1 U4152 ( .B1(n3481), .B2(keyinput84), .C1(n2656), .C2(keyinput86), 
        .A(n3245), .ZN(n3246) );
  NOR4_X1 U4153 ( .A1(n3249), .A2(n3248), .A3(n3247), .A4(n3246), .ZN(n3263)
         );
  INV_X1 U4154 ( .A(IR_REG_21__SCAN_IN), .ZN(n3251) );
  AOI22_X1 U4155 ( .A1(n3251), .A2(keyinput78), .B1(keyinput64), .B2(n3460), 
        .ZN(n3250) );
  OAI221_X1 U4156 ( .B1(n3251), .B2(keyinput78), .C1(n3460), .C2(keyinput64), 
        .A(n3250), .ZN(n3261) );
  INV_X1 U4157 ( .A(ADDR_REG_13__SCAN_IN), .ZN(n3253) );
  INV_X1 U4158 ( .A(DATAO_REG_23__SCAN_IN), .ZN(n3520) );
  AOI22_X1 U4159 ( .A1(n3253), .A2(keyinput54), .B1(keyinput44), .B2(n3520), 
        .ZN(n3252) );
  OAI221_X1 U4160 ( .B1(n3253), .B2(keyinput54), .C1(n3520), .C2(keyinput44), 
        .A(n3252), .ZN(n3260) );
  AOI22_X1 U4161 ( .A1(n3255), .A2(keyinput61), .B1(keyinput52), .B2(n4818), 
        .ZN(n3254) );
  OAI221_X1 U4162 ( .B1(n3255), .B2(keyinput61), .C1(n4818), .C2(keyinput52), 
        .A(n3254), .ZN(n3259) );
  XNOR2_X1 U4163 ( .A(IR_REG_12__SCAN_IN), .B(keyinput80), .ZN(n3257) );
  XNOR2_X1 U4164 ( .A(DATAI_24_), .B(keyinput85), .ZN(n3256) );
  NAND2_X1 U4165 ( .A1(n3257), .A2(n3256), .ZN(n3258) );
  NOR4_X1 U4166 ( .A1(n3261), .A2(n3260), .A3(n3259), .A4(n3258), .ZN(n3262)
         );
  NAND4_X1 U4167 ( .A1(n3265), .A2(n3264), .A3(n3263), .A4(n3262), .ZN(n3362)
         );
  AOI22_X1 U4168 ( .A1(n2510), .A2(keyinput65), .B1(n3267), .B2(keyinput43), 
        .ZN(n3266) );
  OAI221_X1 U4169 ( .B1(n2510), .B2(keyinput65), .C1(n3267), .C2(keyinput43), 
        .A(n3266), .ZN(n3275) );
  AOI22_X1 U4170 ( .A1(n4017), .A2(keyinput46), .B1(keyinput21), .B2(n2473), 
        .ZN(n3268) );
  OAI221_X1 U4171 ( .B1(n4017), .B2(keyinput46), .C1(n2473), .C2(keyinput21), 
        .A(n3268), .ZN(n3274) );
  AOI22_X1 U4172 ( .A1(n4795), .A2(keyinput101), .B1(n4791), .B2(keyinput77), 
        .ZN(n3269) );
  OAI221_X1 U4173 ( .B1(n4795), .B2(keyinput101), .C1(n4791), .C2(keyinput77), 
        .A(n3269), .ZN(n3273) );
  AOI22_X1 U4174 ( .A1(n3271), .A2(keyinput56), .B1(n2617), .B2(keyinput58), 
        .ZN(n3270) );
  OAI221_X1 U4175 ( .B1(n3271), .B2(keyinput56), .C1(n2617), .C2(keyinput58), 
        .A(n3270), .ZN(n3272) );
  NOR4_X1 U4176 ( .A1(n3275), .A2(n3274), .A3(n3273), .A4(n3272), .ZN(n3306)
         );
  AOI22_X1 U4177 ( .A1(n4929), .A2(keyinput100), .B1(keyinput127), .B2(n3993), 
        .ZN(n3276) );
  OAI221_X1 U4178 ( .B1(n4929), .B2(keyinput100), .C1(n3993), .C2(keyinput127), 
        .A(n3276), .ZN(n3284) );
  AOI22_X1 U4179 ( .A1(n3800), .A2(keyinput68), .B1(n3877), .B2(keyinput73), 
        .ZN(n3277) );
  OAI221_X1 U4180 ( .B1(n3800), .B2(keyinput68), .C1(n3877), .C2(keyinput73), 
        .A(n3277), .ZN(n3283) );
  XOR2_X1 U4181 ( .A(n2544), .B(keyinput69), .Z(n3281) );
  XNOR2_X1 U4182 ( .A(REG2_REG_1__SCAN_IN), .B(keyinput3), .ZN(n3280) );
  XNOR2_X1 U4183 ( .A(REG1_REG_2__SCAN_IN), .B(keyinput20), .ZN(n3279) );
  XNOR2_X1 U4184 ( .A(REG1_REG_9__SCAN_IN), .B(keyinput87), .ZN(n3278) );
  NAND4_X1 U4185 ( .A1(n3281), .A2(n3280), .A3(n3279), .A4(n3278), .ZN(n3282)
         );
  NOR3_X1 U4186 ( .A1(n3284), .A2(n3283), .A3(n3282), .ZN(n3305) );
  AOI22_X1 U4187 ( .A1(n4922), .A2(keyinput67), .B1(keyinput107), .B2(n4913), 
        .ZN(n3285) );
  OAI221_X1 U4188 ( .B1(n4922), .B2(keyinput67), .C1(n4913), .C2(keyinput107), 
        .A(n3285), .ZN(n3292) );
  INV_X1 U4189 ( .A(D_REG_11__SCAN_IN), .ZN(n4917) );
  INV_X1 U4190 ( .A(D_REG_12__SCAN_IN), .ZN(n4916) );
  AOI22_X1 U4191 ( .A1(n4917), .A2(keyinput83), .B1(keyinput4), .B2(n4916), 
        .ZN(n3286) );
  OAI221_X1 U4192 ( .B1(n4917), .B2(keyinput83), .C1(n4916), .C2(keyinput4), 
        .A(n3286), .ZN(n3291) );
  AOI22_X1 U4193 ( .A1(n4919), .A2(keyinput17), .B1(keyinput81), .B2(n4911), 
        .ZN(n3287) );
  OAI221_X1 U4194 ( .B1(n4919), .B2(keyinput17), .C1(n4911), .C2(keyinput81), 
        .A(n3287), .ZN(n3290) );
  AOI22_X1 U4195 ( .A1(n4920), .A2(keyinput7), .B1(keyinput90), .B2(n4914), 
        .ZN(n3288) );
  OAI221_X1 U4196 ( .B1(n4920), .B2(keyinput7), .C1(n4914), .C2(keyinput90), 
        .A(n3288), .ZN(n3289) );
  NOR4_X1 U4197 ( .A1(n3292), .A2(n3291), .A3(n3290), .A4(n3289), .ZN(n3304)
         );
  XOR2_X1 U4198 ( .A(n2609), .B(keyinput36), .Z(n3296) );
  XNOR2_X1 U4199 ( .A(IR_REG_11__SCAN_IN), .B(keyinput47), .ZN(n3294) );
  XNOR2_X1 U4200 ( .A(DATAI_9_), .B(keyinput29), .ZN(n3293) );
  NAND4_X1 U4201 ( .A1(n3296), .A2(n3295), .A3(n3294), .A4(n3293), .ZN(n3302)
         );
  XNOR2_X1 U4202 ( .A(IR_REG_3__SCAN_IN), .B(keyinput30), .ZN(n3300) );
  XNOR2_X1 U4203 ( .A(IR_REG_6__SCAN_IN), .B(keyinput39), .ZN(n3299) );
  XNOR2_X1 U4204 ( .A(IR_REG_19__SCAN_IN), .B(keyinput11), .ZN(n3298) );
  XNOR2_X1 U4205 ( .A(DATAI_13_), .B(keyinput50), .ZN(n3297) );
  NAND4_X1 U4206 ( .A1(n3300), .A2(n3299), .A3(n3298), .A4(n3297), .ZN(n3301)
         );
  NOR2_X1 U4207 ( .A1(n3302), .A2(n3301), .ZN(n3303) );
  NAND4_X1 U4208 ( .A1(n3306), .A2(n3305), .A3(n3304), .A4(n3303), .ZN(n3361)
         );
  AOI22_X1 U4209 ( .A1(n4422), .A2(keyinput19), .B1(keyinput97), .B2(n3308), 
        .ZN(n3307) );
  OAI221_X1 U4210 ( .B1(n4422), .B2(keyinput19), .C1(n3308), .C2(keyinput97), 
        .A(n3307), .ZN(n3318) );
  AOI22_X1 U4211 ( .A1(n4062), .A2(keyinput75), .B1(keyinput82), .B2(n4073), 
        .ZN(n3309) );
  OAI221_X1 U4212 ( .B1(n4062), .B2(keyinput75), .C1(n4073), .C2(keyinput82), 
        .A(n3309), .ZN(n3317) );
  AOI22_X1 U4213 ( .A1(n3312), .A2(keyinput9), .B1(keyinput22), .B2(n3311), 
        .ZN(n3310) );
  OAI221_X1 U4214 ( .B1(n3312), .B2(keyinput9), .C1(n3311), .C2(keyinput22), 
        .A(n3310), .ZN(n3316) );
  XNOR2_X1 U4215 ( .A(REG3_REG_0__SCAN_IN), .B(keyinput89), .ZN(n3314) );
  XNOR2_X1 U4216 ( .A(REG3_REG_28__SCAN_IN), .B(keyinput70), .ZN(n3313) );
  NAND2_X1 U4217 ( .A1(n3314), .A2(n3313), .ZN(n3315) );
  NOR4_X1 U4218 ( .A1(n3318), .A2(n3317), .A3(n3316), .A4(n3315), .ZN(n3359)
         );
  AOI22_X1 U4219 ( .A1(keyinput113), .A2(n3320), .B1(keyinput116), .B2(n3469), 
        .ZN(n3319) );
  OAI21_X1 U4220 ( .B1(n3320), .B2(keyinput113), .A(n3319), .ZN(n3330) );
  AOI22_X1 U4221 ( .A1(n4828), .A2(keyinput72), .B1(n3322), .B2(keyinput37), 
        .ZN(n3321) );
  OAI221_X1 U4222 ( .B1(n4828), .B2(keyinput72), .C1(n3322), .C2(keyinput37), 
        .A(n3321), .ZN(n3329) );
  INV_X1 U4223 ( .A(ADDR_REG_3__SCAN_IN), .ZN(n3324) );
  AOI22_X1 U4224 ( .A1(n3126), .A2(keyinput8), .B1(keyinput18), .B2(n3324), 
        .ZN(n3323) );
  OAI221_X1 U4225 ( .B1(n3126), .B2(keyinput8), .C1(n3324), .C2(keyinput18), 
        .A(n3323), .ZN(n3328) );
  INV_X1 U4226 ( .A(ADDR_REG_19__SCAN_IN), .ZN(n3326) );
  AOI22_X1 U4227 ( .A1(n3326), .A2(keyinput102), .B1(n4364), .B2(keyinput24), 
        .ZN(n3325) );
  OAI221_X1 U4228 ( .B1(n3326), .B2(keyinput102), .C1(n4364), .C2(keyinput24), 
        .A(n3325), .ZN(n3327) );
  NOR4_X1 U4229 ( .A1(n3330), .A2(n3329), .A3(n3328), .A4(n3327), .ZN(n3358)
         );
  AOI22_X1 U4230 ( .A1(n3333), .A2(keyinput96), .B1(n3332), .B2(keyinput123), 
        .ZN(n3331) );
  OAI221_X1 U4231 ( .B1(n3333), .B2(keyinput96), .C1(n3332), .C2(keyinput123), 
        .A(n3331), .ZN(n3342) );
  AOI22_X1 U4232 ( .A1(n3335), .A2(keyinput12), .B1(n3819), .B2(keyinput55), 
        .ZN(n3334) );
  OAI221_X1 U4233 ( .B1(n3335), .B2(keyinput12), .C1(n3819), .C2(keyinput55), 
        .A(n3334), .ZN(n3341) );
  AOI22_X1 U4234 ( .A1(n4740), .A2(keyinput94), .B1(keyinput109), .B2(n3954), 
        .ZN(n3336) );
  OAI221_X1 U4235 ( .B1(n4740), .B2(keyinput94), .C1(n3954), .C2(keyinput109), 
        .A(n3336), .ZN(n3340) );
  AOI22_X1 U4236 ( .A1(n2671), .A2(keyinput126), .B1(n3338), .B2(keyinput28), 
        .ZN(n3337) );
  OAI221_X1 U4237 ( .B1(n2671), .B2(keyinput126), .C1(n3338), .C2(keyinput28), 
        .A(n3337), .ZN(n3339) );
  NOR4_X1 U4238 ( .A1(n3342), .A2(n3341), .A3(n3340), .A4(n3339), .ZN(n3357)
         );
  AOI22_X1 U4239 ( .A1(n3587), .A2(keyinput95), .B1(keyinput74), .B2(n3680), 
        .ZN(n3343) );
  OAI221_X1 U4240 ( .B1(n3587), .B2(keyinput95), .C1(n3680), .C2(keyinput74), 
        .A(n3343), .ZN(n3355) );
  AOI22_X1 U4241 ( .A1(n3346), .A2(keyinput98), .B1(keyinput117), .B2(n3345), 
        .ZN(n3344) );
  OAI221_X1 U4242 ( .B1(n3346), .B2(keyinput98), .C1(n3345), .C2(keyinput117), 
        .A(n3344), .ZN(n3354) );
  INV_X1 U4243 ( .A(ADDR_REG_5__SCAN_IN), .ZN(n3349) );
  INV_X1 U4244 ( .A(ADDR_REG_6__SCAN_IN), .ZN(n3348) );
  AOI22_X1 U4245 ( .A1(n3349), .A2(keyinput53), .B1(keyinput66), .B2(n3348), 
        .ZN(n3347) );
  OAI221_X1 U4246 ( .B1(n3349), .B2(keyinput53), .C1(n3348), .C2(keyinput66), 
        .A(n3347), .ZN(n3353) );
  INV_X1 U4247 ( .A(ADDR_REG_0__SCAN_IN), .ZN(n3351) );
  AOI22_X1 U4248 ( .A1(n3351), .A2(keyinput118), .B1(n4830), .B2(keyinput26), 
        .ZN(n3350) );
  OAI221_X1 U4249 ( .B1(n3351), .B2(keyinput118), .C1(n4830), .C2(keyinput26), 
        .A(n3350), .ZN(n3352) );
  NOR4_X1 U4250 ( .A1(n3355), .A2(n3354), .A3(n3353), .A4(n3352), .ZN(n3356)
         );
  NAND4_X1 U4251 ( .A1(n3359), .A2(n3358), .A3(n3357), .A4(n3356), .ZN(n3360)
         );
  NOR4_X1 U4252 ( .A1(n3363), .A2(n3362), .A3(n3361), .A4(n3360), .ZN(n3364)
         );
  OAI221_X1 U4253 ( .B1(keyinput116), .B2(n3469), .C1(keyinput116), .C2(n3365), 
        .A(n3364), .ZN(n3369) );
  NAND2_X1 U4254 ( .A1(U3149), .A2(DATAI_25_), .ZN(n3366) );
  OAI21_X1 U4255 ( .B1(n3367), .B2(U3149), .A(n3366), .ZN(n3368) );
  XNOR2_X1 U4256 ( .A(n3369), .B(n3368), .ZN(U3327) );
  INV_X1 U4257 ( .A(n3531), .ZN(n3370) );
  NAND2_X1 U4258 ( .A1(n3371), .A2(n3370), .ZN(n4921) );
  INV_X1 U4259 ( .A(D_REG_0__SCAN_IN), .ZN(n3375) );
  AND2_X1 U4260 ( .A1(n4924), .A2(n3372), .ZN(n3374) );
  AOI22_X1 U4261 ( .A1(n4921), .A2(n3375), .B1(n3374), .B2(n3373), .ZN(U3458)
         );
  INV_X1 U4262 ( .A(D_REG_1__SCAN_IN), .ZN(n3378) );
  INV_X1 U4263 ( .A(n3376), .ZN(n3377) );
  AOI22_X1 U4264 ( .A1(n4921), .A2(n3378), .B1(n3377), .B2(n4924), .ZN(U3459)
         );
  XNOR2_X1 U4265 ( .A(n3383), .B(REG2_REG_1__SCAN_IN), .ZN(n4298) );
  AND2_X1 U4266 ( .A1(IR_REG_0__SCAN_IN), .A2(REG2_REG_0__SCAN_IN), .ZN(n4308)
         );
  NAND2_X1 U4267 ( .A1(n4298), .A2(n4308), .ZN(n4297) );
  NAND2_X1 U4268 ( .A1(n4299), .A2(REG2_REG_1__SCAN_IN), .ZN(n3379) );
  INV_X1 U4269 ( .A(REG2_REG_2__SCAN_IN), .ZN(n3679) );
  MUX2_X1 U4270 ( .A(n3679), .B(REG2_REG_2__SCAN_IN), .S(n3386), .Z(n4319) );
  NAND2_X1 U4271 ( .A1(n4318), .A2(n4319), .ZN(n4317) );
  OR2_X1 U4272 ( .A1(n3386), .A2(n3679), .ZN(n3380) );
  XNOR2_X1 U4273 ( .A(n3399), .B(REG2_REG_3__SCAN_IN), .ZN(n3398) );
  OR2_X1 U4274 ( .A1(n3381), .A2(U3149), .ZN(n4282) );
  NAND2_X1 U4275 ( .A1(n3531), .A2(n4282), .ZN(n3392) );
  AOI21_X1 U4276 ( .B1(n3382), .B2(n3381), .A(n2518), .ZN(n3390) );
  NOR2_X1 U4277 ( .A1(n4819), .A2(n4305), .ZN(n4309) );
  NAND2_X1 U4278 ( .A1(IR_REG_0__SCAN_IN), .A2(REG1_REG_0__SCAN_IN), .ZN(n4292) );
  AOI21_X1 U4279 ( .B1(n3383), .B2(n4293), .A(n4292), .ZN(n3384) );
  NAND2_X1 U4280 ( .A1(n3385), .A2(n3384), .ZN(n4294) );
  NAND2_X1 U4281 ( .A1(n4294), .A2(n3385), .ZN(n4314) );
  XNOR2_X1 U4282 ( .A(n3386), .B(REG1_REG_2__SCAN_IN), .ZN(n4313) );
  NAND2_X1 U4283 ( .A1(n4314), .A2(n4313), .ZN(n3389) );
  OR2_X1 U4284 ( .A1(n3386), .A2(n3387), .ZN(n3388) );
  XOR2_X1 U4285 ( .A(n3405), .B(REG1_REG_3__SCAN_IN), .Z(n3396) );
  INV_X1 U4286 ( .A(n3390), .ZN(n3391) );
  NOR2_X1 U4287 ( .A1(STATE_REG_SCAN_IN), .A2(n3587), .ZN(n3619) );
  AOI21_X1 U4288 ( .B1(n4883), .B2(ADDR_REG_3__SCAN_IN), .A(n3619), .ZN(n3393)
         );
  OAI21_X1 U4289 ( .B1(n4896), .B2(n3394), .A(n3393), .ZN(n3395) );
  AOI21_X1 U4290 ( .B1(n4877), .B2(n3396), .A(n3395), .ZN(n3397) );
  OAI21_X1 U4291 ( .B1(n3398), .B2(n4856), .A(n3397), .ZN(U3243) );
  NAND2_X1 U4292 ( .A1(n3399), .A2(REG2_REG_3__SCAN_IN), .ZN(n3402) );
  NAND2_X1 U4293 ( .A1(n3400), .A2(n4817), .ZN(n3401) );
  XNOR2_X2 U4294 ( .A(n3403), .B(n3409), .ZN(n4827) );
  MUX2_X1 U4295 ( .A(n2544), .B(REG2_REG_5__SCAN_IN), .S(n4816), .Z(n3433) );
  XNOR2_X1 U4296 ( .A(n3424), .B(REG2_REG_6__SCAN_IN), .ZN(n3418) );
  NAND2_X1 U4297 ( .A1(n3405), .A2(REG1_REG_3__SCAN_IN), .ZN(n3408) );
  NAND2_X1 U4298 ( .A1(n3406), .A2(n4817), .ZN(n3407) );
  NAND2_X1 U4299 ( .A1(n3408), .A2(n3407), .ZN(n3410) );
  MUX2_X1 U4300 ( .A(n2543), .B(REG1_REG_5__SCAN_IN), .S(n4816), .Z(n3436) );
  AND2_X1 U4301 ( .A1(U3149), .A2(REG3_REG_6__SCAN_IN), .ZN(n3829) );
  AOI21_X1 U4302 ( .B1(n4883), .B2(ADDR_REG_6__SCAN_IN), .A(n3829), .ZN(n3414)
         );
  OAI21_X1 U4303 ( .B1(n4896), .B2(n3413), .A(n3414), .ZN(n3415) );
  AOI21_X1 U4304 ( .B1(n3416), .B2(n4877), .A(n3415), .ZN(n3417) );
  OAI21_X1 U4305 ( .B1(n3418), .B2(n4856), .A(n3417), .ZN(U3246) );
  INV_X1 U4306 ( .A(n3446), .ZN(n3447) );
  INV_X1 U4307 ( .A(REG1_REG_7__SCAN_IN), .ZN(n4977) );
  XNOR2_X1 U4308 ( .A(n3447), .B(n4977), .ZN(n3421) );
  XNOR2_X1 U4309 ( .A(n3449), .B(n3421), .ZN(n3431) );
  INV_X1 U4310 ( .A(n4877), .ZN(n4880) );
  INV_X1 U4311 ( .A(n3422), .ZN(n3423) );
  AOI22_X2 U4312 ( .A1(n3424), .A2(REG2_REG_6__SCAN_IN), .B1(n4815), .B2(n3423), .ZN(n3426) );
  MUX2_X1 U4313 ( .A(REG2_REG_7__SCAN_IN), .B(n2587), .S(n3446), .Z(n3425) );
  AOI21_X1 U4314 ( .B1(n3426), .B2(n3425), .A(n4856), .ZN(n3429) );
  OR2_X2 U4315 ( .A1(n3426), .A2(n3425), .ZN(n3443) );
  AND2_X1 U4316 ( .A1(REG3_REG_7__SCAN_IN), .A2(U3149), .ZN(n3576) );
  AOI21_X1 U4317 ( .B1(n4883), .B2(ADDR_REG_7__SCAN_IN), .A(n3576), .ZN(n3427)
         );
  OAI21_X1 U4318 ( .B1(n4896), .B2(n3446), .A(n3427), .ZN(n3428) );
  AOI21_X1 U4319 ( .B1(n3429), .B2(n3443), .A(n3428), .ZN(n3430) );
  OAI21_X1 U4320 ( .B1(n3431), .B2(n4880), .A(n3430), .ZN(U3247) );
  AOI211_X1 U4321 ( .C1(n3434), .C2(n3433), .A(n3432), .B(n4856), .ZN(n3441)
         );
  INV_X1 U4322 ( .A(n4816), .ZN(n3438) );
  AND2_X1 U4323 ( .A1(U3149), .A2(REG3_REG_5__SCAN_IN), .ZN(n3568) );
  AOI21_X1 U4324 ( .B1(n4883), .B2(ADDR_REG_5__SCAN_IN), .A(n3568), .ZN(n3437)
         );
  OAI21_X1 U4325 ( .B1(n4896), .B2(n3438), .A(n3437), .ZN(n3439) );
  OR3_X1 U4326 ( .A1(n3441), .A2(n3440), .A3(n3439), .ZN(U3245) );
  NOR2_X1 U4327 ( .A1(n4883), .A2(U4043), .ZN(U3148) );
  NAND2_X2 U4328 ( .A1(n3443), .A2(n3442), .ZN(n3546) );
  XNOR2_X1 U4329 ( .A(n3547), .B(REG2_REG_8__SCAN_IN), .ZN(n3454) );
  AND2_X1 U4330 ( .A1(REG3_REG_8__SCAN_IN), .A2(U3149), .ZN(n3524) );
  INV_X1 U4331 ( .A(n4814), .ZN(n3444) );
  NOR2_X1 U4332 ( .A1(n4896), .A2(n3444), .ZN(n3445) );
  AOI211_X1 U4333 ( .C1(n4883), .C2(ADDR_REG_8__SCAN_IN), .A(n3524), .B(n3445), 
        .ZN(n3453) );
  NOR2_X1 U4334 ( .A1(n3446), .A2(n4977), .ZN(n3448) );
  INV_X1 U4335 ( .A(n3543), .ZN(n3450) );
  OAI211_X1 U4336 ( .C1(REG1_REG_8__SCAN_IN), .C2(n3451), .A(n3450), .B(n4877), 
        .ZN(n3452) );
  OAI211_X1 U4337 ( .C1(n3454), .C2(n4856), .A(n3453), .B(n3452), .ZN(U3248)
         );
  NAND2_X1 U4338 ( .A1(U4043), .A2(n3620), .ZN(n3455) );
  OAI21_X1 U4339 ( .B1(n3521), .B2(n3456), .A(n3455), .ZN(U3554) );
  NAND2_X1 U4340 ( .A1(U4043), .A2(n3811), .ZN(n3457) );
  OAI21_X1 U4341 ( .B1(U4043), .B2(n3458), .A(n3457), .ZN(U3559) );
  NAND2_X1 U4342 ( .A1(U4043), .A2(n3983), .ZN(n3459) );
  OAI21_X1 U4343 ( .B1(n3521), .B2(n3460), .A(n3459), .ZN(U3563) );
  INV_X1 U4344 ( .A(REG2_REG_30__SCAN_IN), .ZN(n4386) );
  NAND2_X1 U4345 ( .A1(n2525), .A2(REG0_REG_30__SCAN_IN), .ZN(n3464) );
  OR2_X1 U4346 ( .A1(n3462), .A2(n3461), .ZN(n3463) );
  OAI211_X1 U4347 ( .C1(n3465), .C2(n4386), .A(n3464), .B(n3463), .ZN(n4400)
         );
  NAND2_X1 U4348 ( .A1(U4043), .A2(n4400), .ZN(n3466) );
  OAI21_X1 U4349 ( .B1(n3521), .B2(n3467), .A(n3466), .ZN(U3580) );
  NAND2_X1 U4350 ( .A1(U4043), .A2(n3504), .ZN(n3468) );
  OAI21_X1 U4351 ( .B1(U4043), .B2(n3469), .A(n3468), .ZN(U3553) );
  NAND2_X1 U4352 ( .A1(U4043), .A2(n4165), .ZN(n3470) );
  OAI21_X1 U4353 ( .B1(U4043), .B2(n3471), .A(n3470), .ZN(U3581) );
  NAND2_X1 U4354 ( .A1(U4043), .A2(n3796), .ZN(n3472) );
  OAI21_X1 U4355 ( .B1(n3521), .B2(n3473), .A(n3472), .ZN(U3558) );
  NAND2_X1 U4356 ( .A1(U4043), .A2(n3830), .ZN(n3474) );
  OAI21_X1 U4357 ( .B1(n3521), .B2(n3475), .A(n3474), .ZN(U3555) );
  NAND2_X1 U4358 ( .A1(U4043), .A2(n3643), .ZN(n3476) );
  OAI21_X1 U4359 ( .B1(n3521), .B2(n3477), .A(n3476), .ZN(U3552) );
  NAND2_X1 U4360 ( .A1(n4116), .A2(U4043), .ZN(n3478) );
  OAI21_X1 U4361 ( .B1(n3521), .B2(n3479), .A(n3478), .ZN(U3566) );
  NAND2_X1 U4362 ( .A1(n4608), .A2(U4043), .ZN(n3480) );
  OAI21_X1 U4363 ( .B1(n3521), .B2(n3481), .A(n3480), .ZN(U3568) );
  NAND2_X1 U4364 ( .A1(n3482), .A2(U4043), .ZN(n3483) );
  OAI21_X1 U4365 ( .B1(n3521), .B2(n3484), .A(n3483), .ZN(U3569) );
  NAND2_X1 U4366 ( .A1(n4621), .A2(U4043), .ZN(n3485) );
  OAI21_X1 U4367 ( .B1(n3521), .B2(n3486), .A(n3485), .ZN(U3565) );
  NAND2_X1 U4368 ( .A1(n4574), .A2(U4043), .ZN(n3487) );
  OAI21_X1 U4369 ( .B1(n3521), .B2(n3488), .A(n3487), .ZN(U3570) );
  NAND2_X1 U4370 ( .A1(n4532), .A2(U4043), .ZN(n3489) );
  OAI21_X1 U4371 ( .B1(U4043), .B2(n3490), .A(n3489), .ZN(U3572) );
  OR2_X1 U4372 ( .A1(n3491), .A2(n3503), .ZN(n3492) );
  NAND2_X1 U4373 ( .A1(n3493), .A2(n3492), .ZN(n4947) );
  NOR2_X1 U4374 ( .A1(n3495), .A2(n3494), .ZN(n3496) );
  NAND2_X1 U4375 ( .A1(n3497), .A2(n3496), .ZN(n3498) );
  NAND2_X1 U4376 ( .A1(n3498), .A2(n4647), .ZN(n3499) );
  NAND2_X1 U4377 ( .A1(n3500), .A2(n4808), .ZN(n3593) );
  INV_X1 U4378 ( .A(n3593), .ZN(n3501) );
  INV_X1 U4379 ( .A(n4904), .ZN(n3517) );
  INV_X1 U4380 ( .A(n3503), .ZN(n4182) );
  XNOR2_X1 U4381 ( .A(n3502), .B(n4182), .ZN(n3509) );
  AOI22_X1 U4382 ( .A1(n3505), .A2(n4661), .B1(n4622), .B2(n3504), .ZN(n3507)
         );
  NAND2_X1 U4383 ( .A1(n4623), .A2(n3830), .ZN(n3506) );
  OAI211_X1 U4384 ( .C1(n4947), .C2(n3650), .A(n3507), .B(n3506), .ZN(n3508)
         );
  AOI21_X1 U4385 ( .B1(n3509), .B2(n4898), .A(n3508), .ZN(n3510) );
  INV_X1 U4386 ( .A(n3510), .ZN(n4949) );
  INV_X1 U4387 ( .A(n3512), .ZN(n3513) );
  OAI211_X1 U4388 ( .C1(n3511), .C2(n3609), .A(n3513), .B(n4943), .ZN(n4948)
         );
  OAI22_X1 U4389 ( .A1(n4948), .A2(n4808), .B1(n4647), .B2(n3616), .ZN(n3514)
         );
  OAI21_X1 U4390 ( .B1(n4949), .B2(n3514), .A(n4485), .ZN(n3516) );
  NAND2_X1 U4391 ( .A1(n4908), .A2(REG2_REG_4__SCAN_IN), .ZN(n3515) );
  OAI211_X1 U4392 ( .C1(n4947), .C2(n3517), .A(n3516), .B(n3515), .ZN(U3286)
         );
  NAND2_X1 U4393 ( .A1(n3518), .A2(U4043), .ZN(n3519) );
  OAI21_X1 U4394 ( .B1(n3521), .B2(n3520), .A(n3519), .ZN(U3573) );
  XNOR2_X1 U4395 ( .A(n3686), .B(n3687), .ZN(n3523) );
  XNOR2_X1 U4396 ( .A(n3522), .B(n3523), .ZN(n3528) );
  AOI21_X1 U4397 ( .B1(n4117), .B2(n3811), .A(n3524), .ZN(n3526) );
  AOI22_X1 U4398 ( .A1(n3734), .A2(n4119), .B1(n4118), .B2(n4290), .ZN(n3525)
         );
  OAI211_X1 U4399 ( .C1(n4122), .C2(n3735), .A(n3526), .B(n3525), .ZN(n3527)
         );
  AOI21_X1 U4400 ( .B1(n3528), .B2(n2953), .A(n3527), .ZN(n3529) );
  INV_X1 U4401 ( .A(n3529), .ZN(U3218) );
  INV_X1 U4402 ( .A(n3530), .ZN(n3533) );
  NOR3_X1 U4403 ( .A1(n3533), .A2(n3532), .A3(n3531), .ZN(n3631) );
  INV_X1 U4404 ( .A(REG3_REG_0__SCAN_IN), .ZN(n3539) );
  XNOR2_X1 U4405 ( .A(n3535), .B(n3534), .ZN(n4304) );
  OAI22_X1 U4406 ( .A1(n4095), .A2(n2989), .B1(n4304), .B2(n4109), .ZN(n3536)
         );
  AOI21_X1 U4407 ( .B1(n3537), .B2(n4119), .A(n3536), .ZN(n3538) );
  OAI21_X1 U4408 ( .B1(n3631), .B2(n3539), .A(n3538), .ZN(U3229) );
  INV_X1 U4409 ( .A(n3540), .ZN(n3541) );
  XNOR2_X1 U4410 ( .A(n4813), .B(REG1_REG_9__SCAN_IN), .ZN(n3544) );
  AOI211_X1 U4411 ( .C1(n3545), .C2(n3544), .A(n4880), .B(n2192), .ZN(n3554)
         );
  MUX2_X1 U4412 ( .A(n3800), .B(REG2_REG_9__SCAN_IN), .S(n4813), .Z(n3548) );
  AOI211_X1 U4413 ( .C1(n3549), .C2(n3548), .A(n4856), .B(n3657), .ZN(n3553)
         );
  INV_X1 U4414 ( .A(n4813), .ZN(n3551) );
  NOR2_X1 U4415 ( .A1(STATE_REG_SCAN_IN), .A2(n2617), .ZN(n3694) );
  AOI21_X1 U4416 ( .B1(n4883), .B2(ADDR_REG_9__SCAN_IN), .A(n3694), .ZN(n3550)
         );
  OAI21_X1 U4417 ( .B1(n4896), .B2(n3551), .A(n3550), .ZN(n3552) );
  OR3_X1 U4418 ( .A1(n3554), .A2(n3553), .A3(n3552), .ZN(U3249) );
  OAI22_X1 U4419 ( .A1(n3677), .A2(n4095), .B1(n4082), .B2(n2989), .ZN(n3555)
         );
  AOI21_X1 U4420 ( .B1(n2499), .B2(n4119), .A(n3555), .ZN(n3561) );
  OAI21_X1 U4421 ( .B1(n3558), .B2(n3557), .A(n3556), .ZN(n3559) );
  NAND2_X1 U4422 ( .A1(n3559), .A2(n2953), .ZN(n3560) );
  OAI211_X1 U4423 ( .C1(n3631), .C2(n3680), .A(n3561), .B(n3560), .ZN(U3234)
         );
  NAND2_X1 U4424 ( .A1(n3563), .A2(n3564), .ZN(n3565) );
  XOR2_X1 U4425 ( .A(n3562), .B(n3565), .Z(n3566) );
  NAND2_X1 U4426 ( .A1(n3566), .A2(n2953), .ZN(n3570) );
  OAI22_X1 U4427 ( .A1(n4096), .A2(n3602), .B1(n4082), .B2(n3597), .ZN(n3567)
         );
  AOI211_X1 U4428 ( .C1(n4117), .C2(n4291), .A(n3568), .B(n3567), .ZN(n3569)
         );
  OAI211_X1 U4429 ( .C1(n4122), .C2(n3604), .A(n3570), .B(n3569), .ZN(U3224)
         );
  AOI21_X1 U4430 ( .B1(n3572), .B2(n3571), .A(n4109), .ZN(n3574) );
  NAND2_X1 U4431 ( .A1(n3574), .A2(n3573), .ZN(n3578) );
  OAI22_X1 U4432 ( .A1(n4096), .A2(n3700), .B1(n4082), .B2(n3714), .ZN(n3575)
         );
  AOI211_X1 U4433 ( .C1(n4117), .C2(n3796), .A(n3576), .B(n3575), .ZN(n3577)
         );
  OAI211_X1 U4434 ( .C1(n4122), .C2(n3709), .A(n3578), .B(n3577), .ZN(U3210)
         );
  INV_X1 U4435 ( .A(n3650), .ZN(n4899) );
  XNOR2_X1 U4436 ( .A(n3579), .B(n4171), .ZN(n4944) );
  OAI21_X1 U4437 ( .B1(n3582), .B2(n3581), .A(n3580), .ZN(n3583) );
  NAND2_X1 U4438 ( .A1(n3583), .A2(n4898), .ZN(n3585) );
  AOI22_X1 U4439 ( .A1(n4661), .A2(n3590), .B1(n4622), .B2(n3643), .ZN(n3584)
         );
  OAI211_X1 U4440 ( .C1(n3597), .C2(n4901), .A(n3585), .B(n3584), .ZN(n3586)
         );
  AOI21_X1 U4441 ( .B1(n4899), .B2(n4944), .A(n3586), .ZN(n4946) );
  OAI22_X1 U4442 ( .A1(n3499), .A2(n3588), .B1(n4647), .B2(REG3_REG_3__SCAN_IN), .ZN(n3589) );
  AOI21_X1 U4443 ( .B1(n4904), .B2(n4944), .A(n3589), .ZN(n3592) );
  AOI21_X1 U4444 ( .B1(n3590), .B2(n3666), .A(n3511), .ZN(n4942) );
  NAND2_X1 U4445 ( .A1(n4664), .A2(n4942), .ZN(n3591) );
  OAI211_X1 U4446 ( .C1(n4946), .C2(n4908), .A(n3592), .B(n3591), .ZN(U3287)
         );
  NAND2_X1 U4447 ( .A1(n3650), .A2(n3593), .ZN(n3594) );
  NAND2_X1 U4448 ( .A1(n4232), .A2(n4217), .ZN(n4169) );
  XNOR2_X1 U4449 ( .A(n3595), .B(n4169), .ZN(n4955) );
  XOR2_X1 U4450 ( .A(n3596), .B(n4169), .Z(n3600) );
  OAI22_X1 U4451 ( .A1(n4650), .A2(n3597), .B1(n4627), .B2(n3602), .ZN(n3598)
         );
  AOI21_X1 U4452 ( .B1(n4623), .B2(n4291), .A(n3598), .ZN(n3599) );
  OAI21_X1 U4453 ( .B1(n3600), .B2(n4655), .A(n3599), .ZN(n4957) );
  NAND2_X1 U4454 ( .A1(n4957), .A2(n4485), .ZN(n3608) );
  OR2_X1 U4455 ( .A1(n3512), .A2(n3602), .ZN(n3603) );
  NAND2_X1 U4456 ( .A1(n3601), .A2(n3603), .ZN(n4954) );
  INV_X1 U4457 ( .A(n4954), .ZN(n3606) );
  OAI22_X1 U4458 ( .A1(n4485), .A2(n2544), .B1(n3604), .B2(n4647), .ZN(n3605)
         );
  AOI21_X1 U4459 ( .B1(n4664), .B2(n3606), .A(n3605), .ZN(n3607) );
  OAI211_X1 U4460 ( .C1(n4666), .C2(n4955), .A(n3608), .B(n3607), .ZN(U3285)
         );
  AND2_X1 U4461 ( .A1(U3149), .A2(REG3_REG_4__SCAN_IN), .ZN(n4834) );
  OAI22_X1 U4462 ( .A1(n4096), .A2(n3609), .B1(n4082), .B2(n3677), .ZN(n3610)
         );
  AOI211_X1 U4463 ( .C1(n4117), .C2(n3830), .A(n4834), .B(n3610), .ZN(n3615)
         );
  AND2_X1 U4464 ( .A1(n3621), .A2(n3611), .ZN(n3613) );
  OAI211_X1 U4465 ( .C1(n3613), .C2(n3612), .A(n2953), .B(n3563), .ZN(n3614)
         );
  OAI211_X1 U4466 ( .C1(n4122), .C2(n3616), .A(n3615), .B(n3614), .ZN(U3227)
         );
  OAI22_X1 U4467 ( .A1(n4096), .A2(n3617), .B1(n4082), .B2(n2988), .ZN(n3618)
         );
  AOI211_X1 U4468 ( .C1(n4117), .C2(n3620), .A(n3619), .B(n3618), .ZN(n3626)
         );
  OAI21_X1 U4469 ( .B1(n3623), .B2(n3622), .A(n3621), .ZN(n3624) );
  NAND2_X1 U4470 ( .A1(n3624), .A2(n2953), .ZN(n3625) );
  OAI211_X1 U4471 ( .C1(REG3_REG_3__SCAN_IN), .C2(n4122), .A(n3626), .B(n3625), 
        .ZN(U3215) );
  XNOR2_X1 U4472 ( .A(n3628), .B(n3627), .ZN(n3635) );
  OAI22_X1 U4473 ( .A1(n2988), .A2(n4095), .B1(n4082), .B2(n3629), .ZN(n3633)
         );
  NOR2_X1 U4474 ( .A1(n3631), .A2(n3630), .ZN(n3632) );
  AOI211_X1 U4475 ( .C1(n2472), .C2(n4119), .A(n3633), .B(n3632), .ZN(n3634)
         );
  OAI21_X1 U4476 ( .B1(n3635), .B2(n4109), .A(n3634), .ZN(U3219) );
  OAI21_X1 U4477 ( .B1(n3636), .B2(n3646), .A(n3664), .ZN(n4936) );
  OAI21_X1 U4478 ( .B1(n3639), .B2(n3638), .A(n3637), .ZN(n4938) );
  INV_X1 U4479 ( .A(n4938), .ZN(n3655) );
  OAI21_X1 U4480 ( .B1(n3640), .B2(n4208), .A(n3641), .ZN(n3642) );
  NAND2_X1 U4481 ( .A1(n3642), .A2(n4898), .ZN(n3649) );
  NAND2_X1 U4482 ( .A1(n4622), .A2(n2991), .ZN(n3645) );
  NAND2_X1 U4483 ( .A1(n4623), .A2(n3643), .ZN(n3644) );
  OAI211_X1 U4484 ( .C1(n3646), .C2(n4627), .A(n3645), .B(n3644), .ZN(n3647)
         );
  INV_X1 U4485 ( .A(n3647), .ZN(n3648) );
  OAI211_X1 U4486 ( .C1(n4938), .C2(n3650), .A(n3649), .B(n3648), .ZN(n4940)
         );
  NAND2_X1 U4487 ( .A1(n4485), .A2(n4940), .ZN(n3652) );
  INV_X1 U4488 ( .A(n4647), .ZN(n4903) );
  NAND2_X1 U4489 ( .A1(n4903), .A2(REG3_REG_1__SCAN_IN), .ZN(n3651) );
  OAI211_X1 U4490 ( .C1(n3499), .C2(n3653), .A(n3652), .B(n3651), .ZN(n3654)
         );
  AOI21_X1 U4491 ( .B1(n4904), .B2(n3655), .A(n3654), .ZN(n3656) );
  OAI21_X1 U4492 ( .B1(n4639), .B2(n4936), .A(n3656), .ZN(U3289) );
  XNOR2_X1 U4493 ( .A(n3775), .B(REG2_REG_10__SCAN_IN), .ZN(n3663) );
  NAND2_X1 U4494 ( .A1(n3658), .A2(REG1_REG_10__SCAN_IN), .ZN(n3776) );
  OAI211_X1 U4495 ( .C1(n3658), .C2(REG1_REG_10__SCAN_IN), .A(n3776), .B(n4877), .ZN(n3662) );
  NOR2_X1 U4496 ( .A1(STATE_REG_SCAN_IN), .A2(n3659), .ZN(n3768) );
  NOR2_X1 U4497 ( .A1(n4896), .A2(n3777), .ZN(n3660) );
  AOI211_X1 U4498 ( .C1(n4883), .C2(ADDR_REG_10__SCAN_IN), .A(n3768), .B(n3660), .ZN(n3661) );
  OAI211_X1 U4499 ( .C1(n3663), .C2(n4856), .A(n3662), .B(n3661), .ZN(U3250)
         );
  NAND2_X1 U4500 ( .A1(n3664), .A2(n2499), .ZN(n3665) );
  NAND2_X1 U4501 ( .A1(n3666), .A2(n3665), .ZN(n3913) );
  NAND2_X1 U4502 ( .A1(n3637), .A2(n3667), .ZN(n3669) );
  NAND2_X1 U4503 ( .A1(n3669), .A2(n3668), .ZN(n3671) );
  NAND2_X1 U4504 ( .A1(n3671), .A2(n3670), .ZN(n3890) );
  INV_X1 U4505 ( .A(n3672), .ZN(n3674) );
  AND3_X1 U4506 ( .A1(n4209), .A2(n4172), .A3(n3641), .ZN(n3673) );
  OAI21_X1 U4507 ( .B1(n3674), .B2(n3673), .A(n4898), .ZN(n3676) );
  AOI22_X1 U4508 ( .A1(n4661), .A2(n2499), .B1(n4622), .B2(n2990), .ZN(n3675)
         );
  OAI211_X1 U4509 ( .C1(n3677), .C2(n4901), .A(n3676), .B(n3675), .ZN(n3678)
         );
  AOI21_X1 U4510 ( .B1(n4899), .B2(n3890), .A(n3678), .ZN(n3888) );
  MUX2_X1 U4511 ( .A(n3679), .B(n3888), .S(n3499), .Z(n3683) );
  NOR2_X1 U4512 ( .A1(n4647), .A2(n3680), .ZN(n3681) );
  AOI21_X1 U4513 ( .B1(n4904), .B2(n3890), .A(n3681), .ZN(n3682) );
  OAI211_X1 U4514 ( .C1(n4639), .C2(n3913), .A(n3683), .B(n3682), .ZN(U3288)
         );
  XNOR2_X1 U4515 ( .A(n3685), .B(n3684), .ZN(n3692) );
  INV_X1 U4516 ( .A(n3522), .ZN(n3690) );
  OAI21_X1 U4517 ( .B1(n3522), .B2(n3687), .A(n3686), .ZN(n3688) );
  OAI21_X1 U4518 ( .B1(n3690), .B2(n3689), .A(n3688), .ZN(n3691) );
  NOR2_X1 U4519 ( .A1(n3691), .A2(n3692), .ZN(n3761) );
  AOI21_X1 U4520 ( .B1(n3692), .B2(n3691), .A(n3761), .ZN(n3698) );
  OAI22_X1 U4521 ( .A1(n4096), .A2(n3801), .B1(n4095), .B2(n3794), .ZN(n3693)
         );
  AOI211_X1 U4522 ( .C1(n4118), .C2(n3796), .A(n3694), .B(n3693), .ZN(n3697)
         );
  INV_X1 U4523 ( .A(n3695), .ZN(n3804) );
  NAND2_X1 U4524 ( .A1(n4086), .A2(n3804), .ZN(n3696) );
  OAI211_X1 U4525 ( .C1(n3698), .C2(n4109), .A(n3697), .B(n3696), .ZN(U3228)
         );
  XNOR2_X1 U4526 ( .A(n3699), .B(n3716), .ZN(n3703) );
  OAI22_X1 U4527 ( .A1(n4650), .A2(n3714), .B1(n3700), .B2(n4627), .ZN(n3701)
         );
  AOI21_X1 U4528 ( .B1(n4623), .B2(n3796), .A(n3701), .ZN(n3702) );
  OAI21_X1 U4529 ( .B1(n3703), .B2(n4655), .A(n3702), .ZN(n4962) );
  INV_X1 U4530 ( .A(n4962), .ZN(n3721) );
  NAND2_X1 U4531 ( .A1(n3705), .A2(n3706), .ZN(n3707) );
  NAND2_X1 U4532 ( .A1(n3707), .A2(n4943), .ZN(n3708) );
  NOR2_X1 U4533 ( .A1(n3704), .A2(n3708), .ZN(n4963) );
  OAI22_X1 U4534 ( .A1(n4485), .A2(n2587), .B1(n3709), .B2(n4647), .ZN(n3719)
         );
  NAND2_X1 U4535 ( .A1(n3711), .A2(n3710), .ZN(n3741) );
  INV_X1 U4536 ( .A(n3741), .ZN(n3713) );
  AOI21_X1 U4537 ( .B1(n3741), .B2(n4291), .A(n3831), .ZN(n3712) );
  AOI21_X1 U4538 ( .B1(n3714), .B2(n3713), .A(n3712), .ZN(n3715) );
  NOR2_X1 U4539 ( .A1(n3715), .A2(n3716), .ZN(n4961) );
  INV_X1 U4540 ( .A(n3715), .ZN(n3717) );
  INV_X1 U4541 ( .A(n3716), .ZN(n4222) );
  NOR2_X1 U4542 ( .A1(n3717), .A2(n4222), .ZN(n4960) );
  NOR3_X1 U4543 ( .A1(n4961), .A2(n4960), .A3(n4666), .ZN(n3718) );
  AOI211_X1 U4544 ( .C1(n4600), .C2(n4963), .A(n3719), .B(n3718), .ZN(n3720)
         );
  OAI21_X1 U4545 ( .B1(n4908), .B2(n3721), .A(n3720), .ZN(U3283) );
  INV_X1 U4546 ( .A(n3722), .ZN(n3723) );
  NAND2_X1 U4547 ( .A1(n3741), .A2(n3723), .ZN(n3725) );
  NAND2_X1 U4548 ( .A1(n3725), .A2(n3724), .ZN(n3726) );
  NAND2_X1 U4549 ( .A1(n4226), .A2(n4224), .ZN(n3728) );
  INV_X1 U4550 ( .A(n3728), .ZN(n4181) );
  XNOR2_X1 U4551 ( .A(n3726), .B(n4181), .ZN(n3894) );
  INV_X1 U4552 ( .A(n3894), .ZN(n3740) );
  XNOR2_X1 U4553 ( .A(n3727), .B(n3728), .ZN(n3729) );
  NAND2_X1 U4554 ( .A1(n3729), .A2(n4898), .ZN(n3731) );
  AOI22_X1 U4555 ( .A1(n4661), .A2(n3734), .B1(n4623), .B2(n3811), .ZN(n3730)
         );
  OAI211_X1 U4556 ( .C1(n3732), .C2(n4650), .A(n3731), .B(n3730), .ZN(n3893)
         );
  NAND2_X1 U4557 ( .A1(n3893), .A2(n4485), .ZN(n3739) );
  INV_X1 U4558 ( .A(n3704), .ZN(n3733) );
  AOI21_X1 U4559 ( .B1(n3734), .B2(n3733), .A(n3802), .ZN(n3937) );
  OAI22_X1 U4560 ( .A1(n4485), .A2(n3736), .B1(n3735), .B2(n4647), .ZN(n3737)
         );
  AOI21_X1 U4561 ( .B1(n3937), .B2(n4664), .A(n3737), .ZN(n3738) );
  OAI211_X1 U4562 ( .C1(n4666), .C2(n3740), .A(n3739), .B(n3738), .ZN(U3282)
         );
  INV_X1 U4563 ( .A(n4233), .ZN(n4218) );
  AND2_X1 U4564 ( .A1(n4218), .A2(n4221), .ZN(n4186) );
  XNOR2_X1 U4565 ( .A(n3741), .B(n4186), .ZN(n3859) );
  XNOR2_X1 U4566 ( .A(n3742), .B(n4186), .ZN(n3745) );
  AOI22_X1 U4567 ( .A1(n4661), .A2(n3831), .B1(n4622), .B2(n3830), .ZN(n3744)
         );
  NAND2_X1 U4568 ( .A1(n4623), .A2(n4290), .ZN(n3743) );
  OAI211_X1 U4569 ( .C1(n3745), .C2(n4655), .A(n3744), .B(n3743), .ZN(n3746)
         );
  AOI21_X1 U4570 ( .B1(n4899), .B2(n3859), .A(n3746), .ZN(n3860) );
  NAND2_X1 U4571 ( .A1(n3601), .A2(n3831), .ZN(n3747) );
  NAND2_X1 U4572 ( .A1(n3705), .A2(n3747), .ZN(n3948) );
  INV_X1 U4573 ( .A(n3834), .ZN(n3748) );
  AOI22_X1 U4574 ( .A1(n4908), .A2(REG2_REG_6__SCAN_IN), .B1(n3748), .B2(n4903), .ZN(n3749) );
  OAI21_X1 U4575 ( .B1(n4639), .B2(n3948), .A(n3749), .ZN(n3750) );
  AOI21_X1 U4576 ( .B1(n4904), .B2(n3859), .A(n3750), .ZN(n3751) );
  OAI21_X1 U4577 ( .B1(n3860), .B2(n4908), .A(n3751), .ZN(U3284) );
  NAND2_X1 U4578 ( .A1(n3754), .A2(n3753), .ZN(n3755) );
  XNOR2_X1 U4579 ( .A(n3752), .B(n3755), .ZN(n3756) );
  NAND2_X1 U4580 ( .A1(n3756), .A2(n2953), .ZN(n3760) );
  AND2_X1 U4581 ( .A1(U3149), .A2(REG3_REG_11__SCAN_IN), .ZN(n3781) );
  OAI22_X1 U4582 ( .A1(n4096), .A2(n3757), .B1(n4095), .B2(n3848), .ZN(n3758)
         );
  AOI211_X1 U4583 ( .C1(n4118), .C2(n4289), .A(n3781), .B(n3758), .ZN(n3759)
         );
  OAI211_X1 U4584 ( .C1(n4122), .C2(n3854), .A(n3760), .B(n3759), .ZN(U3233)
         );
  AOI21_X1 U4585 ( .B1(n3763), .B2(n3762), .A(n3761), .ZN(n3766) );
  OAI211_X1 U4586 ( .C1(n3766), .C2(n3765), .A(n2953), .B(n3764), .ZN(n3770)
         );
  OAI22_X1 U4587 ( .A1(n4096), .A2(n2237), .B1(n4095), .B2(n3918), .ZN(n3767)
         );
  AOI211_X1 U4588 ( .C1(n4118), .C2(n3811), .A(n3768), .B(n3767), .ZN(n3769)
         );
  OAI211_X1 U4589 ( .C1(n4122), .C2(n3818), .A(n3770), .B(n3769), .ZN(U3214)
         );
  INV_X1 U4590 ( .A(n3772), .ZN(n3774) );
  AOI22_X2 U4591 ( .A1(n3775), .A2(REG2_REG_10__SCAN_IN), .B1(n3774), .B2(
        n3773), .ZN(n3879) );
  XNOR2_X1 U4592 ( .A(n4811), .B(n3877), .ZN(n3878) );
  XNOR2_X1 U4593 ( .A(n3879), .B(n3878), .ZN(n3784) );
  XNOR2_X1 U4594 ( .A(n4811), .B(REG1_REG_11__SCAN_IN), .ZN(n3778) );
  OAI211_X1 U4595 ( .C1(n3779), .C2(n3778), .A(n3881), .B(n4877), .ZN(n3783)
         );
  NOR2_X1 U4596 ( .A1(n4896), .A2(n4811), .ZN(n3780) );
  AOI211_X1 U4597 ( .C1(n4883), .C2(ADDR_REG_11__SCAN_IN), .A(n3781), .B(n3780), .ZN(n3782) );
  OAI211_X1 U4598 ( .C1(n3784), .C2(n4856), .A(n3783), .B(n3782), .ZN(U3251)
         );
  NAND2_X1 U4599 ( .A1(n4443), .A2(U4043), .ZN(n3785) );
  OAI21_X1 U4600 ( .B1(U4043), .B2(n3786), .A(n3785), .ZN(U3577) );
  XNOR2_X1 U4601 ( .A(n3867), .B(n3866), .ZN(n3788) );
  XNOR2_X1 U4602 ( .A(n3787), .B(n3788), .ZN(n3789) );
  NAND2_X1 U4603 ( .A1(n3789), .A2(n2953), .ZN(n3792) );
  AND2_X1 U4604 ( .A1(U3149), .A2(REG3_REG_12__SCAN_IN), .ZN(n3884) );
  OAI22_X1 U4605 ( .A1(n4096), .A2(n3930), .B1(n4095), .B2(n3919), .ZN(n3790)
         );
  AOI211_X1 U4606 ( .C1(n4118), .C2(n4288), .A(n3884), .B(n3790), .ZN(n3791)
         );
  OAI211_X1 U4607 ( .C1(n4122), .C2(n3932), .A(n3792), .B(n3791), .ZN(U3221)
         );
  AND2_X1 U4608 ( .A1(n2373), .A2(n4227), .ZN(n4184) );
  XNOR2_X1 U4609 ( .A(n2154), .B(n4184), .ZN(n3900) );
  INV_X1 U4610 ( .A(n3900), .ZN(n3807) );
  XNOR2_X1 U4611 ( .A(n3793), .B(n4184), .ZN(n3798) );
  OAI22_X1 U4612 ( .A1(n4901), .A2(n3794), .B1(n4627), .B2(n3801), .ZN(n3795)
         );
  AOI21_X1 U4613 ( .B1(n4622), .B2(n3796), .A(n3795), .ZN(n3797) );
  OAI21_X1 U4614 ( .B1(n3798), .B2(n4655), .A(n3797), .ZN(n3899) );
  INV_X1 U4615 ( .A(n3899), .ZN(n3799) );
  MUX2_X1 U4616 ( .A(n3800), .B(n3799), .S(n3499), .Z(n3806) );
  OR2_X1 U4617 ( .A1(n3802), .A2(n3801), .ZN(n3803) );
  AND2_X1 U4618 ( .A1(n3816), .A2(n3803), .ZN(n3940) );
  AOI22_X1 U4619 ( .A1(n3940), .A2(n4664), .B1(n3804), .B2(n4903), .ZN(n3805)
         );
  OAI211_X1 U4620 ( .C1(n4666), .C2(n3807), .A(n3806), .B(n3805), .ZN(U3281)
         );
  NAND2_X1 U4621 ( .A1(n4236), .A2(n4238), .ZN(n4170) );
  XNOR2_X1 U4622 ( .A(n3809), .B(n4170), .ZN(n3897) );
  INV_X1 U4623 ( .A(n3897), .ZN(n3823) );
  XNOR2_X1 U4624 ( .A(n3810), .B(n4170), .ZN(n3814) );
  AOI22_X1 U4625 ( .A1(n3817), .A2(n4661), .B1(n4622), .B2(n3811), .ZN(n3813)
         );
  NAND2_X1 U4626 ( .A1(n4623), .A2(n4288), .ZN(n3812) );
  OAI211_X1 U4627 ( .C1(n3814), .C2(n4655), .A(n3813), .B(n3812), .ZN(n3896)
         );
  NAND2_X1 U4628 ( .A1(n3896), .A2(n4485), .ZN(n3822) );
  AOI21_X1 U4629 ( .B1(n3817), .B2(n3816), .A(n3815), .ZN(n3944) );
  OAI22_X1 U4630 ( .A1(n4485), .A2(n3819), .B1(n3818), .B2(n4647), .ZN(n3820)
         );
  AOI21_X1 U4631 ( .B1(n3944), .B2(n4664), .A(n3820), .ZN(n3821) );
  OAI211_X1 U4632 ( .C1(n4666), .C2(n3823), .A(n3822), .B(n3821), .ZN(U3280)
         );
  AND2_X1 U4633 ( .A1(n3825), .A2(n2188), .ZN(n3828) );
  NAND2_X1 U4634 ( .A1(n2412), .A2(n3826), .ZN(n3827) );
  XNOR2_X1 U4635 ( .A(n3828), .B(n3827), .ZN(n3836) );
  AOI21_X1 U4636 ( .B1(n4117), .B2(n4290), .A(n3829), .ZN(n3833) );
  AOI22_X1 U4637 ( .A1(n3831), .A2(n4119), .B1(n4118), .B2(n3830), .ZN(n3832)
         );
  OAI211_X1 U4638 ( .C1(n4122), .C2(n3834), .A(n3833), .B(n3832), .ZN(n3835)
         );
  AOI21_X1 U4639 ( .B1(n3836), .B2(n2953), .A(n3835), .ZN(n3837) );
  INV_X1 U4640 ( .A(n3837), .ZN(U3236) );
  NAND2_X1 U4641 ( .A1(n4430), .A2(U4043), .ZN(n3838) );
  OAI21_X1 U4642 ( .B1(n3839), .B2(U4043), .A(n3838), .ZN(U3578) );
  XNOR2_X1 U4643 ( .A(n4180), .B(n3840), .ZN(n3851) );
  OR2_X1 U4644 ( .A1(n3809), .A2(n3841), .ZN(n3844) );
  AND2_X1 U4645 ( .A1(n3844), .A2(n3842), .ZN(n3846) );
  NAND2_X1 U4646 ( .A1(n3844), .A2(n3843), .ZN(n3845) );
  OAI21_X1 U4647 ( .B1(n3846), .B2(n4180), .A(n3845), .ZN(n3953) );
  AOI22_X1 U4648 ( .A1(n3852), .A2(n4661), .B1(n4622), .B2(n4289), .ZN(n3847)
         );
  OAI21_X1 U4649 ( .B1(n3848), .B2(n4901), .A(n3847), .ZN(n3849) );
  AOI21_X1 U4650 ( .B1(n3953), .B2(n4899), .A(n3849), .ZN(n3850) );
  OAI21_X1 U4651 ( .B1(n3851), .B2(n4655), .A(n3850), .ZN(n3952) );
  INV_X1 U4652 ( .A(n3952), .ZN(n3858) );
  NAND2_X1 U4653 ( .A1(n2235), .A2(n3852), .ZN(n3853) );
  NAND2_X1 U4654 ( .A1(n3928), .A2(n3853), .ZN(n3959) );
  NOR2_X1 U4655 ( .A1(n3959), .A2(n4639), .ZN(n3856) );
  OAI22_X1 U4656 ( .A1(n4485), .A2(n3877), .B1(n3854), .B2(n4647), .ZN(n3855)
         );
  AOI211_X1 U4657 ( .C1(n3953), .C2(n4904), .A(n3856), .B(n3855), .ZN(n3857)
         );
  OAI21_X1 U4658 ( .B1(n3858), .B2(n4908), .A(n3857), .ZN(U3279) );
  INV_X1 U4659 ( .A(n3859), .ZN(n3861) );
  OAI21_X1 U4660 ( .B1(n4937), .B2(n3861), .A(n3860), .ZN(n3950) );
  OAI22_X1 U4661 ( .A1(n4747), .A2(n3948), .B1(n4975), .B2(n3420), .ZN(n3862)
         );
  AOI21_X1 U4662 ( .B1(n3950), .B2(n4975), .A(n3862), .ZN(n3863) );
  INV_X1 U4663 ( .A(n3863), .ZN(U3524) );
  NAND2_X1 U4664 ( .A1(n3865), .A2(n3864), .ZN(n3872) );
  INV_X1 U4665 ( .A(n3787), .ZN(n3870) );
  OAI21_X1 U4666 ( .B1(n3787), .B2(n3867), .A(n3866), .ZN(n3868) );
  OAI21_X1 U4667 ( .B1(n3870), .B2(n3869), .A(n3868), .ZN(n3871) );
  XOR2_X1 U4668 ( .A(n3872), .B(n3871), .Z(n3876) );
  NOR2_X1 U4669 ( .A1(STATE_REG_SCAN_IN), .A2(n2671), .ZN(n4844) );
  OAI22_X1 U4670 ( .A1(n3973), .A2(n4096), .B1(n4095), .B2(n4651), .ZN(n3873)
         );
  AOI211_X1 U4671 ( .C1(n4118), .C2(n4287), .A(n4844), .B(n3873), .ZN(n3875)
         );
  NAND2_X1 U4672 ( .A1(n4086), .A2(n3976), .ZN(n3874) );
  OAI211_X1 U4673 ( .C1(n3876), .C2(n4109), .A(n3875), .B(n3874), .ZN(U3231)
         );
  OAI22_X2 U4674 ( .A1(n3879), .A2(n3878), .B1(n4811), .B2(n3877), .ZN(n4323)
         );
  XNOR2_X1 U4675 ( .A(n4326), .B(n3332), .ZN(n3887) );
  INV_X1 U4676 ( .A(n4810), .ZN(n4324) );
  XNOR2_X1 U4677 ( .A(n4330), .B(n4324), .ZN(n3882) );
  OAI211_X1 U4678 ( .C1(n3882), .C2(REG1_REG_12__SCAN_IN), .A(n4332), .B(n4877), .ZN(n3886) );
  NOR2_X1 U4679 ( .A1(n4896), .A2(n4324), .ZN(n3883) );
  AOI211_X1 U4680 ( .C1(n4883), .C2(ADDR_REG_12__SCAN_IN), .A(n3884), .B(n3883), .ZN(n3885) );
  OAI211_X1 U4681 ( .C1(n3887), .C2(n4856), .A(n3886), .B(n3885), .ZN(U3252)
         );
  INV_X1 U4682 ( .A(n4937), .ZN(n4951) );
  INV_X1 U4683 ( .A(n3888), .ZN(n3889) );
  AOI21_X1 U4684 ( .B1(n4951), .B2(n3890), .A(n3889), .ZN(n3916) );
  INV_X1 U4685 ( .A(n4747), .ZN(n3901) );
  INV_X1 U4686 ( .A(n3913), .ZN(n3891) );
  AOI22_X1 U4687 ( .A1(n3901), .A2(n3891), .B1(REG1_REG_2__SCAN_IN), .B2(n4976), .ZN(n3892) );
  OAI21_X1 U4688 ( .B1(n3916), .B2(n4976), .A(n3892), .ZN(U3520) );
  AOI21_X1 U4689 ( .B1(n3894), .B2(n4744), .A(n3893), .ZN(n3939) );
  AOI22_X1 U4690 ( .A1(n3937), .A2(n3901), .B1(REG1_REG_8__SCAN_IN), .B2(n4976), .ZN(n3895) );
  OAI21_X1 U4691 ( .B1(n3939), .B2(n4976), .A(n3895), .ZN(U3526) );
  AOI21_X1 U4692 ( .B1(n4744), .B2(n3897), .A(n3896), .ZN(n3946) );
  AOI22_X1 U4693 ( .A1(n3944), .A2(n3901), .B1(REG1_REG_10__SCAN_IN), .B2(
        n4976), .ZN(n3898) );
  OAI21_X1 U4694 ( .B1(n3946), .B2(n4976), .A(n3898), .ZN(U3528) );
  AOI21_X1 U4695 ( .B1(n3900), .B2(n4744), .A(n3899), .ZN(n3942) );
  AOI22_X1 U4696 ( .A1(n3940), .A2(n3901), .B1(REG1_REG_9__SCAN_IN), .B2(n4976), .ZN(n3902) );
  OAI21_X1 U4697 ( .B1(n3942), .B2(n4976), .A(n3902), .ZN(U3527) );
  XNOR2_X1 U4698 ( .A(n3905), .B(n3904), .ZN(n3906) );
  XNOR2_X1 U4699 ( .A(n3903), .B(n3906), .ZN(n3907) );
  NAND2_X1 U4700 ( .A1(n3907), .A2(n2953), .ZN(n3911) );
  AND2_X1 U4701 ( .A1(U3149), .A2(REG3_REG_14__SCAN_IN), .ZN(n4329) );
  INV_X1 U4702 ( .A(n4621), .ZN(n3908) );
  OAI22_X1 U4703 ( .A1(n4096), .A2(n3986), .B1(n4095), .B2(n3908), .ZN(n3909)
         );
  AOI211_X1 U4704 ( .C1(n4118), .C2(n3983), .A(n4329), .B(n3909), .ZN(n3910)
         );
  OAI211_X1 U4705 ( .C1(n4122), .C2(n3992), .A(n3911), .B(n3910), .ZN(U3212)
         );
  INV_X1 U4706 ( .A(REG0_REG_2__SCAN_IN), .ZN(n3912) );
  OAI22_X1 U4707 ( .A1(n4802), .A2(n3913), .B1(n4798), .B2(n3912), .ZN(n3914)
         );
  INV_X1 U4708 ( .A(n3914), .ZN(n3915) );
  OAI21_X1 U4709 ( .B1(n3916), .B2(n4965), .A(n3915), .ZN(U3471) );
  INV_X1 U4710 ( .A(n3960), .ZN(n3917) );
  OR2_X1 U4711 ( .A1(n3917), .A2(n3961), .ZN(n4189) );
  XNOR2_X1 U4712 ( .A(n3962), .B(n4189), .ZN(n3923) );
  OAI22_X1 U4713 ( .A1(n3919), .A2(n4901), .B1(n4650), .B2(n3918), .ZN(n3920)
         );
  AOI21_X1 U4714 ( .B1(n3921), .B2(n4661), .A(n3920), .ZN(n3922) );
  OAI21_X1 U4715 ( .B1(n3923), .B2(n4655), .A(n3922), .ZN(n4742) );
  INV_X1 U4716 ( .A(n4742), .ZN(n3936) );
  OR2_X1 U4717 ( .A1(n3809), .A2(n3924), .ZN(n3926) );
  AND2_X1 U4718 ( .A1(n3926), .A2(n3925), .ZN(n3927) );
  XNOR2_X1 U4719 ( .A(n3927), .B(n4189), .ZN(n4743) );
  INV_X1 U4720 ( .A(n4666), .ZN(n4641) );
  INV_X1 U4721 ( .A(n3928), .ZN(n3931) );
  INV_X1 U4722 ( .A(n3974), .ZN(n3929) );
  OAI21_X1 U4723 ( .B1(n3931), .B2(n3930), .A(n3929), .ZN(n4803) );
  NOR2_X1 U4724 ( .A1(n4803), .A2(n4639), .ZN(n3934) );
  OAI22_X1 U4725 ( .A1(n3499), .A2(n3332), .B1(n3932), .B2(n4647), .ZN(n3933)
         );
  AOI211_X1 U4726 ( .C1(n4743), .C2(n4641), .A(n3934), .B(n3933), .ZN(n3935)
         );
  OAI21_X1 U4727 ( .B1(n3936), .B2(n4908), .A(n3935), .ZN(U3278) );
  INV_X1 U4728 ( .A(n4802), .ZN(n3943) );
  AOI22_X1 U4729 ( .A1(n3937), .A2(n3943), .B1(REG0_REG_8__SCAN_IN), .B2(n4965), .ZN(n3938) );
  OAI21_X1 U4730 ( .B1(n3939), .B2(n4965), .A(n3938), .ZN(U3483) );
  AOI22_X1 U4731 ( .A1(n3940), .A2(n3943), .B1(REG0_REG_9__SCAN_IN), .B2(n4965), .ZN(n3941) );
  OAI21_X1 U4732 ( .B1(n3942), .B2(n4965), .A(n3941), .ZN(U3485) );
  AOI22_X1 U4733 ( .A1(n3944), .A2(n3943), .B1(REG0_REG_10__SCAN_IN), .B2(
        n4965), .ZN(n3945) );
  OAI21_X1 U4734 ( .B1(n3946), .B2(n4965), .A(n3945), .ZN(U3487) );
  INV_X1 U4735 ( .A(REG0_REG_6__SCAN_IN), .ZN(n3947) );
  OAI22_X1 U4736 ( .A1(n4802), .A2(n3948), .B1(n4967), .B2(n3947), .ZN(n3949)
         );
  AOI21_X1 U4737 ( .B1(n3950), .B2(n4798), .A(n3949), .ZN(n3951) );
  INV_X1 U4738 ( .A(n3951), .ZN(U3479) );
  AOI21_X1 U4739 ( .B1(n4951), .B2(n3953), .A(n3952), .ZN(n3956) );
  MUX2_X1 U4740 ( .A(n3954), .B(n3956), .S(n4975), .Z(n3955) );
  OAI21_X1 U4741 ( .B1(n4747), .B2(n3959), .A(n3955), .ZN(U3529) );
  INV_X1 U4742 ( .A(REG0_REG_11__SCAN_IN), .ZN(n3957) );
  MUX2_X1 U4743 ( .A(n3957), .B(n3956), .S(n4967), .Z(n3958) );
  OAI21_X1 U4744 ( .B1(n3959), .B2(n4802), .A(n3958), .ZN(U3489) );
  XNOR2_X1 U4745 ( .A(n3973), .B(n3983), .ZN(n4178) );
  OAI21_X1 U4746 ( .B1(n3962), .B2(n3961), .A(n3960), .ZN(n3963) );
  XOR2_X1 U4747 ( .A(n4178), .B(n3963), .Z(n3971) );
  OR2_X1 U4748 ( .A1(n3809), .A2(n3964), .ZN(n3966) );
  AND2_X1 U4749 ( .A1(n3966), .A2(n3965), .ZN(n3967) );
  XNOR2_X1 U4750 ( .A(n3967), .B(n4178), .ZN(n4739) );
  AOI22_X1 U4751 ( .A1(n4286), .A2(n4623), .B1(n4622), .B2(n4287), .ZN(n3968)
         );
  OAI21_X1 U4752 ( .B1(n3973), .B2(n4627), .A(n3968), .ZN(n3969) );
  AOI21_X1 U4753 ( .B1(n4739), .B2(n4899), .A(n3969), .ZN(n3970) );
  OAI21_X1 U4754 ( .B1(n3971), .B2(n4655), .A(n3970), .ZN(n4738) );
  INV_X1 U4755 ( .A(n4738), .ZN(n3980) );
  OR2_X1 U4756 ( .A1(n3974), .A2(n3973), .ZN(n3975) );
  NAND2_X1 U4757 ( .A1(n3972), .A2(n3975), .ZN(n4797) );
  AOI22_X1 U4758 ( .A1(n4908), .A2(REG2_REG_13__SCAN_IN), .B1(n3976), .B2(
        n4903), .ZN(n3977) );
  OAI21_X1 U4759 ( .B1(n4797), .B2(n4639), .A(n3977), .ZN(n3978) );
  AOI21_X1 U4760 ( .B1(n4739), .B2(n4904), .A(n3978), .ZN(n3979) );
  OAI21_X1 U4761 ( .B1(n3980), .B2(n4908), .A(n3979), .ZN(U3277) );
  XNOR2_X1 U4762 ( .A(n3981), .B(n4176), .ZN(n3982) );
  NAND2_X1 U4763 ( .A1(n3982), .A2(n4898), .ZN(n3985) );
  AOI22_X1 U4764 ( .A1(n4621), .A2(n4623), .B1(n4622), .B2(n3983), .ZN(n3984)
         );
  OAI211_X1 U4765 ( .C1(n4627), .C2(n3986), .A(n3985), .B(n3984), .ZN(n4734)
         );
  INV_X1 U4766 ( .A(n4734), .ZN(n3997) );
  OAI21_X1 U4767 ( .B1(n3987), .B2(n3015), .A(n3988), .ZN(n4735) );
  NAND2_X1 U4768 ( .A1(n3972), .A2(n3990), .ZN(n3991) );
  NAND2_X1 U4769 ( .A1(n4646), .A2(n3991), .ZN(n4793) );
  NOR2_X1 U4770 ( .A1(n4793), .A2(n4639), .ZN(n3995) );
  OAI22_X1 U4771 ( .A1(n3499), .A2(n3993), .B1(n3992), .B2(n4647), .ZN(n3994)
         );
  AOI211_X1 U4772 ( .C1(n4735), .C2(n4641), .A(n3995), .B(n3994), .ZN(n3996)
         );
  OAI21_X1 U4773 ( .B1(n3997), .B2(n4908), .A(n3996), .ZN(U3276) );
  AOI21_X1 U4774 ( .B1(n4113), .B2(n4111), .A(n3998), .ZN(n3999) );
  XOR2_X1 U4775 ( .A(n4000), .B(n3999), .Z(n4005) );
  AND2_X1 U4776 ( .A1(U3149), .A2(REG3_REG_16__SCAN_IN), .ZN(n4868) );
  AOI21_X1 U4777 ( .B1(n4117), .B2(n4624), .A(n4868), .ZN(n4003) );
  AOI22_X1 U4778 ( .A1(n4001), .A2(n4119), .B1(n4118), .B2(n4621), .ZN(n4002)
         );
  OAI211_X1 U4779 ( .C1(n4122), .C2(n4636), .A(n4003), .B(n4002), .ZN(n4004)
         );
  AOI21_X1 U4780 ( .B1(n4005), .B2(n2953), .A(n4004), .ZN(n4006) );
  INV_X1 U4781 ( .A(n4006), .ZN(U3223) );
  XNOR2_X1 U4782 ( .A(n4009), .B(n4008), .ZN(n4010) );
  XNOR2_X1 U4783 ( .A(n4007), .B(n4010), .ZN(n4015) );
  AOI22_X1 U4784 ( .A1(n4011), .A2(n4119), .B1(n4117), .B2(n4608), .ZN(n4012)
         );
  NAND2_X1 U4785 ( .A1(U3149), .A2(REG3_REG_17__SCAN_IN), .ZN(n4360) );
  OAI211_X1 U4786 ( .C1(n4652), .C2(n4082), .A(n4012), .B(n4360), .ZN(n4013)
         );
  AOI21_X1 U4787 ( .B1(n4615), .B2(n4086), .A(n4013), .ZN(n4014) );
  OAI21_X1 U4788 ( .B1(n4015), .B2(n4109), .A(n4014), .ZN(U3225) );
  NAND3_X1 U4789 ( .A1(n4017), .A2(IR_REG_31__SCAN_IN), .A3(STATE_REG_SCAN_IN), 
        .ZN(n4019) );
  INV_X1 U4790 ( .A(DATAI_31_), .ZN(n4018) );
  OAI22_X1 U4791 ( .A1(n4016), .A2(n4019), .B1(STATE_REG_SCAN_IN), .B2(n4018), 
        .ZN(U3321) );
  XNOR2_X1 U4792 ( .A(n4021), .B(n4020), .ZN(n4026) );
  AOI22_X1 U4793 ( .A1(n4119), .A2(n4420), .B1(REG3_REG_27__SCAN_IN), .B2(
        U3149), .ZN(n4023) );
  NAND2_X1 U4794 ( .A1(n4421), .A2(n4086), .ZN(n4022) );
  OAI211_X1 U4795 ( .C1(n4459), .C2(n4082), .A(n4023), .B(n4022), .ZN(n4024)
         );
  AOI21_X1 U4796 ( .B1(n4430), .B2(n4117), .A(n4024), .ZN(n4025) );
  OAI21_X1 U4797 ( .B1(n4026), .B2(n4109), .A(n4025), .ZN(U3211) );
  XOR2_X1 U4798 ( .A(n4027), .B(n4028), .Z(n4035) );
  INV_X1 U4799 ( .A(n4029), .ZN(n4582) );
  AOI22_X1 U4800 ( .A1(n4030), .A2(n4119), .B1(n4118), .B2(n4608), .ZN(n4031)
         );
  NAND2_X1 U4801 ( .A1(U3149), .A2(REG3_REG_19__SCAN_IN), .ZN(n4375) );
  OAI211_X1 U4802 ( .C1(n4032), .C2(n4095), .A(n4031), .B(n4375), .ZN(n4033)
         );
  AOI21_X1 U4803 ( .B1(n4582), .B2(n4086), .A(n4033), .ZN(n4034) );
  OAI21_X1 U4804 ( .B1(n4035), .B2(n4109), .A(n4034), .ZN(U3216) );
  XNOR2_X1 U4805 ( .A(n4038), .B(n4037), .ZN(n4039) );
  XNOR2_X1 U4806 ( .A(n4036), .B(n4039), .ZN(n4046) );
  AOI22_X1 U4807 ( .A1(n4574), .A2(n4118), .B1(REG3_REG_21__SCAN_IN), .B2(
        U3149), .ZN(n4042) );
  NAND2_X1 U4808 ( .A1(n4119), .A2(n4040), .ZN(n4041) );
  OAI211_X1 U4809 ( .C1(n4043), .C2(n4095), .A(n4042), .B(n4041), .ZN(n4044)
         );
  AOI21_X1 U4810 ( .B1(n4538), .B2(n4086), .A(n4044), .ZN(n4045) );
  OAI21_X1 U4811 ( .B1(n4046), .B2(n4109), .A(n4045), .ZN(U3220) );
  NAND2_X1 U4812 ( .A1(n2182), .A2(n4048), .ZN(n4049) );
  XNOR2_X1 U4813 ( .A(n4047), .B(n4049), .ZN(n4055) );
  OAI22_X1 U4814 ( .A1(n4497), .A2(n4082), .B1(STATE_REG_SCAN_IN), .B2(n4050), 
        .ZN(n4051) );
  AOI21_X1 U4815 ( .B1(n4456), .B2(n4119), .A(n4051), .ZN(n4052) );
  OAI21_X1 U4816 ( .B1(n4459), .B2(n4095), .A(n4052), .ZN(n4053) );
  AOI21_X1 U4817 ( .B1(n4465), .B2(n4086), .A(n4053), .ZN(n4054) );
  OAI21_X1 U4818 ( .B1(n4055), .B2(n4109), .A(n4054), .ZN(U3222) );
  INV_X1 U4819 ( .A(n4056), .ZN(n4058) );
  NAND2_X1 U4820 ( .A1(n4058), .A2(n4057), .ZN(n4060) );
  XNOR2_X1 U4821 ( .A(n4060), .B(n4059), .ZN(n4061) );
  NAND2_X1 U4822 ( .A1(n4061), .A2(n2953), .ZN(n4067) );
  OAI22_X1 U4823 ( .A1(n4517), .A2(n4082), .B1(STATE_REG_SCAN_IN), .B2(n4062), 
        .ZN(n4064) );
  NOR2_X1 U4824 ( .A1(n4441), .A2(n4095), .ZN(n4063) );
  AOI211_X1 U4825 ( .C1(n4065), .C2(n4119), .A(n4064), .B(n4063), .ZN(n4066)
         );
  OAI211_X1 U4826 ( .C1(n4122), .C2(n4487), .A(n4067), .B(n4066), .ZN(U3226)
         );
  OR2_X1 U4827 ( .A1(n4070), .A2(n4069), .ZN(n4071) );
  AOI22_X1 U4828 ( .A1(n2168), .A2(n2300), .B1(n4068), .B2(n4071), .ZN(n4077)
         );
  INV_X1 U4829 ( .A(n4072), .ZN(n4560) );
  OAI22_X1 U4830 ( .A1(n4096), .A2(n4558), .B1(n4082), .B2(n4591), .ZN(n4075)
         );
  OAI22_X1 U4831 ( .A1(n4083), .A2(n4095), .B1(STATE_REG_SCAN_IN), .B2(n4073), 
        .ZN(n4074) );
  AOI211_X1 U4832 ( .C1(n4560), .C2(n4086), .A(n4075), .B(n4074), .ZN(n4076)
         );
  OAI21_X1 U4833 ( .B1(n4077), .B2(n4109), .A(n4076), .ZN(U3230) );
  OAI21_X1 U4834 ( .B1(n4079), .B2(n4078), .A(n3096), .ZN(n4080) );
  NAND2_X1 U4835 ( .A1(n4080), .A2(n2953), .ZN(n4088) );
  OAI22_X1 U4836 ( .A1(n4083), .A2(n4082), .B1(STATE_REG_SCAN_IN), .B2(n4081), 
        .ZN(n4085) );
  OAI22_X1 U4837 ( .A1(n4517), .A2(n4095), .B1(n4096), .B2(n4514), .ZN(n4084)
         );
  AOI211_X1 U4838 ( .C1(n4520), .C2(n4086), .A(n4085), .B(n4084), .ZN(n4087)
         );
  NAND2_X1 U4839 ( .A1(n4088), .A2(n4087), .ZN(U3232) );
  INV_X1 U4840 ( .A(n4089), .ZN(n4091) );
  NAND2_X1 U4841 ( .A1(n4091), .A2(n4090), .ZN(n4092) );
  XNOR2_X1 U4842 ( .A(n4093), .B(n4092), .ZN(n4094) );
  NAND2_X1 U4843 ( .A1(n4094), .A2(n2953), .ZN(n4099) );
  AND2_X1 U4844 ( .A1(U3149), .A2(REG3_REG_18__SCAN_IN), .ZN(n4884) );
  OAI22_X1 U4845 ( .A1(n4096), .A2(n4595), .B1(n4095), .B2(n4591), .ZN(n4097)
         );
  AOI211_X1 U4846 ( .C1(n4118), .C2(n4624), .A(n4884), .B(n4097), .ZN(n4098)
         );
  OAI211_X1 U4847 ( .C1(n4122), .C2(n4597), .A(n4099), .B(n4098), .ZN(U3235)
         );
  INV_X1 U4848 ( .A(n4101), .ZN(n4103) );
  NOR2_X1 U4849 ( .A1(n4103), .A2(n4102), .ZN(n4104) );
  XNOR2_X1 U4850 ( .A(n4100), .B(n4104), .ZN(n4110) );
  NAND2_X1 U4851 ( .A1(n4479), .A2(n4118), .ZN(n4106) );
  AOI22_X1 U4852 ( .A1(n4119), .A2(n4446), .B1(REG3_REG_26__SCAN_IN), .B2(
        U3149), .ZN(n4105) );
  OAI211_X1 U4853 ( .C1(n4122), .C2(n4448), .A(n4106), .B(n4105), .ZN(n4107)
         );
  AOI21_X1 U4854 ( .B1(n4443), .B2(n4117), .A(n4107), .ZN(n4108) );
  OAI21_X1 U4855 ( .B1(n4110), .B2(n4109), .A(n4108), .ZN(U3237) );
  INV_X1 U4856 ( .A(n4111), .ZN(n4112) );
  NOR2_X1 U4857 ( .A1(n3998), .A2(n4112), .ZN(n4114) );
  XNOR2_X1 U4858 ( .A(n4114), .B(n4113), .ZN(n4124) );
  NAND2_X1 U4859 ( .A1(U3149), .A2(REG3_REG_15__SCAN_IN), .ZN(n4864) );
  INV_X1 U4860 ( .A(n4864), .ZN(n4115) );
  AOI21_X1 U4861 ( .B1(n4117), .B2(n4116), .A(n4115), .ZN(n4121) );
  AOI22_X1 U4862 ( .A1(n4660), .A2(n4119), .B1(n4118), .B2(n4286), .ZN(n4120)
         );
  OAI211_X1 U4863 ( .C1(n4122), .C2(n4648), .A(n4121), .B(n4120), .ZN(n4123)
         );
  AOI21_X1 U4864 ( .B1(n4124), .B2(n2953), .A(n4123), .ZN(n4125) );
  INV_X1 U4865 ( .A(n4125), .ZN(U3238) );
  INV_X1 U4866 ( .A(n4385), .ZN(n4154) );
  INV_X1 U4867 ( .A(n4165), .ZN(n4153) );
  NAND2_X1 U4868 ( .A1(n4127), .A2(n4126), .ZN(n4244) );
  NAND2_X1 U4869 ( .A1(n4229), .A2(n4230), .ZN(n4128) );
  NAND2_X1 U4870 ( .A1(n4128), .A2(n4127), .ZN(n4246) );
  OAI21_X1 U4871 ( .B1(n3981), .B2(n4244), .A(n4246), .ZN(n4130) );
  INV_X1 U4872 ( .A(n4545), .ZN(n4129) );
  AOI211_X1 U4873 ( .C1(n4130), .C2(n4253), .A(n4129), .B(n4546), .ZN(n4133)
         );
  OAI21_X1 U4874 ( .B1(n4133), .B2(n4132), .A(n4131), .ZN(n4135) );
  INV_X1 U4875 ( .A(n4255), .ZN(n4134) );
  AOI211_X1 U4876 ( .C1(n4135), .C2(n4257), .A(n4134), .B(n4472), .ZN(n4138)
         );
  INV_X1 U4877 ( .A(n4136), .ZN(n4137) );
  NOR2_X1 U4878 ( .A1(n4160), .A2(n2383), .ZN(n4262) );
  OAI21_X1 U4879 ( .B1(n4138), .B2(n4137), .A(n4262), .ZN(n4151) );
  INV_X1 U4880 ( .A(n4139), .ZN(n4140) );
  AND2_X1 U4881 ( .A1(n4140), .A2(n4396), .ZN(n4148) );
  INV_X1 U4882 ( .A(n4148), .ZN(n4144) );
  INV_X1 U4883 ( .A(n4263), .ZN(n4143) );
  INV_X1 U4884 ( .A(n4200), .ZN(n4142) );
  NAND2_X1 U4885 ( .A1(n4165), .A2(n4164), .ZN(n4270) );
  OR2_X1 U4886 ( .A1(n4400), .A2(n4385), .ZN(n4141) );
  AND2_X1 U4887 ( .A1(n4270), .A2(n4141), .ZN(n4146) );
  INV_X1 U4888 ( .A(n4146), .ZN(n4168) );
  NOR4_X1 U4889 ( .A1(n4144), .A2(n4143), .A3(n4142), .A4(n4168), .ZN(n4150)
         );
  NAND2_X1 U4890 ( .A1(n4284), .A2(n4145), .ZN(n4199) );
  NAND2_X1 U4891 ( .A1(n4395), .A2(n4199), .ZN(n4147) );
  NOR2_X1 U4892 ( .A1(n4147), .A2(n4157), .ZN(n4267) );
  OAI211_X1 U4893 ( .C1(n4148), .C2(n4147), .A(n4146), .B(n4200), .ZN(n4205)
         );
  AOI21_X1 U4894 ( .B1(n4426), .B2(n4267), .A(n4205), .ZN(n4149) );
  AOI21_X1 U4895 ( .B1(n4151), .B2(n4150), .A(n4149), .ZN(n4152) );
  AOI21_X1 U4896 ( .B1(n4154), .B2(n4153), .A(n4152), .ZN(n4156) );
  NAND2_X1 U4897 ( .A1(n4400), .A2(n4385), .ZN(n4167) );
  AOI21_X1 U4898 ( .B1(n4167), .B2(n4165), .A(n4164), .ZN(n4155) );
  NOR2_X1 U4899 ( .A1(n4156), .A2(n4155), .ZN(n4277) );
  INV_X1 U4900 ( .A(n4157), .ZN(n4159) );
  NAND2_X1 U4901 ( .A1(n4159), .A2(n4158), .ZN(n4438) );
  NAND2_X1 U4902 ( .A1(n3056), .A2(n4436), .ZN(n4455) );
  NAND2_X1 U4903 ( .A1(n4162), .A2(n4161), .ZN(n4477) );
  INV_X1 U4904 ( .A(n4477), .ZN(n4197) );
  NAND2_X1 U4905 ( .A1(n4473), .A2(n4163), .ZN(n4496) );
  INV_X1 U4906 ( .A(n4496), .ZN(n4196) );
  NAND2_X1 U4907 ( .A1(n4257), .A2(n4255), .ZN(n4528) );
  XNOR2_X1 U4908 ( .A(n4574), .B(n4558), .ZN(n4550) );
  OR2_X1 U4909 ( .A1(n4165), .A2(n4164), .ZN(n4166) );
  NAND2_X1 U4910 ( .A1(n4167), .A2(n4166), .ZN(n4269) );
  NOR2_X1 U4911 ( .A1(n4168), .A2(n4269), .ZN(n4175) );
  NOR2_X1 U4912 ( .A1(n4170), .A2(n4169), .ZN(n4174) );
  NOR2_X1 U4913 ( .A1(n4172), .A2(n4171), .ZN(n4173) );
  NAND4_X1 U4914 ( .A1(n4176), .A2(n4175), .A3(n4174), .A4(n4173), .ZN(n4177)
         );
  NOR3_X1 U4915 ( .A1(n4601), .A2(n4178), .A3(n4177), .ZN(n4193) );
  INV_X1 U4916 ( .A(n4565), .ZN(n4179) );
  AND2_X1 U4917 ( .A1(n4179), .A2(n4566), .ZN(n4611) );
  INV_X1 U4918 ( .A(n4656), .ZN(n4643) );
  INV_X1 U4919 ( .A(n4180), .ZN(n4183) );
  NAND4_X1 U4920 ( .A1(n4184), .A2(n4183), .A3(n4182), .A4(n4181), .ZN(n4188)
         );
  INV_X1 U4921 ( .A(n4208), .ZN(n4185) );
  NAND2_X1 U4922 ( .A1(n3636), .A2(n2991), .ZN(n4207) );
  AND2_X1 U4923 ( .A1(n4185), .A2(n4207), .ZN(n4897) );
  NAND4_X1 U4924 ( .A1(n3640), .A2(n4186), .A3(n4222), .A4(n4897), .ZN(n4187)
         );
  NOR2_X1 U4925 ( .A1(n4188), .A2(n4187), .ZN(n4191) );
  INV_X1 U4926 ( .A(n4189), .ZN(n4190) );
  AND4_X1 U4927 ( .A1(n4611), .A2(n4643), .A3(n4191), .A4(n4190), .ZN(n4192)
         );
  XNOR2_X1 U4928 ( .A(n4591), .B(n4579), .ZN(n4577) );
  NAND4_X1 U4929 ( .A1(n4193), .A2(n4192), .A3(n4577), .A4(n4632), .ZN(n4194)
         );
  NOR3_X1 U4930 ( .A1(n4528), .A2(n4550), .A3(n4194), .ZN(n4195) );
  NAND3_X1 U4931 ( .A1(n4197), .A2(n4196), .A3(n4195), .ZN(n4198) );
  NOR4_X1 U4932 ( .A1(n4438), .A2(n4455), .A3(n4198), .A4(n4511), .ZN(n4201)
         );
  INV_X1 U4933 ( .A(n4677), .ZN(n4674) );
  NAND4_X1 U4934 ( .A1(n4202), .A2(n4201), .A3(n4426), .A4(n4674), .ZN(n4204)
         );
  NAND2_X1 U4935 ( .A1(n4204), .A2(n4203), .ZN(n4274) );
  INV_X1 U4936 ( .A(n4205), .ZN(n4272) );
  OAI211_X1 U4937 ( .C1(n4208), .C2(n2469), .A(n4207), .B(n4206), .ZN(n4210)
         );
  NAND3_X1 U4938 ( .A1(n4210), .A2(n4209), .A3(n3037), .ZN(n4213) );
  NAND3_X1 U4939 ( .A1(n4213), .A2(n4212), .A3(n4211), .ZN(n4216) );
  NAND3_X1 U4940 ( .A1(n4216), .A2(n4215), .A3(n4214), .ZN(n4220) );
  NAND4_X1 U4941 ( .A1(n4220), .A2(n4219), .A3(n4218), .A4(n4217), .ZN(n4223)
         );
  AND3_X1 U4942 ( .A1(n4223), .A2(n4222), .A3(n4221), .ZN(n4228) );
  NAND2_X1 U4943 ( .A1(n4225), .A2(n4224), .ZN(n4234) );
  OAI211_X1 U4944 ( .C1(n4228), .C2(n4234), .A(n4227), .B(n4226), .ZN(n4231)
         );
  NAND4_X1 U4945 ( .A1(n4231), .A2(n4230), .A3(n4229), .A4(n2373), .ZN(n4242)
         );
  NOR4_X1 U4946 ( .A1(n4235), .A2(n4234), .A3(n4233), .A4(n4232), .ZN(n4237)
         );
  OAI21_X1 U4947 ( .B1(n4237), .B2(n2368), .A(n4246), .ZN(n4241) );
  NAND3_X1 U4948 ( .A1(n4245), .A2(n4239), .A3(n4238), .ZN(n4240) );
  AOI21_X1 U4949 ( .B1(n4242), .B2(n4241), .A(n4240), .ZN(n4251) );
  AOI21_X1 U4950 ( .B1(n2377), .B2(n4245), .A(n4244), .ZN(n4249) );
  INV_X1 U4951 ( .A(n4246), .ZN(n4247) );
  AOI21_X1 U4952 ( .B1(n4249), .B2(n4248), .A(n4247), .ZN(n4250) );
  OAI21_X1 U4953 ( .B1(n4251), .B2(n4250), .A(n4545), .ZN(n4254) );
  AOI211_X1 U4954 ( .C1(n4254), .C2(n4253), .A(n4252), .B(n4546), .ZN(n4256)
         );
  OAI21_X1 U4955 ( .B1(n4256), .B2(n2404), .A(n4255), .ZN(n4258) );
  NAND3_X1 U4956 ( .A1(n4258), .A2(n4493), .A3(n4257), .ZN(n4261) );
  INV_X1 U4957 ( .A(n4472), .ZN(n4260) );
  AOI21_X1 U4958 ( .B1(n4261), .B2(n4260), .A(n4259), .ZN(n4265) );
  INV_X1 U4959 ( .A(n4262), .ZN(n4264) );
  OAI21_X1 U4960 ( .B1(n4265), .B2(n4264), .A(n4263), .ZN(n4266) );
  OAI211_X1 U4961 ( .C1(n4420), .C2(n4268), .A(n4267), .B(n4266), .ZN(n4271)
         );
  AOI22_X1 U4962 ( .A1(n4272), .A2(n4271), .B1(n4270), .B2(n4269), .ZN(n4273)
         );
  MUX2_X1 U4963 ( .A(n4274), .B(n4273), .S(n2137), .Z(n4275) );
  OAI21_X1 U4964 ( .B1(n4277), .B2(n4276), .A(n4275), .ZN(n4278) );
  XNOR2_X1 U4965 ( .A(n4278), .B(n4376), .ZN(n4283) );
  NAND2_X1 U4966 ( .A1(n4279), .A2(n4309), .ZN(n4280) );
  OAI211_X1 U4967 ( .C1(n2468), .C2(n4282), .A(n4280), .B(B_REG_SCAN_IN), .ZN(
        n4281) );
  OAI21_X1 U4968 ( .B1(n4283), .B2(n4282), .A(n4281), .ZN(U3239) );
  MUX2_X1 U4969 ( .A(DATAO_REG_29__SCAN_IN), .B(n4284), .S(U4043), .Z(U3579)
         );
  MUX2_X1 U4970 ( .A(DATAO_REG_26__SCAN_IN), .B(n4285), .S(U4043), .Z(U3576)
         );
  MUX2_X1 U4971 ( .A(DATAO_REG_25__SCAN_IN), .B(n4479), .S(U4043), .Z(U3575)
         );
  MUX2_X1 U4972 ( .A(DATAO_REG_24__SCAN_IN), .B(n4457), .S(U4043), .Z(U3574)
         );
  MUX2_X1 U4973 ( .A(DATAO_REG_21__SCAN_IN), .B(n4553), .S(U4043), .Z(U3571)
         );
  MUX2_X1 U4974 ( .A(DATAO_REG_17__SCAN_IN), .B(n4624), .S(U4043), .Z(U3567)
         );
  MUX2_X1 U4975 ( .A(DATAO_REG_14__SCAN_IN), .B(n4286), .S(U4043), .Z(U3564)
         );
  MUX2_X1 U4976 ( .A(DATAO_REG_12__SCAN_IN), .B(n4287), .S(U4043), .Z(U3562)
         );
  MUX2_X1 U4977 ( .A(DATAO_REG_11__SCAN_IN), .B(n4288), .S(U4043), .Z(U3561)
         );
  MUX2_X1 U4978 ( .A(DATAO_REG_10__SCAN_IN), .B(n4289), .S(U4043), .Z(U3560)
         );
  MUX2_X1 U4979 ( .A(DATAO_REG_7__SCAN_IN), .B(n4290), .S(U4043), .Z(U3557) );
  MUX2_X1 U4980 ( .A(DATAO_REG_6__SCAN_IN), .B(n4291), .S(U4043), .Z(U3556) );
  MUX2_X1 U4981 ( .A(DATAO_REG_1__SCAN_IN), .B(n2990), .S(U4043), .Z(U3551) );
  MUX2_X1 U4982 ( .A(DATAO_REG_0__SCAN_IN), .B(n2991), .S(U4043), .Z(U3550) );
  INV_X1 U4983 ( .A(n4292), .ZN(n4296) );
  MUX2_X1 U4984 ( .A(n4293), .B(REG1_REG_1__SCAN_IN), .S(n3383), .Z(n4295) );
  OAI211_X1 U4985 ( .C1(n4296), .C2(n4295), .A(n4877), .B(n4294), .ZN(n4303)
         );
  OAI211_X1 U4986 ( .C1(n4298), .C2(n4308), .A(n4893), .B(n4297), .ZN(n4302)
         );
  AOI22_X1 U4987 ( .A1(n4883), .A2(ADDR_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(U3149), .ZN(n4301) );
  NAND2_X1 U4988 ( .A1(n4863), .A2(n4299), .ZN(n4300) );
  NAND4_X1 U4989 ( .A1(n4303), .A2(n4302), .A3(n4301), .A4(n4300), .ZN(U3241)
         );
  NAND3_X1 U4990 ( .A1(n4304), .A2(n4307), .A3(n4305), .ZN(n4312) );
  INV_X1 U4991 ( .A(REG2_REG_0__SCAN_IN), .ZN(n4906) );
  OR2_X1 U4992 ( .A1(n4305), .A2(REG2_REG_0__SCAN_IN), .ZN(n4306) );
  NAND2_X1 U4993 ( .A1(n4307), .A2(n4306), .ZN(n4822) );
  NAND2_X1 U4994 ( .A1(n4822), .A2(n2443), .ZN(n4311) );
  NAND2_X1 U4995 ( .A1(n4309), .A2(n4308), .ZN(n4310) );
  NAND4_X1 U4996 ( .A1(n4312), .A2(U4043), .A3(n4311), .A4(n4310), .ZN(n4839)
         );
  AOI22_X1 U4997 ( .A1(ADDR_REG_2__SCAN_IN), .A2(n4883), .B1(
        REG3_REG_2__SCAN_IN), .B2(U3149), .ZN(n4322) );
  INV_X1 U4998 ( .A(n3386), .ZN(n4316) );
  XOR2_X1 U4999 ( .A(n4314), .B(n4313), .Z(n4315) );
  AOI22_X1 U5000 ( .A1(n4316), .A2(n4863), .B1(n4877), .B2(n4315), .ZN(n4321)
         );
  OAI211_X1 U5001 ( .C1(n4319), .C2(n4318), .A(n4893), .B(n4317), .ZN(n4320)
         );
  NAND4_X1 U5002 ( .A1(n4839), .A2(n4322), .A3(n4321), .A4(n4320), .ZN(U3242)
         );
  INV_X1 U5003 ( .A(n4323), .ZN(n4325) );
  OAI22_X2 U5004 ( .A1(n4326), .A2(n3332), .B1(n4325), .B2(n4324), .ZN(n4848)
         );
  INV_X1 U5005 ( .A(REG2_REG_13__SCAN_IN), .ZN(n4845) );
  NAND2_X1 U5006 ( .A1(n4845), .A2(n4932), .ZN(n4327) );
  OAI211_X1 U5007 ( .C1(n4328), .C2(REG2_REG_14__SCAN_IN), .A(n4352), .B(n4893), .ZN(n4338) );
  AOI21_X1 U5008 ( .B1(n4883), .B2(ADDR_REG_14__SCAN_IN), .A(n4329), .ZN(n4337) );
  NAND2_X1 U5009 ( .A1(n4330), .A2(n4810), .ZN(n4331) );
  AOI22_X1 U5010 ( .A1(REG1_REG_13__SCAN_IN), .A2(n4932), .B1(n4846), .B2(
        n4740), .ZN(n4842) );
  OAI211_X1 U5011 ( .C1(n4334), .C2(REG1_REG_14__SCAN_IN), .A(n4340), .B(n4877), .ZN(n4336) );
  NAND2_X1 U5012 ( .A1(n4863), .A2(n4809), .ZN(n4335) );
  NAND4_X1 U5013 ( .A1(n4338), .A2(n4337), .A3(n4336), .A4(n4335), .ZN(U3254)
         );
  XNOR2_X1 U5014 ( .A(n4368), .B(n4724), .ZN(n4347) );
  INV_X1 U5015 ( .A(n4862), .ZN(n4930) );
  INV_X1 U5016 ( .A(REG1_REG_15__SCAN_IN), .ZN(n4341) );
  AOI22_X1 U5017 ( .A1(REG1_REG_15__SCAN_IN), .A2(n4930), .B1(n4862), .B2(
        n4341), .ZN(n4854) );
  INV_X1 U5018 ( .A(n4854), .ZN(n4342) );
  NAND2_X1 U5019 ( .A1(n2177), .A2(n4928), .ZN(n4345) );
  OAI21_X1 U5020 ( .B1(n4347), .B2(n4346), .A(n4363), .ZN(n4348) );
  AOI22_X1 U5021 ( .A1(n4368), .A2(n4863), .B1(n4877), .B2(n4348), .ZN(n4361)
         );
  XOR2_X1 U5022 ( .A(REG2_REG_17__SCAN_IN), .B(n4368), .Z(n4356) );
  INV_X1 U5023 ( .A(n4349), .ZN(n4350) );
  NAND2_X1 U5024 ( .A1(n4350), .A2(n4809), .ZN(n4351) );
  AOI22_X1 U5025 ( .A1(REG2_REG_15__SCAN_IN), .A2(n4930), .B1(n4862), .B2(
        n4649), .ZN(n4858) );
  NOR2_X2 U5026 ( .A1(n4857), .A2(n2413), .ZN(n4353) );
  NAND2_X1 U5027 ( .A1(n4353), .A2(n4928), .ZN(n4354) );
  INV_X1 U5028 ( .A(REG2_REG_16__SCAN_IN), .ZN(n4873) );
  NAND2_X1 U5029 ( .A1(n4354), .A2(n4872), .ZN(n4355) );
  OAI21_X1 U5030 ( .B1(n4356), .B2(n4355), .A(n4370), .ZN(n4357) );
  NAND2_X1 U5031 ( .A1(n4893), .A2(n4357), .ZN(n4359) );
  NAND2_X1 U5032 ( .A1(n4883), .A2(ADDR_REG_17__SCAN_IN), .ZN(n4358) );
  NAND4_X1 U5033 ( .A1(n4361), .A2(n4360), .A3(n4359), .A4(n4358), .ZN(U3257)
         );
  OR2_X1 U5034 ( .A1(n4368), .A2(REG1_REG_17__SCAN_IN), .ZN(n4362) );
  AOI22_X1 U5035 ( .A1(REG1_REG_18__SCAN_IN), .A2(n4926), .B1(n4367), .B2(
        n4364), .ZN(n4881) );
  XNOR2_X1 U5036 ( .A(n4376), .B(n4716), .ZN(n4365) );
  XNOR2_X1 U5037 ( .A(n4366), .B(n4365), .ZN(n4380) );
  NAND2_X1 U5038 ( .A1(REG2_REG_18__SCAN_IN), .A2(n4367), .ZN(n4371) );
  OAI21_X1 U5039 ( .B1(REG2_REG_18__SCAN_IN), .B2(n4367), .A(n4371), .ZN(n4891) );
  OR2_X1 U5040 ( .A1(n4368), .A2(REG2_REG_17__SCAN_IN), .ZN(n4369) );
  MUX2_X1 U5041 ( .A(n3126), .B(REG2_REG_19__SCAN_IN), .S(n4376), .Z(n4372) );
  XNOR2_X1 U5042 ( .A(n4373), .B(n4372), .ZN(n4378) );
  NAND2_X1 U5043 ( .A1(n4883), .A2(ADDR_REG_19__SCAN_IN), .ZN(n4374) );
  OAI211_X1 U5044 ( .C1(n4896), .C2(n4376), .A(n4375), .B(n4374), .ZN(n4377)
         );
  OAI21_X1 U5045 ( .B1(n4380), .B2(n4880), .A(n4379), .ZN(U3259) );
  NAND2_X1 U5046 ( .A1(n3499), .A2(n4669), .ZN(n4382) );
  NAND2_X1 U5047 ( .A1(n4908), .A2(REG2_REG_31__SCAN_IN), .ZN(n4381) );
  OAI211_X1 U5048 ( .C1(n4671), .C2(n4639), .A(n4382), .B(n4381), .ZN(U3260)
         );
  OAI21_X1 U5049 ( .B1(n4393), .B2(n4385), .A(n4383), .ZN(n4751) );
  OAI21_X1 U5050 ( .B1(n4385), .B2(n4627), .A(n4384), .ZN(n4748) );
  NOR2_X1 U5051 ( .A1(n3499), .A2(n4386), .ZN(n4387) );
  AOI21_X1 U5052 ( .B1(n3499), .B2(n4748), .A(n4387), .ZN(n4388) );
  OAI21_X1 U5053 ( .B1(n4751), .B2(n4639), .A(n4388), .ZN(U3261) );
  NAND2_X1 U5054 ( .A1(n4430), .A2(n4391), .ZN(n4678) );
  NAND2_X1 U5055 ( .A1(n4679), .A2(n4678), .ZN(n4392) );
  XNOR2_X1 U5056 ( .A(n4392), .B(n4677), .ZN(n4409) );
  AOI21_X1 U5057 ( .B1(n4399), .B2(n4394), .A(n4393), .ZN(n4680) );
  AOI22_X1 U5058 ( .A1(n4680), .A2(n4664), .B1(REG2_REG_29__SCAN_IN), .B2(
        n4908), .ZN(n4408) );
  INV_X1 U5059 ( .A(n4395), .ZN(n4397) );
  NAND2_X1 U5060 ( .A1(n4430), .A2(n4622), .ZN(n4403) );
  AOI22_X1 U5061 ( .A1(n4401), .A2(n4400), .B1(n4661), .B2(n4399), .ZN(n4402)
         );
  NOR2_X1 U5062 ( .A1(n4405), .A2(n4647), .ZN(n4406) );
  OAI21_X1 U5063 ( .B1(n4675), .B2(n4406), .A(n4485), .ZN(n4407) );
  OAI211_X1 U5064 ( .C1(n4409), .C2(n4666), .A(n4408), .B(n4407), .ZN(U3354)
         );
  INV_X1 U5065 ( .A(n4410), .ZN(n4418) );
  NOR2_X1 U5066 ( .A1(n4411), .A2(n4639), .ZN(n4415) );
  INV_X1 U5067 ( .A(REG2_REG_28__SCAN_IN), .ZN(n4412) );
  OAI22_X1 U5068 ( .A1(n4413), .A2(n4647), .B1(n4412), .B2(n4485), .ZN(n4414)
         );
  AOI211_X1 U5069 ( .C1(n4416), .C2(n4485), .A(n4415), .B(n4414), .ZN(n4417)
         );
  OAI21_X1 U5070 ( .B1(n4418), .B2(n4666), .A(n4417), .ZN(U3262) );
  XNOR2_X1 U5071 ( .A(n4419), .B(n4426), .ZN(n4685) );
  AOI21_X1 U5072 ( .B1(n4420), .B2(n2159), .A(n3074), .ZN(n4683) );
  INV_X1 U5073 ( .A(n4421), .ZN(n4423) );
  OAI22_X1 U5074 ( .A1(n4423), .A2(n4647), .B1(n4422), .B2(n4485), .ZN(n4424)
         );
  AOI21_X1 U5075 ( .B1(n4683), .B2(n4664), .A(n4424), .ZN(n4434) );
  XNOR2_X1 U5076 ( .A(n4425), .B(n4426), .ZN(n4427) );
  NAND2_X1 U5077 ( .A1(n4427), .A2(n4898), .ZN(n4432) );
  OAI22_X1 U5078 ( .A1(n4459), .A2(n4650), .B1(n4428), .B2(n4627), .ZN(n4429)
         );
  AOI21_X1 U5079 ( .B1(n4430), .B2(n4623), .A(n4429), .ZN(n4431) );
  NAND2_X1 U5080 ( .A1(n4432), .A2(n4431), .ZN(n4682) );
  NAND2_X1 U5081 ( .A1(n4682), .A2(n4485), .ZN(n4433) );
  OAI211_X1 U5082 ( .C1(n4685), .C2(n4666), .A(n4434), .B(n4433), .ZN(U3263)
         );
  XOR2_X1 U5083 ( .A(n4438), .B(n4435), .Z(n4687) );
  INV_X1 U5084 ( .A(n4687), .ZN(n4452) );
  NAND2_X1 U5085 ( .A1(n4437), .A2(n4436), .ZN(n4439) );
  XNOR2_X1 U5086 ( .A(n4439), .B(n4438), .ZN(n4445) );
  OAI22_X1 U5087 ( .A1(n4441), .A2(n4650), .B1(n4440), .B2(n4627), .ZN(n4442)
         );
  AOI21_X1 U5088 ( .B1(n4623), .B2(n4443), .A(n4442), .ZN(n4444) );
  OAI21_X1 U5089 ( .B1(n4445), .B2(n4655), .A(n4444), .ZN(n4686) );
  NAND2_X1 U5090 ( .A1(n2166), .A2(n4446), .ZN(n4447) );
  NAND2_X1 U5091 ( .A1(n2159), .A2(n4447), .ZN(n4757) );
  NOR2_X1 U5092 ( .A1(n4757), .A2(n4639), .ZN(n4450) );
  OAI22_X1 U5093 ( .A1(n4448), .A2(n4647), .B1(n3186), .B2(n4485), .ZN(n4449)
         );
  AOI211_X1 U5094 ( .C1(n4686), .C2(n4485), .A(n4450), .B(n4449), .ZN(n4451)
         );
  OAI21_X1 U5095 ( .B1(n4452), .B2(n4666), .A(n4451), .ZN(U3264) );
  XOR2_X1 U5096 ( .A(n4455), .B(n4453), .Z(n4691) );
  XNOR2_X1 U5097 ( .A(n4454), .B(n4455), .ZN(n4461) );
  AOI22_X1 U5098 ( .A1(n4457), .A2(n4622), .B1(n4456), .B2(n4661), .ZN(n4458)
         );
  OAI21_X1 U5099 ( .B1(n4459), .B2(n4901), .A(n4458), .ZN(n4460) );
  AOI21_X1 U5100 ( .B1(n4461), .B2(n4898), .A(n4460), .ZN(n4690) );
  INV_X1 U5101 ( .A(n4690), .ZN(n4468) );
  INV_X1 U5102 ( .A(n4483), .ZN(n4464) );
  OAI21_X1 U5103 ( .B1(n4464), .B2(n4463), .A(n2166), .ZN(n4761) );
  AOI22_X1 U5104 ( .A1(n4465), .A2(n4903), .B1(REG2_REG_25__SCAN_IN), .B2(
        n4908), .ZN(n4466) );
  OAI21_X1 U5105 ( .B1(n4761), .B2(n4639), .A(n4466), .ZN(n4467) );
  AOI21_X1 U5106 ( .B1(n4468), .B2(n4485), .A(n4467), .ZN(n4469) );
  OAI21_X1 U5107 ( .B1(n4691), .B2(n4666), .A(n4469), .ZN(U3265) );
  XNOR2_X1 U5108 ( .A(n4470), .B(n4477), .ZN(n4695) );
  INV_X1 U5109 ( .A(n4695), .ZN(n4491) );
  AOI21_X1 U5110 ( .B1(n4471), .B2(n4493), .A(n4472), .ZN(n4475) );
  INV_X1 U5111 ( .A(n4473), .ZN(n4474) );
  NOR2_X1 U5112 ( .A1(n4475), .A2(n4474), .ZN(n4476) );
  XOR2_X1 U5113 ( .A(n4477), .B(n4476), .Z(n4481) );
  OAI22_X1 U5114 ( .A1(n4517), .A2(n4650), .B1(n4484), .B2(n4627), .ZN(n4478)
         );
  AOI21_X1 U5115 ( .B1(n4479), .B2(n4623), .A(n4478), .ZN(n4480) );
  OAI21_X1 U5116 ( .B1(n4481), .B2(n4655), .A(n4480), .ZN(n4694) );
  OAI21_X1 U5117 ( .B1(n4482), .B2(n4484), .A(n4483), .ZN(n4765) );
  NOR2_X1 U5118 ( .A1(n4765), .A2(n4639), .ZN(n4489) );
  INV_X1 U5119 ( .A(REG2_REG_24__SCAN_IN), .ZN(n4486) );
  OAI22_X1 U5120 ( .A1(n4487), .A2(n4647), .B1(n4486), .B2(n4485), .ZN(n4488)
         );
  AOI211_X1 U5121 ( .C1(n4694), .C2(n4485), .A(n4489), .B(n4488), .ZN(n4490)
         );
  OAI21_X1 U5122 ( .B1(n4491), .B2(n4666), .A(n4490), .ZN(U3266) );
  XOR2_X1 U5123 ( .A(n4496), .B(n4492), .Z(n4699) );
  INV_X1 U5124 ( .A(n4699), .ZN(n4509) );
  NOR2_X1 U5125 ( .A1(n4471), .A2(n4511), .ZN(n4512) );
  INV_X1 U5126 ( .A(n4493), .ZN(n4494) );
  NOR2_X1 U5127 ( .A1(n4512), .A2(n4494), .ZN(n4495) );
  XOR2_X1 U5128 ( .A(n4496), .B(n4495), .Z(n4500) );
  OAI22_X1 U5129 ( .A1(n4497), .A2(n4901), .B1(n4627), .B2(n4503), .ZN(n4498)
         );
  AOI21_X1 U5130 ( .B1(n4622), .B2(n4532), .A(n4498), .ZN(n4499) );
  OAI21_X1 U5131 ( .B1(n4500), .B2(n4655), .A(n4499), .ZN(n4698) );
  INV_X1 U5132 ( .A(n4482), .ZN(n4502) );
  OAI21_X1 U5133 ( .B1(n3072), .B2(n4503), .A(n4502), .ZN(n4769) );
  INV_X1 U5134 ( .A(n4504), .ZN(n4505) );
  AOI22_X1 U5135 ( .A1(n4505), .A2(n4903), .B1(REG2_REG_23__SCAN_IN), .B2(
        n4908), .ZN(n4506) );
  OAI21_X1 U5136 ( .B1(n4769), .B2(n4639), .A(n4506), .ZN(n4507) );
  AOI21_X1 U5137 ( .B1(n4698), .B2(n4485), .A(n4507), .ZN(n4508) );
  OAI21_X1 U5138 ( .B1(n4509), .B2(n4666), .A(n4508), .ZN(U3267) );
  OAI21_X1 U5139 ( .B1(n2175), .B2(n4511), .A(n4510), .ZN(n4705) );
  AND2_X1 U5140 ( .A1(n4471), .A2(n4511), .ZN(n4513) );
  OR2_X1 U5141 ( .A1(n4513), .A2(n4512), .ZN(n4519) );
  NOR2_X1 U5142 ( .A1(n4627), .A2(n4514), .ZN(n4515) );
  AOI21_X1 U5143 ( .B1(n4553), .B2(n4622), .A(n4515), .ZN(n4516) );
  OAI21_X1 U5144 ( .B1(n4517), .B2(n4901), .A(n4516), .ZN(n4518) );
  AOI21_X1 U5145 ( .B1(n4519), .B2(n4898), .A(n4518), .ZN(n4704) );
  AOI22_X1 U5146 ( .A1(n4520), .A2(n4903), .B1(REG2_REG_22__SCAN_IN), .B2(
        n4908), .ZN(n4523) );
  NAND2_X1 U5147 ( .A1(n4535), .A2(n4521), .ZN(n4702) );
  NAND3_X1 U5148 ( .A1(n4501), .A2(n4664), .A3(n4702), .ZN(n4522) );
  OAI211_X1 U5149 ( .C1(n4704), .C2(n4908), .A(n4523), .B(n4522), .ZN(n4524)
         );
  INV_X1 U5150 ( .A(n4524), .ZN(n4525) );
  OAI21_X1 U5151 ( .B1(n4705), .B2(n4666), .A(n4525), .ZN(U3268) );
  XOR2_X1 U5152 ( .A(n4528), .B(n4526), .Z(n4707) );
  INV_X1 U5153 ( .A(n4707), .ZN(n4542) );
  XNOR2_X1 U5154 ( .A(n4527), .B(n4528), .ZN(n4529) );
  NAND2_X1 U5155 ( .A1(n4529), .A2(n4898), .ZN(n4534) );
  NAND2_X1 U5156 ( .A1(n4574), .A2(n4622), .ZN(n4530) );
  OAI21_X1 U5157 ( .B1(n4627), .B2(n4536), .A(n4530), .ZN(n4531) );
  AOI21_X1 U5158 ( .B1(n4532), .B2(n4623), .A(n4531), .ZN(n4533) );
  NAND2_X1 U5159 ( .A1(n4534), .A2(n4533), .ZN(n4706) );
  INV_X1 U5160 ( .A(n4557), .ZN(n4537) );
  OAI21_X1 U5161 ( .B1(n4537), .B2(n4536), .A(n4535), .ZN(n4774) );
  AOI22_X1 U5162 ( .A1(n4538), .A2(n4903), .B1(n4908), .B2(
        REG2_REG_21__SCAN_IN), .ZN(n4539) );
  OAI21_X1 U5163 ( .B1(n4774), .B2(n4639), .A(n4539), .ZN(n4540) );
  AOI21_X1 U5164 ( .B1(n4706), .B2(n4485), .A(n4540), .ZN(n4541) );
  OAI21_X1 U5165 ( .B1(n4542), .B2(n4666), .A(n4541), .ZN(U3269) );
  XNOR2_X1 U5166 ( .A(n4543), .B(n4550), .ZN(n4711) );
  INV_X1 U5167 ( .A(n4711), .ZN(n4564) );
  OR2_X1 U5168 ( .A1(n4606), .A2(n4546), .ZN(n4549) );
  INV_X1 U5169 ( .A(n4547), .ZN(n4548) );
  NAND2_X1 U5170 ( .A1(n4549), .A2(n4548), .ZN(n4551) );
  XNOR2_X1 U5171 ( .A(n4551), .B(n4550), .ZN(n4555) );
  OAI22_X1 U5172 ( .A1(n4591), .A2(n4650), .B1(n4558), .B2(n4627), .ZN(n4552)
         );
  AOI21_X1 U5173 ( .B1(n4553), .B2(n4623), .A(n4552), .ZN(n4554) );
  OAI21_X1 U5174 ( .B1(n4555), .B2(n4655), .A(n4554), .ZN(n4710) );
  INV_X1 U5175 ( .A(n4556), .ZN(n4559) );
  OAI21_X1 U5176 ( .B1(n4559), .B2(n4558), .A(n4557), .ZN(n4778) );
  AOI22_X1 U5177 ( .A1(n4908), .A2(REG2_REG_20__SCAN_IN), .B1(n4560), .B2(
        n4903), .ZN(n4561) );
  OAI21_X1 U5178 ( .B1(n4778), .B2(n4639), .A(n4561), .ZN(n4562) );
  AOI21_X1 U5179 ( .B1(n4710), .B2(n4485), .A(n4562), .ZN(n4563) );
  OAI21_X1 U5180 ( .B1(n4564), .B2(n4666), .A(n4563), .ZN(U3270) );
  NAND2_X1 U5181 ( .A1(n4567), .A2(n4566), .ZN(n4588) );
  INV_X1 U5182 ( .A(n4568), .ZN(n4570) );
  OAI21_X1 U5183 ( .B1(n4588), .B2(n4570), .A(n4569), .ZN(n4571) );
  XNOR2_X1 U5184 ( .A(n4571), .B(n4577), .ZN(n4576) );
  OAI22_X1 U5185 ( .A1(n4572), .A2(n4650), .B1(n4627), .B2(n4579), .ZN(n4573)
         );
  AOI21_X1 U5186 ( .B1(n4623), .B2(n4574), .A(n4573), .ZN(n4575) );
  OAI21_X1 U5187 ( .B1(n4576), .B2(n4655), .A(n4575), .ZN(n4714) );
  INV_X1 U5188 ( .A(n4714), .ZN(n4586) );
  XNOR2_X1 U5189 ( .A(n4578), .B(n4577), .ZN(n4715) );
  OR2_X1 U5190 ( .A1(n4580), .A2(n4579), .ZN(n4581) );
  NAND2_X1 U5191 ( .A1(n4556), .A2(n4581), .ZN(n4782) );
  AOI22_X1 U5192 ( .A1(n4908), .A2(REG2_REG_19__SCAN_IN), .B1(n4582), .B2(
        n4903), .ZN(n4583) );
  OAI21_X1 U5193 ( .B1(n4782), .B2(n4639), .A(n4583), .ZN(n4584) );
  AOI21_X1 U5194 ( .B1(n4715), .B2(n4641), .A(n4584), .ZN(n4585) );
  OAI21_X1 U5195 ( .B1(n4908), .B2(n4586), .A(n4585), .ZN(U3271) );
  INV_X1 U5196 ( .A(n4601), .ZN(n4587) );
  XNOR2_X1 U5197 ( .A(n4588), .B(n4587), .ZN(n4593) );
  AOI22_X1 U5198 ( .A1(n4624), .A2(n4622), .B1(n4589), .B2(n4661), .ZN(n4590)
         );
  OAI21_X1 U5199 ( .B1(n4591), .B2(n4901), .A(n4590), .ZN(n4592) );
  AOI21_X1 U5200 ( .B1(n4593), .B2(n4898), .A(n4592), .ZN(n4721) );
  XNOR2_X1 U5201 ( .A(n4594), .B(n4595), .ZN(n4596) );
  AND2_X1 U5202 ( .A1(n4596), .A2(n4943), .ZN(n4718) );
  INV_X1 U5203 ( .A(REG2_REG_18__SCAN_IN), .ZN(n4598) );
  OAI22_X1 U5204 ( .A1(n3499), .A2(n4598), .B1(n4597), .B2(n4647), .ZN(n4599)
         );
  AOI21_X1 U5205 ( .B1(n4718), .B2(n4600), .A(n4599), .ZN(n4605) );
  NOR2_X1 U5206 ( .A1(n2173), .A2(n4601), .ZN(n4602) );
  OR2_X1 U5207 ( .A1(n4603), .A2(n4602), .ZN(n4719) );
  NAND2_X1 U5208 ( .A1(n4719), .A2(n4641), .ZN(n4604) );
  OAI211_X1 U5209 ( .C1(n4721), .C2(n4908), .A(n4605), .B(n4604), .ZN(U3272)
         );
  XNOR2_X1 U5210 ( .A(n4606), .B(n4611), .ZN(n4610) );
  OAI22_X1 U5211 ( .A1(n4652), .A2(n4650), .B1(n4627), .B2(n4613), .ZN(n4607)
         );
  AOI21_X1 U5212 ( .B1(n4623), .B2(n4608), .A(n4607), .ZN(n4609) );
  OAI21_X1 U5213 ( .B1(n4610), .B2(n4655), .A(n4609), .ZN(n4722) );
  INV_X1 U5214 ( .A(n4722), .ZN(n4619) );
  XNOR2_X1 U5215 ( .A(n4612), .B(n4611), .ZN(n4723) );
  OR2_X1 U5216 ( .A1(n4635), .A2(n4613), .ZN(n4614) );
  NAND2_X1 U5217 ( .A1(n4594), .A2(n4614), .ZN(n4787) );
  AOI22_X1 U5218 ( .A1(n4908), .A2(REG2_REG_17__SCAN_IN), .B1(n4615), .B2(
        n4903), .ZN(n4616) );
  OAI21_X1 U5219 ( .B1(n4787), .B2(n4639), .A(n4616), .ZN(n4617) );
  AOI21_X1 U5220 ( .B1(n4723), .B2(n4641), .A(n4617), .ZN(n4618) );
  OAI21_X1 U5221 ( .B1(n4619), .B2(n4908), .A(n4618), .ZN(U3273) );
  OAI211_X1 U5222 ( .C1(n4620), .C2(n4632), .A(n4544), .B(n4898), .ZN(n4626)
         );
  AOI22_X1 U5223 ( .A1(n4624), .A2(n4623), .B1(n4622), .B2(n4621), .ZN(n4625)
         );
  OAI211_X1 U5224 ( .C1(n4627), .C2(n4633), .A(n4626), .B(n4625), .ZN(n4628)
         );
  INV_X1 U5225 ( .A(n4628), .ZN(n4727) );
  INV_X1 U5226 ( .A(n4630), .ZN(n4631) );
  AOI21_X1 U5227 ( .B1(n4632), .B2(n4629), .A(n4631), .ZN(n4726) );
  NOR2_X1 U5228 ( .A1(n2406), .A2(n4633), .ZN(n4634) );
  OR2_X1 U5229 ( .A1(n4635), .A2(n4634), .ZN(n4729) );
  INV_X1 U5230 ( .A(n4636), .ZN(n4637) );
  AOI22_X1 U5231 ( .A1(n4908), .A2(REG2_REG_16__SCAN_IN), .B1(n4637), .B2(
        n4903), .ZN(n4638) );
  OAI21_X1 U5232 ( .B1(n4729), .B2(n4639), .A(n4638), .ZN(n4640) );
  AOI21_X1 U5233 ( .B1(n4726), .B2(n4641), .A(n4640), .ZN(n4642) );
  OAI21_X1 U5234 ( .B1(n4908), .B2(n4727), .A(n4642), .ZN(U3274) );
  XNOR2_X1 U5235 ( .A(n4644), .B(n4643), .ZN(n4733) );
  XNOR2_X1 U5236 ( .A(n4646), .B(n4645), .ZN(n4730) );
  OAI22_X1 U5237 ( .A1(n3499), .A2(n4649), .B1(n4648), .B2(n4647), .ZN(n4663)
         );
  OAI22_X1 U5238 ( .A1(n4652), .A2(n4901), .B1(n4651), .B2(n4650), .ZN(n4659)
         );
  INV_X1 U5239 ( .A(n4653), .ZN(n4654) );
  AOI211_X1 U5240 ( .C1(n4657), .C2(n4656), .A(n4655), .B(n4654), .ZN(n4658)
         );
  AOI211_X1 U5241 ( .C1(n4661), .C2(n4660), .A(n4659), .B(n4658), .ZN(n4732)
         );
  NOR2_X1 U5242 ( .A1(n4732), .A2(n4908), .ZN(n4662) );
  AOI211_X1 U5243 ( .C1(n4664), .C2(n4730), .A(n4663), .B(n4662), .ZN(n4665)
         );
  OAI21_X1 U5244 ( .B1(n4733), .B2(n4666), .A(n4665), .ZN(U3275) );
  NOR2_X1 U5245 ( .A1(n4975), .A2(n4667), .ZN(n4668) );
  AOI21_X1 U5246 ( .B1(n4975), .B2(n4669), .A(n4668), .ZN(n4670) );
  OAI21_X1 U5247 ( .B1(n4671), .B2(n4747), .A(n4670), .ZN(U3549) );
  NAND2_X1 U5248 ( .A1(n4975), .A2(n4748), .ZN(n4673) );
  NAND2_X1 U5249 ( .A1(n4976), .A2(REG1_REG_30__SCAN_IN), .ZN(n4672) );
  OAI211_X1 U5250 ( .C1(n4751), .C2(n4747), .A(n4673), .B(n4672), .ZN(U3548)
         );
  INV_X1 U5251 ( .A(n4744), .ZN(n4959) );
  NAND2_X1 U5252 ( .A1(n4679), .A2(n2409), .ZN(n4681) );
  AOI21_X1 U5253 ( .B1(n4943), .B2(n4683), .A(n4682), .ZN(n4684) );
  OAI21_X1 U5254 ( .B1(n4685), .B2(n4959), .A(n4684), .ZN(n4753) );
  MUX2_X1 U5255 ( .A(REG1_REG_27__SCAN_IN), .B(n4753), .S(n4975), .Z(U3545) );
  AOI21_X1 U5256 ( .B1(n4687), .B2(n4744), .A(n4686), .ZN(n4754) );
  MUX2_X1 U5257 ( .A(n4688), .B(n4754), .S(n4975), .Z(n4689) );
  OAI21_X1 U5258 ( .B1(n4747), .B2(n4757), .A(n4689), .ZN(U3544) );
  OAI21_X1 U5259 ( .B1(n4691), .B2(n4959), .A(n4690), .ZN(n4758) );
  MUX2_X1 U5260 ( .A(REG1_REG_25__SCAN_IN), .B(n4758), .S(n4975), .Z(n4692) );
  INV_X1 U5261 ( .A(n4692), .ZN(n4693) );
  OAI21_X1 U5262 ( .B1(n4747), .B2(n4761), .A(n4693), .ZN(U3543) );
  AOI21_X1 U5263 ( .B1(n4695), .B2(n4744), .A(n4694), .ZN(n4762) );
  MUX2_X1 U5264 ( .A(n4696), .B(n4762), .S(n4975), .Z(n4697) );
  OAI21_X1 U5265 ( .B1(n4747), .B2(n4765), .A(n4697), .ZN(U3542) );
  AOI21_X1 U5266 ( .B1(n4699), .B2(n4744), .A(n4698), .ZN(n4766) );
  MUX2_X1 U5267 ( .A(n4700), .B(n4766), .S(n4975), .Z(n4701) );
  OAI21_X1 U5268 ( .B1(n4747), .B2(n4769), .A(n4701), .ZN(U3541) );
  NAND3_X1 U5269 ( .A1(n4501), .A2(n4943), .A3(n4702), .ZN(n4703) );
  OAI211_X1 U5270 ( .C1(n4705), .C2(n4959), .A(n4704), .B(n4703), .ZN(n4770)
         );
  MUX2_X1 U5271 ( .A(REG1_REG_22__SCAN_IN), .B(n4770), .S(n4975), .Z(U3540) );
  AOI21_X1 U5272 ( .B1(n4707), .B2(n4744), .A(n4706), .ZN(n4771) );
  MUX2_X1 U5273 ( .A(n4708), .B(n4771), .S(n4975), .Z(n4709) );
  OAI21_X1 U5274 ( .B1(n4747), .B2(n4774), .A(n4709), .ZN(U3539) );
  INV_X1 U5275 ( .A(REG1_REG_20__SCAN_IN), .ZN(n4712) );
  AOI21_X1 U5276 ( .B1(n4711), .B2(n4744), .A(n4710), .ZN(n4775) );
  MUX2_X1 U5277 ( .A(n4712), .B(n4775), .S(n4975), .Z(n4713) );
  OAI21_X1 U5278 ( .B1(n4747), .B2(n4778), .A(n4713), .ZN(U3538) );
  AOI21_X1 U5279 ( .B1(n4715), .B2(n4744), .A(n4714), .ZN(n4779) );
  MUX2_X1 U5280 ( .A(n4716), .B(n4779), .S(n4975), .Z(n4717) );
  OAI21_X1 U5281 ( .B1(n4747), .B2(n4782), .A(n4717), .ZN(U3537) );
  AOI21_X1 U5282 ( .B1(n4719), .B2(n4744), .A(n4718), .ZN(n4720) );
  NAND2_X1 U5283 ( .A1(n4721), .A2(n4720), .ZN(n4783) );
  MUX2_X1 U5284 ( .A(REG1_REG_18__SCAN_IN), .B(n4783), .S(n4975), .Z(U3536) );
  AOI21_X1 U5285 ( .B1(n4723), .B2(n4744), .A(n4722), .ZN(n4784) );
  MUX2_X1 U5286 ( .A(n4724), .B(n4784), .S(n4975), .Z(n4725) );
  OAI21_X1 U5287 ( .B1(n4747), .B2(n4787), .A(n4725), .ZN(U3535) );
  NAND2_X1 U5288 ( .A1(n4726), .A2(n4744), .ZN(n4728) );
  OAI211_X1 U5289 ( .C1(n3076), .C2(n4729), .A(n4728), .B(n4727), .ZN(n4788)
         );
  MUX2_X1 U5290 ( .A(REG1_REG_16__SCAN_IN), .B(n4788), .S(n4975), .Z(U3534) );
  NAND2_X1 U5291 ( .A1(n4730), .A2(n4943), .ZN(n4731) );
  OAI211_X1 U5292 ( .C1(n4959), .C2(n4733), .A(n4732), .B(n4731), .ZN(n4789)
         );
  MUX2_X1 U5293 ( .A(REG1_REG_15__SCAN_IN), .B(n4789), .S(n4975), .Z(U3533) );
  AOI21_X1 U5294 ( .B1(n4744), .B2(n4735), .A(n4734), .ZN(n4790) );
  MUX2_X1 U5295 ( .A(n4736), .B(n4790), .S(n4975), .Z(n4737) );
  OAI21_X1 U5296 ( .B1(n4747), .B2(n4793), .A(n4737), .ZN(U3532) );
  AOI21_X1 U5297 ( .B1(n4951), .B2(n4739), .A(n4738), .ZN(n4794) );
  MUX2_X1 U5298 ( .A(n4740), .B(n4794), .S(n4975), .Z(n4741) );
  OAI21_X1 U5299 ( .B1(n4747), .B2(n4797), .A(n4741), .ZN(U3531) );
  AOI21_X1 U5300 ( .B1(n4744), .B2(n4743), .A(n4742), .ZN(n4799) );
  MUX2_X1 U5301 ( .A(n4745), .B(n4799), .S(n4975), .Z(n4746) );
  OAI21_X1 U5302 ( .B1(n4747), .B2(n4803), .A(n4746), .ZN(U3530) );
  NAND2_X1 U5303 ( .A1(n4798), .A2(n4748), .ZN(n4750) );
  NAND2_X1 U5304 ( .A1(n4965), .A2(REG0_REG_30__SCAN_IN), .ZN(n4749) );
  OAI211_X1 U5305 ( .C1(n4751), .C2(n4802), .A(n4750), .B(n4749), .ZN(U3516)
         );
  MUX2_X1 U5306 ( .A(REG0_REG_29__SCAN_IN), .B(n4752), .S(n4967), .Z(U3515) );
  MUX2_X1 U5307 ( .A(REG0_REG_27__SCAN_IN), .B(n4753), .S(n4798), .Z(U3513) );
  INV_X1 U5308 ( .A(REG0_REG_26__SCAN_IN), .ZN(n4755) );
  MUX2_X1 U5309 ( .A(n4755), .B(n4754), .S(n4967), .Z(n4756) );
  OAI21_X1 U5310 ( .B1(n4757), .B2(n4802), .A(n4756), .ZN(U3512) );
  MUX2_X1 U5311 ( .A(REG0_REG_25__SCAN_IN), .B(n4758), .S(n4798), .Z(n4759) );
  INV_X1 U5312 ( .A(n4759), .ZN(n4760) );
  OAI21_X1 U5313 ( .B1(n4761), .B2(n4802), .A(n4760), .ZN(U3511) );
  INV_X1 U5314 ( .A(REG0_REG_24__SCAN_IN), .ZN(n4763) );
  MUX2_X1 U5315 ( .A(n4763), .B(n4762), .S(n4967), .Z(n4764) );
  OAI21_X1 U5316 ( .B1(n4765), .B2(n4802), .A(n4764), .ZN(U3510) );
  INV_X1 U5317 ( .A(REG0_REG_23__SCAN_IN), .ZN(n4767) );
  MUX2_X1 U5318 ( .A(n4767), .B(n4766), .S(n4798), .Z(n4768) );
  OAI21_X1 U5319 ( .B1(n4769), .B2(n4802), .A(n4768), .ZN(U3509) );
  MUX2_X1 U5320 ( .A(REG0_REG_22__SCAN_IN), .B(n4770), .S(n4798), .Z(U3508) );
  INV_X1 U5321 ( .A(REG0_REG_21__SCAN_IN), .ZN(n4772) );
  MUX2_X1 U5322 ( .A(n4772), .B(n4771), .S(n4967), .Z(n4773) );
  OAI21_X1 U5323 ( .B1(n4774), .B2(n4802), .A(n4773), .ZN(U3507) );
  MUX2_X1 U5324 ( .A(n4776), .B(n4775), .S(n4967), .Z(n4777) );
  OAI21_X1 U5325 ( .B1(n4778), .B2(n4802), .A(n4777), .ZN(U3506) );
  INV_X1 U5326 ( .A(REG0_REG_19__SCAN_IN), .ZN(n4780) );
  MUX2_X1 U5327 ( .A(n4780), .B(n4779), .S(n4798), .Z(n4781) );
  OAI21_X1 U5328 ( .B1(n4782), .B2(n4802), .A(n4781), .ZN(U3505) );
  MUX2_X1 U5329 ( .A(REG0_REG_18__SCAN_IN), .B(n4783), .S(n4798), .Z(U3503) );
  INV_X1 U5330 ( .A(REG0_REG_17__SCAN_IN), .ZN(n4785) );
  MUX2_X1 U5331 ( .A(n4785), .B(n4784), .S(n4967), .Z(n4786) );
  OAI21_X1 U5332 ( .B1(n4787), .B2(n4802), .A(n4786), .ZN(U3501) );
  MUX2_X1 U5333 ( .A(REG0_REG_16__SCAN_IN), .B(n4788), .S(n4798), .Z(U3499) );
  MUX2_X1 U5334 ( .A(REG0_REG_15__SCAN_IN), .B(n4789), .S(n4798), .Z(U3497) );
  MUX2_X1 U5335 ( .A(n4791), .B(n4790), .S(n4967), .Z(n4792) );
  OAI21_X1 U5336 ( .B1(n4793), .B2(n4802), .A(n4792), .ZN(U3495) );
  MUX2_X1 U5337 ( .A(n4795), .B(n4794), .S(n4798), .Z(n4796) );
  OAI21_X1 U5338 ( .B1(n4797), .B2(n4802), .A(n4796), .ZN(U3493) );
  INV_X1 U5339 ( .A(REG0_REG_12__SCAN_IN), .ZN(n4800) );
  MUX2_X1 U5340 ( .A(n4800), .B(n4799), .S(n4798), .Z(n4801) );
  OAI21_X1 U5341 ( .B1(n4803), .B2(n4802), .A(n4801), .ZN(U3491) );
  MUX2_X1 U5342 ( .A(DATAI_29_), .B(n4804), .S(STATE_REG_SCAN_IN), .Z(U3323)
         );
  MUX2_X1 U5343 ( .A(DATAI_26_), .B(n4805), .S(STATE_REG_SCAN_IN), .Z(U3326)
         );
  MUX2_X1 U5344 ( .A(DATAI_24_), .B(n4806), .S(STATE_REG_SCAN_IN), .Z(U3328)
         );
  MUX2_X1 U5345 ( .A(n2468), .B(DATAI_22_), .S(U3149), .Z(U3330) );
  MUX2_X1 U5346 ( .A(DATAI_21_), .B(n2469), .S(STATE_REG_SCAN_IN), .Z(U3331)
         );
  MUX2_X1 U5347 ( .A(DATAI_20_), .B(n4807), .S(STATE_REG_SCAN_IN), .Z(U3332)
         );
  MUX2_X1 U5348 ( .A(n4808), .B(DATAI_19_), .S(U3149), .Z(U3333) );
  MUX2_X1 U5349 ( .A(n4809), .B(DATAI_14_), .S(U3149), .Z(U3338) );
  MUX2_X1 U5350 ( .A(n4810), .B(DATAI_12_), .S(U3149), .Z(U3340) );
  INV_X1 U5351 ( .A(n4811), .ZN(n4812) );
  MUX2_X1 U5352 ( .A(n4812), .B(DATAI_11_), .S(U3149), .Z(U3341) );
  MUX2_X1 U5353 ( .A(DATAI_9_), .B(n4813), .S(STATE_REG_SCAN_IN), .Z(U3343) );
  MUX2_X1 U5354 ( .A(DATAI_8_), .B(n4814), .S(STATE_REG_SCAN_IN), .Z(U3344) );
  MUX2_X1 U5355 ( .A(n4815), .B(DATAI_6_), .S(U3149), .Z(U3346) );
  MUX2_X1 U5356 ( .A(n4816), .B(DATAI_5_), .S(U3149), .Z(U3347) );
  MUX2_X1 U5357 ( .A(DATAI_3_), .B(n4817), .S(STATE_REG_SCAN_IN), .Z(U3349) );
  AOI22_X1 U5358 ( .A1(STATE_REG_SCAN_IN), .A2(n4819), .B1(n4818), .B2(U3149), 
        .ZN(U3324) );
  INV_X1 U5359 ( .A(n4822), .ZN(n4820) );
  OAI211_X1 U5360 ( .C1(REG1_REG_0__SCAN_IN), .C2(n4821), .A(n4823), .B(n4820), 
        .ZN(n4826) );
  AOI22_X1 U5361 ( .A1(n4823), .A2(n4822), .B1(n4877), .B2(n4968), .ZN(n4825)
         );
  AOI22_X1 U5362 ( .A1(ADDR_REG_0__SCAN_IN), .A2(n4883), .B1(
        REG3_REG_0__SCAN_IN), .B2(U3149), .ZN(n4824) );
  OAI221_X1 U5363 ( .B1(IR_REG_0__SCAN_IN), .B2(n4826), .C1(n2443), .C2(n4825), 
        .A(n4824), .ZN(U3240) );
  XNOR2_X1 U5364 ( .A(n4827), .B(n4828), .ZN(n4829) );
  NAND2_X1 U5365 ( .A1(n4893), .A2(n4829), .ZN(n4838) );
  XNOR2_X1 U5366 ( .A(n4831), .B(n4830), .ZN(n4832) );
  NAND2_X1 U5367 ( .A1(n4877), .A2(n4832), .ZN(n4837) );
  NAND2_X1 U5368 ( .A1(n4863), .A2(n4833), .ZN(n4836) );
  AOI21_X1 U5369 ( .B1(n4883), .B2(ADDR_REG_4__SCAN_IN), .A(n4834), .ZN(n4835)
         );
  AND4_X1 U5370 ( .A1(n4838), .A2(n4837), .A3(n4836), .A4(n4835), .ZN(n4840)
         );
  NAND2_X1 U5371 ( .A1(n4840), .A2(n4839), .ZN(U3244) );
  AOI211_X1 U5372 ( .C1(n2184), .C2(n4842), .A(n4841), .B(n4880), .ZN(n4843)
         );
  AOI211_X1 U5373 ( .C1(n4883), .C2(ADDR_REG_13__SCAN_IN), .A(n4844), .B(n4843), .ZN(n4851) );
  AOI22_X1 U5374 ( .A1(REG2_REG_13__SCAN_IN), .A2(n4846), .B1(n4932), .B2(
        n4845), .ZN(n4849) );
  AOI21_X1 U5375 ( .B1(n4849), .B2(n4848), .A(n4856), .ZN(n4847) );
  OAI21_X1 U5376 ( .B1(n4849), .B2(n4848), .A(n4847), .ZN(n4850) );
  OAI211_X1 U5377 ( .C1(n4896), .C2(n4932), .A(n4851), .B(n4850), .ZN(U3253)
         );
  INV_X1 U5378 ( .A(n4883), .ZN(n4867) );
  AOI211_X1 U5379 ( .C1(n4855), .C2(n4854), .A(n4853), .B(n4880), .ZN(n4861)
         );
  AOI211_X1 U5380 ( .C1(n4859), .C2(n4858), .A(n4857), .B(n4856), .ZN(n4860)
         );
  AOI211_X1 U5381 ( .C1(n4863), .C2(n4862), .A(n4861), .B(n4860), .ZN(n4865)
         );
  OAI211_X1 U5382 ( .C1(n4867), .C2(n4866), .A(n4865), .B(n4864), .ZN(U3255)
         );
  AOI21_X1 U5383 ( .B1(n4883), .B2(ADDR_REG_16__SCAN_IN), .A(n4868), .ZN(n4879) );
  OAI21_X1 U5384 ( .B1(n4871), .B2(n4870), .A(n4869), .ZN(n4876) );
  OAI21_X1 U5385 ( .B1(n4874), .B2(n4873), .A(n4872), .ZN(n4875) );
  AOI22_X1 U5386 ( .A1(n4877), .A2(n4876), .B1(n4893), .B2(n4875), .ZN(n4878)
         );
  OAI211_X1 U5387 ( .C1(n4928), .C2(n4896), .A(n4879), .B(n4878), .ZN(U3256)
         );
  NAND2_X1 U5388 ( .A1(n4883), .A2(ADDR_REG_18__SCAN_IN), .ZN(n4886) );
  INV_X1 U5389 ( .A(n4884), .ZN(n4885) );
  AOI21_X1 U5390 ( .B1(n4891), .B2(n4890), .A(n4889), .ZN(n4892) );
  NAND2_X1 U5391 ( .A1(n4893), .A2(n4892), .ZN(n4894) );
  OAI211_X1 U5392 ( .C1(n4896), .C2(n4926), .A(n4895), .B(n4894), .ZN(U3258)
         );
  NOR2_X1 U5393 ( .A1(n3636), .A2(n2948), .ZN(n4934) );
  INV_X1 U5394 ( .A(n4897), .ZN(n4935) );
  OAI21_X1 U5395 ( .B1(n4899), .B2(n4898), .A(n4935), .ZN(n4900) );
  OAI21_X1 U5396 ( .B1(n2989), .B2(n4901), .A(n4900), .ZN(n4933) );
  AOI21_X1 U5397 ( .B1(n4934), .B2(n4902), .A(n4933), .ZN(n4907) );
  AOI22_X1 U5398 ( .A1(n4904), .A2(n4935), .B1(REG3_REG_0__SCAN_IN), .B2(n4903), .ZN(n4905) );
  OAI221_X1 U5399 ( .B1(n4908), .B2(n4907), .C1(n3499), .C2(n4906), .A(n4905), 
        .ZN(U3290) );
  AND2_X1 U5400 ( .A1(D_REG_31__SCAN_IN), .A2(n4921), .ZN(U3291) );
  AND2_X1 U5401 ( .A1(D_REG_30__SCAN_IN), .A2(n4921), .ZN(U3292) );
  NOR2_X1 U5402 ( .A1(n4923), .A2(n4909), .ZN(U3293) );
  AND2_X1 U5403 ( .A1(D_REG_28__SCAN_IN), .A2(n4921), .ZN(U3294) );
  AND2_X1 U5404 ( .A1(D_REG_27__SCAN_IN), .A2(n4921), .ZN(U3295) );
  NOR2_X1 U5405 ( .A1(n4923), .A2(n4910), .ZN(U3296) );
  AND2_X1 U5406 ( .A1(D_REG_25__SCAN_IN), .A2(n4921), .ZN(U3297) );
  NOR2_X1 U5407 ( .A1(n4923), .A2(n4911), .ZN(U3298) );
  NOR2_X1 U5408 ( .A1(n4923), .A2(n4912), .ZN(U3299) );
  AND2_X1 U5409 ( .A1(D_REG_22__SCAN_IN), .A2(n4921), .ZN(U3300) );
  NOR2_X1 U5410 ( .A1(n4923), .A2(n4913), .ZN(U3301) );
  AND2_X1 U5411 ( .A1(D_REG_20__SCAN_IN), .A2(n4921), .ZN(U3302) );
  AND2_X1 U5412 ( .A1(D_REG_19__SCAN_IN), .A2(n4921), .ZN(U3303) );
  NOR2_X1 U5413 ( .A1(n4923), .A2(n4914), .ZN(U3304) );
  AND2_X1 U5414 ( .A1(D_REG_17__SCAN_IN), .A2(n4921), .ZN(U3305) );
  NOR2_X1 U5415 ( .A1(n4923), .A2(n4915), .ZN(U3306) );
  AND2_X1 U5416 ( .A1(D_REG_15__SCAN_IN), .A2(n4921), .ZN(U3307) );
  AND2_X1 U5417 ( .A1(D_REG_14__SCAN_IN), .A2(n4921), .ZN(U3308) );
  AND2_X1 U5418 ( .A1(D_REG_13__SCAN_IN), .A2(n4921), .ZN(U3309) );
  NOR2_X1 U5419 ( .A1(n4923), .A2(n4916), .ZN(U3310) );
  NOR2_X1 U5420 ( .A1(n4923), .A2(n4917), .ZN(U3311) );
  AND2_X1 U5421 ( .A1(D_REG_10__SCAN_IN), .A2(n4921), .ZN(U3312) );
  AND2_X1 U5422 ( .A1(D_REG_9__SCAN_IN), .A2(n4921), .ZN(U3313) );
  NOR2_X1 U5423 ( .A1(n4923), .A2(n4918), .ZN(U3314) );
  AND2_X1 U5424 ( .A1(D_REG_7__SCAN_IN), .A2(n4921), .ZN(U3315) );
  NOR2_X1 U5425 ( .A1(n4923), .A2(n4919), .ZN(U3316) );
  NOR2_X1 U5426 ( .A1(n4923), .A2(n4920), .ZN(U3317) );
  AND2_X1 U5427 ( .A1(D_REG_4__SCAN_IN), .A2(n4921), .ZN(U3318) );
  AND2_X1 U5428 ( .A1(D_REG_3__SCAN_IN), .A2(n4921), .ZN(U3319) );
  NOR2_X1 U5429 ( .A1(n4923), .A2(n4922), .ZN(U3320) );
  INV_X1 U5430 ( .A(DATAI_23_), .ZN(n4925) );
  AOI21_X1 U5431 ( .B1(U3149), .B2(n4925), .A(n4924), .ZN(U3329) );
  AOI22_X1 U5432 ( .A1(STATE_REG_SCAN_IN), .A2(n4926), .B1(n2785), .B2(U3149), 
        .ZN(U3334) );
  AOI22_X1 U5433 ( .A1(STATE_REG_SCAN_IN), .A2(n4928), .B1(n4927), .B2(U3149), 
        .ZN(U3336) );
  AOI22_X1 U5434 ( .A1(STATE_REG_SCAN_IN), .A2(n4930), .B1(n4929), .B2(U3149), 
        .ZN(U3337) );
  AOI22_X1 U5435 ( .A1(STATE_REG_SCAN_IN), .A2(n4932), .B1(n4931), .B2(U3149), 
        .ZN(U3339) );
  AOI22_X1 U5436 ( .A1(STATE_REG_SCAN_IN), .A2(n2443), .B1(n2479), .B2(U3149), 
        .ZN(U3352) );
  AOI211_X1 U5437 ( .C1(n4951), .C2(n4935), .A(n4934), .B(n4933), .ZN(n4969)
         );
  AOI22_X1 U5438 ( .A1(n4967), .A2(n4969), .B1(n2473), .B2(n4965), .ZN(U3467)
         );
  OAI22_X1 U5439 ( .A1(n4938), .A2(n4937), .B1(n3076), .B2(n4936), .ZN(n4939)
         );
  NOR2_X1 U5440 ( .A1(n4940), .A2(n4939), .ZN(n4970) );
  INV_X1 U5441 ( .A(REG0_REG_1__SCAN_IN), .ZN(n4941) );
  AOI22_X1 U5442 ( .A1(n4967), .A2(n4970), .B1(n4941), .B2(n4965), .ZN(U3469)
         );
  AOI22_X1 U5443 ( .A1(n4944), .A2(n4951), .B1(n4943), .B2(n4942), .ZN(n4945)
         );
  AND2_X1 U5444 ( .A1(n4946), .A2(n4945), .ZN(n4972) );
  AOI22_X1 U5445 ( .A1(n4967), .A2(n4972), .B1(n2510), .B2(n4965), .ZN(U3473)
         );
  INV_X1 U5446 ( .A(n4947), .ZN(n4952) );
  INV_X1 U5447 ( .A(n4948), .ZN(n4950) );
  AOI211_X1 U5448 ( .C1(n4952), .C2(n4951), .A(n4950), .B(n4949), .ZN(n4973)
         );
  INV_X1 U5449 ( .A(REG0_REG_4__SCAN_IN), .ZN(n4953) );
  AOI22_X1 U5450 ( .A1(n4967), .A2(n4973), .B1(n4953), .B2(n4965), .ZN(U3475)
         );
  OAI22_X1 U5451 ( .A1(n4955), .A2(n4959), .B1(n4954), .B2(n3076), .ZN(n4956)
         );
  NOR2_X1 U5452 ( .A1(n4957), .A2(n4956), .ZN(n4974) );
  INV_X1 U5453 ( .A(REG0_REG_5__SCAN_IN), .ZN(n4958) );
  AOI22_X1 U5454 ( .A1(n4967), .A2(n4974), .B1(n4958), .B2(n4965), .ZN(U3477)
         );
  NOR3_X1 U5455 ( .A1(n4961), .A2(n4960), .A3(n4959), .ZN(n4964) );
  NOR3_X1 U5456 ( .A1(n4964), .A2(n4963), .A3(n4962), .ZN(n4978) );
  INV_X1 U5457 ( .A(REG0_REG_7__SCAN_IN), .ZN(n4966) );
  AOI22_X1 U5458 ( .A1(n4967), .A2(n4978), .B1(n4966), .B2(n4965), .ZN(U3481)
         );
  AOI22_X1 U5459 ( .A1(n4975), .A2(n4969), .B1(n4968), .B2(n4976), .ZN(U3518)
         );
  AOI22_X1 U5460 ( .A1(n4975), .A2(n4970), .B1(n4293), .B2(n4976), .ZN(U3519)
         );
  INV_X1 U5461 ( .A(REG1_REG_3__SCAN_IN), .ZN(n4971) );
  AOI22_X1 U5462 ( .A1(n4975), .A2(n4972), .B1(n4971), .B2(n4976), .ZN(U3521)
         );
  AOI22_X1 U5463 ( .A1(n4975), .A2(n4973), .B1(n4830), .B2(n4976), .ZN(U3522)
         );
  AOI22_X1 U5464 ( .A1(n4975), .A2(n4974), .B1(n2543), .B2(n4976), .ZN(U3523)
         );
  AOI22_X1 U5465 ( .A1(n4975), .A2(n4978), .B1(n4977), .B2(n4976), .ZN(U3525)
         );
  CLKBUF_X2 U2387 ( .A(n2493), .Z(n2133) );
  CLKBUF_X1 U2463 ( .A(n2509), .Z(n3462) );
endmodule

