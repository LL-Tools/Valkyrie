

module b21_C_2inp_gates_syn ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, 
        ADD_1071_U57, ADD_1071_U58, ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, 
        ADD_1071_U62, ADD_1071_U63, ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, 
        ADD_1071_U50, ADD_1071_U51, ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, 
        ADD_1071_U5, ADD_1071_U46, U126, U123, P1_U3353, P1_U3352, P1_U3351, 
        P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, 
        P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, 
        P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, 
        P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, 
        P1_U3322, P1_U3440, P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, 
        P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, 
        P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, 
        P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, 
        P1_U3296, P1_U3295, P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, 
        P1_U3460, P1_U3463, P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, 
        P1_U3481, P1_U3484, P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, 
        P1_U3502, P1_U3505, P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, 
        P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, 
        P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, 
        P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, 
        P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, 
        P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, 
        P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, 
        P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, 
        P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, 
        P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, 
        P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, 
        P1_U3355, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, 
        P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, 
        P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, 
        P1_U3242, P1_U3241, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, 
        P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, 
        P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, 
        P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, 
        P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, 
        P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, 
        P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, 
        P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, 
        P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, 
        P1_U3211, P1_U3084, P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, 
        P2_U3355, P2_U3354, P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, 
        P2_U3348, P2_U3347, P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, 
        P2_U3341, P2_U3340, P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, 
        P2_U3334, P2_U3333, P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, 
        P2_U3327, P2_U3437, P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, 
        P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, 
        P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, 
        P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, 
        P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, 
        P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, 
        P2_U3478, P2_U3481, P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, 
        P2_U3499, P2_U3502, P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, 
        P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, 
        P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, 
        P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, 
        P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, 
        P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, 
        P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, 
        P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, 
        P2_U3564, P2_U3565, P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, 
        P2_U3571, P2_U3572, P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, 
        P2_U3578, P2_U3579, P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, 
        P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3152, P2_U3151, P2_U3966, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283,
         n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293,
         n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303,
         n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313,
         n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323,
         n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333,
         n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343,
         n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353,
         n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363,
         n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373,
         n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383,
         n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393,
         n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403,
         n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413,
         n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423,
         n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433,
         n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443,
         n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453,
         n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463,
         n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473,
         n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483,
         n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493,
         n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503,
         n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513,
         n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523,
         n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533,
         n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543,
         n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553,
         n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563,
         n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573,
         n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583,
         n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593,
         n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603,
         n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613,
         n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623,
         n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633,
         n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643,
         n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653,
         n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663,
         n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673,
         n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683,
         n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693,
         n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703,
         n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713,
         n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723,
         n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733,
         n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743,
         n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753,
         n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763,
         n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773,
         n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783,
         n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793,
         n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803,
         n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813,
         n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823,
         n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833,
         n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843,
         n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853,
         n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863,
         n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873,
         n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883,
         n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893,
         n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903,
         n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913,
         n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923,
         n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4932, n4933, n4934,
         n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944,
         n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954,
         n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964,
         n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974,
         n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984,
         n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994,
         n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004,
         n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014,
         n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024,
         n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034,
         n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044,
         n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054,
         n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064,
         n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074,
         n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084,
         n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094,
         n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104,
         n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114,
         n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124,
         n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134,
         n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144,
         n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154,
         n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164,
         n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174,
         n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184,
         n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194,
         n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204,
         n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214,
         n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224,
         n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234,
         n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244,
         n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254,
         n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264,
         n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274,
         n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284,
         n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294,
         n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304,
         n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314,
         n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324,
         n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334,
         n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344,
         n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354,
         n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364,
         n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374,
         n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384,
         n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394,
         n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404,
         n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414,
         n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424,
         n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434,
         n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444,
         n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454,
         n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464,
         n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474,
         n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484,
         n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494,
         n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504,
         n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514,
         n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524,
         n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534,
         n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544,
         n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554,
         n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564,
         n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574,
         n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584,
         n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594,
         n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604,
         n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614,
         n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624,
         n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634,
         n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644,
         n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654,
         n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664,
         n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674,
         n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684,
         n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694,
         n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704,
         n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714,
         n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724,
         n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734,
         n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744,
         n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754,
         n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764,
         n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774,
         n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784,
         n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794,
         n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804,
         n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814,
         n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824,
         n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834,
         n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844,
         n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854,
         n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864,
         n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874,
         n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884,
         n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894,
         n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904,
         n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914,
         n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924,
         n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934,
         n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944,
         n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954,
         n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964,
         n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974,
         n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984,
         n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994,
         n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004,
         n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014,
         n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024,
         n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034,
         n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044,
         n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054,
         n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064,
         n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074,
         n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084,
         n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094,
         n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104,
         n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114,
         n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124,
         n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134,
         n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144,
         n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154,
         n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164,
         n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174,
         n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184,
         n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194,
         n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204,
         n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214,
         n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224,
         n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234,
         n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244,
         n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254,
         n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264,
         n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274,
         n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284,
         n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294,
         n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304,
         n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314,
         n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324,
         n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334,
         n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344,
         n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354,
         n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364,
         n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374,
         n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384,
         n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394,
         n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404,
         n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414,
         n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424,
         n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434,
         n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444,
         n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454,
         n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464,
         n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474,
         n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484,
         n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494,
         n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504,
         n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514,
         n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524,
         n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534,
         n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544,
         n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554,
         n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564,
         n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574,
         n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584,
         n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594,
         n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604,
         n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614,
         n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624,
         n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634,
         n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644,
         n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654,
         n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664,
         n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674,
         n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684,
         n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694,
         n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704,
         n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714,
         n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724,
         n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734,
         n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744,
         n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754,
         n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764,
         n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774,
         n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784,
         n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794,
         n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804,
         n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814,
         n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824,
         n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834,
         n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844,
         n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854,
         n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864,
         n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874,
         n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884,
         n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894,
         n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904,
         n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914,
         n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924,
         n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934,
         n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944,
         n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954,
         n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964,
         n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974,
         n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984,
         n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994,
         n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004,
         n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014,
         n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024,
         n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034,
         n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044,
         n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054,
         n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064,
         n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074,
         n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084,
         n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094,
         n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104,
         n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114,
         n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124,
         n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134,
         n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144,
         n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154,
         n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164,
         n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174,
         n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184,
         n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194,
         n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204,
         n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214,
         n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224,
         n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234,
         n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244,
         n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254,
         n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264,
         n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274,
         n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284,
         n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294,
         n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304,
         n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314,
         n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324,
         n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334,
         n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344,
         n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354,
         n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364,
         n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374,
         n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384,
         n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394,
         n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404,
         n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414,
         n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424,
         n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434,
         n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444,
         n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454,
         n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464,
         n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474,
         n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484,
         n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494,
         n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504,
         n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514,
         n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524,
         n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534,
         n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544,
         n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554,
         n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564,
         n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574,
         n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584,
         n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594,
         n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604,
         n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614,
         n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624,
         n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634,
         n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644,
         n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654,
         n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664,
         n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674,
         n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684,
         n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694,
         n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704,
         n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714,
         n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724,
         n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734,
         n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744,
         n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754,
         n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764,
         n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774,
         n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784,
         n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794,
         n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804,
         n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814,
         n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824,
         n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834,
         n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844,
         n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854,
         n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864,
         n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874,
         n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884,
         n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894,
         n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904,
         n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914,
         n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924,
         n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934,
         n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944,
         n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954,
         n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964,
         n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974,
         n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984,
         n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994,
         n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004,
         n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014,
         n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024,
         n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034,
         n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044,
         n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054,
         n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064,
         n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074,
         n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084,
         n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094,
         n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104,
         n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114,
         n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124,
         n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134,
         n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144,
         n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154,
         n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164,
         n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174,
         n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184,
         n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194,
         n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204,
         n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214,
         n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224,
         n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234,
         n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244,
         n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254,
         n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264,
         n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274,
         n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284,
         n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294,
         n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304,
         n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314,
         n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324,
         n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334,
         n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344,
         n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354,
         n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364,
         n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374,
         n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384,
         n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394,
         n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404,
         n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414,
         n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424,
         n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434,
         n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444,
         n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454,
         n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464,
         n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474,
         n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484,
         n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494,
         n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504,
         n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514,
         n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524,
         n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534,
         n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544,
         n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554,
         n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564,
         n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574,
         n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584,
         n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594,
         n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604,
         n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614,
         n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624,
         n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634,
         n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644,
         n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654,
         n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664,
         n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674,
         n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684,
         n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694,
         n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704,
         n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714,
         n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724,
         n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734,
         n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744,
         n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754,
         n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764,
         n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774,
         n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784,
         n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794,
         n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804,
         n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814,
         n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824,
         n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834,
         n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844,
         n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854,
         n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864,
         n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874,
         n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884,
         n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894,
         n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904,
         n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914,
         n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924,
         n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934,
         n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944,
         n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954,
         n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964,
         n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974,
         n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984,
         n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994,
         n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004,
         n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014,
         n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024,
         n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034,
         n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044,
         n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054,
         n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064,
         n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074,
         n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084,
         n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094,
         n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104,
         n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114,
         n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124,
         n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134,
         n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144,
         n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154,
         n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164,
         n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174,
         n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184,
         n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194,
         n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204,
         n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214,
         n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224,
         n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234,
         n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244,
         n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254,
         n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264,
         n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274,
         n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284,
         n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294,
         n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304,
         n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314,
         n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324,
         n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334,
         n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344,
         n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354,
         n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364,
         n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374,
         n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384,
         n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394,
         n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404,
         n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414,
         n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424,
         n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434,
         n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444,
         n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454,
         n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464,
         n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474,
         n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484,
         n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494,
         n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504,
         n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514,
         n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524,
         n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534,
         n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544,
         n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554,
         n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564,
         n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574,
         n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584,
         n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594,
         n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604,
         n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614,
         n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624,
         n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634,
         n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644,
         n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654,
         n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664,
         n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674,
         n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684,
         n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694,
         n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704,
         n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714,
         n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724,
         n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734,
         n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744,
         n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754,
         n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764,
         n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774,
         n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784,
         n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794,
         n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804,
         n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814,
         n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824,
         n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834,
         n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844,
         n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854,
         n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864,
         n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874,
         n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884,
         n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894,
         n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904,
         n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914,
         n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924,
         n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934,
         n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944,
         n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954,
         n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964,
         n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974,
         n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984,
         n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994,
         n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003,
         n10004, n10005, n10006, n10007, n10008, n10009, n10010, n10011,
         n10012, n10013, n10014, n10015, n10016, n10017, n10018, n10019,
         n10020, n10021, n10022, n10023, n10024, n10025, n10026, n10027,
         n10028, n10029, n10030, n10031, n10032, n10033, n10034, n10035,
         n10036, n10037, n10038, n10039, n10040, n10041, n10042, n10043,
         n10044, n10045, n10046, n10047, n10048, n10049, n10050, n10051,
         n10052, n10053, n10054, n10055, n10056, n10057, n10058, n10059,
         n10060, n10061, n10062, n10063, n10064, n10065, n10066, n10067,
         n10068, n10069, n10070, n10071, n10072, n10073, n10074, n10075,
         n10076, n10077, n10078, n10079, n10080, n10081, n10082, n10083,
         n10084, n10085, n10086, n10087, n10088, n10089, n10090, n10091,
         n10092, n10093, n10094, n10095, n10096, n10097, n10098, n10099,
         n10100, n10101, n10102, n10103, n10104, n10105, n10106, n10107,
         n10108, n10109, n10110, n10111, n10112, n10113, n10114, n10115,
         n10116, n10117, n10118, n10119, n10120, n10121, n10122, n10123,
         n10124, n10125, n10126, n10127, n10128, n10129, n10130, n10131,
         n10132, n10133, n10134, n10135, n10136, n10137, n10138, n10139,
         n10140, n10141, n10142, n10143, n10144, n10145, n10146, n10147,
         n10148, n10149, n10150, n10151, n10152, n10153, n10154, n10155,
         n10156, n10157, n10158, n10159, n10160, n10161, n10162, n10163,
         n10164, n10165, n10166, n10167, n10168, n10169, n10170, n10171,
         n10172, n10173, n10174, n10175, n10176, n10177, n10178, n10179,
         n10180, n10181, n10182, n10183, n10184, n10185, n10186, n10187,
         n10188, n10189, n10190, n10191, n10192, n10193, n10194, n10195,
         n10196, n10197, n10198, n10199, n10200, n10201, n10202, n10203,
         n10204, n10205, n10206, n10207, n10208, n10209, n10210, n10211,
         n10212, n10213, n10214, n10215, n10216, n10217, n10218, n10219,
         n10220, n10221, n10222, n10223, n10224, n10225, n10226, n10227,
         n10228, n10229, n10230, n10231, n10232, n10233, n10234, n10235,
         n10236, n10237, n10238, n10239, n10240, n10241, n10242, n10243,
         n10244, n10245, n10246, n10247, n10248, n10249, n10250, n10251,
         n10252, n10253, n10254, n10255, n10256, n10257, n10258, n10259,
         n10260, n10261, n10262, n10263, n10264, n10265, n10266, n10267,
         n10268, n10269, n10270, n10271, n10272, n10273, n10274, n10275,
         n10276, n10277, n10278, n10279, n10280, n10281, n10282, n10283,
         n10284, n10285, n10286, n10287, n10288, n10289, n10290, n10291,
         n10292, n10293, n10294, n10295, n10296, n10297, n10298, n10299,
         n10300, n10301, n10302, n10303, n10304;

  CLKBUF_X1 U4779 ( .A(n7036), .Z(n4296) );
  NAND2_X1 U4780 ( .A1(n5986), .A2(n5985), .ZN(n8506) );
  CLKBUF_X2 U4782 ( .A(n6992), .Z(n4285) );
  INV_X1 U4783 ( .A(n7027), .ZN(n10062) );
  CLKBUF_X2 U4784 ( .A(n5743), .Z(n4298) );
  BUF_X2 U4785 ( .A(n5743), .Z(n4297) );
  CLKBUF_X1 U4786 ( .A(n8781), .Z(n4277) );
  INV_X2 U4787 ( .A(n5025), .ZN(n4287) );
  CLKBUF_X1 U4788 ( .A(n5025), .Z(n6562) );
  INV_X2 U4789 ( .A(n9541), .ZN(n9877) );
  AND2_X1 U4790 ( .A1(n9362), .A2(n4528), .ZN(n4527) );
  OAI21_X2 U4791 ( .B1(n7771), .B2(n4866), .A(n4450), .ZN(n8403) );
  NOR2_X1 U4792 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n5783) );
  INV_X1 U4794 ( .A(n7073), .ZN(n8711) );
  INV_X1 U4796 ( .A(n4302), .ZN(n6387) );
  AND3_X1 U4797 ( .A1(n5855), .A2(n5854), .A3(n5853), .ZN(n10056) );
  NAND2_X1 U4798 ( .A1(n5764), .A2(n4861), .ZN(n9299) );
  OAI21_X1 U4799 ( .B1(n4856), .B2(n5159), .A(n4854), .ZN(n5182) );
  INV_X1 U4800 ( .A(n4280), .ZN(n6179) );
  CLKBUF_X2 U4801 ( .A(n5857), .Z(n6076) );
  OR2_X1 U4802 ( .A1(n4288), .A2(n6729), .ZN(n5833) );
  CLKBUF_X3 U4803 ( .A(n5898), .Z(n6182) );
  AND3_X1 U4804 ( .A1(n5444), .A2(n5443), .A3(n5442), .ZN(n9638) );
  NAND2_X1 U4805 ( .A1(n9070), .A2(n9126), .ZN(n9323) );
  INV_X1 U4806 ( .A(n9889), .ZN(n7300) );
  OR2_X1 U4807 ( .A1(n5003), .A2(n9752), .ZN(n5001) );
  INV_X1 U4808 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5615) );
  INV_X1 U4809 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n5200) );
  AND3_X2 U4810 ( .A1(n5822), .A2(n5821), .A3(n5820), .ZN(n10041) );
  INV_X2 U4811 ( .A(n8417), .ZN(n4281) );
  INV_X1 U4812 ( .A(n7282), .ZN(n9896) );
  INV_X1 U4813 ( .A(n9638), .ZN(n9456) );
  NAND4_X2 U4814 ( .A1(n5089), .A2(n5088), .A3(n5087), .A4(n5086), .ZN(n9231)
         );
  CLKBUF_X3 U4815 ( .A(n5856), .Z(n4280) );
  INV_X1 U4816 ( .A(n6724), .ZN(n5870) );
  OR2_X1 U4817 ( .A1(n8206), .A2(n8523), .ZN(n4274) );
  OAI21_X2 U4818 ( .B1(n6245), .B2(n7515), .A(n6246), .ZN(n7571) );
  NAND2_X2 U4819 ( .A1(n4425), .A2(n5081), .ZN(n4453) );
  NAND2_X2 U4820 ( .A1(n8281), .A2(n8287), .ZN(n8280) );
  BUF_X2 U4821 ( .A(n6164), .Z(n4288) );
  NAND2_X2 U4822 ( .A1(n7893), .A2(n4916), .ZN(n7399) );
  INV_X2 U4823 ( .A(n6000), .ZN(n6139) );
  NOR2_X2 U4824 ( .A1(n5253), .A2(n5252), .ZN(n5279) );
  NAND3_X2 U4825 ( .A1(n7540), .A2(n4728), .A3(n4332), .ZN(n4724) );
  OAI22_X2 U4826 ( .A1(n6873), .A2(n6872), .B1(P1_REG2_REG_8__SCAN_IN), .B2(
        n6871), .ZN(n6874) );
  AOI21_X1 U4827 ( .B1(n4527), .B2(n9086), .A(n4525), .ZN(n4524) );
  NAND2_X2 U4828 ( .A1(n8245), .A2(n8178), .ZN(n8230) );
  XNOR2_X2 U4829 ( .A(n5001), .B(n5000), .ZN(n9758) );
  NAND2_X2 U4830 ( .A1(n6171), .A2(n6187), .ZN(n7368) );
  MUX2_X2 U4831 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6169), .S(
        P2_IR_REG_21__SCAN_IN), .Z(n6171) );
  OR2_X1 U4832 ( .A1(n5857), .A2(n6781), .ZN(n5832) );
  NAND2_X1 U4833 ( .A1(n6368), .A2(n6371), .ZN(n4275) );
  NAND2_X1 U4834 ( .A1(n6368), .A2(n6371), .ZN(n4276) );
  NAND2_X1 U4835 ( .A1(n6368), .A2(n6371), .ZN(n6724) );
  BUF_X4 U4838 ( .A(n8781), .Z(n4278) );
  AND2_X2 U4839 ( .A1(n7158), .A2(n6988), .ZN(n8781) );
  AND2_X1 U4840 ( .A1(n4543), .A2(n4542), .ZN(n4279) );
  INV_X2 U4841 ( .A(n5025), .ZN(n6561) );
  NAND2_X2 U4842 ( .A1(n7391), .A2(n7390), .ZN(n7540) );
  NAND2_X2 U4843 ( .A1(n7224), .A2(n4282), .ZN(n7391) );
  NAND2_X1 U4844 ( .A1(n7582), .A2(n7583), .ZN(n4959) );
  OR2_X1 U4845 ( .A1(n9312), .A2(n9515), .ZN(n4534) );
  AOI21_X1 U4846 ( .B1(n4556), .B2(n4576), .A(n8207), .ZN(n4555) );
  NAND2_X1 U4847 ( .A1(n5643), .A2(n9170), .ZN(n9376) );
  INV_X1 U4848 ( .A(n9216), .ZN(n9349) );
  NAND3_X1 U4849 ( .A1(n9136), .A2(n9134), .A3(n7309), .ZN(n7308) );
  AOI21_X1 U4850 ( .B1(n7044), .B2(n6399), .A(n7051), .ZN(n6403) );
  INV_X4 U4851 ( .A(n8779), .ZN(n8774) );
  CLKBUF_X2 U4852 ( .A(n7073), .Z(n4476) );
  CLKBUF_X1 U4853 ( .A(n7323), .Z(n4290) );
  INV_X1 U4854 ( .A(n8067), .ZN(n5868) );
  CLKBUF_X2 U4855 ( .A(n5399), .Z(n5584) );
  NAND4_X1 U4856 ( .A1(n5862), .A2(n5861), .A3(n5860), .A4(n5859), .ZN(n8067)
         );
  XNOR2_X1 U4857 ( .A(n5616), .B(n5615), .ZN(n8993) );
  INV_X1 U4858 ( .A(n6349), .ZN(n6347) );
  NAND4_X1 U4859 ( .A1(n5847), .A2(n5846), .A3(n5845), .A4(n5844), .ZN(n8068)
         );
  INV_X4 U4860 ( .A(n4289), .ZN(n6174) );
  CLKBUF_X2 U4861 ( .A(n5858), .Z(n5892) );
  BUF_X2 U4862 ( .A(n6164), .Z(n4289) );
  INV_X2 U4863 ( .A(n7861), .ZN(n10090) );
  BUF_X1 U4864 ( .A(n7004), .Z(n4300) );
  INV_X2 U4866 ( .A(n5025), .ZN(n4286) );
  AND4_X1 U4867 ( .A1(n6377), .A2(n7507), .A3(n7034), .A4(n10089), .ZN(n4981)
         );
  AOI21_X1 U4868 ( .B1(n6354), .B2(n6353), .A(n6352), .ZN(n6377) );
  OAI21_X1 U4869 ( .B1(n8445), .B2(n8379), .A(n4409), .ZN(n4408) );
  AOI21_X1 U4870 ( .B1(n4578), .B2(n6346), .A(n6345), .ZN(n6186) );
  NAND2_X1 U4871 ( .A1(n8230), .A2(n8237), .ZN(n8229) );
  AOI21_X1 U4872 ( .B1(n4452), .B2(n8186), .A(n8185), .ZN(n8190) );
  AOI21_X1 U4873 ( .B1(n4742), .B2(n10017), .A(n4410), .ZN(n8444) );
  NAND2_X1 U4874 ( .A1(n4553), .A2(n4551), .ZN(n8185) );
  NAND2_X1 U4875 ( .A1(n8855), .A2(n8643), .ZN(n8762) );
  NAND2_X1 U4876 ( .A1(n4807), .A2(n4805), .ZN(n8855) );
  CLKBUF_X1 U4877 ( .A(n8903), .Z(n4490) );
  NAND3_X1 U4878 ( .A1(n8340), .A2(n8332), .A3(n8331), .ZN(n6071) );
  CLKBUF_X1 U4879 ( .A(n4915), .Z(n4447) );
  NAND2_X1 U4880 ( .A1(n4797), .A2(n4800), .ZN(n8878) );
  AOI21_X1 U4881 ( .B1(n4524), .B2(n4526), .A(n4522), .ZN(n4521) );
  NAND2_X1 U4882 ( .A1(n9184), .A2(n9307), .ZN(n5762) );
  OR2_X1 U4883 ( .A1(n9298), .A2(n9591), .ZN(n9184) );
  OR2_X1 U4884 ( .A1(n8447), .A2(n8179), .ZN(n6338) );
  OR2_X1 U4885 ( .A1(n9603), .A2(n8964), .ZN(n9070) );
  NOR2_X1 U4886 ( .A1(n4352), .A2(n4597), .ZN(n4596) );
  XNOR2_X1 U4887 ( .A(n4784), .B(n9263), .ZN(n7674) );
  OR2_X1 U4888 ( .A1(n5464), .A2(n5463), .ZN(n5486) );
  NOR2_X1 U4889 ( .A1(n4350), .A2(n4451), .ZN(n4450) );
  NAND2_X1 U4890 ( .A1(n7132), .A2(n6423), .ZN(n7893) );
  OR2_X2 U4891 ( .A1(n9369), .A2(n9350), .ZN(n9177) );
  INV_X1 U4892 ( .A(n8381), .ZN(n4719) );
  NAND2_X1 U4893 ( .A1(n6052), .A2(n6051), .ZN(n8482) );
  NAND2_X1 U4894 ( .A1(n6029), .A2(n6028), .ZN(n8490) );
  NAND2_X1 U4895 ( .A1(n6017), .A2(n6016), .ZN(n8494) );
  XNOR2_X1 U4896 ( .A(n5398), .B(n5412), .ZN(n7213) );
  NAND2_X1 U4897 ( .A1(n6003), .A2(n6002), .ZN(n8501) );
  NAND2_X1 U4898 ( .A1(n5884), .A2(n6241), .ZN(n7447) );
  NAND2_X1 U4899 ( .A1(n6271), .A2(n7707), .ZN(n7736) );
  OR2_X1 U4900 ( .A1(n7737), .A2(n7846), .ZN(n7841) );
  OAI211_X1 U4901 ( .C1(n7046), .C2(n6404), .A(n6403), .B(n7054), .ZN(n7052)
         );
  AND2_X1 U4902 ( .A1(n7079), .A2(n7152), .ZN(n7084) );
  OR2_X1 U4903 ( .A1(n8506), .A2(n7734), .ZN(n6294) );
  AND4_X2 U4904 ( .A1(n5537), .A2(n5536), .A3(n5535), .A4(n5534), .ZN(n9350)
         );
  NAND2_X1 U4905 ( .A1(n5322), .A2(n5321), .ZN(n9678) );
  NOR2_X1 U4906 ( .A1(n6618), .A2(n4300), .ZN(n9855) );
  INV_X1 U4907 ( .A(n7219), .ZN(n7221) );
  NAND2_X1 U4908 ( .A1(n5973), .A2(n5972), .ZN(n8511) );
  NAND2_X1 U4909 ( .A1(n5936), .A2(n5935), .ZN(n7704) );
  NOR2_X1 U4910 ( .A1(P1_U3083), .A2(n6604), .ZN(n9810) );
  AND2_X1 U4911 ( .A1(n6278), .A2(n7545), .ZN(n7539) );
  INV_X1 U4912 ( .A(n7227), .ZN(n4282) );
  NAND2_X1 U4913 ( .A1(n5922), .A2(n5921), .ZN(n7885) );
  AND2_X1 U4914 ( .A1(n7191), .A2(n6396), .ZN(n7044) );
  NAND2_X1 U4915 ( .A1(n9130), .A2(n5627), .ZN(n9093) );
  OR2_X1 U4916 ( .A1(n7199), .A2(n6401), .ZN(n6402) );
  NAND2_X1 U4917 ( .A1(n4729), .A2(n5912), .ZN(n7389) );
  AND2_X1 U4918 ( .A1(n6262), .A2(n6266), .ZN(n7451) );
  AOI22_X1 U4919 ( .A1(n6867), .A2(n6866), .B1(n6865), .B2(n6870), .ZN(n6881)
         );
  AND2_X1 U4920 ( .A1(n6386), .A2(n7858), .ZN(n6914) );
  AND2_X1 U4921 ( .A1(n4560), .A2(n4559), .ZN(n6873) );
  AND4_X1 U4922 ( .A1(n5176), .A2(n5175), .A3(n5174), .A4(n5173), .ZN(n8953)
         );
  CLKBUF_X2 U4923 ( .A(n7526), .Z(n4284) );
  CLKBUF_X2 U4924 ( .A(n6466), .Z(n4302) );
  XNOR2_X1 U4925 ( .A(n5186), .B(n5185), .ZN(n6579) );
  NAND2_X1 U4926 ( .A1(n5184), .A2(n5183), .ZN(n5186) );
  NAND4_X1 U4927 ( .A1(n5111), .A2(n5110), .A3(n5109), .A4(n5108), .ZN(n9915)
         );
  OR2_X1 U4928 ( .A1(n8993), .A2(n9119), .ZN(n4818) );
  AND4_X2 U4929 ( .A1(n5070), .A2(n5069), .A3(n5068), .A4(n5067), .ZN(n5105)
         );
  AND4_X1 U4930 ( .A1(n5125), .A2(n5124), .A3(n5123), .A4(n5122), .ZN(n9928)
         );
  AND2_X1 U4931 ( .A1(n5867), .A2(n5866), .ZN(n7027) );
  CLKBUF_X3 U4932 ( .A(n5652), .Z(n4467) );
  NAND2_X1 U4933 ( .A1(n4546), .A2(n5057), .ZN(n5060) );
  AND4_X1 U4934 ( .A1(n5908), .A2(n5907), .A3(n5906), .A4(n5905), .ZN(n7135)
         );
  AND2_X1 U4935 ( .A1(n5944), .A2(n5934), .ZN(n8108) );
  CLKBUF_X1 U4936 ( .A(n5399), .Z(n5742) );
  AND4_X1 U4937 ( .A1(n5896), .A2(n5895), .A3(n5894), .A4(n5893), .ZN(n7059)
         );
  INV_X1 U4938 ( .A(n6494), .ZN(n4283) );
  NAND2_X1 U4939 ( .A1(n5614), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5616) );
  CLKBUF_X1 U4940 ( .A(n9198), .Z(n4480) );
  NAND2_X1 U4941 ( .A1(n4430), .A2(n4429), .ZN(n7158) );
  NAND4_X2 U4942 ( .A1(n5834), .A2(n5833), .A3(n5831), .A4(n5832), .ZN(n6388)
         );
  OAI21_X1 U4943 ( .B1(P1_REG2_REG_4__SCAN_IN), .B2(n6630), .A(n6896), .ZN(
        n6651) );
  AND2_X2 U4944 ( .A1(n5009), .A2(n9761), .ZN(n5441) );
  NAND2_X1 U4945 ( .A1(n4294), .A2(n6562), .ZN(n5452) );
  NAND2_X1 U4946 ( .A1(n5126), .A2(n4547), .ZN(n4856) );
  NOR2_X1 U4947 ( .A1(n5417), .A2(n4636), .ZN(n4635) );
  NAND2_X1 U4948 ( .A1(n5613), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5618) );
  INV_X1 U4949 ( .A(n5848), .ZN(n5898) );
  CLKBUF_X2 U4950 ( .A(n7381), .Z(n4301) );
  NAND2_X1 U4951 ( .A1(n5046), .A2(n5045), .ZN(n5126) );
  NAND2_X1 U4952 ( .A1(n8553), .A2(n5805), .ZN(n5858) );
  AND2_X1 U4953 ( .A1(n5803), .A2(n8553), .ZN(n5856) );
  NAND2_X1 U4954 ( .A1(n5004), .A2(n9753), .ZN(n9761) );
  XNOR2_X1 U4955 ( .A(n5620), .B(n5619), .ZN(n9120) );
  NAND2_X1 U4956 ( .A1(n5804), .A2(n5805), .ZN(n5857) );
  INV_X1 U4957 ( .A(n8352), .ZN(n8392) );
  OR2_X1 U4958 ( .A1(n5309), .A2(n8904), .ZN(n5324) );
  NAND2_X1 U4959 ( .A1(n5042), .A2(n5041), .ZN(n5112) );
  NAND2_X1 U4960 ( .A1(n5612), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5620) );
  NOR2_X1 U4961 ( .A1(n5243), .A2(n5242), .ZN(n5265) );
  XNOR2_X1 U4962 ( .A(n5072), .B(n5071), .ZN(n5074) );
  NAND2_X1 U4963 ( .A1(n4817), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5611) );
  XNOR2_X1 U4964 ( .A(n5047), .B(SI_4_), .ZN(n5127) );
  NAND2_X1 U4965 ( .A1(n4448), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6189) );
  NAND2_X1 U4966 ( .A1(n5038), .A2(n5037), .ZN(n5072) );
  NAND2_X1 U4967 ( .A1(n6187), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6194) );
  NAND2_X1 U4968 ( .A1(n5801), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5797) );
  XNOR2_X1 U4969 ( .A(n5051), .B(SI_5_), .ZN(n5159) );
  NAND2_X2 U4970 ( .A1(n4287), .A2(P1_U3084), .ZN(n9763) );
  NAND2_X1 U4971 ( .A1(n4704), .A2(n4703), .ZN(n5044) );
  NAND2_X2 U4972 ( .A1(n6562), .A2(P2_U3152), .ZN(n8550) );
  AND2_X2 U4973 ( .A1(n4543), .A2(n4542), .ZN(n5025) );
  OR2_X1 U4974 ( .A1(n5693), .A2(P1_IR_REG_23__SCAN_IN), .ZN(n4996) );
  INV_X1 U4975 ( .A(n4796), .ZN(n5075) );
  NAND2_X1 U4976 ( .A1(n9752), .A2(n4999), .ZN(n4443) );
  AND3_X1 U4977 ( .A1(n5114), .A2(n5130), .A3(n4744), .ZN(n4743) );
  NAND2_X1 U4978 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n5799), .ZN(n5800) );
  INV_X1 U4979 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n5302) );
  INV_X1 U4980 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5610) );
  INV_X1 U4981 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5619) );
  INV_X1 U4982 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5340) );
  INV_X1 U4983 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n6014) );
  INV_X1 U4984 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n5020) );
  INV_X4 U4985 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  INV_X1 U4986 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n4457) );
  INV_X4 U4987 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  INV_X1 U4988 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n5850) );
  INV_X1 U4989 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n4545) );
  INV_X1 U4990 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n10218) );
  NAND2_X1 U4991 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_28__SCAN_IN), 
        .ZN(n4663) );
  INV_X1 U4992 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n6359) );
  NAND2_X2 U4993 ( .A1(n5557), .A2(n5556), .ZN(n9335) );
  AND2_X1 U4994 ( .A1(n6415), .A2(n6410), .ZN(n4919) );
  NAND2_X1 U4995 ( .A1(n5878), .A2(n5877), .ZN(n7526) );
  BUF_X1 U4996 ( .A(n5016), .Z(n5017) );
  NAND2_X1 U4997 ( .A1(n6988), .A2(n4818), .ZN(n6992) );
  OAI222_X1 U4998 ( .A1(P1_U3084), .A2(n8993), .B1(n9763), .B2(n7896), .C1(
        n7350), .C2(n7782), .ZN(P1_U3331) );
  NOR3_X4 U4999 ( .A1(n4710), .A2(n4709), .A3(n8176), .ZN(n8281) );
  NOR4_X2 U5000 ( .A1(n9206), .A2(n9205), .A3(n9204), .A4(n9203), .ZN(n9207)
         );
  NAND2_X1 U5001 ( .A1(n4550), .A2(n4555), .ZN(n8204) );
  AND2_X1 U5002 ( .A1(n6402), .A2(n6405), .ZN(n7054) );
  OR2_X1 U5003 ( .A1(n6383), .A2(n10041), .ZN(n6246) );
  XNOR2_X1 U5004 ( .A(n4283), .B(n10041), .ZN(n6912) );
  NAND2_X1 U5005 ( .A1(n5804), .A2(n5803), .ZN(n6164) );
  AOI21_X2 U5006 ( .B1(n4959), .B2(n4957), .A(n4372), .ZN(n7452) );
  XNOR2_X1 U5007 ( .A(n5997), .B(P2_IR_REG_14__SCAN_IN), .ZN(n7323) );
  XNOR2_X1 U5008 ( .A(n6189), .B(P2_IR_REG_19__SCAN_IN), .ZN(n8352) );
  OR2_X1 U5009 ( .A1(n5848), .A2(n5835), .ZN(n5839) );
  AOI22_X2 U5010 ( .A1(n8438), .A2(n10019), .B1(n10063), .B2(n8437), .ZN(n8439) );
  OR2_X1 U5011 ( .A1(n6000), .A2(n6564), .ZN(n5840) );
  AOI211_X1 U5012 ( .C1(n5841), .C2(n7574), .A(n4296), .B(n10021), .ZN(n10047)
         );
  MUX2_X2 U5013 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n4333), .S(n10100), .Z(
        P2_U3548) );
  NAND2_X1 U5014 ( .A1(n4733), .A2(n4318), .ZN(n4911) );
  NAND2_X2 U5015 ( .A1(n6421), .A2(n7129), .ZN(n7132) );
  NAND2_X1 U5016 ( .A1(n5751), .A2(n4299), .ZN(n4294) );
  NAND2_X1 U5017 ( .A1(n5751), .A2(n4299), .ZN(n4295) );
  NAND2_X1 U5018 ( .A1(n5751), .A2(n4299), .ZN(n5451) );
  MUX2_X2 U5019 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n4333), .S(n10283), .Z(
        P2_U3516) );
  OR2_X2 U5020 ( .A1(n4411), .A2(n4706), .ZN(n4333) );
  INV_X2 U5021 ( .A(n6494), .ZN(n6510) );
  NOR2_X1 U5022 ( .A1(n5016), .A2(n4998), .ZN(n5014) );
  AND2_X1 U5023 ( .A1(n8217), .A2(n4341), .ZN(n8445) );
  NOR2_X2 U5024 ( .A1(n7427), .A2(n7426), .ZN(n7439) );
  NAND2_X1 U5025 ( .A1(n6512), .A2(n4301), .ZN(n7036) );
  INV_X1 U5026 ( .A(n5452), .ZN(n5743) );
  AND2_X2 U5027 ( .A1(n9319), .A2(n4940), .ZN(n9301) );
  NAND3_X1 U5029 ( .A1(n4444), .A2(n5015), .A3(n4443), .ZN(n7004) );
  OR2_X2 U5030 ( .A1(n7584), .A2(n4284), .ZN(n7455) );
  INV_X2 U5031 ( .A(n6388), .ZN(n5842) );
  NAND4_X2 U5032 ( .A1(n4648), .A2(n5851), .A3(n4647), .A4(n4646), .ZN(n6026)
         );
  NAND2_X1 U5033 ( .A1(n4275), .A2(n4287), .ZN(n6000) );
  OAI21_X1 U5034 ( .B1(n7947), .B2(n4922), .A(n4920), .ZN(n7901) );
  NAND2_X2 U5035 ( .A1(n8229), .A2(n8180), .ZN(n8218) );
  AOI21_X2 U5036 ( .B1(n8403), .B2(n6304), .A(n6024), .ZN(n8384) );
  OAI222_X1 U5037 ( .A1(P1_U3084), .A2(n6584), .B1(n9763), .B2(n5835), .C1(
        n6583), .C2(n7782), .ZN(P1_U3351) );
  OAI222_X1 U5038 ( .A1(n6794), .A2(P2_U3152), .B1(n8550), .B2(n5835), .C1(
        n6564), .C2(n8552), .ZN(P2_U3356) );
  XNOR2_X1 U5039 ( .A(n5074), .B(n5073), .ZN(n5835) );
  NOR2_X2 U5040 ( .A1(n8248), .A2(n8447), .ZN(n8232) );
  OAI21_X2 U5041 ( .B1(n4732), .B2(n8384), .A(n4730), .ZN(n8341) );
  XNOR2_X1 U5042 ( .A(n6192), .B(n6191), .ZN(n7381) );
  NOR2_X2 U5043 ( .A1(n10164), .A2(n5533), .ZN(n5550) );
  NOR3_X4 U5044 ( .A1(n8314), .A2(n4789), .A3(n8456), .ZN(n8265) );
  OR2_X4 U5045 ( .A1(n8346), .A2(n8476), .ZN(n8314) );
  OAI222_X1 U5046 ( .A1(n8552), .A2(n7836), .B1(P2_U3152), .B2(n6371), .C1(
        n8550), .C2(n7835), .ZN(P2_U3330) );
  INV_X1 U5047 ( .A(n5237), .ZN(n4860) );
  OAI21_X1 U5048 ( .B1(n5025), .B2(n4610), .A(n4609), .ZN(n5051) );
  NAND2_X1 U5049 ( .A1(n6334), .A2(n6331), .ZN(n4735) );
  INV_X1 U5050 ( .A(n4577), .ZN(n6126) );
  AND2_X2 U5051 ( .A1(n5836), .A2(n5787), .ZN(n5851) );
  INV_X1 U5052 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n5787) );
  AND2_X1 U5053 ( .A1(n5597), .A2(n5583), .ZN(n5595) );
  INV_X1 U5054 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n4988) );
  OAI21_X1 U5055 ( .B1(n5496), .B2(n5495), .A(n5494), .ZN(n5510) );
  INV_X1 U5056 ( .A(n5892), .ZN(n6175) );
  INV_X1 U5057 ( .A(n6076), .ZN(n6138) );
  NOR2_X1 U5058 ( .A1(n4712), .A2(n4711), .ZN(n4709) );
  AND2_X1 U5059 ( .A1(n4918), .A2(n10142), .ZN(n4917) );
  INV_X1 U5060 ( .A(n9035), .ZN(n4667) );
  AOI21_X1 U5061 ( .B1(n9040), .B2(n9041), .A(n4472), .ZN(n9045) );
  NAND2_X1 U5062 ( .A1(n9497), .A2(n4473), .ZN(n4472) );
  INV_X1 U5063 ( .A(n9048), .ZN(n4697) );
  NOR2_X1 U5064 ( .A1(n6116), .A2(n6115), .ZN(n4577) );
  NOR2_X1 U5065 ( .A1(n6009), .A2(n4868), .ZN(n4867) );
  INV_X1 U5066 ( .A(n6294), .ZN(n4868) );
  AND2_X1 U5067 ( .A1(n5721), .A2(n5720), .ZN(n5727) );
  OR2_X1 U5068 ( .A1(n5733), .A2(n5734), .ZN(n5726) );
  OAI21_X1 U5069 ( .B1(n6561), .B2(n4475), .A(n4474), .ZN(n5047) );
  NAND2_X1 U5070 ( .A1(n6561), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n4474) );
  NAND2_X1 U5071 ( .A1(n5025), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n4703) );
  OR2_X1 U5072 ( .A1(n4279), .A2(n5026), .ZN(n4704) );
  NOR2_X1 U5073 ( .A1(n8026), .A2(n4927), .ZN(n4926) );
  INV_X1 U5074 ( .A(n4929), .ZN(n4927) );
  NOR2_X1 U5075 ( .A1(n4658), .A2(n6232), .ZN(n4657) );
  AND2_X1 U5076 ( .A1(n4291), .A2(n4446), .ZN(n6224) );
  AND2_X1 U5077 ( .A1(n4556), .A2(n4579), .ZN(n4554) );
  NAND2_X1 U5078 ( .A1(n4909), .A2(n4907), .ZN(n4576) );
  NAND2_X1 U5079 ( .A1(n8237), .A2(n6338), .ZN(n4907) );
  NAND2_X1 U5080 ( .A1(n4369), .A2(n6334), .ZN(n4734) );
  NAND2_X1 U5081 ( .A1(n4838), .A2(n6331), .ZN(n4736) );
  NAND2_X1 U5082 ( .A1(n6104), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n6116) );
  INV_X1 U5083 ( .A(n6105), .ZN(n6104) );
  NAND2_X1 U5084 ( .A1(n4888), .A2(n4886), .ZN(n4892) );
  NOR2_X1 U5085 ( .A1(n8307), .A2(n4887), .ZN(n4886) );
  INV_X1 U5086 ( .A(n6320), .ZN(n4887) );
  AOI21_X1 U5087 ( .B1(n4312), .B2(n4720), .A(n4362), .ZN(n4716) );
  OAI21_X1 U5088 ( .B1(n7213), .B2(n4904), .A(n4902), .ZN(n6309) );
  AND2_X1 U5089 ( .A1(n8169), .A2(n4903), .ZN(n4902) );
  NAND2_X1 U5090 ( .A1(n6039), .A2(n5848), .ZN(n4903) );
  NAND2_X1 U5091 ( .A1(n8366), .A2(n6299), .ZN(n8381) );
  AND2_X1 U5092 ( .A1(n6520), .A2(n6519), .ZN(n7015) );
  OR2_X1 U5093 ( .A1(n10030), .A2(P2_D_REG_1__SCAN_IN), .ZN(n6520) );
  OR2_X1 U5094 ( .A1(n10030), .A2(n6530), .ZN(n7013) );
  INV_X1 U5095 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n6049) );
  AND2_X1 U5096 ( .A1(n9115), .A2(n4612), .ZN(n9081) );
  NAND2_X1 U5097 ( .A1(n9249), .A2(n9250), .ZN(n9251) );
  INV_X1 U5098 ( .A(n4784), .ZN(n9248) );
  INV_X1 U5099 ( .A(n4497), .ZN(n4496) );
  OAI21_X1 U5100 ( .B1(n4499), .B2(n4498), .A(n4848), .ZN(n4497) );
  NAND2_X1 U5101 ( .A1(n4516), .A2(n4518), .ZN(n4514) );
  INV_X1 U5102 ( .A(n4516), .ZN(n4515) );
  NAND2_X1 U5103 ( .A1(n7868), .A2(n5637), .ZN(n4530) );
  INV_X1 U5104 ( .A(n4859), .ZN(n4858) );
  OAI21_X1 U5105 ( .B1(n9101), .B2(n4860), .A(n5259), .ZN(n4859) );
  NAND2_X1 U5106 ( .A1(n4313), .A2(n4335), .ZN(n4508) );
  NAND2_X1 U5107 ( .A1(n9944), .A2(n8944), .ZN(n9012) );
  NAND2_X1 U5108 ( .A1(n9227), .A2(n9927), .ZN(n7412) );
  INV_X1 U5109 ( .A(n9758), .ZN(n5009) );
  INV_X1 U5110 ( .A(n9761), .ZN(n5005) );
  NAND2_X1 U5111 ( .A1(n5641), .A2(n4342), .ZN(n9461) );
  NAND2_X1 U5112 ( .A1(n5727), .A2(n5726), .ZN(n5741) );
  NAND2_X1 U5113 ( .A1(n4616), .A2(n4614), .ZN(n5598) );
  AOI21_X1 U5114 ( .B1(n4617), .B2(n4620), .A(n4615), .ZN(n4614) );
  AND2_X1 U5115 ( .A1(n5578), .A2(n5564), .ZN(n5576) );
  INV_X1 U5116 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n4987) );
  AND2_X1 U5117 ( .A1(n5530), .A2(n5516), .ZN(n5528) );
  OAI21_X1 U5118 ( .B1(n4895), .B2(n4634), .A(n4632), .ZN(n5470) );
  INV_X1 U5119 ( .A(n4635), .ZN(n4634) );
  AND2_X1 U5120 ( .A1(n5467), .A2(n4633), .ZN(n4632) );
  AND2_X1 U5121 ( .A1(n5469), .A2(n5432), .ZN(n5466) );
  AOI21_X1 U5122 ( .B1(n4975), .B2(n4899), .A(n4898), .ZN(n4897) );
  INV_X1 U5123 ( .A(n5354), .ZN(n4899) );
  INV_X1 U5124 ( .A(n5376), .ZN(n4898) );
  NAND2_X1 U5125 ( .A1(n4895), .A2(n4894), .ZN(n4893) );
  AOI21_X1 U5126 ( .B1(n4974), .B2(n4884), .A(n4883), .ZN(n4882) );
  INV_X1 U5127 ( .A(n5290), .ZN(n4884) );
  INV_X1 U5128 ( .A(n5317), .ZN(n4883) );
  AOI21_X1 U5129 ( .B1(n5050), .B2(n4701), .A(n4855), .ZN(n4854) );
  INV_X1 U5130 ( .A(n5143), .ZN(n4855) );
  NAND2_X1 U5131 ( .A1(n7213), .A2(n6182), .ZN(n4906) );
  OR2_X1 U5132 ( .A1(n6223), .A2(n8392), .ZN(n7034) );
  AND2_X1 U5133 ( .A1(n6152), .A2(n6151), .ZN(n8182) );
  OR2_X1 U5134 ( .A1(n8210), .A2(n6076), .ZN(n6152) );
  INV_X1 U5135 ( .A(n8429), .ZN(n8159) );
  OR2_X1 U5136 ( .A1(n8437), .A2(n8182), .ZN(n8184) );
  NAND2_X1 U5137 ( .A1(n6172), .A2(n6160), .ZN(n8186) );
  OR2_X1 U5138 ( .A1(n8154), .A2(n8202), .ZN(n6160) );
  XNOR2_X1 U5139 ( .A(n6145), .B(P2_REG3_REG_27__SCAN_IN), .ZN(n8222) );
  AND2_X1 U5140 ( .A1(n6123), .A2(n6122), .ZN(n8273) );
  NOR2_X1 U5141 ( .A1(n8270), .A2(n4971), .ZN(n4970) );
  INV_X1 U5142 ( .A(n4977), .ZN(n4971) );
  NAND2_X1 U5143 ( .A1(n6071), .A2(n4889), .ZN(n4888) );
  NOR2_X1 U5144 ( .A1(n8318), .A2(n4890), .ZN(n4889) );
  INV_X1 U5145 ( .A(n6319), .ZN(n4890) );
  INV_X1 U5146 ( .A(n4713), .ZN(n4712) );
  OAI21_X1 U5147 ( .B1(n4714), .B2(n8326), .A(n4953), .ZN(n4713) );
  OR2_X1 U5148 ( .A1(n8174), .A2(n8175), .ZN(n4953) );
  NOR2_X1 U5149 ( .A1(n8490), .A2(n4771), .ZN(n4769) );
  NAND2_X1 U5150 ( .A1(n6665), .A2(n6371), .ZN(n8407) );
  INV_X1 U5151 ( .A(n8305), .ZN(n10017) );
  OR2_X1 U5152 ( .A1(n7374), .A2(n6518), .ZN(n7068) );
  NAND2_X1 U5153 ( .A1(n6133), .A2(n6132), .ZN(n8441) );
  INV_X1 U5154 ( .A(n5796), .ZN(n4972) );
  AND2_X1 U5155 ( .A1(n4649), .A2(n6014), .ZN(n4646) );
  NAND2_X1 U5156 ( .A1(n8900), .A2(n8901), .ZN(n4812) );
  INV_X1 U5157 ( .A(n5166), .ZN(n5399) );
  NAND2_X1 U5158 ( .A1(n8892), .A2(n8890), .ZN(n4816) );
  INV_X1 U5159 ( .A(n4812), .ZN(n4811) );
  AND2_X1 U5160 ( .A1(n9118), .A2(n4480), .ZN(n9121) );
  CLKBUF_X1 U5161 ( .A(n5021), .Z(n5022) );
  XNOR2_X1 U5162 ( .A(n9251), .B(n9264), .ZN(n9829) );
  NOR2_X1 U5163 ( .A1(n9264), .A2(n9251), .ZN(n9252) );
  INV_X1 U5164 ( .A(n4942), .ZN(n4940) );
  NAND2_X1 U5165 ( .A1(n9761), .A2(n9758), .ZN(n5523) );
  NAND2_X1 U5166 ( .A1(n4495), .A2(n4500), .ZN(n9397) );
  OR2_X1 U5167 ( .A1(n9471), .A2(n4501), .ZN(n4495) );
  NAND2_X1 U5169 ( .A1(n7484), .A2(n9147), .ZN(n5634) );
  AND2_X2 U5170 ( .A1(n5009), .A2(n5005), .ZN(n5652) );
  AND2_X1 U5171 ( .A1(n4300), .A2(n9121), .ZN(n9562) );
  OR2_X1 U5172 ( .A1(n6763), .A2(n5690), .ZN(n6700) );
  INV_X1 U5173 ( .A(n9562), .ZN(n9518) );
  AND2_X1 U5174 ( .A1(n5649), .A2(n5648), .ZN(n9515) );
  AND2_X1 U5175 ( .A1(n5677), .A2(n4430), .ZN(n9878) );
  NOR2_X1 U5176 ( .A1(n7724), .A2(n7784), .ZN(n4429) );
  INV_X1 U5177 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n4992) );
  NOR2_X1 U5178 ( .A1(n5746), .A2(n9535), .ZN(n9289) );
  NAND2_X1 U5179 ( .A1(n4939), .A2(n9115), .ZN(n4938) );
  NOR2_X1 U5180 ( .A1(n4308), .A2(n4644), .ZN(n4643) );
  AOI21_X1 U5181 ( .B1(n4415), .B2(n4337), .A(n4832), .ZN(n4831) );
  NAND2_X1 U5182 ( .A1(n7227), .A2(n6269), .ZN(n4832) );
  AND2_X1 U5183 ( .A1(n6304), .A2(n6301), .ZN(n4824) );
  NAND2_X1 U5184 ( .A1(n4414), .A2(n4412), .ZN(n6306) );
  NAND2_X1 U5185 ( .A1(n4413), .A2(n6349), .ZN(n4412) );
  INV_X1 U5186 ( .A(n6304), .ZN(n4413) );
  AOI21_X1 U5187 ( .B1(n4682), .B2(n9022), .A(n4681), .ZN(n9023) );
  OR2_X1 U5188 ( .A1(n9020), .A2(n9021), .ZN(n4681) );
  NAND2_X1 U5189 ( .A1(n9013), .A2(n4683), .ZN(n4682) );
  AOI21_X1 U5190 ( .B1(n9009), .B2(n9147), .A(n9008), .ZN(n9027) );
  INV_X1 U5191 ( .A(n9149), .ZN(n4665) );
  AOI21_X1 U5192 ( .B1(n8288), .B2(n6349), .A(n4841), .ZN(n4840) );
  NAND2_X1 U5193 ( .A1(n4471), .A2(n4699), .ZN(n4694) );
  INV_X1 U5194 ( .A(n9045), .ZN(n4471) );
  NAND2_X1 U5195 ( .A1(n4690), .A2(n9170), .ZN(n4689) );
  INV_X1 U5196 ( .A(n4692), .ZN(n4690) );
  AOI21_X1 U5197 ( .B1(n4693), .B2(n4696), .A(n9169), .ZN(n4692) );
  INV_X1 U5198 ( .A(n4695), .ZN(n4693) );
  NOR2_X1 U5199 ( .A1(n9098), .A2(n9100), .ZN(n4459) );
  AND2_X1 U5200 ( .A1(n6338), .A2(n4638), .ZN(n4637) );
  OR2_X1 U5201 ( .A1(n6338), .A2(n6347), .ZN(n4835) );
  AND2_X1 U5202 ( .A1(n4879), .A2(n5265), .ZN(n4878) );
  NOR2_X1 U5203 ( .A1(n4588), .A2(n6062), .ZN(n4587) );
  INV_X1 U5204 ( .A(n6063), .ZN(n6061) );
  NAND2_X1 U5205 ( .A1(n4678), .A2(n4677), .ZN(n4676) );
  AOI21_X1 U5206 ( .B1(n9054), .B2(n4671), .A(n9067), .ZN(n4677) );
  AND2_X1 U5207 ( .A1(n9336), .A2(n4674), .ZN(n4673) );
  NAND2_X1 U5208 ( .A1(n4522), .A2(n4671), .ZN(n4674) );
  NOR2_X1 U5209 ( .A1(n9323), .A2(n4461), .ZN(n4460) );
  INV_X1 U5210 ( .A(n9346), .ZN(n4462) );
  AND2_X1 U5211 ( .A1(n4623), .A2(n5576), .ZN(n4622) );
  NAND2_X1 U5212 ( .A1(n5559), .A2(n5558), .ZN(n4623) );
  AND2_X1 U5213 ( .A1(n4631), .A2(n5528), .ZN(n4630) );
  NAND2_X1 U5214 ( .A1(n5509), .A2(n5508), .ZN(n4631) );
  NAND2_X1 U5215 ( .A1(n4635), .A2(n4896), .ZN(n4633) );
  AND2_X1 U5216 ( .A1(n5466), .A2(n5465), .ZN(n5467) );
  INV_X1 U5217 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n5318) );
  AND2_X1 U5218 ( .A1(n5052), .A2(n4700), .ZN(n4428) );
  NAND2_X1 U5219 ( .A1(n5055), .A2(n5054), .ZN(n5058) );
  OR2_X1 U5220 ( .A1(n6561), .A2(n5053), .ZN(n5055) );
  AND2_X1 U5221 ( .A1(n6477), .A2(n6470), .ZN(n4912) );
  AOI21_X1 U5222 ( .B1(n4602), .B2(n4604), .A(n4601), .ZN(n4600) );
  INV_X1 U5223 ( .A(n7937), .ZN(n4601) );
  NAND2_X1 U5224 ( .A1(n7991), .A2(n7992), .ZN(n4915) );
  NOR2_X1 U5225 ( .A1(n6161), .A2(n8186), .ZN(n4579) );
  AND2_X1 U5226 ( .A1(n4574), .A2(n6222), .ZN(n4556) );
  NAND2_X1 U5227 ( .A1(n4575), .A2(n6131), .ZN(n4574) );
  INV_X1 U5228 ( .A(n4576), .ZN(n4575) );
  NOR2_X1 U5229 ( .A1(n8174), .A2(n4955), .ZN(n4954) );
  INV_X1 U5230 ( .A(n4982), .ZN(n4955) );
  NAND2_X1 U5231 ( .A1(n4968), .A2(n4969), .ZN(n4965) );
  INV_X1 U5232 ( .A(n4867), .ZN(n4866) );
  INV_X1 U5233 ( .A(n6302), .ZN(n4451) );
  NOR2_X1 U5234 ( .A1(n4793), .A2(n7737), .ZN(n4791) );
  NAND2_X1 U5235 ( .A1(n10078), .A2(n4794), .ZN(n4793) );
  AOI21_X1 U5236 ( .B1(n6278), .B2(n4874), .A(n4873), .ZN(n4872) );
  INV_X1 U5237 ( .A(n6272), .ZN(n4874) );
  INV_X1 U5238 ( .A(n7028), .ZN(n4958) );
  AND2_X1 U5239 ( .A1(n6383), .A2(n10041), .ZN(n6245) );
  INV_X1 U5240 ( .A(n10029), .ZN(n6518) );
  NOR2_X1 U5241 ( .A1(n8562), .A2(n4799), .ZN(n4798) );
  NAND2_X1 U5242 ( .A1(n8563), .A2(n4802), .ZN(n4801) );
  INV_X1 U5243 ( .A(n7647), .ZN(n4802) );
  NOR2_X1 U5244 ( .A1(n9081), .A2(n9000), .ZN(n9192) );
  AND2_X1 U5245 ( .A1(n6628), .A2(n6627), .ZN(n6899) );
  CLKBUF_X1 U5246 ( .A(n5297), .Z(n5298) );
  OR2_X1 U5247 ( .A1(n9815), .A2(n4785), .ZN(n4784) );
  AND2_X1 U5248 ( .A1(n9820), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n4785) );
  AND2_X1 U5249 ( .A1(n9276), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n4767) );
  NOR2_X1 U5250 ( .A1(n9257), .A2(n4766), .ZN(n4565) );
  NOR2_X1 U5251 ( .A1(n9352), .A2(n9369), .ZN(n4946) );
  NAND2_X1 U5252 ( .A1(n4848), .A2(n4851), .ZN(n4846) );
  NAND2_X1 U5253 ( .A1(n9172), .A2(n9085), .ZN(n4528) );
  AOI21_X1 U5254 ( .B1(n5642), .B2(n4749), .A(n4748), .ZN(n4747) );
  AND2_X1 U5255 ( .A1(n4745), .A2(n4539), .ZN(n4538) );
  NOR2_X1 U5256 ( .A1(n9419), .A2(n4746), .ZN(n4745) );
  NAND2_X1 U5257 ( .A1(n9454), .A2(n4540), .ZN(n4539) );
  INV_X1 U5258 ( .A(n9058), .ZN(n4746) );
  NAND2_X1 U5259 ( .A1(n4368), .A2(n4311), .ZN(n4516) );
  NAND2_X1 U5260 ( .A1(n4329), .A2(n5315), .ZN(n4519) );
  INV_X1 U5261 ( .A(n4508), .ZN(n4505) );
  AND2_X1 U5262 ( .A1(n4858), .A2(n4334), .ZN(n4507) );
  AOI21_X1 U5263 ( .B1(n4858), .B2(n4860), .A(n4357), .ZN(n4857) );
  NOR2_X1 U5264 ( .A1(n5766), .A2(n6557), .ZN(n6707) );
  AND2_X1 U5265 ( .A1(n5727), .A2(n5722), .ZN(n5723) );
  NAND2_X1 U5266 ( .A1(n5718), .A2(n5716), .ZN(n5733) );
  INV_X1 U5267 ( .A(n4622), .ZN(n4620) );
  AOI21_X1 U5268 ( .B1(n4622), .B2(n4619), .A(n4618), .ZN(n4617) );
  INV_X1 U5269 ( .A(n5578), .ZN(n4618) );
  INV_X1 U5270 ( .A(n5558), .ZN(n4619) );
  NAND2_X1 U5271 ( .A1(n5543), .A2(n5542), .ZN(n5560) );
  NAND2_X1 U5272 ( .A1(n4624), .A2(n4316), .ZN(n5543) );
  AOI21_X1 U5273 ( .B1(n4630), .B2(n4627), .A(n4626), .ZN(n4625) );
  INV_X1 U5274 ( .A(n5530), .ZN(n4626) );
  INV_X1 U5275 ( .A(n5508), .ZN(n4627) );
  OR2_X1 U5276 ( .A1(n5510), .A2(n4628), .ZN(n4624) );
  INV_X1 U5277 ( .A(n4630), .ZN(n4628) );
  OR2_X1 U5278 ( .A1(n5425), .A2(n5424), .ZN(n5447) );
  OR2_X1 U5279 ( .A1(n5415), .A2(n5425), .ZN(n5445) );
  NAND2_X1 U5280 ( .A1(n4893), .A2(n4897), .ZN(n5446) );
  INV_X1 U5281 ( .A(n5355), .ZN(n4901) );
  NAND2_X1 U5282 ( .A1(n5337), .A2(n5336), .ZN(n5354) );
  NAND2_X1 U5283 ( .A1(n4549), .A2(n4548), .ZN(n4880) );
  AND2_X1 U5284 ( .A1(n4881), .A2(n5270), .ZN(n4548) );
  NOR2_X1 U5285 ( .A1(n5291), .A2(n4885), .ZN(n4881) );
  INV_X1 U5286 ( .A(n4974), .ZN(n4885) );
  NAND2_X1 U5287 ( .A1(n5272), .A2(n5271), .ZN(n5290) );
  NAND2_X1 U5288 ( .A1(n4549), .A2(n5270), .ZN(n5292) );
  NAND2_X1 U5289 ( .A1(n5060), .A2(n4879), .ZN(n5267) );
  INV_X1 U5290 ( .A(n5127), .ZN(n4547) );
  NAND2_X1 U5291 ( .A1(n4458), .A2(n4457), .ZN(n4796) );
  INV_X1 U5292 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n4458) );
  XNOR2_X1 U5293 ( .A(n5044), .B(n4702), .ZN(n5043) );
  INV_X1 U5294 ( .A(SI_3_), .ZN(n4702) );
  INV_X1 U5295 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4844) );
  NOR2_X1 U5296 ( .A1(n4914), .A2(n4598), .ZN(n4597) );
  NAND2_X1 U5297 ( .A1(n8392), .A2(n4445), .ZN(n6382) );
  NOR2_X1 U5298 ( .A1(n6223), .A2(n4446), .ZN(n4445) );
  NAND2_X1 U5299 ( .A1(n4654), .A2(n6349), .ZN(n4650) );
  OR3_X1 U5300 ( .A1(n7722), .A2(n7819), .A3(n7785), .ZN(n6718) );
  AND2_X1 U5302 ( .A1(n6145), .A2(n6127), .ZN(n8233) );
  NAND2_X1 U5303 ( .A1(n6334), .A2(n6336), .ZN(n8254) );
  AOI21_X1 U5304 ( .B1(n8293), .B2(n6138), .A(n6100), .ZN(n8272) );
  NAND2_X1 U5305 ( .A1(n8269), .A2(n8270), .ZN(n8275) );
  NAND2_X1 U5306 ( .A1(n8327), .A2(n8326), .ZN(n8325) );
  AOI21_X1 U5307 ( .B1(n4309), .B2(n4719), .A(n4366), .ZN(n4718) );
  INV_X1 U5308 ( .A(n4309), .ZN(n4720) );
  AND2_X1 U5310 ( .A1(n4583), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n4582) );
  OR2_X1 U5311 ( .A1(n8490), .A2(n8408), .ZN(n8366) );
  AND2_X1 U5312 ( .A1(n8368), .A2(n8366), .ZN(n6048) );
  AND2_X1 U5313 ( .A1(n7795), .A2(n4376), .ZN(n8360) );
  NAND2_X1 U5314 ( .A1(n4722), .A2(n8408), .ZN(n4721) );
  AND2_X1 U5315 ( .A1(n6315), .A2(n6309), .ZN(n8368) );
  NAND2_X1 U5316 ( .A1(n4454), .A2(n8381), .ZN(n8380) );
  NAND2_X1 U5317 ( .A1(n8384), .A2(n4719), .ZN(n8383) );
  OR2_X1 U5318 ( .A1(n6004), .A2(n8035), .ZN(n6019) );
  OR2_X1 U5319 ( .A1(n5974), .A2(n7996), .ZN(n5991) );
  AND2_X2 U5320 ( .A1(n7775), .A2(n7777), .ZN(n7795) );
  INV_X1 U5321 ( .A(n4865), .ZN(n4869) );
  AND3_X1 U5322 ( .A1(n5995), .A2(n5994), .A3(n5993), .ZN(n7734) );
  NAND2_X1 U5323 ( .A1(n7392), .A2(n6278), .ZN(n7546) );
  XNOR2_X1 U5324 ( .A(n7389), .B(n8063), .ZN(n7227) );
  OR2_X1 U5325 ( .A1(n6384), .A2(n10090), .ZN(n7515) );
  AND2_X1 U5326 ( .A1(n6665), .A2(n6545), .ZN(n7371) );
  AND2_X1 U5327 ( .A1(n4776), .A2(n10019), .ZN(n4773) );
  NAND2_X1 U5328 ( .A1(n6125), .A2(n6124), .ZN(n8447) );
  INV_X1 U5329 ( .A(n10077), .ZN(n10063) );
  NAND2_X1 U5330 ( .A1(n6517), .A2(n10031), .ZN(n7374) );
  OR2_X1 U5331 ( .A1(n10030), .A2(P2_D_REG_0__SCAN_IN), .ZN(n6517) );
  NOR2_X1 U5332 ( .A1(n7015), .A2(n7014), .ZN(n7070) );
  INV_X1 U5333 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5795) );
  NAND2_X1 U5334 ( .A1(n6197), .A2(n10238), .ZN(n6355) );
  NAND2_X1 U5335 ( .A1(n6355), .A2(n6198), .ZN(n6546) );
  OR2_X1 U5336 ( .A1(n6197), .A2(n10238), .ZN(n6198) );
  INV_X1 U5337 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n6195) );
  AND2_X1 U5338 ( .A1(n6168), .A2(n6049), .ZN(n4918) );
  NAND2_X1 U5339 ( .A1(n6050), .A2(n6049), .ZN(n4448) );
  INV_X1 U5340 ( .A(n4456), .ZN(n5919) );
  INV_X1 U5341 ( .A(n5863), .ZN(n5871) );
  NAND2_X1 U5342 ( .A1(n8878), .A2(n8576), .ZN(n8753) );
  XNOR2_X1 U5343 ( .A(n6989), .B(n4285), .ZN(n6998) );
  NAND2_X1 U5344 ( .A1(n8923), .A2(n8596), .ZN(n8821) );
  INV_X1 U5345 ( .A(n4810), .ZN(n4809) );
  OAI21_X1 U5346 ( .B1(n4813), .B2(n4811), .A(n8617), .ZN(n4810) );
  OR2_X1 U5347 ( .A1(n8846), .A2(n8845), .ZN(n8853) );
  AOI22_X1 U5348 ( .A1(n7073), .A2(n7292), .B1(P1_IR_REG_0__SCAN_IN), .B2(
        n8992), .ZN(n4432) );
  INV_X1 U5349 ( .A(n7253), .ZN(n4465) );
  NAND2_X1 U5350 ( .A1(n8753), .A2(n8754), .ZN(n8922) );
  AND4_X1 U5351 ( .A1(n5158), .A2(n5157), .A3(n5156), .A4(n5155), .ZN(n7607)
         );
  INV_X1 U5352 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n4744) );
  OR2_X1 U5353 ( .A1(n6653), .A2(n6654), .ZN(n4560) );
  NOR2_X1 U5354 ( .A1(n6874), .A2(n6875), .ZN(n6882) );
  OR2_X1 U5355 ( .A1(n6882), .A2(n4783), .ZN(n4558) );
  AND2_X1 U5356 ( .A1(n6883), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n4783) );
  NAND2_X1 U5357 ( .A1(n4558), .A2(n4557), .ZN(n4782) );
  INV_X1 U5358 ( .A(n6884), .ZN(n4557) );
  OAI21_X1 U5359 ( .B1(n7245), .B2(P1_REG2_REG_11__SCAN_IN), .A(n7244), .ZN(
        n7246) );
  AND2_X1 U5360 ( .A1(n5303), .A2(n5302), .ZN(n5341) );
  OAI21_X1 U5361 ( .B1(n9829), .B2(n4570), .A(n4568), .ZN(n9840) );
  OR2_X1 U5362 ( .A1(n9841), .A2(n9828), .ZN(n4570) );
  INV_X1 U5363 ( .A(n9841), .ZN(n4569) );
  OR2_X1 U5364 ( .A1(n9829), .A2(n9828), .ZN(n4572) );
  NOR2_X1 U5365 ( .A1(n9851), .A2(n4399), .ZN(n9256) );
  NOR2_X1 U5366 ( .A1(n9270), .A2(n9269), .ZN(n9277) );
  OR2_X1 U5367 ( .A1(n9303), .A2(n9076), .ZN(n9185) );
  NAND2_X1 U5368 ( .A1(n9332), .A2(n9336), .ZN(n9331) );
  INV_X1 U5369 ( .A(n4527), .ZN(n4526) );
  NAND2_X1 U5370 ( .A1(n4307), .A2(n4349), .ZN(n4853) );
  NAND2_X1 U5371 ( .A1(n9461), .A2(n9160), .ZN(n9453) );
  NAND2_X1 U5372 ( .A1(n9453), .A2(n9454), .ZN(n9452) );
  OAI21_X1 U5373 ( .B1(n9479), .B2(n5392), .A(n5393), .ZN(n9471) );
  AND2_X1 U5374 ( .A1(n4310), .A2(n4948), .ZN(n4947) );
  INV_X1 U5375 ( .A(n9657), .ZN(n4948) );
  AND4_X1 U5376 ( .A1(n5353), .A2(n5352), .A3(n5351), .A4(n5350), .ZN(n9502)
         );
  AOI22_X1 U5377 ( .A1(n5638), .A2(n9559), .B1(n9036), .B2(n4530), .ZN(n9514)
         );
  NAND2_X1 U5378 ( .A1(n9565), .A2(n5289), .ZN(n9534) );
  AND4_X1 U5379 ( .A1(n5236), .A2(n5235), .A3(n5234), .A4(n5233), .ZN(n8581)
         );
  NAND2_X1 U5380 ( .A1(n4503), .A2(n4508), .ZN(n7498) );
  NAND2_X1 U5381 ( .A1(n7498), .A2(n9101), .ZN(n7497) );
  NAND2_X1 U5382 ( .A1(n7308), .A2(n4339), .ZN(n7484) );
  NAND2_X1 U5383 ( .A1(n7351), .A2(n5629), .ZN(n9136) );
  INV_X1 U5384 ( .A(n7353), .ZN(n7351) );
  AND2_X1 U5385 ( .A1(n5632), .A2(n5631), .ZN(n9134) );
  NAND2_X1 U5386 ( .A1(n4367), .A2(n5629), .ZN(n5632) );
  AND2_X1 U5387 ( .A1(n9017), .A2(n9133), .ZN(n7309) );
  OAI211_X1 U5388 ( .C1(n6563), .C2(n5166), .A(n5165), .B(n5164), .ZN(n7599)
         );
  OR2_X1 U5389 ( .A1(n6763), .A2(n5663), .ZN(n9535) );
  NAND2_X1 U5390 ( .A1(n5118), .A2(n7352), .ZN(n9090) );
  INV_X1 U5391 ( .A(n9515), .ZN(n9563) );
  NAND2_X1 U5392 ( .A1(n4680), .A2(n4679), .ZN(n7277) );
  INV_X1 U5393 ( .A(n9093), .ZN(n4679) );
  NAND2_X1 U5394 ( .A1(n5743), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n5077) );
  INV_X1 U5395 ( .A(n4453), .ZN(n7297) );
  AND2_X1 U5396 ( .A1(n9121), .A2(n5697), .ZN(n7159) );
  NAND2_X1 U5397 ( .A1(n5586), .A2(n5585), .ZN(n9603) );
  NAND2_X1 U5398 ( .A1(n5455), .A2(n5454), .ZN(n9651) );
  NAND2_X1 U5399 ( .A1(n5641), .A2(n9046), .ZN(n9463) );
  AND2_X1 U5400 ( .A1(n5692), .A2(n5691), .ZN(n6699) );
  NAND2_X1 U5401 ( .A1(n4997), .A2(n4760), .ZN(n4759) );
  AND2_X1 U5402 ( .A1(n4999), .A2(n4761), .ZN(n4760) );
  INV_X1 U5403 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n4761) );
  XNOR2_X1 U5404 ( .A(n5741), .B(n5740), .ZN(n7894) );
  INV_X1 U5405 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5668) );
  NAND2_X1 U5406 ( .A1(n5669), .A2(n5668), .ZN(n5674) );
  XNOR2_X1 U5407 ( .A(n5560), .B(n5559), .ZN(n7781) );
  INV_X1 U5408 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5671) );
  XNOR2_X1 U5409 ( .A(n5694), .B(n10141), .ZN(n8988) );
  NAND2_X1 U5410 ( .A1(n4629), .A2(n5508), .ZN(n5529) );
  OR2_X1 U5411 ( .A1(n5510), .A2(n5509), .ZN(n4629) );
  XNOR2_X1 U5412 ( .A(n5433), .B(n5466), .ZN(n7268) );
  NAND2_X1 U5413 ( .A1(n4893), .A2(n4635), .ZN(n5468) );
  NAND2_X1 U5414 ( .A1(n5397), .A2(n5423), .ZN(n5398) );
  NAND2_X1 U5415 ( .A1(n4893), .A2(n4314), .ZN(n5397) );
  XNOR2_X1 U5416 ( .A(n5292), .B(n5291), .ZN(n6589) );
  INV_X1 U5417 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n5177) );
  NAND2_X1 U5418 ( .A1(n4796), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5129) );
  NOR2_X1 U5419 ( .A1(n9780), .A2(n9779), .ZN(n9781) );
  NAND2_X1 U5420 ( .A1(n9784), .A2(n9785), .ZN(n9786) );
  NAND2_X1 U5421 ( .A1(n7204), .A2(n6410), .ZN(n7063) );
  AOI21_X1 U5422 ( .B1(n4923), .B2(n4925), .A(n4921), .ZN(n4920) );
  INV_X1 U5423 ( .A(n4923), .ZN(n4922) );
  INV_X1 U5424 ( .A(n7897), .ZN(n4921) );
  INV_X1 U5425 ( .A(n8317), .ZN(n8471) );
  NAND2_X1 U5426 ( .A1(n6103), .A2(n6102), .ZN(n8456) );
  AND2_X1 U5427 ( .A1(n6082), .A2(n6081), .ZN(n8173) );
  INV_X1 U5428 ( .A(n8330), .ZN(n8476) );
  AND2_X1 U5429 ( .A1(n6090), .A2(n6089), .ZN(n8009) );
  NOR2_X1 U5430 ( .A1(n6544), .A2(n6545), .ZN(n8005) );
  INV_X1 U5431 ( .A(n6544), .ZN(n6534) );
  NAND2_X1 U5432 ( .A1(n6917), .A2(n10063), .ZN(n8032) );
  NOR2_X1 U5433 ( .A1(n8024), .A2(n8044), .ZN(n4606) );
  NAND2_X1 U5434 ( .A1(n8025), .A2(n8026), .ZN(n4608) );
  AND2_X1 U5435 ( .A1(n8005), .A2(n8370), .ZN(n8033) );
  AND3_X1 U5436 ( .A1(n6023), .A2(n6022), .A3(n6021), .ZN(n8042) );
  OAI22_X1 U5437 ( .A1(n8185), .A2(n6181), .B1(n6180), .B2(n6348), .ZN(n4578)
         );
  NAND2_X1 U5438 ( .A1(n6112), .A2(n6111), .ZN(n8291) );
  OR2_X1 U5439 ( .A1(n7977), .A2(n6076), .ZN(n6112) );
  INV_X1 U5440 ( .A(n8009), .ZN(n8320) );
  NAND2_X1 U5441 ( .A1(n6070), .A2(n6069), .ZN(n8344) );
  OAI21_X1 U5442 ( .B1(n8354), .B2(n6076), .A(n6058), .ZN(n8373) );
  INV_X1 U5443 ( .A(n7734), .ZN(n8057) );
  NOR2_X1 U5444 ( .A1(n6010), .A2(n6011), .ZN(n6012) );
  AND2_X1 U5445 ( .A1(n6740), .A2(n6739), .ZN(n9999) );
  INV_X1 U5446 ( .A(n9999), .ZN(n9987) );
  NAND2_X1 U5447 ( .A1(n4777), .A2(n8423), .ZN(n4776) );
  INV_X1 U5448 ( .A(n4779), .ZN(n4777) );
  AND2_X1 U5449 ( .A1(n4779), .A2(n4656), .ZN(n4778) );
  NAND2_X1 U5450 ( .A1(n8204), .A2(n8184), .ZN(n4452) );
  AOI21_X1 U5451 ( .B1(n4305), .B2(n4963), .A(n4360), .ZN(n4961) );
  AOI21_X1 U5452 ( .B1(n8442), .B2(n8420), .A(n8228), .ZN(n4409) );
  INV_X1 U5453 ( .A(n4740), .ZN(n4410) );
  XNOR2_X1 U5454 ( .A(n4910), .B(n8225), .ZN(n4742) );
  AOI21_X1 U5455 ( .B1(n8226), .B2(n8372), .A(n4741), .ZN(n4740) );
  INV_X1 U5456 ( .A(n4911), .ZN(n8236) );
  OR2_X1 U5457 ( .A1(n4281), .A2(n7377), .ZN(n8379) );
  INV_X1 U5458 ( .A(n8192), .ZN(n8420) );
  OAI21_X1 U5459 ( .B1(n8786), .B2(n4976), .A(n8784), .ZN(n8787) );
  AND4_X1 U5460 ( .A1(n5214), .A2(n5213), .A3(n5212), .A4(n5211), .ZN(n8806)
         );
  NAND2_X1 U5461 ( .A1(n4483), .A2(n4482), .ZN(n4481) );
  INV_X1 U5462 ( .A(n8693), .ZN(n4482) );
  NAND2_X1 U5463 ( .A1(n5308), .A2(n5307), .ZN(n9681) );
  AND4_X1 U5464 ( .A1(n5286), .A2(n5285), .A3(n5284), .A4(n5283), .ZN(n9684)
         );
  INV_X1 U5465 ( .A(n9633), .ZN(n9217) );
  INV_X1 U5466 ( .A(n8830), .ZN(n9561) );
  INV_X1 U5467 ( .A(n8953), .ZN(n9225) );
  AND2_X1 U5468 ( .A1(n6624), .A2(n6623), .ZN(n6898) );
  AND2_X1 U5469 ( .A1(n4405), .A2(n4478), .ZN(n9287) );
  NAND2_X1 U5470 ( .A1(n4406), .A2(n9862), .ZN(n4405) );
  INV_X1 U5471 ( .A(n9286), .ZN(n4423) );
  INV_X1 U5472 ( .A(n9283), .ZN(n9285) );
  INV_X1 U5473 ( .A(n9299), .ZN(n9589) );
  NAND2_X1 U5474 ( .A1(n5770), .A2(n9541), .ZN(n5779) );
  INV_X1 U5475 ( .A(n9722), .ZN(n9388) );
  OR2_X1 U5476 ( .A1(n5771), .A2(n9119), .ZN(n9580) );
  XNOR2_X1 U5477 ( .A(n5611), .B(P1_IR_REG_19__SCAN_IN), .ZN(n9119) );
  NAND2_X1 U5478 ( .A1(n9884), .A2(n5768), .ZN(n9538) );
  NAND2_X1 U5479 ( .A1(n8544), .A2(n5742), .ZN(n5732) );
  INV_X1 U5480 ( .A(n5664), .ZN(n5665) );
  INV_X1 U5481 ( .A(n5770), .ZN(n5666) );
  INV_X1 U5482 ( .A(n9119), .ZN(n9418) );
  NOR2_X1 U5483 ( .A1(n10127), .A2(n4404), .ZN(n10126) );
  NOR2_X1 U5484 ( .A1(n10126), .A2(n10125), .ZN(n10124) );
  OAI21_X1 U5485 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10106), .ZN(n10292) );
  NAND2_X1 U5486 ( .A1(n6264), .A2(n4416), .ZN(n4415) );
  OAI21_X1 U5487 ( .B1(n4330), .B2(n4418), .A(n6290), .ZN(n6293) );
  NAND2_X1 U5488 ( .A1(n4642), .A2(n4643), .ZN(n4418) );
  AND2_X1 U5489 ( .A1(n9017), .A2(n9012), .ZN(n4683) );
  INV_X1 U5490 ( .A(n9547), .ZN(n4668) );
  NAND2_X1 U5491 ( .A1(n4670), .A2(n4669), .ZN(n9032) );
  NAND2_X1 U5492 ( .A1(n9026), .A2(n9077), .ZN(n4669) );
  INV_X1 U5493 ( .A(n9039), .ZN(n4473) );
  AOI21_X1 U5494 ( .B1(n4697), .B2(n4698), .A(n4364), .ZN(n4695) );
  NOR2_X1 U5495 ( .A1(n4839), .A2(n4838), .ZN(n4837) );
  INV_X1 U5496 ( .A(n6329), .ZN(n4839) );
  NAND2_X1 U5497 ( .A1(n9053), .A2(n9077), .ZN(n4678) );
  AND2_X1 U5498 ( .A1(n4691), .A2(n4689), .ZN(n9052) );
  NAND2_X1 U5499 ( .A1(n4331), .A2(n4315), .ZN(n9106) );
  NAND2_X1 U5500 ( .A1(n4909), .A2(n4835), .ZN(n4834) );
  NOR2_X1 U5501 ( .A1(n8167), .A2(n4967), .ZN(n4966) );
  INV_X1 U5502 ( .A(n7793), .ZN(n4967) );
  NOR2_X1 U5503 ( .A1(n4875), .A2(n4282), .ZN(n4871) );
  INV_X1 U5504 ( .A(n6278), .ZN(n4875) );
  INV_X1 U5505 ( .A(n7545), .ZN(n4873) );
  OR2_X1 U5506 ( .A1(n7216), .A2(n7135), .ZN(n6268) );
  INV_X1 U5507 ( .A(n4500), .ZN(n4498) );
  INV_X1 U5508 ( .A(n4501), .ZN(n4499) );
  INV_X1 U5509 ( .A(n9160), .ZN(n4540) );
  NOR2_X1 U5510 ( .A1(n9523), .A2(n9506), .ZN(n4950) );
  INV_X1 U5511 ( .A(n5595), .ZN(n4615) );
  NOR2_X1 U5512 ( .A1(n4996), .A2(n4935), .ZN(n4934) );
  AND2_X1 U5513 ( .A1(n5196), .A2(n5059), .ZN(n4879) );
  INV_X1 U5514 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4544) );
  AND2_X1 U5515 ( .A1(n6453), .A2(n6447), .ZN(n4914) );
  NOR2_X1 U5516 ( .A1(n6345), .A2(n6349), .ZN(n4652) );
  NAND2_X1 U5517 ( .A1(n4656), .A2(n4655), .ZN(n4654) );
  NAND2_X1 U5518 ( .A1(n4577), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n6145) );
  NAND2_X1 U5519 ( .A1(n6061), .A2(n4586), .ZN(n6105) );
  AND2_X1 U5520 ( .A1(n4587), .A2(n4402), .ZN(n4586) );
  NAND2_X1 U5521 ( .A1(n4790), .A2(n8285), .ZN(n4789) );
  INV_X1 U5522 ( .A(n8307), .ZN(n4711) );
  NAND2_X1 U5523 ( .A1(n6061), .A2(n4587), .ZN(n6096) );
  NOR2_X1 U5524 ( .A1(n8466), .A2(n8471), .ZN(n4790) );
  AND2_X1 U5525 ( .A1(n8471), .A2(n8334), .ZN(n8174) );
  NOR2_X1 U5526 ( .A1(n4585), .A2(n4584), .ZN(n4583) );
  INV_X1 U5527 ( .A(n6048), .ZN(n4732) );
  AOI21_X1 U5528 ( .B1(n6048), .B2(n8381), .A(n4731), .ZN(n4730) );
  INV_X1 U5529 ( .A(n6309), .ZN(n4731) );
  OR2_X1 U5530 ( .A1(n8494), .A2(n8042), .ZN(n6304) );
  NAND2_X1 U5531 ( .A1(n6018), .A2(n4583), .ZN(n6041) );
  INV_X1 U5532 ( .A(n6019), .ZN(n6018) );
  NAND2_X1 U5533 ( .A1(n7790), .A2(n7770), .ZN(n4865) );
  OR2_X1 U5534 ( .A1(n8519), .A2(n7735), .ZN(n6286) );
  NOR2_X1 U5535 ( .A1(n7406), .A2(n4581), .ZN(n4580) );
  INV_X1 U5536 ( .A(n5938), .ZN(n5937) );
  NAND2_X1 U5537 ( .A1(n5888), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5903) );
  INV_X1 U5538 ( .A(n5890), .ZN(n5888) );
  NAND2_X1 U5539 ( .A1(n4284), .A2(n4827), .ZN(n6241) );
  NAND2_X1 U5540 ( .A1(n5842), .A2(n5841), .ZN(n6247) );
  NAND2_X1 U5541 ( .A1(n6388), .A2(n10050), .ZN(n6252) );
  INV_X1 U5542 ( .A(SI_10_), .ZN(n10204) );
  NAND2_X1 U5543 ( .A1(n6196), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6197) );
  NAND2_X1 U5544 ( .A1(n6194), .A2(n6195), .ZN(n6196) );
  INV_X1 U5545 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n10238) );
  OAI21_X1 U5546 ( .B1(n5971), .B2(P2_IR_REG_12__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5983) );
  NAND2_X1 U5547 ( .A1(n4738), .A2(n4737), .ZN(n5971) );
  NOR2_X1 U5548 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n4737) );
  NOR2_X1 U5549 ( .A1(n5931), .A2(P2_IR_REG_9__SCAN_IN), .ZN(n4738) );
  NAND2_X1 U5550 ( .A1(n4456), .A2(n4455), .ZN(n5931) );
  INV_X1 U5551 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n4455) );
  NOR2_X1 U5552 ( .A1(n5910), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n4456) );
  OR2_X1 U5553 ( .A1(n5899), .A2(P2_IR_REG_6__SCAN_IN), .ZN(n5910) );
  AND2_X1 U5554 ( .A1(n5851), .A2(n5850), .ZN(n5863) );
  INV_X1 U5555 ( .A(n4277), .ZN(n8709) );
  AND2_X1 U5556 ( .A1(n5439), .A2(n5438), .ZN(n5473) );
  NOR2_X1 U5557 ( .A1(n5406), .A2(n5405), .ZN(n5439) );
  NAND2_X1 U5558 ( .A1(n4277), .A2(n6702), .ZN(n7253) );
  AND3_X1 U5559 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n5136) );
  NOR2_X1 U5560 ( .A1(n5324), .A2(n5323), .ZN(n5346) );
  NAND2_X1 U5561 ( .A1(n4675), .A2(n4673), .ZN(n4672) );
  NOR2_X1 U5562 ( .A1(n9200), .A2(n9125), .ZN(n9116) );
  AND2_X1 U5563 ( .A1(n9111), .A2(n4460), .ZN(n9112) );
  NAND2_X1 U5564 ( .A1(n4943), .A2(n9590), .ZN(n4942) );
  NAND2_X1 U5565 ( .A1(n4304), .A2(n9464), .ZN(n4501) );
  NOR2_X1 U5566 ( .A1(n5170), .A2(n5169), .ZN(n5006) );
  INV_X1 U5567 ( .A(n9004), .ZN(n9018) );
  AND3_X1 U5568 ( .A1(n7414), .A2(n7354), .A3(n9012), .ZN(n5629) );
  NAND2_X1 U5569 ( .A1(n7621), .A2(n9226), .ZN(n9004) );
  NAND2_X1 U5570 ( .A1(n7277), .A2(n4755), .ZN(n7353) );
  NOR2_X1 U5571 ( .A1(n5628), .A2(n4756), .ZN(n4755) );
  INV_X1 U5572 ( .A(n5627), .ZN(n4756) );
  AND2_X1 U5573 ( .A1(n5762), .A2(n5763), .ZN(n4861) );
  NAND2_X1 U5574 ( .A1(n9367), .A2(n9718), .ZN(n9351) );
  NAND2_X1 U5575 ( .A1(n4295), .A2(n4287), .ZN(n5166) );
  NAND2_X1 U5576 ( .A1(n5669), .A2(n5018), .ZN(n5019) );
  NAND2_X1 U5577 ( .A1(n5615), .A2(n5617), .ZN(n5693) );
  INV_X1 U5578 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n10141) );
  XNOR2_X1 U5579 ( .A(n5618), .B(P1_IR_REG_21__SCAN_IN), .ZN(n9198) );
  OR2_X1 U5580 ( .A1(n5428), .A2(n5427), .ZN(n5465) );
  AND2_X1 U5581 ( .A1(n5426), .A2(n5447), .ZN(n5427) );
  INV_X1 U5582 ( .A(n4897), .ZN(n4636) );
  OR2_X1 U5583 ( .A1(n5445), .A2(n5428), .ZN(n5417) );
  XNOR2_X1 U5584 ( .A(n5268), .B(SI_11_), .ZN(n5261) );
  INV_X1 U5585 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n10217) );
  OAI21_X1 U5586 ( .B1(n4856), .B2(n5159), .A(n4428), .ZN(n4546) );
  AND2_X1 U5587 ( .A1(n6509), .A2(n6507), .ZN(n7897) );
  AOI21_X1 U5588 ( .B1(n4926), .B2(n4924), .A(n6508), .ZN(n4923) );
  INV_X1 U5589 ( .A(n4371), .ZN(n4924) );
  INV_X1 U5590 ( .A(n4926), .ZN(n4925) );
  NAND2_X1 U5591 ( .A1(n4447), .A2(n4914), .ZN(n7803) );
  XNOR2_X1 U5592 ( .A(n8482), .B(n6494), .ZN(n6472) );
  OAI21_X1 U5593 ( .B1(n4912), .B2(n4604), .A(n6483), .ZN(n4603) );
  NAND2_X1 U5594 ( .A1(n4605), .A2(n6478), .ZN(n4604) );
  INV_X1 U5595 ( .A(n7984), .ZN(n4605) );
  XNOR2_X1 U5596 ( .A(n4283), .B(n7027), .ZN(n6398) );
  INV_X1 U5597 ( .A(n6398), .ZN(n7049) );
  INV_X1 U5598 ( .A(n7402), .ZN(n6428) );
  AND2_X1 U5599 ( .A1(n4591), .A2(n4590), .ZN(n4589) );
  AND2_X1 U5600 ( .A1(n4306), .A2(n7823), .ZN(n4591) );
  NAND2_X1 U5601 ( .A1(n4596), .A2(n4598), .ZN(n4590) );
  NAND2_X1 U5602 ( .A1(n7945), .A2(n4930), .ZN(n4929) );
  INV_X1 U5603 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n8035) );
  AND2_X1 U5604 ( .A1(n4654), .A2(n6344), .ZN(n6346) );
  AND2_X1 U5605 ( .A1(n8423), .A2(n6695), .ZN(n6345) );
  NAND2_X1 U5606 ( .A1(n4280), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n4829) );
  OR2_X1 U5607 ( .A1(n5892), .A2(n7527), .ZN(n4830) );
  AOI21_X1 U5608 ( .B1(n8092), .B2(n8091), .A(n8090), .ZN(n8089) );
  INV_X1 U5609 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n6723) );
  AOI21_X1 U5610 ( .B1(n6795), .B2(n6736), .A(n6735), .ZN(n6849) );
  OR2_X1 U5611 ( .A1(n6938), .A2(n6937), .ZN(n6962) );
  AOI21_X1 U5612 ( .B1(n8103), .B2(n6942), .A(n6941), .ZN(n7094) );
  OR2_X1 U5613 ( .A1(n6967), .A2(n6966), .ZN(n7122) );
  NAND2_X1 U5614 ( .A1(n7321), .A2(n4486), .ZN(n7691) );
  OR2_X1 U5615 ( .A1(n4290), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n4486) );
  AND2_X1 U5616 ( .A1(n8126), .A2(n8125), .ZN(n10007) );
  NAND2_X1 U5617 ( .A1(n10007), .A2(n10006), .ZN(n10004) );
  NAND2_X1 U5618 ( .A1(n10004), .A2(n4485), .ZN(n8130) );
  OR2_X1 U5619 ( .A1(n8127), .A2(n8128), .ZN(n4485) );
  NOR2_X1 U5620 ( .A1(n8159), .A2(n8154), .ZN(n4779) );
  NAND2_X1 U5621 ( .A1(n4552), .A2(n4579), .ZN(n4551) );
  NAND2_X1 U5622 ( .A1(n8238), .A2(n4554), .ZN(n4553) );
  INV_X1 U5623 ( .A(n4555), .ZN(n4552) );
  NAND2_X1 U5624 ( .A1(n4909), .A2(n8181), .ZN(n4962) );
  NAND2_X1 U5625 ( .A1(n8238), .A2(n4556), .ZN(n4550) );
  NOR2_X1 U5626 ( .A1(n8207), .A2(n4963), .ZN(n4708) );
  NOR2_X1 U5627 ( .A1(n8405), .A2(n8179), .ZN(n4741) );
  NAND2_X1 U5628 ( .A1(n4911), .A2(n6338), .ZN(n4910) );
  AND2_X1 U5629 ( .A1(n6126), .A2(n6117), .ZN(n8251) );
  OR2_X1 U5630 ( .A1(n8456), .A2(n8291), .ZN(n8177) );
  NOR2_X1 U5631 ( .A1(n8287), .A2(n8288), .ZN(n4891) );
  NOR2_X1 U5632 ( .A1(n8314), .A2(n4788), .ZN(n8299) );
  INV_X1 U5633 ( .A(n4790), .ZN(n4788) );
  NOR2_X1 U5634 ( .A1(n8314), .A2(n8471), .ZN(n8313) );
  OR2_X1 U5635 ( .A1(n6053), .A2(n10237), .ZN(n6063) );
  NAND2_X1 U5636 ( .A1(n6018), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n6030) );
  AND2_X1 U5637 ( .A1(n8165), .A2(n8164), .ZN(n8400) );
  NAND2_X1 U5638 ( .A1(n7795), .A2(n7800), .ZN(n8413) );
  NAND2_X1 U5639 ( .A1(n7794), .A2(n7793), .ZN(n8165) );
  NAND2_X1 U5640 ( .A1(n5989), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n6004) );
  INV_X1 U5641 ( .A(n5991), .ZN(n5989) );
  NAND2_X1 U5642 ( .A1(n4795), .A2(n7735), .ZN(n4726) );
  AND2_X1 U5643 ( .A1(n6291), .A2(n7770), .ZN(n7744) );
  NAND2_X1 U5644 ( .A1(n4363), .A2(n4792), .ZN(n7850) );
  AND4_X1 U5645 ( .A1(n5981), .A2(n5980), .A3(n5979), .A4(n5978), .ZN(n7845)
         );
  NAND2_X1 U5646 ( .A1(n4332), .A2(n4725), .ZN(n4723) );
  AND2_X1 U5647 ( .A1(n7539), .A2(n4728), .ZN(n4725) );
  NAND2_X1 U5648 ( .A1(n4792), .A2(n4791), .ZN(n7852) );
  NAND2_X1 U5649 ( .A1(n5937), .A2(n4580), .ZN(n5961) );
  NAND2_X1 U5650 ( .A1(n5937), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5949) );
  NOR2_X1 U5651 ( .A1(n7395), .A2(n4793), .ZN(n7712) );
  AND4_X1 U5652 ( .A1(n5954), .A2(n5953), .A3(n5952), .A4(n5951), .ZN(n7846)
         );
  NOR2_X1 U5653 ( .A1(n7395), .A2(n7885), .ZN(n7551) );
  INV_X1 U5654 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5924) );
  OR2_X1 U5655 ( .A1(n5925), .A2(n5924), .ZN(n5938) );
  NAND2_X1 U5656 ( .A1(n7226), .A2(n7227), .ZN(n4876) );
  INV_X1 U5657 ( .A(n4792), .ZN(n7395) );
  OR2_X1 U5658 ( .A1(n5903), .A2(n6723), .ZN(n5913) );
  INV_X1 U5659 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n6845) );
  OR2_X1 U5660 ( .A1(n5913), .A2(n6845), .ZN(n5925) );
  CLKBUF_X1 U5661 ( .A(n7225), .Z(n7226) );
  NOR2_X1 U5662 ( .A1(n7455), .A2(n7454), .ZN(n7453) );
  NOR2_X1 U5663 ( .A1(n7170), .A2(n4958), .ZN(n4957) );
  NAND2_X1 U5664 ( .A1(n4573), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5890) );
  INV_X1 U5665 ( .A(n5880), .ZN(n4573) );
  AND2_X1 U5666 ( .A1(n6205), .A2(n6240), .ZN(n4863) );
  NAND2_X1 U5667 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n5880) );
  NAND2_X1 U5668 ( .A1(n4765), .A2(n7027), .ZN(n7584) );
  INV_X1 U5669 ( .A(n10020), .ZN(n4765) );
  NAND2_X1 U5670 ( .A1(n10021), .A2(n10056), .ZN(n10020) );
  NOR2_X1 U5671 ( .A1(n7574), .A2(n5841), .ZN(n10021) );
  NAND2_X1 U5672 ( .A1(n7374), .A2(n7373), .ZN(n7380) );
  NAND2_X1 U5673 ( .A1(n6141), .A2(n6140), .ZN(n8437) );
  NAND2_X1 U5674 ( .A1(n6568), .A2(n6182), .ZN(n4729) );
  CLKBUF_X1 U5675 ( .A(n6381), .Z(n10089) );
  NAND2_X1 U5676 ( .A1(n6516), .A2(n6515), .ZN(n10030) );
  NAND2_X1 U5677 ( .A1(n5863), .A2(n4739), .ZN(n5873) );
  NAND2_X1 U5678 ( .A1(n5874), .A2(n5875), .ZN(n5899) );
  INV_X1 U5679 ( .A(n5873), .ZN(n5875) );
  NAND2_X1 U5680 ( .A1(n4803), .A2(n7647), .ZN(n8798) );
  NAND2_X1 U5681 ( .A1(n4449), .A2(n7645), .ZN(n4803) );
  INV_X1 U5682 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n5169) );
  OR2_X1 U5683 ( .A1(n8900), .A2(n8901), .ZN(n4813) );
  INV_X1 U5684 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n5323) );
  AND2_X1 U5685 ( .A1(n5502), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n5519) );
  INV_X1 U5686 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n5230) );
  AND2_X1 U5688 ( .A1(n5473), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n5502) );
  AND2_X1 U5689 ( .A1(n8637), .A2(n4806), .ZN(n4805) );
  NAND2_X1 U5690 ( .A1(n4809), .A2(n4811), .ZN(n4806) );
  NOR2_X1 U5691 ( .A1(n8812), .A2(n4815), .ZN(n4814) );
  INV_X1 U5692 ( .A(n8891), .ZN(n4815) );
  INV_X1 U5693 ( .A(n8865), .ZN(n4483) );
  AND2_X1 U5694 ( .A1(n8682), .A2(n8681), .ZN(n8813) );
  NAND2_X1 U5695 ( .A1(n5519), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n5533) );
  AND2_X1 U5696 ( .A1(n8575), .A2(n4801), .ZN(n4800) );
  OR2_X1 U5697 ( .A1(n5231), .A2(n5230), .ZN(n5253) );
  INV_X1 U5698 ( .A(n7077), .ZN(n4434) );
  CLKBUF_X1 U5699 ( .A(n7646), .Z(n4449) );
  AND2_X1 U5700 ( .A1(n7006), .A2(n7005), .ZN(n8978) );
  NAND2_X1 U5701 ( .A1(n9084), .A2(n4671), .ZN(n4688) );
  NOR2_X1 U5702 ( .A1(n9192), .A2(n9293), .ZN(n9079) );
  INV_X1 U5703 ( .A(n9195), .ZN(n9199) );
  AOI21_X1 U5704 ( .B1(n9192), .B2(n9191), .A(n9200), .ZN(n9193) );
  AND4_X1 U5705 ( .A1(n5656), .A2(n5655), .A3(n5654), .A4(n5653), .ZN(n9076)
         );
  NAND2_X1 U5706 ( .A1(n6639), .A2(n6638), .ZN(n6637) );
  AND2_X1 U5707 ( .A1(n4782), .A2(n4781), .ZN(n6925) );
  NAND2_X1 U5708 ( .A1(n6924), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n4781) );
  NAND2_X1 U5709 ( .A1(n6925), .A2(n6926), .ZN(n7244) );
  AND2_X1 U5710 ( .A1(n7671), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n4786) );
  AOI21_X1 U5711 ( .B1(n7680), .B2(n10253), .A(n7679), .ZN(n7683) );
  NOR2_X1 U5712 ( .A1(n9822), .A2(n9821), .ZN(n7679) );
  NOR2_X1 U5713 ( .A1(n7683), .A2(n7682), .ZN(n9261) );
  NOR2_X1 U5714 ( .A1(n9840), .A2(n4571), .ZN(n9853) );
  AND2_X1 U5715 ( .A1(n9844), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n4571) );
  AOI21_X1 U5716 ( .B1(n9279), .B2(n9278), .A(n9277), .ZN(n9280) );
  OAI21_X1 U5717 ( .B1(n9275), .B2(n4566), .A(n4563), .ZN(n9283) );
  OR2_X1 U5718 ( .A1(n4767), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n4566) );
  AOI21_X1 U5719 ( .B1(n4564), .B2(n4565), .A(n4400), .ZN(n4563) );
  INV_X1 U5720 ( .A(n4941), .ZN(n4939) );
  OR2_X1 U5721 ( .A1(n9319), .A2(n9293), .ZN(n4937) );
  NOR2_X1 U5722 ( .A1(n8999), .A2(n4942), .ZN(n4941) );
  NAND2_X1 U5723 ( .A1(n9367), .A2(n4944), .ZN(n9339) );
  AND2_X1 U5724 ( .A1(n4946), .A2(n4945), .ZN(n4944) );
  OAI22_X1 U5725 ( .A1(n9335), .A2(n5575), .B1(n9349), .B2(n4945), .ZN(n9318)
         );
  AOI21_X1 U5726 ( .B1(n4850), .B2(n4849), .A(n4356), .ZN(n4848) );
  INV_X1 U5727 ( .A(n4325), .ZN(n4849) );
  NAND2_X1 U5728 ( .A1(n4523), .A2(n4527), .ZN(n9360) );
  NAND2_X1 U5729 ( .A1(n9376), .A2(n9085), .ZN(n4523) );
  OAI21_X1 U5730 ( .B1(n9376), .B2(n9172), .A(n9085), .ZN(n9361) );
  AOI21_X1 U5731 ( .B1(n4538), .B2(n4541), .A(n4537), .ZN(n4536) );
  INV_X1 U5732 ( .A(n4747), .ZN(n4537) );
  OR2_X1 U5733 ( .A1(n5489), .A2(n5488), .ZN(n9409) );
  AND2_X1 U5734 ( .A1(n9419), .A2(n9409), .ZN(n9410) );
  AND2_X1 U5735 ( .A1(n5462), .A2(n5461), .ZN(n9466) );
  NAND2_X1 U5736 ( .A1(n9520), .A2(n4310), .ZN(n9487) );
  OR2_X1 U5737 ( .A1(n5386), .A2(n5385), .ZN(n5406) );
  NAND2_X1 U5738 ( .A1(n4511), .A2(n4510), .ZN(n9479) );
  AOI21_X1 U5739 ( .B1(n4513), .B2(n4515), .A(n4365), .ZN(n4510) );
  AND2_X1 U5740 ( .A1(n5374), .A2(n4514), .ZN(n4513) );
  AND2_X1 U5741 ( .A1(n9497), .A2(n4754), .ZN(n4753) );
  NAND2_X1 U5742 ( .A1(n9154), .A2(n9153), .ZN(n4754) );
  OR2_X1 U5743 ( .A1(n9514), .A2(n9154), .ZN(n4752) );
  NAND2_X1 U5744 ( .A1(n4512), .A2(n4516), .ZN(n9530) );
  NAND2_X1 U5745 ( .A1(n9534), .A2(n4517), .ZN(n4512) );
  AND2_X1 U5746 ( .A1(n9520), .A2(n9741), .ZN(n9521) );
  INV_X1 U5747 ( .A(n4530), .ZN(n7866) );
  INV_X1 U5748 ( .A(n9104), .ZN(n9552) );
  NAND2_X1 U5749 ( .A1(n7339), .A2(n4351), .ZN(n9570) );
  NAND2_X1 U5750 ( .A1(n4506), .A2(n4502), .ZN(n9567) );
  AND2_X1 U5751 ( .A1(n4857), .A2(n4504), .ZN(n4502) );
  NAND2_X1 U5752 ( .A1(n4858), .A2(n4505), .ZN(n4504) );
  AND2_X1 U5753 ( .A1(n5635), .A2(n9548), .ZN(n9568) );
  NAND2_X1 U5754 ( .A1(n5634), .A2(n4317), .ZN(n9559) );
  AND2_X1 U5755 ( .A1(n7339), .A2(n4320), .ZN(n9572) );
  NAND2_X1 U5756 ( .A1(n7339), .A2(n4303), .ZN(n7657) );
  OR2_X1 U5757 ( .A1(n5209), .A2(n10248), .ZN(n5231) );
  NAND2_X1 U5758 ( .A1(n8559), .A2(n9224), .ZN(n4509) );
  NAND2_X1 U5759 ( .A1(n5190), .A2(n4845), .ZN(n5192) );
  NOR2_X1 U5760 ( .A1(n7343), .A2(n7336), .ZN(n4845) );
  AND2_X1 U5761 ( .A1(n7419), .A2(n9942), .ZN(n7339) );
  INV_X1 U5762 ( .A(n7309), .ZN(n9098) );
  NOR2_X1 U5763 ( .A1(n7420), .A2(n8944), .ZN(n7419) );
  NAND2_X1 U5764 ( .A1(n4763), .A2(n4762), .ZN(n8944) );
  NAND2_X1 U5765 ( .A1(n6565), .A2(n5399), .ZN(n4762) );
  INV_X1 U5766 ( .A(n4862), .ZN(n4763) );
  OAI21_X1 U5767 ( .B1(n4492), .B2(n6570), .A(n5148), .ZN(n4862) );
  INV_X1 U5768 ( .A(n7414), .ZN(n4469) );
  AND2_X1 U5769 ( .A1(n7411), .A2(n7412), .ZN(n4684) );
  NAND2_X1 U5770 ( .A1(n9004), .A2(n9012), .ZN(n9005) );
  AND2_X1 U5771 ( .A1(n7414), .A2(n7412), .ZN(n9095) );
  OR2_X1 U5772 ( .A1(n7438), .A2(n7599), .ZN(n7420) );
  NAND2_X1 U5773 ( .A1(n5120), .A2(n5119), .ZN(n7437) );
  INV_X1 U5774 ( .A(n9902), .ZN(n7426) );
  NAND3_X1 U5775 ( .A1(n9896), .A2(n9889), .A3(n6715), .ZN(n7427) );
  OR2_X1 U5776 ( .A1(n9593), .A2(n9592), .ZN(n9594) );
  NAND2_X1 U5777 ( .A1(n5549), .A2(n5548), .ZN(n9352) );
  AND3_X1 U5778 ( .A1(n4764), .A2(n5139), .A3(n5142), .ZN(n9944) );
  AND2_X1 U5779 ( .A1(n5140), .A2(n5141), .ZN(n4764) );
  INV_X1 U5780 ( .A(n9950), .ZN(n9966) );
  AND2_X1 U5781 ( .A1(n9887), .A2(n9894), .ZN(n9950) );
  XNOR2_X1 U5782 ( .A(n4611), .B(n5730), .ZN(n8544) );
  OAI211_X1 U5783 ( .C1(n5741), .C2(SI_30_), .A(n5724), .B(n5725), .ZN(n4611)
         );
  XNOR2_X1 U5784 ( .A(n5733), .B(n5736), .ZN(n8551) );
  NAND2_X1 U5786 ( .A1(n4613), .A2(n4617), .ZN(n5596) );
  OR2_X1 U5787 ( .A1(n5560), .A2(n4620), .ZN(n4613) );
  XNOR2_X1 U5788 ( .A(n5676), .B(n5675), .ZN(n7816) );
  INV_X1 U5789 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n5675) );
  NAND2_X1 U5790 ( .A1(n5674), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5676) );
  NAND2_X1 U5791 ( .A1(n4621), .A2(n5558), .ZN(n5577) );
  NAND2_X1 U5792 ( .A1(n4624), .A2(n4625), .ZN(n5539) );
  OR2_X1 U5793 ( .A1(n5446), .A2(n5445), .ZN(n5448) );
  AND2_X1 U5794 ( .A1(n5381), .A2(n5400), .ZN(n9255) );
  NAND2_X1 U5795 ( .A1(n4900), .A2(n5354), .ZN(n5375) );
  NAND2_X1 U5796 ( .A1(n4895), .A2(n4901), .ZN(n4900) );
  NAND2_X1 U5797 ( .A1(n4880), .A2(n4882), .ZN(n5331) );
  OAI21_X1 U5798 ( .B1(n5292), .B2(n5291), .A(n5290), .ZN(n5316) );
  OR2_X1 U5799 ( .A1(n5225), .A2(P1_IR_REG_10__SCAN_IN), .ZN(n5275) );
  AND2_X1 U5800 ( .A1(n5201), .A2(n5200), .ZN(n5204) );
  XNOR2_X1 U5801 ( .A(n5216), .B(n5215), .ZN(n6585) );
  AND2_X1 U5802 ( .A1(n5378), .A2(n5177), .ZN(n5201) );
  XNOR2_X1 U5803 ( .A(n5194), .B(n5195), .ZN(n6568) );
  NAND2_X1 U5804 ( .A1(n5060), .A2(n5059), .ZN(n5194) );
  NOR2_X1 U5805 ( .A1(n5022), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n5378) );
  XNOR2_X1 U5806 ( .A(n5160), .B(n5159), .ZN(n5869) );
  INV_X1 U5807 ( .A(n5043), .ZN(n5113) );
  NOR2_X1 U5808 ( .A1(n9782), .A2(n10287), .ZN(n9783) );
  NAND2_X1 U5809 ( .A1(n9787), .A2(n9788), .ZN(n9789) );
  NAND2_X1 U5810 ( .A1(n4447), .A2(n6447), .ZN(n7805) );
  NAND2_X1 U5811 ( .A1(n6093), .A2(n6092), .ZN(n8461) );
  AND4_X1 U5812 ( .A1(n5930), .A2(n5929), .A3(n5928), .A4(n5927), .ZN(n7565)
         );
  NAND2_X1 U5813 ( .A1(n4913), .A2(n6470), .ZN(n7930) );
  NAND2_X1 U5814 ( .A1(n6114), .A2(n6113), .ZN(n8452) );
  AND3_X1 U5815 ( .A1(n6008), .A2(n6007), .A3(n6006), .ZN(n8406) );
  NAND2_X1 U5816 ( .A1(n4594), .A2(n4306), .ZN(n4593) );
  NAND2_X1 U5817 ( .A1(n4306), .A2(n6454), .ZN(n4595) );
  INV_X1 U5818 ( .A(n4596), .ZN(n4594) );
  OR2_X1 U5819 ( .A1(n5858), .A2(n7518), .ZN(n5806) );
  NAND2_X1 U5820 ( .A1(n7927), .A2(n6478), .ZN(n7985) );
  OR2_X1 U5821 ( .A1(n6549), .A2(P2_U3152), .ZN(n8037) );
  XNOR2_X1 U5822 ( .A(n7704), .B(n6494), .ZN(n7402) );
  AND4_X1 U5823 ( .A1(n5943), .A2(n5942), .A3(n5941), .A4(n5940), .ZN(n7881)
         );
  OR2_X1 U5824 ( .A1(n8044), .A2(n6387), .ZN(n8008) );
  INV_X1 U5825 ( .A(n8033), .ZN(n8020) );
  AND2_X1 U5826 ( .A1(n7205), .A2(n6405), .ZN(n6406) );
  CLKBUF_X1 U5827 ( .A(n7052), .Z(n7053) );
  INV_X1 U5828 ( .A(n8008), .ZN(n8049) );
  OAI21_X1 U5829 ( .B1(n6376), .B2(n6377), .A(n6375), .ZN(n6378) );
  AND2_X1 U5830 ( .A1(n6159), .A2(n6158), .ZN(n8202) );
  OR2_X1 U5831 ( .A1(n8193), .A2(n6076), .ZN(n6159) );
  INV_X1 U5832 ( .A(n8182), .ZN(n8226) );
  INV_X1 U5833 ( .A(n8173), .ZN(n8334) );
  OR2_X1 U5834 ( .A1(n8362), .A2(n6076), .ZN(n6047) );
  OR2_X1 U5835 ( .A1(n6718), .A2(n10032), .ZN(n8056) );
  NAND2_X1 U5836 ( .A1(n5802), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n4431) );
  OR2_X1 U5837 ( .A1(n5858), .A2(n5823), .ZN(n5824) );
  NAND2_X1 U5838 ( .A1(n8071), .A2(n8072), .ZN(n8070) );
  NAND2_X1 U5839 ( .A1(n6748), .A2(n6747), .ZN(n6823) );
  NAND2_X1 U5840 ( .A1(n6757), .A2(n6756), .ZN(n6856) );
  NAND2_X1 U5841 ( .A1(n6839), .A2(n6838), .ZN(n8111) );
  XNOR2_X1 U5842 ( .A(n7691), .B(n7692), .ZN(n7694) );
  OAI21_X1 U5843 ( .B1(n8118), .B2(n8117), .A(n8119), .ZN(n10001) );
  AOI21_X1 U5844 ( .B1(n7894), .B2(n6182), .A(n6162), .ZN(n8429) );
  INV_X1 U5845 ( .A(n8437), .ZN(n8213) );
  NAND2_X1 U5846 ( .A1(n4707), .A2(n8206), .ZN(n8436) );
  NAND2_X1 U5847 ( .A1(n8217), .A2(n4708), .ZN(n4707) );
  NAND2_X1 U5848 ( .A1(n8275), .A2(n6331), .ZN(n8255) );
  NAND2_X1 U5849 ( .A1(n8280), .A2(n4977), .ZN(n8264) );
  INV_X1 U5850 ( .A(n8461), .ZN(n8285) );
  NAND2_X1 U5851 ( .A1(n4888), .A2(n6320), .ZN(n8306) );
  OAI21_X1 U5852 ( .B1(n8327), .B2(n4714), .A(n4712), .ZN(n8298) );
  NAND2_X1 U5853 ( .A1(n6071), .A2(n6319), .ZN(n8319) );
  AND2_X1 U5854 ( .A1(n6073), .A2(n6072), .ZN(n8317) );
  NAND2_X1 U5855 ( .A1(n8325), .A2(n4982), .ZN(n4956) );
  AND2_X1 U5856 ( .A1(n6060), .A2(n6059), .ZN(n8330) );
  NAND2_X1 U5857 ( .A1(n4717), .A2(n4718), .ZN(n8339) );
  OR2_X1 U5858 ( .A1(n4454), .A2(n4720), .ZN(n4717) );
  NAND2_X1 U5859 ( .A1(n8383), .A2(n6048), .ZN(n8367) );
  NAND2_X1 U5860 ( .A1(n7795), .A2(n4769), .ZN(n8361) );
  NAND2_X1 U5861 ( .A1(n8380), .A2(n4721), .ZN(n8359) );
  NAND2_X1 U5862 ( .A1(n7769), .A2(n6294), .ZN(n7787) );
  NAND2_X1 U5863 ( .A1(n7767), .A2(n7766), .ZN(n7789) );
  NAND2_X1 U5864 ( .A1(n4959), .A2(n7028), .ZN(n7171) );
  OR2_X1 U5865 ( .A1(n6000), .A2(n6567), .ZN(n5821) );
  AND2_X2 U5866 ( .A1(n7070), .A2(n7069), .ZN(n10100) );
  NAND2_X1 U5867 ( .A1(n4780), .A2(n4348), .ZN(n8525) );
  INV_X1 U5868 ( .A(n8433), .ZN(n4419) );
  INV_X1 U5869 ( .A(n8434), .ZN(n4420) );
  AND2_X2 U5870 ( .A1(n7070), .A2(n7017), .ZN(n10283) );
  AND3_X1 U5871 ( .A1(n7374), .A2(n10029), .A3(n7016), .ZN(n7017) );
  NAND2_X1 U5872 ( .A1(n10030), .A2(n10029), .ZN(n10035) );
  NAND2_X1 U5873 ( .A1(n6546), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10032) );
  NOR2_X1 U5874 ( .A1(n5796), .A2(P2_IR_REG_29__SCAN_IN), .ZN(n4973) );
  INV_X1 U5875 ( .A(n5804), .ZN(n8553) );
  AND2_X1 U5876 ( .A1(n5813), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5818) );
  CLKBUF_X1 U5877 ( .A(n6368), .Z(n6369) );
  INV_X1 U5878 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7721) );
  XNOR2_X1 U5879 ( .A(n6357), .B(n6356), .ZN(n7722) );
  INV_X1 U5880 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n6356) );
  NAND2_X1 U5881 ( .A1(n6355), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6357) );
  INV_X1 U5882 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n10187) );
  INV_X1 U5883 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7369) );
  NAND2_X1 U5884 ( .A1(n6050), .A2(n4918), .ZN(n6170) );
  INV_X1 U5885 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7290) );
  INV_X1 U5886 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n6191) );
  INV_X1 U5887 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7212) );
  INV_X1 U5888 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n10216) );
  INV_X1 U5889 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n10235) );
  INV_X1 U5890 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6678) );
  INV_X1 U5891 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6602) );
  INV_X1 U5892 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n10144) );
  AND2_X1 U5893 ( .A1(n5604), .A2(n5590), .ZN(n9320) );
  NAND2_X1 U5894 ( .A1(n4808), .A2(n4812), .ZN(n8970) );
  NAND2_X1 U5895 ( .A1(n4490), .A2(n4813), .ZN(n4808) );
  AND4_X1 U5896 ( .A1(n5258), .A2(n5257), .A3(n5256), .A4(n5255), .ZN(n9575)
         );
  NAND2_X1 U5897 ( .A1(n4816), .A2(n8891), .ZN(n8815) );
  AND4_X1 U5898 ( .A1(n5314), .A2(n5313), .A3(n5312), .A4(n5311), .ZN(n8830)
         );
  AND4_X1 U5899 ( .A1(n5391), .A2(n5390), .A3(n5389), .A4(n5388), .ZN(n9503)
         );
  NAND2_X1 U5900 ( .A1(n4804), .A2(n4809), .ZN(n8843) );
  OR2_X1 U5901 ( .A1(n4490), .A2(n4811), .ZN(n4804) );
  AND3_X1 U5902 ( .A1(n5410), .A2(n5409), .A3(n5408), .ZN(n9485) );
  INV_X1 U5903 ( .A(n9912), .ZN(n7442) );
  AND4_X1 U5904 ( .A1(n5329), .A2(n5328), .A3(n5327), .A4(n5326), .ZN(n9519)
         );
  NAND2_X1 U5905 ( .A1(n8922), .A2(n8592), .ZN(n8923) );
  AND2_X1 U5906 ( .A1(n7006), .A2(n6710), .ZN(n8959) );
  INV_X1 U5907 ( .A(n8959), .ZN(n8986) );
  AND4_X1 U5908 ( .A1(n5373), .A2(n5372), .A3(n5371), .A4(n5370), .ZN(n9517)
         );
  OR2_X1 U5909 ( .A1(n6712), .A2(n6711), .ZN(n8980) );
  AND2_X1 U5910 ( .A1(n7163), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8984) );
  AOI21_X1 U5911 ( .B1(n4686), .B2(n4685), .A(n4470), .ZN(n9210) );
  NOR2_X1 U5912 ( .A1(n9079), .A2(n9082), .ZN(n4685) );
  NAND2_X1 U5913 ( .A1(n4688), .A2(n4355), .ZN(n4470) );
  NAND2_X1 U5914 ( .A1(n4687), .A2(n9080), .ZN(n4686) );
  OR2_X1 U5915 ( .A1(n6709), .A2(n5697), .ZN(n8991) );
  INV_X1 U5916 ( .A(n9350), .ZN(n9377) );
  INV_X1 U5917 ( .A(n9575), .ZN(n9689) );
  INV_X1 U5918 ( .A(n7607), .ZN(n9227) );
  INV_X1 U5919 ( .A(n5105), .ZN(n9229) );
  NAND2_X1 U5920 ( .A1(n5652), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n5087) );
  OR2_X1 U5921 ( .A1(n6603), .A2(P1_U3084), .ZN(n9230) );
  AND3_X1 U5922 ( .A1(n5078), .A2(n5079), .A3(n5080), .ZN(n4425) );
  OAI21_X1 U5923 ( .B1(n6642), .B2(n6615), .A(n4484), .ZN(n6645) );
  NAND2_X1 U5924 ( .A1(n6645), .A2(n6644), .ZN(n6643) );
  NAND2_X1 U5925 ( .A1(n4743), .A2(n5075), .ZN(n5161) );
  INV_X1 U5926 ( .A(n4560), .ZN(n6670) );
  OAI21_X1 U5927 ( .B1(n6669), .B2(P1_REG1_REG_7__SCAN_IN), .A(n6668), .ZN(
        n6867) );
  NAND2_X1 U5928 ( .A1(n6671), .A2(n7315), .ZN(n4559) );
  INV_X1 U5929 ( .A(n4558), .ZN(n6885) );
  INV_X1 U5930 ( .A(n4782), .ZN(n6923) );
  AND2_X1 U5931 ( .A1(n5305), .A2(n5304), .ZN(n9820) );
  INV_X1 U5932 ( .A(n9252), .ZN(n4567) );
  NAND2_X1 U5933 ( .A1(n9185), .A2(n9189), .ZN(n9598) );
  NAND2_X1 U5934 ( .A1(n9331), .A2(n9127), .ZN(n9324) );
  AOI22_X1 U5935 ( .A1(n9334), .A2(n9563), .B1(n9562), .B2(n9333), .ZN(n9608)
         );
  AND4_X1 U5936 ( .A1(n5555), .A2(n5554), .A3(n5553), .A4(n5552), .ZN(n9609)
         );
  OAI21_X1 U5937 ( .B1(n9376), .B2(n4526), .A(n4524), .ZN(n9347) );
  NAND2_X1 U5938 ( .A1(n4852), .A2(n4853), .ZN(n9359) );
  NAND2_X1 U5939 ( .A1(n9397), .A2(n4325), .ZN(n4852) );
  NAND2_X1 U5940 ( .A1(n9397), .A2(n5507), .ZN(n9380) );
  AND2_X1 U5941 ( .A1(n5484), .A2(n5483), .ZN(n9633) );
  NAND2_X1 U5942 ( .A1(n5501), .A2(n5500), .ZN(n9405) );
  NAND2_X1 U5943 ( .A1(n4750), .A2(n9089), .ZN(n9420) );
  NAND2_X1 U5944 ( .A1(n9452), .A2(n9058), .ZN(n4750) );
  NAND2_X1 U5945 ( .A1(n5472), .A2(n5471), .ZN(n9641) );
  AND3_X1 U5946 ( .A1(n9441), .A2(n9440), .A3(n9569), .ZN(n9646) );
  NAND2_X1 U5947 ( .A1(n5435), .A2(n5434), .ZN(n9435) );
  OR2_X1 U5948 ( .A1(n9471), .A2(n9470), .ZN(n9659) );
  NAND2_X1 U5949 ( .A1(n5404), .A2(n5403), .ZN(n9657) );
  OAI21_X1 U5950 ( .B1(n9534), .B2(n4329), .A(n5315), .ZN(n7864) );
  NAND2_X1 U5951 ( .A1(n5278), .A2(n5277), .ZN(n9690) );
  NAND2_X1 U5952 ( .A1(n5634), .A2(n9139), .ZN(n7664) );
  NAND2_X1 U5953 ( .A1(n7497), .A2(n5237), .ZN(n7656) );
  AND2_X1 U5954 ( .A1(n7308), .A2(n9017), .ZN(n4984) );
  INV_X1 U5955 ( .A(n9944), .ZN(n9226) );
  INV_X1 U5956 ( .A(n7637), .ZN(n9942) );
  INV_X1 U5957 ( .A(n8944), .ZN(n7621) );
  NAND2_X1 U5958 ( .A1(n9541), .A2(n5772), .ZN(n9526) );
  INV_X1 U5959 ( .A(n9580), .ZN(n9528) );
  NAND2_X1 U5960 ( .A1(n7277), .A2(n5627), .ZN(n4758) );
  INV_X1 U5961 ( .A(n9526), .ZN(n9578) );
  INV_X1 U5962 ( .A(n9538), .ZN(n9874) );
  INV_X1 U5963 ( .A(n9352), .ZN(n9714) );
  AND2_X1 U5964 ( .A1(n5518), .A2(n5517), .ZN(n9722) );
  INV_X1 U5965 ( .A(n9435), .ZN(n9731) );
  AND2_X2 U5966 ( .A1(n5767), .A2(n5706), .ZN(n9970) );
  INV_X1 U5967 ( .A(n9880), .ZN(n9881) );
  AND2_X1 U5968 ( .A1(n7158), .A2(n5695), .ZN(n9884) );
  MUX2_X1 U5969 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5002), .S(
        P1_IR_REG_29__SCAN_IN), .Z(n5004) );
  CLKBUF_X1 U5970 ( .A(n7816), .Z(n4464) );
  INV_X1 U5971 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7783) );
  NAND2_X1 U5972 ( .A1(n5674), .A2(n5670), .ZN(n7784) );
  INV_X1 U5973 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n10232) );
  XNOR2_X1 U5974 ( .A(n5672), .B(n5671), .ZN(n7724) );
  INV_X1 U5975 ( .A(n4996), .ZN(n4933) );
  INV_X1 U5976 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7350) );
  INV_X1 U5977 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7288) );
  INV_X1 U5978 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7269) );
  INV_X1 U5979 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7210) );
  INV_X1 U5980 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n7109) );
  INV_X1 U5981 ( .A(n9255), .ZN(n9858) );
  INV_X1 U5982 ( .A(n9832), .ZN(n9264) );
  INV_X1 U5983 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n6697) );
  INV_X1 U5984 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n6679) );
  INV_X1 U5985 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n6590) );
  INV_X1 U5986 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6592) );
  INV_X1 U5987 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n6594) );
  INV_X1 U5988 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n6586) );
  INV_X1 U5989 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n6581) );
  NAND2_X1 U5990 ( .A1(n4562), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4561) );
  NAND2_X1 U5991 ( .A1(n5129), .A2(n5114), .ZN(n4562) );
  CLKBUF_X1 U5992 ( .A(n9238), .Z(n4477) );
  INV_X1 U5993 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10105) );
  OAI21_X1 U5994 ( .B1(n10101), .B2(n10105), .A(n10103), .ZN(n10299) );
  INV_X1 U5995 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n9774) );
  AND2_X1 U5996 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n9781), .ZN(n10288) );
  XNOR2_X1 U5997 ( .A(n9783), .B(n4442), .ZN(n10286) );
  XNOR2_X1 U5998 ( .A(n9786), .B(n4440), .ZN(n10290) );
  INV_X1 U5999 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n4440) );
  XNOR2_X1 U6000 ( .A(n9789), .B(n4441), .ZN(n10295) );
  INV_X1 U6001 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n4441) );
  NOR2_X1 U6002 ( .A1(n9793), .A2(n10296), .ZN(n10129) );
  NOR2_X1 U6003 ( .A1(n10124), .A2(n4403), .ZN(n10123) );
  NAND2_X1 U6004 ( .A1(n10123), .A2(n10122), .ZN(n10121) );
  OAI21_X1 U6005 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10121), .ZN(n10119) );
  NAND2_X1 U6006 ( .A1(n10119), .A2(n10120), .ZN(n10118) );
  NAND2_X1 U6007 ( .A1(n10118), .A2(n4436), .ZN(n10116) );
  NAND2_X1 U6008 ( .A1(n4438), .A2(n4437), .ZN(n4436) );
  INV_X1 U6009 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n4438) );
  OAI21_X1 U6010 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10115), .ZN(n10113) );
  OAI21_X1 U6011 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n10112), .ZN(n10110) );
  NAND2_X1 U6012 ( .A1(n10110), .A2(n10111), .ZN(n10109) );
  NAND2_X1 U6013 ( .A1(n10109), .A2(n4439), .ZN(n10107) );
  NAND2_X1 U6014 ( .A1(n9850), .A2(n10156), .ZN(n4439) );
  AND2_X1 U6015 ( .A1(n7905), .A2(n4397), .ZN(n4426) );
  NAND2_X1 U6016 ( .A1(n4608), .A2(n4606), .ZN(n8031) );
  NAND2_X1 U6017 ( .A1(n8151), .A2(n8392), .ZN(n4487) );
  NAND2_X1 U6018 ( .A1(n4353), .A2(n4407), .ZN(P2_U3269) );
  INV_X1 U6019 ( .A(n4408), .ZN(n4407) );
  AOI21_X1 U6020 ( .B1(n4423), .B2(n9418), .A(n4422), .ZN(n4421) );
  OR2_X1 U6021 ( .A1(n9287), .A2(n9418), .ZN(n4424) );
  NAND2_X1 U6022 ( .A1(n5779), .A2(n5778), .ZN(n5780) );
  MUX2_X1 U6023 ( .A(n5754), .B(n5757), .S(n9986), .Z(n5756) );
  MUX2_X1 U6024 ( .A(n9586), .B(n9702), .S(n9986), .Z(n9587) );
  AND2_X1 U6025 ( .A1(n5701), .A2(n5700), .ZN(n5702) );
  MUX2_X1 U6026 ( .A(n5758), .B(n5757), .S(n9970), .Z(n5761) );
  MUX2_X1 U6027 ( .A(n9703), .B(n9702), .S(n9970), .Z(n9704) );
  NAND2_X1 U6028 ( .A1(n4533), .A2(n4531), .ZN(P1_U3520) );
  OR2_X1 U6029 ( .A1(n9970), .A2(n4532), .ZN(n4531) );
  INV_X1 U6030 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n4532) );
  AOI21_X1 U6031 ( .B1(n9298), .B2(n5759), .A(n5709), .ZN(n5710) );
  OAI21_X1 U6032 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n9797), .A(n10291), .ZN(
        n9799) );
  AND2_X1 U6033 ( .A1(n5659), .A2(n4952), .ZN(n4303) );
  INV_X1 U6034 ( .A(n8490), .ZN(n4722) );
  INV_X1 U6035 ( .A(n5841), .ZN(n10050) );
  NAND3_X2 U6036 ( .A1(n5840), .A2(n5839), .A3(n5838), .ZN(n5841) );
  OR2_X1 U6037 ( .A1(n8452), .A2(n8273), .ZN(n6334) );
  OR2_X1 U6038 ( .A1(n5490), .A2(n9410), .ZN(n4304) );
  AND2_X1 U6039 ( .A1(n8207), .A2(n4962), .ZN(n4305) );
  AND2_X1 U6040 ( .A1(n6460), .A2(n7960), .ZN(n4306) );
  OR2_X1 U6041 ( .A1(n9388), .A2(n9393), .ZN(n4307) );
  AND2_X1 U6042 ( .A1(n7838), .A2(n6347), .ZN(n4308) );
  AND2_X1 U6043 ( .A1(n4361), .A2(n4721), .ZN(n4309) );
  AND2_X1 U6044 ( .A1(n4950), .A2(n4949), .ZN(n4310) );
  INV_X1 U6045 ( .A(n8181), .ZN(n4963) );
  OR2_X1 U6046 ( .A1(n9678), .A2(n9553), .ZN(n4311) );
  AND2_X1 U6047 ( .A1(n4718), .A2(n4354), .ZN(n4312) );
  NAND2_X1 U6048 ( .A1(n8566), .A2(n9223), .ZN(n4313) );
  AND2_X1 U6049 ( .A1(n4897), .A2(n5394), .ZN(n4314) );
  NAND2_X1 U6050 ( .A1(n5365), .A2(n5364), .ZN(n9506) );
  AND3_X1 U6051 ( .A1(n9103), .A2(n9102), .A3(n4374), .ZN(n4315) );
  AND2_X1 U6052 ( .A1(n4625), .A2(n5538), .ZN(n4316) );
  AND2_X1 U6053 ( .A1(n9139), .A2(n9138), .ZN(n4317) );
  NAND2_X1 U6054 ( .A1(n6184), .A2(n6183), .ZN(n8423) );
  INV_X1 U6055 ( .A(n8423), .ZN(n4656) );
  INV_X1 U6056 ( .A(n7735), .ZN(n8059) );
  AND4_X1 U6057 ( .A1(n5966), .A2(n5965), .A3(n5964), .A4(n5963), .ZN(n7735)
         );
  AND2_X1 U6058 ( .A1(n4734), .A2(n4908), .ZN(n4318) );
  OR2_X1 U6059 ( .A1(n9641), .A2(n9633), .ZN(n9061) );
  INV_X1 U6060 ( .A(n9061), .ZN(n4748) );
  NAND4_X1 U6061 ( .A1(n4933), .A2(n4995), .A3(n5377), .A4(n4932), .ZN(n4319)
         );
  AND2_X1 U6062 ( .A1(n4303), .A2(n4951), .ZN(n4320) );
  AND2_X1 U6063 ( .A1(n4708), .A2(n10086), .ZN(n4321) );
  AND2_X1 U6064 ( .A1(n4580), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n4322) );
  INV_X1 U6065 ( .A(n8270), .ZN(n4838) );
  NAND2_X1 U6066 ( .A1(n5229), .A2(n5228), .ZN(n8580) );
  INV_X1 U6067 ( .A(n8580), .ZN(n4952) );
  NAND2_X1 U6068 ( .A1(n5135), .A2(n5134), .ZN(n7303) );
  AOI21_X1 U6069 ( .B1(n8233), .B2(n6138), .A(n6130), .ZN(n8179) );
  OR2_X2 U6070 ( .A1(n9570), .A2(n9681), .ZN(n4323) );
  NAND2_X1 U6071 ( .A1(n7803), .A2(n6454), .ZN(n7955) );
  INV_X1 U6072 ( .A(n5150), .ZN(n5481) );
  INV_X1 U6073 ( .A(n6039), .ZN(n4904) );
  NAND2_X1 U6074 ( .A1(n6193), .A2(n8392), .ZN(n6466) );
  XNOR2_X1 U6075 ( .A(n8441), .B(n8239), .ZN(n8225) );
  INV_X1 U6076 ( .A(n8225), .ZN(n4909) );
  NAND2_X1 U6077 ( .A1(n9520), .A2(n4950), .ZN(n9486) );
  AND2_X1 U6078 ( .A1(n9367), .A2(n4946), .ZN(n4324) );
  AND2_X1 U6079 ( .A1(n4307), .A2(n5507), .ZN(n4325) );
  AND2_X1 U6080 ( .A1(n9319), .A2(n4941), .ZN(n4326) );
  NAND2_X1 U6081 ( .A1(n8209), .A2(n4779), .ZN(n4327) );
  OR2_X1 U6082 ( .A1(n6266), .A2(n6349), .ZN(n4328) );
  AND2_X1 U6083 ( .A1(n9681), .A2(n9561), .ZN(n4329) );
  AND2_X1 U6084 ( .A1(n4831), .A2(n6282), .ZN(n4330) );
  INV_X2 U6085 ( .A(n7073), .ZN(n8779) );
  NAND2_X1 U6086 ( .A1(n5532), .A2(n5531), .ZN(n9369) );
  NAND2_X1 U6087 ( .A1(n4906), .A2(n6039), .ZN(n8486) );
  INV_X1 U6088 ( .A(n8486), .ZN(n4768) );
  AND4_X1 U6089 ( .A1(n9097), .A2(n9096), .A3(n9095), .A4(n9094), .ZN(n4331)
         );
  OAI21_X1 U6090 ( .B1(n4913), .B2(n4604), .A(n4602), .ZN(n7936) );
  INV_X1 U6091 ( .A(n4851), .ZN(n4850) );
  NAND2_X1 U6092 ( .A1(n4853), .A2(n4347), .ZN(n4851) );
  AND2_X1 U6093 ( .A1(n7736), .A2(n7739), .ZN(n4332) );
  INV_X1 U6094 ( .A(n9089), .ZN(n4749) );
  INV_X1 U6095 ( .A(n6494), .ZN(n6400) );
  INV_X1 U6096 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5617) );
  AND2_X1 U6097 ( .A1(n6294), .A2(n6295), .ZN(n7790) );
  INV_X1 U6098 ( .A(n7790), .ZN(n7768) );
  XNOR2_X1 U6099 ( .A(n8456), .B(n8291), .ZN(n8270) );
  INV_X1 U6100 ( .A(n9050), .ZN(n4525) );
  NAND2_X1 U6101 ( .A1(n4913), .A2(n4912), .ZN(n7927) );
  AND2_X1 U6102 ( .A1(n4509), .A2(n4313), .ZN(n4334) );
  AND2_X1 U6103 ( .A1(n9055), .A2(n9436), .ZN(n9454) );
  INV_X1 U6104 ( .A(n9454), .ZN(n4541) );
  AND2_X1 U6105 ( .A1(n9962), .A2(n8806), .ZN(n4335) );
  AND4_X1 U6106 ( .A1(n5013), .A2(n5012), .A3(n5011), .A4(n5010), .ZN(n8884)
         );
  AND2_X1 U6107 ( .A1(n7740), .A2(n4644), .ZN(n4336) );
  INV_X1 U6108 ( .A(n9523), .ZN(n9741) );
  NAND2_X1 U6109 ( .A1(n5345), .A2(n5344), .ZN(n9523) );
  AND2_X1 U6110 ( .A1(n7221), .A2(n4328), .ZN(n4337) );
  INV_X1 U6111 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n9752) );
  AND2_X1 U6112 ( .A1(n4752), .A2(n9153), .ZN(n4338) );
  AND2_X1 U6113 ( .A1(n5745), .A2(n5744), .ZN(n9705) );
  INV_X1 U6114 ( .A(n9705), .ZN(n8999) );
  AND2_X1 U6115 ( .A1(n7336), .A2(n9017), .ZN(n4339) );
  AND2_X1 U6116 ( .A1(n6036), .A2(n6035), .ZN(n8408) );
  NAND2_X1 U6117 ( .A1(n6084), .A2(n6083), .ZN(n8466) );
  INV_X1 U6118 ( .A(n4699), .ZN(n4698) );
  AND2_X1 U6119 ( .A1(n8184), .A2(n6342), .ZN(n4340) );
  INV_X1 U6120 ( .A(n9464), .ZN(n9470) );
  OR2_X1 U6121 ( .A1(n8218), .A2(n8225), .ZN(n4341) );
  AND2_X1 U6122 ( .A1(n9470), .A2(n9046), .ZN(n4342) );
  AND2_X1 U6123 ( .A1(n9506), .A2(n9220), .ZN(n4343) );
  AND2_X1 U6124 ( .A1(n7768), .A2(n7766), .ZN(n4344) );
  AND2_X1 U6125 ( .A1(n9061), .A2(n9060), .ZN(n5642) );
  INV_X1 U6126 ( .A(n5642), .ZN(n9419) );
  NAND2_X1 U6127 ( .A1(n7620), .A2(n7630), .ZN(n4345) );
  NAND2_X1 U6128 ( .A1(n9408), .A2(n5485), .ZN(n4346) );
  NAND2_X1 U6129 ( .A1(n9369), .A2(n9377), .ZN(n4347) );
  AND2_X1 U6130 ( .A1(n8424), .A2(n8427), .ZN(n4348) );
  NAND2_X1 U6131 ( .A1(n9379), .A2(n5527), .ZN(n4349) );
  AND2_X1 U6132 ( .A1(n4865), .A2(n4867), .ZN(n4350) );
  AND2_X1 U6133 ( .A1(n4320), .A2(n9571), .ZN(n4351) );
  NAND2_X1 U6134 ( .A1(n7961), .A2(n6455), .ZN(n4352) );
  OR2_X1 U6135 ( .A1(n8444), .A2(n4281), .ZN(n4353) );
  NAND2_X1 U6136 ( .A1(n8482), .A2(n8373), .ZN(n4354) );
  NAND2_X1 U6137 ( .A1(n9083), .A2(n9082), .ZN(n4355) );
  NAND2_X1 U6138 ( .A1(n8168), .A2(n8164), .ZN(n4968) );
  INV_X1 U6139 ( .A(n8154), .ZN(n8431) );
  NAND2_X1 U6140 ( .A1(n6154), .A2(n6153), .ZN(n8154) );
  INV_X1 U6141 ( .A(n6454), .ZN(n4598) );
  OR2_X1 U6142 ( .A1(n9352), .A2(n9609), .ZN(n9176) );
  INV_X1 U6143 ( .A(n9176), .ZN(n4522) );
  NOR2_X1 U6144 ( .A1(n9369), .A2(n9377), .ZN(n4356) );
  NOR2_X1 U6145 ( .A1(n8920), .A2(n9689), .ZN(n4357) );
  INV_X1 U6146 ( .A(n4787), .ZN(n8282) );
  NOR2_X1 U6147 ( .A1(n8314), .A2(n4789), .ZN(n4787) );
  INV_X1 U6148 ( .A(n4518), .ZN(n4517) );
  NAND2_X1 U6149 ( .A1(n4311), .A2(n5315), .ZN(n4518) );
  INV_X1 U6150 ( .A(n4896), .ZN(n4894) );
  NAND2_X1 U6151 ( .A1(n4975), .A2(n4901), .ZN(n4896) );
  NAND2_X1 U6152 ( .A1(n5738), .A2(n5737), .ZN(n9303) );
  INV_X1 U6153 ( .A(n9303), .ZN(n4943) );
  INV_X1 U6154 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n5027) );
  OR2_X1 U6155 ( .A1(n8466), .A2(n8009), .ZN(n6091) );
  INV_X1 U6156 ( .A(n8167), .ZN(n4969) );
  AND2_X1 U6157 ( .A1(n8494), .A2(n8166), .ZN(n8167) );
  AND2_X1 U6158 ( .A1(n9588), .A2(n9966), .ZN(n4358) );
  AND2_X1 U6159 ( .A1(n8699), .A2(n8700), .ZN(n4359) );
  AND2_X1 U6160 ( .A1(n8213), .A2(n8182), .ZN(n4360) );
  OR2_X1 U6161 ( .A1(n8486), .A2(n8343), .ZN(n4361) );
  AND2_X1 U6162 ( .A1(n8347), .A2(n8170), .ZN(n4362) );
  INV_X1 U6163 ( .A(n4771), .ZN(n4770) );
  NAND2_X1 U6164 ( .A1(n4772), .A2(n7800), .ZN(n4771) );
  AND2_X1 U6165 ( .A1(n4791), .A2(n4795), .ZN(n4363) );
  NAND2_X1 U6166 ( .A1(n5566), .A2(n5565), .ZN(n9342) );
  INV_X1 U6167 ( .A(n9342), .ZN(n4945) );
  NAND2_X1 U6168 ( .A1(n9436), .A2(n9160), .ZN(n4364) );
  NAND2_X1 U6169 ( .A1(n8184), .A2(n6225), .ZN(n8207) );
  OR2_X1 U6170 ( .A1(n4986), .A2(n4343), .ZN(n4365) );
  INV_X1 U6171 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5799) );
  NAND2_X1 U6172 ( .A1(n4493), .A2(n5189), .ZN(n7342) );
  AND2_X1 U6173 ( .A1(n9155), .A2(n9481), .ZN(n9497) );
  NAND2_X1 U6174 ( .A1(n6338), .A2(n6337), .ZN(n8237) );
  INV_X1 U6175 ( .A(n8237), .ZN(n4908) );
  NOR2_X1 U6176 ( .A1(n4768), .A2(n8169), .ZN(n4366) );
  NAND2_X1 U6177 ( .A1(n7411), .A2(n7352), .ZN(n4367) );
  INV_X1 U6178 ( .A(n4895), .ZN(n5356) );
  AND2_X1 U6179 ( .A1(n5335), .A2(n5334), .ZN(n4895) );
  NAND2_X1 U6180 ( .A1(n4519), .A2(n9105), .ZN(n4368) );
  NAND2_X1 U6181 ( .A1(n6333), .A2(n4736), .ZN(n4369) );
  OR2_X1 U6182 ( .A1(n9678), .A2(n9519), .ZN(n9036) );
  AND2_X1 U6183 ( .A1(n6320), .A2(n6321), .ZN(n4370) );
  OR2_X1 U6184 ( .A1(n7945), .A2(n4930), .ZN(n4371) );
  AND2_X1 U6185 ( .A1(n8066), .A2(n4284), .ZN(n4372) );
  AND2_X1 U6186 ( .A1(n8795), .A2(n8796), .ZN(n4373) );
  AND3_X1 U6187 ( .A1(n7336), .A2(n4459), .A3(n9568), .ZN(n4374) );
  AND2_X1 U6188 ( .A1(n4882), .A2(n5330), .ZN(n4375) );
  AND2_X1 U6189 ( .A1(n4769), .A2(n4768), .ZN(n4376) );
  AND2_X1 U6190 ( .A1(n4846), .A2(n9346), .ZN(n4377) );
  NOR2_X1 U6191 ( .A1(n8717), .A2(n8716), .ZN(n4378) );
  AND2_X1 U6192 ( .A1(n6324), .A2(n6319), .ZN(n4379) );
  AND2_X1 U6193 ( .A1(n6205), .A2(n6241), .ZN(n4380) );
  NOR2_X1 U6194 ( .A1(n6297), .A2(n7793), .ZN(n4381) );
  AND2_X1 U6195 ( .A1(n9069), .A2(n9068), .ZN(n4382) );
  AND2_X1 U6196 ( .A1(n9069), .A2(n9127), .ZN(n4383) );
  AND2_X1 U6197 ( .A1(n9293), .A2(n4941), .ZN(n4384) );
  AND2_X1 U6198 ( .A1(n6292), .A2(n7790), .ZN(n4385) );
  OR2_X1 U6199 ( .A1(n6688), .A2(n6652), .ZN(n4386) );
  AND2_X1 U6200 ( .A1(n5619), .A2(n5610), .ZN(n4387) );
  AND2_X1 U6201 ( .A1(n6343), .A2(n4340), .ZN(n4388) );
  AND2_X1 U6202 ( .A1(n6326), .A2(n4840), .ZN(n4389) );
  AND2_X1 U6203 ( .A1(n6332), .A2(n6333), .ZN(n4390) );
  AND2_X1 U6204 ( .A1(n4572), .A2(n4567), .ZN(n4391) );
  AND2_X1 U6205 ( .A1(n4358), .A2(n4861), .ZN(n4392) );
  INV_X1 U6206 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n10142) );
  INV_X1 U6207 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n4739) );
  INV_X1 U6208 ( .A(n9167), .ZN(n4696) );
  NAND2_X1 U6209 ( .A1(n7380), .A2(n10022), .ZN(n8417) );
  NAND2_X1 U6210 ( .A1(n5601), .A2(n5600), .ZN(n9298) );
  INV_X1 U6211 ( .A(n7681), .ZN(n9263) );
  NAND2_X1 U6212 ( .A1(n7795), .A2(n4770), .ZN(n4393) );
  AND2_X1 U6213 ( .A1(n7339), .A2(n5659), .ZN(n4394) );
  OAI21_X1 U6214 ( .B1(n7540), .B2(n7539), .A(n4728), .ZN(n7741) );
  INV_X1 U6215 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n4610) );
  NAND2_X1 U6216 ( .A1(n4876), .A2(n6272), .ZN(n7392) );
  INV_X1 U6217 ( .A(n7843), .ZN(n4644) );
  OAI21_X1 U6218 ( .B1(n4447), .B2(n4595), .A(n4593), .ZN(n7822) );
  OR2_X1 U6219 ( .A1(n9322), .A2(n8981), .ZN(n4395) );
  NAND2_X1 U6220 ( .A1(n7893), .A2(n6427), .ZN(n7560) );
  INV_X1 U6221 ( .A(n7816), .ZN(n4430) );
  INV_X1 U6222 ( .A(n9115), .ZN(n9293) );
  NAND2_X1 U6223 ( .A1(n5732), .A2(n5731), .ZN(n9115) );
  INV_X1 U6224 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n4581) );
  NAND3_X1 U6225 ( .A1(n4995), .A2(n5377), .A3(n4932), .ZN(n4396) );
  INV_X1 U6226 ( .A(n4935), .ZN(n4932) );
  OR2_X1 U6227 ( .A1(n8224), .A2(n8032), .ZN(n4397) );
  NAND2_X2 U6228 ( .A1(n6223), .A2(n6224), .ZN(n6349) );
  INV_X1 U6229 ( .A(n9077), .ZN(n4671) );
  NAND2_X1 U6230 ( .A1(n5251), .A2(n5250), .ZN(n8920) );
  INV_X1 U6231 ( .A(n8920), .ZN(n4951) );
  INV_X1 U6232 ( .A(n9281), .ZN(n9862) );
  INV_X1 U6233 ( .A(n10086), .ZN(n8523) );
  INV_X1 U6234 ( .A(n9859), .ZN(n4479) );
  NAND2_X1 U6235 ( .A1(n5958), .A2(n5957), .ZN(n8519) );
  INV_X1 U6236 ( .A(n8519), .ZN(n4795) );
  NAND2_X1 U6237 ( .A1(n5384), .A2(n5383), .ZN(n9664) );
  INV_X1 U6238 ( .A(n9664), .ZN(n4949) );
  AND2_X1 U6239 ( .A1(n6665), .A2(n6372), .ZN(n8370) );
  INV_X1 U6240 ( .A(n8370), .ZN(n8405) );
  NAND2_X1 U6241 ( .A1(n4864), .A2(n6240), .ZN(n7578) );
  INV_X1 U6242 ( .A(n7645), .ZN(n4799) );
  INV_X1 U6243 ( .A(n8494), .ZN(n4772) );
  INV_X1 U6244 ( .A(n7885), .ZN(n4794) );
  INV_X1 U6245 ( .A(n4296), .ZN(n10019) );
  INV_X1 U6246 ( .A(n9114), .ZN(n4612) );
  INV_X1 U6247 ( .A(n8066), .ZN(n4827) );
  INV_X1 U6248 ( .A(n6695), .ZN(n4655) );
  OR2_X1 U6249 ( .A1(n9311), .A2(n9310), .ZN(n4398) );
  INV_X1 U6250 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n4584) );
  AND2_X1 U6251 ( .A1(n9255), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n4399) );
  AND2_X1 U6252 ( .A1(n4767), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n4400) );
  OR2_X1 U6253 ( .A1(n9267), .A2(n10240), .ZN(n4401) );
  AND2_X1 U6254 ( .A1(P2_REG3_REG_23__SCAN_IN), .A2(P2_REG3_REG_22__SCAN_IN), 
        .ZN(n4402) );
  AND2_X1 U6255 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n4403) );
  AND2_X1 U6256 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n4404) );
  INV_X1 U6257 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n4437) );
  INV_X1 U6258 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n4475) );
  INV_X1 U6259 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n4442) );
  INV_X1 U6260 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n4766) );
  NOR2_X1 U6261 ( .A1(n6313), .A2(n6349), .ZN(n4841) );
  NAND2_X1 U6262 ( .A1(n8366), .A2(n6349), .ZN(n4819) );
  NOR2_X1 U6263 ( .A1(n6300), .A2(n6349), .ZN(n4821) );
  OR2_X1 U6264 ( .A1(n6265), .A2(n6349), .ZN(n4416) );
  MUX2_X1 U6265 ( .A(n6257), .B(n6256), .S(n6349), .Z(n6259) );
  MUX2_X1 U6266 ( .A(n4380), .B(n6236), .S(n6349), .Z(n6258) );
  NAND2_X1 U6267 ( .A1(n7002), .A2(n7001), .ZN(n7083) );
  NAND2_X1 U6268 ( .A1(n5611), .A2(n5610), .ZN(n5612) );
  INV_X1 U6269 ( .A(n6991), .ZN(n4433) );
  INV_X1 U6270 ( .A(n4480), .ZN(n5662) );
  NAND2_X2 U6271 ( .A1(n9198), .A2(n9120), .ZN(n6988) );
  INV_X1 U6272 ( .A(n9284), .ZN(n4406) );
  NAND2_X1 U6273 ( .A1(n4424), .A2(n4421), .ZN(P1_U3260) );
  NAND2_X1 U6274 ( .A1(n9845), .A2(n4401), .ZN(n9863) );
  AOI22_X1 U6275 ( .A1(n6921), .A2(n6920), .B1(n7764), .B2(n6922), .ZN(n7239)
         );
  NAND2_X1 U6276 ( .A1(n9232), .A2(n6608), .ZN(n6609) );
  NAND2_X1 U6277 ( .A1(n6899), .A2(n6900), .ZN(n6904) );
  NOR2_X1 U6278 ( .A1(n6631), .A2(n6632), .ZN(n6656) );
  NAND2_X1 U6279 ( .A1(n6250), .A2(n10013), .ZN(n4864) );
  NOR2_X1 U6280 ( .A1(n8286), .A2(n6101), .ZN(n8269) );
  NAND2_X1 U6281 ( .A1(n8341), .A2(n8342), .ZN(n8340) );
  OAI21_X1 U6282 ( .B1(n7544), .B2(n7838), .A(n5969), .ZN(n5970) );
  NAND2_X1 U6283 ( .A1(n4274), .A2(n4705), .ZN(n4411) );
  NAND2_X2 U6284 ( .A1(n6252), .A2(n6247), .ZN(n7021) );
  NAND2_X1 U6285 ( .A1(n5970), .A2(n6285), .ZN(n7733) );
  NAND2_X1 U6286 ( .A1(n4870), .A2(n4872), .ZN(n7544) );
  NAND4_X1 U6287 ( .A1(n6303), .A2(n8404), .A3(n6301), .A4(n6302), .ZN(n4414)
         );
  OAI21_X1 U6288 ( .B1(n6311), .B2(n6310), .A(n4379), .ZN(n6312) );
  OAI21_X1 U6289 ( .B1(n6323), .B2(n6322), .A(n4370), .ZN(n6325) );
  AOI21_X1 U6290 ( .B1(n6335), .B2(n6337), .A(n6339), .ZN(n4836) );
  INV_X2 U6292 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5874) );
  NOR2_X4 U6293 ( .A1(n8219), .A2(n8437), .ZN(n8209) );
  NAND2_X1 U6294 ( .A1(n5812), .A2(n5811), .ZN(n6368) );
  NAND3_X1 U6295 ( .A1(n4420), .A2(n8435), .A3(n4419), .ZN(n8527) );
  NOR2_X2 U6296 ( .A1(n7230), .A2(n7389), .ZN(n4792) );
  OAI21_X1 U6297 ( .B1(n6261), .B2(n6347), .A(n6260), .ZN(n6263) );
  NAND2_X1 U6298 ( .A1(n9233), .A2(n9234), .ZN(n9232) );
  OAI21_X1 U6299 ( .B1(n9867), .B2(n5020), .A(n9288), .ZN(n4422) );
  NAND2_X1 U6300 ( .A1(n4433), .A2(n4468), .ZN(n6993) );
  NAND2_X1 U6301 ( .A1(n9863), .A2(n9864), .ZN(n9861) );
  NAND2_X1 U6302 ( .A1(n9847), .A2(n9846), .ZN(n9845) );
  OAI22_X1 U6303 ( .A1(n7239), .A2(n7238), .B1(n7245), .B2(
        P1_REG1_REG_11__SCAN_IN), .ZN(n7678) );
  AOI21_X1 U6304 ( .B1(P1_REG1_REG_5__SCAN_IN), .B2(n6657), .A(n6656), .ZN(
        n6682) );
  NAND2_X1 U6305 ( .A1(n4427), .A2(n4426), .ZN(P2_U3216) );
  NAND2_X1 U6306 ( .A1(n7902), .A2(n7901), .ZN(n4427) );
  NAND2_X1 U6307 ( .A1(n4607), .A2(n4371), .ZN(n4928) );
  INV_X1 U6308 ( .A(n4603), .ZN(n4602) );
  NAND2_X1 U6309 ( .A1(n4877), .A2(n5266), .ZN(n4549) );
  NAND2_X1 U6310 ( .A1(n4880), .A2(n4375), .ZN(n5335) );
  OAI22_X2 U6311 ( .A1(n5105), .A2(n8711), .B1(n9896), .B2(n8709), .ZN(n7074)
         );
  NAND2_X1 U6312 ( .A1(n7140), .A2(n7141), .ZN(n7142) );
  AND2_X2 U6313 ( .A1(n4648), .A2(n4649), .ZN(n4645) );
  AND2_X2 U6314 ( .A1(n5784), .A2(n5786), .ZN(n4648) );
  NAND4_X1 U6315 ( .A1(n4431), .A2(n5825), .A3(n5826), .A4(n5824), .ZN(n6384)
         );
  NAND2_X1 U6316 ( .A1(n4826), .A2(n5800), .ZN(n4825) );
  NAND2_X1 U6317 ( .A1(n6704), .A2(n4432), .ZN(n6990) );
  AND3_X2 U6318 ( .A1(n8171), .A2(n8307), .A3(n4954), .ZN(n4710) );
  NAND2_X1 U6319 ( .A1(n4435), .A2(n4434), .ZN(n7079) );
  INV_X1 U6320 ( .A(n7078), .ZN(n4435) );
  XNOR2_X1 U6321 ( .A(n7074), .B(n4468), .ZN(n7078) );
  OR2_X1 U6322 ( .A1(n5014), .A2(n4663), .ZN(n4444) );
  NAND2_X1 U6323 ( .A1(n4453), .A2(n7073), .ZN(n6706) );
  NAND2_X1 U6324 ( .A1(n8150), .A2(n4291), .ZN(n4488) );
  NAND2_X1 U6325 ( .A1(n4661), .A2(n4381), .ZN(n6303) );
  NAND2_X1 U6326 ( .A1(n6293), .A2(n7744), .ZN(n4662) );
  NAND2_X1 U6327 ( .A1(n4822), .A2(n4821), .ZN(n4820) );
  NAND2_X1 U6328 ( .A1(n4660), .A2(n6298), .ZN(n4823) );
  AND3_X1 U6329 ( .A1(n4830), .A2(n4829), .A3(n5883), .ZN(n4828) );
  NAND2_X1 U6330 ( .A1(n4833), .A2(n4388), .ZN(n4659) );
  NAND3_X1 U6331 ( .A1(n4724), .A2(n4336), .A3(n4723), .ZN(n4727) );
  NAND2_X1 U6332 ( .A1(n7743), .A2(n7742), .ZN(n7767) );
  INV_X2 U6333 ( .A(n7368), .ZN(n4446) );
  NOR2_X2 U6334 ( .A1(n6497), .A2(n6496), .ZN(n7906) );
  INV_X1 U6335 ( .A(n7947), .ZN(n4607) );
  NAND2_X1 U6336 ( .A1(n4964), .A2(n4965), .ZN(n8382) );
  NAND2_X1 U6337 ( .A1(n7052), .A2(n6406), .ZN(n7204) );
  NOR2_X1 U6338 ( .A1(n8836), .A2(n8835), .ZN(n8834) );
  NAND2_X1 U6339 ( .A1(n7258), .A2(n7259), .ZN(n7606) );
  NAND2_X1 U6340 ( .A1(n8826), .A2(n8823), .ZN(n8903) );
  NAND2_X1 U6341 ( .A1(n7635), .A2(n7634), .ZN(n7646) );
  AND4_X2 U6342 ( .A1(n5783), .A2(n5785), .A3(n5782), .A4(n4739), .ZN(n4647)
         );
  NAND2_X1 U6343 ( .A1(n7225), .A2(n4871), .ZN(n4870) );
  NAND2_X1 U6344 ( .A1(n6706), .A2(n6705), .ZN(n6991) );
  AOI21_X2 U6345 ( .B1(n8762), .B2(n8661), .A(n8660), .ZN(n8892) );
  AOI21_X2 U6346 ( .B1(n8736), .B2(n8694), .A(n4481), .ZN(n8867) );
  NAND2_X1 U6347 ( .A1(n7155), .A2(n7154), .ZN(n7257) );
  NAND2_X2 U6348 ( .A1(n4816), .A2(n4814), .ZN(n8736) );
  INV_X4 U6349 ( .A(n6992), .ZN(n4468) );
  NOR2_X2 U6350 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n5836) );
  INV_X1 U6351 ( .A(n8171), .ZN(n8327) );
  INV_X1 U6352 ( .A(n4738), .ZN(n5955) );
  AOI21_X1 U6353 ( .B1(n9283), .B2(n9282), .A(n4479), .ZN(n4478) );
  NAND2_X1 U6354 ( .A1(n6685), .A2(n6686), .ZN(n6684) );
  NOR2_X1 U6355 ( .A1(n7670), .A2(n4786), .ZN(n9817) );
  NOR2_X1 U6356 ( .A1(n9256), .A2(n9257), .ZN(n9275) );
  NAND4_X1 U6357 ( .A1(n4462), .A2(n9396), .A3(n9381), .A4(n9362), .ZN(n4461)
         );
  NOR2_X1 U6358 ( .A1(n9853), .A2(n9852), .ZN(n9851) );
  NAND3_X1 U6359 ( .A1(n4978), .A2(n9116), .A3(n9192), .ZN(n9195) );
  NOR2_X2 U6360 ( .A1(n8867), .A2(n8696), .ZN(n8836) );
  AND2_X2 U6361 ( .A1(n7606), .A2(n7605), .ZN(n7609) );
  NOR2_X2 U6362 ( .A1(n8834), .A2(n4359), .ZN(n8962) );
  NAND2_X1 U6363 ( .A1(n4453), .A2(n4465), .ZN(n6704) );
  NAND2_X1 U6364 ( .A1(n4466), .A2(n4373), .ZN(P1_U3218) );
  NAND2_X1 U6365 ( .A1(n8788), .A2(n8787), .ZN(n4466) );
  NAND2_X1 U6366 ( .A1(n5112), .A2(n5043), .ZN(n5046) );
  AOI21_X2 U6367 ( .B1(n7413), .B2(n4684), .A(n4469), .ZN(n9013) );
  NAND2_X1 U6368 ( .A1(n4666), .A2(n4665), .ZN(n4664) );
  NAND2_X1 U6369 ( .A1(n9027), .A2(n4671), .ZN(n4670) );
  INV_X1 U6370 ( .A(n7275), .ZN(n4680) );
  NAND3_X1 U6371 ( .A1(n5099), .A2(n5100), .A3(n5098), .ZN(n6985) );
  NAND2_X1 U6372 ( .A1(n6990), .A2(n6991), .ZN(n6994) );
  AOI21_X1 U6373 ( .B1(n9263), .B2(n9262), .A(n9261), .ZN(n9265) );
  NAND2_X1 U6374 ( .A1(n4659), .A2(n4657), .ZN(n6351) );
  NAND2_X1 U6375 ( .A1(n4823), .A2(n4719), .ZN(n4822) );
  NAND2_X1 U6376 ( .A1(n4662), .A2(n4385), .ZN(n4661) );
  NAND2_X1 U6377 ( .A1(n6303), .A2(n4824), .ZN(n4660) );
  NAND2_X1 U6378 ( .A1(n4820), .A2(n4819), .ZN(n6308) );
  OAI21_X1 U6379 ( .B1(n4836), .B2(n4834), .A(n6341), .ZN(n4833) );
  NAND2_X1 U6380 ( .A1(n4639), .A2(n4637), .ZN(n6335) );
  AND3_X4 U6381 ( .A1(n4645), .A2(n5851), .A3(n4647), .ZN(n6010) );
  NAND2_X1 U6382 ( .A1(n4653), .A2(n4652), .ZN(n4651) );
  NAND2_X1 U6383 ( .A1(n4727), .A2(n4726), .ZN(n7745) );
  NAND2_X1 U6384 ( .A1(n8262), .A2(n8177), .ZN(n8246) );
  AND2_X2 U6385 ( .A1(n4825), .A2(n5801), .ZN(n5804) );
  NAND2_X1 U6386 ( .A1(n5798), .A2(P2_IR_REG_29__SCAN_IN), .ZN(n4826) );
  OAI21_X1 U6387 ( .B1(n7222), .B2(n7221), .A(n7220), .ZN(n7223) );
  NAND2_X1 U6388 ( .A1(n7000), .A2(n6999), .ZN(n7082) );
  INV_X2 U6389 ( .A(n6985), .ZN(n9889) );
  NAND2_X1 U6390 ( .A1(n6684), .A2(n4386), .ZN(n6653) );
  NOR2_X1 U6391 ( .A1(n9817), .A2(n9816), .ZN(n9815) );
  NAND2_X1 U6392 ( .A1(n6642), .A2(n6615), .ZN(n4484) );
  NAND3_X1 U6393 ( .A1(n4488), .A2(n8153), .A3(n4487), .ZN(P2_U3264) );
  NOR2_X2 U6394 ( .A1(n5852), .A2(n5863), .ZN(n8082) );
  NAND2_X2 U6395 ( .A1(n6010), .A2(n5793), .ZN(n6361) );
  AOI21_X2 U6396 ( .B1(n8205), .B2(n8204), .A(n8203), .ZN(n8440) );
  OAI21_X1 U6397 ( .B1(n8238), .B2(n4576), .A(n4556), .ZN(n8200) );
  NOR2_X2 U6398 ( .A1(n5017), .A2(n4759), .ZN(n5003) );
  NAND2_X1 U6399 ( .A1(n6997), .A2(n6998), .ZN(n7002) );
  NAND3_X1 U6400 ( .A1(n4489), .A2(n8721), .A3(n4395), .ZN(P1_U3212) );
  OAI21_X1 U6401 ( .B1(n8718), .B2(n8786), .A(n8959), .ZN(n4489) );
  NAND2_X1 U6402 ( .A1(n8962), .A2(n8961), .ZN(n8960) );
  OAI21_X1 U6403 ( .B1(n9032), .B2(n4668), .A(n4667), .ZN(n4666) );
  NAND2_X1 U6404 ( .A1(n5014), .A2(n4999), .ZN(n5015) );
  NAND2_X1 U6405 ( .A1(n4672), .A2(n4382), .ZN(n9072) );
  NAND2_X1 U6406 ( .A1(n4664), .A2(n9152), .ZN(n9038) );
  NAND2_X1 U6407 ( .A1(n4676), .A2(n9066), .ZN(n4675) );
  NAND2_X1 U6408 ( .A1(n4694), .A2(n4697), .ZN(n9057) );
  INV_X1 U6409 ( .A(n7342), .ZN(n5190) );
  NAND2_X1 U6410 ( .A1(n7305), .A2(n9098), .ZN(n4493) );
  NAND2_X1 U6411 ( .A1(n5168), .A2(n5167), .ZN(n7305) );
  NAND2_X1 U6412 ( .A1(n4494), .A2(n4496), .ZN(n4847) );
  NAND2_X1 U6413 ( .A1(n9471), .A2(n4500), .ZN(n4494) );
  NAND2_X2 U6414 ( .A1(n4304), .A2(n4346), .ZN(n4500) );
  NAND2_X1 U6415 ( .A1(n9299), .A2(n9597), .ZN(n9300) );
  NAND3_X1 U6416 ( .A1(n5192), .A2(n5193), .A3(n4334), .ZN(n4503) );
  NAND3_X1 U6417 ( .A1(n5192), .A2(n5193), .A3(n4507), .ZN(n4506) );
  NAND3_X1 U6418 ( .A1(n5192), .A2(n5193), .A3(n4509), .ZN(n7486) );
  NAND2_X1 U6419 ( .A1(n9534), .A2(n4513), .ZN(n4511) );
  NAND2_X1 U6420 ( .A1(n9376), .A2(n4524), .ZN(n4520) );
  NAND2_X1 U6421 ( .A1(n4520), .A2(n4521), .ZN(n5644) );
  INV_X1 U6422 ( .A(n9172), .ZN(n4529) );
  NAND2_X1 U6423 ( .A1(n9514), .A2(n9153), .ZN(n4751) );
  NAND2_X1 U6424 ( .A1(n4534), .A2(n4398), .ZN(n9599) );
  NAND2_X1 U6425 ( .A1(n9706), .A2(n9970), .ZN(n4533) );
  NAND4_X1 U6426 ( .A1(n4534), .A2(n9600), .A3(n4398), .A4(n9601), .ZN(n9706)
         );
  NAND2_X1 U6427 ( .A1(n9461), .A2(n4538), .ZN(n4535) );
  NAND2_X1 U6428 ( .A1(n4535), .A2(n4536), .ZN(n9392) );
  MUX2_X1 U6429 ( .A(n6581), .B(n6569), .S(n4279), .Z(n5062) );
  NAND3_X1 U6430 ( .A1(n4844), .A2(P1_ADDR_REG_19__SCAN_IN), .A3(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n4542) );
  NAND3_X1 U6431 ( .A1(n5020), .A2(n4545), .A3(n4544), .ZN(n4543) );
  AND2_X2 U6432 ( .A1(n4892), .A2(n4891), .ZN(n8286) );
  NAND2_X2 U6433 ( .A1(n4733), .A2(n4734), .ZN(n8238) );
  XNOR2_X2 U6434 ( .A(n4561), .B(P1_IR_REG_3__SCAN_IN), .ZN(n6626) );
  INV_X1 U6435 ( .A(n9256), .ZN(n4564) );
  NAND2_X1 U6436 ( .A1(n9252), .A2(n4569), .ZN(n4568) );
  INV_X1 U6437 ( .A(n4572), .ZN(n9827) );
  AOI21_X2 U6438 ( .B1(n8222), .B2(n6138), .A(n6137), .ZN(n8239) );
  NAND2_X1 U6439 ( .A1(n5937), .A2(n4322), .ZN(n5974) );
  NAND2_X1 U6440 ( .A1(n6018), .A2(n4582), .ZN(n6053) );
  INV_X1 U6441 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n4585) );
  NAND2_X1 U6442 ( .A1(n6061), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n6074) );
  INV_X1 U6443 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n4588) );
  NAND2_X1 U6444 ( .A1(n4915), .A2(n4596), .ZN(n4592) );
  NAND2_X1 U6445 ( .A1(n4592), .A2(n4589), .ZN(n6465) );
  NAND2_X1 U6446 ( .A1(n4913), .A2(n4602), .ZN(n4599) );
  NAND2_X1 U6447 ( .A1(n4599), .A2(n4600), .ZN(n6488) );
  NAND2_X1 U6448 ( .A1(n7402), .A2(n6430), .ZN(n6431) );
  AND2_X2 U6449 ( .A1(n4928), .A2(n4926), .ZN(n8024) );
  NAND2_X1 U6450 ( .A1(n4279), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n4609) );
  NAND2_X1 U6451 ( .A1(n5560), .A2(n4617), .ZN(n4616) );
  OR2_X1 U6452 ( .A1(n5560), .A2(n5559), .ZN(n4621) );
  OR2_X1 U6453 ( .A1(n6334), .A2(n6349), .ZN(n4638) );
  NAND2_X1 U6454 ( .A1(n4640), .A2(n4390), .ZN(n4639) );
  NAND2_X1 U6455 ( .A1(n4641), .A2(n4837), .ZN(n4640) );
  NAND3_X1 U6456 ( .A1(n4843), .A2(n4842), .A3(n4389), .ZN(n4641) );
  NAND3_X1 U6457 ( .A1(n6282), .A2(n6273), .A3(n6274), .ZN(n4642) );
  NAND2_X1 U6458 ( .A1(n4651), .A2(n4650), .ZN(n6354) );
  NAND2_X1 U6459 ( .A1(n6351), .A2(n6346), .ZN(n4653) );
  NAND2_X1 U6460 ( .A1(n6348), .A2(n6344), .ZN(n4658) );
  NAND3_X1 U6461 ( .A1(n9075), .A2(n9073), .A3(n9074), .ZN(n4687) );
  NAND4_X1 U6462 ( .A1(n9045), .A2(n9170), .A3(n4697), .A4(n4696), .ZN(n4691)
         );
  NOR2_X1 U6463 ( .A1(n9044), .A2(n9482), .ZN(n4699) );
  NAND2_X1 U6464 ( .A1(n5050), .A2(n4701), .ZN(n4700) );
  NAND2_X1 U6465 ( .A1(n4856), .A2(n5048), .ZN(n5160) );
  INV_X1 U6466 ( .A(n5048), .ZN(n4701) );
  NAND2_X1 U6467 ( .A1(n8217), .A2(n4321), .ZN(n4705) );
  NAND2_X1 U6468 ( .A1(n8440), .A2(n8439), .ZN(n4706) );
  INV_X1 U6469 ( .A(n4954), .ZN(n4714) );
  NAND2_X1 U6470 ( .A1(n4715), .A2(n4716), .ZN(n8171) );
  NAND2_X1 U6471 ( .A1(n8382), .A2(n4312), .ZN(n4715) );
  NAND3_X1 U6472 ( .A1(n4724), .A2(n7740), .A3(n4723), .ZN(n7837) );
  INV_X1 U6473 ( .A(n7745), .ZN(n7743) );
  OR2_X1 U6474 ( .A1(n7885), .A2(n8062), .ZN(n4728) );
  OR2_X2 U6475 ( .A1(n8269), .A2(n4735), .ZN(n4733) );
  NAND3_X1 U6476 ( .A1(n4743), .A2(n5075), .A3(n4987), .ZN(n5021) );
  NAND2_X1 U6477 ( .A1(n4751), .A2(n4753), .ZN(n9480) );
  XNOR2_X1 U6478 ( .A(n4758), .B(n4757), .ZN(n7425) );
  INV_X1 U6479 ( .A(n9090), .ZN(n4757) );
  NAND2_X1 U6480 ( .A1(n9331), .A2(n4383), .ZN(n9326) );
  NAND2_X1 U6481 ( .A1(n7297), .A2(n7292), .ZN(n7295) );
  NAND2_X1 U6482 ( .A1(n8209), .A2(n8431), .ZN(n8191) );
  NAND3_X1 U6483 ( .A1(n4774), .A2(n4775), .A3(n4776), .ZN(n8425) );
  NAND3_X1 U6484 ( .A1(n4775), .A2(n4774), .A3(n4773), .ZN(n4780) );
  OR2_X1 U6485 ( .A1(n8209), .A2(n4656), .ZN(n4774) );
  NAND2_X1 U6486 ( .A1(n8209), .A2(n4778), .ZN(n4775) );
  XNOR2_X1 U6487 ( .A(n5129), .B(P1_IR_REG_2__SCAN_IN), .ZN(n9238) );
  NAND2_X1 U6488 ( .A1(n7646), .A2(n4798), .ZN(n4797) );
  NAND2_X1 U6489 ( .A1(n8903), .A2(n4809), .ZN(n4807) );
  AND2_X2 U6490 ( .A1(n8960), .A2(n4378), .ZN(n8786) );
  NAND3_X1 U6491 ( .A1(n4995), .A2(n4994), .A3(n5377), .ZN(n4817) );
  NOR2_X2 U6492 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n5785) );
  NAND3_X1 U6493 ( .A1(n5793), .A2(n6010), .A3(n4972), .ZN(n5815) );
  NAND2_X2 U6494 ( .A1(n4828), .A2(n5882), .ZN(n8066) );
  NAND4_X1 U6495 ( .A1(n6325), .A2(n6324), .A3(n6347), .A4(n6091), .ZN(n4842)
         );
  NAND4_X1 U6496 ( .A1(n6312), .A2(n6313), .A3(n6349), .A4(n6320), .ZN(n4843)
         );
  OAI21_X1 U6497 ( .B1(n9397), .B2(n4851), .A(n4848), .ZN(n9345) );
  NAND2_X1 U6498 ( .A1(n4847), .A2(n4377), .ZN(n5557) );
  NAND2_X1 U6499 ( .A1(n5764), .A2(n4392), .ZN(n9596) );
  OR2_X2 U6500 ( .A1(n9318), .A2(n9069), .ZN(n5764) );
  NAND2_X1 U6501 ( .A1(n4864), .A2(n4863), .ZN(n7029) );
  NOR2_X2 U6502 ( .A1(n6358), .A2(n5792), .ZN(n5793) );
  NAND4_X1 U6503 ( .A1(n5788), .A2(n5789), .A3(n5790), .A4(n5791), .ZN(n6358)
         );
  NAND2_X1 U6504 ( .A1(n7771), .A2(n4869), .ZN(n7769) );
  NAND2_X1 U6506 ( .A1(n5060), .A2(n4878), .ZN(n4877) );
  INV_X1 U6507 ( .A(n4892), .ZN(n8304) );
  NAND2_X1 U6508 ( .A1(n4906), .A2(n4905), .ZN(n6315) );
  NOR2_X1 U6509 ( .A1(n8169), .A2(n4904), .ZN(n4905) );
  NAND2_X2 U6510 ( .A1(n8015), .A2(n8016), .ZN(n4913) );
  AND2_X1 U6511 ( .A1(n6432), .A2(n6427), .ZN(n4916) );
  NAND2_X1 U6512 ( .A1(n6050), .A2(n4917), .ZN(n6187) );
  NAND2_X1 U6513 ( .A1(n7204), .A2(n4919), .ZN(n7064) );
  NAND2_X1 U6514 ( .A1(n7064), .A2(n6416), .ZN(n6421) );
  NAND2_X1 U6515 ( .A1(n6223), .A2(n7368), .ZN(n6381) );
  XNOR2_X2 U6516 ( .A(n6194), .B(n6195), .ZN(n6223) );
  INV_X1 U6517 ( .A(n6223), .ZN(n6370) );
  NAND2_X1 U6518 ( .A1(n4928), .A2(n4929), .ZN(n8025) );
  INV_X1 U6519 ( .A(n7944), .ZN(n4930) );
  NAND2_X1 U6520 ( .A1(n4994), .A2(n4387), .ZN(n4935) );
  NAND4_X1 U6522 ( .A1(n4995), .A2(n4934), .A3(n5671), .A4(n5377), .ZN(n5016)
         );
  NAND3_X1 U6523 ( .A1(n4937), .A2(n4936), .A3(n4938), .ZN(n5746) );
  NAND2_X1 U6524 ( .A1(n9319), .A2(n4384), .ZN(n4936) );
  NAND2_X1 U6525 ( .A1(n9319), .A2(n9590), .ZN(n9302) );
  AND2_X2 U6526 ( .A1(n9520), .A2(n4947), .ZN(n9474) );
  XNOR2_X1 U6527 ( .A(n4956), .B(n8318), .ZN(n8475) );
  NAND2_X1 U6528 ( .A1(n4960), .A2(n4961), .ZN(n8183) );
  NAND2_X1 U6529 ( .A1(n8218), .A2(n4305), .ZN(n4960) );
  NAND2_X1 U6530 ( .A1(n8218), .A2(n8225), .ZN(n8217) );
  OAI21_X2 U6531 ( .B1(n8218), .B2(n4963), .A(n4305), .ZN(n8206) );
  NAND2_X1 U6532 ( .A1(n7794), .A2(n4966), .ZN(n4964) );
  NAND2_X1 U6533 ( .A1(n8280), .A2(n4970), .ZN(n8262) );
  NAND2_X1 U6534 ( .A1(n7767), .A2(n4344), .ZN(n7792) );
  NAND3_X1 U6535 ( .A1(n6010), .A2(n4973), .A3(n5793), .ZN(n5801) );
  XNOR2_X1 U6536 ( .A(n5713), .B(n5712), .ZN(n7833) );
  XNOR2_X2 U6537 ( .A(n5097), .B(P1_IR_REG_1__SCAN_IN), .ZN(n6642) );
  OR2_X1 U6538 ( .A1(n5764), .A2(n5762), .ZN(n5623) );
  NAND2_X1 U6539 ( .A1(n5707), .A2(n9986), .ZN(n5703) );
  NAND2_X1 U6540 ( .A1(n6994), .A2(n6993), .ZN(n6997) );
  OAI211_X2 U6541 ( .C1(n5835), .C2(n5166), .A(n5077), .B(n5076), .ZN(n7282)
         );
  AND2_X1 U6542 ( .A1(n9596), .A2(n4979), .ZN(n9601) );
  XNOR2_X1 U6543 ( .A(n9309), .B(n9598), .ZN(n9312) );
  AND2_X1 U6544 ( .A1(n7034), .A2(n7033), .ZN(n8305) );
  XNOR2_X1 U6545 ( .A(n4283), .B(n7923), .ZN(n6394) );
  OR2_X1 U6546 ( .A1(n4492), .A2(n4610), .ZN(n5165) );
  NAND2_X1 U6547 ( .A1(n6384), .A2(n7861), .ZN(n7018) );
  OR2_X1 U6548 ( .A1(n6000), .A2(n5027), .ZN(n5854) );
  INV_X1 U6549 ( .A(n5803), .ZN(n5805) );
  MUX2_X1 U6550 ( .A(P1_IR_REG_0__SCAN_IN), .B(n9766), .S(n5451), .Z(n7292) );
  AOI22_X2 U6551 ( .A1(n6500), .A2(n7970), .B1(n7972), .B2(n7974), .ZN(n7947)
         );
  INV_X1 U6552 ( .A(n9701), .ZN(n5698) );
  AND2_X1 U6553 ( .A1(n5317), .A2(n5296), .ZN(n4974) );
  AND2_X1 U6554 ( .A1(n5376), .A2(n5361), .ZN(n4975) );
  OR2_X1 U6555 ( .A1(n8793), .A2(n8986), .ZN(n4976) );
  NAND2_X2 U6556 ( .A1(n5771), .A2(n9538), .ZN(n9541) );
  OR2_X1 U6557 ( .A1(n8285), .A2(n8272), .ZN(n4977) );
  AND4_X1 U6558 ( .A1(n9588), .A2(n9113), .A3(n9112), .A4(n9336), .ZN(n4978)
         );
  NAND2_X1 U6559 ( .A1(n9970), .A2(n9913), .ZN(n9751) );
  INV_X1 U6560 ( .A(n9751), .ZN(n5759) );
  INV_X1 U6561 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n5053) );
  INV_X1 U6562 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n5049) );
  INV_X1 U6563 ( .A(n10024), .ZN(n8396) );
  OR3_X1 U6564 ( .A1(n4281), .A2(n10089), .A3(n4301), .ZN(n10024) );
  NOR2_X1 U6565 ( .A1(n9595), .A2(n9594), .ZN(n4979) );
  OR2_X1 U6566 ( .A1(n8202), .A2(n8041), .ZN(n4980) );
  OR2_X1 U6567 ( .A1(n8330), .A2(n8172), .ZN(n4982) );
  NAND2_X1 U6568 ( .A1(n9435), .A2(n9456), .ZN(n4983) );
  INV_X1 U6569 ( .A(n7451), .ZN(n7172) );
  AND3_X1 U6570 ( .A1(n9598), .A2(n9966), .A3(n9597), .ZN(n4985) );
  INV_X1 U6571 ( .A(n9298), .ZN(n9590) );
  NOR2_X1 U6572 ( .A1(n9497), .A2(n9495), .ZN(n4986) );
  INV_X1 U6573 ( .A(n7412), .ZN(n5630) );
  INV_X1 U6574 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n4991) );
  INV_X1 U6575 ( .A(n7562), .ZN(n6432) );
  INV_X1 U6576 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5794) );
  OAI21_X1 U6577 ( .B1(n8876), .B2(n8800), .A(n8797), .ZN(n8562) );
  NOR2_X1 U6578 ( .A1(n8999), .A2(n9311), .ZN(n9000) );
  INV_X1 U6579 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n5357) );
  AND2_X1 U6580 ( .A1(n5183), .A2(n5143), .ZN(n5052) );
  INV_X1 U6581 ( .A(n7062), .ZN(n6415) );
  INV_X1 U6582 ( .A(n8562), .ZN(n8563) );
  NOR2_X1 U6583 ( .A1(n9915), .A2(n9902), .ZN(n5628) );
  INV_X1 U6584 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n4999) );
  INV_X1 U6585 ( .A(SI_22_), .ZN(n10251) );
  NOR2_X1 U6586 ( .A1(n5414), .A2(n5413), .ZN(n5425) );
  NAND2_X1 U6587 ( .A1(n4287), .A2(P2_DATAO_REG_7__SCAN_IN), .ZN(n5054) );
  INV_X1 U6588 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5114) );
  AND2_X1 U6589 ( .A1(n6498), .A2(n6499), .ZN(n6495) );
  INV_X1 U6590 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n10237) );
  NAND2_X1 U6591 ( .A1(n5868), .A2(n10062), .ZN(n6205) );
  INV_X1 U6592 ( .A(n6381), .ZN(n6512) );
  INV_X1 U6593 ( .A(n7744), .ZN(n7742) );
  INV_X1 U6594 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n10248) );
  INV_X1 U6595 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n5252) );
  NAND2_X1 U6596 ( .A1(n7609), .A2(n4345), .ZN(n7635) );
  AND2_X1 U6597 ( .A1(n5346), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n5366) );
  INV_X1 U6598 ( .A(n9497), .ZN(n9500) );
  NAND2_X1 U6599 ( .A1(n9029), .A2(n9151), .ZN(n9104) );
  NAND2_X1 U6600 ( .A1(n5430), .A2(n5429), .ZN(n5469) );
  NAND2_X1 U6601 ( .A1(n5359), .A2(n5358), .ZN(n5376) );
  OR2_X1 U6602 ( .A1(n6538), .A2(n6537), .ZN(n6539) );
  OR2_X1 U6603 ( .A1(n7068), .A2(n7370), .ZN(n6544) );
  OR2_X1 U6604 ( .A1(n7938), .A2(n6076), .ZN(n6082) );
  INV_X1 U6605 ( .A(n6958), .ZN(n6383) );
  INV_X1 U6606 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n7406) );
  INV_X1 U6607 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n7996) );
  INV_X1 U6608 ( .A(n8452), .ZN(n8253) );
  AND2_X1 U6609 ( .A1(n6370), .A2(n4446), .ZN(n6665) );
  AND2_X1 U6610 ( .A1(n10029), .A2(n7372), .ZN(n7373) );
  NAND2_X1 U6611 ( .A1(n4301), .A2(n8392), .ZN(n6545) );
  INV_X1 U6612 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n8545) );
  NAND2_X1 U6613 ( .A1(n5366), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n5386) );
  AND2_X1 U6614 ( .A1(n6708), .A2(n6707), .ZN(n7006) );
  INV_X1 U6615 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n8904) );
  OR2_X1 U6616 ( .A1(n9603), .A2(n9333), .ZN(n5763) );
  AND2_X1 U6617 ( .A1(n9177), .A2(n9050), .ZN(n9362) );
  AND2_X1 U6618 ( .A1(n9170), .A2(n9087), .ZN(n9396) );
  INV_X1 U6619 ( .A(n9544), .ZN(n9576) );
  INV_X1 U6620 ( .A(n9986), .ZN(n5699) );
  AND2_X1 U6621 ( .A1(n9114), .A2(n5753), .ZN(n9584) );
  INV_X1 U6622 ( .A(n9535), .ZN(n9569) );
  INV_X1 U6623 ( .A(n8559), .ZN(n9953) );
  NAND2_X1 U6624 ( .A1(n8989), .A2(n9121), .ZN(n9943) );
  NOR2_X1 U6625 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n10288), .ZN(n9782) );
  INV_X1 U6626 ( .A(n8041), .ZN(n8018) );
  INV_X1 U6627 ( .A(n8032), .ZN(n8048) );
  OR2_X1 U6628 ( .A1(n5858), .A2(n8083), .ZN(n5845) );
  AND2_X1 U6629 ( .A1(n6726), .A2(n6725), .ZN(n10005) );
  INV_X1 U6630 ( .A(n9988), .ZN(n10003) );
  INV_X1 U6631 ( .A(n8407), .ZN(n8372) );
  AND2_X1 U6632 ( .A1(n6286), .A2(n6285), .ZN(n7843) );
  NAND2_X1 U6633 ( .A1(n10029), .A2(n6532), .ZN(n10022) );
  NOR2_X1 U6634 ( .A1(n7068), .A2(n7371), .ZN(n7069) );
  NAND2_X1 U6635 ( .A1(n6512), .A2(n6545), .ZN(n10077) );
  INV_X1 U6636 ( .A(n7557), .ZN(n10083) );
  AND2_X1 U6637 ( .A1(n6223), .A2(n6531), .ZN(n10084) );
  NAND2_X1 U6638 ( .A1(n10014), .A2(n8518), .ZN(n10086) );
  AND2_X1 U6639 ( .A1(n6718), .A2(n10038), .ZN(n10029) );
  AND2_X1 U6640 ( .A1(n9313), .A2(n5605), .ZN(n8792) );
  INV_X1 U6641 ( .A(n8980), .ZN(n8894) );
  INV_X1 U6642 ( .A(n8981), .ZN(n8941) );
  INV_X1 U6643 ( .A(n8993), .ZN(n9118) );
  INV_X1 U6644 ( .A(n5777), .ZN(n5778) );
  INV_X1 U6645 ( .A(n9943), .ZN(n9914) );
  INV_X1 U6646 ( .A(n9513), .ZN(n9582) );
  INV_X1 U6647 ( .A(n9882), .ZN(n6708) );
  INV_X1 U6648 ( .A(n9961), .ZN(n9913) );
  AND2_X1 U6649 ( .A1(n5704), .A2(n9884), .ZN(n5767) );
  INV_X1 U6650 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n5000) );
  XNOR2_X1 U6651 ( .A(n5182), .B(n5180), .ZN(n6565) );
  INV_X1 U6652 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n9772) );
  AND2_X1 U6653 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n9792), .ZN(n9793) );
  NAND2_X1 U6654 ( .A1(n6667), .A2(n6666), .ZN(n9997) );
  INV_X1 U6655 ( .A(n8441), .ZN(n8224) );
  OR2_X1 U6656 ( .A1(n7826), .A2(n8407), .ZN(n8041) );
  NAND2_X2 U6657 ( .A1(n6534), .A2(n6533), .ZN(n8044) );
  NOR2_X1 U6658 ( .A1(n6378), .A2(n4981), .ZN(n6379) );
  INV_X1 U6659 ( .A(n8408), .ZN(n8371) );
  INV_X1 U6660 ( .A(n7881), .ZN(n8061) );
  INV_X1 U6661 ( .A(n10005), .ZN(n9989) );
  OR2_X1 U6662 ( .A1(n10023), .A2(n4296), .ZN(n8192) );
  OR2_X1 U6663 ( .A1(n7705), .A2(n7541), .ZN(n7557) );
  INV_X1 U6664 ( .A(n10100), .ZN(n10098) );
  OR2_X1 U6665 ( .A1(n8499), .A2(n8498), .ZN(n8539) );
  INV_X1 U6666 ( .A(n10283), .ZN(n10281) );
  INV_X1 U6667 ( .A(n10035), .ZN(n10033) );
  INV_X1 U6668 ( .A(n10032), .ZN(n10038) );
  INV_X1 U6669 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n10263) );
  INV_X1 U6670 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n7108) );
  INV_X1 U6671 ( .A(n8566), .ZN(n9962) );
  OR2_X1 U6672 ( .A1(n8958), .A2(n9961), .ZN(n8981) );
  INV_X1 U6673 ( .A(n9609), .ZN(n9364) );
  INV_X1 U6674 ( .A(n9684), .ZN(n9543) );
  INV_X1 U6675 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n9773) );
  INV_X1 U6676 ( .A(n9855), .ZN(n9839) );
  OR2_X1 U6677 ( .A1(n9802), .A2(n6605), .ZN(n9281) );
  INV_X1 U6678 ( .A(n9810), .ZN(n9867) );
  NAND2_X1 U6679 ( .A1(n9541), .A2(n7299), .ZN(n9513) );
  NAND2_X1 U6680 ( .A1(n9986), .A2(n9913), .ZN(n9701) );
  AND2_X2 U6681 ( .A1(n5696), .A2(n6708), .ZN(n9986) );
  INV_X1 U6682 ( .A(n9369), .ZN(n9718) );
  INV_X1 U6683 ( .A(n9506), .ZN(n9737) );
  AND4_X1 U6684 ( .A1(n9909), .A2(n9908), .A3(n9907), .A4(n9906), .ZN(n9975)
         );
  INV_X1 U6685 ( .A(n9970), .ZN(n9968) );
  AND2_X1 U6686 ( .A1(n9884), .A2(n9879), .ZN(n9880) );
  INV_X1 U6687 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n6863) );
  CLKBUF_X1 U6688 ( .A(n9765), .Z(n7782) );
  NOR2_X1 U6689 ( .A1(n10298), .A2(n10297), .ZN(n10296) );
  NOR2_X1 U6690 ( .A1(n10129), .A2(n10128), .ZN(n10127) );
  INV_X2 U6691 ( .A(n8056), .ZN(P2_U3966) );
  INV_X2 U6692 ( .A(n9230), .ZN(P1_U4006) );
  OR2_X1 U6693 ( .A1(n5781), .A2(n5780), .ZN(P1_U3263) );
  NAND2_X1 U6694 ( .A1(n5703), .A2(n5702), .ZN(P1_U3551) );
  INV_X1 U6695 ( .A(n5021), .ZN(n4995) );
  NOR2_X1 U6696 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n4990) );
  NOR2_X2 U6697 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n4989) );
  NAND4_X1 U6698 ( .A1(n4990), .A2(n4989), .A3(n4988), .A4(n5200), .ZN(n5297)
         );
  NAND4_X1 U6699 ( .A1(n4992), .A2(n5340), .A3(n5302), .A4(n4991), .ZN(n4993)
         );
  NOR2_X2 U6700 ( .A1(n5297), .A2(n4993), .ZN(n5377) );
  NOR3_X2 U6701 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .A3(
        P1_IR_REG_17__SCAN_IN), .ZN(n4994) );
  NOR3_X1 U6702 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(P1_IR_REG_25__SCAN_IN), .A3(
        P1_IR_REG_27__SCAN_IN), .ZN(n4997) );
  INV_X1 U6703 ( .A(n4997), .ZN(n4998) );
  NAND2_X1 U6704 ( .A1(n5015), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5002) );
  INV_X1 U6705 ( .A(n5003), .ZN(n9753) );
  AND2_X2 U6706 ( .A1(n9758), .A2(n5005), .ZN(n5150) );
  NAND2_X1 U6707 ( .A1(n8994), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5013) );
  NAND2_X1 U6708 ( .A1(n8995), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n5012) );
  NAND2_X1 U6709 ( .A1(n5136), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5170) );
  NAND2_X1 U6710 ( .A1(n5006), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n5209) );
  INV_X1 U6711 ( .A(n5006), .ZN(n5172) );
  INV_X1 U6712 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n5007) );
  NAND2_X1 U6713 ( .A1(n5172), .A2(n5007), .ZN(n5008) );
  AND2_X1 U6714 ( .A1(n5209), .A2(n5008), .ZN(n8809) );
  NAND2_X1 U6715 ( .A1(n4467), .A2(n8809), .ZN(n5011) );
  BUF_X2 U6716 ( .A(n5441), .Z(n5747) );
  NAND2_X1 U6717 ( .A1(n5747), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n5010) );
  NAND2_X2 U6718 ( .A1(n5017), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5669) );
  OAI21_X1 U6719 ( .B1(P1_IR_REG_26__SCAN_IN), .B2(P1_IR_REG_25__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5018) );
  XNOR2_X2 U6720 ( .A(n5019), .B(P1_IR_REG_27__SCAN_IN), .ZN(n5751) );
  OR2_X1 U6721 ( .A1(n5201), .A2(n9752), .ZN(n5023) );
  XNOR2_X1 U6722 ( .A(n5023), .B(n5200), .ZN(n6870) );
  OAI22_X1 U6723 ( .A1(n4492), .A2(n6581), .B1(n4491), .B2(n6870), .ZN(n5024)
         );
  INV_X1 U6724 ( .A(n5024), .ZN(n5066) );
  INV_X1 U6725 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n5026) );
  INV_X1 U6726 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6564) );
  NAND2_X1 U6727 ( .A1(n4286), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n5028) );
  INV_X1 U6728 ( .A(SI_2_), .ZN(n5071) );
  OAI211_X1 U6729 ( .C1(n6561), .C2(n6564), .A(n5028), .B(n5071), .ZN(n5039)
         );
  AND2_X1 U6730 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n5084) );
  INV_X1 U6731 ( .A(n5084), .ZN(n5031) );
  INV_X1 U6732 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6572) );
  NAND2_X1 U6733 ( .A1(n5031), .A2(n6572), .ZN(n5029) );
  NAND2_X1 U6734 ( .A1(n5029), .A2(SI_1_), .ZN(n5030) );
  OAI21_X1 U6735 ( .B1(n5031), .B2(n6572), .A(n5030), .ZN(n5032) );
  NAND2_X1 U6736 ( .A1(n4286), .A2(n5032), .ZN(n5038) );
  AND2_X1 U6737 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n5090) );
  INV_X1 U6738 ( .A(n5090), .ZN(n5035) );
  INV_X1 U6739 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6567) );
  NAND2_X1 U6740 ( .A1(n5035), .A2(n6567), .ZN(n5033) );
  NAND2_X1 U6741 ( .A1(n5033), .A2(SI_1_), .ZN(n5034) );
  OAI21_X1 U6742 ( .B1(n5035), .B2(n6567), .A(n5034), .ZN(n5036) );
  NAND2_X1 U6743 ( .A1(n5025), .A2(n5036), .ZN(n5037) );
  NAND2_X1 U6744 ( .A1(n5039), .A2(n5072), .ZN(n5042) );
  INV_X1 U6745 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6583) );
  NAND2_X1 U6746 ( .A1(n4286), .A2(n6583), .ZN(n5040) );
  OAI211_X1 U6747 ( .C1(n6561), .C2(P1_DATAO_REG_2__SCAN_IN), .A(n5040), .B(
        SI_2_), .ZN(n5041) );
  NAND2_X1 U6748 ( .A1(n5044), .A2(SI_3_), .ZN(n5045) );
  NAND2_X1 U6749 ( .A1(n5047), .A2(SI_4_), .ZN(n5048) );
  INV_X1 U6750 ( .A(n5159), .ZN(n5050) );
  MUX2_X1 U6751 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n6561), .Z(n5144) );
  NAND2_X1 U6752 ( .A1(n5144), .A2(SI_6_), .ZN(n5183) );
  NAND2_X1 U6753 ( .A1(n5051), .A2(SI_5_), .ZN(n5143) );
  XNOR2_X1 U6754 ( .A(n5058), .B(SI_7_), .ZN(n5185) );
  NOR2_X1 U6755 ( .A1(n5144), .A2(SI_6_), .ZN(n5056) );
  NOR2_X1 U6756 ( .A1(n5185), .A2(n5056), .ZN(n5057) );
  NAND2_X1 U6757 ( .A1(n5058), .A2(SI_7_), .ZN(n5059) );
  INV_X1 U6758 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6569) );
  INV_X1 U6759 ( .A(SI_8_), .ZN(n5061) );
  NAND2_X1 U6760 ( .A1(n5062), .A2(n5061), .ZN(n5239) );
  INV_X1 U6761 ( .A(n5062), .ZN(n5063) );
  NAND2_X1 U6762 ( .A1(n5063), .A2(SI_8_), .ZN(n5064) );
  NAND2_X1 U6763 ( .A1(n5239), .A2(n5064), .ZN(n5195) );
  NAND2_X1 U6764 ( .A1(n6568), .A2(n5584), .ZN(n5065) );
  NAND2_X1 U6765 ( .A1(n5066), .A2(n5065), .ZN(n8559) );
  INV_X2 U6766 ( .A(n5523), .ZN(n5149) );
  NAND2_X1 U6767 ( .A1(n5149), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5070) );
  NAND2_X1 U6768 ( .A1(n5150), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5069) );
  NAND2_X1 U6769 ( .A1(n5652), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n5068) );
  NAND2_X1 U6770 ( .A1(n5441), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5067) );
  MUX2_X1 U6771 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .S(n6561), .Z(n5073) );
  INV_X2 U6772 ( .A(n5451), .ZN(n6555) );
  NAND2_X1 U6773 ( .A1(n6555), .A2(n4477), .ZN(n5076) );
  NAND2_X1 U6774 ( .A1(n5105), .A2(n7282), .ZN(n5627) );
  NAND2_X1 U6775 ( .A1(n9229), .A2(n9896), .ZN(n9130) );
  NAND2_X1 U6776 ( .A1(n5149), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5081) );
  NAND2_X1 U6777 ( .A1(n5150), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5080) );
  NAND2_X1 U6778 ( .A1(n5652), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n5079) );
  NAND2_X1 U6779 ( .A1(n5441), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n5078) );
  INV_X1 U6780 ( .A(SI_0_), .ZN(n5083) );
  INV_X1 U6781 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5082) );
  OAI21_X1 U6782 ( .B1(n6562), .B2(n5083), .A(n5082), .ZN(n5085) );
  NAND2_X1 U6783 ( .A1(n4286), .A2(n5084), .ZN(n5091) );
  AND2_X1 U6784 ( .A1(n5085), .A2(n5091), .ZN(n9766) );
  NAND2_X1 U6785 ( .A1(n4453), .A2(n7292), .ZN(n5102) );
  NAND2_X1 U6786 ( .A1(n5149), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n5089) );
  NAND2_X1 U6787 ( .A1(n5150), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n5088) );
  NAND2_X1 U6788 ( .A1(n5441), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5086) );
  INV_X1 U6789 ( .A(n9231), .ZN(n7274) );
  NAND2_X1 U6790 ( .A1(n5102), .A2(n7274), .ZN(n5101) );
  NAND2_X1 U6791 ( .A1(n4297), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n5100) );
  NAND2_X1 U6792 ( .A1(n4279), .A2(n5090), .ZN(n5829) );
  NAND2_X1 U6793 ( .A1(n5091), .A2(n5829), .ZN(n5093) );
  INV_X1 U6794 ( .A(SI_1_), .ZN(n5092) );
  XNOR2_X1 U6795 ( .A(n5093), .B(n5092), .ZN(n5095) );
  MUX2_X1 U6796 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .S(n6561), .Z(n5094) );
  XNOR2_X1 U6797 ( .A(n5095), .B(n5094), .ZN(n6573) );
  INV_X1 U6798 ( .A(n6573), .ZN(n5096) );
  NAND2_X1 U6799 ( .A1(n5399), .A2(n5096), .ZN(n5099) );
  NAND2_X1 U6800 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5097) );
  NAND2_X1 U6801 ( .A1(n6555), .A2(n6642), .ZN(n5098) );
  NAND2_X1 U6802 ( .A1(n5101), .A2(n7300), .ZN(n5104) );
  INV_X1 U6803 ( .A(n5102), .ZN(n7291) );
  NAND2_X1 U6804 ( .A1(n7291), .A2(n9231), .ZN(n5103) );
  NAND3_X1 U6805 ( .A1(n9093), .A2(n5104), .A3(n5103), .ZN(n5107) );
  NAND2_X1 U6806 ( .A1(n5105), .A2(n9896), .ZN(n5106) );
  NAND2_X1 U6807 ( .A1(n5107), .A2(n5106), .ZN(n7432) );
  NAND2_X1 U6808 ( .A1(n5149), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n5111) );
  NAND2_X1 U6809 ( .A1(n5150), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n5110) );
  INV_X1 U6810 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n7167) );
  NAND2_X1 U6811 ( .A1(n5652), .A2(n7167), .ZN(n5109) );
  NAND2_X1 U6812 ( .A1(n5441), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5108) );
  NAND2_X1 U6813 ( .A1(n4298), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n5117) );
  XNOR2_X1 U6814 ( .A(n5113), .B(n5112), .ZN(n6575) );
  NAND2_X1 U6815 ( .A1(n5399), .A2(n6575), .ZN(n5116) );
  NAND2_X1 U6816 ( .A1(n6555), .A2(n6626), .ZN(n5115) );
  AND3_X2 U6817 ( .A1(n5117), .A2(n5116), .A3(n5115), .ZN(n9902) );
  INV_X1 U6818 ( .A(n5628), .ZN(n5118) );
  NAND2_X1 U6819 ( .A1(n9915), .A2(n9902), .ZN(n7352) );
  NAND2_X1 U6820 ( .A1(n7432), .A2(n9090), .ZN(n5120) );
  INV_X1 U6821 ( .A(n9915), .ZN(n7273) );
  NAND2_X1 U6822 ( .A1(n7273), .A2(n9902), .ZN(n5119) );
  NAND2_X1 U6823 ( .A1(n5150), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5125) );
  NAND2_X1 U6824 ( .A1(n5441), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n5124) );
  INV_X1 U6825 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n5121) );
  XNOR2_X1 U6826 ( .A(n5121), .B(P1_REG3_REG_3__SCAN_IN), .ZN(n7440) );
  NAND2_X1 U6827 ( .A1(n5652), .A2(n7440), .ZN(n5123) );
  INV_X2 U6828 ( .A(n5523), .ZN(n8995) );
  NAND2_X1 U6829 ( .A1(n8995), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5122) );
  XNOR2_X1 U6830 ( .A(n5126), .B(n5127), .ZN(n5865) );
  INV_X1 U6831 ( .A(n5865), .ZN(n6577) );
  NAND2_X1 U6832 ( .A1(n4297), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n5133) );
  OAI21_X1 U6833 ( .B1(P1_IR_REG_2__SCAN_IN), .B2(P1_IR_REG_3__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5128) );
  NAND2_X1 U6834 ( .A1(n5129), .A2(n5128), .ZN(n5131) );
  INV_X1 U6835 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n5130) );
  XNOR2_X1 U6836 ( .A(n5131), .B(n5130), .ZN(n6630) );
  NAND2_X1 U6837 ( .A1(n6555), .A2(n6630), .ZN(n5132) );
  OAI211_X1 U6838 ( .C1(n6577), .C2(n5166), .A(n5133), .B(n5132), .ZN(n9912)
         );
  NAND2_X1 U6839 ( .A1(n9928), .A2(n9912), .ZN(n7354) );
  INV_X1 U6840 ( .A(n9928), .ZN(n9228) );
  NAND2_X1 U6841 ( .A1(n9228), .A2(n7442), .ZN(n7411) );
  NAND2_X1 U6842 ( .A1(n7354), .A2(n7411), .ZN(n9091) );
  NAND2_X1 U6843 ( .A1(n7437), .A2(n9091), .ZN(n5135) );
  NAND2_X1 U6844 ( .A1(n9928), .A2(n7442), .ZN(n5134) );
  INV_X1 U6845 ( .A(n7303), .ZN(n5191) );
  NAND2_X1 U6846 ( .A1(n8884), .A2(n8559), .ZN(n9019) );
  INV_X1 U6847 ( .A(n8884), .ZN(n9224) );
  NAND2_X1 U6848 ( .A1(n9224), .A2(n9953), .ZN(n9014) );
  NAND2_X1 U6849 ( .A1(n9019), .A2(n9014), .ZN(n9099) );
  INV_X1 U6850 ( .A(n5136), .ZN(n5154) );
  INV_X1 U6851 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n5137) );
  NAND2_X1 U6852 ( .A1(n5154), .A2(n5137), .ZN(n5138) );
  AND2_X1 U6853 ( .A1(n5170), .A2(n5138), .ZN(n8955) );
  NAND2_X1 U6854 ( .A1(n4467), .A2(n8955), .ZN(n5139) );
  NAND2_X1 U6855 ( .A1(n5149), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5142) );
  NAND2_X1 U6856 ( .A1(n5150), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n5141) );
  NAND2_X1 U6857 ( .A1(n5441), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n5140) );
  INV_X1 U6858 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6570) );
  XNOR2_X1 U6859 ( .A(n5144), .B(SI_6_), .ZN(n5180) );
  NAND2_X1 U6860 ( .A1(n5022), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5145) );
  MUX2_X1 U6861 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5145), .S(
        P1_IR_REG_6__SCAN_IN), .Z(n5146) );
  INV_X1 U6862 ( .A(n5146), .ZN(n5147) );
  NOR2_X1 U6863 ( .A1(n5147), .A2(n5378), .ZN(n6658) );
  NAND2_X1 U6864 ( .A1(n6555), .A2(n6658), .ZN(n5148) );
  NAND2_X1 U6865 ( .A1(n5149), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n5158) );
  NAND2_X1 U6866 ( .A1(n5150), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5157) );
  INV_X1 U6867 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n5152) );
  NAND2_X1 U6868 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n5151) );
  NAND2_X1 U6869 ( .A1(n5152), .A2(n5151), .ZN(n5153) );
  AND2_X1 U6870 ( .A1(n5154), .A2(n5153), .ZN(n7612) );
  NAND2_X1 U6871 ( .A1(n4467), .A2(n7612), .ZN(n5156) );
  NAND2_X1 U6872 ( .A1(n5441), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n5155) );
  INV_X1 U6873 ( .A(n5869), .ZN(n6563) );
  NAND2_X1 U6874 ( .A1(n5161), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5162) );
  MUX2_X1 U6875 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5162), .S(
        P1_IR_REG_5__SCAN_IN), .Z(n5163) );
  AND2_X1 U6876 ( .A1(n5163), .A2(n5022), .ZN(n6657) );
  NAND2_X1 U6877 ( .A1(n6555), .A2(n6657), .ZN(n5164) );
  NAND2_X1 U6878 ( .A1(n7607), .A2(n7599), .ZN(n7414) );
  INV_X1 U6879 ( .A(n7599), .ZN(n9927) );
  NAND2_X1 U6880 ( .A1(n9227), .A2(n7599), .ZN(n7416) );
  NAND3_X1 U6881 ( .A1(n9005), .A2(n9095), .A3(n7416), .ZN(n5168) );
  NAND2_X1 U6882 ( .A1(n9944), .A2(n7621), .ZN(n5167) );
  NAND2_X1 U6883 ( .A1(n8994), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n5176) );
  NAND2_X1 U6884 ( .A1(n8995), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5175) );
  NAND2_X1 U6885 ( .A1(n5170), .A2(n5169), .ZN(n5171) );
  AND2_X1 U6886 ( .A1(n5172), .A2(n5171), .ZN(n7653) );
  NAND2_X1 U6887 ( .A1(n4467), .A2(n7653), .ZN(n5174) );
  NAND2_X1 U6888 ( .A1(n5441), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n5173) );
  INV_X1 U6889 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6580) );
  OR2_X1 U6890 ( .A1(n5378), .A2(n9752), .ZN(n5178) );
  XNOR2_X1 U6891 ( .A(n5178), .B(n5177), .ZN(n6671) );
  OAI22_X1 U6892 ( .A1(n4492), .A2(n6580), .B1(n4491), .B2(n6671), .ZN(n5179)
         );
  INV_X1 U6893 ( .A(n5179), .ZN(n5188) );
  INV_X1 U6894 ( .A(n5180), .ZN(n5181) );
  NAND2_X1 U6895 ( .A1(n5182), .A2(n5181), .ZN(n5184) );
  NAND2_X1 U6896 ( .A1(n6579), .A2(n5399), .ZN(n5187) );
  NAND2_X1 U6897 ( .A1(n5188), .A2(n5187), .ZN(n7637) );
  NAND2_X1 U6898 ( .A1(n8953), .A2(n7637), .ZN(n9017) );
  NAND2_X1 U6899 ( .A1(n9225), .A2(n9942), .ZN(n9133) );
  NAND2_X1 U6900 ( .A1(n8953), .A2(n9942), .ZN(n5189) );
  NAND3_X1 U6901 ( .A1(n5191), .A2(n9099), .A3(n5190), .ZN(n5193) );
  INV_X1 U6902 ( .A(n9099), .ZN(n7336) );
  NAND2_X1 U6903 ( .A1(n9005), .A2(n7416), .ZN(n7304) );
  NOR2_X1 U6904 ( .A1(n7304), .A2(n7309), .ZN(n7343) );
  INV_X1 U6905 ( .A(n5195), .ZN(n5196) );
  NAND2_X1 U6906 ( .A1(n5267), .A2(n5239), .ZN(n5216) );
  INV_X1 U6907 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6598) );
  MUX2_X1 U6908 ( .A(n6598), .B(n6586), .S(n4286), .Z(n5198) );
  INV_X1 U6909 ( .A(SI_9_), .ZN(n5197) );
  NAND2_X1 U6910 ( .A1(n5198), .A2(n5197), .ZN(n5238) );
  INV_X1 U6911 ( .A(n5198), .ZN(n5199) );
  NAND2_X1 U6912 ( .A1(n5199), .A2(SI_9_), .ZN(n5241) );
  AND2_X1 U6913 ( .A1(n5238), .A2(n5241), .ZN(n5215) );
  NAND2_X1 U6914 ( .A1(n6585), .A2(n5584), .ZN(n5208) );
  NOR2_X1 U6915 ( .A1(n5204), .A2(n9752), .ZN(n5202) );
  MUX2_X1 U6916 ( .A(n9752), .B(n5202), .S(P1_IR_REG_9__SCAN_IN), .Z(n5203) );
  INV_X1 U6917 ( .A(n5203), .ZN(n5205) );
  NAND2_X1 U6918 ( .A1(n5204), .A2(n10217), .ZN(n5225) );
  NAND2_X1 U6919 ( .A1(n5205), .A2(n5225), .ZN(n6869) );
  OAI22_X1 U6920 ( .A1(n4492), .A2(n6586), .B1(n4491), .B2(n6869), .ZN(n5206)
         );
  INV_X1 U6921 ( .A(n5206), .ZN(n5207) );
  NAND2_X1 U6922 ( .A1(n5208), .A2(n5207), .ZN(n8566) );
  NAND2_X1 U6923 ( .A1(n8994), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n5214) );
  NAND2_X1 U6924 ( .A1(n5747), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n5213) );
  NAND2_X1 U6925 ( .A1(n5209), .A2(n10248), .ZN(n5210) );
  AND2_X1 U6926 ( .A1(n5231), .A2(n5210), .ZN(n8887) );
  NAND2_X1 U6927 ( .A1(n4467), .A2(n8887), .ZN(n5212) );
  NAND2_X1 U6928 ( .A1(n8995), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5211) );
  INV_X1 U6929 ( .A(n8806), .ZN(n9223) );
  NAND2_X1 U6930 ( .A1(n5216), .A2(n5215), .ZN(n5217) );
  NAND2_X1 U6931 ( .A1(n5217), .A2(n5238), .ZN(n5223) );
  INV_X1 U6932 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n5218) );
  MUX2_X1 U6933 ( .A(n5218), .B(n6594), .S(n6561), .Z(n5219) );
  NAND2_X1 U6934 ( .A1(n5219), .A2(n10204), .ZN(n5260) );
  INV_X1 U6935 ( .A(n5219), .ZN(n5220) );
  NAND2_X1 U6936 ( .A1(n5220), .A2(SI_10_), .ZN(n5221) );
  NAND2_X1 U6937 ( .A1(n5260), .A2(n5221), .ZN(n5243) );
  INV_X1 U6938 ( .A(n5243), .ZN(n5222) );
  XNOR2_X1 U6939 ( .A(n5223), .B(n5222), .ZN(n6587) );
  NAND2_X1 U6940 ( .A1(n6587), .A2(n5584), .ZN(n5229) );
  NAND2_X1 U6941 ( .A1(n5225), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5224) );
  MUX2_X1 U6942 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5224), .S(
        P1_IR_REG_10__SCAN_IN), .Z(n5226) );
  NAND2_X1 U6943 ( .A1(n5226), .A2(n5275), .ZN(n6922) );
  OAI22_X1 U6944 ( .A1(n4492), .A2(n6594), .B1(n4491), .B2(n6922), .ZN(n5227)
         );
  INV_X1 U6945 ( .A(n5227), .ZN(n5228) );
  NAND2_X1 U6946 ( .A1(n8994), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n5236) );
  NAND2_X1 U6947 ( .A1(n5747), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n5235) );
  NAND2_X1 U6948 ( .A1(n5231), .A2(n5230), .ZN(n5232) );
  AND2_X1 U6949 ( .A1(n5253), .A2(n5232), .ZN(n8759) );
  NAND2_X1 U6950 ( .A1(n4467), .A2(n8759), .ZN(n5234) );
  NAND2_X1 U6951 ( .A1(n8995), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5233) );
  OR2_X1 U6952 ( .A1(n8580), .A2(n8581), .ZN(n9011) );
  NAND2_X1 U6953 ( .A1(n8580), .A2(n8581), .ZN(n9025) );
  NAND2_X1 U6954 ( .A1(n9011), .A2(n9025), .ZN(n9101) );
  INV_X1 U6955 ( .A(n8581), .ZN(n9222) );
  OR2_X1 U6956 ( .A1(n8580), .A2(n9222), .ZN(n5237) );
  NAND2_X1 U6957 ( .A1(n5239), .A2(n5238), .ZN(n5264) );
  INV_X1 U6958 ( .A(n5264), .ZN(n5240) );
  NAND2_X1 U6959 ( .A1(n5267), .A2(n5240), .ZN(n5244) );
  INV_X1 U6960 ( .A(n5241), .ZN(n5242) );
  NAND2_X1 U6961 ( .A1(n5244), .A2(n5265), .ZN(n5245) );
  NAND2_X1 U6962 ( .A1(n5245), .A2(n5260), .ZN(n5246) );
  MUX2_X1 U6963 ( .A(n10144), .B(n6592), .S(n4286), .Z(n5268) );
  XNOR2_X1 U6964 ( .A(n5246), .B(n5261), .ZN(n6591) );
  NAND2_X1 U6965 ( .A1(n6591), .A2(n5584), .ZN(n5251) );
  NAND2_X1 U6966 ( .A1(n5275), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5248) );
  INV_X1 U6967 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n5247) );
  XNOR2_X1 U6968 ( .A(n5248), .B(n5247), .ZN(n7237) );
  OAI22_X1 U6969 ( .A1(n4492), .A2(n6592), .B1(n4491), .B2(n7237), .ZN(n5249)
         );
  INV_X1 U6970 ( .A(n5249), .ZN(n5250) );
  NAND2_X1 U6971 ( .A1(n8995), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5258) );
  NAND2_X1 U6972 ( .A1(n8994), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n5257) );
  INV_X1 U6973 ( .A(n5279), .ZN(n5281) );
  NAND2_X1 U6974 ( .A1(n5253), .A2(n5252), .ZN(n5254) );
  AND2_X1 U6975 ( .A1(n5281), .A2(n5254), .ZN(n8929) );
  NAND2_X1 U6976 ( .A1(n4467), .A2(n8929), .ZN(n5256) );
  NAND2_X1 U6977 ( .A1(n5747), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n5255) );
  NAND2_X1 U6978 ( .A1(n8920), .A2(n9689), .ZN(n5259) );
  INV_X1 U6979 ( .A(n9567), .ZN(n5288) );
  INV_X1 U6980 ( .A(n5260), .ZN(n5263) );
  INV_X1 U6981 ( .A(n5261), .ZN(n5262) );
  AOI211_X1 U6982 ( .C1(n5265), .C2(n5264), .A(n5263), .B(n5262), .ZN(n5266)
         );
  INV_X1 U6983 ( .A(n5268), .ZN(n5269) );
  NAND2_X1 U6984 ( .A1(n5269), .A2(SI_11_), .ZN(n5270) );
  MUX2_X1 U6985 ( .A(n6602), .B(n6590), .S(n4287), .Z(n5272) );
  INV_X1 U6986 ( .A(SI_12_), .ZN(n5271) );
  INV_X1 U6987 ( .A(n5272), .ZN(n5273) );
  NAND2_X1 U6988 ( .A1(n5273), .A2(SI_12_), .ZN(n5274) );
  NAND2_X1 U6989 ( .A1(n5290), .A2(n5274), .ZN(n5291) );
  NAND2_X1 U6990 ( .A1(n6589), .A2(n5584), .ZN(n5278) );
  OAI21_X1 U6991 ( .B1(n5275), .B2(P1_IR_REG_11__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5276) );
  XNOR2_X1 U6992 ( .A(n5276), .B(P1_IR_REG_12__SCAN_IN), .ZN(n7671) );
  AOI22_X1 U6993 ( .A1(n4298), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n6555), .B2(
        n7671), .ZN(n5277) );
  NAND2_X1 U6994 ( .A1(n8994), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n5286) );
  NAND2_X1 U6995 ( .A1(n8995), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5285) );
  NAND2_X1 U6996 ( .A1(n5279), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n5309) );
  INV_X1 U6997 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n5280) );
  NAND2_X1 U6998 ( .A1(n5281), .A2(n5280), .ZN(n5282) );
  AND2_X1 U6999 ( .A1(n5309), .A2(n5282), .ZN(n9573) );
  NAND2_X1 U7000 ( .A1(n4467), .A2(n9573), .ZN(n5284) );
  NAND2_X1 U7001 ( .A1(n5747), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n5283) );
  OR2_X1 U7002 ( .A1(n9690), .A2(n9684), .ZN(n5635) );
  NAND2_X1 U7003 ( .A1(n9690), .A2(n9684), .ZN(n9548) );
  INV_X1 U7004 ( .A(n9568), .ZN(n5287) );
  NAND2_X1 U7005 ( .A1(n5288), .A2(n5287), .ZN(n9565) );
  NAND2_X1 U7006 ( .A1(n9690), .A2(n9543), .ZN(n5289) );
  MUX2_X1 U7007 ( .A(n6678), .B(n6679), .S(n4286), .Z(n5294) );
  INV_X1 U7008 ( .A(SI_13_), .ZN(n5293) );
  NAND2_X1 U7009 ( .A1(n5294), .A2(n5293), .ZN(n5317) );
  INV_X1 U7010 ( .A(n5294), .ZN(n5295) );
  NAND2_X1 U7011 ( .A1(n5295), .A2(SI_13_), .ZN(n5296) );
  XNOR2_X1 U7012 ( .A(n5316), .B(n4974), .ZN(n6677) );
  NAND2_X1 U7013 ( .A1(n6677), .A2(n5584), .ZN(n5308) );
  INV_X1 U7014 ( .A(n5298), .ZN(n5299) );
  AND2_X1 U7015 ( .A1(n5378), .A2(n5299), .ZN(n5303) );
  NOR2_X1 U7016 ( .A1(n5303), .A2(n9752), .ZN(n5300) );
  MUX2_X1 U7017 ( .A(n9752), .B(n5300), .S(P1_IR_REG_13__SCAN_IN), .Z(n5301)
         );
  INV_X1 U7018 ( .A(n5301), .ZN(n5305) );
  INV_X1 U7019 ( .A(n5341), .ZN(n5304) );
  INV_X1 U7020 ( .A(n9820), .ZN(n7680) );
  OAI22_X1 U7021 ( .A1(n4492), .A2(n6679), .B1(n4491), .B2(n7680), .ZN(n5306)
         );
  INV_X1 U7022 ( .A(n5306), .ZN(n5307) );
  NAND2_X1 U7023 ( .A1(n8994), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n5314) );
  NAND2_X1 U7024 ( .A1(n8995), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n5313) );
  NAND2_X1 U7025 ( .A1(n5309), .A2(n8904), .ZN(n5310) );
  AND2_X1 U7026 ( .A1(n5324), .A2(n5310), .ZN(n9537) );
  NAND2_X1 U7027 ( .A1(n4467), .A2(n9537), .ZN(n5312) );
  NAND2_X1 U7028 ( .A1(n5747), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n5311) );
  OR2_X1 U7029 ( .A1(n9681), .A2(n9561), .ZN(n5315) );
  MUX2_X1 U7030 ( .A(n5318), .B(n6697), .S(n4287), .Z(n5332) );
  XNOR2_X1 U7031 ( .A(n5332), .B(SI_14_), .ZN(n5330) );
  XNOR2_X1 U7032 ( .A(n5331), .B(n5330), .ZN(n6693) );
  NAND2_X1 U7033 ( .A1(n6693), .A2(n5584), .ZN(n5322) );
  OR2_X1 U7034 ( .A1(n5341), .A2(n9752), .ZN(n5319) );
  XNOR2_X1 U7035 ( .A(n5319), .B(P1_IR_REG_14__SCAN_IN), .ZN(n7681) );
  OAI22_X1 U7036 ( .A1(n4492), .A2(n6697), .B1(n4491), .B2(n9263), .ZN(n5320)
         );
  INV_X1 U7037 ( .A(n5320), .ZN(n5321) );
  NAND2_X1 U7038 ( .A1(n8995), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5329) );
  NAND2_X1 U7039 ( .A1(n8994), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n5328) );
  INV_X1 U7040 ( .A(n5346), .ZN(n5348) );
  NAND2_X1 U7041 ( .A1(n5324), .A2(n5323), .ZN(n5325) );
  AND2_X1 U7042 ( .A1(n5348), .A2(n5325), .ZN(n8727) );
  NAND2_X1 U7043 ( .A1(n4467), .A2(n8727), .ZN(n5327) );
  NAND2_X1 U7044 ( .A1(n5747), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n5326) );
  NAND2_X1 U7045 ( .A1(n9678), .A2(n9519), .ZN(n9152) );
  NAND2_X1 U7046 ( .A1(n9036), .A2(n9152), .ZN(n9105) );
  INV_X1 U7047 ( .A(n9519), .ZN(n9553) );
  INV_X1 U7048 ( .A(n5332), .ZN(n5333) );
  NAND2_X1 U7049 ( .A1(n5333), .A2(SI_14_), .ZN(n5334) );
  MUX2_X1 U7050 ( .A(n10235), .B(n6863), .S(n4287), .Z(n5337) );
  INV_X1 U7051 ( .A(SI_15_), .ZN(n5336) );
  INV_X1 U7052 ( .A(n5337), .ZN(n5338) );
  NAND2_X1 U7053 ( .A1(n5338), .A2(SI_15_), .ZN(n5339) );
  NAND2_X1 U7054 ( .A1(n5354), .A2(n5339), .ZN(n5355) );
  XNOR2_X1 U7055 ( .A(n5356), .B(n5355), .ZN(n6862) );
  NAND2_X1 U7056 ( .A1(n6862), .A2(n5584), .ZN(n5345) );
  NAND2_X1 U7057 ( .A1(n5341), .A2(n5340), .ZN(n5362) );
  NAND2_X1 U7058 ( .A1(n5362), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5342) );
  XNOR2_X1 U7059 ( .A(n5342), .B(P1_IR_REG_15__SCAN_IN), .ZN(n9832) );
  OAI22_X1 U7060 ( .A1(n4492), .A2(n6863), .B1(n4491), .B2(n9264), .ZN(n5343)
         );
  INV_X1 U7061 ( .A(n5343), .ZN(n5344) );
  NAND2_X1 U7062 ( .A1(n8995), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n5353) );
  NAND2_X1 U7063 ( .A1(n8994), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n5352) );
  INV_X1 U7064 ( .A(n5366), .ZN(n5368) );
  INV_X1 U7065 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n5347) );
  NAND2_X1 U7066 ( .A1(n5348), .A2(n5347), .ZN(n5349) );
  AND2_X1 U7067 ( .A1(n5368), .A2(n5349), .ZN(n9524) );
  NAND2_X1 U7068 ( .A1(n4467), .A2(n9524), .ZN(n5351) );
  NAND2_X1 U7069 ( .A1(n5747), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n5350) );
  INV_X1 U7070 ( .A(n9502), .ZN(n9221) );
  OR2_X1 U7071 ( .A1(n9523), .A2(n9221), .ZN(n9494) );
  MUX2_X1 U7072 ( .A(n10216), .B(n5357), .S(n6561), .Z(n5359) );
  INV_X1 U7073 ( .A(SI_16_), .ZN(n5358) );
  INV_X1 U7074 ( .A(n5359), .ZN(n5360) );
  NAND2_X1 U7075 ( .A1(n5360), .A2(SI_16_), .ZN(n5361) );
  XNOR2_X1 U7076 ( .A(n5375), .B(n4975), .ZN(n6983) );
  NAND2_X1 U7077 ( .A1(n6983), .A2(n5584), .ZN(n5365) );
  OAI21_X1 U7078 ( .B1(n5362), .B2(P1_IR_REG_15__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5363) );
  XNOR2_X1 U7079 ( .A(n5363), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9844) );
  AOI22_X1 U7080 ( .A1(n4297), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n6555), .B2(
        n9844), .ZN(n5364) );
  INV_X2 U7081 ( .A(n5481), .ZN(n8994) );
  NAND2_X1 U7082 ( .A1(n8994), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n5373) );
  NAND2_X1 U7083 ( .A1(n5747), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n5372) );
  INV_X1 U7084 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n5367) );
  NAND2_X1 U7085 ( .A1(n5368), .A2(n5367), .ZN(n5369) );
  AND2_X1 U7086 ( .A1(n5386), .A2(n5369), .ZN(n9507) );
  NAND2_X1 U7087 ( .A1(n4467), .A2(n9507), .ZN(n5371) );
  INV_X1 U7088 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n10257) );
  OR2_X1 U7089 ( .A1(n5523), .A2(n10257), .ZN(n5370) );
  OR2_X1 U7090 ( .A1(n9506), .A2(n9517), .ZN(n9155) );
  NAND2_X1 U7091 ( .A1(n9506), .A2(n9517), .ZN(n9481) );
  AND2_X1 U7092 ( .A1(n9494), .A2(n9500), .ZN(n5374) );
  NAND2_X1 U7093 ( .A1(n9523), .A2(n9221), .ZN(n9495) );
  INV_X1 U7094 ( .A(n9517), .ZN(n9220) );
  MUX2_X1 U7095 ( .A(n7108), .B(n7109), .S(n6561), .Z(n5395) );
  XNOR2_X1 U7096 ( .A(n5395), .B(SI_17_), .ZN(n5394) );
  XNOR2_X1 U7097 ( .A(n5446), .B(n5394), .ZN(n7107) );
  NAND2_X1 U7098 ( .A1(n7107), .A2(n5584), .ZN(n5384) );
  NAND2_X1 U7099 ( .A1(n5378), .A2(n5377), .ZN(n5380) );
  NAND2_X1 U7100 ( .A1(n5380), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5379) );
  MUX2_X1 U7101 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5379), .S(
        P1_IR_REG_17__SCAN_IN), .Z(n5381) );
  OR2_X1 U7102 ( .A1(n5380), .A2(P1_IR_REG_17__SCAN_IN), .ZN(n5400) );
  OAI22_X1 U7103 ( .A1(n4492), .A2(n7109), .B1(n4491), .B2(n9858), .ZN(n5382)
         );
  INV_X1 U7104 ( .A(n5382), .ZN(n5383) );
  INV_X1 U7105 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n5385) );
  NAND2_X1 U7106 ( .A1(n5386), .A2(n5385), .ZN(n5387) );
  AND2_X1 U7107 ( .A1(n5406), .A2(n5387), .ZN(n9489) );
  NAND2_X1 U7108 ( .A1(n9489), .A2(n4467), .ZN(n5391) );
  NAND2_X1 U7109 ( .A1(n8994), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n5390) );
  NAND2_X1 U7110 ( .A1(n5747), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n5389) );
  NAND2_X1 U7111 ( .A1(n8995), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n5388) );
  INV_X1 U7112 ( .A(n9503), .ZN(n9219) );
  AND2_X1 U7113 ( .A1(n9664), .A2(n9219), .ZN(n5392) );
  OR2_X1 U7114 ( .A1(n9664), .A2(n9219), .ZN(n5393) );
  INV_X1 U7115 ( .A(n5394), .ZN(n5415) );
  INV_X1 U7116 ( .A(n5395), .ZN(n5396) );
  NAND2_X1 U7117 ( .A1(n5396), .A2(SI_17_), .ZN(n5423) );
  MUX2_X1 U7118 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n6561), .Z(n5411) );
  XNOR2_X1 U7119 ( .A(n5411), .B(SI_18_), .ZN(n5412) );
  NAND2_X1 U7120 ( .A1(n7213), .A2(n5742), .ZN(n5404) );
  INV_X1 U7121 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n7214) );
  NAND2_X1 U7122 ( .A1(n5400), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5401) );
  XNOR2_X1 U7123 ( .A(n5401), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9276) );
  INV_X1 U7124 ( .A(n9276), .ZN(n9279) );
  OAI22_X1 U7125 ( .A1(n4492), .A2(n7214), .B1(n4491), .B2(n9279), .ZN(n5402)
         );
  INV_X1 U7126 ( .A(n5402), .ZN(n5403) );
  INV_X1 U7127 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n5405) );
  INV_X1 U7128 ( .A(n5439), .ZN(n5456) );
  NAND2_X1 U7129 ( .A1(n5406), .A2(n5405), .ZN(n5407) );
  NAND2_X1 U7130 ( .A1(n5456), .A2(n5407), .ZN(n9467) );
  INV_X1 U7131 ( .A(n4467), .ZN(n5478) );
  OR2_X1 U7132 ( .A1(n9467), .A2(n5478), .ZN(n5410) );
  AOI22_X1 U7133 ( .A1(n8995), .A2(P1_REG0_REG_18__SCAN_IN), .B1(n8994), .B2(
        P1_REG1_REG_18__SCAN_IN), .ZN(n5409) );
  NAND2_X1 U7134 ( .A1(n5747), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n5408) );
  OR2_X1 U7135 ( .A1(n9657), .A2(n9485), .ZN(n9056) );
  NAND2_X1 U7136 ( .A1(n9657), .A2(n9485), .ZN(n9160) );
  NAND2_X1 U7137 ( .A1(n9056), .A2(n9160), .ZN(n9464) );
  INV_X1 U7138 ( .A(n9485), .ZN(n9455) );
  NAND2_X1 U7139 ( .A1(n9657), .A2(n9455), .ZN(n9427) );
  NAND2_X1 U7140 ( .A1(n5411), .A2(SI_18_), .ZN(n5422) );
  INV_X1 U7141 ( .A(n5422), .ZN(n5414) );
  INV_X1 U7142 ( .A(n5412), .ZN(n5413) );
  MUX2_X1 U7143 ( .A(n7212), .B(n7210), .S(n4287), .Z(n5418) );
  INV_X1 U7144 ( .A(SI_19_), .ZN(n5416) );
  NAND2_X1 U7145 ( .A1(n5418), .A2(n5416), .ZN(n5421) );
  INV_X1 U7146 ( .A(n5421), .ZN(n5428) );
  INV_X1 U7147 ( .A(n5418), .ZN(n5419) );
  NAND2_X1 U7148 ( .A1(n5419), .A2(SI_19_), .ZN(n5420) );
  NAND2_X1 U7149 ( .A1(n5421), .A2(n5420), .ZN(n5449) );
  INV_X1 U7150 ( .A(n5449), .ZN(n5426) );
  AND2_X1 U7151 ( .A1(n5423), .A2(n5422), .ZN(n5424) );
  AND2_X1 U7152 ( .A1(n5468), .A2(n5465), .ZN(n5433) );
  MUX2_X1 U7153 ( .A(n7290), .B(n7269), .S(n4287), .Z(n5430) );
  INV_X1 U7154 ( .A(SI_20_), .ZN(n5429) );
  INV_X1 U7155 ( .A(n5430), .ZN(n5431) );
  NAND2_X1 U7156 ( .A1(n5431), .A2(SI_20_), .ZN(n5432) );
  NAND2_X1 U7157 ( .A1(n7268), .A2(n5742), .ZN(n5435) );
  NAND2_X1 U7158 ( .A1(n4298), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n5434) );
  INV_X1 U7159 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n5437) );
  INV_X1 U7160 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n5436) );
  OAI21_X1 U7161 ( .B1(n5456), .B2(n5437), .A(n5436), .ZN(n5440) );
  AND2_X1 U7162 ( .A1(P1_REG3_REG_20__SCAN_IN), .A2(P1_REG3_REG_19__SCAN_IN), 
        .ZN(n5438) );
  INV_X1 U7163 ( .A(n5473), .ZN(n5475) );
  NAND2_X1 U7164 ( .A1(n5440), .A2(n5475), .ZN(n9432) );
  OR2_X1 U7165 ( .A1(n9432), .A2(n5478), .ZN(n5444) );
  AOI22_X1 U7166 ( .A1(n8994), .A2(P1_REG1_REG_20__SCAN_IN), .B1(n5441), .B2(
        P1_REG2_REG_20__SCAN_IN), .ZN(n5443) );
  NAND2_X1 U7167 ( .A1(n8995), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n5442) );
  NAND2_X1 U7168 ( .A1(n9731), .A2(n9638), .ZN(n5487) );
  INV_X1 U7169 ( .A(n5487), .ZN(n5464) );
  NAND2_X1 U7170 ( .A1(n5448), .A2(n5447), .ZN(n5450) );
  XNOR2_X1 U7171 ( .A(n5450), .B(n5449), .ZN(n7209) );
  NAND2_X1 U7172 ( .A1(n7209), .A2(n5742), .ZN(n5455) );
  OAI22_X1 U7173 ( .A1(n4492), .A2(n7210), .B1(n9418), .B2(n4491), .ZN(n5453)
         );
  INV_X1 U7174 ( .A(n5453), .ZN(n5454) );
  XNOR2_X1 U7175 ( .A(n5456), .B(P1_REG3_REG_19__SCAN_IN), .ZN(n9449) );
  NAND2_X1 U7176 ( .A1(n9449), .A2(n4467), .ZN(n5462) );
  INV_X1 U7177 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n5459) );
  NAND2_X1 U7178 ( .A1(n5747), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n5458) );
  NAND2_X1 U7179 ( .A1(n8995), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n5457) );
  OAI211_X1 U7180 ( .C1(n5481), .C2(n5459), .A(n5458), .B(n5457), .ZN(n5460)
         );
  INV_X1 U7181 ( .A(n5460), .ZN(n5461) );
  INV_X1 U7182 ( .A(n9466), .ZN(n9218) );
  NAND2_X1 U7183 ( .A1(n9651), .A2(n9218), .ZN(n9429) );
  AND2_X1 U7184 ( .A1(n9429), .A2(n4983), .ZN(n5463) );
  AND2_X1 U7185 ( .A1(n9427), .A2(n5486), .ZN(n9408) );
  NAND2_X1 U7186 ( .A1(n5470), .A2(n5469), .ZN(n5496) );
  MUX2_X1 U7187 ( .A(n7369), .B(n7288), .S(n4287), .Z(n5492) );
  XNOR2_X1 U7188 ( .A(n5492), .B(SI_21_), .ZN(n5491) );
  XNOR2_X1 U7189 ( .A(n5496), .B(n5491), .ZN(n7287) );
  NAND2_X1 U7190 ( .A1(n7287), .A2(n5742), .ZN(n5472) );
  NAND2_X1 U7191 ( .A1(n4297), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n5471) );
  INV_X1 U7192 ( .A(n5502), .ZN(n5477) );
  INV_X1 U7193 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n5474) );
  NAND2_X1 U7194 ( .A1(n5475), .A2(n5474), .ZN(n5476) );
  NAND2_X1 U7195 ( .A1(n5477), .A2(n5476), .ZN(n9416) );
  OR2_X1 U7196 ( .A1(n9416), .A2(n5478), .ZN(n5484) );
  INV_X1 U7197 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n10254) );
  NAND2_X1 U7198 ( .A1(n8995), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n5480) );
  NAND2_X1 U7199 ( .A1(n5747), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n5479) );
  OAI211_X1 U7200 ( .C1(n5481), .C2(n10254), .A(n5480), .B(n5479), .ZN(n5482)
         );
  INV_X1 U7201 ( .A(n5482), .ZN(n5483) );
  NAND2_X1 U7202 ( .A1(n9641), .A2(n9217), .ZN(n5485) );
  INV_X1 U7203 ( .A(n5485), .ZN(n5490) );
  NAND2_X1 U7204 ( .A1(n9641), .A2(n9633), .ZN(n9060) );
  INV_X1 U7205 ( .A(n5486), .ZN(n5489) );
  OR2_X1 U7206 ( .A1(n9651), .A2(n9218), .ZN(n9428) );
  AND2_X1 U7207 ( .A1(n9428), .A2(n5487), .ZN(n5488) );
  INV_X1 U7208 ( .A(n5491), .ZN(n5495) );
  INV_X1 U7209 ( .A(n5492), .ZN(n5493) );
  NAND2_X1 U7210 ( .A1(n5493), .A2(SI_21_), .ZN(n5494) );
  MUX2_X1 U7211 ( .A(n10187), .B(n7350), .S(n4287), .Z(n5497) );
  NAND2_X1 U7212 ( .A1(n5497), .A2(n10251), .ZN(n5508) );
  INV_X1 U7213 ( .A(n5497), .ZN(n5498) );
  NAND2_X1 U7214 ( .A1(n5498), .A2(SI_22_), .ZN(n5499) );
  NAND2_X1 U7215 ( .A1(n5508), .A2(n5499), .ZN(n5509) );
  XNOR2_X1 U7216 ( .A(n5510), .B(n5509), .ZN(n7349) );
  NAND2_X1 U7217 ( .A1(n7349), .A2(n5742), .ZN(n5501) );
  NAND2_X1 U7218 ( .A1(n4297), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n5500) );
  NOR2_X1 U7219 ( .A1(n5502), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n5503) );
  NOR2_X1 U7220 ( .A1(n5519), .A2(n5503), .ZN(n9398) );
  INV_X1 U7221 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n9723) );
  NAND2_X1 U7222 ( .A1(n5747), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n5505) );
  NAND2_X1 U7223 ( .A1(n8994), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n5504) );
  OAI211_X1 U7224 ( .C1(n5523), .C2(n9723), .A(n5505), .B(n5504), .ZN(n5506)
         );
  AOI21_X1 U7225 ( .B1(n9398), .B2(n4467), .A(n5506), .ZN(n9626) );
  INV_X1 U7226 ( .A(n9626), .ZN(n9421) );
  OR2_X1 U7227 ( .A1(n9405), .A2(n9421), .ZN(n5507) );
  NAND2_X1 U7228 ( .A1(n9405), .A2(n9421), .ZN(n9379) );
  INV_X1 U7229 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n5512) );
  INV_X1 U7230 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n5511) );
  MUX2_X1 U7231 ( .A(n5512), .B(n5511), .S(n4287), .Z(n5514) );
  INV_X1 U7232 ( .A(SI_23_), .ZN(n5513) );
  NAND2_X1 U7233 ( .A1(n5514), .A2(n5513), .ZN(n5530) );
  INV_X1 U7234 ( .A(n5514), .ZN(n5515) );
  NAND2_X1 U7235 ( .A1(n5515), .A2(SI_23_), .ZN(n5516) );
  XNOR2_X1 U7236 ( .A(n5529), .B(n5528), .ZN(n7506) );
  NAND2_X1 U7237 ( .A1(n7506), .A2(n5742), .ZN(n5518) );
  NAND2_X1 U7238 ( .A1(n4298), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n5517) );
  OR2_X1 U7239 ( .A1(n5519), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n5520) );
  AND2_X1 U7240 ( .A1(n5520), .A2(n5533), .ZN(n9383) );
  NAND2_X1 U7241 ( .A1(n9383), .A2(n4467), .ZN(n5526) );
  INV_X1 U7242 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n9720) );
  NAND2_X1 U7243 ( .A1(n5747), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n5522) );
  NAND2_X1 U7244 ( .A1(n8994), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n5521) );
  OAI211_X1 U7245 ( .C1(n5523), .C2(n9720), .A(n5522), .B(n5521), .ZN(n5524)
         );
  INV_X1 U7246 ( .A(n5524), .ZN(n5525) );
  NAND2_X1 U7247 ( .A1(n5526), .A2(n5525), .ZN(n9393) );
  NAND2_X1 U7248 ( .A1(n9388), .A2(n9393), .ZN(n5527) );
  MUX2_X1 U7249 ( .A(n7721), .B(n10232), .S(n4287), .Z(n5540) );
  XNOR2_X1 U7250 ( .A(n5540), .B(SI_24_), .ZN(n5538) );
  XNOR2_X1 U7251 ( .A(n5539), .B(n5538), .ZN(n7720) );
  NAND2_X1 U7252 ( .A1(n7720), .A2(n5742), .ZN(n5532) );
  NAND2_X1 U7253 ( .A1(n4298), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n5531) );
  NAND2_X1 U7254 ( .A1(n8994), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n5537) );
  NAND2_X1 U7255 ( .A1(n5747), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n5536) );
  INV_X1 U7256 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n10164) );
  AOI21_X1 U7257 ( .B1(n10164), .B2(n5533), .A(n5550), .ZN(n9370) );
  NAND2_X1 U7258 ( .A1(n4467), .A2(n9370), .ZN(n5535) );
  NAND2_X1 U7259 ( .A1(n8995), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n5534) );
  INV_X1 U7260 ( .A(n5540), .ZN(n5541) );
  NAND2_X1 U7261 ( .A1(n5541), .A2(SI_24_), .ZN(n5542) );
  MUX2_X1 U7262 ( .A(n10263), .B(n7783), .S(n4287), .Z(n5545) );
  INV_X1 U7263 ( .A(SI_25_), .ZN(n5544) );
  NAND2_X1 U7264 ( .A1(n5545), .A2(n5544), .ZN(n5558) );
  INV_X1 U7265 ( .A(n5545), .ZN(n5546) );
  NAND2_X1 U7266 ( .A1(n5546), .A2(SI_25_), .ZN(n5547) );
  NAND2_X1 U7267 ( .A1(n5558), .A2(n5547), .ZN(n5559) );
  NAND2_X1 U7268 ( .A1(n7781), .A2(n5584), .ZN(n5549) );
  NAND2_X1 U7269 ( .A1(n4297), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n5548) );
  NAND2_X1 U7270 ( .A1(n8994), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n5555) );
  NAND2_X1 U7271 ( .A1(n5747), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n5554) );
  NAND2_X1 U7272 ( .A1(n5550), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n5568) );
  OAI21_X1 U7273 ( .B1(n5550), .B2(P1_REG3_REG_25__SCAN_IN), .A(n5568), .ZN(
        n5551) );
  INV_X1 U7274 ( .A(n5551), .ZN(n9353) );
  NAND2_X1 U7275 ( .A1(n4467), .A2(n9353), .ZN(n5553) );
  NAND2_X1 U7276 ( .A1(n8995), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n5552) );
  NAND2_X1 U7277 ( .A1(n9352), .A2(n9609), .ZN(n9179) );
  NAND2_X1 U7278 ( .A1(n9176), .A2(n9179), .ZN(n9346) );
  OR2_X1 U7279 ( .A1(n9352), .A2(n9364), .ZN(n5556) );
  INV_X1 U7280 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n7817) );
  INV_X1 U7281 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n7815) );
  MUX2_X1 U7282 ( .A(n7817), .B(n7815), .S(n4287), .Z(n5562) );
  INV_X1 U7283 ( .A(SI_26_), .ZN(n5561) );
  NAND2_X1 U7284 ( .A1(n5562), .A2(n5561), .ZN(n5578) );
  INV_X1 U7285 ( .A(n5562), .ZN(n5563) );
  NAND2_X1 U7286 ( .A1(n5563), .A2(SI_26_), .ZN(n5564) );
  XNOR2_X1 U7287 ( .A(n5577), .B(n5576), .ZN(n7814) );
  NAND2_X1 U7288 ( .A1(n7814), .A2(n5742), .ZN(n5566) );
  NAND2_X1 U7289 ( .A1(n4298), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n5565) );
  NAND2_X1 U7290 ( .A1(n8995), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n5574) );
  NAND2_X1 U7291 ( .A1(n8994), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n5573) );
  INV_X1 U7292 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n5567) );
  NAND2_X1 U7293 ( .A1(n5567), .A2(n5568), .ZN(n5570) );
  INV_X1 U7294 ( .A(n5568), .ZN(n5569) );
  NAND2_X1 U7295 ( .A1(P1_REG3_REG_26__SCAN_IN), .A2(n5569), .ZN(n5589) );
  AND2_X1 U7296 ( .A1(n5570), .A2(n5589), .ZN(n9337) );
  NAND2_X1 U7297 ( .A1(n4467), .A2(n9337), .ZN(n5572) );
  NAND2_X1 U7298 ( .A1(n5747), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n5571) );
  NAND4_X1 U7299 ( .A1(n5574), .A2(n5573), .A3(n5572), .A4(n5571), .ZN(n9216)
         );
  NOR2_X1 U7300 ( .A1(n9342), .A2(n9216), .ZN(n5575) );
  INV_X1 U7301 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n7832) );
  INV_X1 U7302 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n5579) );
  MUX2_X1 U7303 ( .A(n7832), .B(n5579), .S(n4287), .Z(n5581) );
  INV_X1 U7304 ( .A(SI_27_), .ZN(n5580) );
  NAND2_X1 U7305 ( .A1(n5581), .A2(n5580), .ZN(n5597) );
  INV_X1 U7306 ( .A(n5581), .ZN(n5582) );
  NAND2_X1 U7307 ( .A1(n5582), .A2(SI_27_), .ZN(n5583) );
  XNOR2_X1 U7308 ( .A(n5596), .B(n5595), .ZN(n7820) );
  NAND2_X1 U7309 ( .A1(n7820), .A2(n5584), .ZN(n5586) );
  NAND2_X1 U7310 ( .A1(n4297), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n5585) );
  NAND2_X1 U7311 ( .A1(n8994), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n5594) );
  NAND2_X1 U7312 ( .A1(n8995), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n5593) );
  INV_X1 U7313 ( .A(n5589), .ZN(n5587) );
  NAND2_X1 U7314 ( .A1(n5587), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n5604) );
  INV_X1 U7315 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n5588) );
  NAND2_X1 U7316 ( .A1(n5589), .A2(n5588), .ZN(n5590) );
  NAND2_X1 U7317 ( .A1(n4467), .A2(n9320), .ZN(n5592) );
  NAND2_X1 U7318 ( .A1(n5747), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n5591) );
  AND4_X2 U7319 ( .A1(n5594), .A2(n5593), .A3(n5592), .A4(n5591), .ZN(n8964)
         );
  NAND2_X1 U7320 ( .A1(n9603), .A2(n8964), .ZN(n9126) );
  INV_X1 U7321 ( .A(n9323), .ZN(n9069) );
  NAND2_X1 U7322 ( .A1(n5598), .A2(n5597), .ZN(n5713) );
  INV_X1 U7323 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n7836) );
  INV_X1 U7324 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n5599) );
  MUX2_X1 U7325 ( .A(n7836), .B(n5599), .S(n4287), .Z(n5715) );
  XNOR2_X1 U7326 ( .A(n5715), .B(SI_28_), .ZN(n5712) );
  NAND2_X1 U7327 ( .A1(n7833), .A2(n5742), .ZN(n5601) );
  NAND2_X1 U7328 ( .A1(n4298), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n5600) );
  NAND2_X1 U7329 ( .A1(n8995), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n5609) );
  NAND2_X1 U7330 ( .A1(n8994), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n5608) );
  INV_X1 U7331 ( .A(n5604), .ZN(n5602) );
  NAND2_X1 U7332 ( .A1(n5602), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n9313) );
  INV_X1 U7333 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n5603) );
  NAND2_X1 U7334 ( .A1(n5604), .A2(n5603), .ZN(n5605) );
  NAND2_X1 U7335 ( .A1(n4467), .A2(n8792), .ZN(n5607) );
  NAND2_X1 U7336 ( .A1(n5747), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n5606) );
  AND4_X2 U7337 ( .A1(n5609), .A2(n5608), .A3(n5607), .A4(n5606), .ZN(n9591)
         );
  NAND2_X1 U7338 ( .A1(n9298), .A2(n9591), .ZN(n9307) );
  INV_X1 U7339 ( .A(n8964), .ZN(n9333) );
  NAND2_X1 U7340 ( .A1(n5620), .A2(n5619), .ZN(n5613) );
  NAND2_X1 U7341 ( .A1(n5618), .A2(n5617), .ZN(n5614) );
  INV_X1 U7342 ( .A(n9121), .ZN(n6709) );
  NAND2_X1 U7343 ( .A1(n9120), .A2(n9418), .ZN(n5697) );
  AOI21_X1 U7344 ( .B1(n8993), .B2(n6988), .A(n9119), .ZN(n5621) );
  NAND2_X1 U7345 ( .A1(n8991), .A2(n5621), .ZN(n9887) );
  NAND2_X1 U7346 ( .A1(n9120), .A2(n9119), .ZN(n5690) );
  INV_X1 U7347 ( .A(n5690), .ZN(n9869) );
  NAND2_X1 U7348 ( .A1(n8993), .A2(n9869), .ZN(n9894) );
  OAI21_X1 U7349 ( .B1(n5762), .B2(n5763), .A(n9966), .ZN(n5622) );
  INV_X1 U7350 ( .A(n5622), .ZN(n5624) );
  NAND3_X1 U7351 ( .A1(n9299), .A2(n5624), .A3(n5623), .ZN(n5667) );
  OAI21_X1 U7352 ( .B1(n7295), .B2(n9231), .A(n9889), .ZN(n5626) );
  NAND2_X1 U7353 ( .A1(n7295), .A2(n9231), .ZN(n5625) );
  NAND2_X1 U7354 ( .A1(n5626), .A2(n5625), .ZN(n7275) );
  AOI21_X1 U7355 ( .B1(n9012), .B2(n5630), .A(n9018), .ZN(n5631) );
  OR2_X1 U7356 ( .A1(n8806), .A2(n8566), .ZN(n9010) );
  AND2_X1 U7357 ( .A1(n9010), .A2(n9014), .ZN(n5633) );
  AND2_X1 U7358 ( .A1(n5633), .A2(n9011), .ZN(n9147) );
  NAND2_X1 U7359 ( .A1(n8806), .A2(n8566), .ZN(n7492) );
  NAND2_X1 U7360 ( .A1(n9025), .A2(n7492), .ZN(n9020) );
  NAND2_X1 U7361 ( .A1(n9020), .A2(n9011), .ZN(n9139) );
  AND2_X1 U7362 ( .A1(n8920), .A2(n9575), .ZN(n9033) );
  OR2_X1 U7363 ( .A1(n8920), .A2(n9575), .ZN(n9558) );
  AND2_X1 U7364 ( .A1(n5635), .A2(n9558), .ZN(n9547) );
  OR2_X1 U7365 ( .A1(n9681), .A2(n8830), .ZN(n9029) );
  NAND2_X1 U7366 ( .A1(n9681), .A2(n8830), .ZN(n9151) );
  AND2_X1 U7367 ( .A1(n9547), .A2(n9552), .ZN(n7865) );
  AND2_X1 U7368 ( .A1(n7865), .A2(n9036), .ZN(n5638) );
  INV_X1 U7369 ( .A(n9151), .ZN(n5636) );
  NOR2_X1 U7370 ( .A1(n9105), .A2(n5636), .ZN(n5637) );
  OR2_X1 U7371 ( .A1(n9104), .A2(n9548), .ZN(n7868) );
  NOR2_X1 U7372 ( .A1(n9523), .A2(n9502), .ZN(n9154) );
  INV_X1 U7373 ( .A(n9154), .ZN(n5639) );
  NAND2_X1 U7374 ( .A1(n9523), .A2(n9502), .ZN(n9153) );
  OR2_X1 U7375 ( .A1(n9664), .A2(n9503), .ZN(n9046) );
  NAND2_X1 U7376 ( .A1(n9664), .A2(n9503), .ZN(n9158) );
  NAND2_X1 U7377 ( .A1(n9046), .A2(n9158), .ZN(n9482) );
  INV_X1 U7378 ( .A(n9481), .ZN(n9042) );
  NOR2_X1 U7379 ( .A1(n9482), .A2(n9042), .ZN(n5640) );
  NAND2_X1 U7380 ( .A1(n9480), .A2(n5640), .ZN(n5641) );
  OR2_X1 U7381 ( .A1(n9651), .A2(n9466), .ZN(n9055) );
  NAND2_X1 U7382 ( .A1(n9651), .A2(n9466), .ZN(n9436) );
  NAND2_X1 U7383 ( .A1(n9435), .A2(n9638), .ZN(n9088) );
  AND2_X1 U7384 ( .A1(n9088), .A2(n9436), .ZN(n9058) );
  NAND2_X1 U7385 ( .A1(n9731), .A2(n9456), .ZN(n9089) );
  NAND2_X1 U7386 ( .A1(n9405), .A2(n9626), .ZN(n9087) );
  NAND2_X1 U7387 ( .A1(n9392), .A2(n9087), .ZN(n5643) );
  OR2_X1 U7388 ( .A1(n9405), .A2(n9626), .ZN(n9170) );
  AND2_X1 U7389 ( .A1(n9722), .A2(n9393), .ZN(n9172) );
  INV_X1 U7390 ( .A(n9393), .ZN(n8916) );
  NAND2_X1 U7391 ( .A1(n9388), .A2(n8916), .ZN(n9085) );
  NAND2_X1 U7392 ( .A1(n9369), .A2(n9350), .ZN(n9050) );
  NAND2_X1 U7393 ( .A1(n5644), .A2(n9179), .ZN(n9332) );
  XNOR2_X1 U7394 ( .A(n9342), .B(n9216), .ZN(n9336) );
  NAND2_X1 U7395 ( .A1(n9342), .A2(n9349), .ZN(n9127) );
  NAND2_X1 U7396 ( .A1(n9326), .A2(n9070), .ZN(n5645) );
  NAND2_X1 U7397 ( .A1(n5645), .A2(n5762), .ZN(n5647) );
  INV_X1 U7398 ( .A(n9070), .ZN(n9128) );
  NOR2_X1 U7399 ( .A1(n5762), .A2(n9128), .ZN(n5646) );
  NAND2_X1 U7400 ( .A1(n9326), .A2(n5646), .ZN(n9308) );
  NAND2_X1 U7401 ( .A1(n5647), .A2(n9308), .ZN(n5650) );
  NAND2_X1 U7402 ( .A1(n9118), .A2(n9119), .ZN(n5649) );
  INV_X1 U7403 ( .A(n9120), .ZN(n5663) );
  NAND2_X1 U7404 ( .A1(n4480), .A2(n5663), .ZN(n5648) );
  NAND2_X1 U7405 ( .A1(n5650), .A2(n9563), .ZN(n5658) );
  NAND2_X1 U7406 ( .A1(n8995), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n5656) );
  NAND2_X1 U7407 ( .A1(n8994), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n5655) );
  INV_X1 U7408 ( .A(n9313), .ZN(n5651) );
  NAND2_X1 U7409 ( .A1(n4467), .A2(n5651), .ZN(n5654) );
  NAND2_X1 U7410 ( .A1(n5747), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n5653) );
  OR2_X1 U7411 ( .A1(n9076), .A2(n9518), .ZN(n5657) );
  NAND2_X1 U7412 ( .A1(n5658), .A2(n5657), .ZN(n5770) );
  INV_X1 U7413 ( .A(n4300), .ZN(n8989) );
  INV_X1 U7414 ( .A(n7292), .ZN(n6715) );
  NAND2_X1 U7415 ( .A1(n7439), .A2(n7442), .ZN(n7438) );
  AND2_X1 U7416 ( .A1(n9953), .A2(n9962), .ZN(n5659) );
  INV_X1 U7417 ( .A(n9690), .ZN(n9571) );
  NOR2_X4 U7418 ( .A1(n4323), .A2(n9678), .ZN(n9520) );
  INV_X1 U7419 ( .A(n9651), .ZN(n9451) );
  AND2_X2 U7420 ( .A1(n9474), .A2(n9451), .ZN(n9447) );
  INV_X1 U7421 ( .A(n9641), .ZN(n5660) );
  AND2_X1 U7422 ( .A1(n9731), .A2(n5660), .ZN(n5661) );
  NAND2_X1 U7423 ( .A1(n9447), .A2(n5661), .ZN(n9400) );
  NOR2_X2 U7424 ( .A1(n9400), .A2(n9405), .ZN(n9401) );
  AND2_X2 U7425 ( .A1(n9401), .A2(n9722), .ZN(n9367) );
  NOR2_X4 U7426 ( .A1(n9339), .A2(n9603), .ZN(n9319) );
  NAND2_X1 U7427 ( .A1(n8993), .A2(n5662), .ZN(n6763) );
  OAI211_X1 U7428 ( .C1(n9319), .C2(n9590), .A(n9302), .B(n9569), .ZN(n5776)
         );
  OAI21_X1 U7429 ( .B1(n8964), .B2(n9943), .A(n5776), .ZN(n5664) );
  NAND3_X1 U7430 ( .A1(n5667), .A2(n5666), .A3(n5665), .ZN(n5707) );
  OR2_X1 U7431 ( .A1(n5669), .A2(n5668), .ZN(n5670) );
  NAND2_X1 U7432 ( .A1(n7784), .A2(P1_B_REG_SCAN_IN), .ZN(n5673) );
  NAND2_X1 U7433 ( .A1(n4319), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5672) );
  MUX2_X1 U7434 ( .A(P1_B_REG_SCAN_IN), .B(n5673), .S(n7724), .Z(n5677) );
  INV_X1 U7435 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n6560) );
  NAND2_X1 U7436 ( .A1(n9878), .A2(n6560), .ZN(n5679) );
  NAND2_X1 U7437 ( .A1(n4464), .A2(n7784), .ZN(n5678) );
  NAND2_X1 U7438 ( .A1(n5679), .A2(n5678), .ZN(n6557) );
  NOR4_X1 U7439 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        P1_D_REG_6__SCAN_IN), .A4(P1_D_REG_7__SCAN_IN), .ZN(n5688) );
  NOR4_X1 U7440 ( .A1(P1_D_REG_8__SCAN_IN), .A2(P1_D_REG_9__SCAN_IN), .A3(
        P1_D_REG_10__SCAN_IN), .A4(P1_D_REG_11__SCAN_IN), .ZN(n5687) );
  INV_X1 U7441 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n10173) );
  INV_X1 U7442 ( .A(P1_D_REG_21__SCAN_IN), .ZN(n10199) );
  INV_X1 U7443 ( .A(P1_D_REG_5__SCAN_IN), .ZN(n10227) );
  INV_X1 U7444 ( .A(P1_D_REG_15__SCAN_IN), .ZN(n10247) );
  NAND4_X1 U7445 ( .A1(n10173), .A2(n10199), .A3(n10227), .A4(n10247), .ZN(
        n5685) );
  NOR4_X1 U7446 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_18__SCAN_IN), .A3(
        P1_D_REG_19__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n5683) );
  NOR4_X1 U7447 ( .A1(P1_D_REG_14__SCAN_IN), .A2(P1_D_REG_12__SCAN_IN), .A3(
        P1_D_REG_13__SCAN_IN), .A4(P1_D_REG_16__SCAN_IN), .ZN(n5682) );
  NOR4_X1 U7448 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n5681) );
  NOR4_X1 U7449 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n5680) );
  NAND4_X1 U7450 ( .A1(n5683), .A2(n5682), .A3(n5681), .A4(n5680), .ZN(n5684)
         );
  NOR4_X1 U7451 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        n5685), .A4(n5684), .ZN(n5686) );
  NAND3_X1 U7452 ( .A1(n5688), .A2(n5687), .A3(n5686), .ZN(n5689) );
  NAND2_X1 U7453 ( .A1(n9878), .A2(n5689), .ZN(n5765) );
  NAND3_X1 U7454 ( .A1(n6557), .A2(n5765), .A3(n6700), .ZN(n5705) );
  NOR2_X1 U7455 ( .A1(n5705), .A2(n7159), .ZN(n5696) );
  INV_X1 U7456 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n9883) );
  NAND2_X1 U7457 ( .A1(n9878), .A2(n9883), .ZN(n5692) );
  NAND2_X1 U7458 ( .A1(n4464), .A2(n7724), .ZN(n5691) );
  OAI21_X1 U7459 ( .B1(n4396), .B2(n5693), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n5694) );
  AND2_X1 U7460 ( .A1(n8988), .A2(P1_STATE_REG_SCAN_IN), .ZN(n5695) );
  NAND2_X1 U7461 ( .A1(n6699), .A2(n9884), .ZN(n9882) );
  INV_X1 U7462 ( .A(n5697), .ZN(n9194) );
  OR2_X1 U7463 ( .A1(n6763), .A2(n9194), .ZN(n9961) );
  NAND2_X1 U7464 ( .A1(n9298), .A2(n5698), .ZN(n5701) );
  NAND2_X1 U7465 ( .A1(n5699), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n5700) );
  NOR2_X1 U7466 ( .A1(n6699), .A2(n7159), .ZN(n5704) );
  INV_X1 U7467 ( .A(n5705), .ZN(n5706) );
  NAND2_X1 U7468 ( .A1(n5707), .A2(n9970), .ZN(n5711) );
  INV_X1 U7469 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n5708) );
  NOR2_X1 U7470 ( .A1(n9970), .A2(n5708), .ZN(n5709) );
  NAND2_X1 U7471 ( .A1(n5711), .A2(n5710), .ZN(P1_U3519) );
  INV_X1 U7472 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n5754) );
  NAND2_X1 U7473 ( .A1(n5713), .A2(n5712), .ZN(n5718) );
  INV_X1 U7474 ( .A(SI_28_), .ZN(n5714) );
  NAND2_X1 U7475 ( .A1(n5715), .A2(n5714), .ZN(n5716) );
  INV_X1 U7476 ( .A(SI_29_), .ZN(n5734) );
  MUX2_X1 U7477 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .S(n4287), .Z(n5735) );
  AND2_X1 U7478 ( .A1(n5716), .A2(n5735), .ZN(n5717) );
  NAND2_X1 U7479 ( .A1(n5718), .A2(n5717), .ZN(n5721) );
  INV_X1 U7480 ( .A(n5735), .ZN(n5719) );
  OR2_X1 U7481 ( .A1(n5719), .A2(n5734), .ZN(n5720) );
  MUX2_X1 U7482 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n6562), .Z(n5739) );
  INV_X1 U7483 ( .A(n5739), .ZN(n5722) );
  NAND2_X1 U7484 ( .A1(n5726), .A2(n5723), .ZN(n5725) );
  OR2_X1 U7485 ( .A1(n5739), .A2(SI_30_), .ZN(n5724) );
  INV_X1 U7486 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n5728) );
  INV_X1 U7487 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n8546) );
  MUX2_X1 U7488 ( .A(n5728), .B(n8546), .S(n6562), .Z(n5729) );
  XNOR2_X1 U7489 ( .A(n5729), .B(SI_31_), .ZN(n5730) );
  NAND2_X1 U7490 ( .A1(n4297), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n5731) );
  XNOR2_X1 U7491 ( .A(n5735), .B(n5734), .ZN(n5736) );
  NAND2_X1 U7492 ( .A1(n8551), .A2(n5742), .ZN(n5738) );
  NAND2_X1 U7493 ( .A1(n4297), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n5737) );
  XNOR2_X1 U7494 ( .A(n5739), .B(SI_30_), .ZN(n5740) );
  NAND2_X1 U7495 ( .A1(n7894), .A2(n5742), .ZN(n5745) );
  NAND2_X1 U7496 ( .A1(n4298), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n5744) );
  NAND2_X1 U7497 ( .A1(n8994), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n5750) );
  NAND2_X1 U7498 ( .A1(n5747), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n5749) );
  NAND2_X1 U7499 ( .A1(n8995), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n5748) );
  NAND3_X1 U7500 ( .A1(n5750), .A2(n5749), .A3(n5748), .ZN(n9114) );
  INV_X1 U7501 ( .A(n6893), .ZN(n6890) );
  NAND2_X1 U7502 ( .A1(n6890), .A2(P1_B_REG_SCAN_IN), .ZN(n5752) );
  NAND2_X1 U7503 ( .A1(n9562), .A2(n5752), .ZN(n9310) );
  INV_X1 U7504 ( .A(n9310), .ZN(n5753) );
  NOR2_X1 U7505 ( .A1(n9289), .A2(n9584), .ZN(n5757) );
  NAND2_X1 U7506 ( .A1(n9115), .A2(n5698), .ZN(n5755) );
  NAND2_X1 U7507 ( .A1(n5756), .A2(n5755), .ZN(P1_U3554) );
  INV_X1 U7508 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n5758) );
  NAND2_X1 U7509 ( .A1(n9115), .A2(n5759), .ZN(n5760) );
  NAND2_X1 U7510 ( .A1(n5761), .A2(n5760), .ZN(P1_U3522) );
  INV_X1 U7511 ( .A(n5762), .ZN(n9113) );
  NAND2_X1 U7512 ( .A1(n5764), .A2(n5763), .ZN(n5769) );
  INV_X1 U7513 ( .A(n5765), .ZN(n5766) );
  NAND2_X1 U7514 ( .A1(n5767), .A2(n6707), .ZN(n5771) );
  INV_X1 U7515 ( .A(n6700), .ZN(n5768) );
  OR2_X1 U7516 ( .A1(n6988), .A2(n9418), .ZN(n7271) );
  NAND2_X1 U7517 ( .A1(n9887), .A2(n7271), .ZN(n7299) );
  AOI211_X1 U7518 ( .C1(n9113), .C2(n5769), .A(n9513), .B(n9589), .ZN(n5781)
         );
  NOR2_X1 U7519 ( .A1(n6763), .A2(n9120), .ZN(n5772) );
  AND2_X1 U7520 ( .A1(n9541), .A2(n9914), .ZN(n9544) );
  AOI22_X1 U7521 ( .A1(n9877), .A2(P1_REG2_REG_28__SCAN_IN), .B1(n8792), .B2(
        n9874), .ZN(n5773) );
  OAI21_X1 U7522 ( .B1(n9576), .B2(n8964), .A(n5773), .ZN(n5774) );
  AOI21_X1 U7523 ( .B1(n9298), .B2(n9578), .A(n5774), .ZN(n5775) );
  OAI21_X1 U7524 ( .B1(n5776), .B2(n9580), .A(n5775), .ZN(n5777) );
  NOR2_X2 U7525 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n5784) );
  NOR2_X2 U7526 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_13__SCAN_IN), .ZN(
        n5782) );
  NOR2_X2 U7527 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n5786) );
  NOR2_X1 U7528 ( .A1(P2_IR_REG_23__SCAN_IN), .A2(P2_IR_REG_22__SCAN_IN), .ZN(
        n5791) );
  NOR2_X1 U7529 ( .A1(P2_IR_REG_24__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), .ZN(
        n5790) );
  NOR2_X1 U7530 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n5789) );
  NOR2_X1 U7531 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), .ZN(
        n5788) );
  NAND3_X1 U7532 ( .A1(n6014), .A2(n10218), .A3(n6359), .ZN(n5792) );
  NAND2_X1 U7533 ( .A1(n5795), .A2(n5794), .ZN(n5796) );
  XNOR2_X2 U7534 ( .A(n5797), .B(n8545), .ZN(n5803) );
  NAND2_X1 U7535 ( .A1(n5815), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5798) );
  NAND2_X1 U7536 ( .A1(n5856), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n5809) );
  INV_X1 U7537 ( .A(n4288), .ZN(n5802) );
  NAND2_X1 U7538 ( .A1(n5802), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5808) );
  INV_X1 U7539 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n7511) );
  OR2_X1 U7540 ( .A1(n5857), .A2(n7511), .ZN(n5807) );
  INV_X1 U7541 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n7518) );
  AND4_X2 U7542 ( .A1(n5808), .A2(n5809), .A3(n5807), .A4(n5806), .ZN(n6958)
         );
  NAND2_X1 U7543 ( .A1(n6361), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5810) );
  MUX2_X2 U7544 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5810), .S(
        P2_IR_REG_27__SCAN_IN), .Z(n5812) );
  OR2_X2 U7545 ( .A1(n6361), .A2(P2_IR_REG_27__SCAN_IN), .ZN(n5811) );
  NAND2_X1 U7546 ( .A1(P2_IR_REG_27__SCAN_IN), .A2(P2_IR_REG_28__SCAN_IN), 
        .ZN(n5813) );
  AND2_X1 U7547 ( .A1(n6011), .A2(P2_IR_REG_28__SCAN_IN), .ZN(n5817) );
  AND2_X1 U7548 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_28__SCAN_IN), .ZN(
        n5814) );
  NAND2_X1 U7549 ( .A1(n6361), .A2(n5814), .ZN(n5816) );
  OAI211_X2 U7550 ( .C1(n5818), .C2(n5817), .A(n5816), .B(n5815), .ZN(n6371)
         );
  NAND2_X1 U7551 ( .A1(n4276), .A2(n6562), .ZN(n5848) );
  OR2_X1 U7552 ( .A1(n5848), .A2(n6573), .ZN(n5822) );
  NAND2_X1 U7553 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5819) );
  XNOR2_X1 U7554 ( .A(n5819), .B(P2_IR_REG_1__SCAN_IN), .ZN(n8069) );
  NAND2_X1 U7555 ( .A1(n5870), .A2(n8069), .ZN(n5820) );
  NAND2_X1 U7556 ( .A1(n5856), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5826) );
  INV_X1 U7557 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n7534) );
  OR2_X1 U7558 ( .A1(n5857), .A2(n7534), .ZN(n5825) );
  INV_X1 U7559 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n5823) );
  NAND2_X1 U7560 ( .A1(n6562), .A2(SI_0_), .ZN(n5828) );
  INV_X1 U7561 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5827) );
  NAND2_X1 U7562 ( .A1(n5828), .A2(n5827), .ZN(n5830) );
  AND2_X1 U7563 ( .A1(n5830), .A2(n5829), .ZN(n8554) );
  MUX2_X1 U7564 ( .A(P2_IR_REG_0__SCAN_IN), .B(n8554), .S(n6724), .Z(n7861) );
  NAND2_X1 U7565 ( .A1(n5856), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5834) );
  INV_X1 U7566 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n6729) );
  INV_X1 U7567 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n6781) );
  INV_X1 U7568 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n6741) );
  OR2_X1 U7569 ( .A1(n5858), .A2(n6741), .ZN(n5831) );
  INV_X1 U7570 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n6011) );
  OR2_X1 U7571 ( .A1(n5836), .A2(n6011), .ZN(n5837) );
  XNOR2_X1 U7572 ( .A(n5837), .B(P2_IR_REG_2__SCAN_IN), .ZN(n6788) );
  NAND2_X1 U7573 ( .A1(n5870), .A2(n6788), .ZN(n5838) );
  INV_X1 U7574 ( .A(n7021), .ZN(n7570) );
  NAND2_X1 U7575 ( .A1(n7571), .A2(n7570), .ZN(n5843) );
  NAND2_X1 U7576 ( .A1(n5843), .A2(n6247), .ZN(n6250) );
  NAND2_X1 U7577 ( .A1(n5856), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5847) );
  INV_X1 U7578 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n6730) );
  OR2_X1 U7579 ( .A1(n4289), .A2(n6730), .ZN(n5846) );
  OR2_X1 U7580 ( .A1(n5857), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n5844) );
  NAND2_X1 U7581 ( .A1(n5898), .A2(n6575), .ZN(n5855) );
  NOR2_X1 U7582 ( .A1(n5851), .A2(n6011), .ZN(n5849) );
  MUX2_X1 U7583 ( .A(n6011), .B(n5849), .S(P2_IR_REG_3__SCAN_IN), .Z(n5852) );
  NAND2_X1 U7584 ( .A1(n5870), .A2(n8082), .ZN(n5853) );
  OR2_X1 U7585 ( .A1(n8068), .A2(n10056), .ZN(n6240) );
  NAND2_X1 U7586 ( .A1(n8068), .A2(n10056), .ZN(n6235) );
  NAND2_X1 U7587 ( .A1(n6240), .A2(n6235), .ZN(n7024) );
  INV_X1 U7588 ( .A(n7024), .ZN(n10013) );
  NAND2_X1 U7589 ( .A1(n4280), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n5862) );
  NAND2_X1 U7590 ( .A1(n6174), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5861) );
  OAI21_X1 U7591 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(P2_REG3_REG_4__SCAN_IN), 
        .A(n5880), .ZN(n7586) );
  OR2_X1 U7592 ( .A1(n6076), .A2(n7586), .ZN(n5860) );
  INV_X1 U7593 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n6746) );
  OR2_X1 U7594 ( .A1(n5892), .A2(n6746), .ZN(n5859) );
  NAND2_X1 U7595 ( .A1(n5871), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5864) );
  XNOR2_X1 U7596 ( .A(n5864), .B(P2_IR_REG_4__SCAN_IN), .ZN(n6819) );
  AOI22_X1 U7597 ( .A1(n6139), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n4292), .B2(
        n6819), .ZN(n5867) );
  NAND2_X1 U7598 ( .A1(n5865), .A2(n5898), .ZN(n5866) );
  NAND2_X1 U7599 ( .A1(n5869), .A2(n5898), .ZN(n5878) );
  NAND2_X1 U7600 ( .A1(n5873), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5872) );
  MUX2_X1 U7601 ( .A(n5872), .B(P2_IR_REG_31__SCAN_IN), .S(n5874), .Z(n5876)
         );
  NAND2_X1 U7602 ( .A1(n5876), .A2(n5899), .ZN(n6780) );
  INV_X1 U7603 ( .A(n6780), .ZN(n6751) );
  AOI22_X1 U7604 ( .A1(n6139), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n4293), .B2(
        n6751), .ZN(n5877) );
  INV_X1 U7605 ( .A(n4284), .ZN(n7058) );
  INV_X1 U7606 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n6733) );
  OR2_X1 U7607 ( .A1(n4289), .A2(n6733), .ZN(n5883) );
  INV_X1 U7608 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n7527) );
  INV_X1 U7609 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5879) );
  NAND2_X1 U7610 ( .A1(n5880), .A2(n5879), .ZN(n5881) );
  NAND2_X1 U7611 ( .A1(n5890), .A2(n5881), .ZN(n7522) );
  OR2_X1 U7612 ( .A1(n6076), .A2(n7522), .ZN(n5882) );
  NAND2_X1 U7613 ( .A1(n7058), .A2(n8066), .ZN(n6233) );
  NAND2_X1 U7614 ( .A1(n8067), .A2(n7027), .ZN(n7030) );
  AND2_X1 U7615 ( .A1(n6233), .A2(n7030), .ZN(n6236) );
  NAND2_X1 U7616 ( .A1(n7029), .A2(n6236), .ZN(n5884) );
  NAND2_X1 U7617 ( .A1(n6565), .A2(n6182), .ZN(n5887) );
  NAND2_X1 U7618 ( .A1(n5899), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5885) );
  XNOR2_X1 U7619 ( .A(n5885), .B(P2_IR_REG_6__SCAN_IN), .ZN(n6803) );
  AOI22_X1 U7620 ( .A1(n6139), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n4292), .B2(
        n6803), .ZN(n5886) );
  NAND2_X2 U7621 ( .A1(n5887), .A2(n5886), .ZN(n7454) );
  NAND2_X1 U7622 ( .A1(n4280), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5896) );
  INV_X1 U7623 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n6734) );
  OR2_X1 U7624 ( .A1(n4289), .A2(n6734), .ZN(n5895) );
  INV_X1 U7625 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n5889) );
  NAND2_X1 U7626 ( .A1(n5890), .A2(n5889), .ZN(n5891) );
  NAND2_X1 U7627 ( .A1(n5903), .A2(n5891), .ZN(n7196) );
  OR2_X1 U7628 ( .A1(n6076), .A2(n7196), .ZN(n5894) );
  INV_X1 U7629 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n6752) );
  OR2_X1 U7630 ( .A1(n5892), .A2(n6752), .ZN(n5893) );
  OR2_X1 U7631 ( .A1(n7454), .A2(n7059), .ZN(n6262) );
  NAND2_X1 U7632 ( .A1(n7454), .A2(n7059), .ZN(n6266) );
  NAND2_X1 U7633 ( .A1(n7447), .A2(n7451), .ZN(n5897) );
  NAND2_X1 U7634 ( .A1(n5897), .A2(n6266), .ZN(n7175) );
  NAND2_X1 U7635 ( .A1(n6579), .A2(n6182), .ZN(n5902) );
  NAND2_X1 U7636 ( .A1(n5910), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5900) );
  XNOR2_X1 U7637 ( .A(n5900), .B(P2_IR_REG_7__SCAN_IN), .ZN(n6835) );
  AOI22_X1 U7638 ( .A1(n6139), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n6835), .B2(
        n4292), .ZN(n5901) );
  NAND2_X1 U7639 ( .A1(n5902), .A2(n5901), .ZN(n7216) );
  NAND2_X1 U7640 ( .A1(n4280), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5908) );
  INV_X1 U7641 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n6827) );
  OR2_X1 U7642 ( .A1(n4289), .A2(n6827), .ZN(n5907) );
  NAND2_X1 U7643 ( .A1(n5903), .A2(n6723), .ZN(n5904) );
  NAND2_X1 U7644 ( .A1(n5913), .A2(n5904), .ZN(n7475) );
  OR2_X1 U7645 ( .A1(n6076), .A2(n7475), .ZN(n5906) );
  INV_X1 U7646 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n6755) );
  OR2_X1 U7647 ( .A1(n5892), .A2(n6755), .ZN(n5905) );
  NAND2_X1 U7648 ( .A1(n7175), .A2(n6268), .ZN(n5909) );
  NAND2_X1 U7649 ( .A1(n7216), .A2(n7135), .ZN(n6267) );
  NAND2_X1 U7650 ( .A1(n5909), .A2(n6267), .ZN(n7225) );
  NAND2_X1 U7651 ( .A1(n5919), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5911) );
  XNOR2_X1 U7652 ( .A(n5911), .B(P2_IR_REG_8__SCAN_IN), .ZN(n6853) );
  AOI22_X1 U7653 ( .A1(n6853), .A2(n4293), .B1(n6139), .B2(
        P1_DATAO_REG_8__SCAN_IN), .ZN(n5912) );
  NAND2_X1 U7654 ( .A1(n4280), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n5918) );
  INV_X1 U7655 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n6829) );
  OR2_X1 U7656 ( .A1(n4289), .A2(n6829), .ZN(n5917) );
  INV_X1 U7657 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7379) );
  OR2_X1 U7658 ( .A1(n5892), .A2(n7379), .ZN(n5916) );
  NAND2_X1 U7659 ( .A1(n5913), .A2(n6845), .ZN(n5914) );
  NAND2_X1 U7660 ( .A1(n5925), .A2(n5914), .ZN(n7382) );
  OR2_X1 U7661 ( .A1(n6076), .A2(n7382), .ZN(n5915) );
  NAND4_X1 U7662 ( .A1(n5918), .A2(n5917), .A3(n5916), .A4(n5915), .ZN(n8063)
         );
  INV_X1 U7663 ( .A(n8063), .ZN(n7882) );
  NAND2_X1 U7664 ( .A1(n7389), .A2(n7882), .ZN(n6272) );
  NAND2_X1 U7665 ( .A1(n6585), .A2(n6182), .ZN(n5922) );
  NAND2_X1 U7666 ( .A1(n5931), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5920) );
  XNOR2_X1 U7667 ( .A(n5920), .B(P2_IR_REG_9__SCAN_IN), .ZN(n6932) );
  AOI22_X1 U7668 ( .A1(n6932), .A2(n4292), .B1(n6139), .B2(
        P1_DATAO_REG_9__SCAN_IN), .ZN(n5921) );
  NAND2_X1 U7669 ( .A1(n4280), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5930) );
  INV_X1 U7670 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n5923) );
  OR2_X1 U7671 ( .A1(n4289), .A2(n5923), .ZN(n5929) );
  NAND2_X1 U7672 ( .A1(n5925), .A2(n5924), .ZN(n5926) );
  NAND2_X1 U7673 ( .A1(n5938), .A2(n5926), .ZN(n7880) );
  OR2_X1 U7674 ( .A1(n6076), .A2(n7880), .ZN(n5928) );
  INV_X1 U7675 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n7394) );
  OR2_X1 U7676 ( .A1(n5892), .A2(n7394), .ZN(n5927) );
  OR2_X2 U7677 ( .A1(n7885), .A2(n7565), .ZN(n6278) );
  NAND2_X1 U7678 ( .A1(n7885), .A2(n7565), .ZN(n7545) );
  NAND2_X1 U7679 ( .A1(n6587), .A2(n6182), .ZN(n5936) );
  NAND2_X1 U7680 ( .A1(n5955), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5933) );
  INV_X1 U7681 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5932) );
  NAND2_X1 U7682 ( .A1(n5933), .A2(n5932), .ZN(n5944) );
  OR2_X1 U7683 ( .A1(n5933), .A2(n5932), .ZN(n5934) );
  AOI22_X1 U7684 ( .A1(n8108), .A2(n4293), .B1(n6139), .B2(
        P1_DATAO_REG_10__SCAN_IN), .ZN(n5935) );
  NAND2_X1 U7685 ( .A1(n4280), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5943) );
  INV_X1 U7686 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n6940) );
  OR2_X1 U7687 ( .A1(n4289), .A2(n6940), .ZN(n5942) );
  NAND2_X1 U7688 ( .A1(n5938), .A2(n4581), .ZN(n5939) );
  NAND2_X1 U7689 ( .A1(n5949), .A2(n5939), .ZN(n7564) );
  OR2_X1 U7690 ( .A1(n6076), .A2(n7564), .ZN(n5941) );
  INV_X1 U7691 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7550) );
  OR2_X1 U7692 ( .A1(n5892), .A2(n7550), .ZN(n5940) );
  NAND2_X1 U7693 ( .A1(n7704), .A2(n7881), .ZN(n7707) );
  NAND2_X1 U7694 ( .A1(n6591), .A2(n6182), .ZN(n5947) );
  NAND2_X1 U7695 ( .A1(n5944), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5945) );
  XNOR2_X1 U7696 ( .A(n5945), .B(P2_IR_REG_11__SCAN_IN), .ZN(n6968) );
  AOI22_X1 U7697 ( .A1(n6968), .A2(n4293), .B1(n6139), .B2(
        P1_DATAO_REG_11__SCAN_IN), .ZN(n5946) );
  NAND2_X1 U7698 ( .A1(n4280), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5954) );
  INV_X1 U7699 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n5948) );
  OR2_X1 U7700 ( .A1(n4289), .A2(n5948), .ZN(n5953) );
  NAND2_X1 U7701 ( .A1(n5949), .A2(n7406), .ZN(n5950) );
  NAND2_X1 U7702 ( .A1(n5961), .A2(n5950), .ZN(n7715) );
  OR2_X1 U7703 ( .A1(n6076), .A2(n7715), .ZN(n5952) );
  INV_X1 U7704 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n7711) );
  OR2_X1 U7705 ( .A1(n5892), .A2(n7711), .ZN(n5951) );
  NAND2_X1 U7706 ( .A1(n7737), .A2(n7846), .ZN(n6284) );
  NAND2_X1 U7707 ( .A1(n7707), .A2(n6284), .ZN(n7838) );
  OR2_X1 U7708 ( .A1(n7704), .A2(n7881), .ZN(n6271) );
  NAND2_X1 U7709 ( .A1(n6589), .A2(n6182), .ZN(n5958) );
  NAND2_X1 U7710 ( .A1(n5971), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5956) );
  XNOR2_X1 U7711 ( .A(n5956), .B(P2_IR_REG_12__SCAN_IN), .ZN(n7101) );
  AOI22_X1 U7712 ( .A1(n7101), .A2(n4292), .B1(n6139), .B2(
        P1_DATAO_REG_12__SCAN_IN), .ZN(n5957) );
  NAND2_X1 U7713 ( .A1(n6174), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n5966) );
  INV_X1 U7714 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n5959) );
  OR2_X1 U7715 ( .A1(n6179), .A2(n5959), .ZN(n5965) );
  INV_X1 U7716 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n5960) );
  NAND2_X1 U7717 ( .A1(n5961), .A2(n5960), .ZN(n5962) );
  NAND2_X1 U7718 ( .A1(n5974), .A2(n5962), .ZN(n7853) );
  OR2_X1 U7719 ( .A1(n6076), .A2(n7853), .ZN(n5964) );
  INV_X1 U7720 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n7849) );
  OR2_X1 U7721 ( .A1(n5892), .A2(n7849), .ZN(n5963) );
  OAI21_X1 U7722 ( .B1(n6271), .B2(n7846), .A(n6286), .ZN(n5968) );
  AOI21_X1 U7723 ( .B1(n6271), .B2(n7846), .A(n7737), .ZN(n5967) );
  NOR2_X1 U7724 ( .A1(n5968), .A2(n5967), .ZN(n5969) );
  NAND2_X1 U7725 ( .A1(n8519), .A2(n7735), .ZN(n6285) );
  NAND2_X1 U7726 ( .A1(n6677), .A2(n6182), .ZN(n5973) );
  INV_X1 U7727 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5982) );
  XNOR2_X1 U7728 ( .A(n5983), .B(P2_IR_REG_13__SCAN_IN), .ZN(n7116) );
  AOI22_X1 U7729 ( .A1(n7116), .A2(n4293), .B1(n6139), .B2(
        P1_DATAO_REG_13__SCAN_IN), .ZN(n5972) );
  NAND2_X1 U7730 ( .A1(n5974), .A2(n7996), .ZN(n5975) );
  AND2_X1 U7731 ( .A1(n5991), .A2(n5975), .ZN(n7995) );
  NAND2_X1 U7732 ( .A1(n6138), .A2(n7995), .ZN(n5981) );
  INV_X1 U7733 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n5976) );
  OR2_X1 U7734 ( .A1(n4289), .A2(n5976), .ZN(n5980) );
  INV_X1 U7735 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n6964) );
  OR2_X1 U7736 ( .A1(n5892), .A2(n6964), .ZN(n5979) );
  INV_X1 U7737 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n5977) );
  OR2_X1 U7738 ( .A1(n6179), .A2(n5977), .ZN(n5978) );
  OR2_X1 U7739 ( .A1(n8511), .A2(n7845), .ZN(n6291) );
  NAND2_X1 U7740 ( .A1(n8511), .A2(n7845), .ZN(n7770) );
  NAND2_X1 U7741 ( .A1(n6693), .A2(n6182), .ZN(n5986) );
  NAND2_X1 U7742 ( .A1(n5983), .A2(n5982), .ZN(n5984) );
  NAND2_X1 U7743 ( .A1(n5984), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5997) );
  AOI22_X1 U7744 ( .A1(n7323), .A2(n4292), .B1(n6139), .B2(
        P1_DATAO_REG_14__SCAN_IN), .ZN(n5985) );
  INV_X1 U7745 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n10233) );
  OR2_X1 U7746 ( .A1(n6179), .A2(n10233), .ZN(n5988) );
  INV_X1 U7747 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n7111) );
  OR2_X1 U7748 ( .A1(n4289), .A2(n7111), .ZN(n5987) );
  AND2_X1 U7749 ( .A1(n5988), .A2(n5987), .ZN(n5995) );
  INV_X1 U7750 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n5990) );
  NAND2_X1 U7751 ( .A1(n5991), .A2(n5990), .ZN(n5992) );
  NAND2_X1 U7752 ( .A1(n6004), .A2(n5992), .ZN(n7810) );
  OR2_X1 U7753 ( .A1(n7810), .A2(n6076), .ZN(n5994) );
  NAND2_X1 U7754 ( .A1(n6175), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n5993) );
  NAND2_X1 U7755 ( .A1(n8506), .A2(n7734), .ZN(n6295) );
  NAND2_X1 U7756 ( .A1(n6862), .A2(n6182), .ZN(n6003) );
  INV_X1 U7757 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5996) );
  NAND2_X1 U7758 ( .A1(n5997), .A2(n5996), .ZN(n5998) );
  NAND2_X1 U7759 ( .A1(n5998), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5999) );
  XNOR2_X1 U7760 ( .A(n5999), .B(P2_IR_REG_15__SCAN_IN), .ZN(n7322) );
  NOR2_X1 U7761 ( .A1(n4417), .A2(n10235), .ZN(n6001) );
  AOI21_X1 U7762 ( .B1(n7322), .B2(n4293), .A(n6001), .ZN(n6002) );
  NAND2_X1 U7763 ( .A1(n6004), .A2(n8035), .ZN(n6005) );
  AND2_X1 U7764 ( .A1(n6019), .A2(n6005), .ZN(n8034) );
  NAND2_X1 U7765 ( .A1(n8034), .A2(n6138), .ZN(n6008) );
  AOI22_X1 U7766 ( .A1(n4280), .A2(P2_REG0_REG_15__SCAN_IN), .B1(n6174), .B2(
        P2_REG1_REG_15__SCAN_IN), .ZN(n6007) );
  NAND2_X1 U7767 ( .A1(n6175), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n6006) );
  OR2_X1 U7768 ( .A1(n8501), .A2(n8406), .ZN(n6201) );
  INV_X1 U7769 ( .A(n6201), .ZN(n6009) );
  NAND2_X1 U7770 ( .A1(n8501), .A2(n8406), .ZN(n6302) );
  NAND2_X1 U7771 ( .A1(n6983), .A2(n6182), .ZN(n6017) );
  MUX2_X1 U7772 ( .A(n6011), .B(n6012), .S(P2_IR_REG_16__SCAN_IN), .Z(n6013)
         );
  INV_X1 U7773 ( .A(n6013), .ZN(n6015) );
  AND2_X1 U7774 ( .A1(n6015), .A2(n6026), .ZN(n8123) );
  AOI22_X1 U7775 ( .A1(n6139), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n4292), .B2(
        n8123), .ZN(n6016) );
  NAND2_X1 U7776 ( .A1(n6019), .A2(n4584), .ZN(n6020) );
  NAND2_X1 U7777 ( .A1(n6030), .A2(n6020), .ZN(n8415) );
  OR2_X1 U7778 ( .A1(n8415), .A2(n6076), .ZN(n6023) );
  AOI22_X1 U7779 ( .A1(n4280), .A2(P2_REG0_REG_16__SCAN_IN), .B1(n6174), .B2(
        P2_REG1_REG_16__SCAN_IN), .ZN(n6022) );
  INV_X1 U7780 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8416) );
  OR2_X1 U7781 ( .A1(n5892), .A2(n8416), .ZN(n6021) );
  NAND2_X1 U7782 ( .A1(n8494), .A2(n8042), .ZN(n6298) );
  INV_X1 U7783 ( .A(n6298), .ZN(n6024) );
  NAND2_X1 U7784 ( .A1(n7107), .A2(n6182), .ZN(n6029) );
  NAND2_X1 U7785 ( .A1(n6026), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6025) );
  MUX2_X1 U7786 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6025), .S(
        P2_IR_REG_17__SCAN_IN), .Z(n6027) );
  NOR2_X2 U7787 ( .A1(n6026), .A2(P2_IR_REG_17__SCAN_IN), .ZN(n6050) );
  INV_X1 U7788 ( .A(n6050), .ZN(n6037) );
  NAND2_X1 U7789 ( .A1(n6027), .A2(n6037), .ZN(n8127) );
  INV_X1 U7790 ( .A(n8127), .ZN(n10002) );
  AOI22_X1 U7791 ( .A1(n6139), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n4293), .B2(
        n10002), .ZN(n6028) );
  NAND2_X1 U7792 ( .A1(n6030), .A2(n4585), .ZN(n6031) );
  NAND2_X1 U7793 ( .A1(n6041), .A2(n6031), .ZN(n8393) );
  OR2_X1 U7794 ( .A1(n8393), .A2(n6076), .ZN(n6036) );
  INV_X1 U7795 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n8128) );
  NAND2_X1 U7796 ( .A1(n4280), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n6033) );
  INV_X1 U7797 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8394) );
  OR2_X1 U7798 ( .A1(n5892), .A2(n8394), .ZN(n6032) );
  OAI211_X1 U7799 ( .C1(n4289), .C2(n8128), .A(n6033), .B(n6032), .ZN(n6034)
         );
  INV_X1 U7800 ( .A(n6034), .ZN(n6035) );
  NAND2_X1 U7801 ( .A1(n8490), .A2(n8408), .ZN(n6299) );
  NAND2_X1 U7802 ( .A1(n6037), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6038) );
  XNOR2_X1 U7803 ( .A(n6038), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8137) );
  AOI22_X1 U7804 ( .A1(n6139), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n4292), .B2(
        n8137), .ZN(n6039) );
  INV_X1 U7805 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n6040) );
  NAND2_X1 U7806 ( .A1(n6041), .A2(n6040), .ZN(n6042) );
  NAND2_X1 U7807 ( .A1(n6053), .A2(n6042), .ZN(n8362) );
  INV_X1 U7808 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8142) );
  NAND2_X1 U7809 ( .A1(n4280), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n6044) );
  NAND2_X1 U7810 ( .A1(n6175), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n6043) );
  OAI211_X1 U7811 ( .C1(n4289), .C2(n8142), .A(n6044), .B(n6043), .ZN(n6045)
         );
  INV_X1 U7812 ( .A(n6045), .ZN(n6046) );
  NAND2_X1 U7813 ( .A1(n6047), .A2(n6046), .ZN(n8343) );
  INV_X1 U7814 ( .A(n8343), .ZN(n8169) );
  NAND2_X1 U7815 ( .A1(n7209), .A2(n6182), .ZN(n6052) );
  AOI22_X1 U7816 ( .A1(n4293), .A2(n4291), .B1(n6139), .B2(
        P1_DATAO_REG_19__SCAN_IN), .ZN(n6051) );
  NAND2_X1 U7817 ( .A1(n6053), .A2(n10237), .ZN(n6054) );
  NAND2_X1 U7818 ( .A1(n6063), .A2(n6054), .ZN(n8354) );
  INV_X1 U7819 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n8145) );
  NAND2_X1 U7820 ( .A1(n4280), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n6056) );
  INV_X1 U7821 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n8355) );
  OR2_X1 U7822 ( .A1(n5892), .A2(n8355), .ZN(n6055) );
  OAI211_X1 U7823 ( .C1(n4289), .C2(n8145), .A(n6056), .B(n6055), .ZN(n6057)
         );
  INV_X1 U7824 ( .A(n6057), .ZN(n6058) );
  INV_X1 U7825 ( .A(n8373), .ZN(n8170) );
  NOR2_X1 U7826 ( .A1(n8482), .A2(n8170), .ZN(n6317) );
  AND2_X1 U7827 ( .A1(n8482), .A2(n8170), .ZN(n6314) );
  NOR2_X1 U7828 ( .A1(n6317), .A2(n6314), .ZN(n8342) );
  NAND2_X1 U7829 ( .A1(n7268), .A2(n6182), .ZN(n6060) );
  NAND2_X1 U7830 ( .A1(n6139), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n6059) );
  INV_X1 U7831 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n6062) );
  NAND2_X1 U7832 ( .A1(n6063), .A2(n6062), .ZN(n6064) );
  AND2_X1 U7833 ( .A1(n6074), .A2(n6064), .ZN(n8328) );
  NAND2_X1 U7834 ( .A1(n8328), .A2(n6138), .ZN(n6070) );
  INV_X1 U7835 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n6067) );
  NAND2_X1 U7836 ( .A1(n6175), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n6066) );
  NAND2_X1 U7837 ( .A1(n6174), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n6065) );
  OAI211_X1 U7838 ( .C1(n6179), .C2(n6067), .A(n6066), .B(n6065), .ZN(n6068)
         );
  INV_X1 U7839 ( .A(n6068), .ZN(n6069) );
  NAND2_X1 U7840 ( .A1(n8330), .A2(n8344), .ZN(n6319) );
  INV_X1 U7841 ( .A(n8344), .ZN(n8172) );
  NAND2_X1 U7842 ( .A1(n8476), .A2(n8172), .ZN(n6321) );
  NAND2_X1 U7843 ( .A1(n6319), .A2(n6321), .ZN(n8326) );
  INV_X1 U7844 ( .A(n8326), .ZN(n8332) );
  INV_X1 U7845 ( .A(n6314), .ZN(n8331) );
  NAND2_X1 U7846 ( .A1(n7287), .A2(n6182), .ZN(n6073) );
  NAND2_X1 U7847 ( .A1(n6139), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n6072) );
  NAND2_X1 U7848 ( .A1(n6074), .A2(n4588), .ZN(n6075) );
  NAND2_X1 U7849 ( .A1(n6096), .A2(n6075), .ZN(n7938) );
  INV_X1 U7850 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n6079) );
  NAND2_X1 U7851 ( .A1(n6175), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n6078) );
  NAND2_X1 U7852 ( .A1(n6174), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n6077) );
  OAI211_X1 U7853 ( .C1(n6179), .C2(n6079), .A(n6078), .B(n6077), .ZN(n6080)
         );
  INV_X1 U7854 ( .A(n6080), .ZN(n6081) );
  OR2_X1 U7855 ( .A1(n8471), .A2(n8173), .ZN(n6324) );
  NAND2_X1 U7856 ( .A1(n8471), .A2(n8173), .ZN(n6320) );
  NAND2_X1 U7857 ( .A1(n6324), .A2(n6320), .ZN(n8318) );
  NAND2_X1 U7858 ( .A1(n7349), .A2(n6182), .ZN(n6084) );
  OR2_X1 U7859 ( .A1(n4417), .A2(n10187), .ZN(n6083) );
  XNOR2_X1 U7860 ( .A(n6096), .B(P2_REG3_REG_22__SCAN_IN), .ZN(n8301) );
  NAND2_X1 U7861 ( .A1(n8301), .A2(n6138), .ZN(n6090) );
  INV_X1 U7862 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n6087) );
  NAND2_X1 U7863 ( .A1(n6174), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n6086) );
  NAND2_X1 U7864 ( .A1(n6175), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n6085) );
  OAI211_X1 U7865 ( .C1(n6179), .C2(n6087), .A(n6086), .B(n6085), .ZN(n6088)
         );
  INV_X1 U7866 ( .A(n6088), .ZN(n6089) );
  NAND2_X1 U7867 ( .A1(n8466), .A2(n8009), .ZN(n6313) );
  NAND2_X1 U7868 ( .A1(n6091), .A2(n6313), .ZN(n8307) );
  INV_X1 U7869 ( .A(n6091), .ZN(n8288) );
  NAND2_X1 U7870 ( .A1(n7506), .A2(n6182), .ZN(n6093) );
  NAND2_X1 U7871 ( .A1(n6139), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n6092) );
  INV_X1 U7872 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n6095) );
  INV_X1 U7873 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n6094) );
  OAI21_X1 U7874 ( .B1(n6096), .B2(n6095), .A(n6094), .ZN(n6097) );
  AND2_X1 U7875 ( .A1(n6097), .A2(n6105), .ZN(n8293) );
  INV_X1 U7876 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n8284) );
  NAND2_X1 U7877 ( .A1(n6174), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n6099) );
  NAND2_X1 U7878 ( .A1(n4280), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n6098) );
  OAI211_X1 U7879 ( .C1(n5892), .C2(n8284), .A(n6099), .B(n6098), .ZN(n6100)
         );
  OR2_X1 U7880 ( .A1(n8461), .A2(n8272), .ZN(n6328) );
  NAND2_X1 U7881 ( .A1(n8461), .A2(n8272), .ZN(n6327) );
  NAND2_X1 U7882 ( .A1(n6328), .A2(n6327), .ZN(n8287) );
  INV_X1 U7883 ( .A(n6327), .ZN(n6101) );
  NAND2_X1 U7884 ( .A1(n7720), .A2(n6182), .ZN(n6103) );
  NAND2_X1 U7885 ( .A1(n6139), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n6102) );
  INV_X1 U7886 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n10265) );
  NAND2_X1 U7887 ( .A1(n6105), .A2(n10265), .ZN(n6106) );
  NAND2_X1 U7888 ( .A1(n6116), .A2(n6106), .ZN(n7977) );
  INV_X1 U7889 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n6109) );
  NAND2_X1 U7890 ( .A1(n6175), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n6108) );
  NAND2_X1 U7891 ( .A1(n6174), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n6107) );
  OAI211_X1 U7892 ( .C1(n6179), .C2(n6109), .A(n6108), .B(n6107), .ZN(n6110)
         );
  INV_X1 U7893 ( .A(n6110), .ZN(n6111) );
  INV_X1 U7894 ( .A(n8291), .ZN(n7912) );
  OR2_X1 U7895 ( .A1(n8456), .A2(n7912), .ZN(n6331) );
  NAND2_X1 U7896 ( .A1(n7781), .A2(n6182), .ZN(n6114) );
  OR2_X1 U7897 ( .A1(n4417), .A2(n10263), .ZN(n6113) );
  INV_X1 U7898 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n6115) );
  NAND2_X1 U7899 ( .A1(n6116), .A2(n6115), .ZN(n6117) );
  NAND2_X1 U7900 ( .A1(n8251), .A2(n6138), .ZN(n6123) );
  INV_X1 U7901 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n6120) );
  NAND2_X1 U7902 ( .A1(n6175), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n6119) );
  NAND2_X1 U7903 ( .A1(n6174), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n6118) );
  OAI211_X1 U7904 ( .C1(n6179), .C2(n6120), .A(n6119), .B(n6118), .ZN(n6121)
         );
  INV_X1 U7905 ( .A(n6121), .ZN(n6122) );
  NAND2_X1 U7906 ( .A1(n8452), .A2(n8273), .ZN(n6336) );
  INV_X1 U7907 ( .A(n8254), .ZN(n6333) );
  NAND2_X1 U7908 ( .A1(n7814), .A2(n6182), .ZN(n6125) );
  NAND2_X1 U7909 ( .A1(n6139), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n6124) );
  INV_X1 U7910 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n10241) );
  NAND2_X1 U7911 ( .A1(n6126), .A2(n10241), .ZN(n6127) );
  INV_X1 U7912 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n10256) );
  NAND2_X1 U7913 ( .A1(n6175), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n6129) );
  NAND2_X1 U7914 ( .A1(n6174), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n6128) );
  OAI211_X1 U7915 ( .C1(n6179), .C2(n10256), .A(n6129), .B(n6128), .ZN(n6130)
         );
  NAND2_X1 U7916 ( .A1(n8447), .A2(n8179), .ZN(n6337) );
  INV_X1 U7917 ( .A(n6338), .ZN(n6131) );
  NAND2_X1 U7918 ( .A1(n7820), .A2(n6182), .ZN(n6133) );
  NAND2_X1 U7919 ( .A1(n6139), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n6132) );
  INV_X1 U7920 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n6136) );
  NAND2_X1 U7921 ( .A1(n6174), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n6135) );
  NAND2_X1 U7922 ( .A1(n6175), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n6134) );
  OAI211_X1 U7923 ( .C1(n6136), .C2(n6179), .A(n6135), .B(n6134), .ZN(n6137)
         );
  OR2_X1 U7924 ( .A1(n8441), .A2(n8239), .ZN(n6222) );
  NAND2_X1 U7925 ( .A1(n7833), .A2(n6182), .ZN(n6141) );
  NAND2_X1 U7926 ( .A1(n6139), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n6140) );
  INV_X1 U7927 ( .A(n6145), .ZN(n6143) );
  AND2_X1 U7928 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(P2_REG3_REG_28__SCAN_IN), 
        .ZN(n6142) );
  NAND2_X1 U7929 ( .A1(n6143), .A2(n6142), .ZN(n8193) );
  INV_X1 U7930 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n6144) );
  INV_X1 U7931 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n6550) );
  OAI21_X1 U7932 ( .B1(n6145), .B2(n6144), .A(n6550), .ZN(n6146) );
  NAND2_X1 U7933 ( .A1(n8193), .A2(n6146), .ZN(n8210) );
  INV_X1 U7934 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n6149) );
  NAND2_X1 U7935 ( .A1(n6175), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n6148) );
  NAND2_X1 U7936 ( .A1(n6174), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n6147) );
  OAI211_X1 U7937 ( .C1(n6179), .C2(n6149), .A(n6148), .B(n6147), .ZN(n6150)
         );
  INV_X1 U7938 ( .A(n6150), .ZN(n6151) );
  NAND2_X1 U7939 ( .A1(n8437), .A2(n8182), .ZN(n6225) );
  INV_X1 U7940 ( .A(n8184), .ZN(n6161) );
  NAND2_X1 U7941 ( .A1(n8551), .A2(n6182), .ZN(n6154) );
  INV_X1 U7942 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n10165) );
  OR2_X1 U7943 ( .A1(n4417), .A2(n10165), .ZN(n6153) );
  INV_X1 U7944 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n10161) );
  NAND2_X1 U7945 ( .A1(n4280), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n6156) );
  NAND2_X1 U7946 ( .A1(n6175), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n6155) );
  OAI211_X1 U7947 ( .C1(n4289), .C2(n10161), .A(n6156), .B(n6155), .ZN(n6157)
         );
  INV_X1 U7948 ( .A(n6157), .ZN(n6158) );
  NAND2_X1 U7949 ( .A1(n8154), .A2(n8202), .ZN(n6172) );
  INV_X1 U7950 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n7895) );
  NOR2_X1 U7951 ( .A1(n4417), .A2(n7895), .ZN(n6162) );
  NAND2_X1 U7952 ( .A1(n4280), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n6167) );
  INV_X1 U7953 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n6163) );
  OR2_X1 U7954 ( .A1(n4289), .A2(n6163), .ZN(n6166) );
  INV_X1 U7955 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n8155) );
  OR2_X1 U7956 ( .A1(n5892), .A2(n8155), .ZN(n6165) );
  AND3_X1 U7957 ( .A1(n6167), .A2(n6166), .A3(n6165), .ZN(n6695) );
  NOR2_X1 U7958 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), .ZN(
        n6168) );
  NAND2_X1 U7959 ( .A1(n6170), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6169) );
  NAND2_X1 U7960 ( .A1(n6695), .A2(n4446), .ZN(n6173) );
  OAI21_X1 U7961 ( .B1(n8429), .B2(n6173), .A(n6172), .ZN(n6181) );
  INV_X1 U7962 ( .A(n6173), .ZN(n6180) );
  INV_X1 U7963 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n6178) );
  NAND2_X1 U7964 ( .A1(n6174), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n6177) );
  NAND2_X1 U7965 ( .A1(n6175), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n6176) );
  OAI211_X1 U7966 ( .C1(n6179), .C2(n6178), .A(n6177), .B(n6176), .ZN(n8187)
         );
  INV_X1 U7967 ( .A(n8187), .ZN(n6185) );
  OR2_X1 U7968 ( .A1(n8159), .A2(n6185), .ZN(n6348) );
  NAND2_X1 U7969 ( .A1(n8544), .A2(n6182), .ZN(n6184) );
  OR2_X1 U7970 ( .A1(n4417), .A2(n8546), .ZN(n6183) );
  NAND2_X1 U7971 ( .A1(n8159), .A2(n6185), .ZN(n6344) );
  XNOR2_X1 U7972 ( .A(n6186), .B(n8392), .ZN(n6200) );
  INV_X1 U7973 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n6188) );
  NAND2_X1 U7974 ( .A1(n6189), .A2(n6188), .ZN(n6190) );
  NAND2_X1 U7975 ( .A1(n6190), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6192) );
  INV_X1 U7976 ( .A(n7036), .ZN(n6193) );
  INV_X1 U7977 ( .A(n6387), .ZN(n6471) );
  INV_X1 U7978 ( .A(n4301), .ZN(n6352) );
  NAND2_X1 U7979 ( .A1(n4446), .A2(n6352), .ZN(n7033) );
  NOR2_X1 U7980 ( .A1(n6546), .A2(P2_U3152), .ZN(n7507) );
  INV_X1 U7981 ( .A(n7507), .ZN(n6717) );
  AOI21_X1 U7982 ( .B1(n6471), .B2(n7033), .A(n6717), .ZN(n6199) );
  NAND2_X1 U7983 ( .A1(n6200), .A2(n6199), .ZN(n6380) );
  INV_X1 U7984 ( .A(n6346), .ZN(n6218) );
  INV_X1 U7985 ( .A(n6345), .ZN(n6350) );
  INV_X1 U7986 ( .A(n8186), .ZN(n6343) );
  INV_X1 U7987 ( .A(n8287), .ZN(n6326) );
  NAND2_X1 U7988 ( .A1(n6304), .A2(n6298), .ZN(n8168) );
  NAND2_X1 U7989 ( .A1(n6201), .A2(n6302), .ZN(n7793) );
  NAND2_X1 U7990 ( .A1(n7841), .A2(n6284), .ZN(n7739) );
  INV_X1 U7991 ( .A(n7739), .ZN(n7708) );
  NAND2_X1 U7992 ( .A1(n6268), .A2(n6267), .ZN(n7219) );
  INV_X1 U7993 ( .A(n6245), .ZN(n6202) );
  AND2_X1 U7994 ( .A1(n6246), .A2(n6202), .ZN(n7514) );
  AND2_X1 U7995 ( .A1(n6384), .A2(n10090), .ZN(n6244) );
  INV_X1 U7996 ( .A(n6244), .ZN(n6203) );
  NAND2_X1 U7997 ( .A1(n7515), .A2(n6203), .ZN(n10085) );
  NOR2_X1 U7998 ( .A1(n7021), .A2(n10085), .ZN(n6204) );
  NAND4_X1 U7999 ( .A1(n7514), .A2(n6204), .A3(n6352), .A4(n10013), .ZN(n6206)
         );
  NAND2_X1 U8000 ( .A1(n6205), .A2(n7030), .ZN(n7583) );
  NOR2_X1 U8001 ( .A1(n6206), .A2(n7583), .ZN(n6207) );
  XNOR2_X1 U8002 ( .A(n8066), .B(n4284), .ZN(n7032) );
  AND4_X1 U8003 ( .A1(n7221), .A2(n6207), .A3(n7451), .A4(n7032), .ZN(n6208)
         );
  NAND3_X1 U8004 ( .A1(n7539), .A2(n6208), .A3(n7227), .ZN(n6209) );
  NOR2_X1 U8005 ( .A1(n6209), .A2(n7736), .ZN(n6210) );
  NAND4_X1 U8006 ( .A1(n7744), .A2(n7843), .A3(n7708), .A4(n6210), .ZN(n6211)
         );
  NOR4_X1 U8007 ( .A1(n8168), .A2(n7793), .A3(n7768), .A4(n6211), .ZN(n6212)
         );
  NAND4_X1 U8008 ( .A1(n8342), .A2(n4719), .A3(n8368), .A4(n6212), .ZN(n6213)
         );
  NOR4_X1 U8009 ( .A1(n8307), .A2(n8326), .A3(n8318), .A4(n6213), .ZN(n6214)
         );
  NAND4_X1 U8010 ( .A1(n6333), .A2(n6326), .A3(n6214), .A4(n8270), .ZN(n6215)
         );
  NOR4_X1 U8011 ( .A1(n8207), .A2(n8225), .A3(n8237), .A4(n6215), .ZN(n6216)
         );
  NAND4_X1 U8012 ( .A1(n6350), .A2(n6343), .A3(n6216), .A4(n6348), .ZN(n6217)
         );
  NOR2_X1 U8013 ( .A1(n6218), .A2(n6217), .ZN(n6219) );
  XNOR2_X1 U8014 ( .A(n6219), .B(n4291), .ZN(n6220) );
  OAI22_X1 U8015 ( .A1(n6220), .A2(n4446), .B1(n6352), .B2(n7034), .ZN(n6221)
         );
  NAND2_X1 U8016 ( .A1(n6221), .A2(n7507), .ZN(n6376) );
  NAND2_X1 U8017 ( .A1(n8184), .A2(n6222), .ZN(n6226) );
  NAND3_X1 U8018 ( .A1(n6226), .A2(n6347), .A3(n6225), .ZN(n6231) );
  NOR2_X1 U8019 ( .A1(n8202), .A2(n6349), .ZN(n6229) );
  NAND2_X1 U8020 ( .A1(n8202), .A2(n6349), .ZN(n6227) );
  NAND2_X1 U8021 ( .A1(n8154), .A2(n6227), .ZN(n6228) );
  OAI21_X1 U8022 ( .B1(n8154), .B2(n6229), .A(n6228), .ZN(n6230) );
  OAI21_X1 U8023 ( .B1(n8186), .B2(n6231), .A(n6230), .ZN(n6232) );
  INV_X1 U8024 ( .A(n6258), .ZN(n6234) );
  NAND2_X1 U8025 ( .A1(n6234), .A2(n6233), .ZN(n6239) );
  NAND2_X1 U8026 ( .A1(n6236), .A2(n6235), .ZN(n6238) );
  INV_X1 U8027 ( .A(n6262), .ZN(n6237) );
  AOI21_X1 U8028 ( .B1(n6239), .B2(n6238), .A(n6237), .ZN(n6265) );
  NAND2_X1 U8029 ( .A1(n6205), .A2(n6240), .ZN(n6243) );
  NAND2_X1 U8030 ( .A1(n6266), .A2(n6241), .ZN(n6242) );
  AOI21_X1 U8031 ( .B1(n6258), .B2(n6243), .A(n6242), .ZN(n6261) );
  NOR2_X1 U8032 ( .A1(n6245), .A2(n6244), .ZN(n6253) );
  INV_X1 U8033 ( .A(n6253), .ZN(n6248) );
  NAND3_X1 U8034 ( .A1(n6248), .A2(n6247), .A3(n6246), .ZN(n6249) );
  NAND2_X1 U8035 ( .A1(n6249), .A2(n6252), .ZN(n6257) );
  CLKBUF_X1 U8036 ( .A(n6250), .Z(n6251) );
  INV_X1 U8037 ( .A(n6251), .ZN(n6255) );
  NAND3_X1 U8038 ( .A1(n6253), .A2(n4446), .A3(n6252), .ZN(n6254) );
  NAND2_X1 U8039 ( .A1(n6255), .A2(n6254), .ZN(n6256) );
  NAND3_X1 U8040 ( .A1(n6259), .A2(n6258), .A3(n10013), .ZN(n6260) );
  NAND2_X1 U8041 ( .A1(n6263), .A2(n6262), .ZN(n6264) );
  MUX2_X1 U8042 ( .A(n6268), .B(n6267), .S(n6349), .Z(n6269) );
  INV_X1 U8043 ( .A(n7389), .ZN(n7383) );
  AOI21_X1 U8044 ( .B1(n7383), .B2(n8063), .A(n6347), .ZN(n6270) );
  NAND4_X1 U8045 ( .A1(n6271), .A2(n6270), .A3(n7841), .A4(n6278), .ZN(n6274)
         );
  NAND3_X1 U8046 ( .A1(n7545), .A2(n6347), .A3(n6272), .ZN(n6273) );
  NAND2_X1 U8047 ( .A1(n7881), .A2(n6349), .ZN(n6277) );
  OAI21_X1 U8048 ( .B1(n7545), .B2(n6347), .A(n8061), .ZN(n6275) );
  NAND2_X1 U8049 ( .A1(n6275), .A2(n7704), .ZN(n6276) );
  OAI21_X1 U8050 ( .B1(n6277), .B2(n7545), .A(n6276), .ZN(n6281) );
  AOI21_X1 U8051 ( .B1(n6278), .B2(n7881), .A(n6349), .ZN(n6280) );
  NAND2_X1 U8052 ( .A1(n7704), .A2(n6278), .ZN(n6279) );
  AOI22_X1 U8053 ( .A1(n6281), .A2(n7841), .B1(n6280), .B2(n6279), .ZN(n6282)
         );
  NAND2_X1 U8054 ( .A1(n6286), .A2(n7841), .ZN(n6283) );
  NAND2_X1 U8055 ( .A1(n6283), .A2(n6285), .ZN(n6289) );
  NAND2_X1 U8056 ( .A1(n6285), .A2(n6284), .ZN(n6287) );
  NAND2_X1 U8057 ( .A1(n6287), .A2(n6286), .ZN(n6288) );
  MUX2_X1 U8058 ( .A(n6289), .B(n6288), .S(n6349), .Z(n6290) );
  MUX2_X1 U8059 ( .A(n6291), .B(n7770), .S(n6349), .Z(n6292) );
  MUX2_X1 U8060 ( .A(n6295), .B(n6294), .S(n6349), .Z(n6296) );
  INV_X1 U8061 ( .A(n6296), .ZN(n6297) );
  OR3_X1 U8062 ( .A1(n8501), .A2(n8406), .A3(n6349), .ZN(n6301) );
  NAND2_X1 U8063 ( .A1(n6309), .A2(n6299), .ZN(n6300) );
  INV_X1 U8064 ( .A(n8168), .ZN(n8404) );
  INV_X1 U8065 ( .A(n6315), .ZN(n6305) );
  AOI21_X1 U8066 ( .B1(n6306), .B2(n4719), .A(n6305), .ZN(n6307) );
  NAND2_X1 U8067 ( .A1(n6308), .A2(n6307), .ZN(n6316) );
  AOI21_X1 U8068 ( .B1(n6316), .B2(n6309), .A(n6317), .ZN(n6311) );
  NAND2_X1 U8069 ( .A1(n6321), .A2(n8331), .ZN(n6310) );
  AOI21_X1 U8070 ( .B1(n6316), .B2(n6315), .A(n6314), .ZN(n6323) );
  INV_X1 U8071 ( .A(n6317), .ZN(n6318) );
  NAND2_X1 U8072 ( .A1(n6319), .A2(n6318), .ZN(n6322) );
  MUX2_X1 U8073 ( .A(n6328), .B(n6327), .S(n6349), .Z(n6329) );
  NAND2_X1 U8074 ( .A1(n8456), .A2(n7912), .ZN(n6330) );
  MUX2_X1 U8075 ( .A(n6331), .B(n6330), .S(n6347), .Z(n6332) );
  AOI21_X1 U8076 ( .B1(n6337), .B2(n6336), .A(n6347), .ZN(n6339) );
  AND2_X1 U8077 ( .A1(n8441), .A2(n8239), .ZN(n6340) );
  OAI21_X1 U8078 ( .B1(n8207), .B2(n6340), .A(n6349), .ZN(n6341) );
  NAND3_X1 U8079 ( .A1(n8437), .A2(n8182), .A3(n6347), .ZN(n6342) );
  NAND4_X1 U8080 ( .A1(n6351), .A2(n6350), .A3(n6349), .A4(n6348), .ZN(n6353)
         );
  INV_X1 U8081 ( .A(P2_B_REG_SCAN_IN), .ZN(n10176) );
  NOR2_X1 U8082 ( .A1(n6026), .A2(n6358), .ZN(n6363) );
  NAND2_X1 U8083 ( .A1(n6363), .A2(n6359), .ZN(n6366) );
  NAND2_X1 U8084 ( .A1(n6366), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6360) );
  MUX2_X1 U8085 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6360), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n6362) );
  NAND2_X1 U8086 ( .A1(n6362), .A2(n6361), .ZN(n7819) );
  INV_X1 U8087 ( .A(n6363), .ZN(n6364) );
  NAND2_X1 U8088 ( .A1(n6364), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6365) );
  MUX2_X1 U8089 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6365), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n6367) );
  NAND2_X1 U8090 ( .A1(n6367), .A2(n6366), .ZN(n7785) );
  INV_X1 U8091 ( .A(n6371), .ZN(n6372) );
  NOR4_X1 U8092 ( .A1(n6518), .A2(n6369), .A3(n6545), .A4(n8405), .ZN(n6373)
         );
  AOI211_X1 U8093 ( .C1(n7507), .C2(n6223), .A(n10176), .B(n6373), .ZN(n6374)
         );
  INV_X1 U8094 ( .A(n6374), .ZN(n6375) );
  NAND2_X1 U8095 ( .A1(n6380), .A2(n6379), .ZN(P2_U3244) );
  NAND2_X1 U8096 ( .A1(n4446), .A2(n7381), .ZN(n7375) );
  AND2_X4 U8097 ( .A1(n6382), .A2(n7375), .ZN(n6494) );
  NAND2_X1 U8098 ( .A1(n4302), .A2(n6383), .ZN(n6913) );
  NAND2_X1 U8099 ( .A1(n6494), .A2(n10090), .ZN(n6386) );
  INV_X1 U8100 ( .A(n7018), .ZN(n6385) );
  NAND2_X1 U8101 ( .A1(n6466), .A2(n6385), .ZN(n7858) );
  OAI21_X1 U8102 ( .B1(n6912), .B2(n6913), .A(n6914), .ZN(n6389) );
  NAND2_X1 U8103 ( .A1(n6912), .A2(n6913), .ZN(n6951) );
  XNOR2_X1 U8104 ( .A(n6494), .B(n5841), .ZN(n7917) );
  NAND2_X1 U8105 ( .A1(n4302), .A2(n6388), .ZN(n6390) );
  NAND2_X1 U8106 ( .A1(n7917), .A2(n6390), .ZN(n6953) );
  NAND3_X1 U8107 ( .A1(n6389), .A2(n6951), .A3(n6953), .ZN(n6393) );
  INV_X1 U8108 ( .A(n7917), .ZN(n6392) );
  INV_X1 U8109 ( .A(n6390), .ZN(n6391) );
  NAND2_X1 U8110 ( .A1(n6392), .A2(n6391), .ZN(n6954) );
  NAND2_X1 U8111 ( .A1(n6393), .A2(n6954), .ZN(n7046) );
  INV_X1 U8112 ( .A(n10056), .ZN(n7923) );
  AND2_X1 U8113 ( .A1(n4302), .A2(n8068), .ZN(n6395) );
  NAND2_X1 U8114 ( .A1(n6394), .A2(n6395), .ZN(n7050) );
  AND2_X1 U8115 ( .A1(n4302), .A2(n8067), .ZN(n6397) );
  NAND2_X1 U8116 ( .A1(n7049), .A2(n6397), .ZN(n6399) );
  NAND2_X1 U8117 ( .A1(n7050), .A2(n6399), .ZN(n6404) );
  INV_X1 U8118 ( .A(n6394), .ZN(n7191) );
  INV_X1 U8119 ( .A(n6395), .ZN(n6396) );
  INV_X1 U8120 ( .A(n6397), .ZN(n7048) );
  AND2_X1 U8121 ( .A1(n7048), .A2(n6398), .ZN(n7051) );
  XNOR2_X1 U8122 ( .A(n6400), .B(n7526), .ZN(n7199) );
  AND2_X1 U8123 ( .A1(n4302), .A2(n8066), .ZN(n6401) );
  NAND2_X1 U8124 ( .A1(n7199), .A2(n6401), .ZN(n6405) );
  XNOR2_X1 U8125 ( .A(n6510), .B(n7454), .ZN(n6409) );
  INV_X1 U8126 ( .A(n7059), .ZN(n8065) );
  NAND2_X1 U8127 ( .A1(n4302), .A2(n8065), .ZN(n6407) );
  XNOR2_X1 U8128 ( .A(n6409), .B(n6407), .ZN(n7205) );
  INV_X1 U8129 ( .A(n6407), .ZN(n6408) );
  OR2_X1 U8130 ( .A1(n6409), .A2(n6408), .ZN(n6410) );
  XNOR2_X1 U8131 ( .A(n7216), .B(n6510), .ZN(n6411) );
  INV_X1 U8132 ( .A(n7135), .ZN(n8064) );
  AND2_X1 U8133 ( .A1(n4302), .A2(n8064), .ZN(n6412) );
  NAND2_X1 U8134 ( .A1(n6411), .A2(n6412), .ZN(n6416) );
  INV_X1 U8135 ( .A(n6411), .ZN(n7131) );
  INV_X1 U8136 ( .A(n6412), .ZN(n6413) );
  NAND2_X1 U8137 ( .A1(n7131), .A2(n6413), .ZN(n6414) );
  NAND2_X1 U8138 ( .A1(n6416), .A2(n6414), .ZN(n7062) );
  XNOR2_X1 U8139 ( .A(n7389), .B(n6510), .ZN(n7886) );
  AND2_X1 U8140 ( .A1(n6471), .A2(n8063), .ZN(n6417) );
  NAND2_X1 U8141 ( .A1(n7886), .A2(n6417), .ZN(n6422) );
  INV_X1 U8142 ( .A(n7886), .ZN(n6419) );
  INV_X1 U8143 ( .A(n6417), .ZN(n6418) );
  NAND2_X1 U8144 ( .A1(n6419), .A2(n6418), .ZN(n6420) );
  AND2_X1 U8145 ( .A1(n6422), .A2(n6420), .ZN(n7129) );
  XNOR2_X1 U8146 ( .A(n7885), .B(n6510), .ZN(n6424) );
  INV_X1 U8147 ( .A(n7565), .ZN(n8062) );
  NAND2_X1 U8148 ( .A1(n4302), .A2(n8062), .ZN(n6425) );
  XNOR2_X1 U8149 ( .A(n6424), .B(n6425), .ZN(n7888) );
  AND2_X1 U8150 ( .A1(n7888), .A2(n6422), .ZN(n6423) );
  INV_X1 U8151 ( .A(n6424), .ZN(n6426) );
  NAND2_X1 U8152 ( .A1(n6426), .A2(n6425), .ZN(n6427) );
  AND2_X1 U8153 ( .A1(n6471), .A2(n8061), .ZN(n6429) );
  NAND2_X1 U8154 ( .A1(n6428), .A2(n6429), .ZN(n6433) );
  INV_X1 U8155 ( .A(n6429), .ZN(n6430) );
  NAND2_X1 U8156 ( .A1(n6433), .A2(n6431), .ZN(n7562) );
  NAND2_X1 U8157 ( .A1(n7399), .A2(n6433), .ZN(n6434) );
  XNOR2_X1 U8158 ( .A(n7737), .B(n6510), .ZN(n6437) );
  INV_X1 U8159 ( .A(n7846), .ZN(n8060) );
  NAND2_X1 U8160 ( .A1(n6471), .A2(n8060), .ZN(n6435) );
  XNOR2_X1 U8161 ( .A(n6437), .B(n6435), .ZN(n7400) );
  NAND2_X1 U8162 ( .A1(n6434), .A2(n7400), .ZN(n7403) );
  INV_X1 U8163 ( .A(n6435), .ZN(n6436) );
  NAND2_X1 U8164 ( .A1(n6437), .A2(n6436), .ZN(n6438) );
  NAND2_X1 U8165 ( .A1(n7403), .A2(n6438), .ZN(n7592) );
  XNOR2_X1 U8166 ( .A(n8519), .B(n6494), .ZN(n6439) );
  NAND2_X1 U8167 ( .A1(n6471), .A2(n8059), .ZN(n6440) );
  NAND2_X1 U8168 ( .A1(n6439), .A2(n6440), .ZN(n7591) );
  NAND2_X1 U8169 ( .A1(n7592), .A2(n7591), .ZN(n6443) );
  INV_X1 U8170 ( .A(n6439), .ZN(n6442) );
  INV_X1 U8171 ( .A(n6440), .ZN(n6441) );
  NAND2_X1 U8172 ( .A1(n6442), .A2(n6441), .ZN(n7590) );
  NAND2_X1 U8173 ( .A1(n6443), .A2(n7590), .ZN(n7991) );
  XNOR2_X1 U8174 ( .A(n8511), .B(n6510), .ZN(n6446) );
  INV_X1 U8175 ( .A(n7845), .ZN(n8058) );
  NAND2_X1 U8176 ( .A1(n6471), .A2(n8058), .ZN(n6444) );
  XNOR2_X1 U8177 ( .A(n6446), .B(n6444), .ZN(n7992) );
  INV_X1 U8178 ( .A(n6444), .ZN(n6445) );
  NAND2_X1 U8179 ( .A1(n6446), .A2(n6445), .ZN(n6447) );
  XNOR2_X1 U8180 ( .A(n8506), .B(n6494), .ZN(n6448) );
  NAND2_X1 U8181 ( .A1(n8057), .A2(n4302), .ZN(n6449) );
  NAND2_X1 U8182 ( .A1(n6448), .A2(n6449), .ZN(n6454) );
  INV_X1 U8183 ( .A(n6448), .ZN(n6451) );
  INV_X1 U8184 ( .A(n6449), .ZN(n6450) );
  NAND2_X1 U8185 ( .A1(n6451), .A2(n6450), .ZN(n6452) );
  NAND2_X1 U8186 ( .A1(n6454), .A2(n6452), .ZN(n7806) );
  INV_X1 U8187 ( .A(n7806), .ZN(n6453) );
  XNOR2_X1 U8188 ( .A(n8494), .B(n6510), .ZN(n6456) );
  NOR2_X1 U8189 ( .A1(n8042), .A2(n6387), .ZN(n6457) );
  NAND2_X1 U8190 ( .A1(n6456), .A2(n6457), .ZN(n7961) );
  XNOR2_X1 U8191 ( .A(n8501), .B(n6494), .ZN(n8043) );
  INV_X1 U8192 ( .A(n8043), .ZN(n7958) );
  OR2_X1 U8193 ( .A1(n8406), .A2(n6387), .ZN(n7956) );
  INV_X1 U8194 ( .A(n7956), .ZN(n8045) );
  NAND2_X1 U8195 ( .A1(n7958), .A2(n8045), .ZN(n6455) );
  NAND3_X1 U8196 ( .A1(n7961), .A2(n8043), .A3(n7956), .ZN(n6460) );
  INV_X1 U8197 ( .A(n6456), .ZN(n6459) );
  INV_X1 U8198 ( .A(n6457), .ZN(n6458) );
  NAND2_X1 U8199 ( .A1(n6459), .A2(n6458), .ZN(n7960) );
  XNOR2_X1 U8200 ( .A(n8490), .B(n6494), .ZN(n6461) );
  NOR2_X1 U8201 ( .A1(n8408), .A2(n6387), .ZN(n6462) );
  XNOR2_X1 U8202 ( .A(n6461), .B(n6462), .ZN(n7823) );
  INV_X1 U8203 ( .A(n6461), .ZN(n6463) );
  NAND2_X1 U8204 ( .A1(n6463), .A2(n6462), .ZN(n6464) );
  NAND2_X1 U8205 ( .A1(n6465), .A2(n6464), .ZN(n8015) );
  XNOR2_X1 U8206 ( .A(n8486), .B(n6510), .ZN(n6469) );
  NAND2_X1 U8207 ( .A1(n8343), .A2(n4302), .ZN(n6467) );
  XNOR2_X1 U8208 ( .A(n6469), .B(n6467), .ZN(n8016) );
  INV_X1 U8209 ( .A(n6467), .ZN(n6468) );
  NAND2_X1 U8210 ( .A1(n6469), .A2(n6468), .ZN(n6470) );
  NAND2_X1 U8211 ( .A1(n8373), .A2(n6471), .ZN(n6473) );
  NAND2_X1 U8212 ( .A1(n6472), .A2(n6473), .ZN(n6478) );
  INV_X1 U8213 ( .A(n6472), .ZN(n6475) );
  INV_X1 U8214 ( .A(n6473), .ZN(n6474) );
  NAND2_X1 U8215 ( .A1(n6475), .A2(n6474), .ZN(n6476) );
  NAND2_X1 U8216 ( .A1(n6478), .A2(n6476), .ZN(n7929) );
  INV_X1 U8217 ( .A(n7929), .ZN(n6477) );
  XNOR2_X1 U8218 ( .A(n8330), .B(n6400), .ZN(n6479) );
  NAND2_X1 U8219 ( .A1(n8344), .A2(n6471), .ZN(n6480) );
  XNOR2_X1 U8220 ( .A(n6479), .B(n6480), .ZN(n7984) );
  INV_X1 U8221 ( .A(n6479), .ZN(n6482) );
  INV_X1 U8222 ( .A(n6480), .ZN(n6481) );
  NAND2_X1 U8223 ( .A1(n6482), .A2(n6481), .ZN(n6483) );
  XNOR2_X1 U8224 ( .A(n8317), .B(n4283), .ZN(n6484) );
  NOR2_X1 U8225 ( .A1(n8173), .A2(n6387), .ZN(n6485) );
  XNOR2_X1 U8226 ( .A(n6484), .B(n6485), .ZN(n7937) );
  INV_X1 U8227 ( .A(n6484), .ZN(n6486) );
  NAND2_X1 U8228 ( .A1(n6486), .A2(n6485), .ZN(n6487) );
  NAND2_X1 U8229 ( .A1(n6488), .A2(n6487), .ZN(n6492) );
  XNOR2_X1 U8230 ( .A(n8466), .B(n6494), .ZN(n6490) );
  XNOR2_X1 U8231 ( .A(n6492), .B(n6490), .ZN(n8010) );
  OR2_X1 U8232 ( .A1(n8009), .A2(n6387), .ZN(n6489) );
  NAND2_X1 U8233 ( .A1(n8010), .A2(n6489), .ZN(n8014) );
  INV_X1 U8234 ( .A(n6490), .ZN(n6491) );
  OR2_X1 U8235 ( .A1(n6492), .A2(n6491), .ZN(n6493) );
  NAND2_X1 U8236 ( .A1(n8014), .A2(n6493), .ZN(n6497) );
  XNOR2_X1 U8237 ( .A(n8461), .B(n6494), .ZN(n6496) );
  XNOR2_X1 U8238 ( .A(n8456), .B(n6510), .ZN(n6498) );
  AND2_X1 U8239 ( .A1(n8291), .A2(n6471), .ZN(n6499) );
  NOR2_X1 U8240 ( .A1(n7906), .A2(n6495), .ZN(n6500) );
  NAND2_X1 U8241 ( .A1(n6497), .A2(n6496), .ZN(n7907) );
  NOR2_X1 U8242 ( .A1(n8272), .A2(n6387), .ZN(n7908) );
  NAND2_X1 U8243 ( .A1(n7907), .A2(n7908), .ZN(n7970) );
  INV_X1 U8244 ( .A(n6498), .ZN(n7972) );
  INV_X1 U8245 ( .A(n6499), .ZN(n7974) );
  XNOR2_X1 U8246 ( .A(n8253), .B(n6510), .ZN(n7945) );
  NOR2_X1 U8247 ( .A1(n8273), .A2(n6387), .ZN(n7944) );
  XNOR2_X1 U8248 ( .A(n8447), .B(n6400), .ZN(n7898) );
  NOR2_X1 U8249 ( .A1(n8179), .A2(n6387), .ZN(n6501) );
  NAND2_X1 U8250 ( .A1(n7898), .A2(n6501), .ZN(n6502) );
  OAI21_X1 U8251 ( .B1(n7898), .B2(n6501), .A(n6502), .ZN(n8026) );
  INV_X1 U8252 ( .A(n6502), .ZN(n6508) );
  XNOR2_X1 U8253 ( .A(n8441), .B(n6400), .ZN(n6503) );
  NOR2_X1 U8254 ( .A1(n8239), .A2(n6387), .ZN(n6504) );
  NAND2_X1 U8255 ( .A1(n6503), .A2(n6504), .ZN(n6509) );
  INV_X1 U8256 ( .A(n6503), .ZN(n6506) );
  INV_X1 U8257 ( .A(n6504), .ZN(n6505) );
  NAND2_X1 U8258 ( .A1(n6506), .A2(n6505), .ZN(n6507) );
  NAND2_X1 U8259 ( .A1(n7901), .A2(n6509), .ZN(n6543) );
  NOR2_X1 U8260 ( .A1(n8182), .A2(n6387), .ZN(n6511) );
  XNOR2_X1 U8261 ( .A(n6511), .B(n6510), .ZN(n6535) );
  INV_X1 U8262 ( .A(n6535), .ZN(n6536) );
  NOR3_X1 U8263 ( .A1(n8213), .A2(n10063), .A3(n6536), .ZN(n6513) );
  AOI21_X1 U8264 ( .B1(n8213), .B2(n6536), .A(n6513), .ZN(n6542) );
  XNOR2_X1 U8265 ( .A(n7722), .B(P2_B_REG_SCAN_IN), .ZN(n6514) );
  NAND2_X1 U8266 ( .A1(n6514), .A2(n7785), .ZN(n6516) );
  INV_X1 U8267 ( .A(n7819), .ZN(n6515) );
  NAND2_X1 U8268 ( .A1(n7722), .A2(n7819), .ZN(n10031) );
  AND2_X1 U8269 ( .A1(n7819), .A2(n7785), .ZN(n10037) );
  INV_X1 U8270 ( .A(n10037), .ZN(n6519) );
  NOR2_X1 U8271 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_5__SCAN_IN), .ZN(
        n10150) );
  NOR4_X1 U8272 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_31__SCAN_IN), .A3(
        P2_D_REG_2__SCAN_IN), .A4(P2_D_REG_30__SCAN_IN), .ZN(n6523) );
  NOR4_X1 U8273 ( .A1(P2_D_REG_6__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_8__SCAN_IN), .A4(P2_D_REG_10__SCAN_IN), .ZN(n6522) );
  NOR4_X1 U8274 ( .A1(P2_D_REG_23__SCAN_IN), .A2(P2_D_REG_9__SCAN_IN), .A3(
        P2_D_REG_3__SCAN_IN), .A4(P2_D_REG_4__SCAN_IN), .ZN(n6521) );
  NAND4_X1 U8275 ( .A1(n10150), .A2(n6523), .A3(n6522), .A4(n6521), .ZN(n6529)
         );
  NOR4_X1 U8276 ( .A1(P2_D_REG_14__SCAN_IN), .A2(P2_D_REG_17__SCAN_IN), .A3(
        P2_D_REG_18__SCAN_IN), .A4(P2_D_REG_19__SCAN_IN), .ZN(n6527) );
  NOR4_X1 U8277 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_12__SCAN_IN), .A3(
        P2_D_REG_16__SCAN_IN), .A4(P2_D_REG_13__SCAN_IN), .ZN(n6526) );
  NOR4_X1 U8278 ( .A1(P2_D_REG_25__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_27__SCAN_IN), .A4(P2_D_REG_28__SCAN_IN), .ZN(n6525) );
  NOR4_X1 U8279 ( .A1(P2_D_REG_20__SCAN_IN), .A2(P2_D_REG_24__SCAN_IN), .A3(
        P2_D_REG_21__SCAN_IN), .A4(P2_D_REG_22__SCAN_IN), .ZN(n6524) );
  NAND4_X1 U8280 ( .A1(n6527), .A2(n6526), .A3(n6525), .A4(n6524), .ZN(n6528)
         );
  NOR2_X1 U8281 ( .A1(n6529), .A2(n6528), .ZN(n6530) );
  NAND2_X1 U8282 ( .A1(n7015), .A2(n7013), .ZN(n7370) );
  AND2_X1 U8283 ( .A1(n4301), .A2(n4291), .ZN(n6531) );
  NAND2_X1 U8284 ( .A1(n10084), .A2(n7368), .ZN(n7012) );
  INV_X1 U8285 ( .A(n7012), .ZN(n6532) );
  NAND2_X1 U8286 ( .A1(n6544), .A2(n10022), .ZN(n6917) );
  INV_X1 U8287 ( .A(n6665), .ZN(n6716) );
  AND2_X1 U8288 ( .A1(n10077), .A2(n6716), .ZN(n6533) );
  OAI21_X1 U8289 ( .B1(n8213), .B2(n8032), .A(n8044), .ZN(n6541) );
  NOR3_X1 U8290 ( .A1(n8213), .A2(n10063), .A3(n6535), .ZN(n6538) );
  NOR2_X1 U8291 ( .A1(n8437), .A2(n6536), .ZN(n6537) );
  NAND2_X1 U8292 ( .A1(n6543), .A2(n6539), .ZN(n6540) );
  OAI211_X1 U8293 ( .C1(n6543), .C2(n6542), .A(n6541), .B(n6540), .ZN(n6553)
         );
  INV_X1 U8294 ( .A(n8239), .ZN(n8053) );
  OR2_X1 U8295 ( .A1(n7374), .A2(n7370), .ZN(n6548) );
  INV_X1 U8296 ( .A(n7371), .ZN(n7016) );
  NAND3_X1 U8297 ( .A1(n6718), .A2(n6546), .A3(n7016), .ZN(n6547) );
  AOI21_X1 U8298 ( .B1(n6548), .B2(n7012), .A(n6547), .ZN(n6549) );
  OAI22_X1 U8299 ( .A1(n8210), .A2(n8037), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6550), .ZN(n6551) );
  AOI21_X1 U8300 ( .B1(n8053), .B2(n8033), .A(n6551), .ZN(n6552) );
  INV_X1 U8301 ( .A(n8005), .ZN(n7826) );
  NAND3_X1 U8302 ( .A1(n6553), .A2(n6552), .A3(n4980), .ZN(P2_U3222) );
  INV_X1 U8303 ( .A(n7158), .ZN(n8992) );
  NAND2_X1 U8304 ( .A1(n8992), .A2(n8988), .ZN(n6603) );
  NAND2_X1 U8305 ( .A1(n9121), .A2(n8988), .ZN(n6554) );
  NAND2_X1 U8306 ( .A1(n6603), .A2(n6554), .ZN(n9802) );
  OR2_X1 U8307 ( .A1(n9802), .A2(n6555), .ZN(n6556) );
  NAND2_X1 U8308 ( .A1(n6556), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U3083) );
  INV_X1 U8309 ( .A(n6657), .ZN(n6649) );
  NAND2_X1 U8310 ( .A1(n6562), .A2(P1_U3084), .ZN(n9765) );
  OAI222_X1 U8311 ( .A1(n6649), .A2(P1_U3084), .B1(n9763), .B2(n6563), .C1(
        n4610), .C2(n9765), .ZN(P1_U3348) );
  INV_X1 U8312 ( .A(n6557), .ZN(n6558) );
  NAND2_X1 U8313 ( .A1(n6558), .A2(n9884), .ZN(n6559) );
  OAI21_X1 U8314 ( .B1(n9884), .B2(n6560), .A(n6559), .ZN(P1_U3441) );
  AND2_X1 U8315 ( .A1(n4287), .A2(P2_U3152), .ZN(n7508) );
  INV_X2 U8316 ( .A(n7508), .ZN(n8552) );
  OAI222_X1 U8317 ( .A1(n8552), .A2(n5049), .B1(n8550), .B2(n6563), .C1(
        P2_U3152), .C2(n6780), .ZN(P2_U3353) );
  INV_X1 U8318 ( .A(n6788), .ZN(n6794) );
  INV_X1 U8319 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6566) );
  INV_X1 U8320 ( .A(n6565), .ZN(n6571) );
  INV_X1 U8321 ( .A(n6803), .ZN(n6811) );
  OAI222_X1 U8322 ( .A1(n8552), .A2(n6566), .B1(n8550), .B2(n6571), .C1(
        P2_U3152), .C2(n6811), .ZN(P2_U3352) );
  INV_X1 U8323 ( .A(n6819), .ZN(n6826) );
  OAI222_X1 U8324 ( .A1(n8552), .A2(n4475), .B1(n8550), .B2(n6577), .C1(
        P2_U3152), .C2(n6826), .ZN(P2_U3354) );
  INV_X1 U8325 ( .A(n8069), .ZN(n6728) );
  OAI222_X1 U8326 ( .A1(n6728), .A2(P2_U3152), .B1(n8550), .B2(n6573), .C1(
        n6567), .C2(n8552), .ZN(P2_U3357) );
  INV_X1 U8327 ( .A(n6568), .ZN(n6582) );
  INV_X1 U8328 ( .A(n6853), .ZN(n6861) );
  OAI222_X1 U8329 ( .A1(n8552), .A2(n6569), .B1(n8550), .B2(n6582), .C1(
        P2_U3152), .C2(n6861), .ZN(P2_U3350) );
  INV_X1 U8330 ( .A(n6658), .ZN(n6688) );
  OAI222_X1 U8331 ( .A1(n6688), .A2(P1_U3084), .B1(n9763), .B2(n6571), .C1(
        n6570), .C2(n9765), .ZN(P1_U3347) );
  INV_X1 U8332 ( .A(n6642), .ZN(n6574) );
  OAI222_X1 U8333 ( .A1(P1_U3084), .A2(n6574), .B1(n9763), .B2(n6573), .C1(
        n6572), .C2(n9765), .ZN(P1_U3352) );
  INV_X1 U8334 ( .A(n6575), .ZN(n6600) );
  INV_X1 U8335 ( .A(n9765), .ZN(n9755) );
  AOI22_X1 U8336 ( .A1(n6626), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_3__SCAN_IN), .B2(n9755), .ZN(n6576) );
  OAI21_X1 U8337 ( .B1(n6600), .B2(n9763), .A(n6576), .ZN(P1_U3350) );
  INV_X1 U8338 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6578) );
  INV_X1 U8339 ( .A(n6630), .ZN(n6907) );
  OAI222_X1 U8340 ( .A1(n7782), .A2(n6578), .B1(n9763), .B2(n6577), .C1(
        P1_U3084), .C2(n6907), .ZN(P1_U3349) );
  INV_X1 U8341 ( .A(n6579), .ZN(n6596) );
  OAI222_X1 U8342 ( .A1(n6671), .A2(P1_U3084), .B1(n9763), .B2(n6596), .C1(
        n6580), .C2(n7782), .ZN(P1_U3346) );
  OAI222_X1 U8343 ( .A1(n6870), .A2(P1_U3084), .B1(n9763), .B2(n6582), .C1(
        n6581), .C2(n7782), .ZN(P1_U3345) );
  INV_X1 U8344 ( .A(n4477), .ZN(n6584) );
  INV_X1 U8345 ( .A(n6585), .ZN(n6597) );
  OAI222_X1 U8346 ( .A1(P1_U3084), .A2(n6869), .B1(n9763), .B2(n6597), .C1(
        n6586), .C2(n9765), .ZN(P1_U3344) );
  INV_X1 U8347 ( .A(n6587), .ZN(n6595) );
  AOI22_X1 U8348 ( .A1(n8108), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_10__SCAN_IN), .B2(n7508), .ZN(n6588) );
  OAI21_X1 U8349 ( .B1(n6595), .B2(n8550), .A(n6588), .ZN(P2_U3348) );
  INV_X1 U8350 ( .A(n7671), .ZN(n7242) );
  INV_X1 U8351 ( .A(n6589), .ZN(n6601) );
  OAI222_X1 U8352 ( .A1(n7242), .A2(P1_U3084), .B1(n9763), .B2(n6601), .C1(
        n6590), .C2(n7782), .ZN(P1_U3341) );
  INV_X1 U8353 ( .A(n6591), .ZN(n6599) );
  OAI222_X1 U8354 ( .A1(P1_U3084), .A2(n7237), .B1(n9763), .B2(n6599), .C1(
        n6592), .C2(n9765), .ZN(P1_U3342) );
  NAND2_X1 U8355 ( .A1(n9114), .A2(P1_U4006), .ZN(n6593) );
  OAI21_X1 U8356 ( .B1(P1_U4006), .B2(n8546), .A(n6593), .ZN(P1_U3586) );
  OAI222_X1 U8357 ( .A1(P1_U3084), .A2(n6922), .B1(n9763), .B2(n6595), .C1(
        n6594), .C2(n7782), .ZN(P1_U3343) );
  INV_X1 U8358 ( .A(n6835), .ZN(n6828) );
  OAI222_X1 U8359 ( .A1(n8552), .A2(n5053), .B1(n8550), .B2(n6596), .C1(
        P2_U3152), .C2(n6828), .ZN(P2_U3351) );
  INV_X1 U8360 ( .A(n6932), .ZN(n6939) );
  OAI222_X1 U8361 ( .A1(n8552), .A2(n6598), .B1(n8550), .B2(n6597), .C1(n6939), 
        .C2(P2_U3152), .ZN(P2_U3349) );
  INV_X1 U8362 ( .A(n6968), .ZN(n6945) );
  OAI222_X1 U8363 ( .A1(n8552), .A2(n10144), .B1(n8550), .B2(n6599), .C1(n6945), .C2(P2_U3152), .ZN(P2_U3347) );
  INV_X1 U8364 ( .A(n8082), .ZN(n6731) );
  OAI222_X1 U8365 ( .A1(n8552), .A2(n5027), .B1(n8550), .B2(n6600), .C1(
        P2_U3152), .C2(n6731), .ZN(P2_U3355) );
  INV_X1 U8366 ( .A(n7101), .ZN(n6970) );
  OAI222_X1 U8367 ( .A1(n8552), .A2(n6602), .B1(n8550), .B2(n6601), .C1(
        P2_U3152), .C2(n6970), .ZN(P2_U3346) );
  INV_X1 U8368 ( .A(n6603), .ZN(n6604) );
  OR2_X1 U8369 ( .A1(n6893), .A2(P1_U3084), .ZN(n9806) );
  NOR2_X1 U8370 ( .A1(n9802), .A2(n9806), .ZN(n9282) );
  NAND2_X1 U8371 ( .A1(n9282), .A2(n4300), .ZN(n9859) );
  AND2_X1 U8372 ( .A1(P1_U3084), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n7164) );
  NOR2_X1 U8373 ( .A1(n4300), .A2(P1_U3084), .ZN(n9805) );
  NAND2_X1 U8374 ( .A1(n9805), .A2(n6893), .ZN(n6605) );
  INV_X1 U8375 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6606) );
  XNOR2_X1 U8376 ( .A(n6626), .B(n6606), .ZN(n6610) );
  INV_X1 U8377 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n9973) );
  MUX2_X1 U8378 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n9973), .S(n9238), .Z(n9234)
         );
  INV_X1 U8379 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n9971) );
  MUX2_X1 U8380 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n9971), .S(n6642), .Z(n6639)
         );
  AND2_X1 U8381 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n6638) );
  NAND2_X1 U8382 ( .A1(n6642), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6607) );
  NAND2_X1 U8383 ( .A1(n6637), .A2(n6607), .ZN(n9233) );
  NAND2_X1 U8384 ( .A1(n4477), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6608) );
  NAND2_X1 U8385 ( .A1(n6609), .A2(n6610), .ZN(n6628) );
  OAI21_X1 U8386 ( .B1(n6610), .B2(n6609), .A(n6628), .ZN(n6611) );
  NOR2_X1 U8387 ( .A1(n9281), .A2(n6611), .ZN(n6612) );
  AOI211_X1 U8388 ( .C1(n4479), .C2(n6626), .A(n7164), .B(n6612), .ZN(n6622)
         );
  INV_X1 U8389 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n6613) );
  XNOR2_X1 U8390 ( .A(n6626), .B(n6613), .ZN(n6620) );
  INV_X1 U8391 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n6614) );
  MUX2_X1 U8392 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n6614), .S(n9238), .Z(n9241)
         );
  INV_X1 U8393 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n6615) );
  NAND2_X1 U8394 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n6891) );
  INV_X1 U8395 ( .A(n6891), .ZN(n6644) );
  NAND2_X1 U8396 ( .A1(n6642), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6616) );
  NAND2_X1 U8397 ( .A1(n6643), .A2(n6616), .ZN(n9240) );
  NAND2_X1 U8398 ( .A1(n9241), .A2(n9240), .ZN(n9239) );
  NAND2_X1 U8399 ( .A1(n4477), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6617) );
  NAND2_X1 U8400 ( .A1(n9239), .A2(n6617), .ZN(n6619) );
  INV_X1 U8401 ( .A(n9282), .ZN(n6618) );
  NAND2_X1 U8402 ( .A1(n6619), .A2(n6620), .ZN(n6624) );
  OAI211_X1 U8403 ( .C1(n6620), .C2(n6619), .A(n9855), .B(n6624), .ZN(n6621)
         );
  OAI211_X1 U8404 ( .C1(n9773), .C2(n9867), .A(n6622), .B(n6621), .ZN(P1_U3244) );
  INV_X1 U8405 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n7359) );
  XNOR2_X1 U8406 ( .A(n6657), .B(n7359), .ZN(n6650) );
  NAND2_X1 U8407 ( .A1(n6626), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6623) );
  INV_X1 U8408 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6625) );
  XNOR2_X1 U8409 ( .A(n6630), .B(n6625), .ZN(n6897) );
  NAND2_X1 U8410 ( .A1(n6898), .A2(n6897), .ZN(n6896) );
  XOR2_X1 U8411 ( .A(n6650), .B(n6651), .Z(n6636) );
  AND2_X1 U8412 ( .A1(P1_U3084), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n7611) );
  XNOR2_X1 U8413 ( .A(n6657), .B(P1_REG1_REG_5__SCAN_IN), .ZN(n6632) );
  NAND2_X1 U8414 ( .A1(n6626), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6627) );
  INV_X1 U8415 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n6629) );
  XNOR2_X1 U8416 ( .A(n6630), .B(n6629), .ZN(n6900) );
  OAI21_X1 U8417 ( .B1(P1_REG1_REG_4__SCAN_IN), .B2(n6630), .A(n6904), .ZN(
        n6631) );
  AOI211_X1 U8418 ( .C1(n6632), .C2(n6631), .A(n6656), .B(n9281), .ZN(n6633)
         );
  AOI211_X1 U8419 ( .C1(n4479), .C2(n6657), .A(n7611), .B(n6633), .ZN(n6635)
         );
  NAND2_X1 U8420 ( .A1(n9810), .A2(P1_ADDR_REG_5__SCAN_IN), .ZN(n6634) );
  OAI211_X1 U8421 ( .C1(n9839), .C2(n6636), .A(n6635), .B(n6634), .ZN(P1_U3246) );
  INV_X1 U8422 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n6648) );
  INV_X1 U8423 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n7294) );
  OAI211_X1 U8424 ( .C1(n6639), .C2(n6638), .A(n9862), .B(n6637), .ZN(n6640)
         );
  OAI21_X1 U8425 ( .B1(P1_STATE_REG_SCAN_IN), .B2(n7294), .A(n6640), .ZN(n6641) );
  AOI21_X1 U8426 ( .B1(n6642), .B2(n4479), .A(n6641), .ZN(n6647) );
  OAI211_X1 U8427 ( .C1(n6645), .C2(n6644), .A(n9855), .B(n6643), .ZN(n6646)
         );
  OAI211_X1 U8428 ( .C1(n6648), .C2(n9867), .A(n6647), .B(n6646), .ZN(P1_U3242) );
  INV_X1 U8429 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n7315) );
  XNOR2_X1 U8430 ( .A(n6671), .B(n7315), .ZN(n6654) );
  INV_X1 U8431 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n6652) );
  AOI22_X1 U8432 ( .A1(n6651), .A2(n6650), .B1(n6649), .B2(n7359), .ZN(n6685)
         );
  XOR2_X1 U8433 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n6658), .Z(n6686) );
  AOI21_X1 U8434 ( .B1(n6654), .B2(n6653), .A(n6670), .ZN(n6664) );
  AND2_X1 U8435 ( .A1(P1_U3084), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n7650) );
  NOR2_X1 U8436 ( .A1(n9859), .A2(n6671), .ZN(n6655) );
  AOI211_X1 U8437 ( .C1(n9810), .C2(P1_ADDR_REG_7__SCAN_IN), .A(n7650), .B(
        n6655), .ZN(n6663) );
  XNOR2_X1 U8438 ( .A(n6671), .B(P1_REG1_REG_7__SCAN_IN), .ZN(n6660) );
  XNOR2_X1 U8439 ( .A(n6688), .B(P1_REG1_REG_6__SCAN_IN), .ZN(n6683) );
  NAND2_X1 U8440 ( .A1(n6682), .A2(n6683), .ZN(n6681) );
  OAI21_X1 U8441 ( .B1(n6658), .B2(P1_REG1_REG_6__SCAN_IN), .A(n6681), .ZN(
        n6659) );
  NAND2_X1 U8442 ( .A1(n6659), .A2(n6660), .ZN(n6668) );
  OAI21_X1 U8443 ( .B1(n6660), .B2(n6659), .A(n6668), .ZN(n6661) );
  NAND2_X1 U8444 ( .A1(n6661), .A2(n9862), .ZN(n6662) );
  OAI211_X1 U8445 ( .C1(n6664), .C2(n9839), .A(n6663), .B(n6662), .ZN(P1_U3248) );
  OAI21_X1 U8446 ( .B1(n10029), .B2(n7507), .A(n4293), .ZN(n6667) );
  NAND2_X1 U8447 ( .A1(n10029), .A2(n6665), .ZN(n6666) );
  NOR2_X1 U8448 ( .A1(n9997), .A2(P2_U3966), .ZN(P2_U3151) );
  XNOR2_X1 U8449 ( .A(n6870), .B(P1_REG1_REG_8__SCAN_IN), .ZN(n6866) );
  INV_X1 U8450 ( .A(n6671), .ZN(n6669) );
  XOR2_X1 U8451 ( .A(n6867), .B(n6866), .Z(n6676) );
  XOR2_X1 U8452 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n6870), .Z(n6872) );
  XNOR2_X1 U8453 ( .A(n6873), .B(n6872), .ZN(n6674) );
  NAND2_X1 U8454 ( .A1(n9810), .A2(P1_ADDR_REG_8__SCAN_IN), .ZN(n6672) );
  NAND2_X1 U8455 ( .A1(P1_U3084), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n8804) );
  OAI211_X1 U8456 ( .C1(n9859), .C2(n6870), .A(n6672), .B(n8804), .ZN(n6673)
         );
  AOI21_X1 U8457 ( .B1(n6674), .B2(n9855), .A(n6673), .ZN(n6675) );
  OAI21_X1 U8458 ( .B1(n9281), .B2(n6676), .A(n6675), .ZN(P1_U3249) );
  INV_X1 U8459 ( .A(n6677), .ZN(n6680) );
  INV_X1 U8460 ( .A(n7116), .ZN(n6977) );
  OAI222_X1 U8461 ( .A1(n8552), .A2(n6678), .B1(n8550), .B2(n6680), .C1(n6977), 
        .C2(P2_U3152), .ZN(P2_U3345) );
  OAI222_X1 U8462 ( .A1(P1_U3084), .A2(n7680), .B1(n9763), .B2(n6680), .C1(
        n6679), .C2(n9765), .ZN(P1_U3340) );
  OAI21_X1 U8463 ( .B1(n6683), .B2(n6682), .A(n6681), .ZN(n6691) );
  NAND2_X1 U8464 ( .A1(P1_U3084), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n8951) );
  INV_X1 U8465 ( .A(n8951), .ZN(n6690) );
  OAI211_X1 U8466 ( .C1(n6686), .C2(n6685), .A(n9855), .B(n6684), .ZN(n6687)
         );
  OAI21_X1 U8467 ( .B1(n9859), .B2(n6688), .A(n6687), .ZN(n6689) );
  AOI211_X1 U8468 ( .C1(n9862), .C2(n6691), .A(n6690), .B(n6689), .ZN(n6692)
         );
  OAI21_X1 U8469 ( .B1(n9867), .B2(n4442), .A(n6692), .ZN(P1_U3247) );
  INV_X1 U8470 ( .A(n6693), .ZN(n6698) );
  AOI22_X1 U8471 ( .A1(n4290), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_14__SCAN_IN), .B2(n7508), .ZN(n6694) );
  OAI21_X1 U8472 ( .B1(n6698), .B2(n8550), .A(n6694), .ZN(P2_U3344) );
  NAND2_X1 U8473 ( .A1(P2_U3966), .A2(n4655), .ZN(n6696) );
  OAI21_X1 U8474 ( .B1(P2_U3966), .B2(n5728), .A(n6696), .ZN(P2_U3583) );
  OAI222_X1 U8475 ( .A1(P1_U3084), .A2(n9263), .B1(n9763), .B2(n6698), .C1(
        n6697), .C2(n9765), .ZN(P1_U3339) );
  NAND2_X1 U8476 ( .A1(n6707), .A2(n6699), .ZN(n6701) );
  NAND2_X1 U8477 ( .A1(n6701), .A2(n6700), .ZN(n7162) );
  NAND2_X1 U8478 ( .A1(n7162), .A2(n9884), .ZN(n8958) );
  NAND2_X1 U8479 ( .A1(n8993), .A2(n9194), .ZN(n6702) );
  INV_X1 U8480 ( .A(n6988), .ZN(n6703) );
  AND2_X2 U8481 ( .A1(n7158), .A2(n6703), .ZN(n7073) );
  AOI22_X1 U8482 ( .A1(n7292), .A2(n4278), .B1(n8992), .B2(
        P1_REG1_REG_0__SCAN_IN), .ZN(n6705) );
  XOR2_X1 U8483 ( .A(n6990), .B(n6991), .Z(n6892) );
  AND2_X1 U8484 ( .A1(n6709), .A2(n9961), .ZN(n6710) );
  NAND2_X1 U8485 ( .A1(n6892), .A2(n8959), .ZN(n6714) );
  OR2_X1 U8486 ( .A1(n8958), .A2(n7159), .ZN(n7088) );
  INV_X1 U8487 ( .A(n7006), .ZN(n6712) );
  INV_X1 U8488 ( .A(n8991), .ZN(n6764) );
  NAND2_X1 U8489 ( .A1(n6764), .A2(n4300), .ZN(n6711) );
  AOI22_X1 U8490 ( .A1(n7088), .A2(P1_REG3_REG_0__SCAN_IN), .B1(n8894), .B2(
        n9231), .ZN(n6713) );
  OAI211_X1 U8491 ( .C1(n8981), .C2(n6715), .A(n6714), .B(n6713), .ZN(P1_U3230) );
  NAND2_X1 U8492 ( .A1(n10029), .A2(n6716), .ZN(n6721) );
  OAI21_X1 U8493 ( .B1(n6718), .B2(P2_U3152), .A(n6717), .ZN(n6719) );
  INV_X1 U8494 ( .A(n6719), .ZN(n6720) );
  NAND2_X1 U8495 ( .A1(n6721), .A2(n6720), .ZN(n6726) );
  NAND2_X1 U8496 ( .A1(n6726), .A2(n6724), .ZN(n6722) );
  NAND2_X1 U8497 ( .A1(n6722), .A2(n8056), .ZN(n6740) );
  NAND2_X1 U8498 ( .A1(n6740), .A2(n6371), .ZN(n9988) );
  NOR2_X1 U8499 ( .A1(n6723), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7061) );
  AND2_X1 U8500 ( .A1(n6724), .A2(n6369), .ZN(n6725) );
  INV_X1 U8501 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n10092) );
  MUX2_X1 U8502 ( .A(n10092), .B(P2_REG1_REG_1__SCAN_IN), .S(n8069), .Z(n8074)
         );
  INV_X1 U8503 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n6727) );
  INV_X1 U8504 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n8075) );
  NOR3_X1 U8505 ( .A1(n8074), .A2(n6727), .A3(n8075), .ZN(n8073) );
  NOR2_X1 U8506 ( .A1(n6728), .A2(n10092), .ZN(n6783) );
  MUX2_X1 U8507 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n6729), .S(n6788), .Z(n6782)
         );
  OAI21_X1 U8508 ( .B1(n8073), .B2(n6783), .A(n6782), .ZN(n8092) );
  NAND2_X1 U8509 ( .A1(n6788), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n8091) );
  MUX2_X1 U8510 ( .A(n6730), .B(P2_REG1_REG_3__SCAN_IN), .S(n8082), .Z(n8090)
         );
  NOR2_X1 U8511 ( .A1(n6731), .A2(n6730), .ZN(n6814) );
  INV_X1 U8512 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n6732) );
  MUX2_X1 U8513 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n6732), .S(n6819), .Z(n6813)
         );
  OAI21_X1 U8514 ( .B1(n8089), .B2(n6814), .A(n6813), .ZN(n6812) );
  NAND2_X1 U8515 ( .A1(n6819), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n6772) );
  MUX2_X1 U8516 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n6733), .S(n6780), .Z(n6771)
         );
  AOI21_X1 U8517 ( .B1(n6812), .B2(n6772), .A(n6771), .ZN(n6798) );
  NOR2_X1 U8518 ( .A1(n6780), .A2(n6733), .ZN(n6797) );
  MUX2_X1 U8519 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n6734), .S(n6803), .Z(n6796)
         );
  OAI21_X1 U8520 ( .B1(n6798), .B2(n6797), .A(n6796), .ZN(n6795) );
  NAND2_X1 U8521 ( .A1(n6803), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6736) );
  MUX2_X1 U8522 ( .A(n6827), .B(P2_REG1_REG_7__SCAN_IN), .S(n6835), .Z(n6735)
         );
  AND3_X1 U8523 ( .A1(n6795), .A2(n6736), .A3(n6735), .ZN(n6737) );
  NOR3_X1 U8524 ( .A1(n9989), .A2(n6849), .A3(n6737), .ZN(n6738) );
  AOI211_X1 U8525 ( .C1(P2_ADDR_REG_7__SCAN_IN), .C2(n9997), .A(n7061), .B(
        n6738), .ZN(n6762) );
  NOR2_X1 U8526 ( .A1(n6369), .A2(n6371), .ZN(n6739) );
  MUX2_X1 U8527 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n8083), .S(n8082), .Z(n6745)
         );
  MUX2_X1 U8528 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n6741), .S(n6788), .Z(n6743)
         );
  MUX2_X1 U8529 ( .A(P2_REG2_REG_1__SCAN_IN), .B(n7518), .S(n8069), .Z(n8071)
         );
  AND2_X1 U8530 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(
        n8072) );
  NAND2_X1 U8531 ( .A1(n8069), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n6789) );
  NAND2_X1 U8532 ( .A1(n8070), .A2(n6789), .ZN(n6742) );
  NAND2_X1 U8533 ( .A1(n6743), .A2(n6742), .ZN(n8085) );
  NAND2_X1 U8534 ( .A1(n6788), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n8084) );
  NAND2_X1 U8535 ( .A1(n8085), .A2(n8084), .ZN(n6744) );
  NAND2_X1 U8536 ( .A1(n6745), .A2(n6744), .ZN(n8088) );
  NAND2_X1 U8537 ( .A1(n8082), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n6821) );
  NAND2_X1 U8538 ( .A1(n8088), .A2(n6821), .ZN(n6748) );
  MUX2_X1 U8539 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n6746), .S(n6819), .Z(n6747)
         );
  NAND2_X1 U8540 ( .A1(n6819), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n6776) );
  NAND2_X1 U8541 ( .A1(n6823), .A2(n6776), .ZN(n6750) );
  MUX2_X1 U8542 ( .A(n7527), .B(P2_REG2_REG_5__SCAN_IN), .S(n6780), .Z(n6749)
         );
  NAND2_X1 U8543 ( .A1(n6750), .A2(n6749), .ZN(n6806) );
  NAND2_X1 U8544 ( .A1(n6751), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n6805) );
  NAND2_X1 U8545 ( .A1(n6806), .A2(n6805), .ZN(n6754) );
  MUX2_X1 U8546 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n6752), .S(n6803), .Z(n6753)
         );
  NAND2_X1 U8547 ( .A1(n6754), .A2(n6753), .ZN(n6808) );
  NAND2_X1 U8548 ( .A1(n6803), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n6759) );
  NAND2_X1 U8549 ( .A1(n6808), .A2(n6759), .ZN(n6757) );
  MUX2_X1 U8550 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n6755), .S(n6835), .Z(n6756)
         );
  MUX2_X1 U8551 ( .A(n6755), .B(P2_REG2_REG_7__SCAN_IN), .S(n6835), .Z(n6758)
         );
  NAND3_X1 U8552 ( .A1(n6808), .A2(n6759), .A3(n6758), .ZN(n6760) );
  NAND3_X1 U8553 ( .A1(n9999), .A2(n6856), .A3(n6760), .ZN(n6761) );
  OAI211_X1 U8554 ( .C1(n9988), .C2(n6828), .A(n6762), .B(n6761), .ZN(P2_U3252) );
  INV_X1 U8555 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n6768) );
  OR2_X1 U8556 ( .A1(n7297), .A2(n7292), .ZN(n9132) );
  NAND2_X1 U8557 ( .A1(n9132), .A2(n7295), .ZN(n9092) );
  INV_X1 U8558 ( .A(n6763), .ZN(n6766) );
  NOR2_X1 U8559 ( .A1(n6764), .A2(n6766), .ZN(n6765) );
  AOI22_X1 U8560 ( .A1(n9092), .A2(n6765), .B1(n9562), .B2(n9231), .ZN(n9871)
         );
  NAND2_X1 U8561 ( .A1(n7292), .A2(n6766), .ZN(n9870) );
  NAND2_X1 U8562 ( .A1(n9871), .A2(n9870), .ZN(n6769) );
  NAND2_X1 U8563 ( .A1(n6769), .A2(n9970), .ZN(n6767) );
  OAI21_X1 U8564 ( .B1(n9970), .B2(n6768), .A(n6767), .ZN(P1_U3454) );
  INV_X1 U8565 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n9811) );
  NAND2_X1 U8566 ( .A1(n6769), .A2(n9986), .ZN(n6770) );
  OAI21_X1 U8567 ( .B1(n9986), .B2(n9811), .A(n6770), .ZN(P1_U3523) );
  AND2_X1 U8568 ( .A1(P2_U3152), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n7042) );
  AND3_X1 U8569 ( .A1(n6812), .A2(n6772), .A3(n6771), .ZN(n6773) );
  NOR3_X1 U8570 ( .A1(n9989), .A2(n6798), .A3(n6773), .ZN(n6774) );
  AOI211_X1 U8571 ( .C1(P2_ADDR_REG_5__SCAN_IN), .C2(n9997), .A(n7042), .B(
        n6774), .ZN(n6779) );
  MUX2_X1 U8572 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n7527), .S(n6780), .Z(n6775)
         );
  NAND3_X1 U8573 ( .A1(n6823), .A2(n6776), .A3(n6775), .ZN(n6777) );
  NAND3_X1 U8574 ( .A1(n9999), .A2(n6806), .A3(n6777), .ZN(n6778) );
  OAI211_X1 U8575 ( .C1(n9988), .C2(n6780), .A(n6779), .B(n6778), .ZN(P2_U3250) );
  NOR2_X1 U8576 ( .A1(n6781), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6787) );
  INV_X1 U8577 ( .A(n8092), .ZN(n6785) );
  NOR3_X1 U8578 ( .A1(n8073), .A2(n6783), .A3(n6782), .ZN(n6784) );
  NOR3_X1 U8579 ( .A1(n9989), .A2(n6785), .A3(n6784), .ZN(n6786) );
  AOI211_X1 U8580 ( .C1(P2_ADDR_REG_2__SCAN_IN), .C2(n9997), .A(n6787), .B(
        n6786), .ZN(n6793) );
  MUX2_X1 U8581 ( .A(n6741), .B(P2_REG2_REG_2__SCAN_IN), .S(n6788), .Z(n6790)
         );
  NAND3_X1 U8582 ( .A1(n6790), .A2(n8070), .A3(n6789), .ZN(n6791) );
  NAND3_X1 U8583 ( .A1(n9999), .A2(n8085), .A3(n6791), .ZN(n6792) );
  OAI211_X1 U8584 ( .C1(n9988), .C2(n6794), .A(n6793), .B(n6792), .ZN(P2_U3247) );
  NAND2_X1 U8585 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3152), .ZN(n7197) );
  INV_X1 U8586 ( .A(n7197), .ZN(n6802) );
  INV_X1 U8587 ( .A(n6795), .ZN(n6800) );
  NOR3_X1 U8588 ( .A1(n6798), .A2(n6797), .A3(n6796), .ZN(n6799) );
  NOR3_X1 U8589 ( .A1(n9989), .A2(n6800), .A3(n6799), .ZN(n6801) );
  AOI211_X1 U8590 ( .C1(P2_ADDR_REG_6__SCAN_IN), .C2(n9997), .A(n6802), .B(
        n6801), .ZN(n6810) );
  MUX2_X1 U8591 ( .A(n6752), .B(P2_REG2_REG_6__SCAN_IN), .S(n6803), .Z(n6804)
         );
  NAND3_X1 U8592 ( .A1(n6806), .A2(n6805), .A3(n6804), .ZN(n6807) );
  NAND3_X1 U8593 ( .A1(n9999), .A2(n6808), .A3(n6807), .ZN(n6809) );
  OAI211_X1 U8594 ( .C1(n9988), .C2(n6811), .A(n6810), .B(n6809), .ZN(P2_U3251) );
  NAND2_X1 U8595 ( .A1(P2_U3152), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n7187) );
  INV_X1 U8596 ( .A(n7187), .ZN(n6818) );
  INV_X1 U8597 ( .A(n6812), .ZN(n6816) );
  NOR3_X1 U8598 ( .A1(n8089), .A2(n6814), .A3(n6813), .ZN(n6815) );
  NOR3_X1 U8599 ( .A1(n9989), .A2(n6816), .A3(n6815), .ZN(n6817) );
  AOI211_X1 U8600 ( .C1(P2_ADDR_REG_4__SCAN_IN), .C2(n9997), .A(n6818), .B(
        n6817), .ZN(n6825) );
  MUX2_X1 U8601 ( .A(n6746), .B(P2_REG2_REG_4__SCAN_IN), .S(n6819), .Z(n6820)
         );
  NAND3_X1 U8602 ( .A1(n8088), .A2(n6821), .A3(n6820), .ZN(n6822) );
  NAND3_X1 U8603 ( .A1(n9999), .A2(n6823), .A3(n6822), .ZN(n6824) );
  OAI211_X1 U8604 ( .C1(n9988), .C2(n6826), .A(n6825), .B(n6824), .ZN(P2_U3249) );
  NAND2_X1 U8605 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3152), .ZN(n7879) );
  INV_X1 U8606 ( .A(n7879), .ZN(n6834) );
  NOR2_X1 U8607 ( .A1(n6828), .A2(n6827), .ZN(n6848) );
  MUX2_X1 U8608 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n6829), .S(n6853), .Z(n6847)
         );
  OAI21_X1 U8609 ( .B1(n6849), .B2(n6848), .A(n6847), .ZN(n6846) );
  NAND2_X1 U8610 ( .A1(n6853), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n6831) );
  MUX2_X1 U8611 ( .A(n5923), .B(P2_REG1_REG_9__SCAN_IN), .S(n6932), .Z(n6830)
         );
  AOI21_X1 U8612 ( .B1(n6846), .B2(n6831), .A(n6830), .ZN(n8101) );
  AND3_X1 U8613 ( .A1(n6846), .A2(n6831), .A3(n6830), .ZN(n6832) );
  NOR3_X1 U8614 ( .A1(n8101), .A2(n6832), .A3(n9989), .ZN(n6833) );
  AOI211_X1 U8615 ( .C1(P2_ADDR_REG_9__SCAN_IN), .C2(n9997), .A(n6834), .B(
        n6833), .ZN(n6844) );
  NAND2_X1 U8616 ( .A1(n6835), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n6855) );
  NAND2_X1 U8617 ( .A1(n6856), .A2(n6855), .ZN(n6837) );
  MUX2_X1 U8618 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n7379), .S(n6853), .Z(n6836)
         );
  NAND2_X1 U8619 ( .A1(n6837), .A2(n6836), .ZN(n6858) );
  NAND2_X1 U8620 ( .A1(n6853), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n6841) );
  NAND2_X1 U8621 ( .A1(n6858), .A2(n6841), .ZN(n6839) );
  MUX2_X1 U8622 ( .A(P2_REG2_REG_9__SCAN_IN), .B(n7394), .S(n6932), .Z(n6838)
         );
  MUX2_X1 U8623 ( .A(n7394), .B(P2_REG2_REG_9__SCAN_IN), .S(n6932), .Z(n6840)
         );
  NAND3_X1 U8624 ( .A1(n6858), .A2(n6841), .A3(n6840), .ZN(n6842) );
  NAND3_X1 U8625 ( .A1(n9999), .A2(n8111), .A3(n6842), .ZN(n6843) );
  OAI211_X1 U8626 ( .C1(n9988), .C2(n6939), .A(n6844), .B(n6843), .ZN(P2_U3254) );
  NOR2_X1 U8627 ( .A1(n6845), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7137) );
  INV_X1 U8628 ( .A(n6846), .ZN(n6851) );
  NOR3_X1 U8629 ( .A1(n6849), .A2(n6848), .A3(n6847), .ZN(n6850) );
  NOR3_X1 U8630 ( .A1(n6851), .A2(n9989), .A3(n6850), .ZN(n6852) );
  AOI211_X1 U8631 ( .C1(P2_ADDR_REG_8__SCAN_IN), .C2(n9997), .A(n7137), .B(
        n6852), .ZN(n6860) );
  MUX2_X1 U8632 ( .A(n7379), .B(P2_REG2_REG_8__SCAN_IN), .S(n6853), .Z(n6854)
         );
  NAND3_X1 U8633 ( .A1(n6856), .A2(n6855), .A3(n6854), .ZN(n6857) );
  NAND3_X1 U8634 ( .A1(n9999), .A2(n6858), .A3(n6857), .ZN(n6859) );
  OAI211_X1 U8635 ( .C1(n9988), .C2(n6861), .A(n6860), .B(n6859), .ZN(P2_U3253) );
  INV_X1 U8636 ( .A(n6862), .ZN(n6864) );
  INV_X1 U8637 ( .A(n7322), .ZN(n7692) );
  OAI222_X1 U8638 ( .A1(n8552), .A2(n10235), .B1(n8550), .B2(n6864), .C1(
        P2_U3152), .C2(n7692), .ZN(P2_U3343) );
  OAI222_X1 U8639 ( .A1(n9264), .A2(P1_U3084), .B1(n9763), .B2(n6864), .C1(
        n6863), .C2(n9765), .ZN(P1_U3338) );
  INV_X1 U8640 ( .A(n6869), .ZN(n6883) );
  XNOR2_X1 U8641 ( .A(n6883), .B(P1_REG1_REG_9__SCAN_IN), .ZN(n6880) );
  INV_X1 U8642 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n6865) );
  XOR2_X1 U8643 ( .A(n6881), .B(n6880), .Z(n6879) );
  NOR2_X1 U8644 ( .A1(n10248), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8882) );
  INV_X1 U8645 ( .A(n8882), .ZN(n6868) );
  OAI21_X1 U8646 ( .B1(n9859), .B2(n6869), .A(n6868), .ZN(n6877) );
  XOR2_X1 U8647 ( .A(P1_REG2_REG_9__SCAN_IN), .B(n6869), .Z(n6875) );
  INV_X1 U8648 ( .A(n6870), .ZN(n6871) );
  AOI211_X1 U8649 ( .C1(n6875), .C2(n6874), .A(n9839), .B(n6882), .ZN(n6876)
         );
  AOI211_X1 U8650 ( .C1(n9810), .C2(P1_ADDR_REG_9__SCAN_IN), .A(n6877), .B(
        n6876), .ZN(n6878) );
  OAI21_X1 U8651 ( .B1(n9281), .B2(n6879), .A(n6878), .ZN(P1_U3250) );
  XNOR2_X1 U8652 ( .A(n6922), .B(P1_REG1_REG_10__SCAN_IN), .ZN(n6920) );
  OAI22_X1 U8653 ( .A1(n6881), .A2(n6880), .B1(n6883), .B2(
        P1_REG1_REG_9__SCAN_IN), .ZN(n6921) );
  XOR2_X1 U8654 ( .A(n6920), .B(n6921), .Z(n6889) );
  NAND2_X1 U8655 ( .A1(P1_U3084), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n8756) );
  OAI21_X1 U8656 ( .B1(n9859), .B2(n6922), .A(n8756), .ZN(n6887) );
  XOR2_X1 U8657 ( .A(P1_REG2_REG_10__SCAN_IN), .B(n6922), .Z(n6884) );
  AOI211_X1 U8658 ( .C1(n6885), .C2(n6884), .A(n9839), .B(n6923), .ZN(n6886)
         );
  AOI211_X1 U8659 ( .C1(n9810), .C2(P1_ADDR_REG_10__SCAN_IN), .A(n6887), .B(
        n6886), .ZN(n6888) );
  OAI21_X1 U8660 ( .B1(n9281), .B2(n6889), .A(n6888), .ZN(P1_U3251) );
  MUX2_X1 U8661 ( .A(n6892), .B(n6891), .S(n6890), .Z(n6895) );
  OR2_X1 U8662 ( .A1(n6893), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n6894) );
  NAND2_X1 U8663 ( .A1(n8989), .A2(n6894), .ZN(n9800) );
  NAND2_X1 U8664 ( .A1(n9800), .A2(n4457), .ZN(n9801) );
  OAI211_X1 U8665 ( .C1(n6895), .C2(n4300), .A(P1_U4006), .B(n9801), .ZN(n9245) );
  OAI21_X1 U8666 ( .B1(n6898), .B2(n6897), .A(n6896), .ZN(n6910) );
  INV_X1 U8667 ( .A(n6899), .ZN(n6902) );
  INV_X1 U8668 ( .A(n6900), .ZN(n6901) );
  NAND2_X1 U8669 ( .A1(n6902), .A2(n6901), .ZN(n6903) );
  NAND2_X1 U8670 ( .A1(n6904), .A2(n6903), .ZN(n6905) );
  AND2_X1 U8671 ( .A1(P1_U3084), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n7260) );
  AOI21_X1 U8672 ( .B1(n9862), .B2(n6905), .A(n7260), .ZN(n6906) );
  OAI21_X1 U8673 ( .B1(n9859), .B2(n6907), .A(n6906), .ZN(n6909) );
  NOR2_X1 U8674 ( .A1(n9867), .A2(n9772), .ZN(n6908) );
  AOI211_X1 U8675 ( .C1(n9855), .C2(n6910), .A(n6909), .B(n6908), .ZN(n6911)
         );
  NAND2_X1 U8676 ( .A1(n9245), .A2(n6911), .ZN(P1_U3245) );
  INV_X1 U8677 ( .A(n8044), .ZN(n7993) );
  XOR2_X1 U8678 ( .A(n6912), .B(n6913), .Z(n6915) );
  NAND2_X1 U8679 ( .A1(n6915), .A2(n6914), .ZN(n6952) );
  OAI21_X1 U8680 ( .B1(n6915), .B2(n6914), .A(n6952), .ZN(n6916) );
  INV_X1 U8681 ( .A(n6384), .ZN(n7857) );
  OAI22_X1 U8682 ( .A1(n8405), .A2(n7857), .B1(n5842), .B2(n8407), .ZN(n7516)
         );
  AOI22_X1 U8683 ( .A1(n7993), .A2(n6916), .B1(n8005), .B2(n7516), .ZN(n6919)
         );
  NAND2_X1 U8684 ( .A1(n6917), .A2(n7016), .ZN(n7860) );
  NAND2_X1 U8685 ( .A1(n7860), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n6918) );
  OAI211_X1 U8686 ( .C1(n10041), .C2(n8032), .A(n6919), .B(n6918), .ZN(
        P2_U3224) );
  INV_X1 U8687 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n9699) );
  XNOR2_X1 U8688 ( .A(n7237), .B(n9699), .ZN(n7238) );
  INV_X1 U8689 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n7764) );
  XOR2_X1 U8690 ( .A(n7238), .B(n7239), .Z(n6931) );
  XNOR2_X1 U8691 ( .A(n7237), .B(P1_REG2_REG_11__SCAN_IN), .ZN(n6926) );
  INV_X1 U8692 ( .A(n6922), .ZN(n6924) );
  OAI21_X1 U8693 ( .B1(n6926), .B2(n6925), .A(n7244), .ZN(n6929) );
  NAND2_X1 U8694 ( .A1(n9810), .A2(P1_ADDR_REG_11__SCAN_IN), .ZN(n6927) );
  NAND2_X1 U8695 ( .A1(P1_U3084), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n8926) );
  OAI211_X1 U8696 ( .C1(n9859), .C2(n7237), .A(n6927), .B(n8926), .ZN(n6928)
         );
  AOI21_X1 U8697 ( .B1(n6929), .B2(n9855), .A(n6928), .ZN(n6930) );
  OAI21_X1 U8698 ( .B1(n9281), .B2(n6931), .A(n6930), .ZN(P1_U3252) );
  NAND2_X1 U8699 ( .A1(n6932), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n8110) );
  NAND2_X1 U8700 ( .A1(n8111), .A2(n8110), .ZN(n6934) );
  MUX2_X1 U8701 ( .A(P2_REG2_REG_10__SCAN_IN), .B(n7550), .S(n8108), .Z(n6933)
         );
  NAND2_X1 U8702 ( .A1(n6934), .A2(n6933), .ZN(n8113) );
  NAND2_X1 U8703 ( .A1(n8108), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n6935) );
  NAND2_X1 U8704 ( .A1(n8113), .A2(n6935), .ZN(n6938) );
  MUX2_X1 U8705 ( .A(n7711), .B(P2_REG2_REG_11__SCAN_IN), .S(n6968), .Z(n6937)
         );
  INV_X1 U8706 ( .A(n6962), .ZN(n6936) );
  AOI21_X1 U8707 ( .B1(n6938), .B2(n6937), .A(n6936), .ZN(n6950) );
  NOR2_X1 U8708 ( .A1(n6939), .A2(n5923), .ZN(n8100) );
  MUX2_X1 U8709 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n6940), .S(n8108), .Z(n8099)
         );
  OAI21_X1 U8710 ( .B1(n8101), .B2(n8100), .A(n8099), .ZN(n8103) );
  NAND2_X1 U8711 ( .A1(n8108), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n6942) );
  MUX2_X1 U8712 ( .A(n5948), .B(P2_REG1_REG_11__SCAN_IN), .S(n6968), .Z(n6941)
         );
  INV_X1 U8713 ( .A(n7094), .ZN(n6944) );
  NAND3_X1 U8714 ( .A1(n8103), .A2(n6942), .A3(n6941), .ZN(n6943) );
  NAND3_X1 U8715 ( .A1(n6944), .A2(n10005), .A3(n6943), .ZN(n6949) );
  NOR2_X1 U8716 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7406), .ZN(n6947) );
  NOR2_X1 U8717 ( .A1(n9988), .A2(n6945), .ZN(n6946) );
  AOI211_X1 U8718 ( .C1(P2_ADDR_REG_11__SCAN_IN), .C2(n9997), .A(n6947), .B(
        n6946), .ZN(n6948) );
  OAI211_X1 U8719 ( .C1(n6950), .C2(n9987), .A(n6949), .B(n6948), .ZN(P2_U3256) );
  NAND2_X1 U8720 ( .A1(n6952), .A2(n6951), .ZN(n6956) );
  NAND2_X1 U8721 ( .A1(n6954), .A2(n6953), .ZN(n6955) );
  OR2_X1 U8722 ( .A1(n6956), .A2(n6955), .ZN(n7919) );
  AOI21_X1 U8723 ( .B1(n6956), .B2(n6955), .A(n8044), .ZN(n6957) );
  NAND2_X1 U8724 ( .A1(n7919), .A2(n6957), .ZN(n6960) );
  INV_X1 U8725 ( .A(n8068), .ZN(n7190) );
  OAI22_X1 U8726 ( .A1(n8405), .A2(n6958), .B1(n7190), .B2(n8407), .ZN(n7572)
         );
  AOI22_X1 U8727 ( .A1(n8005), .A2(n7572), .B1(n7860), .B2(
        P2_REG3_REG_2__SCAN_IN), .ZN(n6959) );
  OAI211_X1 U8728 ( .C1(n10050), .C2(n8032), .A(n6960), .B(n6959), .ZN(
        P2_U3239) );
  OR2_X1 U8729 ( .A1(n6968), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n6961) );
  NAND2_X1 U8730 ( .A1(n6962), .A2(n6961), .ZN(n7100) );
  MUX2_X1 U8731 ( .A(n7849), .B(P2_REG2_REG_12__SCAN_IN), .S(n7101), .Z(n7099)
         );
  OR2_X1 U8732 ( .A1(n7100), .A2(n7099), .ZN(n7097) );
  NAND2_X1 U8733 ( .A1(n7101), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n6963) );
  NAND2_X1 U8734 ( .A1(n7097), .A2(n6963), .ZN(n6967) );
  MUX2_X1 U8735 ( .A(n6964), .B(P2_REG2_REG_13__SCAN_IN), .S(n7116), .Z(n6966)
         );
  INV_X1 U8736 ( .A(n7122), .ZN(n6965) );
  AOI21_X1 U8737 ( .B1(n6967), .B2(n6966), .A(n6965), .ZN(n6982) );
  AND2_X1 U8738 ( .A1(n6968), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n7093) );
  INV_X1 U8739 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n6969) );
  NAND2_X1 U8740 ( .A1(n6970), .A2(n6969), .ZN(n6971) );
  OAI21_X1 U8741 ( .B1(n6970), .B2(n6969), .A(n6971), .ZN(n7092) );
  NOR3_X1 U8742 ( .A1(n7094), .A2(n7093), .A3(n7092), .ZN(n7091) );
  INV_X1 U8743 ( .A(n6971), .ZN(n6974) );
  OR2_X1 U8744 ( .A1(n7116), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n7112) );
  NAND2_X1 U8745 ( .A1(n7116), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n6972) );
  AND2_X1 U8746 ( .A1(n7112), .A2(n6972), .ZN(n6973) );
  OAI21_X1 U8747 ( .B1(n7091), .B2(n6974), .A(n6973), .ZN(n7113) );
  INV_X1 U8748 ( .A(n7113), .ZN(n6976) );
  NOR3_X1 U8749 ( .A1(n7091), .A2(n6974), .A3(n6973), .ZN(n6975) );
  OAI21_X1 U8750 ( .B1(n6976), .B2(n6975), .A(n10005), .ZN(n6981) );
  NOR2_X1 U8751 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7996), .ZN(n6979) );
  NOR2_X1 U8752 ( .A1(n9988), .A2(n6977), .ZN(n6978) );
  AOI211_X1 U8753 ( .C1(P2_ADDR_REG_13__SCAN_IN), .C2(n9997), .A(n6979), .B(
        n6978), .ZN(n6980) );
  OAI211_X1 U8754 ( .C1(n6982), .C2(n9987), .A(n6981), .B(n6980), .ZN(P2_U3258) );
  INV_X1 U8755 ( .A(n6983), .ZN(n7011) );
  AOI22_X1 U8756 ( .A1(n9844), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n9755), .ZN(n6984) );
  OAI21_X1 U8757 ( .B1(n7011), .B2(n9763), .A(n6984), .ZN(P1_U3337) );
  NAND2_X1 U8758 ( .A1(n6985), .A2(n4278), .ZN(n6987) );
  NAND2_X1 U8759 ( .A1(n9231), .A2(n7073), .ZN(n6986) );
  NAND2_X1 U8760 ( .A1(n6987), .A2(n6986), .ZN(n6989) );
  NAND2_X1 U8761 ( .A1(n7300), .A2(n4476), .ZN(n6996) );
  INV_X1 U8762 ( .A(n7253), .ZN(n8704) );
  NAND2_X1 U8763 ( .A1(n9231), .A2(n8704), .ZN(n6995) );
  AND2_X1 U8764 ( .A1(n6996), .A2(n6995), .ZN(n7001) );
  INV_X1 U8765 ( .A(n7083), .ZN(n7081) );
  INV_X1 U8766 ( .A(n6997), .ZN(n7000) );
  INV_X1 U8767 ( .A(n6998), .ZN(n6999) );
  AOI21_X1 U8768 ( .B1(n7082), .B2(n7002), .A(n7001), .ZN(n7003) );
  AOI21_X1 U8769 ( .B1(n7081), .B2(n7082), .A(n7003), .ZN(n7010) );
  NOR2_X1 U8770 ( .A1(n8981), .A2(n9889), .ZN(n7008) );
  NOR2_X1 U8771 ( .A1(n8991), .A2(n4300), .ZN(n7005) );
  INV_X1 U8772 ( .A(n8978), .ZN(n8885) );
  OAI22_X1 U8773 ( .A1(n8885), .A2(n7297), .B1(n5105), .B2(n8980), .ZN(n7007)
         );
  AOI211_X1 U8774 ( .C1(P1_REG3_REG_1__SCAN_IN), .C2(n7088), .A(n7008), .B(
        n7007), .ZN(n7009) );
  OAI21_X1 U8775 ( .B1(n7010), .B2(n8986), .A(n7009), .ZN(P1_U3220) );
  INV_X1 U8776 ( .A(n8123), .ZN(n7695) );
  OAI222_X1 U8777 ( .A1(n8552), .A2(n10216), .B1(n8550), .B2(n7011), .C1(n7695), .C2(P2_U3152), .ZN(P2_U3342) );
  NAND2_X1 U8778 ( .A1(n7013), .A2(n7012), .ZN(n7014) );
  INV_X1 U8779 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n7040) );
  XNOR2_X1 U8780 ( .A(n6370), .B(n7375), .ZN(n8387) );
  NAND2_X1 U8781 ( .A1(n8387), .A2(n8392), .ZN(n10014) );
  INV_X1 U8782 ( .A(n10084), .ZN(n8518) );
  OAI21_X1 U8783 ( .B1(n7018), .B2(n10041), .A(n6958), .ZN(n7020) );
  NAND2_X1 U8784 ( .A1(n7018), .A2(n10041), .ZN(n7019) );
  NAND2_X1 U8785 ( .A1(n7020), .A2(n7019), .ZN(n7569) );
  NAND2_X1 U8786 ( .A1(n7569), .A2(n7021), .ZN(n7023) );
  OR2_X1 U8787 ( .A1(n6388), .A2(n5841), .ZN(n7022) );
  NAND2_X1 U8788 ( .A1(n7023), .A2(n7022), .ZN(n10012) );
  NAND2_X1 U8789 ( .A1(n10012), .A2(n7024), .ZN(n7026) );
  OR2_X1 U8790 ( .A1(n8068), .A2(n7923), .ZN(n7025) );
  NAND2_X1 U8791 ( .A1(n7026), .A2(n7025), .ZN(n7582) );
  OR2_X1 U8792 ( .A1(n8067), .A2(n10062), .ZN(n7028) );
  XNOR2_X1 U8793 ( .A(n7171), .B(n7032), .ZN(n7531) );
  NAND2_X1 U8794 ( .A1(n7029), .A2(n7030), .ZN(n7031) );
  XOR2_X1 U8795 ( .A(n7032), .B(n7031), .Z(n7035) );
  OAI22_X1 U8796 ( .A1(n8405), .A2(n5868), .B1(n7059), .B2(n8407), .ZN(n7043)
         );
  AOI21_X1 U8797 ( .B1(n7035), .B2(n10017), .A(n7043), .ZN(n7528) );
  NAND2_X1 U8798 ( .A1(n10041), .A2(n10090), .ZN(n7574) );
  INV_X1 U8799 ( .A(n7455), .ZN(n7037) );
  AOI211_X1 U8800 ( .C1(n4284), .C2(n7584), .A(n4296), .B(n7037), .ZN(n7521)
         );
  AOI21_X1 U8801 ( .B1(n10063), .B2(n4284), .A(n7521), .ZN(n7038) );
  OAI211_X1 U8802 ( .C1(n8523), .C2(n7531), .A(n7528), .B(n7038), .ZN(n7071)
         );
  NAND2_X1 U8803 ( .A1(n7071), .A2(n10283), .ZN(n7039) );
  OAI21_X1 U8804 ( .B1(n10283), .B2(n7040), .A(n7039), .ZN(P2_U3466) );
  NOR2_X1 U8805 ( .A1(n8037), .A2(n7522), .ZN(n7041) );
  AOI211_X1 U8806 ( .C1(n8005), .C2(n7043), .A(n7042), .B(n7041), .ZN(n7057)
         );
  INV_X1 U8807 ( .A(n7044), .ZN(n7045) );
  NAND2_X1 U8808 ( .A1(n7045), .A2(n7050), .ZN(n7918) );
  INV_X1 U8809 ( .A(n7918), .ZN(n7047) );
  NAND2_X1 U8810 ( .A1(n7047), .A2(n7046), .ZN(n7920) );
  XNOR2_X1 U8811 ( .A(n7049), .B(n7048), .ZN(n7189) );
  AND3_X1 U8812 ( .A1(n7920), .A2(n7050), .A3(n7189), .ZN(n7182) );
  NOR2_X1 U8813 ( .A1(n7182), .A2(n7051), .ZN(n7055) );
  OAI211_X1 U8814 ( .C1(n7055), .C2(n7054), .A(n7993), .B(n7053), .ZN(n7056)
         );
  OAI211_X1 U8815 ( .C1(n7058), .C2(n8032), .A(n7057), .B(n7056), .ZN(P2_U3229) );
  INV_X1 U8816 ( .A(n7216), .ZN(n7478) );
  OAI22_X1 U8817 ( .A1(n8405), .A2(n7059), .B1(n7882), .B2(n8407), .ZN(n7176)
         );
  NOR2_X1 U8818 ( .A1(n8037), .A2(n7475), .ZN(n7060) );
  AOI211_X1 U8819 ( .C1(n8005), .C2(n7176), .A(n7061), .B(n7060), .ZN(n7067)
         );
  AOI21_X1 U8820 ( .B1(n7063), .B2(n7062), .A(n8044), .ZN(n7065) );
  NAND2_X1 U8821 ( .A1(n7065), .A2(n7064), .ZN(n7066) );
  OAI211_X1 U8822 ( .C1(n7478), .C2(n8032), .A(n7067), .B(n7066), .ZN(P2_U3215) );
  NAND2_X1 U8823 ( .A1(n7071), .A2(n10100), .ZN(n7072) );
  OAI21_X1 U8824 ( .B1(n10100), .B2(n6733), .A(n7072), .ZN(P2_U3525) );
  INV_X1 U8825 ( .A(n7082), .ZN(n7080) );
  OR2_X1 U8826 ( .A1(n5105), .A2(n7253), .ZN(n7076) );
  NAND2_X1 U8827 ( .A1(n7282), .A2(n7073), .ZN(n7075) );
  AND2_X1 U8828 ( .A1(n7076), .A2(n7075), .ZN(n7077) );
  NAND2_X1 U8829 ( .A1(n7078), .A2(n7077), .ZN(n7152) );
  NOR3_X1 U8830 ( .A1(n7081), .A2(n7080), .A3(n7084), .ZN(n7086) );
  NAND2_X1 U8831 ( .A1(n7083), .A2(n7082), .ZN(n7085) );
  NAND2_X1 U8832 ( .A1(n7085), .A2(n7084), .ZN(n7153) );
  INV_X1 U8833 ( .A(n7153), .ZN(n7151) );
  OAI21_X1 U8834 ( .B1(n7086), .B2(n7151), .A(n8959), .ZN(n7090) );
  OAI22_X1 U8835 ( .A1(n8885), .A2(n7274), .B1(n7273), .B2(n8980), .ZN(n7087)
         );
  AOI21_X1 U8836 ( .B1(P1_REG3_REG_2__SCAN_IN), .B2(n7088), .A(n7087), .ZN(
        n7089) );
  OAI211_X1 U8837 ( .C1(n9896), .C2(n8981), .A(n7090), .B(n7089), .ZN(P1_U3235) );
  INV_X1 U8838 ( .A(n7091), .ZN(n7096) );
  OAI21_X1 U8839 ( .B1(n7094), .B2(n7093), .A(n7092), .ZN(n7095) );
  AOI21_X1 U8840 ( .B1(n7096), .B2(n7095), .A(n9989), .ZN(n7106) );
  INV_X1 U8841 ( .A(n7097), .ZN(n7098) );
  AOI211_X1 U8842 ( .C1(n7100), .C2(n7099), .A(n9987), .B(n7098), .ZN(n7105)
         );
  INV_X1 U8843 ( .A(n9997), .ZN(n8106) );
  INV_X1 U8844 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n7103) );
  NAND2_X1 U8845 ( .A1(n10003), .A2(n7101), .ZN(n7102) );
  NAND2_X1 U8846 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3152), .ZN(n7594) );
  OAI211_X1 U8847 ( .C1(n8106), .C2(n7103), .A(n7102), .B(n7594), .ZN(n7104)
         );
  OR3_X1 U8848 ( .A1(n7106), .A2(n7105), .A3(n7104), .ZN(P2_U3257) );
  INV_X1 U8849 ( .A(n7107), .ZN(n7110) );
  OAI222_X1 U8850 ( .A1(n8552), .A2(n7108), .B1(n8550), .B2(n7110), .C1(n8127), 
        .C2(P2_U3152), .ZN(P2_U3341) );
  OAI222_X1 U8851 ( .A1(P1_U3084), .A2(n9858), .B1(n9763), .B2(n7110), .C1(
        n7109), .C2(n9765), .ZN(P1_U3336) );
  XNOR2_X1 U8852 ( .A(n4290), .B(n7111), .ZN(n7115) );
  NAND2_X1 U8853 ( .A1(n7113), .A2(n7112), .ZN(n7114) );
  NAND2_X1 U8854 ( .A1(n7114), .A2(n7115), .ZN(n7321) );
  OAI21_X1 U8855 ( .B1(n7115), .B2(n7114), .A(n7321), .ZN(n7127) );
  OR2_X1 U8856 ( .A1(n7116), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n7120) );
  NAND2_X1 U8857 ( .A1(n7122), .A2(n7120), .ZN(n7118) );
  INV_X1 U8858 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n7117) );
  MUX2_X1 U8859 ( .A(P2_REG2_REG_14__SCAN_IN), .B(n7117), .S(n4290), .Z(n7119)
         );
  NAND2_X1 U8860 ( .A1(n7118), .A2(n7119), .ZN(n7325) );
  INV_X1 U8861 ( .A(n7119), .ZN(n7121) );
  NAND3_X1 U8862 ( .A1(n7122), .A2(n7121), .A3(n7120), .ZN(n7123) );
  AOI21_X1 U8863 ( .B1(n7325), .B2(n7123), .A(n9987), .ZN(n7126) );
  INV_X1 U8864 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n10157) );
  NAND2_X1 U8865 ( .A1(n10003), .A2(n4290), .ZN(n7124) );
  NAND2_X1 U8866 ( .A1(P2_U3152), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n7808) );
  OAI211_X1 U8867 ( .C1(n8106), .C2(n10157), .A(n7124), .B(n7808), .ZN(n7125)
         );
  AOI211_X1 U8868 ( .C1(n7127), .C2(n10005), .A(n7126), .B(n7125), .ZN(n7128)
         );
  INV_X1 U8869 ( .A(n7128), .ZN(P2_U3259) );
  INV_X1 U8870 ( .A(n7129), .ZN(n7130) );
  AOI21_X1 U8871 ( .B1(n7064), .B2(n7130), .A(n8044), .ZN(n7134) );
  NOR3_X1 U8872 ( .A1(n8008), .A2(n7131), .A3(n7135), .ZN(n7133) );
  OAI21_X1 U8873 ( .B1(n7134), .B2(n7133), .A(n7132), .ZN(n7139) );
  OAI22_X1 U8874 ( .A1(n8405), .A2(n7135), .B1(n7565), .B2(n8407), .ZN(n7228)
         );
  NOR2_X1 U8875 ( .A1(n8037), .A2(n7382), .ZN(n7136) );
  AOI211_X1 U8876 ( .C1(n8005), .C2(n7228), .A(n7137), .B(n7136), .ZN(n7138)
         );
  OAI211_X1 U8877 ( .C1(n7383), .C2(n8032), .A(n7139), .B(n7138), .ZN(P2_U3223) );
  INV_X1 U8878 ( .A(n7152), .ZN(n7150) );
  NAND2_X1 U8879 ( .A1(n7426), .A2(n4278), .ZN(n7141) );
  NAND2_X1 U8880 ( .A1(n9915), .A2(n8774), .ZN(n7140) );
  XNOR2_X1 U8881 ( .A(n7142), .B(n4468), .ZN(n7145) );
  NAND2_X1 U8882 ( .A1(n7426), .A2(n8774), .ZN(n7144) );
  NAND2_X1 U8883 ( .A1(n9915), .A2(n8704), .ZN(n7143) );
  AND2_X1 U8884 ( .A1(n7144), .A2(n7143), .ZN(n7146) );
  NAND2_X1 U8885 ( .A1(n7145), .A2(n7146), .ZN(n7256) );
  INV_X1 U8886 ( .A(n7145), .ZN(n7148) );
  INV_X1 U8887 ( .A(n7146), .ZN(n7147) );
  NAND2_X1 U8888 ( .A1(n7148), .A2(n7147), .ZN(n7149) );
  AND2_X1 U8889 ( .A1(n7256), .A2(n7149), .ZN(n7154) );
  NOR3_X1 U8890 ( .A1(n7151), .A2(n7150), .A3(n7154), .ZN(n7157) );
  NAND2_X1 U8891 ( .A1(n7153), .A2(n7152), .ZN(n7155) );
  INV_X1 U8892 ( .A(n7257), .ZN(n7156) );
  OAI21_X1 U8893 ( .B1(n7157), .B2(n7156), .A(n8959), .ZN(n7169) );
  NAND2_X1 U8894 ( .A1(n7158), .A2(n8988), .ZN(n7160) );
  NOR2_X1 U8895 ( .A1(n7160), .A2(n7159), .ZN(n7161) );
  NAND2_X1 U8896 ( .A1(n7162), .A2(n7161), .ZN(n7163) );
  AOI21_X1 U8897 ( .B1(n8978), .B2(n9229), .A(n7164), .ZN(n7165) );
  OAI21_X1 U8898 ( .B1(n9928), .B2(n8980), .A(n7165), .ZN(n7166) );
  AOI21_X1 U8899 ( .B1(n8984), .B2(n7167), .A(n7166), .ZN(n7168) );
  OAI211_X1 U8900 ( .C1(n9902), .C2(n8981), .A(n7169), .B(n7168), .ZN(P1_U3216) );
  NOR2_X1 U8901 ( .A1(n8066), .A2(n4284), .ZN(n7170) );
  NAND2_X1 U8902 ( .A1(n7452), .A2(n7172), .ZN(n7222) );
  INV_X1 U8903 ( .A(n7222), .ZN(n7173) );
  NOR2_X1 U8904 ( .A1(n7454), .A2(n8065), .ZN(n7218) );
  NOR2_X1 U8905 ( .A1(n7173), .A2(n7218), .ZN(n7174) );
  XNOR2_X1 U8906 ( .A(n7174), .B(n7221), .ZN(n7472) );
  XNOR2_X1 U8907 ( .A(n7175), .B(n7221), .ZN(n7177) );
  AOI21_X1 U8908 ( .B1(n7177), .B2(n10017), .A(n7176), .ZN(n7473) );
  NAND2_X1 U8909 ( .A1(n7453), .A2(n7478), .ZN(n7230) );
  OAI211_X1 U8910 ( .C1(n7453), .C2(n7478), .A(n10019), .B(n7230), .ZN(n7474)
         );
  OAI211_X1 U8911 ( .C1(n7478), .C2(n10077), .A(n7473), .B(n7474), .ZN(n7178)
         );
  AOI21_X1 U8912 ( .B1(n10086), .B2(n7472), .A(n7178), .ZN(n7181) );
  OR2_X1 U8913 ( .A1(n10100), .A2(n6827), .ZN(n7179) );
  OAI21_X1 U8914 ( .B1(n7181), .B2(n10098), .A(n7179), .ZN(P2_U3527) );
  INV_X1 U8915 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n10177) );
  NAND2_X1 U8916 ( .A1(n10281), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n7180) );
  OAI21_X1 U8917 ( .B1(n7181), .B2(n10281), .A(n7180), .ZN(P2_U3472) );
  INV_X1 U8918 ( .A(n7189), .ZN(n7184) );
  INV_X1 U8919 ( .A(n7920), .ZN(n7183) );
  AOI21_X1 U8920 ( .B1(n7184), .B2(n7183), .A(n7182), .ZN(n7195) );
  NAND2_X1 U8921 ( .A1(n8372), .A2(n8066), .ZN(n7186) );
  NAND2_X1 U8922 ( .A1(n8370), .A2(n8068), .ZN(n7185) );
  NAND2_X1 U8923 ( .A1(n7186), .A2(n7185), .ZN(n7580) );
  NAND2_X1 U8924 ( .A1(n8005), .A2(n7580), .ZN(n7188) );
  OAI211_X1 U8925 ( .C1(n8037), .C2(n7586), .A(n7188), .B(n7187), .ZN(n7193)
         );
  NOR4_X1 U8926 ( .A1(n8008), .A2(n7191), .A3(n7190), .A4(n7189), .ZN(n7192)
         );
  AOI211_X1 U8927 ( .C1(n8048), .C2(n10062), .A(n7193), .B(n7192), .ZN(n7194)
         );
  OAI21_X1 U8928 ( .B1(n7195), .B2(n8044), .A(n7194), .ZN(P2_U3232) );
  INV_X1 U8929 ( .A(n7454), .ZN(n10071) );
  INV_X1 U8930 ( .A(n8037), .ZN(n8027) );
  INV_X1 U8931 ( .A(n7196), .ZN(n7458) );
  NAND2_X1 U8932 ( .A1(n8027), .A2(n7458), .ZN(n7198) );
  OAI211_X1 U8933 ( .C1(n8032), .C2(n10071), .A(n7198), .B(n7197), .ZN(n7203)
         );
  INV_X1 U8934 ( .A(n7205), .ZN(n7200) );
  NAND3_X1 U8935 ( .A1(n8049), .A2(n7200), .A3(n7199), .ZN(n7201) );
  AOI21_X1 U8936 ( .B1(n7201), .B2(n8020), .A(n4827), .ZN(n7202) );
  AOI211_X1 U8937 ( .C1(n8018), .C2(n8064), .A(n7203), .B(n7202), .ZN(n7208)
         );
  OAI21_X1 U8938 ( .B1(n7053), .B2(n7205), .A(n7204), .ZN(n7206) );
  NAND2_X1 U8939 ( .A1(n7206), .A2(n7993), .ZN(n7207) );
  NAND2_X1 U8940 ( .A1(n7208), .A2(n7207), .ZN(P2_U3241) );
  INV_X1 U8941 ( .A(n7209), .ZN(n7211) );
  OAI222_X1 U8942 ( .A1(P1_U3084), .A2(n9418), .B1(n9763), .B2(n7211), .C1(
        n7210), .C2(n7782), .ZN(P1_U3334) );
  OAI222_X1 U8943 ( .A1(n8552), .A2(n7212), .B1(n8550), .B2(n7211), .C1(n8392), 
        .C2(P2_U3152), .ZN(P2_U3339) );
  INV_X1 U8944 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n10205) );
  INV_X1 U8945 ( .A(n7213), .ZN(n7215) );
  INV_X1 U8946 ( .A(n8137), .ZN(n8143) );
  OAI222_X1 U8947 ( .A1(n8552), .A2(n10205), .B1(n8550), .B2(n7215), .C1(
        P2_U3152), .C2(n8143), .ZN(P2_U3340) );
  OAI222_X1 U8948 ( .A1(n9279), .A2(P1_U3084), .B1(n9763), .B2(n7215), .C1(
        n7214), .C2(n7782), .ZN(P1_U3335) );
  INV_X1 U8949 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n7234) );
  NOR2_X1 U8950 ( .A1(n7216), .A2(n8064), .ZN(n7217) );
  AOI21_X1 U8951 ( .B1(n7219), .B2(n7218), .A(n7217), .ZN(n7220) );
  INV_X1 U8952 ( .A(n7223), .ZN(n7224) );
  OAI21_X1 U8953 ( .B1(n7224), .B2(n4282), .A(n7391), .ZN(n7388) );
  XNOR2_X1 U8954 ( .A(n7226), .B(n7227), .ZN(n7229) );
  AOI21_X1 U8955 ( .B1(n7229), .B2(n10017), .A(n7228), .ZN(n7378) );
  AOI21_X1 U8956 ( .B1(n7230), .B2(n7389), .A(n4296), .ZN(n7231) );
  AND2_X1 U8957 ( .A1(n7231), .A2(n7395), .ZN(n7385) );
  AOI21_X1 U8958 ( .B1(n10063), .B2(n7389), .A(n7385), .ZN(n7232) );
  OAI211_X1 U8959 ( .C1(n7388), .C2(n8523), .A(n7378), .B(n7232), .ZN(n7235)
         );
  NAND2_X1 U8960 ( .A1(n7235), .A2(n10283), .ZN(n7233) );
  OAI21_X1 U8961 ( .B1(n10283), .B2(n7234), .A(n7233), .ZN(P2_U3475) );
  NAND2_X1 U8962 ( .A1(n7235), .A2(n10100), .ZN(n7236) );
  OAI21_X1 U8963 ( .B1(n10100), .B2(n6829), .A(n7236), .ZN(P2_U3528) );
  INV_X1 U8964 ( .A(n7237), .ZN(n7245) );
  NOR2_X1 U8965 ( .A1(n7671), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n7677) );
  INV_X1 U8966 ( .A(n7677), .ZN(n7240) );
  NAND2_X1 U8967 ( .A1(n7671), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n7676) );
  NAND2_X1 U8968 ( .A1(n7240), .A2(n7676), .ZN(n7241) );
  XNOR2_X1 U8969 ( .A(n7678), .B(n7241), .ZN(n7251) );
  NAND2_X1 U8970 ( .A1(P1_U3084), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n8828) );
  OAI21_X1 U8971 ( .B1(n9859), .B2(n7242), .A(n8828), .ZN(n7249) );
  NAND2_X1 U8972 ( .A1(n7671), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n7243) );
  OAI21_X1 U8973 ( .B1(n7671), .B2(P1_REG2_REG_12__SCAN_IN), .A(n7243), .ZN(
        n7247) );
  NOR2_X1 U8974 ( .A1(n7246), .A2(n7247), .ZN(n7670) );
  AOI211_X1 U8975 ( .C1(n7247), .C2(n7246), .A(n9839), .B(n7670), .ZN(n7248)
         );
  AOI211_X1 U8976 ( .C1(n9810), .C2(P1_ADDR_REG_12__SCAN_IN), .A(n7249), .B(
        n7248), .ZN(n7250) );
  OAI21_X1 U8977 ( .B1(n9281), .B2(n7251), .A(n7250), .ZN(P1_U3253) );
  OAI22_X1 U8978 ( .A1(n9928), .A2(n8711), .B1(n7442), .B2(n4463), .ZN(n7252)
         );
  XNOR2_X1 U8979 ( .A(n7252), .B(n4468), .ZN(n7604) );
  OR2_X1 U8980 ( .A1(n9928), .A2(n8775), .ZN(n7255) );
  NAND2_X1 U8981 ( .A1(n9912), .A2(n8774), .ZN(n7254) );
  NAND2_X1 U8982 ( .A1(n7255), .A2(n7254), .ZN(n7602) );
  XNOR2_X1 U8983 ( .A(n7604), .B(n7602), .ZN(n7259) );
  NAND2_X1 U8984 ( .A1(n7257), .A2(n7256), .ZN(n7258) );
  OAI21_X1 U8985 ( .B1(n7259), .B2(n7258), .A(n7606), .ZN(n7266) );
  NOR2_X1 U8986 ( .A1(n8981), .A2(n7442), .ZN(n7265) );
  AOI21_X1 U8987 ( .B1(n8978), .B2(n9915), .A(n7260), .ZN(n7263) );
  NAND2_X1 U8988 ( .A1(n8984), .A2(n7440), .ZN(n7262) );
  NAND2_X1 U8989 ( .A1(n8894), .A2(n9227), .ZN(n7261) );
  NAND3_X1 U8990 ( .A1(n7263), .A2(n7262), .A3(n7261), .ZN(n7264) );
  AOI211_X1 U8991 ( .C1(n7266), .C2(n8959), .A(n7265), .B(n7264), .ZN(n7267)
         );
  INV_X1 U8992 ( .A(n7267), .ZN(P1_U3228) );
  INV_X1 U8993 ( .A(n7268), .ZN(n7289) );
  OAI222_X1 U8994 ( .A1(n9120), .A2(P1_U3084), .B1(n9763), .B2(n7289), .C1(
        n7269), .C2(n7782), .ZN(P1_U3333) );
  XNOR2_X1 U8995 ( .A(n9231), .B(n7300), .ZN(n9094) );
  OAI22_X1 U8996 ( .A1(n9094), .A2(n7291), .B1(n9231), .B2(n7300), .ZN(n7270)
         );
  XNOR2_X1 U8997 ( .A(n7270), .B(n9093), .ZN(n9900) );
  INV_X1 U8998 ( .A(n9900), .ZN(n7286) );
  INV_X1 U8999 ( .A(n7271), .ZN(n7272) );
  NAND2_X1 U9000 ( .A1(n9541), .A2(n7272), .ZN(n7285) );
  INV_X1 U9001 ( .A(n9887), .ZN(n9923) );
  OAI22_X1 U9002 ( .A1(n7274), .A2(n9943), .B1(n7273), .B2(n9518), .ZN(n7279)
         );
  NAND2_X1 U9003 ( .A1(n7275), .A2(n9093), .ZN(n7276) );
  AOI21_X1 U9004 ( .B1(n7277), .B2(n7276), .A(n9515), .ZN(n7278) );
  AOI211_X1 U9005 ( .C1(n9923), .C2(n9900), .A(n7279), .B(n7278), .ZN(n9897)
         );
  MUX2_X1 U9006 ( .A(n6614), .B(n9897), .S(n9541), .Z(n7284) );
  OAI21_X1 U9007 ( .B1(n7300), .B2(n7292), .A(n7282), .ZN(n7280) );
  NAND3_X1 U9008 ( .A1(n7280), .A2(n9569), .A3(n7427), .ZN(n9895) );
  INV_X1 U9009 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n9235) );
  OAI22_X1 U9010 ( .A1(n9895), .A2(n9580), .B1(n9235), .B2(n9538), .ZN(n7281)
         );
  AOI21_X1 U9011 ( .B1(n9578), .B2(n7282), .A(n7281), .ZN(n7283) );
  OAI211_X1 U9012 ( .C1(n7286), .C2(n7285), .A(n7284), .B(n7283), .ZN(P1_U3289) );
  INV_X1 U9013 ( .A(n7287), .ZN(n7367) );
  OAI222_X1 U9014 ( .A1(n5662), .A2(P1_U3084), .B1(n9763), .B2(n7367), .C1(
        n7288), .C2(n9765), .ZN(P1_U3332) );
  OAI222_X1 U9015 ( .A1(n8552), .A2(n7290), .B1(P2_U3152), .B2(n4301), .C1(
        n8550), .C2(n7289), .ZN(P2_U3338) );
  XNOR2_X1 U9016 ( .A(n9094), .B(n7291), .ZN(n9885) );
  XNOR2_X1 U9017 ( .A(n9889), .B(n7292), .ZN(n7293) );
  NAND2_X1 U9018 ( .A1(n7293), .A2(n9569), .ZN(n9888) );
  OAI22_X1 U9019 ( .A1(n9888), .A2(n9119), .B1(n9538), .B2(n7294), .ZN(n7298)
         );
  XNOR2_X1 U9020 ( .A(n9094), .B(n7295), .ZN(n7296) );
  OAI222_X1 U9021 ( .A1(n9518), .A2(n5105), .B1(n9943), .B2(n7297), .C1(n7296), 
        .C2(n9515), .ZN(n9891) );
  AOI211_X1 U9022 ( .C1(n9885), .C2(n7299), .A(n7298), .B(n9891), .ZN(n7302)
         );
  AOI22_X1 U9023 ( .A1(n9578), .A2(n7300), .B1(n9877), .B2(
        P1_REG2_REG_1__SCAN_IN), .ZN(n7301) );
  OAI21_X1 U9024 ( .B1(n7302), .B2(n9877), .A(n7301), .ZN(P1_U3290) );
  INV_X1 U9025 ( .A(n7304), .ZN(n7306) );
  AOI21_X1 U9026 ( .B1(n7303), .B2(n7306), .A(n7305), .ZN(n7307) );
  XNOR2_X1 U9027 ( .A(n7307), .B(n9098), .ZN(n9941) );
  INV_X1 U9028 ( .A(n7308), .ZN(n7311) );
  AOI21_X1 U9029 ( .B1(n9136), .B2(n9134), .A(n7309), .ZN(n7310) );
  OAI21_X1 U9030 ( .B1(n7311), .B2(n7310), .A(n9563), .ZN(n7312) );
  OAI21_X1 U9031 ( .B1(n8884), .B2(n9518), .A(n7312), .ZN(n9948) );
  OAI21_X1 U9032 ( .B1(n7419), .B2(n9942), .A(n9569), .ZN(n7313) );
  NOR2_X1 U9033 ( .A1(n7313), .A2(n7339), .ZN(n9946) );
  NAND2_X1 U9034 ( .A1(n9946), .A2(n9528), .ZN(n7318) );
  INV_X1 U9035 ( .A(n7653), .ZN(n7314) );
  OAI22_X1 U9036 ( .A1(n9541), .A2(n7315), .B1(n7314), .B2(n9538), .ZN(n7316)
         );
  AOI21_X1 U9037 ( .B1(n9544), .B2(n9226), .A(n7316), .ZN(n7317) );
  OAI211_X1 U9038 ( .C1(n9942), .C2(n9526), .A(n7318), .B(n7317), .ZN(n7319)
         );
  AOI21_X1 U9039 ( .B1(n9948), .B2(n9541), .A(n7319), .ZN(n7320) );
  OAI21_X1 U9040 ( .B1(n9941), .B2(n9513), .A(n7320), .ZN(P1_U3284) );
  XOR2_X1 U9041 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n7694), .Z(n7335) );
  OR2_X1 U9042 ( .A1(n4290), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n7324) );
  NAND2_X1 U9043 ( .A1(n7325), .A2(n7324), .ZN(n7326) );
  NAND2_X1 U9044 ( .A1(n7326), .A2(n7692), .ZN(n7689) );
  OR2_X1 U9045 ( .A1(n7326), .A2(n7692), .ZN(n7327) );
  AND2_X1 U9046 ( .A1(n7689), .A2(n7327), .ZN(n7329) );
  INV_X1 U9047 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n7328) );
  NAND2_X1 U9048 ( .A1(n7329), .A2(n7328), .ZN(n7690) );
  OAI21_X1 U9049 ( .B1(n7329), .B2(n7328), .A(n7690), .ZN(n7333) );
  AND2_X1 U9050 ( .A1(P2_U3152), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n7330) );
  AOI21_X1 U9051 ( .B1(n9997), .B2(P2_ADDR_REG_15__SCAN_IN), .A(n7330), .ZN(
        n7331) );
  OAI21_X1 U9052 ( .B1(n9988), .B2(n7692), .A(n7331), .ZN(n7332) );
  AOI21_X1 U9053 ( .B1(n7333), .B2(n9999), .A(n7332), .ZN(n7334) );
  OAI21_X1 U9054 ( .B1(n7335), .B2(n9989), .A(n7334), .ZN(P2_U3260) );
  OAI211_X1 U9055 ( .C1(n4984), .C2(n7336), .A(n9563), .B(n7484), .ZN(n7338)
         );
  AOI22_X1 U9056 ( .A1(n9562), .A2(n9223), .B1(n9225), .B2(n9914), .ZN(n7337)
         );
  NAND2_X1 U9057 ( .A1(n7338), .A2(n7337), .ZN(n9954) );
  NAND2_X1 U9058 ( .A1(n7339), .A2(n9953), .ZN(n7487) );
  OAI211_X1 U9059 ( .C1(n7339), .C2(n9953), .A(n9569), .B(n7487), .ZN(n9952)
         );
  AOI22_X1 U9060 ( .A1(n9877), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n8809), .B2(
        n9874), .ZN(n7341) );
  NAND2_X1 U9061 ( .A1(n9578), .A2(n8559), .ZN(n7340) );
  OAI211_X1 U9062 ( .C1(n9952), .C2(n9580), .A(n7341), .B(n7340), .ZN(n7347)
         );
  AOI21_X1 U9063 ( .B1(n7303), .B2(n7343), .A(n7342), .ZN(n7344) );
  NOR2_X1 U9064 ( .A1(n7344), .A2(n9099), .ZN(n9951) );
  NAND2_X1 U9065 ( .A1(n7344), .A2(n9099), .ZN(n9956) );
  INV_X1 U9066 ( .A(n9956), .ZN(n7345) );
  NOR3_X1 U9067 ( .A1(n9951), .A2(n7345), .A3(n9513), .ZN(n7346) );
  AOI211_X1 U9068 ( .C1(n9541), .C2(n9954), .A(n7347), .B(n7346), .ZN(n7348)
         );
  INV_X1 U9069 ( .A(n7348), .ZN(P1_U3283) );
  INV_X1 U9070 ( .A(n7349), .ZN(n7896) );
  NAND2_X1 U9071 ( .A1(n7353), .A2(n7352), .ZN(n7435) );
  NAND2_X1 U9072 ( .A1(n7435), .A2(n7354), .ZN(n7413) );
  NAND2_X1 U9073 ( .A1(n7413), .A2(n7411), .ZN(n7355) );
  XNOR2_X1 U9074 ( .A(n7355), .B(n9095), .ZN(n7356) );
  OAI22_X1 U9075 ( .A1(n7356), .A2(n9515), .B1(n9944), .B2(n9518), .ZN(n9932)
         );
  INV_X1 U9076 ( .A(n9932), .ZN(n7366) );
  INV_X1 U9077 ( .A(n7420), .ZN(n7357) );
  AOI211_X1 U9078 ( .C1(n7599), .C2(n7438), .A(n9535), .B(n7357), .ZN(n9930)
         );
  INV_X1 U9079 ( .A(n7612), .ZN(n7358) );
  OAI22_X1 U9080 ( .A1(n9541), .A2(n7359), .B1(n7358), .B2(n9538), .ZN(n7360)
         );
  AOI21_X1 U9081 ( .B1(n9578), .B2(n7599), .A(n7360), .ZN(n7361) );
  OAI21_X1 U9082 ( .B1(n9928), .B2(n9576), .A(n7361), .ZN(n7364) );
  INV_X1 U9083 ( .A(n9095), .ZN(n7362) );
  NOR2_X1 U9084 ( .A1(n5191), .A2(n7362), .ZN(n9926) );
  NAND2_X1 U9085 ( .A1(n5191), .A2(n7362), .ZN(n7417) );
  INV_X1 U9086 ( .A(n7417), .ZN(n9925) );
  NOR3_X1 U9087 ( .A1(n9926), .A2(n9925), .A3(n9513), .ZN(n7363) );
  AOI211_X1 U9088 ( .C1(n9528), .C2(n9930), .A(n7364), .B(n7363), .ZN(n7365)
         );
  OAI21_X1 U9089 ( .B1(n9877), .B2(n7366), .A(n7365), .ZN(P1_U3286) );
  OAI222_X1 U9090 ( .A1(n8552), .A2(n7369), .B1(P2_U3152), .B2(n7368), .C1(
        n8550), .C2(n7367), .ZN(P2_U3337) );
  NOR2_X1 U9091 ( .A1(n7371), .A2(n7370), .ZN(n7372) );
  INV_X1 U9092 ( .A(n7375), .ZN(n7376) );
  NAND2_X1 U9093 ( .A1(n7376), .A2(n4291), .ZN(n7542) );
  AND2_X1 U9094 ( .A1(n10014), .A2(n7542), .ZN(n7377) );
  MUX2_X1 U9095 ( .A(n7379), .B(n7378), .S(n8417), .Z(n7387) );
  OR2_X1 U9096 ( .A1(n7380), .A2(n4291), .ZN(n10023) );
  INV_X1 U9097 ( .A(n10023), .ZN(n8377) );
  OAI22_X1 U9098 ( .A1(n10024), .A2(n7383), .B1(n10022), .B2(n7382), .ZN(n7384) );
  AOI21_X1 U9099 ( .B1(n8377), .B2(n7385), .A(n7384), .ZN(n7386) );
  OAI211_X1 U9100 ( .C1(n8379), .C2(n7388), .A(n7387), .B(n7386), .ZN(P2_U3288) );
  NAND2_X1 U9101 ( .A1(n7389), .A2(n8063), .ZN(n7390) );
  XOR2_X1 U9102 ( .A(n7540), .B(n7539), .Z(n7467) );
  XNOR2_X1 U9103 ( .A(n7392), .B(n7539), .ZN(n7393) );
  AOI222_X1 U9104 ( .A1(n10017), .A2(n7393), .B1(n8061), .B2(n8372), .C1(n8063), .C2(n8370), .ZN(n7466) );
  MUX2_X1 U9105 ( .A(n7394), .B(n7466), .S(n8417), .Z(n7398) );
  AOI21_X1 U9106 ( .B1(n7885), .B2(n7395), .A(n7551), .ZN(n7464) );
  OAI22_X1 U9107 ( .A1(n10024), .A2(n4794), .B1(n10022), .B2(n7880), .ZN(n7396) );
  AOI21_X1 U9108 ( .B1(n7464), .B2(n8420), .A(n7396), .ZN(n7397) );
  OAI211_X1 U9109 ( .C1(n8379), .C2(n7467), .A(n7398), .B(n7397), .ZN(P2_U3287) );
  INV_X1 U9110 ( .A(n7400), .ZN(n7401) );
  AOI21_X1 U9111 ( .B1(n7399), .B2(n7401), .A(n8044), .ZN(n7405) );
  NOR3_X1 U9112 ( .A1(n8008), .A2(n7402), .A3(n7881), .ZN(n7404) );
  OAI21_X1 U9113 ( .B1(n7405), .B2(n7404), .A(n7403), .ZN(n7410) );
  OAI22_X1 U9114 ( .A1(n8037), .A2(n7715), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7406), .ZN(n7408) );
  OAI22_X1 U9115 ( .A1(n8020), .A2(n7881), .B1(n7735), .B2(n8041), .ZN(n7407)
         );
  AOI211_X1 U9116 ( .C1(n8048), .C2(n7737), .A(n7408), .B(n7407), .ZN(n7409)
         );
  NAND2_X1 U9117 ( .A1(n7410), .A2(n7409), .ZN(P2_U3238) );
  XNOR2_X1 U9118 ( .A(n9013), .B(n9005), .ZN(n7415) );
  AOI222_X1 U9119 ( .A1(n9563), .A2(n7415), .B1(n9227), .B2(n9914), .C1(n9225), 
        .C2(n9562), .ZN(n9939) );
  NAND2_X1 U9120 ( .A1(n7417), .A2(n7416), .ZN(n7418) );
  INV_X1 U9121 ( .A(n9005), .ZN(n9096) );
  XNOR2_X1 U9122 ( .A(n7418), .B(n9096), .ZN(n9937) );
  AOI211_X1 U9123 ( .C1(n8944), .C2(n7420), .A(n9535), .B(n7419), .ZN(n9935)
         );
  NAND2_X1 U9124 ( .A1(n9935), .A2(n9528), .ZN(n7422) );
  AOI22_X1 U9125 ( .A1(n9877), .A2(P1_REG2_REG_6__SCAN_IN), .B1(n8955), .B2(
        n9874), .ZN(n7421) );
  OAI211_X1 U9126 ( .C1(n7621), .C2(n9526), .A(n7422), .B(n7421), .ZN(n7423)
         );
  AOI21_X1 U9127 ( .B1(n9582), .B2(n9937), .A(n7423), .ZN(n7424) );
  OAI21_X1 U9128 ( .B1(n9939), .B2(n9877), .A(n7424), .ZN(P1_U3285) );
  AOI22_X1 U9129 ( .A1(n7425), .A2(n9563), .B1(n9562), .B2(n9228), .ZN(n9909)
         );
  NAND2_X1 U9130 ( .A1(n7427), .A2(n7426), .ZN(n7428) );
  NAND2_X1 U9131 ( .A1(n7428), .A2(n9569), .ZN(n7429) );
  NOR2_X1 U9132 ( .A1(n7439), .A2(n7429), .ZN(n9904) );
  OAI22_X1 U9133 ( .A1(n9541), .A2(n6613), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        n9538), .ZN(n7431) );
  OAI22_X1 U9134 ( .A1(n9576), .A2(n5105), .B1(n9902), .B2(n9526), .ZN(n7430)
         );
  AOI211_X1 U9135 ( .C1(n9528), .C2(n9904), .A(n7431), .B(n7430), .ZN(n7434)
         );
  XNOR2_X1 U9136 ( .A(n7432), .B(n9090), .ZN(n9905) );
  NAND2_X1 U9137 ( .A1(n9905), .A2(n9582), .ZN(n7433) );
  OAI211_X1 U9138 ( .C1(n9909), .C2(n9877), .A(n7434), .B(n7433), .ZN(P1_U3288) );
  XNOR2_X1 U9139 ( .A(n7435), .B(n9091), .ZN(n7436) );
  AOI22_X1 U9140 ( .A1(n7436), .A2(n9563), .B1(n9562), .B2(n9227), .ZN(n9919)
         );
  XNOR2_X1 U9141 ( .A(n7437), .B(n9091), .ZN(n9922) );
  OAI211_X1 U9142 ( .C1(n7439), .C2(n7442), .A(n9569), .B(n7438), .ZN(n9916)
         );
  AOI22_X1 U9143 ( .A1(n9877), .A2(P1_REG2_REG_4__SCAN_IN), .B1(n7440), .B2(
        n9874), .ZN(n7441) );
  OAI21_X1 U9144 ( .B1(n7442), .B2(n9526), .A(n7441), .ZN(n7443) );
  AOI21_X1 U9145 ( .B1(n9544), .B2(n9915), .A(n7443), .ZN(n7444) );
  OAI21_X1 U9146 ( .B1(n9580), .B2(n9916), .A(n7444), .ZN(n7445) );
  AOI21_X1 U9147 ( .B1(n9582), .B2(n9922), .A(n7445), .ZN(n7446) );
  OAI21_X1 U9148 ( .B1(n9919), .B2(n9877), .A(n7446), .ZN(P1_U3287) );
  XNOR2_X1 U9149 ( .A(n7447), .B(n7451), .ZN(n7448) );
  NAND2_X1 U9150 ( .A1(n7448), .A2(n10017), .ZN(n7450) );
  AOI22_X1 U9151 ( .A1(n8064), .A2(n8372), .B1(n8370), .B2(n8066), .ZN(n7449)
         );
  NAND2_X1 U9152 ( .A1(n7450), .A2(n7449), .ZN(n10073) );
  INV_X1 U9153 ( .A(n10073), .ZN(n7463) );
  OAI21_X1 U9154 ( .B1(n7452), .B2(n7172), .A(n7222), .ZN(n10075) );
  INV_X1 U9155 ( .A(n8379), .ZN(n8208) );
  NOR2_X1 U9156 ( .A1(n10024), .A2(n10071), .ZN(n7461) );
  INV_X1 U9157 ( .A(n7453), .ZN(n7457) );
  NAND2_X1 U9158 ( .A1(n7455), .A2(n7454), .ZN(n7456) );
  NAND2_X1 U9159 ( .A1(n7457), .A2(n7456), .ZN(n10072) );
  INV_X1 U9160 ( .A(n10022), .ZN(n8363) );
  AOI22_X1 U9161 ( .A1(n4281), .A2(P2_REG2_REG_6__SCAN_IN), .B1(n7458), .B2(
        n8363), .ZN(n7459) );
  OAI21_X1 U9162 ( .B1(n8192), .B2(n10072), .A(n7459), .ZN(n7460) );
  AOI211_X1 U9163 ( .C1(n10075), .C2(n8208), .A(n7461), .B(n7460), .ZN(n7462)
         );
  OAI21_X1 U9164 ( .B1(n4281), .B2(n7463), .A(n7462), .ZN(P2_U3290) );
  INV_X1 U9165 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n7469) );
  AOI22_X1 U9166 ( .A1(n7464), .A2(n10019), .B1(n10063), .B2(n7885), .ZN(n7465) );
  OAI211_X1 U9167 ( .C1(n8523), .C2(n7467), .A(n7466), .B(n7465), .ZN(n7470)
         );
  NAND2_X1 U9168 ( .A1(n7470), .A2(n10283), .ZN(n7468) );
  OAI21_X1 U9169 ( .B1(n10283), .B2(n7469), .A(n7468), .ZN(P2_U3478) );
  NAND2_X1 U9170 ( .A1(n7470), .A2(n10100), .ZN(n7471) );
  OAI21_X1 U9171 ( .B1(n10100), .B2(n5923), .A(n7471), .ZN(P2_U3529) );
  INV_X1 U9172 ( .A(n7472), .ZN(n7483) );
  INV_X1 U9173 ( .A(n7473), .ZN(n7481) );
  NOR2_X1 U9174 ( .A1(n10023), .A2(n7474), .ZN(n7480) );
  NOR2_X1 U9175 ( .A1(n10022), .A2(n7475), .ZN(n7476) );
  AOI21_X1 U9176 ( .B1(n4281), .B2(P2_REG2_REG_7__SCAN_IN), .A(n7476), .ZN(
        n7477) );
  OAI21_X1 U9177 ( .B1(n10024), .B2(n7478), .A(n7477), .ZN(n7479) );
  AOI211_X1 U9178 ( .C1(n7481), .C2(n8417), .A(n7480), .B(n7479), .ZN(n7482)
         );
  OAI21_X1 U9179 ( .B1(n7483), .B2(n8379), .A(n7482), .ZN(P2_U3289) );
  NAND2_X1 U9180 ( .A1(n7484), .A2(n9014), .ZN(n7494) );
  NAND2_X1 U9181 ( .A1(n9010), .A2(n7492), .ZN(n9100) );
  XNOR2_X1 U9182 ( .A(n7494), .B(n9100), .ZN(n7485) );
  AOI222_X1 U9183 ( .A1(n9563), .A2(n7485), .B1(n9224), .B2(n9914), .C1(n9222), 
        .C2(n9562), .ZN(n9963) );
  XOR2_X1 U9184 ( .A(n7486), .B(n9100), .Z(n9967) );
  AOI211_X1 U9185 ( .C1(n8566), .C2(n7487), .A(n9535), .B(n4394), .ZN(n9959)
         );
  NAND2_X1 U9186 ( .A1(n9959), .A2(n9528), .ZN(n7489) );
  AOI22_X1 U9187 ( .A1(n9877), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n8887), .B2(
        n9874), .ZN(n7488) );
  OAI211_X1 U9188 ( .C1(n9962), .C2(n9526), .A(n7489), .B(n7488), .ZN(n7490)
         );
  AOI21_X1 U9189 ( .B1(n9582), .B2(n9967), .A(n7490), .ZN(n7491) );
  OAI21_X1 U9190 ( .B1(n9963), .B2(n9877), .A(n7491), .ZN(P1_U3282) );
  INV_X1 U9191 ( .A(n9010), .ZN(n7493) );
  OAI21_X1 U9192 ( .B1(n7494), .B2(n7493), .A(n7492), .ZN(n7495) );
  XNOR2_X1 U9193 ( .A(n7495), .B(n9101), .ZN(n7496) );
  OAI22_X1 U9194 ( .A1(n7496), .A2(n9515), .B1(n9575), .B2(n9518), .ZN(n7758)
         );
  INV_X1 U9195 ( .A(n7758), .ZN(n7504) );
  OAI21_X1 U9196 ( .B1(n7498), .B2(n9101), .A(n7497), .ZN(n7760) );
  OAI211_X1 U9197 ( .C1(n4394), .C2(n4952), .A(n9569), .B(n7657), .ZN(n7757)
         );
  AOI22_X1 U9198 ( .A1(n9877), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n8759), .B2(
        n9874), .ZN(n7499) );
  OAI21_X1 U9199 ( .B1(n9576), .B2(n8806), .A(n7499), .ZN(n7500) );
  AOI21_X1 U9200 ( .B1(n9578), .B2(n8580), .A(n7500), .ZN(n7501) );
  OAI21_X1 U9201 ( .B1(n7757), .B2(n9580), .A(n7501), .ZN(n7502) );
  AOI21_X1 U9202 ( .B1(n9582), .B2(n7760), .A(n7502), .ZN(n7503) );
  OAI21_X1 U9203 ( .B1(n7504), .B2(n9877), .A(n7503), .ZN(P1_U3281) );
  NAND2_X1 U9204 ( .A1(n8056), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n7505) );
  OAI21_X1 U9205 ( .B1(n8202), .B2(n8056), .A(n7505), .ZN(P2_U3581) );
  INV_X1 U9206 ( .A(n7506), .ZN(n7559) );
  AOI21_X1 U9207 ( .B1(P1_DATAO_REG_23__SCAN_IN), .B2(n7508), .A(n7507), .ZN(
        n7509) );
  OAI21_X1 U9208 ( .B1(n7559), .B2(n8550), .A(n7509), .ZN(P2_U3335) );
  XNOR2_X1 U9209 ( .A(n7018), .B(n7514), .ZN(n10039) );
  INV_X1 U9210 ( .A(n10041), .ZN(n7513) );
  OAI21_X1 U9211 ( .B1(n10090), .B2(n10041), .A(n7574), .ZN(n7510) );
  OR2_X1 U9212 ( .A1(n4296), .A2(n7510), .ZN(n10040) );
  OAI22_X1 U9213 ( .A1(n10023), .A2(n10040), .B1(n7511), .B2(n10022), .ZN(
        n7512) );
  AOI21_X1 U9214 ( .B1(n8396), .B2(n7513), .A(n7512), .ZN(n7520) );
  XOR2_X1 U9215 ( .A(n7515), .B(n7514), .Z(n7517) );
  AOI21_X1 U9216 ( .B1(n7517), .B2(n10017), .A(n7516), .ZN(n10042) );
  MUX2_X1 U9217 ( .A(n10042), .B(n7518), .S(n4281), .Z(n7519) );
  OAI211_X1 U9218 ( .C1(n10039), .C2(n8379), .A(n7520), .B(n7519), .ZN(
        P2_U3295) );
  NOR2_X1 U9219 ( .A1(n4281), .A2(n4291), .ZN(n8260) );
  INV_X1 U9220 ( .A(n8260), .ZN(n7524) );
  INV_X1 U9221 ( .A(n7521), .ZN(n7523) );
  OAI22_X1 U9222 ( .A1(n7524), .A2(n7523), .B1(n7522), .B2(n10022), .ZN(n7525)
         );
  AOI21_X1 U9223 ( .B1(n8396), .B2(n4284), .A(n7525), .ZN(n7530) );
  MUX2_X1 U9224 ( .A(n7528), .B(n7527), .S(n4281), .Z(n7529) );
  OAI211_X1 U9225 ( .C1(n8379), .C2(n7531), .A(n7530), .B(n7529), .ZN(P2_U3291) );
  INV_X1 U9226 ( .A(n10085), .ZN(n7538) );
  NAND2_X1 U9227 ( .A1(n10085), .A2(n10017), .ZN(n7533) );
  OR2_X1 U9228 ( .A1(n8407), .A2(n6958), .ZN(n7532) );
  AND2_X1 U9229 ( .A1(n7533), .A2(n7532), .ZN(n10088) );
  OAI22_X1 U9230 ( .A1(n4281), .A2(n10088), .B1(n7534), .B2(n10022), .ZN(n7535) );
  AOI21_X1 U9231 ( .B1(P2_REG2_REG_0__SCAN_IN), .B2(n4281), .A(n7535), .ZN(
        n7537) );
  OAI21_X1 U9232 ( .B1(n8396), .B2(n8420), .A(n7861), .ZN(n7536) );
  OAI211_X1 U9233 ( .C1(n7538), .C2(n8379), .A(n7537), .B(n7536), .ZN(P2_U3296) );
  INV_X1 U9234 ( .A(n7736), .ZN(n7543) );
  NOR2_X1 U9235 ( .A1(n7741), .A2(n7543), .ZN(n7705) );
  AND2_X1 U9236 ( .A1(n7741), .A2(n7543), .ZN(n7541) );
  NOR2_X1 U9237 ( .A1(n4281), .A2(n7542), .ZN(n7754) );
  INV_X1 U9238 ( .A(n7754), .ZN(n10025) );
  INV_X1 U9239 ( .A(n10014), .ZN(n8401) );
  NAND2_X1 U9240 ( .A1(n7544), .A2(n7543), .ZN(n7840) );
  NAND3_X1 U9241 ( .A1(n7546), .A2(n7545), .A3(n7736), .ZN(n7547) );
  AOI21_X1 U9242 ( .B1(n7840), .B2(n7547), .A(n8305), .ZN(n7549) );
  OAI22_X1 U9243 ( .A1(n8405), .A2(n7565), .B1(n7846), .B2(n8407), .ZN(n7548)
         );
  AOI211_X1 U9244 ( .C1(n10083), .C2(n8401), .A(n7549), .B(n7548), .ZN(n10080)
         );
  MUX2_X1 U9245 ( .A(n7550), .B(n10080), .S(n8417), .Z(n7556) );
  INV_X1 U9246 ( .A(n7704), .ZN(n10078) );
  NOR2_X1 U9247 ( .A1(n7551), .A2(n10078), .ZN(n7552) );
  OR2_X1 U9248 ( .A1(n7712), .A2(n7552), .ZN(n10079) );
  INV_X1 U9249 ( .A(n10079), .ZN(n7554) );
  OAI22_X1 U9250 ( .A1(n10024), .A2(n10078), .B1(n10022), .B2(n7564), .ZN(
        n7553) );
  AOI21_X1 U9251 ( .B1(n7554), .B2(n8420), .A(n7553), .ZN(n7555) );
  OAI211_X1 U9252 ( .C1(n7557), .C2(n10025), .A(n7556), .B(n7555), .ZN(
        P2_U3286) );
  OR2_X1 U9253 ( .A1(n8988), .A2(P1_U3084), .ZN(n9203) );
  NAND2_X1 U9254 ( .A1(n9755), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n7558) );
  OAI211_X1 U9255 ( .C1(n7559), .C2(n9763), .A(n9203), .B(n7558), .ZN(P1_U3330) );
  INV_X1 U9256 ( .A(n7399), .ZN(n7561) );
  AOI211_X1 U9257 ( .C1(n7562), .C2(n7560), .A(n8044), .B(n7561), .ZN(n7568)
         );
  NAND2_X1 U9258 ( .A1(n8018), .A2(n8060), .ZN(n7563) );
  NAND2_X1 U9259 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3152), .ZN(n8104) );
  OAI211_X1 U9260 ( .C1(n8037), .C2(n7564), .A(n7563), .B(n8104), .ZN(n7567)
         );
  OAI22_X1 U9261 ( .A1(n8020), .A2(n7565), .B1(n10078), .B2(n8032), .ZN(n7566)
         );
  OR3_X1 U9262 ( .A1(n7568), .A2(n7567), .A3(n7566), .ZN(P2_U3219) );
  XNOR2_X1 U9263 ( .A(n7021), .B(n7569), .ZN(n10052) );
  AOI22_X1 U9264 ( .A1(n8208), .A2(n10052), .B1(n8396), .B2(n5841), .ZN(n7577)
         );
  XNOR2_X1 U9265 ( .A(n7570), .B(n7571), .ZN(n7573) );
  AOI21_X1 U9266 ( .B1(n7573), .B2(n10017), .A(n7572), .ZN(n10049) );
  OAI21_X1 U9267 ( .B1(n6781), .B2(n10022), .A(n10049), .ZN(n7575) );
  AOI22_X1 U9268 ( .A1(n8417), .A2(n7575), .B1(n8377), .B2(n10047), .ZN(n7576)
         );
  OAI211_X1 U9269 ( .C1(n6741), .C2(n8417), .A(n7577), .B(n7576), .ZN(P2_U3294) );
  INV_X1 U9270 ( .A(n7583), .ZN(n7579) );
  XNOR2_X1 U9271 ( .A(n7578), .B(n7579), .ZN(n7581) );
  AOI21_X1 U9272 ( .B1(n7581), .B2(n10017), .A(n7580), .ZN(n10069) );
  XNOR2_X1 U9273 ( .A(n7582), .B(n7583), .ZN(n10066) );
  AOI22_X1 U9274 ( .A1(n8208), .A2(n10066), .B1(n8396), .B2(n10062), .ZN(n7589) );
  AOI21_X1 U9275 ( .B1(n10020), .B2(n10062), .A(n4296), .ZN(n7585) );
  NAND2_X1 U9276 ( .A1(n7585), .A2(n7584), .ZN(n10065) );
  OAI22_X1 U9277 ( .A1(n10023), .A2(n10065), .B1(n7586), .B2(n10022), .ZN(
        n7587) );
  AOI21_X1 U9278 ( .B1(n4281), .B2(P2_REG2_REG_4__SCAN_IN), .A(n7587), .ZN(
        n7588) );
  OAI211_X1 U9279 ( .C1(n4281), .C2(n10069), .A(n7589), .B(n7588), .ZN(
        P2_U3292) );
  NAND2_X1 U9280 ( .A1(n7591), .A2(n7590), .ZN(n7593) );
  XOR2_X1 U9281 ( .A(n7593), .B(n7592), .Z(n7598) );
  OAI21_X1 U9282 ( .B1(n8037), .B2(n7853), .A(n7594), .ZN(n7596) );
  OAI22_X1 U9283 ( .A1(n8020), .A2(n7846), .B1(n4795), .B2(n8032), .ZN(n7595)
         );
  AOI211_X1 U9284 ( .C1(n8018), .C2(n8058), .A(n7596), .B(n7595), .ZN(n7597)
         );
  OAI21_X1 U9285 ( .B1(n7598), .B2(n8044), .A(n7597), .ZN(P2_U3226) );
  OR2_X1 U9286 ( .A1(n7607), .A2(n8775), .ZN(n7601) );
  NAND2_X1 U9287 ( .A1(n7599), .A2(n8774), .ZN(n7600) );
  AND2_X1 U9288 ( .A1(n7601), .A2(n7600), .ZN(n7630) );
  INV_X1 U9289 ( .A(n7602), .ZN(n7603) );
  NAND2_X1 U9290 ( .A1(n7604), .A2(n7603), .ZN(n7605) );
  OAI22_X1 U9291 ( .A1(n7607), .A2(n8711), .B1(n9927), .B2(n4463), .ZN(n7608)
         );
  XNOR2_X1 U9292 ( .A(n7608), .B(n4468), .ZN(n7620) );
  INV_X1 U9293 ( .A(n7620), .ZN(n7632) );
  NOR2_X1 U9294 ( .A1(n7609), .A2(n7632), .ZN(n8945) );
  AOI21_X1 U9295 ( .B1(n7609), .B2(n7632), .A(n8945), .ZN(n7610) );
  NAND2_X1 U9296 ( .A1(n7610), .A2(n7630), .ZN(n8948) );
  OAI21_X1 U9297 ( .B1(n7630), .B2(n7610), .A(n8948), .ZN(n7618) );
  NOR2_X1 U9298 ( .A1(n8981), .A2(n9927), .ZN(n7617) );
  AOI21_X1 U9299 ( .B1(n8978), .B2(n9228), .A(n7611), .ZN(n7615) );
  NAND2_X1 U9300 ( .A1(n8984), .A2(n7612), .ZN(n7614) );
  NAND2_X1 U9301 ( .A1(n8894), .A2(n9226), .ZN(n7613) );
  NAND3_X1 U9302 ( .A1(n7615), .A2(n7614), .A3(n7613), .ZN(n7616) );
  AOI211_X1 U9303 ( .C1(n7618), .C2(n8959), .A(n7617), .B(n7616), .ZN(n7619)
         );
  INV_X1 U9304 ( .A(n7619), .ZN(P1_U3225) );
  OAI22_X1 U9305 ( .A1(n9944), .A2(n8711), .B1(n7621), .B2(n4463), .ZN(n7622)
         );
  XNOR2_X1 U9306 ( .A(n7622), .B(n4468), .ZN(n7625) );
  OR2_X1 U9307 ( .A1(n9944), .A2(n8775), .ZN(n7624) );
  NAND2_X1 U9308 ( .A1(n8944), .A2(n8774), .ZN(n7623) );
  AND2_X1 U9309 ( .A1(n7624), .A2(n7623), .ZN(n7626) );
  NAND2_X1 U9310 ( .A1(n7625), .A2(n7626), .ZN(n7645) );
  INV_X1 U9311 ( .A(n7625), .ZN(n7628) );
  INV_X1 U9312 ( .A(n7626), .ZN(n7627) );
  NAND2_X1 U9313 ( .A1(n7628), .A2(n7627), .ZN(n7629) );
  NAND2_X1 U9314 ( .A1(n7645), .A2(n7629), .ZN(n8947) );
  INV_X1 U9315 ( .A(n7630), .ZN(n7631) );
  AND2_X1 U9316 ( .A1(n7632), .A2(n7631), .ZN(n7633) );
  NOR2_X1 U9317 ( .A1(n8947), .A2(n7633), .ZN(n7634) );
  INV_X1 U9318 ( .A(n4449), .ZN(n8949) );
  OAI22_X1 U9319 ( .A1(n8953), .A2(n8711), .B1(n9942), .B2(n4463), .ZN(n7636)
         );
  XNOR2_X1 U9320 ( .A(n7636), .B(n4468), .ZN(n7640) );
  OR2_X1 U9321 ( .A1(n8953), .A2(n8775), .ZN(n7639) );
  NAND2_X1 U9322 ( .A1(n7637), .A2(n8774), .ZN(n7638) );
  AND2_X1 U9323 ( .A1(n7639), .A2(n7638), .ZN(n7641) );
  NAND2_X1 U9324 ( .A1(n7640), .A2(n7641), .ZN(n8797) );
  INV_X1 U9325 ( .A(n7640), .ZN(n7643) );
  INV_X1 U9326 ( .A(n7641), .ZN(n7642) );
  NAND2_X1 U9327 ( .A1(n7643), .A2(n7642), .ZN(n7644) );
  AND2_X1 U9328 ( .A1(n8797), .A2(n7644), .ZN(n7647) );
  NOR3_X1 U9329 ( .A1(n8949), .A2(n4799), .A3(n7647), .ZN(n7649) );
  INV_X1 U9330 ( .A(n8798), .ZN(n7648) );
  OAI21_X1 U9331 ( .B1(n7649), .B2(n7648), .A(n8959), .ZN(n7655) );
  AOI21_X1 U9332 ( .B1(n8978), .B2(n9226), .A(n7650), .ZN(n7651) );
  OAI21_X1 U9333 ( .B1(n8884), .B2(n8980), .A(n7651), .ZN(n7652) );
  AOI21_X1 U9334 ( .B1(n7653), .B2(n8984), .A(n7652), .ZN(n7654) );
  OAI211_X1 U9335 ( .C1(n9942), .C2(n8981), .A(n7655), .B(n7654), .ZN(P1_U3211) );
  INV_X1 U9336 ( .A(n9033), .ZN(n9138) );
  NAND2_X1 U9337 ( .A1(n9138), .A2(n9558), .ZN(n9028) );
  XNOR2_X1 U9338 ( .A(n7656), .B(n9028), .ZN(n9695) );
  INV_X1 U9339 ( .A(n9572), .ZN(n7659) );
  AOI21_X1 U9340 ( .B1(n7657), .B2(n8920), .A(n9535), .ZN(n7658) );
  NAND2_X1 U9341 ( .A1(n7659), .A2(n7658), .ZN(n9696) );
  INV_X1 U9342 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n7661) );
  INV_X1 U9343 ( .A(n8929), .ZN(n7660) );
  OAI22_X1 U9344 ( .A1(n9541), .A2(n7661), .B1(n7660), .B2(n9538), .ZN(n7662)
         );
  AOI21_X1 U9345 ( .B1(n9578), .B2(n8920), .A(n7662), .ZN(n7663) );
  OAI21_X1 U9346 ( .B1(n9696), .B2(n9580), .A(n7663), .ZN(n7668) );
  INV_X1 U9347 ( .A(n9028), .ZN(n9103) );
  XNOR2_X1 U9348 ( .A(n7664), .B(n9103), .ZN(n7666) );
  OAI22_X1 U9349 ( .A1(n8581), .A2(n9943), .B1(n9684), .B2(n9518), .ZN(n7665)
         );
  AOI21_X1 U9350 ( .B1(n7666), .B2(n9563), .A(n7665), .ZN(n9698) );
  NOR2_X1 U9351 ( .A1(n9698), .A2(n9877), .ZN(n7667) );
  AOI211_X1 U9352 ( .C1(n9582), .C2(n9695), .A(n7668), .B(n7667), .ZN(n7669)
         );
  INV_X1 U9353 ( .A(n7669), .ZN(P1_U3280) );
  NAND2_X1 U9354 ( .A1(n9820), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n7672) );
  OAI21_X1 U9355 ( .B1(n9820), .B2(P1_REG2_REG_13__SCAN_IN), .A(n7672), .ZN(
        n9816) );
  INV_X1 U9356 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n7673) );
  NAND2_X1 U9357 ( .A1(n7674), .A2(n7673), .ZN(n9249) );
  OAI21_X1 U9358 ( .B1(n7674), .B2(n7673), .A(n9249), .ZN(n7687) );
  NAND2_X1 U9359 ( .A1(n9810), .A2(P1_ADDR_REG_14__SCAN_IN), .ZN(n7675) );
  NAND2_X1 U9360 ( .A1(P1_U3084), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n8724) );
  OAI211_X1 U9361 ( .C1(n9859), .C2(n9263), .A(n7675), .B(n8724), .ZN(n7686)
         );
  INV_X1 U9362 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n10253) );
  OAI21_X1 U9363 ( .B1(n7678), .B2(n7677), .A(n7676), .ZN(n9822) );
  XNOR2_X1 U9364 ( .A(n9820), .B(P1_REG1_REG_13__SCAN_IN), .ZN(n9821) );
  INV_X1 U9365 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n9262) );
  AOI22_X1 U9366 ( .A1(n7681), .A2(n9262), .B1(P1_REG1_REG_14__SCAN_IN), .B2(
        n9263), .ZN(n7682) );
  AOI21_X1 U9367 ( .B1(n7683), .B2(n7682), .A(n9261), .ZN(n7684) );
  NOR2_X1 U9368 ( .A1(n7684), .A2(n9281), .ZN(n7685) );
  AOI211_X1 U9369 ( .C1(n7687), .C2(n9855), .A(n7686), .B(n7685), .ZN(n7688)
         );
  INV_X1 U9370 ( .A(n7688), .ZN(P1_U3255) );
  NAND2_X1 U9371 ( .A1(n7690), .A2(n7689), .ZN(n8118) );
  XNOR2_X1 U9372 ( .A(n8123), .B(P2_REG2_REG_16__SCAN_IN), .ZN(n8117) );
  XNOR2_X1 U9373 ( .A(n8118), .B(n8117), .ZN(n7703) );
  INV_X1 U9374 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n10156) );
  NAND2_X1 U9375 ( .A1(P2_U3152), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n7964) );
  OAI21_X1 U9376 ( .B1(n8106), .B2(n10156), .A(n7964), .ZN(n7701) );
  INV_X1 U9377 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n7693) );
  OAI22_X1 U9378 ( .A1(n7694), .A2(n7693), .B1(n7692), .B2(n7691), .ZN(n7698)
         );
  INV_X1 U9379 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n7696) );
  AOI22_X1 U9380 ( .A1(n8123), .A2(n7696), .B1(P2_REG1_REG_16__SCAN_IN), .B2(
        n7695), .ZN(n7697) );
  NOR2_X1 U9381 ( .A1(n7697), .A2(n7698), .ZN(n8124) );
  AOI21_X1 U9382 ( .B1(n7698), .B2(n7697), .A(n8124), .ZN(n7699) );
  NOR2_X1 U9383 ( .A1(n7699), .A2(n9989), .ZN(n7700) );
  AOI211_X1 U9384 ( .C1(n10003), .C2(n8123), .A(n7701), .B(n7700), .ZN(n7702)
         );
  OAI21_X1 U9385 ( .B1(n9987), .B2(n7703), .A(n7702), .ZN(P2_U3261) );
  AND2_X1 U9386 ( .A1(n7704), .A2(n8061), .ZN(n7738) );
  NOR2_X1 U9387 ( .A1(n7705), .A2(n7738), .ZN(n7706) );
  XNOR2_X1 U9388 ( .A(n7706), .B(n7708), .ZN(n7728) );
  NAND2_X1 U9389 ( .A1(n7840), .A2(n7707), .ZN(n7709) );
  XNOR2_X1 U9390 ( .A(n7709), .B(n7708), .ZN(n7710) );
  AOI222_X1 U9391 ( .A1(n10017), .A2(n7710), .B1(n8061), .B2(n8370), .C1(n8059), .C2(n8372), .ZN(n7727) );
  MUX2_X1 U9392 ( .A(n7711), .B(n7727), .S(n8417), .Z(n7719) );
  INV_X1 U9393 ( .A(n7712), .ZN(n7714) );
  INV_X1 U9394 ( .A(n7737), .ZN(n7716) );
  INV_X1 U9395 ( .A(n7852), .ZN(n7713) );
  AOI21_X1 U9396 ( .B1(n7737), .B2(n7714), .A(n7713), .ZN(n7725) );
  OAI22_X1 U9397 ( .A1(n10024), .A2(n7716), .B1(n7715), .B2(n10022), .ZN(n7717) );
  AOI21_X1 U9398 ( .B1(n7725), .B2(n8420), .A(n7717), .ZN(n7718) );
  OAI211_X1 U9399 ( .C1(n8379), .C2(n7728), .A(n7719), .B(n7718), .ZN(P2_U3285) );
  INV_X1 U9400 ( .A(n7720), .ZN(n7723) );
  OAI222_X1 U9401 ( .A1(P2_U3152), .A2(n7722), .B1(n8550), .B2(n7723), .C1(
        n7721), .C2(n8552), .ZN(P2_U3334) );
  OAI222_X1 U9402 ( .A1(n7724), .A2(P1_U3084), .B1(n9763), .B2(n7723), .C1(
        n10232), .C2(n9765), .ZN(P1_U3329) );
  INV_X1 U9403 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n7730) );
  AOI22_X1 U9404 ( .A1(n7725), .A2(n10019), .B1(n10063), .B2(n7737), .ZN(n7726) );
  OAI211_X1 U9405 ( .C1(n7728), .C2(n8523), .A(n7727), .B(n7726), .ZN(n7731)
         );
  NAND2_X1 U9406 ( .A1(n7731), .A2(n10283), .ZN(n7729) );
  OAI21_X1 U9407 ( .B1(n10283), .B2(n7730), .A(n7729), .ZN(P2_U3484) );
  NAND2_X1 U9408 ( .A1(n7731), .A2(n10100), .ZN(n7732) );
  OAI21_X1 U9409 ( .B1(n10100), .B2(n5948), .A(n7732), .ZN(P2_U3531) );
  OAI21_X1 U9410 ( .B1(n7744), .B2(n7733), .A(n7771), .ZN(n7749) );
  OAI22_X1 U9411 ( .A1(n8405), .A2(n7735), .B1(n7734), .B2(n8407), .ZN(n7748)
         );
  AOI22_X1 U9412 ( .A1(n7739), .A2(n7738), .B1(n8060), .B2(n7737), .ZN(n7740)
         );
  NAND2_X1 U9413 ( .A1(n7745), .A2(n7744), .ZN(n7746) );
  NAND2_X1 U9414 ( .A1(n7767), .A2(n7746), .ZN(n8517) );
  NOR2_X1 U9415 ( .A1(n8517), .A2(n10014), .ZN(n7747) );
  AOI211_X1 U9416 ( .C1(n10017), .C2(n7749), .A(n7748), .B(n7747), .ZN(n8516)
         );
  INV_X1 U9417 ( .A(n8517), .ZN(n7755) );
  AND2_X1 U9418 ( .A1(n7850), .A2(n8511), .ZN(n7750) );
  NOR2_X2 U9419 ( .A1(n7850), .A2(n8511), .ZN(n7775) );
  OR2_X1 U9420 ( .A1(n7750), .A2(n7775), .ZN(n8513) );
  AOI22_X1 U9421 ( .A1(n4281), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n7995), .B2(
        n8363), .ZN(n7752) );
  NAND2_X1 U9422 ( .A1(n8396), .A2(n8511), .ZN(n7751) );
  OAI211_X1 U9423 ( .C1(n8513), .C2(n8192), .A(n7752), .B(n7751), .ZN(n7753)
         );
  AOI21_X1 U9424 ( .B1(n7755), .B2(n7754), .A(n7753), .ZN(n7756) );
  OAI21_X1 U9425 ( .B1(n8516), .B2(n4281), .A(n7756), .ZN(P2_U3283) );
  INV_X1 U9426 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n7761) );
  OAI21_X1 U9427 ( .B1(n8806), .B2(n9943), .A(n7757), .ZN(n7759) );
  AOI211_X1 U9428 ( .C1(n9966), .C2(n7760), .A(n7759), .B(n7758), .ZN(n7763)
         );
  MUX2_X1 U9429 ( .A(n7761), .B(n7763), .S(n9970), .Z(n7762) );
  OAI21_X1 U9430 ( .B1(n4952), .B2(n9751), .A(n7762), .ZN(P1_U3484) );
  MUX2_X1 U9431 ( .A(n7764), .B(n7763), .S(n9986), .Z(n7765) );
  OAI21_X1 U9432 ( .B1(n4952), .B2(n9701), .A(n7765), .ZN(P1_U3533) );
  NAND2_X1 U9433 ( .A1(n8511), .A2(n8058), .ZN(n7766) );
  XNOR2_X1 U9434 ( .A(n7789), .B(n7768), .ZN(n8510) );
  INV_X1 U9435 ( .A(n7769), .ZN(n7773) );
  AOI21_X1 U9436 ( .B1(n7771), .B2(n7770), .A(n7790), .ZN(n7772) );
  NOR3_X1 U9437 ( .A1(n7773), .A2(n7772), .A3(n8305), .ZN(n7774) );
  OAI22_X1 U9438 ( .A1(n8406), .A2(n8407), .B1(n7845), .B2(n8405), .ZN(n7807)
         );
  NOR2_X1 U9439 ( .A1(n7774), .A2(n7807), .ZN(n8509) );
  MUX2_X1 U9440 ( .A(n7117), .B(n8509), .S(n8417), .Z(n7780) );
  INV_X1 U9441 ( .A(n7775), .ZN(n7776) );
  INV_X1 U9442 ( .A(n8506), .ZN(n7777) );
  AOI21_X1 U9443 ( .B1(n8506), .B2(n7776), .A(n7795), .ZN(n8507) );
  OAI22_X1 U9444 ( .A1(n7777), .A2(n10024), .B1(n10022), .B2(n7810), .ZN(n7778) );
  AOI21_X1 U9445 ( .B1(n8507), .B2(n8420), .A(n7778), .ZN(n7779) );
  OAI211_X1 U9446 ( .C1(n8510), .C2(n8379), .A(n7780), .B(n7779), .ZN(P2_U3282) );
  INV_X1 U9447 ( .A(n7781), .ZN(n7786) );
  OAI222_X1 U9448 ( .A1(P1_U3084), .A2(n7784), .B1(n9763), .B2(n7786), .C1(
        n7783), .C2(n7782), .ZN(P1_U3328) );
  OAI222_X1 U9449 ( .A1(n8552), .A2(n10263), .B1(n8550), .B2(n7786), .C1(
        P2_U3152), .C2(n7785), .ZN(P2_U3333) );
  XNOR2_X1 U9450 ( .A(n7787), .B(n7793), .ZN(n7788) );
  INV_X1 U9451 ( .A(n8042), .ZN(n8166) );
  AOI222_X1 U9452 ( .A1(n10017), .A2(n7788), .B1(n8057), .B2(n8370), .C1(n8166), .C2(n8372), .ZN(n8504) );
  OR2_X1 U9453 ( .A1(n8506), .A2(n8057), .ZN(n7791) );
  NAND2_X1 U9454 ( .A1(n7792), .A2(n7791), .ZN(n7794) );
  OAI21_X1 U9455 ( .B1(n7794), .B2(n7793), .A(n8165), .ZN(n8500) );
  INV_X1 U9456 ( .A(n8501), .ZN(n7800) );
  INV_X1 U9457 ( .A(n7795), .ZN(n7797) );
  INV_X1 U9458 ( .A(n8413), .ZN(n7796) );
  AOI21_X1 U9459 ( .B1(n8501), .B2(n7797), .A(n7796), .ZN(n8502) );
  NAND2_X1 U9460 ( .A1(n8502), .A2(n8420), .ZN(n7799) );
  AOI22_X1 U9461 ( .A1(n4281), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n8034), .B2(
        n8363), .ZN(n7798) );
  OAI211_X1 U9462 ( .C1(n7800), .C2(n10024), .A(n7799), .B(n7798), .ZN(n7801)
         );
  AOI21_X1 U9463 ( .B1(n8500), .B2(n8208), .A(n7801), .ZN(n7802) );
  OAI21_X1 U9464 ( .B1(n8504), .B2(n4281), .A(n7802), .ZN(P2_U3281) );
  INV_X1 U9465 ( .A(n7803), .ZN(n7804) );
  AOI21_X1 U9466 ( .B1(n7806), .B2(n7805), .A(n7804), .ZN(n7813) );
  NAND2_X1 U9467 ( .A1(n8005), .A2(n7807), .ZN(n7809) );
  OAI211_X1 U9468 ( .C1(n8037), .C2(n7810), .A(n7809), .B(n7808), .ZN(n7811)
         );
  AOI21_X1 U9469 ( .B1(n8048), .B2(n8506), .A(n7811), .ZN(n7812) );
  OAI21_X1 U9470 ( .B1(n7813), .B2(n8044), .A(n7812), .ZN(P2_U3217) );
  INV_X1 U9471 ( .A(n7814), .ZN(n7818) );
  OAI222_X1 U9472 ( .A1(n4464), .A2(P1_U3084), .B1(n9763), .B2(n7818), .C1(
        n7815), .C2(n9765), .ZN(P1_U3327) );
  OAI222_X1 U9473 ( .A1(P2_U3152), .A2(n7819), .B1(n8550), .B2(n7818), .C1(
        n7817), .C2(n8552), .ZN(P2_U3332) );
  INV_X1 U9474 ( .A(n7820), .ZN(n7831) );
  NAND2_X1 U9475 ( .A1(n9755), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n7821) );
  OAI211_X1 U9476 ( .C1(n7831), .C2(n9763), .A(n9806), .B(n7821), .ZN(P1_U3326) );
  XNOR2_X1 U9477 ( .A(n7822), .B(n7823), .ZN(n7830) );
  NOR2_X1 U9478 ( .A1(n8037), .A2(n8393), .ZN(n7828) );
  NAND2_X1 U9479 ( .A1(n8343), .A2(n8372), .ZN(n7825) );
  NAND2_X1 U9480 ( .A1(n8166), .A2(n8370), .ZN(n7824) );
  AND2_X1 U9481 ( .A1(n7825), .A2(n7824), .ZN(n8385) );
  NAND2_X1 U9482 ( .A1(P2_U3152), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n9995) );
  OAI21_X1 U9483 ( .B1(n7826), .B2(n8385), .A(n9995), .ZN(n7827) );
  AOI211_X1 U9484 ( .C1(n8490), .C2(n8048), .A(n7828), .B(n7827), .ZN(n7829)
         );
  OAI21_X1 U9485 ( .B1(n7830), .B2(n8044), .A(n7829), .ZN(P2_U3230) );
  OAI222_X1 U9486 ( .A1(n8552), .A2(n7832), .B1(n8550), .B2(n7831), .C1(n6369), 
        .C2(P2_U3152), .ZN(P2_U3331) );
  INV_X1 U9487 ( .A(n7833), .ZN(n7835) );
  AOI21_X1 U9488 ( .B1(n9755), .B2(P2_DATAO_REG_28__SCAN_IN), .A(n9805), .ZN(
        n7834) );
  OAI21_X1 U9489 ( .B1(n7835), .B2(n9763), .A(n7834), .ZN(P1_U3325) );
  XOR2_X1 U9490 ( .A(n7837), .B(n7843), .Z(n8524) );
  INV_X1 U9491 ( .A(n7838), .ZN(n7839) );
  NAND2_X1 U9492 ( .A1(n7840), .A2(n7839), .ZN(n7842) );
  NAND2_X1 U9493 ( .A1(n7842), .A2(n7841), .ZN(n7844) );
  XNOR2_X1 U9494 ( .A(n7844), .B(n4644), .ZN(n7848) );
  OAI22_X1 U9495 ( .A1(n8405), .A2(n7846), .B1(n7845), .B2(n8407), .ZN(n7847)
         );
  AOI21_X1 U9496 ( .B1(n7848), .B2(n10017), .A(n7847), .ZN(n8522) );
  MUX2_X1 U9497 ( .A(n7849), .B(n8522), .S(n8417), .Z(n7856) );
  INV_X1 U9498 ( .A(n7850), .ZN(n7851) );
  AOI21_X1 U9499 ( .B1(n8519), .B2(n7852), .A(n7851), .ZN(n8520) );
  OAI22_X1 U9500 ( .A1(n10024), .A2(n4795), .B1(n10022), .B2(n7853), .ZN(n7854) );
  AOI21_X1 U9501 ( .B1(n8520), .B2(n8420), .A(n7854), .ZN(n7855) );
  OAI211_X1 U9502 ( .C1(n8524), .C2(n8379), .A(n7856), .B(n7855), .ZN(P2_U3284) );
  OAI22_X1 U9503 ( .A1(n8008), .A2(n7857), .B1(n10090), .B2(n8044), .ZN(n7859)
         );
  NAND2_X1 U9504 ( .A1(n7859), .A2(n7858), .ZN(n7863) );
  AOI22_X1 U9505 ( .A1(n8048), .A2(n7861), .B1(P2_REG3_REG_0__SCAN_IN), .B2(
        n7860), .ZN(n7862) );
  OAI211_X1 U9506 ( .C1(n6958), .C2(n8041), .A(n7863), .B(n7862), .ZN(P2_U3234) );
  XOR2_X1 U9507 ( .A(n9105), .B(n7864), .Z(n9680) );
  NAND2_X1 U9508 ( .A1(n9559), .A2(n7865), .ZN(n7869) );
  NAND2_X1 U9509 ( .A1(n7869), .A2(n7866), .ZN(n7867) );
  NAND2_X1 U9510 ( .A1(n7867), .A2(n9563), .ZN(n7873) );
  AND2_X1 U9511 ( .A1(n7869), .A2(n7868), .ZN(n9550) );
  INV_X1 U9512 ( .A(n9105), .ZN(n7870) );
  AOI21_X1 U9513 ( .B1(n9550), .B2(n9151), .A(n7870), .ZN(n7872) );
  AOI22_X1 U9514 ( .A1(n9562), .A2(n9221), .B1(n9561), .B2(n9914), .ZN(n7871)
         );
  OAI21_X1 U9515 ( .B1(n7873), .B2(n7872), .A(n7871), .ZN(n9677) );
  INV_X1 U9516 ( .A(n9678), .ZN(n7876) );
  AOI211_X1 U9517 ( .C1(n9678), .C2(n4323), .A(n9535), .B(n9520), .ZN(n9676)
         );
  NAND2_X1 U9518 ( .A1(n9676), .A2(n9528), .ZN(n7875) );
  AOI22_X1 U9519 ( .A1(n9877), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n8727), .B2(
        n9874), .ZN(n7874) );
  OAI211_X1 U9520 ( .C1(n7876), .C2(n9526), .A(n7875), .B(n7874), .ZN(n7877)
         );
  AOI21_X1 U9521 ( .B1(n9541), .B2(n9677), .A(n7877), .ZN(n7878) );
  OAI21_X1 U9522 ( .B1(n9680), .B2(n9513), .A(n7878), .ZN(P1_U3277) );
  OAI21_X1 U9523 ( .B1(n8037), .B2(n7880), .A(n7879), .ZN(n7884) );
  OAI22_X1 U9524 ( .A1(n8020), .A2(n7882), .B1(n7881), .B2(n8041), .ZN(n7883)
         );
  AOI211_X1 U9525 ( .C1(n8048), .C2(n7885), .A(n7884), .B(n7883), .ZN(n7892)
         );
  NAND3_X1 U9526 ( .A1(n8049), .A2(n7886), .A3(n8063), .ZN(n7887) );
  OAI21_X1 U9527 ( .B1(n7132), .B2(n8044), .A(n7887), .ZN(n7890) );
  INV_X1 U9528 ( .A(n7888), .ZN(n7889) );
  NAND2_X1 U9529 ( .A1(n7890), .A2(n7889), .ZN(n7891) );
  OAI211_X1 U9530 ( .C1(n8044), .C2(n7893), .A(n7892), .B(n7891), .ZN(P2_U3233) );
  INV_X1 U9531 ( .A(n7894), .ZN(n9759) );
  OAI222_X1 U9532 ( .A1(n8552), .A2(n7895), .B1(n8550), .B2(n9759), .C1(n5803), 
        .C2(P2_U3152), .ZN(P2_U3328) );
  OAI222_X1 U9533 ( .A1(n8552), .A2(n10187), .B1(n8550), .B2(n7896), .C1(n6223), .C2(P2_U3152), .ZN(P2_U3336) );
  NOR2_X1 U9534 ( .A1(n8024), .A2(n7897), .ZN(n7900) );
  INV_X1 U9535 ( .A(n8179), .ZN(n8227) );
  NAND3_X1 U9536 ( .A1(n7898), .A2(n8049), .A3(n8227), .ZN(n7899) );
  OAI21_X1 U9537 ( .B1(n7900), .B2(n8044), .A(n7899), .ZN(n7902) );
  AOI22_X1 U9538 ( .A1(n8222), .A2(n8027), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3152), .ZN(n7903) );
  OAI21_X1 U9539 ( .B1(n8182), .B2(n8041), .A(n7903), .ZN(n7904) );
  AOI21_X1 U9540 ( .B1(n8033), .B2(n8227), .A(n7904), .ZN(n7905) );
  INV_X1 U9541 ( .A(n7906), .ZN(n7971) );
  NAND2_X1 U9542 ( .A1(n7971), .A2(n7907), .ZN(n7909) );
  OR3_X1 U9543 ( .A1(n7909), .A2(n7908), .A3(n8044), .ZN(n7916) );
  INV_X1 U9544 ( .A(n8272), .ZN(n8055) );
  NAND3_X1 U9545 ( .A1(n7909), .A2(n8049), .A3(n8055), .ZN(n7915) );
  AOI22_X1 U9546 ( .A1(n8027), .A2(n8293), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3152), .ZN(n7911) );
  NAND2_X1 U9547 ( .A1(n8320), .A2(n8033), .ZN(n7910) );
  OAI211_X1 U9548 ( .C1(n7912), .C2(n8041), .A(n7911), .B(n7910), .ZN(n7913)
         );
  AOI21_X1 U9549 ( .B1(n8461), .B2(n8048), .A(n7913), .ZN(n7914) );
  NAND3_X1 U9550 ( .A1(n7916), .A2(n7915), .A3(n7914), .ZN(P2_U3218) );
  NOR3_X1 U9551 ( .A1(n8008), .A2(n7917), .A3(n5842), .ZN(n7922) );
  AOI21_X1 U9552 ( .B1(n7919), .B2(n7918), .A(n8044), .ZN(n7921) );
  OAI21_X1 U9553 ( .B1(n7922), .B2(n7921), .A(n7920), .ZN(n7926) );
  OAI22_X1 U9554 ( .A1(n8405), .A2(n5842), .B1(n5868), .B2(n8407), .ZN(n10016)
         );
  AOI22_X1 U9555 ( .A1(n8048), .A2(n7923), .B1(n8005), .B2(n10016), .ZN(n7925)
         );
  MUX2_X1 U9556 ( .A(n8037), .B(P2_STATE_REG_SCAN_IN), .S(
        P2_REG3_REG_3__SCAN_IN), .Z(n7924) );
  NAND3_X1 U9557 ( .A1(n7926), .A2(n7925), .A3(n7924), .ZN(P2_U3220) );
  INV_X1 U9558 ( .A(n7927), .ZN(n7928) );
  AOI21_X1 U9559 ( .B1(n7930), .B2(n7929), .A(n7928), .ZN(n7935) );
  AND2_X1 U9560 ( .A1(P2_U3152), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8152) );
  NOR2_X1 U9561 ( .A1(n8037), .A2(n8354), .ZN(n7931) );
  AOI211_X1 U9562 ( .C1(n8018), .C2(n8344), .A(n8152), .B(n7931), .ZN(n7932)
         );
  OAI21_X1 U9563 ( .B1(n8020), .B2(n8169), .A(n7932), .ZN(n7933) );
  AOI21_X1 U9564 ( .B1(n8482), .B2(n8048), .A(n7933), .ZN(n7934) );
  OAI21_X1 U9565 ( .B1(n7935), .B2(n8044), .A(n7934), .ZN(P2_U3221) );
  XNOR2_X1 U9566 ( .A(n7936), .B(n7937), .ZN(n7943) );
  NAND2_X1 U9567 ( .A1(n8033), .A2(n8344), .ZN(n7940) );
  INV_X1 U9568 ( .A(n7938), .ZN(n8315) );
  AOI22_X1 U9569 ( .A1(n8027), .A2(n8315), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3152), .ZN(n7939) );
  OAI211_X1 U9570 ( .C1(n8009), .C2(n8041), .A(n7940), .B(n7939), .ZN(n7941)
         );
  AOI21_X1 U9571 ( .B1(n8471), .B2(n8048), .A(n7941), .ZN(n7942) );
  OAI21_X1 U9572 ( .B1(n7943), .B2(n8044), .A(n7942), .ZN(P2_U3225) );
  XNOR2_X1 U9573 ( .A(n7945), .B(n7944), .ZN(n7946) );
  XNOR2_X1 U9574 ( .A(n7947), .B(n7946), .ZN(n7954) );
  INV_X1 U9575 ( .A(n8251), .ZN(n7951) );
  OR2_X1 U9576 ( .A1(n8179), .A2(n8407), .ZN(n7949) );
  NAND2_X1 U9577 ( .A1(n8291), .A2(n8370), .ZN(n7948) );
  NAND2_X1 U9578 ( .A1(n7949), .A2(n7948), .ZN(n8256) );
  AOI22_X1 U9579 ( .A1(n8256), .A2(n8005), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3152), .ZN(n7950) );
  OAI21_X1 U9580 ( .B1(n7951), .B2(n8037), .A(n7950), .ZN(n7952) );
  AOI21_X1 U9581 ( .B1(n8452), .B2(n8048), .A(n7952), .ZN(n7953) );
  OAI21_X1 U9582 ( .B1(n7954), .B2(n8044), .A(n7953), .ZN(P2_U3227) );
  INV_X1 U9583 ( .A(n7955), .ZN(n7959) );
  AOI21_X1 U9584 ( .B1(n7955), .B2(n8043), .A(n7956), .ZN(n7957) );
  AOI21_X1 U9585 ( .B1(n7959), .B2(n7958), .A(n7957), .ZN(n7963) );
  NAND2_X1 U9586 ( .A1(n7961), .A2(n7960), .ZN(n7962) );
  XNOR2_X1 U9587 ( .A(n7963), .B(n7962), .ZN(n7969) );
  OAI21_X1 U9588 ( .B1(n8037), .B2(n8415), .A(n7964), .ZN(n7965) );
  AOI21_X1 U9589 ( .B1(n8018), .B2(n8371), .A(n7965), .ZN(n7966) );
  OAI21_X1 U9590 ( .B1(n8406), .B2(n8020), .A(n7966), .ZN(n7967) );
  AOI21_X1 U9591 ( .B1(n8048), .B2(n8494), .A(n7967), .ZN(n7968) );
  OAI21_X1 U9592 ( .B1(n7969), .B2(n8044), .A(n7968), .ZN(P2_U3228) );
  NAND2_X1 U9593 ( .A1(n7971), .A2(n7970), .ZN(n7973) );
  XNOR2_X1 U9594 ( .A(n7973), .B(n7972), .ZN(n7975) );
  NAND3_X1 U9595 ( .A1(n7975), .A2(n7993), .A3(n7974), .ZN(n7983) );
  INV_X1 U9596 ( .A(n7975), .ZN(n7976) );
  NAND3_X1 U9597 ( .A1(n7976), .A2(n8049), .A3(n8291), .ZN(n7982) );
  NOR2_X1 U9598 ( .A1(n8273), .A2(n8041), .ZN(n7980) );
  INV_X1 U9599 ( .A(n7977), .ZN(n8266) );
  AOI22_X1 U9600 ( .A1(n8266), .A2(n8027), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3152), .ZN(n7978) );
  OAI21_X1 U9601 ( .B1(n8020), .B2(n8272), .A(n7978), .ZN(n7979) );
  AOI211_X1 U9602 ( .C1(n8456), .C2(n8048), .A(n7980), .B(n7979), .ZN(n7981)
         );
  NAND3_X1 U9603 ( .A1(n7983), .A2(n7982), .A3(n7981), .ZN(P2_U3231) );
  XNOR2_X1 U9604 ( .A(n7985), .B(n7984), .ZN(n7990) );
  NAND2_X1 U9605 ( .A1(n8033), .A2(n8373), .ZN(n7987) );
  AOI22_X1 U9606 ( .A1(n8027), .A2(n8328), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3152), .ZN(n7986) );
  OAI211_X1 U9607 ( .C1(n8173), .C2(n8041), .A(n7987), .B(n7986), .ZN(n7988)
         );
  AOI21_X1 U9608 ( .B1(n8476), .B2(n8048), .A(n7988), .ZN(n7989) );
  OAI21_X1 U9609 ( .B1(n7990), .B2(n8044), .A(n7989), .ZN(P2_U3235) );
  XOR2_X1 U9610 ( .A(n7991), .B(n7992), .Z(n7994) );
  NAND2_X1 U9611 ( .A1(n7994), .A2(n7993), .ZN(n8002) );
  INV_X1 U9612 ( .A(n7995), .ZN(n7997) );
  OAI22_X1 U9613 ( .A1(n8037), .A2(n7997), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7996), .ZN(n7998) );
  AOI21_X1 U9614 ( .B1(n8018), .B2(n8057), .A(n7998), .ZN(n8001) );
  NAND2_X1 U9615 ( .A1(n8048), .A2(n8511), .ZN(n8000) );
  NAND2_X1 U9616 ( .A1(n8033), .A2(n8059), .ZN(n7999) );
  NAND4_X1 U9617 ( .A1(n8002), .A2(n8001), .A3(n8000), .A4(n7999), .ZN(
        P2_U3236) );
  INV_X1 U9618 ( .A(n8301), .ZN(n8007) );
  OR2_X1 U9619 ( .A1(n8272), .A2(n8407), .ZN(n8004) );
  NAND2_X1 U9620 ( .A1(n8334), .A2(n8370), .ZN(n8003) );
  NAND2_X1 U9621 ( .A1(n8004), .A2(n8003), .ZN(n8308) );
  AOI22_X1 U9622 ( .A1(n8308), .A2(n8005), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3152), .ZN(n8006) );
  OAI21_X1 U9623 ( .B1(n8007), .B2(n8037), .A(n8006), .ZN(n8012) );
  NOR3_X1 U9624 ( .A1(n8010), .A2(n8009), .A3(n8008), .ZN(n8011) );
  AOI211_X1 U9625 ( .C1(n8048), .C2(n8466), .A(n8012), .B(n8011), .ZN(n8013)
         );
  OAI21_X1 U9626 ( .B1(n8014), .B2(n8044), .A(n8013), .ZN(P2_U3237) );
  XNOR2_X1 U9627 ( .A(n8015), .B(n8016), .ZN(n8023) );
  NAND2_X1 U9628 ( .A1(P2_U3152), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8121) );
  OAI21_X1 U9629 ( .B1(n8037), .B2(n8362), .A(n8121), .ZN(n8017) );
  AOI21_X1 U9630 ( .B1(n8018), .B2(n8373), .A(n8017), .ZN(n8019) );
  OAI21_X1 U9631 ( .B1(n8408), .B2(n8020), .A(n8019), .ZN(n8021) );
  AOI21_X1 U9632 ( .B1(n8486), .B2(n8048), .A(n8021), .ZN(n8022) );
  OAI21_X1 U9633 ( .B1(n8023), .B2(n8044), .A(n8022), .ZN(P2_U3240) );
  INV_X1 U9634 ( .A(n8447), .ZN(n8235) );
  INV_X1 U9635 ( .A(n8273), .ZN(n8054) );
  AOI22_X1 U9636 ( .A1(n8233), .A2(n8027), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3152), .ZN(n8028) );
  OAI21_X1 U9637 ( .B1(n8239), .B2(n8041), .A(n8028), .ZN(n8029) );
  AOI21_X1 U9638 ( .B1(n8033), .B2(n8054), .A(n8029), .ZN(n8030) );
  OAI211_X1 U9639 ( .C1(n8235), .C2(n8032), .A(n8031), .B(n8030), .ZN(P2_U3242) );
  NAND2_X1 U9640 ( .A1(n8033), .A2(n8057), .ZN(n8040) );
  INV_X1 U9641 ( .A(n8034), .ZN(n8036) );
  OAI22_X1 U9642 ( .A1(n8037), .A2(n8036), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8035), .ZN(n8038) );
  INV_X1 U9643 ( .A(n8038), .ZN(n8039) );
  OAI211_X1 U9644 ( .C1(n8042), .C2(n8041), .A(n8040), .B(n8039), .ZN(n8047)
         );
  XNOR2_X1 U9645 ( .A(n7955), .B(n8043), .ZN(n8050) );
  NOR3_X1 U9646 ( .A1(n8050), .A2(n8045), .A3(n8044), .ZN(n8046) );
  AOI211_X1 U9647 ( .C1(n8048), .C2(n8501), .A(n8047), .B(n8046), .ZN(n8052)
         );
  INV_X1 U9648 ( .A(n8406), .ZN(n8163) );
  NAND3_X1 U9649 ( .A1(n8050), .A2(n8049), .A3(n8163), .ZN(n8051) );
  NAND2_X1 U9650 ( .A1(n8052), .A2(n8051), .ZN(P2_U3243) );
  MUX2_X1 U9651 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n8187), .S(P2_U3966), .Z(
        P2_U3582) );
  MUX2_X1 U9652 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n8226), .S(P2_U3966), .Z(
        P2_U3580) );
  MUX2_X1 U9653 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8053), .S(P2_U3966), .Z(
        P2_U3579) );
  MUX2_X1 U9654 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n8227), .S(P2_U3966), .Z(
        P2_U3578) );
  MUX2_X1 U9655 ( .A(n8054), .B(P2_DATAO_REG_25__SCAN_IN), .S(n8056), .Z(
        P2_U3577) );
  MUX2_X1 U9656 ( .A(n8291), .B(P2_DATAO_REG_24__SCAN_IN), .S(n8056), .Z(
        P2_U3576) );
  MUX2_X1 U9657 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(n8055), .S(P2_U3966), .Z(
        P2_U3575) );
  MUX2_X1 U9658 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8320), .S(P2_U3966), .Z(
        P2_U3574) );
  MUX2_X1 U9659 ( .A(n8334), .B(P2_DATAO_REG_21__SCAN_IN), .S(n8056), .Z(
        P2_U3573) );
  MUX2_X1 U9660 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8344), .S(P2_U3966), .Z(
        P2_U3572) );
  MUX2_X1 U9661 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n8373), .S(P2_U3966), .Z(
        P2_U3571) );
  MUX2_X1 U9662 ( .A(n8343), .B(P2_DATAO_REG_18__SCAN_IN), .S(n8056), .Z(
        P2_U3570) );
  MUX2_X1 U9663 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8371), .S(P2_U3966), .Z(
        P2_U3569) );
  MUX2_X1 U9664 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n8166), .S(P2_U3966), .Z(
        P2_U3568) );
  MUX2_X1 U9665 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n8163), .S(P2_U3966), .Z(
        P2_U3567) );
  MUX2_X1 U9666 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n8057), .S(P2_U3966), .Z(
        P2_U3566) );
  MUX2_X1 U9667 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n8058), .S(P2_U3966), .Z(
        P2_U3565) );
  MUX2_X1 U9668 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n8059), .S(P2_U3966), .Z(
        P2_U3564) );
  MUX2_X1 U9669 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n8060), .S(P2_U3966), .Z(
        P2_U3563) );
  MUX2_X1 U9670 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n8061), .S(P2_U3966), .Z(
        P2_U3562) );
  MUX2_X1 U9671 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n8062), .S(P2_U3966), .Z(
        P2_U3561) );
  MUX2_X1 U9672 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n8063), .S(P2_U3966), .Z(
        P2_U3560) );
  MUX2_X1 U9673 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n8064), .S(P2_U3966), .Z(
        P2_U3559) );
  MUX2_X1 U9674 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n8065), .S(P2_U3966), .Z(
        P2_U3558) );
  MUX2_X1 U9675 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(n8066), .S(P2_U3966), .Z(
        P2_U3557) );
  MUX2_X1 U9676 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n8067), .S(P2_U3966), .Z(
        P2_U3556) );
  MUX2_X1 U9677 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(n8068), .S(P2_U3966), .Z(
        P2_U3555) );
  MUX2_X1 U9678 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(n6388), .S(P2_U3966), .Z(
        P2_U3554) );
  MUX2_X1 U9679 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n6383), .S(P2_U3966), .Z(
        P2_U3553) );
  MUX2_X1 U9680 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(n6384), .S(P2_U3966), .Z(
        P2_U3552) );
  NAND2_X1 U9681 ( .A1(n10003), .A2(n8069), .ZN(n8081) );
  OAI211_X1 U9682 ( .C1(n8072), .C2(n8071), .A(n9999), .B(n8070), .ZN(n8080)
         );
  AOI22_X1 U9683 ( .A1(n9997), .A2(P2_ADDR_REG_1__SCAN_IN), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(P2_U3152), .ZN(n8079) );
  INV_X1 U9684 ( .A(n8073), .ZN(n8077) );
  OAI21_X1 U9685 ( .B1(n6727), .B2(n8075), .A(n8074), .ZN(n8076) );
  NAND3_X1 U9686 ( .A1(n10005), .A2(n8077), .A3(n8076), .ZN(n8078) );
  NAND4_X1 U9687 ( .A1(n8081), .A2(n8080), .A3(n8079), .A4(n8078), .ZN(
        P2_U3246) );
  NAND2_X1 U9688 ( .A1(n10003), .A2(n8082), .ZN(n8098) );
  AOI22_X1 U9689 ( .A1(n9997), .A2(P2_ADDR_REG_3__SCAN_IN), .B1(
        P2_REG3_REG_3__SCAN_IN), .B2(P2_U3152), .ZN(n8097) );
  INV_X1 U9690 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n8083) );
  MUX2_X1 U9691 ( .A(n8083), .B(P2_REG2_REG_3__SCAN_IN), .S(n8082), .Z(n8086)
         );
  NAND3_X1 U9692 ( .A1(n8086), .A2(n8085), .A3(n8084), .ZN(n8087) );
  NAND3_X1 U9693 ( .A1(n9999), .A2(n8088), .A3(n8087), .ZN(n8096) );
  INV_X1 U9694 ( .A(n8089), .ZN(n8094) );
  NAND3_X1 U9695 ( .A1(n8092), .A2(n8091), .A3(n8090), .ZN(n8093) );
  NAND3_X1 U9696 ( .A1(n10005), .A2(n8094), .A3(n8093), .ZN(n8095) );
  NAND4_X1 U9697 ( .A1(n8098), .A2(n8097), .A3(n8096), .A4(n8095), .ZN(
        P2_U3248) );
  OR3_X1 U9698 ( .A1(n8101), .A2(n8100), .A3(n8099), .ZN(n8102) );
  NAND3_X1 U9699 ( .A1(n8103), .A2(n10005), .A3(n8102), .ZN(n8116) );
  INV_X1 U9700 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n8105) );
  OAI21_X1 U9701 ( .B1(n8106), .B2(n8105), .A(n8104), .ZN(n8107) );
  AOI21_X1 U9702 ( .B1(n8108), .B2(n10003), .A(n8107), .ZN(n8115) );
  MUX2_X1 U9703 ( .A(n7550), .B(P2_REG2_REG_10__SCAN_IN), .S(n8108), .Z(n8109)
         );
  NAND3_X1 U9704 ( .A1(n8111), .A2(n8110), .A3(n8109), .ZN(n8112) );
  NAND3_X1 U9705 ( .A1(n9999), .A2(n8113), .A3(n8112), .ZN(n8114) );
  NAND3_X1 U9706 ( .A1(n8116), .A2(n8115), .A3(n8114), .ZN(P2_U3255) );
  XNOR2_X1 U9707 ( .A(n8127), .B(P2_REG2_REG_17__SCAN_IN), .ZN(n10000) );
  NAND2_X1 U9708 ( .A1(n8123), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n8119) );
  NAND2_X1 U9709 ( .A1(n10000), .A2(n10001), .ZN(n9998) );
  OAI21_X1 U9710 ( .B1(n8394), .B2(n8127), .A(n9998), .ZN(n8136) );
  XNOR2_X1 U9711 ( .A(n8136), .B(n8143), .ZN(n8120) );
  NAND2_X1 U9712 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n8120), .ZN(n8139) );
  OAI21_X1 U9713 ( .B1(P2_REG2_REG_18__SCAN_IN), .B2(n8120), .A(n8139), .ZN(
        n8135) );
  NAND2_X1 U9714 ( .A1(n9997), .A2(P2_ADDR_REG_18__SCAN_IN), .ZN(n8122) );
  NAND2_X1 U9715 ( .A1(n8122), .A2(n8121), .ZN(n8133) );
  XNOR2_X1 U9716 ( .A(n8127), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n10006) );
  OR2_X1 U9717 ( .A1(n8123), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n8126) );
  INV_X1 U9718 ( .A(n8124), .ZN(n8125) );
  AOI22_X1 U9719 ( .A1(n8137), .A2(n8142), .B1(P2_REG1_REG_18__SCAN_IN), .B2(
        n8143), .ZN(n8129) );
  NOR2_X1 U9720 ( .A1(n8130), .A2(n8129), .ZN(n8141) );
  AOI21_X1 U9721 ( .B1(n8130), .B2(n8129), .A(n8141), .ZN(n8131) );
  NOR2_X1 U9722 ( .A1(n8131), .A2(n9989), .ZN(n8132) );
  AOI211_X1 U9723 ( .C1(n10003), .C2(n8137), .A(n8133), .B(n8132), .ZN(n8134)
         );
  OAI21_X1 U9724 ( .B1(n8135), .B2(n9987), .A(n8134), .ZN(P2_U3263) );
  NAND2_X1 U9725 ( .A1(n8137), .A2(n8136), .ZN(n8138) );
  NAND2_X1 U9726 ( .A1(n8139), .A2(n8138), .ZN(n8140) );
  XOR2_X1 U9727 ( .A(n8140), .B(n8355), .Z(n8147) );
  AOI21_X1 U9728 ( .B1(n8143), .B2(n8142), .A(n8141), .ZN(n8144) );
  XOR2_X1 U9729 ( .A(n8145), .B(n8144), .Z(n8146) );
  OAI22_X1 U9730 ( .A1(n8147), .A2(n9987), .B1(n8146), .B2(n9989), .ZN(n8151)
         );
  NAND2_X1 U9731 ( .A1(n8146), .A2(n10005), .ZN(n8149) );
  NAND2_X1 U9732 ( .A1(n8147), .A2(n9999), .ZN(n8148) );
  NAND3_X1 U9733 ( .A1(n8149), .A2(n8148), .A3(n9988), .ZN(n8150) );
  AOI21_X1 U9734 ( .B1(n9997), .B2(P2_ADDR_REG_19__SCAN_IN), .A(n8152), .ZN(
        n8153) );
  INV_X1 U9735 ( .A(n8482), .ZN(n8347) );
  NAND2_X1 U9736 ( .A1(n8360), .A2(n8347), .ZN(n8346) );
  INV_X1 U9737 ( .A(n8466), .ZN(n8303) );
  NAND2_X1 U9738 ( .A1(n8253), .A2(n8265), .ZN(n8248) );
  NAND2_X1 U9739 ( .A1(n8224), .A2(n8232), .ZN(n8219) );
  NOR2_X1 U9740 ( .A1(n8417), .A2(n8155), .ZN(n8157) );
  NOR2_X1 U9741 ( .A1(n6369), .A2(n10176), .ZN(n8156) );
  NOR2_X1 U9742 ( .A1(n8407), .A2(n8156), .ZN(n8188) );
  NAND2_X1 U9743 ( .A1(n8188), .A2(n4655), .ZN(n8427) );
  NOR2_X1 U9744 ( .A1(n4281), .A2(n8427), .ZN(n8160) );
  AOI211_X1 U9745 ( .C1(n8423), .C2(n8396), .A(n8157), .B(n8160), .ZN(n8158)
         );
  OAI21_X1 U9746 ( .B1(n8425), .B2(n8192), .A(n8158), .ZN(P2_U3265) );
  NAND2_X1 U9747 ( .A1(n8159), .A2(n8191), .ZN(n8426) );
  NAND3_X1 U9748 ( .A1(n4327), .A2(n8420), .A3(n8426), .ZN(n8162) );
  AOI21_X1 U9749 ( .B1(n4281), .B2(P2_REG2_REG_30__SCAN_IN), .A(n8160), .ZN(
        n8161) );
  OAI211_X1 U9750 ( .C1(n8429), .C2(n10024), .A(n8162), .B(n8161), .ZN(
        P2_U3266) );
  OR2_X1 U9751 ( .A1(n8501), .A2(n8163), .ZN(n8164) );
  NAND2_X1 U9752 ( .A1(n8317), .A2(n8173), .ZN(n8175) );
  NOR2_X1 U9753 ( .A1(n8466), .A2(n8320), .ZN(n8176) );
  NAND2_X1 U9754 ( .A1(n8246), .A2(n8254), .ZN(n8245) );
  NAND2_X1 U9755 ( .A1(n8253), .A2(n8273), .ZN(n8178) );
  NAND2_X1 U9756 ( .A1(n8235), .A2(n8179), .ZN(n8180) );
  NAND2_X1 U9757 ( .A1(n8224), .A2(n8239), .ZN(n8181) );
  XNOR2_X1 U9758 ( .A(n8183), .B(n8186), .ZN(n8430) );
  INV_X1 U9759 ( .A(n8430), .ZN(n8199) );
  AOI22_X1 U9760 ( .A1(n8226), .A2(n8370), .B1(n8188), .B2(n8187), .ZN(n8189)
         );
  OAI21_X1 U9761 ( .B1(n8190), .B2(n8305), .A(n8189), .ZN(n8434) );
  OAI21_X1 U9762 ( .B1(n8209), .B2(n8431), .A(n8191), .ZN(n8432) );
  NOR2_X1 U9763 ( .A1(n8432), .A2(n8192), .ZN(n8197) );
  INV_X1 U9764 ( .A(n8193), .ZN(n8194) );
  AOI22_X1 U9765 ( .A1(n8194), .A2(n8363), .B1(P2_REG2_REG_29__SCAN_IN), .B2(
        n4281), .ZN(n8195) );
  OAI21_X1 U9766 ( .B1(n8431), .B2(n10024), .A(n8195), .ZN(n8196) );
  AOI211_X1 U9767 ( .C1(n8434), .C2(n8417), .A(n8197), .B(n8196), .ZN(n8198)
         );
  OAI21_X1 U9768 ( .B1(n8199), .B2(n8379), .A(n8198), .ZN(P2_U3267) );
  INV_X1 U9769 ( .A(n8200), .ZN(n8201) );
  AOI21_X1 U9770 ( .B1(n8201), .B2(n8207), .A(n8305), .ZN(n8205) );
  OAI22_X1 U9771 ( .A1(n8239), .A2(n8405), .B1(n8202), .B2(n8407), .ZN(n8203)
         );
  NAND2_X1 U9772 ( .A1(n8436), .A2(n8208), .ZN(n8216) );
  AOI21_X1 U9773 ( .B1(n8437), .B2(n8219), .A(n8209), .ZN(n8438) );
  INV_X1 U9774 ( .A(n8210), .ZN(n8211) );
  AOI22_X1 U9775 ( .A1(n8211), .A2(n8363), .B1(P2_REG2_REG_28__SCAN_IN), .B2(
        n4281), .ZN(n8212) );
  OAI21_X1 U9776 ( .B1(n8213), .B2(n10024), .A(n8212), .ZN(n8214) );
  AOI21_X1 U9777 ( .B1(n8438), .B2(n8420), .A(n8214), .ZN(n8215) );
  OAI211_X1 U9778 ( .C1(n4281), .C2(n8440), .A(n8216), .B(n8215), .ZN(P2_U3268) );
  INV_X1 U9779 ( .A(n8232), .ZN(n8221) );
  INV_X1 U9780 ( .A(n8219), .ZN(n8220) );
  AOI21_X1 U9781 ( .B1(n8441), .B2(n8221), .A(n8220), .ZN(n8442) );
  AOI22_X1 U9782 ( .A1(n8222), .A2(n8363), .B1(P2_REG2_REG_27__SCAN_IN), .B2(
        n4281), .ZN(n8223) );
  OAI21_X1 U9783 ( .B1(n8224), .B2(n10024), .A(n8223), .ZN(n8228) );
  OAI21_X1 U9784 ( .B1(n8230), .B2(n8237), .A(n8229), .ZN(n8231) );
  INV_X1 U9785 ( .A(n8231), .ZN(n8450) );
  AOI211_X1 U9786 ( .C1(n8447), .C2(n8248), .A(n4296), .B(n8232), .ZN(n8446)
         );
  AOI22_X1 U9787 ( .A1(n8233), .A2(n8363), .B1(P2_REG2_REG_26__SCAN_IN), .B2(
        n4281), .ZN(n8234) );
  OAI21_X1 U9788 ( .B1(n8235), .B2(n10024), .A(n8234), .ZN(n8243) );
  AOI211_X1 U9789 ( .C1(n8238), .C2(n8237), .A(n8305), .B(n8236), .ZN(n8241)
         );
  OAI22_X1 U9790 ( .A1(n8239), .A2(n8407), .B1(n8273), .B2(n8405), .ZN(n8240)
         );
  NOR2_X1 U9791 ( .A1(n8241), .A2(n8240), .ZN(n8449) );
  NOR2_X1 U9792 ( .A1(n8449), .A2(n4281), .ZN(n8242) );
  AOI211_X1 U9793 ( .C1(n8446), .C2(n8260), .A(n8243), .B(n8242), .ZN(n8244)
         );
  OAI21_X1 U9794 ( .B1(n8450), .B2(n8379), .A(n8244), .ZN(P2_U3270) );
  OAI21_X1 U9795 ( .B1(n8246), .B2(n8254), .A(n8245), .ZN(n8247) );
  INV_X1 U9796 ( .A(n8247), .ZN(n8455) );
  INV_X1 U9797 ( .A(n8265), .ZN(n8250) );
  INV_X1 U9798 ( .A(n8248), .ZN(n8249) );
  AOI211_X1 U9799 ( .C1(n8452), .C2(n8250), .A(n4296), .B(n8249), .ZN(n8451)
         );
  AOI22_X1 U9800 ( .A1(n8251), .A2(n8363), .B1(P2_REG2_REG_25__SCAN_IN), .B2(
        n4281), .ZN(n8252) );
  OAI21_X1 U9801 ( .B1(n8253), .B2(n10024), .A(n8252), .ZN(n8259) );
  XNOR2_X1 U9802 ( .A(n8255), .B(n8254), .ZN(n8257) );
  AOI21_X1 U9803 ( .B1(n8257), .B2(n10017), .A(n8256), .ZN(n8454) );
  NOR2_X1 U9804 ( .A1(n8454), .A2(n4281), .ZN(n8258) );
  AOI211_X1 U9805 ( .C1(n8260), .C2(n8451), .A(n8259), .B(n8258), .ZN(n8261)
         );
  OAI21_X1 U9806 ( .B1(n8455), .B2(n8379), .A(n8261), .ZN(P2_U3271) );
  INV_X1 U9807 ( .A(n8262), .ZN(n8263) );
  AOI21_X1 U9808 ( .B1(n8270), .B2(n8264), .A(n8263), .ZN(n8460) );
  AOI21_X1 U9809 ( .B1(n8456), .B2(n8282), .A(n8265), .ZN(n8457) );
  INV_X1 U9810 ( .A(n8456), .ZN(n8268) );
  AOI22_X1 U9811 ( .A1(n8266), .A2(n8363), .B1(P2_REG2_REG_24__SCAN_IN), .B2(
        n4281), .ZN(n8267) );
  OAI21_X1 U9812 ( .B1(n8268), .B2(n10024), .A(n8267), .ZN(n8278) );
  INV_X1 U9813 ( .A(n8269), .ZN(n8271) );
  AOI21_X1 U9814 ( .B1(n8271), .B2(n4838), .A(n8305), .ZN(n8276) );
  OAI22_X1 U9815 ( .A1(n8273), .A2(n8407), .B1(n8272), .B2(n8405), .ZN(n8274)
         );
  AOI21_X1 U9816 ( .B1(n8276), .B2(n8275), .A(n8274), .ZN(n8459) );
  NOR2_X1 U9817 ( .A1(n8459), .A2(n4281), .ZN(n8277) );
  AOI211_X1 U9818 ( .C1(n8457), .C2(n8420), .A(n8278), .B(n8277), .ZN(n8279)
         );
  OAI21_X1 U9819 ( .B1(n8460), .B2(n8379), .A(n8279), .ZN(P2_U3272) );
  OAI21_X1 U9820 ( .B1(n8281), .B2(n8287), .A(n8280), .ZN(n8465) );
  INV_X1 U9821 ( .A(n8299), .ZN(n8283) );
  AOI21_X1 U9822 ( .B1(n8461), .B2(n8283), .A(n4787), .ZN(n8462) );
  OAI22_X1 U9823 ( .A1(n8285), .A2(n10024), .B1(n8417), .B2(n8284), .ZN(n8296)
         );
  INV_X1 U9824 ( .A(n8286), .ZN(n8290) );
  OAI21_X1 U9825 ( .B1(n8304), .B2(n8288), .A(n8287), .ZN(n8289) );
  NAND2_X1 U9826 ( .A1(n8290), .A2(n8289), .ZN(n8292) );
  AOI222_X1 U9827 ( .A1(n10017), .A2(n8292), .B1(n8291), .B2(n8372), .C1(n8320), .C2(n8370), .ZN(n8464) );
  NAND2_X1 U9828 ( .A1(n8293), .A2(n8363), .ZN(n8294) );
  AOI21_X1 U9829 ( .B1(n8464), .B2(n8294), .A(n4281), .ZN(n8295) );
  AOI211_X1 U9830 ( .C1(n8462), .C2(n8420), .A(n8296), .B(n8295), .ZN(n8297)
         );
  OAI21_X1 U9831 ( .B1(n8379), .B2(n8465), .A(n8297), .ZN(P2_U3273) );
  XOR2_X1 U9832 ( .A(n8298), .B(n8307), .Z(n8470) );
  INV_X1 U9833 ( .A(n8313), .ZN(n8300) );
  AOI21_X1 U9834 ( .B1(n8466), .B2(n8300), .A(n8299), .ZN(n8467) );
  AOI22_X1 U9835 ( .A1(n8301), .A2(n8363), .B1(n4281), .B2(
        P2_REG2_REG_22__SCAN_IN), .ZN(n8302) );
  OAI21_X1 U9836 ( .B1(n8303), .B2(n10024), .A(n8302), .ZN(n8311) );
  AOI211_X1 U9837 ( .C1(n8307), .C2(n8306), .A(n8305), .B(n8304), .ZN(n8309)
         );
  NOR2_X1 U9838 ( .A1(n8309), .A2(n8308), .ZN(n8469) );
  NOR2_X1 U9839 ( .A1(n8469), .A2(n4281), .ZN(n8310) );
  AOI211_X1 U9840 ( .C1(n8467), .C2(n8420), .A(n8311), .B(n8310), .ZN(n8312)
         );
  OAI21_X1 U9841 ( .B1(n8470), .B2(n8379), .A(n8312), .ZN(P2_U3274) );
  AOI21_X1 U9842 ( .B1(n8471), .B2(n8314), .A(n8313), .ZN(n8472) );
  AOI22_X1 U9843 ( .A1(n4281), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n8315), .B2(
        n8363), .ZN(n8316) );
  OAI21_X1 U9844 ( .B1(n8317), .B2(n10024), .A(n8316), .ZN(n8323) );
  XNOR2_X1 U9845 ( .A(n8319), .B(n8318), .ZN(n8321) );
  AOI222_X1 U9846 ( .A1(n10017), .A2(n8321), .B1(n8344), .B2(n8370), .C1(n8320), .C2(n8372), .ZN(n8474) );
  NOR2_X1 U9847 ( .A1(n8474), .A2(n4281), .ZN(n8322) );
  AOI211_X1 U9848 ( .C1(n8472), .C2(n8420), .A(n8323), .B(n8322), .ZN(n8324)
         );
  OAI21_X1 U9849 ( .B1(n8475), .B2(n8379), .A(n8324), .ZN(P2_U3275) );
  OAI21_X1 U9850 ( .B1(n8327), .B2(n8326), .A(n8325), .ZN(n8480) );
  XNOR2_X1 U9851 ( .A(n8346), .B(n8330), .ZN(n8477) );
  AOI22_X1 U9852 ( .A1(n4281), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n8328), .B2(
        n8363), .ZN(n8329) );
  OAI21_X1 U9853 ( .B1(n8330), .B2(n10024), .A(n8329), .ZN(n8337) );
  NAND2_X1 U9854 ( .A1(n8340), .A2(n8331), .ZN(n8333) );
  XNOR2_X1 U9855 ( .A(n8333), .B(n8332), .ZN(n8335) );
  AOI222_X1 U9856 ( .A1(n10017), .A2(n8335), .B1(n8334), .B2(n8372), .C1(n8373), .C2(n8370), .ZN(n8479) );
  NOR2_X1 U9857 ( .A1(n8479), .A2(n4281), .ZN(n8336) );
  AOI211_X1 U9858 ( .C1(n8477), .C2(n8420), .A(n8337), .B(n8336), .ZN(n8338)
         );
  OAI21_X1 U9859 ( .B1(n8480), .B2(n8379), .A(n8338), .ZN(P2_U3276) );
  XOR2_X1 U9860 ( .A(n8342), .B(n8339), .Z(n8484) );
  OAI21_X1 U9861 ( .B1(n8342), .B2(n8341), .A(n8340), .ZN(n8345) );
  AOI222_X1 U9862 ( .A1(n10017), .A2(n8345), .B1(n8344), .B2(n8372), .C1(n8343), .C2(n8370), .ZN(n8351) );
  INV_X1 U9863 ( .A(n8484), .ZN(n8349) );
  OAI211_X1 U9864 ( .C1(n8347), .C2(n8360), .A(n8346), .B(n10019), .ZN(n8348)
         );
  NAND2_X1 U9865 ( .A1(n8351), .A2(n8348), .ZN(n8481) );
  AOI21_X1 U9866 ( .B1(n8349), .B2(n8387), .A(n8481), .ZN(n8350) );
  AOI211_X1 U9867 ( .C1(n4291), .C2(n8351), .A(n4281), .B(n8350), .ZN(n8353)
         );
  INV_X1 U9868 ( .A(n8353), .ZN(n8358) );
  OAI22_X1 U9869 ( .A1(n8417), .A2(n8355), .B1(n8354), .B2(n10022), .ZN(n8356)
         );
  AOI21_X1 U9870 ( .B1(n8482), .B2(n8396), .A(n8356), .ZN(n8357) );
  OAI211_X1 U9871 ( .C1(n8484), .C2(n10025), .A(n8358), .B(n8357), .ZN(
        P2_U3277) );
  XNOR2_X1 U9872 ( .A(n8359), .B(n8368), .ZN(n8489) );
  AOI211_X1 U9873 ( .C1(n8486), .C2(n8361), .A(n4296), .B(n8360), .ZN(n8485)
         );
  INV_X1 U9874 ( .A(n8362), .ZN(n8364) );
  AOI22_X1 U9875 ( .A1(n4281), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n8364), .B2(
        n8363), .ZN(n8365) );
  OAI21_X1 U9876 ( .B1(n4768), .B2(n10024), .A(n8365), .ZN(n8376) );
  AND2_X1 U9877 ( .A1(n8383), .A2(n8366), .ZN(n8369) );
  OAI21_X1 U9878 ( .B1(n8369), .B2(n8368), .A(n8367), .ZN(n8374) );
  AOI222_X1 U9879 ( .A1(n10017), .A2(n8374), .B1(n8373), .B2(n8372), .C1(n8371), .C2(n8370), .ZN(n8488) );
  NOR2_X1 U9880 ( .A1(n8488), .A2(n4281), .ZN(n8375) );
  AOI211_X1 U9881 ( .C1(n8485), .C2(n8377), .A(n8376), .B(n8375), .ZN(n8378)
         );
  OAI21_X1 U9882 ( .B1(n8489), .B2(n8379), .A(n8378), .ZN(P2_U3278) );
  OAI21_X1 U9883 ( .B1(n4454), .B2(n8381), .A(n8380), .ZN(n8491) );
  INV_X1 U9884 ( .A(n8491), .ZN(n8399) );
  OAI211_X1 U9885 ( .C1(n8384), .C2(n4719), .A(n8383), .B(n10017), .ZN(n8386)
         );
  NAND2_X1 U9886 ( .A1(n8386), .A2(n8385), .ZN(n8391) );
  INV_X1 U9887 ( .A(n8387), .ZN(n8389) );
  XOR2_X1 U9888 ( .A(n4393), .B(n8490), .Z(n8388) );
  AOI21_X1 U9889 ( .B1(n10019), .B2(n8388), .A(n8391), .ZN(n8492) );
  OAI21_X1 U9890 ( .B1(n8399), .B2(n8389), .A(n8492), .ZN(n8390) );
  OAI211_X1 U9891 ( .C1(n8392), .C2(n8391), .A(n8390), .B(n8417), .ZN(n8398)
         );
  OAI22_X1 U9892 ( .A1(n8417), .A2(n8394), .B1(n8393), .B2(n10022), .ZN(n8395)
         );
  AOI21_X1 U9893 ( .B1(n8490), .B2(n8396), .A(n8395), .ZN(n8397) );
  OAI211_X1 U9894 ( .C1(n8399), .C2(n10025), .A(n8398), .B(n8397), .ZN(
        P2_U3279) );
  XNOR2_X1 U9895 ( .A(n8400), .B(n8404), .ZN(n8402) );
  INV_X1 U9896 ( .A(n8402), .ZN(n8497) );
  NAND2_X1 U9897 ( .A1(n8402), .A2(n8401), .ZN(n8412) );
  XNOR2_X1 U9898 ( .A(n8403), .B(n8404), .ZN(n8410) );
  OAI22_X1 U9899 ( .A1(n8408), .A2(n8407), .B1(n8406), .B2(n8405), .ZN(n8409)
         );
  AOI21_X1 U9900 ( .B1(n8410), .B2(n10017), .A(n8409), .ZN(n8411) );
  NAND2_X1 U9901 ( .A1(n8412), .A2(n8411), .ZN(n8499) );
  NAND2_X1 U9902 ( .A1(n8499), .A2(n8417), .ZN(n8422) );
  NAND2_X1 U9903 ( .A1(n8413), .A2(n8494), .ZN(n8414) );
  AND2_X1 U9904 ( .A1(n4393), .A2(n8414), .ZN(n8495) );
  NOR2_X1 U9905 ( .A1(n4772), .A2(n10024), .ZN(n8419) );
  OAI22_X1 U9906 ( .A1(n8417), .A2(n8416), .B1(n8415), .B2(n10022), .ZN(n8418)
         );
  AOI211_X1 U9907 ( .C1(n8495), .C2(n8420), .A(n8419), .B(n8418), .ZN(n8421)
         );
  OAI211_X1 U9908 ( .C1(n8497), .C2(n10025), .A(n8422), .B(n8421), .ZN(
        P2_U3280) );
  NAND2_X1 U9909 ( .A1(n8423), .A2(n10063), .ZN(n8424) );
  MUX2_X1 U9910 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n8525), .S(n10100), .Z(
        P2_U3551) );
  NAND3_X1 U9911 ( .A1(n4327), .A2(n10019), .A3(n8426), .ZN(n8428) );
  OAI211_X1 U9912 ( .C1(n8429), .C2(n10077), .A(n8428), .B(n8427), .ZN(n8526)
         );
  MUX2_X1 U9913 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n8526), .S(n10100), .Z(
        P2_U3550) );
  NAND2_X1 U9914 ( .A1(n8430), .A2(n10086), .ZN(n8435) );
  OAI22_X1 U9915 ( .A1(n8432), .A2(n4296), .B1(n8431), .B2(n10077), .ZN(n8433)
         );
  MUX2_X1 U9916 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n8527), .S(n10100), .Z(
        P2_U3549) );
  AOI22_X1 U9917 ( .A1(n8442), .A2(n10019), .B1(n10063), .B2(n8441), .ZN(n8443) );
  OAI211_X1 U9918 ( .C1(n8445), .C2(n8523), .A(n8444), .B(n8443), .ZN(n8528)
         );
  MUX2_X1 U9919 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n8528), .S(n10100), .Z(
        P2_U3547) );
  AOI21_X1 U9920 ( .B1(n10063), .B2(n8447), .A(n8446), .ZN(n8448) );
  OAI211_X1 U9921 ( .C1(n8450), .C2(n8523), .A(n8449), .B(n8448), .ZN(n8529)
         );
  MUX2_X1 U9922 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n8529), .S(n10100), .Z(
        P2_U3546) );
  AOI21_X1 U9923 ( .B1(n10063), .B2(n8452), .A(n8451), .ZN(n8453) );
  OAI211_X1 U9924 ( .C1(n8455), .C2(n8523), .A(n8454), .B(n8453), .ZN(n8530)
         );
  MUX2_X1 U9925 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n8530), .S(n10100), .Z(
        P2_U3545) );
  AOI22_X1 U9926 ( .A1(n8457), .A2(n10019), .B1(n10063), .B2(n8456), .ZN(n8458) );
  OAI211_X1 U9927 ( .C1(n8460), .C2(n8523), .A(n8459), .B(n8458), .ZN(n8531)
         );
  MUX2_X1 U9928 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n8531), .S(n10100), .Z(
        P2_U3544) );
  AOI22_X1 U9929 ( .A1(n8462), .A2(n10019), .B1(n10063), .B2(n8461), .ZN(n8463) );
  OAI211_X1 U9930 ( .C1(n8465), .C2(n8523), .A(n8464), .B(n8463), .ZN(n8532)
         );
  MUX2_X1 U9931 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n8532), .S(n10100), .Z(
        P2_U3543) );
  AOI22_X1 U9932 ( .A1(n8467), .A2(n10019), .B1(n10063), .B2(n8466), .ZN(n8468) );
  OAI211_X1 U9933 ( .C1(n8470), .C2(n8523), .A(n8469), .B(n8468), .ZN(n8533)
         );
  MUX2_X1 U9934 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n8533), .S(n10100), .Z(
        P2_U3542) );
  AOI22_X1 U9935 ( .A1(n8472), .A2(n10019), .B1(n10063), .B2(n8471), .ZN(n8473) );
  OAI211_X1 U9936 ( .C1(n8475), .C2(n8523), .A(n8474), .B(n8473), .ZN(n8534)
         );
  MUX2_X1 U9937 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n8534), .S(n10100), .Z(
        P2_U3541) );
  AOI22_X1 U9938 ( .A1(n8477), .A2(n10019), .B1(n10063), .B2(n8476), .ZN(n8478) );
  OAI211_X1 U9939 ( .C1(n8480), .C2(n8523), .A(n8479), .B(n8478), .ZN(n8535)
         );
  MUX2_X1 U9940 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n8535), .S(n10100), .Z(
        P2_U3540) );
  AOI21_X1 U9941 ( .B1(n10063), .B2(n8482), .A(n8481), .ZN(n8483) );
  OAI21_X1 U9942 ( .B1(n8484), .B2(n8523), .A(n8483), .ZN(n8536) );
  MUX2_X1 U9943 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n8536), .S(n10100), .Z(
        P2_U3539) );
  AOI21_X1 U9944 ( .B1(n10063), .B2(n8486), .A(n8485), .ZN(n8487) );
  OAI211_X1 U9945 ( .C1(n8489), .C2(n8523), .A(n8488), .B(n8487), .ZN(n8537)
         );
  MUX2_X1 U9946 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n8537), .S(n10100), .Z(
        P2_U3538) );
  NAND2_X1 U9947 ( .A1(n8491), .A2(n10086), .ZN(n8493) );
  OAI211_X1 U9948 ( .C1(n4722), .C2(n10077), .A(n8493), .B(n8492), .ZN(n8538)
         );
  MUX2_X1 U9949 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n8538), .S(n10100), .Z(
        P2_U3537) );
  AOI22_X1 U9950 ( .A1(n8495), .A2(n10019), .B1(n10063), .B2(n8494), .ZN(n8496) );
  OAI21_X1 U9951 ( .B1(n8497), .B2(n8518), .A(n8496), .ZN(n8498) );
  MUX2_X1 U9952 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n8539), .S(n10100), .Z(
        P2_U3536) );
  INV_X1 U9953 ( .A(n8500), .ZN(n8505) );
  AOI22_X1 U9954 ( .A1(n8502), .A2(n10019), .B1(n10063), .B2(n8501), .ZN(n8503) );
  OAI211_X1 U9955 ( .C1(n8505), .C2(n8523), .A(n8504), .B(n8503), .ZN(n8540)
         );
  MUX2_X1 U9956 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n8540), .S(n10100), .Z(
        P2_U3535) );
  AOI22_X1 U9957 ( .A1(n8507), .A2(n10019), .B1(n10063), .B2(n8506), .ZN(n8508) );
  OAI211_X1 U9958 ( .C1(n8510), .C2(n8523), .A(n8509), .B(n8508), .ZN(n8541)
         );
  MUX2_X1 U9959 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n8541), .S(n10100), .Z(
        P2_U3534) );
  INV_X1 U9960 ( .A(n8511), .ZN(n8512) );
  OAI22_X1 U9961 ( .A1(n8513), .A2(n4296), .B1(n8512), .B2(n10077), .ZN(n8514)
         );
  INV_X1 U9962 ( .A(n8514), .ZN(n8515) );
  OAI211_X1 U9963 ( .C1(n8518), .C2(n8517), .A(n8516), .B(n8515), .ZN(n8542)
         );
  MUX2_X1 U9964 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n8542), .S(n10100), .Z(
        P2_U3533) );
  AOI22_X1 U9965 ( .A1(n8520), .A2(n10019), .B1(n10063), .B2(n8519), .ZN(n8521) );
  OAI211_X1 U9966 ( .C1(n8524), .C2(n8523), .A(n8522), .B(n8521), .ZN(n8543)
         );
  MUX2_X1 U9967 ( .A(n8543), .B(P2_REG1_REG_12__SCAN_IN), .S(n10098), .Z(
        P2_U3532) );
  MUX2_X1 U9968 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n8525), .S(n10283), .Z(
        P2_U3519) );
  MUX2_X1 U9969 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n8526), .S(n10283), .Z(
        P2_U3518) );
  MUX2_X1 U9970 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n8527), .S(n10283), .Z(
        P2_U3517) );
  MUX2_X1 U9971 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n8528), .S(n10283), .Z(
        P2_U3515) );
  MUX2_X1 U9972 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n8529), .S(n10283), .Z(
        P2_U3514) );
  MUX2_X1 U9973 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n8530), .S(n10283), .Z(
        P2_U3513) );
  MUX2_X1 U9974 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n8531), .S(n10283), .Z(
        P2_U3512) );
  MUX2_X1 U9975 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n8532), .S(n10283), .Z(
        P2_U3511) );
  MUX2_X1 U9976 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n8533), .S(n10283), .Z(
        P2_U3510) );
  MUX2_X1 U9977 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n8534), .S(n10283), .Z(
        P2_U3509) );
  MUX2_X1 U9978 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n8535), .S(n10283), .Z(
        P2_U3508) );
  MUX2_X1 U9979 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n8536), .S(n10283), .Z(
        P2_U3507) );
  MUX2_X1 U9980 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n8537), .S(n10283), .Z(
        P2_U3505) );
  MUX2_X1 U9981 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n8538), .S(n10283), .Z(
        P2_U3502) );
  MUX2_X1 U9982 ( .A(n8539), .B(P2_REG0_REG_16__SCAN_IN), .S(n10281), .Z(
        P2_U3499) );
  MUX2_X1 U9983 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n8540), .S(n10283), .Z(
        P2_U3496) );
  MUX2_X1 U9984 ( .A(P2_REG0_REG_14__SCAN_IN), .B(n8541), .S(n10283), .Z(
        P2_U3493) );
  MUX2_X1 U9985 ( .A(P2_REG0_REG_13__SCAN_IN), .B(n8542), .S(n10283), .Z(
        P2_U3490) );
  MUX2_X1 U9986 ( .A(n8543), .B(P2_REG0_REG_12__SCAN_IN), .S(n10281), .Z(
        P2_U3487) );
  INV_X1 U9987 ( .A(n8544), .ZN(n9757) );
  NAND3_X1 U9988 ( .A1(n8545), .A2(P2_IR_REG_31__SCAN_IN), .A3(
        P2_STATE_REG_SCAN_IN), .ZN(n8547) );
  OAI22_X1 U9989 ( .A1(n5801), .A2(n8547), .B1(n8546), .B2(n8552), .ZN(n8548)
         );
  INV_X1 U9990 ( .A(n8548), .ZN(n8549) );
  OAI21_X1 U9991 ( .B1(n9757), .B2(n8550), .A(n8549), .ZN(P2_U3327) );
  INV_X1 U9992 ( .A(n8551), .ZN(n9762) );
  OAI222_X1 U9993 ( .A1(n8550), .A2(n9762), .B1(P2_U3152), .B2(n8553), .C1(
        n10165), .C2(n8552), .ZN(P2_U3329) );
  MUX2_X1 U9994 ( .A(n8554), .B(P2_IR_REG_0__SCAN_IN), .S(P2_STATE_REG_SCAN_IN), .Z(P2_U3358) );
  INV_X1 U9995 ( .A(n9603), .ZN(n9322) );
  OAI22_X1 U9996 ( .A1(n9714), .A2(n8711), .B1(n9609), .B2(n8775), .ZN(n8697)
         );
  INV_X1 U9997 ( .A(n8697), .ZN(n8700) );
  NAND2_X1 U9998 ( .A1(n9352), .A2(n4278), .ZN(n8556) );
  OR2_X1 U9999 ( .A1(n9609), .A2(n8779), .ZN(n8555) );
  NAND2_X1 U10000 ( .A1(n8556), .A2(n8555), .ZN(n8557) );
  XNOR2_X1 U10001 ( .A(n8557), .B(n4285), .ZN(n8698) );
  INV_X1 U10002 ( .A(n8698), .ZN(n8699) );
  OAI22_X1 U10003 ( .A1(n8884), .A2(n8711), .B1(n9953), .B2(n4463), .ZN(n8558)
         );
  XNOR2_X1 U10004 ( .A(n8558), .B(n4285), .ZN(n8876) );
  OR2_X1 U10005 ( .A1(n8884), .A2(n8775), .ZN(n8561) );
  NAND2_X1 U10006 ( .A1(n8559), .A2(n8774), .ZN(n8560) );
  NAND2_X1 U10007 ( .A1(n8561), .A2(n8560), .ZN(n8800) );
  NAND2_X1 U10008 ( .A1(n8566), .A2(n4278), .ZN(n8564) );
  OAI21_X1 U10009 ( .B1(n8806), .B2(n8711), .A(n8564), .ZN(n8565) );
  XNOR2_X1 U10010 ( .A(n8565), .B(n4468), .ZN(n8569) );
  OR2_X1 U10011 ( .A1(n8806), .A2(n8775), .ZN(n8568) );
  NAND2_X1 U10012 ( .A1(n8566), .A2(n8774), .ZN(n8567) );
  AND2_X1 U10013 ( .A1(n8568), .A2(n8567), .ZN(n8570) );
  NAND2_X1 U10014 ( .A1(n8569), .A2(n8570), .ZN(n8576) );
  INV_X1 U10015 ( .A(n8569), .ZN(n8572) );
  INV_X1 U10016 ( .A(n8570), .ZN(n8571) );
  NAND2_X1 U10017 ( .A1(n8572), .A2(n8571), .ZN(n8573) );
  NAND2_X1 U10018 ( .A1(n8576), .A2(n8573), .ZN(n8877) );
  AND2_X1 U10019 ( .A1(n8876), .A2(n8800), .ZN(n8574) );
  NOR2_X1 U10020 ( .A1(n8877), .A2(n8574), .ZN(n8575) );
  NAND2_X1 U10021 ( .A1(n8580), .A2(n4278), .ZN(n8578) );
  OR2_X1 U10022 ( .A1(n8581), .A2(n8779), .ZN(n8577) );
  NAND2_X1 U10023 ( .A1(n8578), .A2(n8577), .ZN(n8579) );
  XNOR2_X1 U10024 ( .A(n8579), .B(n4468), .ZN(n8591) );
  NAND2_X1 U10025 ( .A1(n8580), .A2(n4476), .ZN(n8583) );
  OR2_X1 U10026 ( .A1(n8581), .A2(n8775), .ZN(n8582) );
  NAND2_X1 U10027 ( .A1(n8583), .A2(n8582), .ZN(n8589) );
  XNOR2_X1 U10028 ( .A(n8591), .B(n8589), .ZN(n8754) );
  NAND2_X1 U10029 ( .A1(n8920), .A2(n4278), .ZN(n8585) );
  OR2_X1 U10030 ( .A1(n9575), .A2(n8779), .ZN(n8584) );
  NAND2_X1 U10031 ( .A1(n8585), .A2(n8584), .ZN(n8586) );
  XNOR2_X1 U10032 ( .A(n8586), .B(n4468), .ZN(n8593) );
  NAND2_X1 U10033 ( .A1(n8920), .A2(n4476), .ZN(n8588) );
  OR2_X1 U10034 ( .A1(n9575), .A2(n8775), .ZN(n8587) );
  NAND2_X1 U10035 ( .A1(n8588), .A2(n8587), .ZN(n8594) );
  XNOR2_X1 U10036 ( .A(n8593), .B(n8594), .ZN(n8924) );
  INV_X1 U10037 ( .A(n8589), .ZN(n8590) );
  NAND2_X1 U10038 ( .A1(n8591), .A2(n8590), .ZN(n8921) );
  AND2_X1 U10039 ( .A1(n8924), .A2(n8921), .ZN(n8592) );
  INV_X1 U10040 ( .A(n8593), .ZN(n8595) );
  NAND2_X1 U10041 ( .A1(n8595), .A2(n8594), .ZN(n8596) );
  NAND2_X1 U10042 ( .A1(n9690), .A2(n4278), .ZN(n8598) );
  OR2_X1 U10043 ( .A1(n9684), .A2(n8779), .ZN(n8597) );
  NAND2_X1 U10044 ( .A1(n8598), .A2(n8597), .ZN(n8599) );
  XNOR2_X1 U10045 ( .A(n8599), .B(n4468), .ZN(n8600) );
  AOI22_X1 U10046 ( .A1(n9690), .A2(n4476), .B1(n9543), .B2(n8704), .ZN(n8601)
         );
  NAND2_X1 U10047 ( .A1(n8600), .A2(n8601), .ZN(n8822) );
  NAND2_X1 U10048 ( .A1(n8821), .A2(n8822), .ZN(n8826) );
  INV_X1 U10049 ( .A(n8600), .ZN(n8603) );
  INV_X1 U10050 ( .A(n8601), .ZN(n8602) );
  NAND2_X1 U10051 ( .A1(n8603), .A2(n8602), .ZN(n8823) );
  NAND2_X1 U10052 ( .A1(n9681), .A2(n4278), .ZN(n8605) );
  OR2_X1 U10053 ( .A1(n8830), .A2(n8779), .ZN(n8604) );
  NAND2_X1 U10054 ( .A1(n8605), .A2(n8604), .ZN(n8606) );
  XNOR2_X1 U10055 ( .A(n8606), .B(n4285), .ZN(n8900) );
  NAND2_X1 U10056 ( .A1(n9681), .A2(n4476), .ZN(n8608) );
  OR2_X1 U10057 ( .A1(n8830), .A2(n8775), .ZN(n8607) );
  NAND2_X1 U10058 ( .A1(n8608), .A2(n8607), .ZN(n8901) );
  NAND2_X1 U10059 ( .A1(n9523), .A2(n4278), .ZN(n8610) );
  OR2_X1 U10060 ( .A1(n9502), .A2(n8779), .ZN(n8609) );
  NAND2_X1 U10061 ( .A1(n8610), .A2(n8609), .ZN(n8611) );
  XNOR2_X1 U10062 ( .A(n8611), .B(n4468), .ZN(n8975) );
  NOR2_X1 U10063 ( .A1(n9502), .A2(n8775), .ZN(n8612) );
  AOI21_X1 U10064 ( .B1(n9523), .B2(n4476), .A(n8612), .ZN(n8632) );
  NAND2_X1 U10065 ( .A1(n9678), .A2(n4278), .ZN(n8614) );
  OR2_X1 U10066 ( .A1(n9519), .A2(n8779), .ZN(n8613) );
  NAND2_X1 U10067 ( .A1(n8614), .A2(n8613), .ZN(n8615) );
  XNOR2_X1 U10068 ( .A(n8615), .B(n4468), .ZN(n8722) );
  NOR2_X1 U10069 ( .A1(n9519), .A2(n8775), .ZN(n8616) );
  AOI21_X1 U10070 ( .B1(n9678), .B2(n4476), .A(n8616), .ZN(n8972) );
  AOI22_X1 U10071 ( .A1(n8975), .A2(n8632), .B1(n8722), .B2(n8972), .ZN(n8617)
         );
  NAND2_X1 U10072 ( .A1(n9506), .A2(n4278), .ZN(n8619) );
  NAND2_X1 U10073 ( .A1(n9220), .A2(n4476), .ZN(n8618) );
  NAND2_X1 U10074 ( .A1(n8619), .A2(n8618), .ZN(n8620) );
  XNOR2_X1 U10075 ( .A(n8620), .B(n4468), .ZN(n8622) );
  NOR2_X1 U10076 ( .A1(n9517), .A2(n8775), .ZN(n8621) );
  AOI21_X1 U10077 ( .B1(n9506), .B2(n4476), .A(n8621), .ZN(n8623) );
  NAND2_X1 U10078 ( .A1(n8622), .A2(n8623), .ZN(n8852) );
  INV_X1 U10079 ( .A(n8622), .ZN(n8625) );
  INV_X1 U10080 ( .A(n8623), .ZN(n8624) );
  NAND2_X1 U10081 ( .A1(n8625), .A2(n8624), .ZN(n8626) );
  NAND2_X1 U10082 ( .A1(n8852), .A2(n8626), .ZN(n8845) );
  NAND2_X1 U10083 ( .A1(n9664), .A2(n4278), .ZN(n8628) );
  OR2_X1 U10084 ( .A1(n9503), .A2(n8779), .ZN(n8627) );
  NAND2_X1 U10085 ( .A1(n8628), .A2(n8627), .ZN(n8629) );
  XNOR2_X1 U10086 ( .A(n8629), .B(n4285), .ZN(n8639) );
  NOR2_X1 U10087 ( .A1(n9503), .A2(n8775), .ZN(n8630) );
  AOI21_X1 U10088 ( .B1(n9664), .B2(n4476), .A(n8630), .ZN(n8640) );
  XNOR2_X1 U10089 ( .A(n8639), .B(n8640), .ZN(n8858) );
  INV_X1 U10090 ( .A(n8858), .ZN(n8638) );
  NOR2_X1 U10091 ( .A1(n8845), .A2(n8638), .ZN(n8636) );
  INV_X1 U10092 ( .A(n8975), .ZN(n8635) );
  INV_X1 U10093 ( .A(n8722), .ZN(n8968) );
  INV_X1 U10094 ( .A(n8972), .ZN(n8969) );
  NAND2_X1 U10095 ( .A1(n8968), .A2(n8969), .ZN(n8631) );
  NAND2_X1 U10096 ( .A1(n8631), .A2(n8632), .ZN(n8634) );
  INV_X1 U10097 ( .A(n8631), .ZN(n8633) );
  INV_X1 U10098 ( .A(n8632), .ZN(n8974) );
  AOI22_X1 U10099 ( .A1(n8635), .A2(n8634), .B1(n8633), .B2(n8974), .ZN(n8842)
         );
  AND2_X1 U10100 ( .A1(n8636), .A2(n8842), .ZN(n8637) );
  OR2_X1 U10101 ( .A1(n8638), .A2(n8852), .ZN(n8854) );
  INV_X1 U10102 ( .A(n8639), .ZN(n8641) );
  NAND2_X1 U10103 ( .A1(n8641), .A2(n8640), .ZN(n8642) );
  AND2_X1 U10104 ( .A1(n8854), .A2(n8642), .ZN(n8643) );
  NAND2_X1 U10105 ( .A1(n9651), .A2(n4278), .ZN(n8645) );
  OR2_X1 U10106 ( .A1(n9466), .A2(n8779), .ZN(n8644) );
  NAND2_X1 U10107 ( .A1(n8645), .A2(n8644), .ZN(n8646) );
  XNOR2_X1 U10108 ( .A(n8646), .B(n4285), .ZN(n8655) );
  NAND2_X1 U10109 ( .A1(n9651), .A2(n8774), .ZN(n8648) );
  OR2_X1 U10110 ( .A1(n9466), .A2(n8775), .ZN(n8647) );
  NAND2_X1 U10111 ( .A1(n8648), .A2(n8647), .ZN(n8656) );
  NAND2_X1 U10112 ( .A1(n8655), .A2(n8656), .ZN(n8766) );
  NAND2_X1 U10113 ( .A1(n9657), .A2(n4278), .ZN(n8650) );
  OR2_X1 U10114 ( .A1(n9485), .A2(n8779), .ZN(n8649) );
  NAND2_X1 U10115 ( .A1(n8650), .A2(n8649), .ZN(n8651) );
  XNOR2_X1 U10116 ( .A(n8651), .B(n4468), .ZN(n8763) );
  INV_X1 U10117 ( .A(n8763), .ZN(n8653) );
  NOR2_X1 U10118 ( .A1(n9485), .A2(n8775), .ZN(n8652) );
  AOI21_X1 U10119 ( .B1(n9657), .B2(n8774), .A(n8652), .ZN(n8935) );
  INV_X1 U10120 ( .A(n8935), .ZN(n8764) );
  NAND2_X1 U10121 ( .A1(n8653), .A2(n8764), .ZN(n8654) );
  AND2_X1 U10122 ( .A1(n8766), .A2(n8654), .ZN(n8661) );
  NAND3_X1 U10123 ( .A1(n8766), .A2(n8935), .A3(n8763), .ZN(n8659) );
  INV_X1 U10124 ( .A(n8655), .ZN(n8658) );
  INV_X1 U10125 ( .A(n8656), .ZN(n8657) );
  NAND2_X1 U10126 ( .A1(n8658), .A2(n8657), .ZN(n8765) );
  NAND2_X1 U10127 ( .A1(n8659), .A2(n8765), .ZN(n8660) );
  NAND2_X1 U10128 ( .A1(n9435), .A2(n4278), .ZN(n8663) );
  NAND2_X1 U10129 ( .A1(n9456), .A2(n8774), .ZN(n8662) );
  NAND2_X1 U10130 ( .A1(n8663), .A2(n8662), .ZN(n8664) );
  XNOR2_X1 U10131 ( .A(n8664), .B(n4468), .ZN(n8666) );
  NOR2_X1 U10132 ( .A1(n9638), .A2(n8775), .ZN(n8665) );
  AOI21_X1 U10133 ( .B1(n9435), .B2(n4476), .A(n8665), .ZN(n8667) );
  NAND2_X1 U10134 ( .A1(n8666), .A2(n8667), .ZN(n8890) );
  INV_X1 U10135 ( .A(n8666), .ZN(n8669) );
  INV_X1 U10136 ( .A(n8667), .ZN(n8668) );
  NAND2_X1 U10137 ( .A1(n8669), .A2(n8668), .ZN(n8891) );
  NAND2_X1 U10138 ( .A1(n9641), .A2(n4278), .ZN(n8671) );
  NAND2_X1 U10139 ( .A1(n9217), .A2(n4476), .ZN(n8670) );
  NAND2_X1 U10140 ( .A1(n8671), .A2(n8670), .ZN(n8672) );
  XNOR2_X1 U10141 ( .A(n8672), .B(n4285), .ZN(n8679) );
  NAND2_X1 U10142 ( .A1(n9641), .A2(n4476), .ZN(n8674) );
  NAND2_X1 U10143 ( .A1(n9217), .A2(n8704), .ZN(n8673) );
  NAND2_X1 U10144 ( .A1(n8674), .A2(n8673), .ZN(n8680) );
  AND2_X1 U10145 ( .A1(n8679), .A2(n8680), .ZN(n8812) );
  NAND2_X1 U10146 ( .A1(n9405), .A2(n4278), .ZN(n8676) );
  OR2_X1 U10147 ( .A1(n9626), .A2(n8779), .ZN(n8675) );
  NAND2_X1 U10148 ( .A1(n8676), .A2(n8675), .ZN(n8677) );
  XNOR2_X1 U10149 ( .A(n8677), .B(n4468), .ZN(n8912) );
  NOR2_X1 U10150 ( .A1(n9626), .A2(n8775), .ZN(n8678) );
  AOI21_X1 U10151 ( .B1(n9405), .B2(n8774), .A(n8678), .ZN(n8734) );
  INV_X1 U10152 ( .A(n8679), .ZN(n8682) );
  INV_X1 U10153 ( .A(n8680), .ZN(n8681) );
  OAI22_X1 U10154 ( .A1(n9722), .A2(n4463), .B1(n8916), .B2(n8711), .ZN(n8683)
         );
  XNOR2_X1 U10155 ( .A(n8683), .B(n4285), .ZN(n8737) );
  OR2_X1 U10156 ( .A1(n9722), .A2(n8779), .ZN(n8685) );
  NAND2_X1 U10157 ( .A1(n9393), .A2(n8704), .ZN(n8684) );
  NAND2_X1 U10158 ( .A1(n8685), .A2(n8684), .ZN(n8690) );
  NOR2_X1 U10159 ( .A1(n8737), .A2(n8690), .ZN(n8692) );
  AOI211_X1 U10160 ( .C1(n8912), .C2(n8734), .A(n8813), .B(n8692), .ZN(n8694)
         );
  OAI22_X1 U10161 ( .A1(n9718), .A2(n4463), .B1(n9350), .B2(n8711), .ZN(n8686)
         );
  XOR2_X1 U10162 ( .A(n4285), .B(n8686), .Z(n8688) );
  AOI22_X1 U10163 ( .A1(n9369), .A2(n4476), .B1(n8704), .B2(n9377), .ZN(n8687)
         );
  NAND2_X1 U10164 ( .A1(n8688), .A2(n8687), .ZN(n8695) );
  OAI21_X1 U10165 ( .B1(n8688), .B2(n8687), .A(n8695), .ZN(n8865) );
  INV_X1 U10166 ( .A(n8912), .ZN(n8733) );
  INV_X1 U10167 ( .A(n8734), .ZN(n8689) );
  NAND2_X1 U10168 ( .A1(n8733), .A2(n8689), .ZN(n8691) );
  INV_X1 U10169 ( .A(n8737), .ZN(n8740) );
  INV_X1 U10170 ( .A(n8690), .ZN(n8744) );
  OAI22_X1 U10171 ( .A1(n8692), .A2(n8691), .B1(n8740), .B2(n8744), .ZN(n8693)
         );
  INV_X1 U10172 ( .A(n8695), .ZN(n8696) );
  XNOR2_X1 U10173 ( .A(n8698), .B(n8697), .ZN(n8835) );
  NAND2_X1 U10174 ( .A1(n9342), .A2(n4278), .ZN(n8702) );
  NAND2_X1 U10175 ( .A1(n9216), .A2(n8774), .ZN(n8701) );
  NAND2_X1 U10176 ( .A1(n8702), .A2(n8701), .ZN(n8703) );
  XNOR2_X1 U10177 ( .A(n8703), .B(n4285), .ZN(n8708) );
  AND2_X1 U10178 ( .A1(n9216), .A2(n8704), .ZN(n8705) );
  AOI21_X1 U10179 ( .B1(n9342), .B2(n4476), .A(n8705), .ZN(n8706) );
  XNOR2_X1 U10180 ( .A(n8708), .B(n8706), .ZN(n8961) );
  INV_X1 U10181 ( .A(n8706), .ZN(n8707) );
  NAND2_X1 U10182 ( .A1(n8708), .A2(n8707), .ZN(n8715) );
  OAI22_X1 U10183 ( .A1(n9322), .A2(n4463), .B1(n8964), .B2(n8711), .ZN(n8710)
         );
  XNOR2_X1 U10184 ( .A(n8710), .B(n4285), .ZN(n8713) );
  OAI22_X1 U10185 ( .A1(n9322), .A2(n8711), .B1(n8964), .B2(n8775), .ZN(n8712)
         );
  NOR2_X1 U10186 ( .A1(n8713), .A2(n8712), .ZN(n8793) );
  AOI21_X1 U10187 ( .B1(n8713), .B2(n8712), .A(n8793), .ZN(n8714) );
  AOI21_X1 U10188 ( .B1(n8960), .B2(n8715), .A(n8714), .ZN(n8718) );
  INV_X1 U10189 ( .A(n8714), .ZN(n8717) );
  INV_X1 U10190 ( .A(n8715), .ZN(n8716) );
  AOI22_X1 U10191 ( .A1(n8978), .A2(n9216), .B1(P1_REG3_REG_27__SCAN_IN), .B2(
        P1_U3084), .ZN(n8719) );
  OAI21_X1 U10192 ( .B1(n9591), .B2(n8980), .A(n8719), .ZN(n8720) );
  AOI21_X1 U10193 ( .B1(n9320), .B2(n8984), .A(n8720), .ZN(n8721) );
  XNOR2_X1 U10194 ( .A(n8722), .B(n8969), .ZN(n8723) );
  XNOR2_X1 U10195 ( .A(n8970), .B(n8723), .ZN(n8730) );
  NAND2_X1 U10196 ( .A1(n8978), .A2(n9561), .ZN(n8725) );
  OAI211_X1 U10197 ( .C1(n9502), .C2(n8980), .A(n8725), .B(n8724), .ZN(n8726)
         );
  AOI21_X1 U10198 ( .B1(n8727), .B2(n8984), .A(n8726), .ZN(n8729) );
  NAND2_X1 U10199 ( .A1(n9678), .A2(n8941), .ZN(n8728) );
  OAI211_X1 U10200 ( .C1(n8730), .C2(n8986), .A(n8729), .B(n8728), .ZN(
        P1_U3213) );
  INV_X1 U10201 ( .A(n8813), .ZN(n8731) );
  NAND2_X1 U10202 ( .A1(n8736), .A2(n8731), .ZN(n8732) );
  NAND2_X1 U10203 ( .A1(n8732), .A2(n8734), .ZN(n8910) );
  AND2_X1 U10204 ( .A1(n8910), .A2(n8733), .ZN(n8738) );
  NOR2_X1 U10205 ( .A1(n8813), .A2(n8734), .ZN(n8735) );
  AND2_X1 U10206 ( .A1(n8736), .A2(n8735), .ZN(n8739) );
  OAI21_X1 U10207 ( .B1(n8738), .B2(n8739), .A(n8737), .ZN(n8745) );
  NAND2_X1 U10208 ( .A1(n8745), .A2(n8744), .ZN(n8866) );
  INV_X1 U10209 ( .A(n8738), .ZN(n8742) );
  INV_X1 U10210 ( .A(n8739), .ZN(n8911) );
  AND2_X1 U10211 ( .A1(n8911), .A2(n8740), .ZN(n8741) );
  NAND2_X1 U10212 ( .A1(n8742), .A2(n8741), .ZN(n8864) );
  INV_X1 U10213 ( .A(n8864), .ZN(n8743) );
  NOR2_X1 U10214 ( .A1(n8866), .A2(n8743), .ZN(n8747) );
  AOI21_X1 U10215 ( .B1(n8745), .B2(n8864), .A(n8744), .ZN(n8746) );
  OAI21_X1 U10216 ( .B1(n8747), .B2(n8746), .A(n8959), .ZN(n8752) );
  INV_X1 U10217 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n8748) );
  OAI22_X1 U10218 ( .A1(n8980), .A2(n9350), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8748), .ZN(n8750) );
  NOR2_X1 U10219 ( .A1(n9626), .A2(n8885), .ZN(n8749) );
  AOI211_X1 U10220 ( .C1(n8984), .C2(n9383), .A(n8750), .B(n8749), .ZN(n8751)
         );
  OAI211_X1 U10221 ( .C1(n9722), .C2(n8981), .A(n8752), .B(n8751), .ZN(
        P1_U3214) );
  OAI21_X1 U10222 ( .B1(n8754), .B2(n8753), .A(n8922), .ZN(n8755) );
  NAND2_X1 U10223 ( .A1(n8755), .A2(n8959), .ZN(n8761) );
  NAND2_X1 U10224 ( .A1(n8978), .A2(n9223), .ZN(n8757) );
  OAI211_X1 U10225 ( .C1(n9575), .C2(n8980), .A(n8757), .B(n8756), .ZN(n8758)
         );
  AOI21_X1 U10226 ( .B1(n8759), .B2(n8984), .A(n8758), .ZN(n8760) );
  OAI211_X1 U10227 ( .C1(n4952), .C2(n8981), .A(n8761), .B(n8760), .ZN(
        P1_U3215) );
  NAND2_X1 U10228 ( .A1(n8762), .A2(n8763), .ZN(n8933) );
  NOR2_X1 U10229 ( .A1(n8762), .A2(n8763), .ZN(n8932) );
  AOI21_X1 U10230 ( .B1(n8764), .B2(n8933), .A(n8932), .ZN(n8768) );
  NAND2_X1 U10231 ( .A1(n8766), .A2(n8765), .ZN(n8767) );
  XNOR2_X1 U10232 ( .A(n8768), .B(n8767), .ZN(n8773) );
  NAND2_X1 U10233 ( .A1(n8978), .A2(n9455), .ZN(n8769) );
  NAND2_X1 U10234 ( .A1(P1_U3084), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9288) );
  OAI211_X1 U10235 ( .C1(n9638), .C2(n8980), .A(n8769), .B(n9288), .ZN(n8771)
         );
  NOR2_X1 U10236 ( .A1(n9451), .A2(n8981), .ZN(n8770) );
  AOI211_X1 U10237 ( .C1(n8984), .C2(n9449), .A(n8771), .B(n8770), .ZN(n8772)
         );
  OAI21_X1 U10238 ( .B1(n8773), .B2(n8986), .A(n8772), .ZN(P1_U3217) );
  NAND2_X1 U10239 ( .A1(n8786), .A2(n8959), .ZN(n8785) );
  NAND2_X1 U10240 ( .A1(n9298), .A2(n8774), .ZN(n8777) );
  OR2_X1 U10241 ( .A1(n9591), .A2(n8775), .ZN(n8776) );
  NAND2_X1 U10242 ( .A1(n8777), .A2(n8776), .ZN(n8778) );
  XNOR2_X1 U10243 ( .A(n8778), .B(n4468), .ZN(n8783) );
  NOR2_X1 U10244 ( .A1(n9591), .A2(n8779), .ZN(n8780) );
  AOI21_X1 U10245 ( .B1(n9298), .B2(n4278), .A(n8780), .ZN(n8782) );
  XNOR2_X1 U10246 ( .A(n8783), .B(n8782), .ZN(n8784) );
  INV_X1 U10247 ( .A(n8784), .ZN(n8794) );
  NAND2_X1 U10248 ( .A1(n8785), .A2(n8794), .ZN(n8788) );
  INV_X1 U10249 ( .A(n9076), .ZN(n9215) );
  AOI22_X1 U10250 ( .A1(n8894), .A2(n9215), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3084), .ZN(n8789) );
  OAI21_X1 U10251 ( .B1(n8964), .B2(n8885), .A(n8789), .ZN(n8791) );
  NOR2_X1 U10252 ( .A1(n9590), .A2(n8981), .ZN(n8790) );
  AOI211_X1 U10253 ( .C1(n8792), .C2(n8984), .A(n8791), .B(n8790), .ZN(n8796)
         );
  NAND3_X1 U10254 ( .A1(n8794), .A2(n8793), .A3(n8959), .ZN(n8795) );
  AND2_X1 U10255 ( .A1(n8798), .A2(n8797), .ZN(n8799) );
  NAND2_X1 U10256 ( .A1(n8799), .A2(n8800), .ZN(n8873) );
  INV_X1 U10257 ( .A(n8799), .ZN(n8802) );
  INV_X1 U10258 ( .A(n8800), .ZN(n8801) );
  NAND2_X1 U10259 ( .A1(n8802), .A2(n8801), .ZN(n8875) );
  NAND2_X1 U10260 ( .A1(n8873), .A2(n8875), .ZN(n8803) );
  XOR2_X1 U10261 ( .A(n8876), .B(n8803), .Z(n8811) );
  NAND2_X1 U10262 ( .A1(n8978), .A2(n9225), .ZN(n8805) );
  OAI211_X1 U10263 ( .C1(n8806), .C2(n8980), .A(n8805), .B(n8804), .ZN(n8808)
         );
  NOR2_X1 U10264 ( .A1(n8981), .A2(n9953), .ZN(n8807) );
  AOI211_X1 U10265 ( .C1(n8984), .C2(n8809), .A(n8808), .B(n8807), .ZN(n8810)
         );
  OAI21_X1 U10266 ( .B1(n8811), .B2(n8986), .A(n8810), .ZN(P1_U3219) );
  NOR2_X1 U10267 ( .A1(n8813), .A2(n8812), .ZN(n8814) );
  XNOR2_X1 U10268 ( .A(n8815), .B(n8814), .ZN(n8820) );
  INV_X1 U10269 ( .A(n8984), .ZN(n8939) );
  NAND2_X1 U10270 ( .A1(n9421), .A2(n8894), .ZN(n8817) );
  AOI22_X1 U10271 ( .A1(n9456), .A2(n8978), .B1(P1_REG3_REG_21__SCAN_IN), .B2(
        P1_U3084), .ZN(n8816) );
  OAI211_X1 U10272 ( .C1(n8939), .C2(n9416), .A(n8817), .B(n8816), .ZN(n8818)
         );
  AOI21_X1 U10273 ( .B1(n9641), .B2(n8941), .A(n8818), .ZN(n8819) );
  OAI21_X1 U10274 ( .B1(n8820), .B2(n8986), .A(n8819), .ZN(P1_U3221) );
  INV_X1 U10275 ( .A(n8823), .ZN(n8827) );
  AOI21_X1 U10276 ( .B1(n8823), .B2(n8822), .A(n8821), .ZN(n8824) );
  NOR2_X1 U10277 ( .A1(n8824), .A2(n8986), .ZN(n8825) );
  OAI21_X1 U10278 ( .B1(n8827), .B2(n8826), .A(n8825), .ZN(n8833) );
  NAND2_X1 U10279 ( .A1(n8978), .A2(n9689), .ZN(n8829) );
  OAI211_X1 U10280 ( .C1(n8830), .C2(n8980), .A(n8829), .B(n8828), .ZN(n8831)
         );
  AOI21_X1 U10281 ( .B1(n9573), .B2(n8984), .A(n8831), .ZN(n8832) );
  OAI211_X1 U10282 ( .C1(n9571), .C2(n8981), .A(n8833), .B(n8832), .ZN(
        P1_U3222) );
  AOI21_X1 U10283 ( .B1(n8836), .B2(n8835), .A(n8834), .ZN(n8841) );
  AOI22_X1 U10284 ( .A1(n8894), .A2(n9216), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3084), .ZN(n8837) );
  OAI21_X1 U10285 ( .B1(n9350), .B2(n8885), .A(n8837), .ZN(n8839) );
  NOR2_X1 U10286 ( .A1(n9714), .A2(n8981), .ZN(n8838) );
  AOI211_X1 U10287 ( .C1(n8984), .C2(n9353), .A(n8839), .B(n8838), .ZN(n8840)
         );
  OAI21_X1 U10288 ( .B1(n8841), .B2(n8986), .A(n8840), .ZN(P1_U3223) );
  NAND2_X1 U10289 ( .A1(n8843), .A2(n8842), .ZN(n8846) );
  INV_X1 U10290 ( .A(n8853), .ZN(n8844) );
  AOI21_X1 U10291 ( .B1(n8846), .B2(n8845), .A(n8844), .ZN(n8851) );
  NAND2_X1 U10292 ( .A1(n8978), .A2(n9221), .ZN(n8847) );
  NAND2_X1 U10293 ( .A1(P1_U3084), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9838) );
  OAI211_X1 U10294 ( .C1(n9503), .C2(n8980), .A(n8847), .B(n9838), .ZN(n8849)
         );
  NOR2_X1 U10295 ( .A1(n9737), .A2(n8981), .ZN(n8848) );
  AOI211_X1 U10296 ( .C1(n8984), .C2(n9507), .A(n8849), .B(n8848), .ZN(n8850)
         );
  OAI21_X1 U10297 ( .B1(n8851), .B2(n8986), .A(n8850), .ZN(P1_U3224) );
  NAND2_X1 U10298 ( .A1(n8853), .A2(n8852), .ZN(n8857) );
  AND2_X1 U10299 ( .A1(n8855), .A2(n8854), .ZN(n8856) );
  OAI21_X1 U10300 ( .B1(n8858), .B2(n8857), .A(n8856), .ZN(n8859) );
  NAND2_X1 U10301 ( .A1(n8859), .A2(n8959), .ZN(n8863) );
  NAND2_X1 U10302 ( .A1(n8978), .A2(n9220), .ZN(n8860) );
  NAND2_X1 U10303 ( .A1(P1_U3084), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9856) );
  OAI211_X1 U10304 ( .C1(n9485), .C2(n8980), .A(n8860), .B(n9856), .ZN(n8861)
         );
  AOI21_X1 U10305 ( .B1(n9489), .B2(n8984), .A(n8861), .ZN(n8862) );
  OAI211_X1 U10306 ( .C1(n4949), .C2(n8981), .A(n8863), .B(n8862), .ZN(
        P1_U3226) );
  AND3_X1 U10307 ( .A1(n8866), .A2(n8865), .A3(n8864), .ZN(n8868) );
  OAI21_X1 U10308 ( .B1(n8868), .B2(n8867), .A(n8959), .ZN(n8872) );
  AOI22_X1 U10309 ( .A1(n8894), .A2(n9364), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3084), .ZN(n8869) );
  OAI21_X1 U10310 ( .B1(n8916), .B2(n8885), .A(n8869), .ZN(n8870) );
  AOI21_X1 U10311 ( .B1(n9370), .B2(n8984), .A(n8870), .ZN(n8871) );
  OAI211_X1 U10312 ( .C1(n9718), .C2(n8981), .A(n8872), .B(n8871), .ZN(
        P1_U3227) );
  INV_X1 U10313 ( .A(n8873), .ZN(n8874) );
  AOI21_X1 U10314 ( .B1(n8876), .B2(n8875), .A(n8874), .ZN(n8880) );
  INV_X1 U10315 ( .A(n8877), .ZN(n8879) );
  OAI21_X1 U10316 ( .B1(n8880), .B2(n8879), .A(n8878), .ZN(n8881) );
  NAND2_X1 U10317 ( .A1(n8881), .A2(n8959), .ZN(n8889) );
  AOI21_X1 U10318 ( .B1(n8894), .B2(n9222), .A(n8882), .ZN(n8883) );
  OAI21_X1 U10319 ( .B1(n8885), .B2(n8884), .A(n8883), .ZN(n8886) );
  AOI21_X1 U10320 ( .B1(n8887), .B2(n8984), .A(n8886), .ZN(n8888) );
  OAI211_X1 U10321 ( .C1(n9962), .C2(n8981), .A(n8889), .B(n8888), .ZN(
        P1_U3229) );
  NAND2_X1 U10322 ( .A1(n8891), .A2(n8890), .ZN(n8893) );
  XOR2_X1 U10323 ( .A(n8893), .B(n8892), .Z(n8899) );
  NAND2_X1 U10324 ( .A1(n9217), .A2(n8894), .ZN(n8896) );
  AOI22_X1 U10325 ( .A1(n9218), .A2(n8978), .B1(P1_REG3_REG_20__SCAN_IN), .B2(
        P1_U3084), .ZN(n8895) );
  OAI211_X1 U10326 ( .C1(n8939), .C2(n9432), .A(n8896), .B(n8895), .ZN(n8897)
         );
  AOI21_X1 U10327 ( .B1(n9435), .B2(n8941), .A(n8897), .ZN(n8898) );
  OAI21_X1 U10328 ( .B1(n8899), .B2(n8986), .A(n8898), .ZN(P1_U3231) );
  XOR2_X1 U10329 ( .A(n8901), .B(n8900), .Z(n8902) );
  XNOR2_X1 U10330 ( .A(n4490), .B(n8902), .ZN(n8909) );
  NOR2_X1 U10331 ( .A1(n8904), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9819) );
  AOI21_X1 U10332 ( .B1(n8978), .B2(n9543), .A(n9819), .ZN(n8906) );
  NAND2_X1 U10333 ( .A1(n8984), .A2(n9537), .ZN(n8905) );
  OAI211_X1 U10334 ( .C1(n9519), .C2(n8980), .A(n8906), .B(n8905), .ZN(n8907)
         );
  AOI21_X1 U10335 ( .B1(n8941), .B2(n9681), .A(n8907), .ZN(n8908) );
  OAI21_X1 U10336 ( .B1(n8909), .B2(n8986), .A(n8908), .ZN(P1_U3232) );
  NAND2_X1 U10337 ( .A1(n8911), .A2(n8910), .ZN(n8913) );
  XNOR2_X1 U10338 ( .A(n8913), .B(n8912), .ZN(n8919) );
  AOI22_X1 U10339 ( .A1(n9217), .A2(n8978), .B1(P1_REG3_REG_22__SCAN_IN), .B2(
        P1_U3084), .ZN(n8915) );
  NAND2_X1 U10340 ( .A1(n9398), .A2(n8984), .ZN(n8914) );
  OAI211_X1 U10341 ( .C1(n8916), .C2(n8980), .A(n8915), .B(n8914), .ZN(n8917)
         );
  AOI21_X1 U10342 ( .B1(n9405), .B2(n8941), .A(n8917), .ZN(n8918) );
  OAI21_X1 U10343 ( .B1(n8919), .B2(n8986), .A(n8918), .ZN(P1_U3233) );
  AND2_X1 U10344 ( .A1(n8922), .A2(n8921), .ZN(n8925) );
  OAI211_X1 U10345 ( .C1(n8925), .C2(n8924), .A(n8959), .B(n8923), .ZN(n8931)
         );
  NAND2_X1 U10346 ( .A1(n8978), .A2(n9222), .ZN(n8927) );
  OAI211_X1 U10347 ( .C1(n9684), .C2(n8980), .A(n8927), .B(n8926), .ZN(n8928)
         );
  AOI21_X1 U10348 ( .B1(n8929), .B2(n8984), .A(n8928), .ZN(n8930) );
  OAI211_X1 U10349 ( .C1(n4951), .C2(n8981), .A(n8931), .B(n8930), .ZN(
        P1_U3234) );
  INV_X1 U10350 ( .A(n8932), .ZN(n8934) );
  NAND2_X1 U10351 ( .A1(n8934), .A2(n8933), .ZN(n8936) );
  XNOR2_X1 U10352 ( .A(n8936), .B(n8935), .ZN(n8943) );
  NAND2_X1 U10353 ( .A1(P1_U3084), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9259) );
  OAI21_X1 U10354 ( .B1(n9466), .B2(n8980), .A(n9259), .ZN(n8937) );
  AOI21_X1 U10355 ( .B1(n8978), .B2(n9219), .A(n8937), .ZN(n8938) );
  OAI21_X1 U10356 ( .B1(n9467), .B2(n8939), .A(n8938), .ZN(n8940) );
  AOI21_X1 U10357 ( .B1(n9657), .B2(n8941), .A(n8940), .ZN(n8942) );
  OAI21_X1 U10358 ( .B1(n8943), .B2(n8986), .A(n8942), .ZN(P1_U3236) );
  NAND2_X1 U10359 ( .A1(n8944), .A2(n9913), .ZN(n9934) );
  INV_X1 U10360 ( .A(n8945), .ZN(n8946) );
  AND3_X1 U10361 ( .A1(n8948), .A2(n8947), .A3(n8946), .ZN(n8950) );
  OAI21_X1 U10362 ( .B1(n8950), .B2(n8949), .A(n8959), .ZN(n8957) );
  NAND2_X1 U10363 ( .A1(n8978), .A2(n9227), .ZN(n8952) );
  OAI211_X1 U10364 ( .C1(n8953), .C2(n8980), .A(n8952), .B(n8951), .ZN(n8954)
         );
  AOI21_X1 U10365 ( .B1(n8955), .B2(n8984), .A(n8954), .ZN(n8956) );
  OAI211_X1 U10366 ( .C1(n8958), .C2(n9934), .A(n8957), .B(n8956), .ZN(
        P1_U3237) );
  OAI211_X1 U10367 ( .C1(n8962), .C2(n8961), .A(n8960), .B(n8959), .ZN(n8967)
         );
  AOI22_X1 U10368 ( .A1(n8978), .A2(n9364), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3084), .ZN(n8963) );
  OAI21_X1 U10369 ( .B1(n8964), .B2(n8980), .A(n8963), .ZN(n8965) );
  AOI21_X1 U10370 ( .B1(n9337), .B2(n8984), .A(n8965), .ZN(n8966) );
  OAI211_X1 U10371 ( .C1(n4945), .C2(n8981), .A(n8967), .B(n8966), .ZN(
        P1_U3238) );
  INV_X1 U10372 ( .A(n8970), .ZN(n8973) );
  OAI21_X1 U10373 ( .B1(n8970), .B2(n8969), .A(n8968), .ZN(n8971) );
  OAI21_X1 U10374 ( .B1(n8973), .B2(n8972), .A(n8971), .ZN(n8977) );
  XNOR2_X1 U10375 ( .A(n8975), .B(n8974), .ZN(n8976) );
  XNOR2_X1 U10376 ( .A(n8977), .B(n8976), .ZN(n8987) );
  NAND2_X1 U10377 ( .A1(n8978), .A2(n9553), .ZN(n8979) );
  NAND2_X1 U10378 ( .A1(P1_U3084), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9826) );
  OAI211_X1 U10379 ( .C1(n9517), .C2(n8980), .A(n8979), .B(n9826), .ZN(n8983)
         );
  NOR2_X1 U10380 ( .A1(n9741), .A2(n8981), .ZN(n8982) );
  AOI211_X1 U10381 ( .C1(n8984), .C2(n9524), .A(n8983), .B(n8982), .ZN(n8985)
         );
  OAI21_X1 U10382 ( .B1(n8987), .B2(n8986), .A(n8985), .ZN(P1_U3239) );
  NAND2_X1 U10383 ( .A1(n8989), .A2(n8988), .ZN(n8990) );
  NOR4_X1 U10384 ( .A1(n8992), .A2(n8991), .A3(n8990), .A4(n9806), .ZN(n9213)
         );
  OAI21_X1 U10385 ( .B1(n9118), .B2(n9203), .A(P1_B_REG_SCAN_IN), .ZN(n9212)
         );
  NAND2_X1 U10386 ( .A1(n8993), .A2(n9119), .ZN(n9077) );
  NAND2_X1 U10387 ( .A1(n8994), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n8998) );
  NAND2_X1 U10388 ( .A1(n5747), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n8997) );
  NAND2_X1 U10389 ( .A1(n8995), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n8996) );
  AND3_X1 U10390 ( .A1(n8998), .A2(n8997), .A3(n8996), .ZN(n9311) );
  INV_X1 U10391 ( .A(n9311), .ZN(n9214) );
  AOI21_X1 U10392 ( .B1(n9214), .B2(n9114), .A(n9705), .ZN(n9082) );
  INV_X1 U10393 ( .A(n9079), .ZN(n9001) );
  OAI21_X1 U10394 ( .B1(n9082), .B2(n9185), .A(n9001), .ZN(n9084) );
  AND2_X1 U10395 ( .A1(n9050), .A2(n9085), .ZN(n9173) );
  INV_X1 U10396 ( .A(n9173), .ZN(n9003) );
  INV_X1 U10397 ( .A(n9179), .ZN(n9002) );
  AOI21_X1 U10398 ( .B1(n9177), .B2(n9003), .A(n9002), .ZN(n9054) );
  INV_X1 U10399 ( .A(n9013), .ZN(n9006) );
  OAI211_X1 U10400 ( .C1(n9006), .C2(n9005), .A(n9133), .B(n9004), .ZN(n9007)
         );
  AND2_X1 U10401 ( .A1(n9017), .A2(n9019), .ZN(n9141) );
  NAND2_X1 U10402 ( .A1(n9007), .A2(n9141), .ZN(n9009) );
  INV_X1 U10403 ( .A(n9139), .ZN(n9008) );
  NAND2_X1 U10404 ( .A1(n9011), .A2(n9010), .ZN(n9024) );
  INV_X1 U10405 ( .A(n9014), .ZN(n9016) );
  INV_X1 U10406 ( .A(n9133), .ZN(n9015) );
  AOI211_X1 U10407 ( .C1(n9018), .C2(n9017), .A(n9016), .B(n9015), .ZN(n9022)
         );
  INV_X1 U10408 ( .A(n9019), .ZN(n9021) );
  AOI21_X1 U10409 ( .B1(n9025), .B2(n9024), .A(n9023), .ZN(n9026) );
  OAI21_X1 U10410 ( .B1(n9032), .B2(n9028), .A(n9547), .ZN(n9030) );
  NAND2_X1 U10411 ( .A1(n9036), .A2(n9029), .ZN(n9149) );
  AOI211_X1 U10412 ( .C1(n9030), .C2(n9548), .A(n4671), .B(n9149), .ZN(n9031)
         );
  XNOR2_X1 U10413 ( .A(n9523), .B(n9502), .ZN(n9107) );
  NOR2_X1 U10414 ( .A1(n9031), .A2(n9107), .ZN(n9041) );
  OAI21_X1 U10415 ( .B1(n9033), .B2(n9684), .A(n9690), .ZN(n9034) );
  OAI211_X1 U10416 ( .C1(n9138), .C2(n9543), .A(n9151), .B(n9034), .ZN(n9035)
         );
  NAND2_X1 U10417 ( .A1(n9152), .A2(n9151), .ZN(n9137) );
  NAND2_X1 U10418 ( .A1(n9137), .A2(n9036), .ZN(n9037) );
  MUX2_X1 U10419 ( .A(n9038), .B(n9037), .S(n9077), .Z(n9040) );
  INV_X1 U10420 ( .A(n9153), .ZN(n9143) );
  MUX2_X1 U10421 ( .A(n9143), .B(n9154), .S(n9077), .Z(n9039) );
  INV_X1 U10422 ( .A(n9155), .ZN(n9043) );
  MUX2_X1 U10423 ( .A(n9043), .B(n9042), .S(n9077), .Z(n9044) );
  NAND2_X1 U10424 ( .A1(n9160), .A2(n9158), .ZN(n9047) );
  NAND2_X1 U10425 ( .A1(n9056), .A2(n9046), .ZN(n9129) );
  MUX2_X1 U10426 ( .A(n9047), .B(n9129), .S(n9077), .Z(n9048) );
  AND2_X1 U10427 ( .A1(n9089), .A2(n9055), .ZN(n9049) );
  NAND2_X1 U10428 ( .A1(n9061), .A2(n9049), .ZN(n9167) );
  OAI211_X1 U10429 ( .C1(n4748), .C2(n9088), .A(n9087), .B(n9060), .ZN(n9169)
         );
  OAI211_X1 U10430 ( .C1(n4525), .C2(n4529), .A(n9176), .B(n9177), .ZN(n9051)
         );
  AOI21_X1 U10431 ( .B1(n9052), .B2(n9173), .A(n9051), .ZN(n9053) );
  NOR2_X1 U10432 ( .A1(n9179), .A2(n4671), .ZN(n9067) );
  NAND3_X1 U10433 ( .A1(n9057), .A2(n9056), .A3(n9055), .ZN(n9059) );
  AOI21_X1 U10434 ( .B1(n9059), .B2(n9058), .A(n4749), .ZN(n9063) );
  INV_X1 U10435 ( .A(n9060), .ZN(n9062) );
  OAI211_X1 U10436 ( .C1(n9063), .C2(n9062), .A(n9061), .B(n9170), .ZN(n9064)
         );
  NAND2_X1 U10437 ( .A1(n9064), .A2(n9087), .ZN(n9065) );
  NAND4_X1 U10438 ( .A1(n9065), .A2(n4671), .A3(n9177), .A4(n4529), .ZN(n9066)
         );
  OR2_X1 U10439 ( .A1(n9342), .A2(n9349), .ZN(n9182) );
  MUX2_X1 U10440 ( .A(n9127), .B(n9182), .S(n9077), .Z(n9068) );
  MUX2_X1 U10441 ( .A(n9070), .B(n9126), .S(n9077), .Z(n9071) );
  NAND3_X1 U10442 ( .A1(n9072), .A2(n9113), .A3(n9071), .ZN(n9075) );
  XNOR2_X1 U10443 ( .A(n9303), .B(n9215), .ZN(n9074) );
  MUX2_X1 U10444 ( .A(n9307), .B(n9184), .S(n9077), .Z(n9073) );
  NAND2_X1 U10445 ( .A1(n9303), .A2(n9076), .ZN(n9189) );
  INV_X1 U10446 ( .A(n9189), .ZN(n9078) );
  NAND2_X1 U10447 ( .A1(n9078), .A2(n9077), .ZN(n9080) );
  NOR2_X1 U10448 ( .A1(n9081), .A2(n4671), .ZN(n9083) );
  INV_X1 U10449 ( .A(n9598), .ZN(n9588) );
  INV_X1 U10450 ( .A(n9085), .ZN(n9086) );
  NOR2_X1 U10451 ( .A1(n9172), .A2(n9086), .ZN(n9381) );
  NAND2_X1 U10452 ( .A1(n9089), .A2(n9088), .ZN(n9437) );
  NOR4_X1 U10453 ( .A1(n9093), .A2(n9092), .A3(n9091), .A4(n9090), .ZN(n9097)
         );
  INV_X1 U10454 ( .A(n9101), .ZN(n9102) );
  NOR4_X1 U10455 ( .A1(n9500), .A2(n9106), .A3(n9105), .A4(n9104), .ZN(n9109)
         );
  INV_X1 U10456 ( .A(n9482), .ZN(n9108) );
  INV_X1 U10457 ( .A(n9107), .ZN(n9529) );
  NAND4_X1 U10458 ( .A1(n9109), .A2(n9470), .A3(n9108), .A4(n9529), .ZN(n9110)
         );
  NOR4_X1 U10459 ( .A1(n9419), .A2(n9437), .A3(n4541), .A4(n9110), .ZN(n9111)
         );
  NOR2_X1 U10460 ( .A1(n9115), .A2(n4612), .ZN(n9200) );
  NOR2_X1 U10461 ( .A1(n9705), .A2(n9214), .ZN(n9125) );
  NAND2_X1 U10462 ( .A1(n9195), .A2(n5662), .ZN(n9124) );
  OR2_X1 U10463 ( .A1(n9120), .A2(n9418), .ZN(n9201) );
  INV_X1 U10464 ( .A(n9201), .ZN(n9117) );
  OAI211_X1 U10465 ( .C1(n9118), .C2(n5662), .A(n9124), .B(n9117), .ZN(n9209)
         );
  NOR2_X1 U10466 ( .A1(n9120), .A2(n9119), .ZN(n9196) );
  NAND2_X1 U10467 ( .A1(n4480), .A2(n9196), .ZN(n9122) );
  OAI22_X1 U10468 ( .A1(n9200), .A2(n9122), .B1(n9121), .B2(n9201), .ZN(n9123)
         );
  NAND3_X1 U10469 ( .A1(n9210), .A2(n9124), .A3(n9123), .ZN(n9208) );
  INV_X1 U10470 ( .A(n9125), .ZN(n9190) );
  OAI211_X1 U10471 ( .C1(n9128), .C2(n9127), .A(n9307), .B(n9126), .ZN(n9187)
         );
  INV_X1 U10472 ( .A(n9129), .ZN(n9165) );
  AOI21_X1 U10473 ( .B1(n9231), .B2(n9889), .A(n5662), .ZN(n9131) );
  AND3_X1 U10474 ( .A1(n9132), .A2(n9131), .A3(n9130), .ZN(n9135) );
  OAI211_X1 U10475 ( .C1(n9136), .C2(n9135), .A(n9134), .B(n9133), .ZN(n9142)
         );
  INV_X1 U10476 ( .A(n9137), .ZN(n9140) );
  AND3_X1 U10477 ( .A1(n9139), .A2(n9138), .A3(n9548), .ZN(n9145) );
  NAND4_X1 U10478 ( .A1(n9142), .A2(n9141), .A3(n9140), .A4(n9145), .ZN(n9144)
         );
  NOR2_X1 U10479 ( .A1(n9144), .A2(n9143), .ZN(n9163) );
  INV_X1 U10480 ( .A(n9145), .ZN(n9148) );
  INV_X1 U10481 ( .A(n9548), .ZN(n9146) );
  OAI22_X1 U10482 ( .A1(n9148), .A2(n9147), .B1(n9547), .B2(n9146), .ZN(n9150)
         );
  AOI21_X1 U10483 ( .B1(n9151), .B2(n9150), .A(n9149), .ZN(n9157) );
  NAND2_X1 U10484 ( .A1(n9153), .A2(n9152), .ZN(n9156) );
  OAI211_X1 U10485 ( .C1(n9157), .C2(n9156), .A(n9155), .B(n5639), .ZN(n9162)
         );
  AND2_X1 U10486 ( .A1(n9158), .A2(n9481), .ZN(n9159) );
  AND2_X1 U10487 ( .A1(n9160), .A2(n9159), .ZN(n9161) );
  OAI211_X1 U10488 ( .C1(n9163), .C2(n9162), .A(n9436), .B(n9161), .ZN(n9164)
         );
  OAI21_X1 U10489 ( .B1(n4364), .B2(n9165), .A(n9164), .ZN(n9166) );
  NOR2_X1 U10490 ( .A1(n9167), .A2(n9166), .ZN(n9168) );
  NOR2_X1 U10491 ( .A1(n9169), .A2(n9168), .ZN(n9175) );
  INV_X1 U10492 ( .A(n9170), .ZN(n9171) );
  OR2_X1 U10493 ( .A1(n9172), .A2(n9171), .ZN(n9174) );
  OAI21_X1 U10494 ( .B1(n9175), .B2(n9174), .A(n9173), .ZN(n9178) );
  NAND3_X1 U10495 ( .A1(n9178), .A2(n9177), .A3(n9176), .ZN(n9180) );
  NAND2_X1 U10496 ( .A1(n9180), .A2(n9179), .ZN(n9181) );
  NAND2_X1 U10497 ( .A1(n9182), .A2(n9181), .ZN(n9183) );
  NOR2_X1 U10498 ( .A1(n9323), .A2(n9183), .ZN(n9186) );
  OAI211_X1 U10499 ( .C1(n9187), .C2(n9186), .A(n9185), .B(n9184), .ZN(n9188)
         );
  NAND3_X1 U10500 ( .A1(n9190), .A2(n9189), .A3(n9188), .ZN(n9191) );
  MUX2_X1 U10501 ( .A(n9869), .B(n9194), .S(n9193), .Z(n9206) );
  INV_X1 U10502 ( .A(n9196), .ZN(n9197) );
  NOR3_X1 U10503 ( .A1(n9199), .A2(n4480), .A3(n9197), .ZN(n9205) );
  INV_X1 U10504 ( .A(n9200), .ZN(n9202) );
  NOR3_X1 U10505 ( .A1(n9202), .A2(n5662), .A3(n9201), .ZN(n9204) );
  OAI211_X1 U10506 ( .C1(n9210), .C2(n9209), .A(n9208), .B(n9207), .ZN(n9211)
         );
  OAI21_X1 U10507 ( .B1(n9213), .B2(n9212), .A(n9211), .ZN(P1_U3240) );
  MUX2_X1 U10508 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9214), .S(P1_U4006), .Z(
        P1_U3585) );
  MUX2_X1 U10509 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n9215), .S(P1_U4006), .Z(
        P1_U3584) );
  INV_X1 U10510 ( .A(n9591), .ZN(n9304) );
  MUX2_X1 U10511 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9304), .S(P1_U4006), .Z(
        P1_U3583) );
  MUX2_X1 U10512 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9333), .S(P1_U4006), .Z(
        P1_U3582) );
  MUX2_X1 U10513 ( .A(n9216), .B(P1_DATAO_REG_26__SCAN_IN), .S(n9230), .Z(
        P1_U3581) );
  MUX2_X1 U10514 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9364), .S(P1_U4006), .Z(
        P1_U3580) );
  MUX2_X1 U10515 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9377), .S(P1_U4006), .Z(
        P1_U3579) );
  MUX2_X1 U10516 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9393), .S(P1_U4006), .Z(
        P1_U3578) );
  MUX2_X1 U10517 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9421), .S(P1_U4006), .Z(
        P1_U3577) );
  MUX2_X1 U10518 ( .A(n9217), .B(P1_DATAO_REG_21__SCAN_IN), .S(n9230), .Z(
        P1_U3576) );
  MUX2_X1 U10519 ( .A(n9456), .B(P1_DATAO_REG_20__SCAN_IN), .S(n9230), .Z(
        P1_U3575) );
  MUX2_X1 U10520 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9218), .S(P1_U4006), .Z(
        P1_U3574) );
  MUX2_X1 U10521 ( .A(n9455), .B(P1_DATAO_REG_18__SCAN_IN), .S(n9230), .Z(
        P1_U3573) );
  MUX2_X1 U10522 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9219), .S(P1_U4006), .Z(
        P1_U3572) );
  MUX2_X1 U10523 ( .A(n9220), .B(P1_DATAO_REG_16__SCAN_IN), .S(n9230), .Z(
        P1_U3571) );
  MUX2_X1 U10524 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n9221), .S(P1_U4006), .Z(
        P1_U3570) );
  MUX2_X1 U10525 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n9553), .S(P1_U4006), .Z(
        P1_U3569) );
  MUX2_X1 U10526 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9561), .S(P1_U4006), .Z(
        P1_U3568) );
  MUX2_X1 U10527 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n9543), .S(P1_U4006), .Z(
        P1_U3567) );
  MUX2_X1 U10528 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n9689), .S(P1_U4006), .Z(
        P1_U3566) );
  MUX2_X1 U10529 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n9222), .S(P1_U4006), .Z(
        P1_U3565) );
  MUX2_X1 U10530 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n9223), .S(P1_U4006), .Z(
        P1_U3564) );
  MUX2_X1 U10531 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n9224), .S(P1_U4006), .Z(
        P1_U3563) );
  MUX2_X1 U10532 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n9225), .S(P1_U4006), .Z(
        P1_U3562) );
  MUX2_X1 U10533 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n9226), .S(P1_U4006), .Z(
        P1_U3561) );
  MUX2_X1 U10534 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n9227), .S(P1_U4006), .Z(
        P1_U3560) );
  MUX2_X1 U10535 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n9228), .S(P1_U4006), .Z(
        P1_U3559) );
  MUX2_X1 U10536 ( .A(n9915), .B(P1_DATAO_REG_3__SCAN_IN), .S(n9230), .Z(
        P1_U3558) );
  MUX2_X1 U10537 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n9229), .S(P1_U4006), .Z(
        P1_U3557) );
  MUX2_X1 U10538 ( .A(n9231), .B(P1_DATAO_REG_1__SCAN_IN), .S(n9230), .Z(
        P1_U3556) );
  MUX2_X1 U10539 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n4453), .S(P1_U4006), .Z(
        P1_U3555) );
  OAI21_X1 U10540 ( .B1(n9234), .B2(n9233), .A(n9232), .ZN(n9236) );
  OAI22_X1 U10541 ( .A1(n9281), .A2(n9236), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9235), .ZN(n9237) );
  AOI21_X1 U10542 ( .B1(n4479), .B2(n4477), .A(n9237), .ZN(n9244) );
  NAND2_X1 U10543 ( .A1(n9810), .A2(P1_ADDR_REG_2__SCAN_IN), .ZN(n9243) );
  OAI211_X1 U10544 ( .C1(n9241), .C2(n9240), .A(n9855), .B(n9239), .ZN(n9242)
         );
  NAND4_X1 U10545 ( .A1(n9245), .A2(n9244), .A3(n9243), .A4(n9242), .ZN(
        P1_U3243) );
  INV_X1 U10546 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n9468) );
  OR2_X1 U10547 ( .A1(n9276), .A2(n9468), .ZN(n9247) );
  NAND2_X1 U10548 ( .A1(n9276), .A2(n9468), .ZN(n9246) );
  AND2_X1 U10549 ( .A1(n9247), .A2(n9246), .ZN(n9257) );
  NAND2_X1 U10550 ( .A1(n9248), .A2(n9263), .ZN(n9250) );
  INV_X1 U10551 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n9828) );
  NAND2_X1 U10552 ( .A1(n9844), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n9253) );
  OAI21_X1 U10553 ( .B1(n9844), .B2(P1_REG2_REG_16__SCAN_IN), .A(n9253), .ZN(
        n9841) );
  NAND2_X1 U10554 ( .A1(P1_REG2_REG_17__SCAN_IN), .A2(n9255), .ZN(n9254) );
  OAI21_X1 U10555 ( .B1(n9255), .B2(P1_REG2_REG_17__SCAN_IN), .A(n9254), .ZN(
        n9852) );
  AOI21_X1 U10556 ( .B1(n9257), .B2(n9256), .A(n9275), .ZN(n9258) );
  NAND2_X1 U10557 ( .A1(n9855), .A2(n9258), .ZN(n9260) );
  OAI211_X1 U10558 ( .C1(n9859), .C2(n9279), .A(n9260), .B(n9259), .ZN(n9273)
         );
  INV_X1 U10559 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9278) );
  AOI22_X1 U10560 ( .A1(P1_REG1_REG_18__SCAN_IN), .A2(n9279), .B1(n9276), .B2(
        n9278), .ZN(n9270) );
  INV_X1 U10561 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n9268) );
  XNOR2_X1 U10562 ( .A(n9858), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n9864) );
  INV_X1 U10563 ( .A(n9844), .ZN(n9267) );
  INV_X1 U10564 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n10240) );
  XNOR2_X1 U10565 ( .A(n9844), .B(n10240), .ZN(n9846) );
  NAND2_X1 U10566 ( .A1(n9832), .A2(n9265), .ZN(n9266) );
  XNOR2_X1 U10567 ( .A(n9265), .B(n9264), .ZN(n9834) );
  NAND2_X1 U10568 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(n9834), .ZN(n9833) );
  NAND2_X1 U10569 ( .A1(n9266), .A2(n9833), .ZN(n9847) );
  OAI21_X1 U10570 ( .B1(n9858), .B2(n9268), .A(n9861), .ZN(n9269) );
  AOI21_X1 U10571 ( .B1(n9270), .B2(n9269), .A(n9277), .ZN(n9271) );
  NOR2_X1 U10572 ( .A1(n9271), .A2(n9281), .ZN(n9272) );
  AOI211_X1 U10573 ( .C1(n9810), .C2(P1_ADDR_REG_18__SCAN_IN), .A(n9273), .B(
        n9272), .ZN(n9274) );
  INV_X1 U10574 ( .A(n9274), .ZN(P1_U3259) );
  XOR2_X1 U10575 ( .A(n9280), .B(P1_REG1_REG_19__SCAN_IN), .Z(n9284) );
  AOI22_X1 U10576 ( .A1(n9285), .A2(n9855), .B1(n9862), .B2(n9284), .ZN(n9286)
         );
  NAND2_X1 U10577 ( .A1(n9289), .A2(n9528), .ZN(n9292) );
  INV_X1 U10578 ( .A(n9584), .ZN(n9290) );
  NOR2_X1 U10579 ( .A1(n9877), .A2(n9290), .ZN(n9295) );
  AOI21_X1 U10580 ( .B1(n9877), .B2(P1_REG2_REG_31__SCAN_IN), .A(n9295), .ZN(
        n9291) );
  OAI211_X1 U10581 ( .C1(n9293), .C2(n9526), .A(n9292), .B(n9291), .ZN(
        P1_U3261) );
  INV_X1 U10582 ( .A(n9301), .ZN(n9294) );
  AOI211_X2 U10583 ( .C1(n8999), .C2(n9294), .A(n9535), .B(n4326), .ZN(n9585)
         );
  NAND2_X1 U10584 ( .A1(n9585), .A2(n9528), .ZN(n9297) );
  AOI21_X1 U10585 ( .B1(n9877), .B2(P1_REG2_REG_30__SCAN_IN), .A(n9295), .ZN(
        n9296) );
  OAI211_X1 U10586 ( .C1(n9705), .C2(n9526), .A(n9297), .B(n9296), .ZN(
        P1_U3262) );
  NAND2_X1 U10587 ( .A1(n9298), .A2(n9304), .ZN(n9597) );
  XNOR2_X1 U10588 ( .A(n9300), .B(n9598), .ZN(n9317) );
  AOI211_X1 U10589 ( .C1(n9303), .C2(n9302), .A(n9535), .B(n9301), .ZN(n9595)
         );
  AOI22_X1 U10590 ( .A1(n9544), .A2(n9304), .B1(n9877), .B2(
        P1_REG2_REG_29__SCAN_IN), .ZN(n9305) );
  OAI21_X1 U10591 ( .B1(n4943), .B2(n9526), .A(n9305), .ZN(n9306) );
  AOI21_X1 U10592 ( .B1(n9595), .B2(n9528), .A(n9306), .ZN(n9316) );
  NAND2_X1 U10593 ( .A1(n9308), .A2(n9307), .ZN(n9309) );
  NOR2_X1 U10594 ( .A1(n9538), .A2(n9313), .ZN(n9314) );
  OAI21_X1 U10595 ( .B1(n9599), .B2(n9314), .A(n9541), .ZN(n9315) );
  OAI211_X1 U10596 ( .C1(n9317), .C2(n9513), .A(n9316), .B(n9315), .ZN(
        P1_U3355) );
  XNOR2_X1 U10597 ( .A(n9318), .B(n9323), .ZN(n9606) );
  AOI211_X1 U10598 ( .C1(n9603), .C2(n9339), .A(n9535), .B(n9319), .ZN(n9602)
         );
  AOI22_X1 U10599 ( .A1(n9877), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n9320), .B2(
        n9874), .ZN(n9321) );
  OAI21_X1 U10600 ( .B1(n9322), .B2(n9526), .A(n9321), .ZN(n9329) );
  AOI21_X1 U10601 ( .B1(n9324), .B2(n9323), .A(n9515), .ZN(n9327) );
  OAI22_X1 U10602 ( .A1(n9349), .A2(n9943), .B1(n9591), .B2(n9518), .ZN(n9325)
         );
  AOI21_X1 U10603 ( .B1(n9327), .B2(n9326), .A(n9325), .ZN(n9605) );
  NOR2_X1 U10604 ( .A1(n9605), .A2(n9877), .ZN(n9328) );
  AOI211_X1 U10605 ( .C1(n9528), .C2(n9602), .A(n9329), .B(n9328), .ZN(n9330)
         );
  OAI21_X1 U10606 ( .B1(n9606), .B2(n9513), .A(n9330), .ZN(P1_U3264) );
  OAI21_X1 U10607 ( .B1(n9332), .B2(n9336), .A(n9331), .ZN(n9334) );
  XOR2_X1 U10608 ( .A(n9336), .B(n9335), .Z(n9611) );
  NAND2_X1 U10609 ( .A1(n9611), .A2(n9582), .ZN(n9344) );
  AOI22_X1 U10610 ( .A1(n9877), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n9337), .B2(
        n9874), .ZN(n9338) );
  OAI21_X1 U10611 ( .B1(n9576), .B2(n9609), .A(n9338), .ZN(n9341) );
  OAI211_X1 U10612 ( .C1(n4945), .C2(n4324), .A(n9339), .B(n9569), .ZN(n9607)
         );
  NOR2_X1 U10613 ( .A1(n9607), .A2(n9580), .ZN(n9340) );
  AOI211_X1 U10614 ( .C1(n9578), .C2(n9342), .A(n9341), .B(n9340), .ZN(n9343)
         );
  OAI211_X1 U10615 ( .C1(n9877), .C2(n9608), .A(n9344), .B(n9343), .ZN(
        P1_U3265) );
  XNOR2_X1 U10616 ( .A(n9345), .B(n9346), .ZN(n9616) );
  INV_X1 U10617 ( .A(n9616), .ZN(n9358) );
  XNOR2_X1 U10618 ( .A(n9347), .B(n9346), .ZN(n9348) );
  OAI222_X1 U10619 ( .A1(n9943), .A2(n9350), .B1(n9518), .B2(n9349), .C1(n9348), .C2(n9515), .ZN(n9614) );
  AOI211_X1 U10620 ( .C1(n9352), .C2(n9351), .A(n9535), .B(n4324), .ZN(n9615)
         );
  NAND2_X1 U10621 ( .A1(n9615), .A2(n9528), .ZN(n9355) );
  AOI22_X1 U10622 ( .A1(n9877), .A2(P1_REG2_REG_25__SCAN_IN), .B1(n9874), .B2(
        n9353), .ZN(n9354) );
  OAI211_X1 U10623 ( .C1(n9714), .C2(n9526), .A(n9355), .B(n9354), .ZN(n9356)
         );
  AOI21_X1 U10624 ( .B1(n9614), .B2(n9541), .A(n9356), .ZN(n9357) );
  OAI21_X1 U10625 ( .B1(n9358), .B2(n9513), .A(n9357), .ZN(P1_U3266) );
  XNOR2_X1 U10626 ( .A(n9359), .B(n9362), .ZN(n9621) );
  INV_X1 U10627 ( .A(n9621), .ZN(n9375) );
  OAI21_X1 U10628 ( .B1(n9362), .B2(n9361), .A(n9360), .ZN(n9363) );
  NAND2_X1 U10629 ( .A1(n9363), .A2(n9563), .ZN(n9366) );
  AOI22_X1 U10630 ( .A1(n9393), .A2(n9914), .B1(n9562), .B2(n9364), .ZN(n9365)
         );
  NAND2_X1 U10631 ( .A1(n9366), .A2(n9365), .ZN(n9619) );
  INV_X1 U10632 ( .A(n9367), .ZN(n9385) );
  INV_X1 U10633 ( .A(n9351), .ZN(n9368) );
  AOI211_X1 U10634 ( .C1(n9369), .C2(n9385), .A(n9535), .B(n9368), .ZN(n9620)
         );
  NAND2_X1 U10635 ( .A1(n9620), .A2(n9528), .ZN(n9372) );
  AOI22_X1 U10636 ( .A1(n9877), .A2(P1_REG2_REG_24__SCAN_IN), .B1(n9370), .B2(
        n9874), .ZN(n9371) );
  OAI211_X1 U10637 ( .C1(n9718), .C2(n9526), .A(n9372), .B(n9371), .ZN(n9373)
         );
  AOI21_X1 U10638 ( .B1(n9541), .B2(n9619), .A(n9373), .ZN(n9374) );
  OAI21_X1 U10639 ( .B1(n9375), .B2(n9513), .A(n9374), .ZN(P1_U3267) );
  XOR2_X1 U10640 ( .A(n9376), .B(n9381), .Z(n9378) );
  AOI22_X1 U10641 ( .A1(n9378), .A2(n9563), .B1(n9562), .B2(n9377), .ZN(n9625)
         );
  NAND2_X1 U10642 ( .A1(n9380), .A2(n9379), .ZN(n9382) );
  XNOR2_X1 U10643 ( .A(n9382), .B(n9381), .ZN(n9628) );
  NAND2_X1 U10644 ( .A1(n9628), .A2(n9582), .ZN(n9390) );
  AOI22_X1 U10645 ( .A1(n9383), .A2(n9874), .B1(P1_REG2_REG_23__SCAN_IN), .B2(
        n9877), .ZN(n9384) );
  OAI21_X1 U10646 ( .B1(n9626), .B2(n9576), .A(n9384), .ZN(n9387) );
  OAI211_X1 U10647 ( .C1(n9722), .C2(n9401), .A(n9385), .B(n9569), .ZN(n9624)
         );
  NOR2_X1 U10648 ( .A1(n9624), .A2(n9580), .ZN(n9386) );
  AOI211_X1 U10649 ( .C1(n9578), .C2(n9388), .A(n9387), .B(n9386), .ZN(n9389)
         );
  OAI211_X1 U10650 ( .C1(n9877), .C2(n9625), .A(n9390), .B(n9389), .ZN(
        P1_U3268) );
  INV_X1 U10651 ( .A(n9396), .ZN(n9391) );
  XNOR2_X1 U10652 ( .A(n9392), .B(n9391), .ZN(n9395) );
  AND2_X1 U10653 ( .A1(n9393), .A2(n9562), .ZN(n9394) );
  AOI21_X1 U10654 ( .B1(n9395), .B2(n9563), .A(n9394), .ZN(n9632) );
  XNOR2_X1 U10655 ( .A(n9397), .B(n9396), .ZN(n9635) );
  NAND2_X1 U10656 ( .A1(n9635), .A2(n9582), .ZN(n9407) );
  AOI22_X1 U10657 ( .A1(n9398), .A2(n9874), .B1(P1_REG2_REG_22__SCAN_IN), .B2(
        n9877), .ZN(n9399) );
  OAI21_X1 U10658 ( .B1(n9633), .B2(n9576), .A(n9399), .ZN(n9404) );
  INV_X1 U10659 ( .A(n9405), .ZN(n9726) );
  INV_X1 U10660 ( .A(n9400), .ZN(n9415) );
  INV_X1 U10661 ( .A(n9401), .ZN(n9402) );
  OAI211_X1 U10662 ( .C1(n9726), .C2(n9415), .A(n9402), .B(n9569), .ZN(n9631)
         );
  NOR2_X1 U10663 ( .A1(n9631), .A2(n9580), .ZN(n9403) );
  AOI211_X1 U10664 ( .C1(n9578), .C2(n9405), .A(n9404), .B(n9403), .ZN(n9406)
         );
  OAI211_X1 U10665 ( .C1(n9877), .C2(n9632), .A(n9407), .B(n9406), .ZN(
        P1_U3269) );
  NAND2_X1 U10666 ( .A1(n9659), .A2(n9408), .ZN(n9411) );
  AND2_X1 U10667 ( .A1(n9411), .A2(n9409), .ZN(n9413) );
  NAND2_X1 U10668 ( .A1(n9411), .A2(n9410), .ZN(n9412) );
  OAI21_X1 U10669 ( .B1(n9413), .B2(n9419), .A(n9412), .ZN(n9644) );
  INV_X1 U10670 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n9414) );
  OAI22_X1 U10671 ( .A1(n9576), .A2(n9638), .B1(n9414), .B2(n9541), .ZN(n9425)
         );
  NAND2_X1 U10672 ( .A1(n9447), .A2(n9731), .ZN(n9441) );
  AOI211_X1 U10673 ( .C1(n9641), .C2(n9441), .A(n9535), .B(n9415), .ZN(n9639)
         );
  INV_X1 U10674 ( .A(n9416), .ZN(n9417) );
  AOI22_X1 U10675 ( .A1(n9639), .A2(n9418), .B1(n9874), .B2(n9417), .ZN(n9423)
         );
  XNOR2_X1 U10676 ( .A(n9420), .B(n9419), .ZN(n9422) );
  AOI22_X1 U10677 ( .A1(n9422), .A2(n9563), .B1(n9562), .B2(n9421), .ZN(n9642)
         );
  AOI21_X1 U10678 ( .B1(n9423), .B2(n9642), .A(n9877), .ZN(n9424) );
  AOI211_X1 U10679 ( .C1(n9578), .C2(n9641), .A(n9425), .B(n9424), .ZN(n9426)
         );
  OAI21_X1 U10680 ( .B1(n9513), .B2(n9644), .A(n9426), .ZN(P1_U3270) );
  NAND2_X1 U10681 ( .A1(n9659), .A2(n9427), .ZN(n9446) );
  NAND2_X1 U10682 ( .A1(n9446), .A2(n9428), .ZN(n9430) );
  NAND2_X1 U10683 ( .A1(n9430), .A2(n9429), .ZN(n9431) );
  XOR2_X1 U10684 ( .A(n9437), .B(n9431), .Z(n9647) );
  NAND2_X1 U10685 ( .A1(n9647), .A2(n9582), .ZN(n9445) );
  INV_X1 U10686 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n9433) );
  OAI22_X1 U10687 ( .A1(n9541), .A2(n9433), .B1(n9432), .B2(n9538), .ZN(n9434)
         );
  AOI21_X1 U10688 ( .B1(n9435), .B2(n9578), .A(n9434), .ZN(n9444) );
  NAND2_X1 U10689 ( .A1(n9452), .A2(n9436), .ZN(n9438) );
  XNOR2_X1 U10690 ( .A(n9438), .B(n9437), .ZN(n9439) );
  OAI222_X1 U10691 ( .A1(n9518), .A2(n9633), .B1(n9943), .B2(n9466), .C1(n9439), .C2(n9515), .ZN(n9645) );
  NAND2_X1 U10692 ( .A1(n9645), .A2(n9541), .ZN(n9443) );
  OR2_X1 U10693 ( .A1(n9447), .A2(n9731), .ZN(n9440) );
  NAND2_X1 U10694 ( .A1(n9646), .A2(n9528), .ZN(n9442) );
  NAND4_X1 U10695 ( .A1(n9445), .A2(n9444), .A3(n9443), .A4(n9442), .ZN(
        P1_U3271) );
  XNOR2_X1 U10696 ( .A(n9446), .B(n4541), .ZN(n9654) );
  INV_X1 U10697 ( .A(n9474), .ZN(n9448) );
  AOI211_X1 U10698 ( .C1(n9651), .C2(n9448), .A(n9535), .B(n9447), .ZN(n9650)
         );
  AOI22_X1 U10699 ( .A1(n9877), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9449), .B2(
        n9874), .ZN(n9450) );
  OAI21_X1 U10700 ( .B1(n9451), .B2(n9526), .A(n9450), .ZN(n9459) );
  OAI21_X1 U10701 ( .B1(n9454), .B2(n9453), .A(n9452), .ZN(n9457) );
  AOI222_X1 U10702 ( .A1(n9563), .A2(n9457), .B1(n9456), .B2(n9562), .C1(n9455), .C2(n9914), .ZN(n9653) );
  NOR2_X1 U10703 ( .A1(n9653), .A2(n9877), .ZN(n9458) );
  AOI211_X1 U10704 ( .C1(n9650), .C2(n9528), .A(n9459), .B(n9458), .ZN(n9460)
         );
  OAI21_X1 U10705 ( .B1(n9513), .B2(n9654), .A(n9460), .ZN(P1_U3272) );
  INV_X1 U10706 ( .A(n9461), .ZN(n9462) );
  AOI21_X1 U10707 ( .B1(n9464), .B2(n9463), .A(n9462), .ZN(n9465) );
  OAI222_X1 U10708 ( .A1(n9518), .A2(n9466), .B1(n9943), .B2(n9503), .C1(n9515), .C2(n9465), .ZN(n9655) );
  NAND2_X1 U10709 ( .A1(n9655), .A2(n9541), .ZN(n9478) );
  OAI22_X1 U10710 ( .A1(n9541), .A2(n9468), .B1(n9467), .B2(n9538), .ZN(n9469)
         );
  AOI21_X1 U10711 ( .B1(n9657), .B2(n9578), .A(n9469), .ZN(n9477) );
  NAND2_X1 U10712 ( .A1(n9471), .A2(n9470), .ZN(n9658) );
  NAND3_X1 U10713 ( .A1(n9659), .A2(n9658), .A3(n9582), .ZN(n9476) );
  NAND2_X1 U10714 ( .A1(n9487), .A2(n9657), .ZN(n9472) );
  NAND2_X1 U10715 ( .A1(n9472), .A2(n9569), .ZN(n9473) );
  NOR2_X1 U10716 ( .A1(n9474), .A2(n9473), .ZN(n9656) );
  NAND2_X1 U10717 ( .A1(n9656), .A2(n9528), .ZN(n9475) );
  NAND4_X1 U10718 ( .A1(n9478), .A2(n9477), .A3(n9476), .A4(n9475), .ZN(
        P1_U3273) );
  XNOR2_X1 U10719 ( .A(n9479), .B(n9482), .ZN(n9666) );
  NAND2_X1 U10720 ( .A1(n9480), .A2(n9481), .ZN(n9483) );
  XNOR2_X1 U10721 ( .A(n9483), .B(n9482), .ZN(n9484) );
  OAI222_X1 U10722 ( .A1(n9518), .A2(n9485), .B1(n9943), .B2(n9517), .C1(n9484), .C2(n9515), .ZN(n9662) );
  INV_X1 U10723 ( .A(n9487), .ZN(n9488) );
  AOI211_X1 U10724 ( .C1(n9664), .C2(n9486), .A(n9535), .B(n9488), .ZN(n9663)
         );
  NAND2_X1 U10725 ( .A1(n9663), .A2(n9528), .ZN(n9491) );
  AOI22_X1 U10726 ( .A1(n9877), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9489), .B2(
        n9874), .ZN(n9490) );
  OAI211_X1 U10727 ( .C1(n4949), .C2(n9526), .A(n9491), .B(n9490), .ZN(n9492)
         );
  AOI21_X1 U10728 ( .B1(n9541), .B2(n9662), .A(n9492), .ZN(n9493) );
  OAI21_X1 U10729 ( .B1(n9513), .B2(n9666), .A(n9493), .ZN(P1_U3274) );
  NAND2_X1 U10730 ( .A1(n9530), .A2(n9494), .ZN(n9496) );
  NAND2_X1 U10731 ( .A1(n9496), .A2(n9495), .ZN(n9498) );
  XNOR2_X1 U10732 ( .A(n9498), .B(n9497), .ZN(n9669) );
  INV_X1 U10733 ( .A(n9669), .ZN(n9512) );
  INV_X1 U10734 ( .A(n9480), .ZN(n9499) );
  AOI21_X1 U10735 ( .B1(n4338), .B2(n9500), .A(n9499), .ZN(n9501) );
  OAI222_X1 U10736 ( .A1(n9518), .A2(n9503), .B1(n9943), .B2(n9502), .C1(n9515), .C2(n9501), .ZN(n9667) );
  INV_X1 U10737 ( .A(n9521), .ZN(n9505) );
  INV_X1 U10738 ( .A(n9486), .ZN(n9504) );
  AOI211_X1 U10739 ( .C1(n9506), .C2(n9505), .A(n9535), .B(n9504), .ZN(n9668)
         );
  NAND2_X1 U10740 ( .A1(n9668), .A2(n9528), .ZN(n9509) );
  AOI22_X1 U10741 ( .A1(n9877), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n9507), .B2(
        n9874), .ZN(n9508) );
  OAI211_X1 U10742 ( .C1(n9737), .C2(n9526), .A(n9509), .B(n9508), .ZN(n9510)
         );
  AOI21_X1 U10743 ( .B1(n9667), .B2(n9541), .A(n9510), .ZN(n9511) );
  OAI21_X1 U10744 ( .B1(n9513), .B2(n9512), .A(n9511), .ZN(P1_U3275) );
  XNOR2_X1 U10745 ( .A(n9514), .B(n9529), .ZN(n9516) );
  OAI222_X1 U10746 ( .A1(n9943), .A2(n9519), .B1(n9518), .B2(n9517), .C1(n9516), .C2(n9515), .ZN(n9671) );
  INV_X1 U10747 ( .A(n9671), .ZN(n9533) );
  INV_X1 U10748 ( .A(n9520), .ZN(n9522) );
  AOI211_X1 U10749 ( .C1(n9523), .C2(n9522), .A(n9535), .B(n9521), .ZN(n9672)
         );
  AOI22_X1 U10750 ( .A1(n9877), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n9524), .B2(
        n9874), .ZN(n9525) );
  OAI21_X1 U10751 ( .B1(n9741), .B2(n9526), .A(n9525), .ZN(n9527) );
  AOI21_X1 U10752 ( .B1(n9672), .B2(n9528), .A(n9527), .ZN(n9532) );
  XNOR2_X1 U10753 ( .A(n9530), .B(n9529), .ZN(n9673) );
  NAND2_X1 U10754 ( .A1(n9673), .A2(n9582), .ZN(n9531) );
  OAI211_X1 U10755 ( .C1(n9533), .C2(n9877), .A(n9532), .B(n9531), .ZN(
        P1_U3276) );
  XNOR2_X1 U10756 ( .A(n9534), .B(n9552), .ZN(n9686) );
  AOI21_X1 U10757 ( .B1(n9570), .B2(n9681), .A(n9535), .ZN(n9536) );
  NAND2_X1 U10758 ( .A1(n9536), .A2(n4323), .ZN(n9682) );
  INV_X1 U10759 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n9540) );
  INV_X1 U10760 ( .A(n9537), .ZN(n9539) );
  OAI22_X1 U10761 ( .A1(n9541), .A2(n9540), .B1(n9539), .B2(n9538), .ZN(n9542)
         );
  AOI21_X1 U10762 ( .B1(n9544), .B2(n9543), .A(n9542), .ZN(n9546) );
  NAND2_X1 U10763 ( .A1(n9578), .A2(n9681), .ZN(n9545) );
  OAI211_X1 U10764 ( .C1(n9682), .C2(n9580), .A(n9546), .B(n9545), .ZN(n9556)
         );
  NAND2_X1 U10765 ( .A1(n9559), .A2(n9547), .ZN(n9549) );
  NAND2_X1 U10766 ( .A1(n9549), .A2(n9548), .ZN(n9551) );
  OAI21_X1 U10767 ( .B1(n9552), .B2(n9551), .A(n9550), .ZN(n9554) );
  AOI22_X1 U10768 ( .A1(n9554), .A2(n9563), .B1(n9562), .B2(n9553), .ZN(n9683)
         );
  NOR2_X1 U10769 ( .A1(n9683), .A2(n9877), .ZN(n9555) );
  AOI211_X1 U10770 ( .C1(n9686), .C2(n9582), .A(n9556), .B(n9555), .ZN(n9557)
         );
  INV_X1 U10771 ( .A(n9557), .ZN(P1_U3278) );
  NAND2_X1 U10772 ( .A1(n9559), .A2(n9558), .ZN(n9560) );
  XOR2_X1 U10773 ( .A(n9568), .B(n9560), .Z(n9564) );
  AOI22_X1 U10774 ( .A1(n9564), .A2(n9563), .B1(n9562), .B2(n9561), .ZN(n9694)
         );
  INV_X1 U10775 ( .A(n9565), .ZN(n9566) );
  AOI21_X1 U10776 ( .B1(n9568), .B2(n9567), .A(n9566), .ZN(n9688) );
  OAI211_X1 U10777 ( .C1(n9572), .C2(n9571), .A(n9570), .B(n9569), .ZN(n9691)
         );
  AOI22_X1 U10778 ( .A1(n9877), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n9573), .B2(
        n9874), .ZN(n9574) );
  OAI21_X1 U10779 ( .B1(n9576), .B2(n9575), .A(n9574), .ZN(n9577) );
  AOI21_X1 U10780 ( .B1(n9578), .B2(n9690), .A(n9577), .ZN(n9579) );
  OAI21_X1 U10781 ( .B1(n9691), .B2(n9580), .A(n9579), .ZN(n9581) );
  AOI21_X1 U10782 ( .B1(n9688), .B2(n9582), .A(n9581), .ZN(n9583) );
  OAI21_X1 U10783 ( .B1(n9694), .B2(n9877), .A(n9583), .ZN(P1_U3279) );
  INV_X1 U10784 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n9586) );
  NOR2_X1 U10785 ( .A1(n9585), .A2(n9584), .ZN(n9702) );
  OAI21_X1 U10786 ( .B1(n9705), .B2(n9701), .A(n9587), .ZN(P1_U3553) );
  NOR4_X1 U10787 ( .A1(n9598), .A2(n9590), .A3(n9591), .A4(n9950), .ZN(n9593)
         );
  OAI22_X1 U10788 ( .A1(n4943), .A2(n9961), .B1(n9591), .B2(n9943), .ZN(n9592)
         );
  NAND2_X1 U10789 ( .A1(n9299), .A2(n4985), .ZN(n9600) );
  MUX2_X1 U10790 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n9706), .S(n9986), .Z(
        P1_U3552) );
  AOI21_X1 U10791 ( .B1(n9913), .B2(n9603), .A(n9602), .ZN(n9604) );
  OAI211_X1 U10792 ( .C1(n9606), .C2(n9950), .A(n9605), .B(n9604), .ZN(n9707)
         );
  MUX2_X1 U10793 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9707), .S(n9986), .Z(
        P1_U3550) );
  INV_X1 U10794 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n9612) );
  OAI211_X1 U10795 ( .C1(n9609), .C2(n9943), .A(n9608), .B(n9607), .ZN(n9610)
         );
  AOI21_X1 U10796 ( .B1(n9611), .B2(n9966), .A(n9610), .ZN(n9708) );
  MUX2_X1 U10797 ( .A(n9612), .B(n9708), .S(n9986), .Z(n9613) );
  OAI21_X1 U10798 ( .B1(n4945), .B2(n9701), .A(n9613), .ZN(P1_U3549) );
  INV_X1 U10799 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n9617) );
  AOI211_X1 U10800 ( .C1(n9966), .C2(n9616), .A(n9615), .B(n9614), .ZN(n9711)
         );
  MUX2_X1 U10801 ( .A(n9617), .B(n9711), .S(n9986), .Z(n9618) );
  OAI21_X1 U10802 ( .B1(n9714), .B2(n9701), .A(n9618), .ZN(P1_U3548) );
  INV_X1 U10803 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n9622) );
  AOI211_X1 U10804 ( .C1(n9621), .C2(n9966), .A(n9620), .B(n9619), .ZN(n9715)
         );
  MUX2_X1 U10805 ( .A(n9622), .B(n9715), .S(n9986), .Z(n9623) );
  OAI21_X1 U10806 ( .B1(n9718), .B2(n9701), .A(n9623), .ZN(P1_U3547) );
  INV_X1 U10807 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n9629) );
  OAI211_X1 U10808 ( .C1(n9626), .C2(n9943), .A(n9625), .B(n9624), .ZN(n9627)
         );
  AOI21_X1 U10809 ( .B1(n9628), .B2(n9966), .A(n9627), .ZN(n9719) );
  MUX2_X1 U10810 ( .A(n9629), .B(n9719), .S(n9986), .Z(n9630) );
  OAI21_X1 U10811 ( .B1(n9722), .B2(n9701), .A(n9630), .ZN(P1_U3546) );
  OAI211_X1 U10812 ( .C1(n9633), .C2(n9943), .A(n9632), .B(n9631), .ZN(n9634)
         );
  AOI21_X1 U10813 ( .B1(n9635), .B2(n9966), .A(n9634), .ZN(n9724) );
  INV_X1 U10814 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n9636) );
  MUX2_X1 U10815 ( .A(n9724), .B(n9636), .S(n5699), .Z(n9637) );
  OAI21_X1 U10816 ( .B1(n9726), .B2(n9701), .A(n9637), .ZN(P1_U3545) );
  NOR2_X1 U10817 ( .A1(n9638), .A2(n9943), .ZN(n9640) );
  AOI211_X1 U10818 ( .C1(n9913), .C2(n9641), .A(n9640), .B(n9639), .ZN(n9643)
         );
  OAI211_X1 U10819 ( .C1(n9950), .C2(n9644), .A(n9643), .B(n9642), .ZN(n9727)
         );
  MUX2_X1 U10820 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9727), .S(n9986), .Z(
        P1_U3544) );
  INV_X1 U10821 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n9648) );
  AOI211_X1 U10822 ( .C1(n9647), .C2(n9966), .A(n9646), .B(n9645), .ZN(n9728)
         );
  MUX2_X1 U10823 ( .A(n9648), .B(n9728), .S(n9986), .Z(n9649) );
  OAI21_X1 U10824 ( .B1(n9731), .B2(n9701), .A(n9649), .ZN(P1_U3543) );
  AOI21_X1 U10825 ( .B1(n9913), .B2(n9651), .A(n9650), .ZN(n9652) );
  OAI211_X1 U10826 ( .C1(n9950), .C2(n9654), .A(n9653), .B(n9652), .ZN(n9732)
         );
  MUX2_X1 U10827 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9732), .S(n9986), .Z(
        P1_U3542) );
  AOI211_X1 U10828 ( .C1(n9913), .C2(n9657), .A(n9656), .B(n9655), .ZN(n9661)
         );
  NAND3_X1 U10829 ( .A1(n9659), .A2(n9966), .A3(n9658), .ZN(n9660) );
  NAND2_X1 U10830 ( .A1(n9661), .A2(n9660), .ZN(n9733) );
  MUX2_X1 U10831 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9733), .S(n9986), .Z(
        P1_U3541) );
  AOI211_X1 U10832 ( .C1(n9913), .C2(n9664), .A(n9663), .B(n9662), .ZN(n9665)
         );
  OAI21_X1 U10833 ( .B1(n9950), .B2(n9666), .A(n9665), .ZN(n9734) );
  MUX2_X1 U10834 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9734), .S(n9986), .Z(
        P1_U3540) );
  AOI211_X1 U10835 ( .C1(n9669), .C2(n9966), .A(n9668), .B(n9667), .ZN(n9735)
         );
  MUX2_X1 U10836 ( .A(n10240), .B(n9735), .S(n9986), .Z(n9670) );
  OAI21_X1 U10837 ( .B1(n9737), .B2(n9701), .A(n9670), .ZN(P1_U3539) );
  INV_X1 U10838 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n9674) );
  AOI211_X1 U10839 ( .C1(n9673), .C2(n9966), .A(n9672), .B(n9671), .ZN(n9738)
         );
  MUX2_X1 U10840 ( .A(n9674), .B(n9738), .S(n9986), .Z(n9675) );
  OAI21_X1 U10841 ( .B1(n9741), .B2(n9701), .A(n9675), .ZN(P1_U3538) );
  AOI211_X1 U10842 ( .C1(n9913), .C2(n9678), .A(n9677), .B(n9676), .ZN(n9679)
         );
  OAI21_X1 U10843 ( .B1(n9950), .B2(n9680), .A(n9679), .ZN(n9742) );
  MUX2_X1 U10844 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n9742), .S(n9986), .Z(
        P1_U3537) );
  INV_X1 U10845 ( .A(n9681), .ZN(n9746) );
  OAI211_X1 U10846 ( .C1(n9684), .C2(n9943), .A(n9683), .B(n9682), .ZN(n9685)
         );
  AOI21_X1 U10847 ( .B1(n9686), .B2(n9966), .A(n9685), .ZN(n9743) );
  MUX2_X1 U10848 ( .A(n10253), .B(n9743), .S(n9986), .Z(n9687) );
  OAI21_X1 U10849 ( .B1(n9746), .B2(n9701), .A(n9687), .ZN(P1_U3536) );
  NAND2_X1 U10850 ( .A1(n9688), .A2(n9966), .ZN(n9693) );
  AOI22_X1 U10851 ( .A1(n9690), .A2(n9913), .B1(n9689), .B2(n9914), .ZN(n9692)
         );
  NAND4_X1 U10852 ( .A1(n9694), .A2(n9693), .A3(n9692), .A4(n9691), .ZN(n9747)
         );
  MUX2_X1 U10853 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n9747), .S(n9986), .Z(
        P1_U3535) );
  NAND2_X1 U10854 ( .A1(n9695), .A2(n9966), .ZN(n9697) );
  AND3_X1 U10855 ( .A1(n9698), .A2(n9697), .A3(n9696), .ZN(n9748) );
  MUX2_X1 U10856 ( .A(n9699), .B(n9748), .S(n9986), .Z(n9700) );
  OAI21_X1 U10857 ( .B1(n4951), .B2(n9701), .A(n9700), .ZN(P1_U3534) );
  INV_X1 U10858 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n9703) );
  OAI21_X1 U10859 ( .B1(n9705), .B2(n9751), .A(n9704), .ZN(P1_U3521) );
  MUX2_X1 U10860 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9707), .S(n9970), .Z(
        P1_U3518) );
  INV_X1 U10861 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n9709) );
  MUX2_X1 U10862 ( .A(n9709), .B(n9708), .S(n9970), .Z(n9710) );
  OAI21_X1 U10863 ( .B1(n4945), .B2(n9751), .A(n9710), .ZN(P1_U3517) );
  INV_X1 U10864 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n9712) );
  MUX2_X1 U10865 ( .A(n9712), .B(n9711), .S(n9970), .Z(n9713) );
  OAI21_X1 U10866 ( .B1(n9714), .B2(n9751), .A(n9713), .ZN(P1_U3516) );
  INV_X1 U10867 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n9716) );
  MUX2_X1 U10868 ( .A(n9716), .B(n9715), .S(n9970), .Z(n9717) );
  OAI21_X1 U10869 ( .B1(n9718), .B2(n9751), .A(n9717), .ZN(P1_U3515) );
  MUX2_X1 U10870 ( .A(n9720), .B(n9719), .S(n9970), .Z(n9721) );
  OAI21_X1 U10871 ( .B1(n9722), .B2(n9751), .A(n9721), .ZN(P1_U3514) );
  MUX2_X1 U10872 ( .A(n9724), .B(n9723), .S(n9968), .Z(n9725) );
  OAI21_X1 U10873 ( .B1(n9726), .B2(n9751), .A(n9725), .ZN(P1_U3513) );
  MUX2_X1 U10874 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9727), .S(n9970), .Z(
        P1_U3512) );
  INV_X1 U10875 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n9729) );
  MUX2_X1 U10876 ( .A(n9729), .B(n9728), .S(n9970), .Z(n9730) );
  OAI21_X1 U10877 ( .B1(n9731), .B2(n9751), .A(n9730), .ZN(P1_U3511) );
  MUX2_X1 U10878 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9732), .S(n9970), .Z(
        P1_U3510) );
  MUX2_X1 U10879 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9733), .S(n9970), .Z(
        P1_U3508) );
  MUX2_X1 U10880 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9734), .S(n9970), .Z(
        P1_U3505) );
  MUX2_X1 U10881 ( .A(n10257), .B(n9735), .S(n9970), .Z(n9736) );
  OAI21_X1 U10882 ( .B1(n9737), .B2(n9751), .A(n9736), .ZN(P1_U3502) );
  INV_X1 U10883 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n9739) );
  MUX2_X1 U10884 ( .A(n9739), .B(n9738), .S(n9970), .Z(n9740) );
  OAI21_X1 U10885 ( .B1(n9741), .B2(n9751), .A(n9740), .ZN(P1_U3499) );
  MUX2_X1 U10886 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n9742), .S(n9970), .Z(
        P1_U3496) );
  INV_X1 U10887 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n9744) );
  MUX2_X1 U10888 ( .A(n9744), .B(n9743), .S(n9970), .Z(n9745) );
  OAI21_X1 U10889 ( .B1(n9746), .B2(n9751), .A(n9745), .ZN(P1_U3493) );
  MUX2_X1 U10890 ( .A(P1_REG0_REG_12__SCAN_IN), .B(n9747), .S(n9970), .Z(
        P1_U3490) );
  INV_X1 U10891 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n9749) );
  MUX2_X1 U10892 ( .A(n9749), .B(n9748), .S(n9970), .Z(n9750) );
  OAI21_X1 U10893 ( .B1(n4951), .B2(n9751), .A(n9750), .ZN(P1_U3487) );
  NOR4_X1 U10894 ( .A1(n9753), .A2(P1_IR_REG_30__SCAN_IN), .A3(P1_U3084), .A4(
        n9752), .ZN(n9754) );
  AOI21_X1 U10895 ( .B1(n9755), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9754), .ZN(
        n9756) );
  OAI21_X1 U10896 ( .B1(n9757), .B2(n9763), .A(n9756), .ZN(P1_U3322) );
  INV_X1 U10897 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n9760) );
  OAI222_X1 U10898 ( .A1(n9765), .A2(n9760), .B1(n9763), .B2(n9759), .C1(
        P1_U3084), .C2(n9758), .ZN(P1_U3323) );
  INV_X1 U10899 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n9764) );
  OAI222_X1 U10900 ( .A1(n9765), .A2(n9764), .B1(n9763), .B2(n9762), .C1(
        P1_U3084), .C2(n9761), .ZN(P1_U3324) );
  MUX2_X1 U10901 ( .A(n9766), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3353) );
  INV_X1 U10902 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n10293) );
  NOR2_X1 U10903 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n9767) );
  AOI21_X1 U10904 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n9767), .ZN(n10108) );
  NOR2_X1 U10905 ( .A1(P1_ADDR_REG_16__SCAN_IN), .A2(P2_ADDR_REG_16__SCAN_IN), 
        .ZN(n9768) );
  AOI21_X1 U10906 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n9768), .ZN(n10111) );
  NOR2_X1 U10907 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n9769) );
  AOI21_X1 U10908 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n9769), .ZN(n10114) );
  NOR2_X1 U10909 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n9770) );
  AOI21_X1 U10910 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n9770), .ZN(n10117) );
  NOR2_X1 U10911 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n9771) );
  AOI21_X1 U10912 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n9771), .ZN(n10120) );
  NOR2_X1 U10913 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n9780) );
  XOR2_X1 U10914 ( .A(n9772), .B(P2_ADDR_REG_4__SCAN_IN), .Z(n10304) );
  NAND2_X1 U10915 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n9778) );
  XNOR2_X1 U10916 ( .A(n9773), .B(P2_ADDR_REG_3__SCAN_IN), .ZN(n10302) );
  NAND2_X1 U10917 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n9776) );
  XNOR2_X1 U10918 ( .A(P2_ADDR_REG_2__SCAN_IN), .B(n9774), .ZN(n10300) );
  AOI21_X1 U10919 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10101) );
  NAND3_X1 U10920 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_1__SCAN_IN), .ZN(n10103) );
  NAND2_X1 U10921 ( .A1(n10300), .A2(n10299), .ZN(n9775) );
  NAND2_X1 U10922 ( .A1(n9776), .A2(n9775), .ZN(n10301) );
  NAND2_X1 U10923 ( .A1(n10302), .A2(n10301), .ZN(n9777) );
  NAND2_X1 U10924 ( .A1(n9778), .A2(n9777), .ZN(n10303) );
  NOR2_X1 U10925 ( .A1(n10304), .A2(n10303), .ZN(n9779) );
  NOR2_X1 U10926 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n9781), .ZN(n10287) );
  NAND2_X1 U10927 ( .A1(n9783), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n9785) );
  NAND2_X1 U10928 ( .A1(n10286), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n9784) );
  NAND2_X1 U10929 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n9786), .ZN(n9788) );
  NAND2_X1 U10930 ( .A1(n10290), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n9787) );
  NAND2_X1 U10931 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n9789), .ZN(n9791) );
  NAND2_X1 U10932 ( .A1(n10295), .A2(P2_ADDR_REG_8__SCAN_IN), .ZN(n9790) );
  NAND2_X1 U10933 ( .A1(n9791), .A2(n9790), .ZN(n9792) );
  INV_X1 U10934 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n10298) );
  XNOR2_X1 U10935 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n9792), .ZN(n10297) );
  NAND2_X1 U10936 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n9794) );
  OAI21_X1 U10937 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n9794), .ZN(n10128) );
  NAND2_X1 U10938 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n9795) );
  OAI21_X1 U10939 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n9795), .ZN(n10125) );
  NOR2_X1 U10940 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n9796) );
  AOI21_X1 U10941 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n9796), .ZN(n10122) );
  NAND2_X1 U10942 ( .A1(n10117), .A2(n10116), .ZN(n10115) );
  NAND2_X1 U10943 ( .A1(n10114), .A2(n10113), .ZN(n10112) );
  NAND2_X1 U10944 ( .A1(n10108), .A2(n10107), .ZN(n10106) );
  NOR2_X1 U10945 ( .A1(n10293), .A2(n10292), .ZN(n9797) );
  NAND2_X1 U10946 ( .A1(n10293), .A2(n10292), .ZN(n10291) );
  XNOR2_X1 U10947 ( .A(n4545), .B(P1_ADDR_REG_19__SCAN_IN), .ZN(n9798) );
  XNOR2_X1 U10948 ( .A(n9799), .B(n9798), .ZN(ADD_1071_U4) );
  XNOR2_X1 U10949 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U10950 ( .A(P2_RD_REG_SCAN_IN), .B(P1_RD_REG_SCAN_IN), .ZN(U126) );
  INV_X1 U10951 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n9814) );
  INV_X1 U10952 ( .A(n9800), .ZN(n9804) );
  INV_X1 U10953 ( .A(n9801), .ZN(n9803) );
  AOI211_X1 U10954 ( .C1(P1_IR_REG_0__SCAN_IN), .C2(n9804), .A(n9803), .B(
        n9802), .ZN(n9809) );
  INV_X1 U10955 ( .A(n9805), .ZN(n9807) );
  OAI21_X1 U10956 ( .B1(n9807), .B2(n9811), .A(n9806), .ZN(n9808) );
  AOI22_X1 U10957 ( .A1(n9810), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(n9809), .B2(
        n9808), .ZN(n9813) );
  NAND3_X1 U10958 ( .A1(n9862), .A2(P1_IR_REG_0__SCAN_IN), .A3(n9811), .ZN(
        n9812) );
  OAI211_X1 U10959 ( .C1(P1_STATE_REG_SCAN_IN), .C2(n9814), .A(n9813), .B(
        n9812), .ZN(P1_U3241) );
  AOI211_X1 U10960 ( .C1(n9817), .C2(n9816), .A(n9815), .B(n9839), .ZN(n9818)
         );
  AOI211_X1 U10961 ( .C1(n4479), .C2(n9820), .A(n9819), .B(n9818), .ZN(n9825)
         );
  XNOR2_X1 U10962 ( .A(n9822), .B(n9821), .ZN(n9823) );
  NAND2_X1 U10963 ( .A1(n9823), .A2(n9862), .ZN(n9824) );
  OAI211_X1 U10964 ( .C1(n4437), .C2(n9867), .A(n9825), .B(n9824), .ZN(
        P1_U3254) );
  INV_X1 U10965 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n9837) );
  INV_X1 U10966 ( .A(n9826), .ZN(n9831) );
  AOI211_X1 U10967 ( .C1(n9829), .C2(n9828), .A(n9827), .B(n9839), .ZN(n9830)
         );
  AOI211_X1 U10968 ( .C1(n4479), .C2(n9832), .A(n9831), .B(n9830), .ZN(n9836)
         );
  OAI211_X1 U10969 ( .C1(n9834), .C2(P1_REG1_REG_15__SCAN_IN), .A(n9862), .B(
        n9833), .ZN(n9835) );
  OAI211_X1 U10970 ( .C1(n9837), .C2(n9867), .A(n9836), .B(n9835), .ZN(
        P1_U3256) );
  INV_X1 U10971 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n9850) );
  INV_X1 U10972 ( .A(n9838), .ZN(n9843) );
  AOI211_X1 U10973 ( .C1(n4391), .C2(n9841), .A(n9840), .B(n9839), .ZN(n9842)
         );
  AOI211_X1 U10974 ( .C1(n4479), .C2(n9844), .A(n9843), .B(n9842), .ZN(n9849)
         );
  OAI211_X1 U10975 ( .C1(n9847), .C2(n9846), .A(n9862), .B(n9845), .ZN(n9848)
         );
  OAI211_X1 U10976 ( .C1(n9850), .C2(n9867), .A(n9849), .B(n9848), .ZN(
        P1_U3257) );
  INV_X1 U10977 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n9868) );
  AOI21_X1 U10978 ( .B1(n9853), .B2(n9852), .A(n9851), .ZN(n9854) );
  NAND2_X1 U10979 ( .A1(n9855), .A2(n9854), .ZN(n9857) );
  OAI211_X1 U10980 ( .C1(n9859), .C2(n9858), .A(n9857), .B(n9856), .ZN(n9860)
         );
  INV_X1 U10981 ( .A(n9860), .ZN(n9866) );
  OAI211_X1 U10982 ( .C1(n9864), .C2(n9863), .A(n9862), .B(n9861), .ZN(n9865)
         );
  OAI211_X1 U10983 ( .C1(n9868), .C2(n9867), .A(n9866), .B(n9865), .ZN(
        P1_U3258) );
  INV_X1 U10984 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n9876) );
  NOR2_X1 U10985 ( .A1(n9870), .A2(n9869), .ZN(n9873) );
  INV_X1 U10986 ( .A(n9871), .ZN(n9872) );
  AOI211_X1 U10987 ( .C1(n9874), .C2(P1_REG3_REG_0__SCAN_IN), .A(n9873), .B(
        n9872), .ZN(n9875) );
  AOI22_X1 U10988 ( .A1(n9877), .A2(n9876), .B1(n9875), .B2(n9541), .ZN(
        P1_U3291) );
  INV_X1 U10989 ( .A(n9878), .ZN(n9879) );
  AND2_X1 U10990 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n9881), .ZN(P1_U3292) );
  AND2_X1 U10991 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n9881), .ZN(P1_U3293) );
  AND2_X1 U10992 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n9881), .ZN(P1_U3294) );
  AND2_X1 U10993 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n9881), .ZN(P1_U3295) );
  AND2_X1 U10994 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n9881), .ZN(P1_U3296) );
  AND2_X1 U10995 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n9881), .ZN(P1_U3297) );
  AND2_X1 U10996 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n9881), .ZN(P1_U3298) );
  AND2_X1 U10997 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n9881), .ZN(P1_U3299) );
  AND2_X1 U10998 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n9881), .ZN(P1_U3300) );
  AND2_X1 U10999 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n9881), .ZN(P1_U3301) );
  NOR2_X1 U11000 ( .A1(n9880), .A2(n10199), .ZN(P1_U3302) );
  AND2_X1 U11001 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n9881), .ZN(P1_U3303) );
  AND2_X1 U11002 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n9881), .ZN(P1_U3304) );
  AND2_X1 U11003 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n9881), .ZN(P1_U3305) );
  AND2_X1 U11004 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n9881), .ZN(P1_U3306) );
  AND2_X1 U11005 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n9881), .ZN(P1_U3307) );
  NOR2_X1 U11006 ( .A1(n9880), .A2(n10247), .ZN(P1_U3308) );
  AND2_X1 U11007 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n9881), .ZN(P1_U3309) );
  AND2_X1 U11008 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n9881), .ZN(P1_U3310) );
  AND2_X1 U11009 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n9881), .ZN(P1_U3311) );
  AND2_X1 U11010 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n9881), .ZN(P1_U3312) );
  AND2_X1 U11011 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n9881), .ZN(P1_U3313) );
  AND2_X1 U11012 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n9881), .ZN(P1_U3314) );
  AND2_X1 U11013 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n9881), .ZN(P1_U3315) );
  AND2_X1 U11014 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n9881), .ZN(P1_U3316) );
  AND2_X1 U11015 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n9881), .ZN(P1_U3317) );
  NOR2_X1 U11016 ( .A1(n9880), .A2(n10227), .ZN(P1_U3318) );
  NOR2_X1 U11017 ( .A1(n9880), .A2(n10173), .ZN(P1_U3319) );
  AND2_X1 U11018 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n9881), .ZN(P1_U3320) );
  AND2_X1 U11019 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n9881), .ZN(P1_U3321) );
  OAI21_X1 U11020 ( .B1(n9884), .B2(n9883), .A(n9882), .ZN(P1_U3440) );
  INV_X1 U11021 ( .A(n9885), .ZN(n9886) );
  AOI21_X1 U11022 ( .B1(n9887), .B2(n9894), .A(n9886), .ZN(n9892) );
  OAI21_X1 U11023 ( .B1(n9889), .B2(n9961), .A(n9888), .ZN(n9890) );
  NOR3_X1 U11024 ( .A1(n9892), .A2(n9891), .A3(n9890), .ZN(n9972) );
  INV_X1 U11025 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n9893) );
  AOI22_X1 U11026 ( .A1(n9970), .A2(n9972), .B1(n9893), .B2(n9968), .ZN(
        P1_U3457) );
  INV_X1 U11027 ( .A(n9894), .ZN(n9911) );
  OAI21_X1 U11028 ( .B1(n9896), .B2(n9961), .A(n9895), .ZN(n9899) );
  INV_X1 U11029 ( .A(n9897), .ZN(n9898) );
  AOI211_X1 U11030 ( .C1(n9911), .C2(n9900), .A(n9899), .B(n9898), .ZN(n9974)
         );
  INV_X1 U11031 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n9901) );
  AOI22_X1 U11032 ( .A1(n9970), .A2(n9974), .B1(n9901), .B2(n9968), .ZN(
        P1_U3460) );
  OAI22_X1 U11033 ( .A1(n5105), .A2(n9943), .B1(n9902), .B2(n9961), .ZN(n9903)
         );
  NOR2_X1 U11034 ( .A1(n9904), .A2(n9903), .ZN(n9908) );
  NAND2_X1 U11035 ( .A1(n9905), .A2(n9911), .ZN(n9907) );
  NAND2_X1 U11036 ( .A1(n9905), .A2(n9923), .ZN(n9906) );
  INV_X1 U11037 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n9910) );
  AOI22_X1 U11038 ( .A1(n9970), .A2(n9975), .B1(n9910), .B2(n9968), .ZN(
        P1_U3463) );
  NAND2_X1 U11039 ( .A1(n9922), .A2(n9911), .ZN(n9918) );
  AOI22_X1 U11040 ( .A1(n9915), .A2(n9914), .B1(n9913), .B2(n9912), .ZN(n9917)
         );
  NAND3_X1 U11041 ( .A1(n9918), .A2(n9917), .A3(n9916), .ZN(n9921) );
  INV_X1 U11042 ( .A(n9919), .ZN(n9920) );
  AOI211_X1 U11043 ( .C1(n9923), .C2(n9922), .A(n9921), .B(n9920), .ZN(n9976)
         );
  INV_X1 U11044 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n9924) );
  AOI22_X1 U11045 ( .A1(n9970), .A2(n9976), .B1(n9924), .B2(n9968), .ZN(
        P1_U3466) );
  NOR3_X1 U11046 ( .A1(n9926), .A2(n9925), .A3(n9950), .ZN(n9931) );
  OAI22_X1 U11047 ( .A1(n9928), .A2(n9943), .B1(n9927), .B2(n9961), .ZN(n9929)
         );
  NOR4_X1 U11048 ( .A1(n9932), .A2(n9931), .A3(n9930), .A4(n9929), .ZN(n9978)
         );
  INV_X1 U11049 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n9933) );
  AOI22_X1 U11050 ( .A1(n9970), .A2(n9978), .B1(n9933), .B2(n9968), .ZN(
        P1_U3469) );
  INV_X1 U11051 ( .A(n9934), .ZN(n9936) );
  AOI211_X1 U11052 ( .C1(n9937), .C2(n9966), .A(n9936), .B(n9935), .ZN(n9938)
         );
  AND2_X1 U11053 ( .A1(n9939), .A2(n9938), .ZN(n9980) );
  INV_X1 U11054 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n9940) );
  AOI22_X1 U11055 ( .A1(n9970), .A2(n9980), .B1(n9940), .B2(n9968), .ZN(
        P1_U3472) );
  NOR2_X1 U11056 ( .A1(n9941), .A2(n9950), .ZN(n9947) );
  OAI22_X1 U11057 ( .A1(n9944), .A2(n9943), .B1(n9942), .B2(n9961), .ZN(n9945)
         );
  NOR4_X1 U11058 ( .A1(n9948), .A2(n9947), .A3(n9946), .A4(n9945), .ZN(n9982)
         );
  INV_X1 U11059 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n9949) );
  AOI22_X1 U11060 ( .A1(n9970), .A2(n9982), .B1(n9949), .B2(n9968), .ZN(
        P1_U3475) );
  NOR2_X1 U11061 ( .A1(n9951), .A2(n9950), .ZN(n9957) );
  OAI21_X1 U11062 ( .B1(n9953), .B2(n9961), .A(n9952), .ZN(n9955) );
  AOI211_X1 U11063 ( .C1(n9957), .C2(n9956), .A(n9955), .B(n9954), .ZN(n9983)
         );
  INV_X1 U11064 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n9958) );
  AOI22_X1 U11065 ( .A1(n9970), .A2(n9983), .B1(n9958), .B2(n9968), .ZN(
        P1_U3478) );
  INV_X1 U11066 ( .A(n9959), .ZN(n9960) );
  OAI21_X1 U11067 ( .B1(n9962), .B2(n9961), .A(n9960), .ZN(n9965) );
  INV_X1 U11068 ( .A(n9963), .ZN(n9964) );
  AOI211_X1 U11069 ( .C1(n9967), .C2(n9966), .A(n9965), .B(n9964), .ZN(n9985)
         );
  INV_X1 U11070 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n9969) );
  AOI22_X1 U11071 ( .A1(n9970), .A2(n9985), .B1(n9969), .B2(n9968), .ZN(
        P1_U3481) );
  AOI22_X1 U11072 ( .A1(n9986), .A2(n9972), .B1(n9971), .B2(n5699), .ZN(
        P1_U3524) );
  AOI22_X1 U11073 ( .A1(n9986), .A2(n9974), .B1(n9973), .B2(n5699), .ZN(
        P1_U3525) );
  AOI22_X1 U11074 ( .A1(n9986), .A2(n9975), .B1(n6606), .B2(n5699), .ZN(
        P1_U3526) );
  AOI22_X1 U11075 ( .A1(n9986), .A2(n9976), .B1(n6629), .B2(n5699), .ZN(
        P1_U3527) );
  INV_X1 U11076 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n9977) );
  AOI22_X1 U11077 ( .A1(n9986), .A2(n9978), .B1(n9977), .B2(n5699), .ZN(
        P1_U3528) );
  INV_X1 U11078 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n9979) );
  AOI22_X1 U11079 ( .A1(n9986), .A2(n9980), .B1(n9979), .B2(n5699), .ZN(
        P1_U3529) );
  INV_X1 U11080 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n9981) );
  AOI22_X1 U11081 ( .A1(n9986), .A2(n9982), .B1(n9981), .B2(n5699), .ZN(
        P1_U3530) );
  AOI22_X1 U11082 ( .A1(n9986), .A2(n9983), .B1(n6865), .B2(n5699), .ZN(
        P1_U3531) );
  INV_X1 U11083 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n9984) );
  AOI22_X1 U11084 ( .A1(n9986), .A2(n9985), .B1(n9984), .B2(n5699), .ZN(
        P1_U3532) );
  AOI22_X1 U11085 ( .A1(n9999), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n10005), .ZN(n9994) );
  AOI22_X1 U11086 ( .A1(n9997), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3152), .ZN(n9993) );
  NOR2_X1 U11087 ( .A1(n9987), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n9991) );
  OAI21_X1 U11088 ( .B1(n9989), .B2(P2_REG1_REG_0__SCAN_IN), .A(n9988), .ZN(
        n9990) );
  OAI21_X1 U11089 ( .B1(n9991), .B2(n9990), .A(P2_IR_REG_0__SCAN_IN), .ZN(
        n9992) );
  OAI211_X1 U11090 ( .C1(P2_IR_REG_0__SCAN_IN), .C2(n9994), .A(n9993), .B(
        n9992), .ZN(P2_U3245) );
  INV_X1 U11091 ( .A(n9995), .ZN(n9996) );
  AOI21_X1 U11092 ( .B1(n9997), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n9996), .ZN(
        n10011) );
  OAI211_X1 U11093 ( .C1(n10001), .C2(n10000), .A(n9999), .B(n9998), .ZN(
        n10010) );
  NAND2_X1 U11094 ( .A1(n10003), .A2(n10002), .ZN(n10009) );
  OAI211_X1 U11095 ( .C1(n10007), .C2(n10006), .A(n10005), .B(n10004), .ZN(
        n10008) );
  NAND4_X1 U11096 ( .A1(n10011), .A2(n10010), .A3(n10009), .A4(n10008), .ZN(
        P2_U3262) );
  XNOR2_X1 U11097 ( .A(n6251), .B(n10013), .ZN(n10018) );
  XNOR2_X1 U11098 ( .A(n10012), .B(n10013), .ZN(n10054) );
  NOR2_X1 U11099 ( .A1(n10054), .A2(n10014), .ZN(n10015) );
  AOI211_X1 U11100 ( .C1(n10018), .C2(n10017), .A(n10016), .B(n10015), .ZN(
        n10057) );
  OAI211_X1 U11101 ( .C1(n10021), .C2(n10056), .A(n10020), .B(n10019), .ZN(
        n10055) );
  OAI22_X1 U11102 ( .A1(n10023), .A2(n10055), .B1(P2_REG3_REG_3__SCAN_IN), 
        .B2(n10022), .ZN(n10027) );
  OAI22_X1 U11103 ( .A1(n10025), .A2(n10054), .B1(n10056), .B2(n10024), .ZN(
        n10026) );
  AOI211_X1 U11104 ( .C1(n4281), .C2(P2_REG2_REG_3__SCAN_IN), .A(n10027), .B(
        n10026), .ZN(n10028) );
  OAI21_X1 U11105 ( .B1(n4281), .B2(n10057), .A(n10028), .ZN(P2_U3293) );
  AND2_X1 U11106 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n10035), .ZN(P2_U3297) );
  INV_X1 U11107 ( .A(P2_D_REG_30__SCAN_IN), .ZN(n10174) );
  NOR2_X1 U11108 ( .A1(n10033), .A2(n10174), .ZN(P2_U3298) );
  AND2_X1 U11109 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n10035), .ZN(P2_U3299) );
  AND2_X1 U11110 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n10035), .ZN(P2_U3300) );
  AND2_X1 U11111 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n10035), .ZN(P2_U3301) );
  AND2_X1 U11112 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n10035), .ZN(P2_U3302) );
  AND2_X1 U11113 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n10035), .ZN(P2_U3303) );
  AND2_X1 U11114 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n10035), .ZN(P2_U3304) );
  INV_X1 U11115 ( .A(P2_D_REG_23__SCAN_IN), .ZN(n10198) );
  NOR2_X1 U11116 ( .A1(n10033), .A2(n10198), .ZN(P2_U3305) );
  AND2_X1 U11117 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n10035), .ZN(P2_U3306) );
  AND2_X1 U11118 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n10035), .ZN(P2_U3307) );
  AND2_X1 U11119 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n10035), .ZN(P2_U3308) );
  AND2_X1 U11120 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n10035), .ZN(P2_U3309) );
  AND2_X1 U11121 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n10035), .ZN(P2_U3310) );
  AND2_X1 U11122 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n10035), .ZN(P2_U3311) );
  AND2_X1 U11123 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n10035), .ZN(P2_U3312) );
  INV_X1 U11124 ( .A(P2_D_REG_15__SCAN_IN), .ZN(n10189) );
  NOR2_X1 U11125 ( .A1(n10033), .A2(n10189), .ZN(P2_U3313) );
  AND2_X1 U11126 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n10035), .ZN(P2_U3314) );
  AND2_X1 U11127 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n10035), .ZN(P2_U3315) );
  AND2_X1 U11128 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n10035), .ZN(P2_U3316) );
  AND2_X1 U11129 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n10035), .ZN(P2_U3317) );
  AND2_X1 U11130 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n10035), .ZN(P2_U3318) );
  INV_X1 U11131 ( .A(P2_D_REG_9__SCAN_IN), .ZN(n10226) );
  NOR2_X1 U11132 ( .A1(n10033), .A2(n10226), .ZN(P2_U3319) );
  AND2_X1 U11133 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n10035), .ZN(P2_U3320) );
  AND2_X1 U11134 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n10035), .ZN(P2_U3321) );
  AND2_X1 U11135 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n10035), .ZN(P2_U3322) );
  INV_X1 U11136 ( .A(P2_D_REG_5__SCAN_IN), .ZN(n10185) );
  NOR2_X1 U11137 ( .A1(n10033), .A2(n10185), .ZN(P2_U3323) );
  AND2_X1 U11138 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n10035), .ZN(P2_U3324) );
  AND2_X1 U11139 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n10035), .ZN(P2_U3325) );
  INV_X1 U11140 ( .A(P2_D_REG_2__SCAN_IN), .ZN(n10159) );
  NOR2_X1 U11141 ( .A1(n10033), .A2(n10159), .ZN(P2_U3326) );
  OAI22_X1 U11142 ( .A1(P2_D_REG_0__SCAN_IN), .A2(n10033), .B1(n10032), .B2(
        n10031), .ZN(n10034) );
  INV_X1 U11143 ( .A(n10034), .ZN(P2_U3437) );
  INV_X1 U11144 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n10036) );
  AOI22_X1 U11145 ( .A1(n10038), .A2(n10037), .B1(n10036), .B2(n10035), .ZN(
        P2_U3438) );
  INV_X1 U11146 ( .A(n10039), .ZN(n10045) );
  OAI21_X1 U11147 ( .B1(n10041), .B2(n10077), .A(n10040), .ZN(n10044) );
  INV_X1 U11148 ( .A(n10042), .ZN(n10043) );
  AOI211_X1 U11149 ( .C1(n10086), .C2(n10045), .A(n10044), .B(n10043), .ZN(
        n10093) );
  INV_X1 U11150 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n10046) );
  AOI22_X1 U11151 ( .A1(n10283), .A2(n10093), .B1(n10046), .B2(n10281), .ZN(
        P2_U3454) );
  INV_X1 U11152 ( .A(n10047), .ZN(n10048) );
  OAI211_X1 U11153 ( .C1(n10050), .C2(n10077), .A(n10049), .B(n10048), .ZN(
        n10051) );
  AOI21_X1 U11154 ( .B1(n10086), .B2(n10052), .A(n10051), .ZN(n10094) );
  INV_X1 U11155 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n10053) );
  AOI22_X1 U11156 ( .A1(n10283), .A2(n10094), .B1(n10053), .B2(n10281), .ZN(
        P2_U3457) );
  INV_X1 U11157 ( .A(n10054), .ZN(n10060) );
  OAI21_X1 U11158 ( .B1(n10056), .B2(n10077), .A(n10055), .ZN(n10059) );
  INV_X1 U11159 ( .A(n10057), .ZN(n10058) );
  AOI211_X1 U11160 ( .C1(n10084), .C2(n10060), .A(n10059), .B(n10058), .ZN(
        n10095) );
  INV_X1 U11161 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n10061) );
  AOI22_X1 U11162 ( .A1(n10283), .A2(n10095), .B1(n10061), .B2(n10281), .ZN(
        P2_U3460) );
  NAND2_X1 U11163 ( .A1(n10063), .A2(n10062), .ZN(n10064) );
  AND2_X1 U11164 ( .A1(n10065), .A2(n10064), .ZN(n10068) );
  NAND2_X1 U11165 ( .A1(n10066), .A2(n10086), .ZN(n10067) );
  AND3_X1 U11166 ( .A1(n10069), .A2(n10068), .A3(n10067), .ZN(n10096) );
  INV_X1 U11167 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n10070) );
  AOI22_X1 U11168 ( .A1(n10283), .A2(n10096), .B1(n10070), .B2(n10281), .ZN(
        P2_U3463) );
  OAI22_X1 U11169 ( .A1(n10072), .A2(n4296), .B1(n10071), .B2(n10077), .ZN(
        n10074) );
  AOI211_X1 U11170 ( .C1(n10086), .C2(n10075), .A(n10074), .B(n10073), .ZN(
        n10097) );
  INV_X1 U11171 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10076) );
  AOI22_X1 U11172 ( .A1(n10283), .A2(n10097), .B1(n10076), .B2(n10281), .ZN(
        P2_U3469) );
  OAI22_X1 U11173 ( .A1(n10079), .A2(n4296), .B1(n10078), .B2(n10077), .ZN(
        n10082) );
  INV_X1 U11174 ( .A(n10080), .ZN(n10081) );
  AOI211_X1 U11175 ( .C1(n10084), .C2(n10083), .A(n10082), .B(n10081), .ZN(
        n10099) );
  INV_X1 U11176 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n10188) );
  AOI22_X1 U11177 ( .A1(n10283), .A2(n10099), .B1(n10188), .B2(n10281), .ZN(
        P2_U3481) );
  NAND2_X1 U11178 ( .A1(n10086), .A2(n10085), .ZN(n10087) );
  OAI211_X1 U11179 ( .C1(n10090), .C2(n10089), .A(n10088), .B(n10087), .ZN(
        n10282) );
  OAI22_X1 U11180 ( .A1(n10098), .A2(n10282), .B1(P2_REG1_REG_0__SCAN_IN), 
        .B2(n10100), .ZN(n10091) );
  INV_X1 U11181 ( .A(n10091), .ZN(P2_U3520) );
  AOI22_X1 U11182 ( .A1(n10100), .A2(n10093), .B1(n10092), .B2(n10098), .ZN(
        P2_U3521) );
  AOI22_X1 U11183 ( .A1(n10100), .A2(n10094), .B1(n6729), .B2(n10098), .ZN(
        P2_U3522) );
  AOI22_X1 U11184 ( .A1(n10100), .A2(n10095), .B1(n6730), .B2(n10098), .ZN(
        P2_U3523) );
  AOI22_X1 U11185 ( .A1(n10100), .A2(n10096), .B1(n6732), .B2(n10098), .ZN(
        P2_U3524) );
  AOI22_X1 U11186 ( .A1(n10100), .A2(n10097), .B1(n6734), .B2(n10098), .ZN(
        P2_U3526) );
  AOI22_X1 U11187 ( .A1(n10100), .A2(n10099), .B1(n6940), .B2(n10098), .ZN(
        P2_U3530) );
  INV_X1 U11188 ( .A(n10101), .ZN(n10102) );
  NAND2_X1 U11189 ( .A1(n10103), .A2(n10102), .ZN(n10104) );
  XOR2_X1 U11190 ( .A(n10105), .B(n10104), .Z(ADD_1071_U5) );
  XOR2_X1 U11191 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1071_U46) );
  OAI21_X1 U11192 ( .B1(n10108), .B2(n10107), .A(n10106), .ZN(ADD_1071_U56) );
  OAI21_X1 U11193 ( .B1(n10111), .B2(n10110), .A(n10109), .ZN(ADD_1071_U57) );
  OAI21_X1 U11194 ( .B1(n10114), .B2(n10113), .A(n10112), .ZN(ADD_1071_U58) );
  OAI21_X1 U11195 ( .B1(n10117), .B2(n10116), .A(n10115), .ZN(ADD_1071_U59) );
  OAI21_X1 U11196 ( .B1(n10120), .B2(n10119), .A(n10118), .ZN(ADD_1071_U60) );
  OAI21_X1 U11197 ( .B1(n10123), .B2(n10122), .A(n10121), .ZN(ADD_1071_U61) );
  AOI21_X1 U11198 ( .B1(n10126), .B2(n10125), .A(n10124), .ZN(ADD_1071_U62) );
  AOI21_X1 U11199 ( .B1(n10129), .B2(n10128), .A(n10127), .ZN(ADD_1071_U63) );
  NAND4_X1 U11200 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_D_REG_5__SCAN_IN), .A3(
        P1_ADDR_REG_19__SCAN_IN), .A4(P1_DATAO_REG_16__SCAN_IN), .ZN(n10134)
         );
  NAND4_X1 U11201 ( .A1(P1_DATAO_REG_15__SCAN_IN), .A2(SI_10_), .A3(
        P2_REG0_REG_14__SCAN_IN), .A4(P2_REG2_REG_23__SCAN_IN), .ZN(n10131) );
  NAND4_X1 U11202 ( .A1(P2_DATAO_REG_24__SCAN_IN), .A2(P1_REG1_REG_16__SCAN_IN), .A3(P2_REG3_REG_26__SCAN_IN), .A4(P2_REG3_REG_19__SCAN_IN), .ZN(n10130) );
  NOR3_X1 U11203 ( .A1(P2_REG1_REG_6__SCAN_IN), .A2(n10131), .A3(n10130), .ZN(
        n10132) );
  NAND4_X1 U11204 ( .A1(n10218), .A2(P2_DATAO_REG_27__SCAN_IN), .A3(n10132), 
        .A4(P2_D_REG_9__SCAN_IN), .ZN(n10133) );
  NOR2_X1 U11205 ( .A1(n10134), .A2(n10133), .ZN(n10280) );
  NAND4_X1 U11206 ( .A1(P1_D_REG_4__SCAN_IN), .A2(P2_B_REG_SCAN_IN), .A3(
        P2_REG0_REG_16__SCAN_IN), .A4(P2_REG0_REG_7__SCAN_IN), .ZN(n10137) );
  NAND4_X1 U11207 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(n7711), .A3(n10187), .A4(
        n10188), .ZN(n10136) );
  NAND3_X1 U11208 ( .A1(P1_D_REG_21__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .A3(n6730), .ZN(n10135) );
  NOR4_X1 U11209 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(n10137), .A3(n10136), .A4(
        n10135), .ZN(n10154) );
  NAND3_X1 U11210 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(P1_REG2_REG_7__SCAN_IN), 
        .A3(n10263), .ZN(n10140) );
  INV_X1 U11211 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n10250) );
  NAND4_X1 U11212 ( .A1(SI_22_), .A2(P1_D_REG_15__SCAN_IN), .A3(
        P1_REG3_REG_9__SCAN_IN), .A4(n10250), .ZN(n10139) );
  NAND4_X1 U11213 ( .A1(P2_REG0_REG_26__SCAN_IN), .A2(n10254), .A3(n10257), 
        .A4(n10253), .ZN(n10138) );
  NOR4_X1 U11214 ( .A1(SI_1_), .A2(n10140), .A3(n10139), .A4(n10138), .ZN(
        n10153) );
  NOR4_X1 U11215 ( .A1(P2_D_REG_23__SCAN_IN), .A2(SI_11_), .A3(
        P2_REG2_REG_16__SCAN_IN), .A4(n10205), .ZN(n10151) );
  NAND4_X1 U11216 ( .A1(n10141), .A2(n10238), .A3(n10164), .A4(SI_13_), .ZN(
        n10147) );
  NAND4_X1 U11217 ( .A1(n10142), .A2(P2_IR_REG_31__SCAN_IN), .A3(
        P2_REG3_REG_24__SCAN_IN), .A4(P2_REG3_REG_17__SCAN_IN), .ZN(n10146) );
  NOR4_X1 U11218 ( .A1(P1_REG1_REG_29__SCAN_IN), .A2(P2_REG1_REG_29__SCAN_IN), 
        .A3(n6827), .A4(n10165), .ZN(n10143) );
  NAND3_X1 U11219 ( .A1(n10144), .A2(P2_D_REG_30__SCAN_IN), .A3(n10143), .ZN(
        n10145) );
  NOR3_X1 U11220 ( .A1(n10147), .A2(n10146), .A3(n10145), .ZN(n10149) );
  AND4_X1 U11221 ( .A1(P2_D_REG_2__SCAN_IN), .A2(P1_ADDR_REG_5__SCAN_IN), .A3(
        n10157), .A4(n10156), .ZN(n10148) );
  AND4_X1 U11222 ( .A1(n10151), .A2(n10150), .A3(n10149), .A4(n10148), .ZN(
        n10152) );
  AND3_X1 U11223 ( .A1(n10154), .A2(n10153), .A3(n10152), .ZN(n10279) );
  AOI22_X1 U11224 ( .A1(n10157), .A2(keyinput47), .B1(n10156), .B2(keyinput59), 
        .ZN(n10155) );
  OAI221_X1 U11225 ( .B1(n10157), .B2(keyinput47), .C1(n10156), .C2(keyinput59), .A(n10155), .ZN(n10169) );
  AOI22_X1 U11226 ( .A1(n10159), .A2(keyinput62), .B1(keyinput51), .B2(n6827), 
        .ZN(n10158) );
  OAI221_X1 U11227 ( .B1(n10159), .B2(keyinput62), .C1(n6827), .C2(keyinput51), 
        .A(n10158), .ZN(n10168) );
  INV_X1 U11228 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n10162) );
  AOI22_X1 U11229 ( .A1(n10162), .A2(keyinput55), .B1(keyinput19), .B2(n10161), 
        .ZN(n10160) );
  OAI221_X1 U11230 ( .B1(n10162), .B2(keyinput55), .C1(n10161), .C2(keyinput19), .A(n10160), .ZN(n10167) );
  AOI22_X1 U11231 ( .A1(n10165), .A2(keyinput3), .B1(n10164), .B2(keyinput39), 
        .ZN(n10163) );
  OAI221_X1 U11232 ( .B1(n10165), .B2(keyinput3), .C1(n10164), .C2(keyinput39), 
        .A(n10163), .ZN(n10166) );
  NOR4_X1 U11233 ( .A1(n10169), .A2(n10168), .A3(n10167), .A4(n10166), .ZN(
        n10215) );
  INV_X1 U11234 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n10171) );
  AOI22_X1 U11235 ( .A1(n10171), .A2(keyinput2), .B1(keyinput61), .B2(n7711), 
        .ZN(n10170) );
  OAI221_X1 U11236 ( .B1(n10171), .B2(keyinput2), .C1(n7711), .C2(keyinput61), 
        .A(n10170), .ZN(n10183) );
  AOI22_X1 U11237 ( .A1(n10174), .A2(keyinput23), .B1(n10173), .B2(keyinput38), 
        .ZN(n10172) );
  OAI221_X1 U11238 ( .B1(n10174), .B2(keyinput23), .C1(n10173), .C2(keyinput38), .A(n10172), .ZN(n10182) );
  AOI22_X1 U11239 ( .A1(n10177), .A2(keyinput20), .B1(n10176), .B2(keyinput15), 
        .ZN(n10175) );
  OAI221_X1 U11240 ( .B1(n10177), .B2(keyinput20), .C1(n10176), .C2(keyinput15), .A(n10175), .ZN(n10181) );
  XNOR2_X1 U11241 ( .A(P1_IR_REG_23__SCAN_IN), .B(keyinput56), .ZN(n10179) );
  XNOR2_X1 U11242 ( .A(SI_13_), .B(keyinput26), .ZN(n10178) );
  NAND2_X1 U11243 ( .A1(n10179), .A2(n10178), .ZN(n10180) );
  NOR4_X1 U11244 ( .A1(n10183), .A2(n10182), .A3(n10181), .A4(n10180), .ZN(
        n10214) );
  AOI22_X1 U11245 ( .A1(n10185), .A2(keyinput6), .B1(keyinput40), .B2(n6727), 
        .ZN(n10184) );
  OAI221_X1 U11246 ( .B1(n10185), .B2(keyinput6), .C1(n6727), .C2(keyinput40), 
        .A(n10184), .ZN(n10196) );
  AOI22_X1 U11247 ( .A1(n10188), .A2(keyinput8), .B1(n10187), .B2(keyinput13), 
        .ZN(n10186) );
  OAI221_X1 U11248 ( .B1(n10188), .B2(keyinput8), .C1(n10187), .C2(keyinput13), 
        .A(n10186), .ZN(n10195) );
  XNOR2_X1 U11249 ( .A(n10189), .B(keyinput28), .ZN(n10194) );
  XOR2_X1 U11250 ( .A(n6730), .B(keyinput50), .Z(n10192) );
  XNOR2_X1 U11251 ( .A(P1_IR_REG_22__SCAN_IN), .B(keyinput4), .ZN(n10191) );
  XNOR2_X1 U11252 ( .A(P1_IR_REG_5__SCAN_IN), .B(keyinput36), .ZN(n10190) );
  NAND3_X1 U11253 ( .A1(n10192), .A2(n10191), .A3(n10190), .ZN(n10193) );
  NOR4_X1 U11254 ( .A1(n10196), .A2(n10195), .A3(n10194), .A4(n10193), .ZN(
        n10213) );
  AOI22_X1 U11255 ( .A1(n10199), .A2(keyinput63), .B1(keyinput21), .B2(n10198), 
        .ZN(n10197) );
  OAI221_X1 U11256 ( .B1(n10199), .B2(keyinput63), .C1(n10198), .C2(keyinput21), .A(n10197), .ZN(n10211) );
  INV_X1 U11257 ( .A(SI_11_), .ZN(n10202) );
  INV_X1 U11258 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n10201) );
  AOI22_X1 U11259 ( .A1(n10202), .A2(keyinput57), .B1(keyinput14), .B2(n10201), 
        .ZN(n10200) );
  OAI221_X1 U11260 ( .B1(n10202), .B2(keyinput57), .C1(n10201), .C2(keyinput14), .A(n10200), .ZN(n10210) );
  AOI22_X1 U11261 ( .A1(n10205), .A2(keyinput53), .B1(keyinput27), .B2(n10204), 
        .ZN(n10203) );
  OAI221_X1 U11262 ( .B1(n10205), .B2(keyinput53), .C1(n10204), .C2(keyinput27), .A(n10203), .ZN(n10209) );
  XNOR2_X1 U11263 ( .A(P2_REG2_REG_16__SCAN_IN), .B(keyinput35), .ZN(n10207)
         );
  XNOR2_X1 U11264 ( .A(P2_IR_REG_21__SCAN_IN), .B(keyinput41), .ZN(n10206) );
  NAND2_X1 U11265 ( .A1(n10207), .A2(n10206), .ZN(n10208) );
  NOR4_X1 U11266 ( .A1(n10211), .A2(n10210), .A3(n10209), .A4(n10208), .ZN(
        n10212) );
  NAND4_X1 U11267 ( .A1(n10215), .A2(n10214), .A3(n10213), .A4(n10212), .ZN(
        n10278) );
  XNOR2_X1 U11268 ( .A(n10216), .B(keyinput43), .ZN(n10221) );
  XNOR2_X1 U11269 ( .A(n10217), .B(keyinput7), .ZN(n10220) );
  XNOR2_X1 U11270 ( .A(n10218), .B(keyinput1), .ZN(n10219) );
  NOR3_X1 U11271 ( .A1(n10221), .A2(n10220), .A3(n10219), .ZN(n10224) );
  XNOR2_X1 U11272 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(keyinput25), .ZN(n10223)
         );
  XNOR2_X1 U11273 ( .A(P1_ADDR_REG_19__SCAN_IN), .B(keyinput58), .ZN(n10222)
         );
  NAND3_X1 U11274 ( .A1(n10224), .A2(n10223), .A3(n10222), .ZN(n10230) );
  AOI22_X1 U11275 ( .A1(n10226), .A2(keyinput22), .B1(keyinput60), .B2(n6734), 
        .ZN(n10225) );
  OAI221_X1 U11276 ( .B1(n10226), .B2(keyinput22), .C1(n6734), .C2(keyinput60), 
        .A(n10225), .ZN(n10229) );
  XNOR2_X1 U11277 ( .A(n10227), .B(keyinput42), .ZN(n10228) );
  NOR3_X1 U11278 ( .A1(n10230), .A2(n10229), .A3(n10228), .ZN(n10276) );
  AOI22_X1 U11279 ( .A1(n10233), .A2(keyinput52), .B1(n10232), .B2(keyinput29), 
        .ZN(n10231) );
  OAI221_X1 U11280 ( .B1(n10233), .B2(keyinput52), .C1(n10232), .C2(keyinput29), .A(n10231), .ZN(n10245) );
  AOI22_X1 U11281 ( .A1(n10235), .A2(keyinput34), .B1(keyinput44), .B2(n8284), 
        .ZN(n10234) );
  OAI221_X1 U11282 ( .B1(n10235), .B2(keyinput34), .C1(n8284), .C2(keyinput44), 
        .A(n10234), .ZN(n10244) );
  AOI22_X1 U11283 ( .A1(n10238), .A2(keyinput37), .B1(keyinput33), .B2(n10237), 
        .ZN(n10236) );
  OAI221_X1 U11284 ( .B1(n10238), .B2(keyinput37), .C1(n10237), .C2(keyinput33), .A(n10236), .ZN(n10243) );
  AOI22_X1 U11285 ( .A1(n10241), .A2(keyinput16), .B1(n10240), .B2(keyinput30), 
        .ZN(n10239) );
  OAI221_X1 U11286 ( .B1(n10241), .B2(keyinput16), .C1(n10240), .C2(keyinput30), .A(n10239), .ZN(n10242) );
  NOR4_X1 U11287 ( .A1(n10245), .A2(n10244), .A3(n10243), .A4(n10242), .ZN(
        n10275) );
  AOI22_X1 U11288 ( .A1(n10248), .A2(keyinput0), .B1(n10247), .B2(keyinput9), 
        .ZN(n10246) );
  OAI221_X1 U11289 ( .B1(n10248), .B2(keyinput0), .C1(n10247), .C2(keyinput9), 
        .A(n10246), .ZN(n10261) );
  AOI22_X1 U11290 ( .A1(n10251), .A2(keyinput11), .B1(keyinput46), .B2(n10250), 
        .ZN(n10249) );
  OAI221_X1 U11291 ( .B1(n10251), .B2(keyinput11), .C1(n10250), .C2(keyinput46), .A(n10249), .ZN(n10260) );
  AOI22_X1 U11292 ( .A1(n10254), .A2(keyinput18), .B1(keyinput45), .B2(n10253), 
        .ZN(n10252) );
  OAI221_X1 U11293 ( .B1(n10254), .B2(keyinput18), .C1(n10253), .C2(keyinput45), .A(n10252), .ZN(n10259) );
  AOI22_X1 U11294 ( .A1(n10257), .A2(keyinput24), .B1(keyinput49), .B2(n10256), 
        .ZN(n10255) );
  OAI221_X1 U11295 ( .B1(n10257), .B2(keyinput24), .C1(n10256), .C2(keyinput49), .A(n10255), .ZN(n10258) );
  NOR4_X1 U11296 ( .A1(n10261), .A2(n10260), .A3(n10259), .A4(n10258), .ZN(
        n10274) );
  AOI22_X1 U11297 ( .A1(n7315), .A2(keyinput31), .B1(n10263), .B2(keyinput48), 
        .ZN(n10262) );
  OAI221_X1 U11298 ( .B1(n7315), .B2(keyinput31), .C1(n10263), .C2(keyinput48), 
        .A(n10262), .ZN(n10272) );
  AOI22_X1 U11299 ( .A1(n10265), .A2(keyinput12), .B1(keyinput17), .B2(n4585), 
        .ZN(n10264) );
  OAI221_X1 U11300 ( .B1(n10265), .B2(keyinput12), .C1(n4585), .C2(keyinput17), 
        .A(n10264), .ZN(n10271) );
  XNOR2_X1 U11301 ( .A(SI_1_), .B(keyinput32), .ZN(n10269) );
  XNOR2_X1 U11302 ( .A(P1_IR_REG_28__SCAN_IN), .B(keyinput54), .ZN(n10268) );
  XNOR2_X1 U11303 ( .A(P2_IR_REG_31__SCAN_IN), .B(keyinput5), .ZN(n10267) );
  XNOR2_X1 U11304 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(keyinput10), .ZN(n10266)
         );
  NAND4_X1 U11305 ( .A1(n10269), .A2(n10268), .A3(n10267), .A4(n10266), .ZN(
        n10270) );
  NOR3_X1 U11306 ( .A1(n10272), .A2(n10271), .A3(n10270), .ZN(n10273) );
  NAND4_X1 U11307 ( .A1(n10276), .A2(n10275), .A3(n10274), .A4(n10273), .ZN(
        n10277) );
  AOI211_X1 U11308 ( .C1(n10280), .C2(n10279), .A(n10278), .B(n10277), .ZN(
        n10285) );
  AOI22_X1 U11309 ( .A1(n10283), .A2(n10282), .B1(P2_REG0_REG_0__SCAN_IN), 
        .B2(n10281), .ZN(n10284) );
  XNOR2_X1 U11310 ( .A(n10285), .B(n10284), .ZN(P2_U3451) );
  XOR2_X1 U11311 ( .A(n10286), .B(P2_ADDR_REG_6__SCAN_IN), .Z(ADD_1071_U50) );
  NOR2_X1 U11312 ( .A1(n10288), .A2(n10287), .ZN(n10289) );
  XOR2_X1 U11313 ( .A(n10289), .B(P1_ADDR_REG_5__SCAN_IN), .Z(ADD_1071_U51) );
  XOR2_X1 U11314 ( .A(n10290), .B(P2_ADDR_REG_7__SCAN_IN), .Z(ADD_1071_U49) );
  OAI21_X1 U11315 ( .B1(n10293), .B2(n10292), .A(n10291), .ZN(n10294) );
  XNOR2_X1 U11316 ( .A(n10294), .B(P1_ADDR_REG_18__SCAN_IN), .ZN(ADD_1071_U55)
         );
  XOR2_X1 U11317 ( .A(n10295), .B(P2_ADDR_REG_8__SCAN_IN), .Z(ADD_1071_U48) );
  AOI21_X1 U11318 ( .B1(n10298), .B2(n10297), .A(n10296), .ZN(ADD_1071_U47) );
  XOR2_X1 U11319 ( .A(n10300), .B(n10299), .Z(ADD_1071_U54) );
  XOR2_X1 U11320 ( .A(n10301), .B(n10302), .Z(ADD_1071_U53) );
  XNOR2_X1 U11321 ( .A(n10304), .B(n10303), .ZN(ADD_1071_U52) );
  NAND2_X1 U4781 ( .A1(n5946), .A2(n5947), .ZN(n7737) );
  AND2_X1 U4793 ( .A1(n5874), .A2(n5850), .ZN(n4649) );
  CLKBUF_X1 U4795 ( .A(n5451), .Z(n4491) );
  CLKBUF_X1 U4836 ( .A(n5452), .Z(n4492) );
  CLKBUF_X2 U4837 ( .A(n5870), .Z(n4292) );
  CLKBUF_X1 U4865 ( .A(n8709), .Z(n4463) );
  CLKBUF_X1 U5028 ( .A(n7004), .Z(n4299) );
  CLKBUF_X1 U5168 ( .A(n7253), .Z(n8775) );
  CLKBUF_X2 U5301 ( .A(n5870), .Z(n4293) );
  CLKBUF_X1 U5309 ( .A(n6000), .Z(n4417) );
  CLKBUF_X1 U5687 ( .A(n8382), .Z(n4454) );
  NAND2_X1 U5785 ( .A1(n7733), .A2(n7744), .ZN(n7771) );
  CLKBUF_X1 U6291 ( .A(n8352), .Z(n4291) );
  CLKBUF_X1 U6505 ( .A(n5751), .Z(n6893) );
endmodule

