

module b20_C_gen_AntiSAT_k_128_10 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, keyinput_f0, 
        keyinput_f1, keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5, 
        keyinput_f6, keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10, 
        keyinput_f11, keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15, 
        keyinput_f16, keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20, 
        keyinput_f21, keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25, 
        keyinput_f26, keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30, 
        keyinput_f31, keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35, 
        keyinput_f36, keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40, 
        keyinput_f41, keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45, 
        keyinput_f46, keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50, 
        keyinput_f51, keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55, 
        keyinput_f56, keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60, 
        keyinput_f61, keyinput_f62, keyinput_f63, keyinput_g0, keyinput_g1, 
        keyinput_g2, keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, 
        keyinput_g7, keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, 
        keyinput_g12, keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, 
        keyinput_g17, keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, 
        keyinput_g22, keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, 
        keyinput_g27, keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, 
        keyinput_g32, keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, 
        keyinput_g37, keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, 
        keyinput_g42, keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, 
        keyinput_g47, keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, 
        keyinput_g52, keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, 
        keyinput_g57, keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, 
        keyinput_g62, keyinput_g63, ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, 
        ADD_1068_U57, ADD_1068_U58, ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, 
        ADD_1068_U62, ADD_1068_U63, ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, 
        ADD_1068_U50, ADD_1068_U51, ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, 
        ADD_1068_U5, ADD_1068_U46, U126, U123, P1_U3355, P1_U3354, P1_U3353, 
        P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, 
        P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, 
        P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, 
        P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, 
        P1_U3324, P1_U3439, P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, 
        P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, 
        P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, 
        P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, 
        P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, 
        P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, 
        P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, 
        P1_U3501, P1_U3504, P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, 
        P1_U3513, P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, 
        P1_U3520, P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, 
        P1_U3527, P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, 
        P1_U3534, P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, 
        P1_U3541, P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, 
        P1_U3548, P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, 
        P1_U3292, P1_U3291, P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, 
        P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, 
        P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, 
        P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, 
        P1_U3356, P1_U3264, P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, 
        P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, 
        P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, 
        P1_U3244, P1_U3243, P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, 
        P1_U3559, P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, 
        P1_U3566, P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, 
        P1_U3573, P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, 
        P1_U3580, P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, 
        P1_U3241, P1_U3240, P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, 
        P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, 
        P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, 
        P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, 
        P1_U3213, P1_U3086, P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, 
        P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, 
        P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, 
        P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, 
        P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, 
        P2_U3264, P2_U3376, P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, 
        P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, 
        P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, 
        P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, 
        P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, 
        P2_U3396, P2_U3399, P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, 
        P2_U3417, P2_U3420, P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, 
        P2_U3438, P2_U3441, P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, 
        P2_U3450, P2_U3451, P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, 
        P2_U3457, P2_U3458, P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, 
        P2_U3464, P2_U3465, P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, 
        P2_U3471, P2_U3472, P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, 
        P2_U3478, P2_U3479, P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, 
        P2_U3485, P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, 
        P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, 
        P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, 
        P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, 
        P2_U3211, P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, 
        P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, 
        P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, 
        P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, 
        P2_U3183, P2_U3182, P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, 
        P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, 
        P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, 
        P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, 
        P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, 
        P2_U3181, P2_U3180, P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, 
        P2_U3174, P2_U3173, P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, 
        P2_U3167, P2_U3166, P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, 
        P2_U3160, P2_U3159, P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, 
        P2_U3153, P2_U3151, P2_U3150, P2_U3893 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, keyinput_f0, keyinput_f1, keyinput_f2,
         keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, keyinput_f7,
         keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, keyinput_f12,
         keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, keyinput_f17,
         keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, keyinput_f22,
         keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, keyinput_f27,
         keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, keyinput_f32,
         keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, keyinput_f37,
         keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, keyinput_f42,
         keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, keyinput_f47,
         keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, keyinput_f52,
         keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, keyinput_f57,
         keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, keyinput_f62,
         keyinput_f63, keyinput_g0, keyinput_g1, keyinput_g2, keyinput_g3,
         keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7, keyinput_g8,
         keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12, keyinput_g13,
         keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17, keyinput_g18,
         keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22, keyinput_g23,
         keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27, keyinput_g28,
         keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32, keyinput_g33,
         keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37, keyinput_g38,
         keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42, keyinput_g43,
         keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47, keyinput_g48,
         keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52, keyinput_g53,
         keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57, keyinput_g58,
         keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62, keyinput_g63;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354,
         n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364,
         n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374,
         n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384,
         n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394,
         n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404,
         n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414,
         n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424,
         n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434,
         n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444,
         n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454,
         n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464,
         n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474,
         n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484,
         n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494,
         n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504,
         n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514,
         n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524,
         n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534,
         n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544,
         n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554,
         n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564,
         n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574,
         n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584,
         n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594,
         n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604,
         n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614,
         n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624,
         n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634,
         n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644,
         n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654,
         n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664,
         n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674,
         n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684,
         n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694,
         n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704,
         n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714,
         n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724,
         n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734,
         n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744,
         n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754,
         n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764,
         n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774,
         n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784,
         n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794,
         n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804,
         n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814,
         n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824,
         n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834,
         n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844,
         n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854,
         n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864,
         n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874,
         n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884,
         n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894,
         n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904,
         n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914,
         n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924,
         n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934,
         n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944,
         n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954,
         n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964,
         n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974,
         n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984,
         n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994,
         n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004,
         n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014,
         n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024,
         n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034,
         n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044,
         n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054,
         n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064,
         n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074,
         n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084,
         n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094,
         n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104,
         n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114,
         n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124,
         n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134,
         n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144,
         n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154,
         n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164,
         n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174,
         n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184,
         n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194,
         n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204,
         n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214,
         n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224,
         n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234,
         n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244,
         n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254,
         n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264,
         n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274,
         n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284,
         n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294,
         n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304,
         n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314,
         n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324,
         n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334,
         n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344,
         n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354,
         n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364,
         n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374,
         n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384,
         n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394,
         n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404,
         n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414,
         n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424,
         n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434,
         n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444,
         n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454,
         n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464,
         n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474,
         n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484,
         n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494,
         n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504,
         n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514,
         n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524,
         n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534,
         n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544,
         n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554,
         n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564,
         n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574,
         n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584,
         n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594,
         n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604,
         n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614,
         n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624,
         n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634,
         n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644,
         n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654,
         n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664,
         n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674,
         n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684,
         n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694,
         n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704,
         n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714,
         n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724,
         n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734,
         n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744,
         n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754,
         n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764,
         n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774,
         n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784,
         n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794,
         n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804,
         n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814,
         n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824,
         n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834,
         n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844,
         n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854,
         n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864,
         n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874,
         n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884,
         n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894,
         n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904,
         n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914,
         n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924,
         n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934,
         n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944,
         n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954,
         n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964,
         n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974,
         n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984,
         n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994,
         n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004,
         n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014,
         n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024,
         n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034,
         n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044,
         n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054,
         n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064,
         n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074,
         n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084,
         n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094,
         n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104,
         n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114,
         n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124,
         n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134,
         n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144,
         n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154,
         n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164,
         n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174,
         n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184,
         n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194,
         n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204,
         n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214,
         n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224,
         n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234,
         n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244,
         n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254,
         n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264,
         n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274,
         n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284,
         n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294,
         n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304,
         n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314,
         n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324,
         n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334,
         n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344,
         n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354,
         n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364,
         n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374,
         n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384,
         n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394,
         n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404,
         n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414,
         n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424,
         n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434,
         n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444,
         n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454,
         n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464,
         n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474,
         n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484,
         n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494,
         n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504,
         n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514,
         n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524,
         n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534,
         n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544,
         n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554,
         n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564,
         n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574,
         n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584,
         n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594,
         n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604,
         n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614,
         n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624,
         n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634,
         n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644,
         n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654,
         n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664,
         n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674,
         n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684,
         n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694,
         n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704,
         n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714,
         n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724,
         n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734,
         n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744,
         n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754,
         n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764,
         n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774,
         n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784,
         n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794,
         n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804,
         n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814,
         n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824,
         n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834,
         n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844,
         n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854,
         n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864,
         n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874,
         n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884,
         n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894,
         n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904,
         n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914,
         n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924,
         n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934,
         n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944,
         n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954,
         n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964,
         n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974,
         n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984,
         n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994,
         n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004,
         n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014,
         n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024,
         n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034,
         n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044,
         n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054,
         n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064,
         n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074,
         n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084,
         n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094,
         n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104,
         n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114,
         n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124,
         n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134,
         n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144,
         n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154,
         n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164,
         n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174,
         n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184,
         n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194,
         n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204,
         n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214,
         n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224,
         n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234,
         n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244,
         n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254,
         n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264,
         n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274,
         n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284,
         n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294,
         n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304,
         n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314,
         n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324,
         n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334,
         n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344,
         n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354,
         n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364,
         n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374,
         n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384,
         n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394,
         n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404,
         n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414,
         n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424,
         n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434,
         n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444,
         n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454,
         n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464,
         n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474,
         n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484,
         n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494,
         n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504,
         n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514,
         n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524,
         n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534,
         n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544,
         n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554,
         n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564,
         n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574,
         n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584,
         n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594,
         n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604,
         n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614,
         n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624,
         n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634,
         n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644,
         n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654,
         n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664,
         n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674,
         n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684,
         n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694,
         n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704,
         n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714,
         n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724,
         n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734,
         n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744,
         n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754,
         n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764,
         n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774,
         n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784,
         n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794,
         n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804,
         n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814,
         n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824,
         n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834,
         n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844,
         n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854,
         n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864,
         n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874,
         n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884,
         n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894,
         n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904,
         n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914,
         n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924,
         n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934,
         n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944,
         n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954,
         n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964,
         n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974,
         n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984,
         n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994,
         n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004,
         n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014,
         n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024,
         n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034,
         n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044,
         n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054,
         n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064,
         n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074,
         n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084,
         n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094,
         n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104,
         n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114,
         n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124,
         n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134,
         n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144,
         n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154,
         n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164,
         n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174,
         n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184,
         n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194,
         n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204,
         n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214,
         n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224,
         n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234,
         n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244,
         n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254,
         n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264,
         n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274,
         n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284,
         n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294,
         n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304,
         n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314,
         n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324,
         n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334,
         n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344,
         n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354,
         n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364,
         n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374,
         n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384,
         n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394,
         n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404,
         n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414,
         n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424,
         n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434,
         n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444,
         n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454,
         n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464,
         n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474,
         n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484,
         n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494,
         n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504,
         n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514,
         n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524,
         n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534,
         n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544,
         n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554,
         n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564,
         n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574,
         n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584,
         n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594,
         n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604,
         n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614,
         n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624,
         n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634,
         n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644,
         n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654,
         n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664,
         n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674,
         n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684,
         n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694,
         n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704,
         n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714,
         n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724,
         n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734,
         n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744,
         n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754,
         n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764,
         n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774,
         n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784,
         n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794,
         n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804,
         n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814,
         n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824,
         n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834,
         n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844,
         n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854,
         n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864,
         n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874,
         n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884,
         n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894,
         n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904,
         n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914,
         n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924,
         n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934,
         n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944,
         n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954,
         n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964,
         n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974,
         n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984,
         n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994,
         n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004,
         n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014,
         n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024,
         n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034,
         n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044,
         n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054,
         n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064,
         n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074,
         n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084,
         n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094,
         n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104,
         n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114,
         n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124,
         n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134,
         n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144,
         n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154,
         n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164,
         n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174,
         n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184,
         n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194,
         n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204,
         n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214,
         n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224,
         n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234,
         n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244,
         n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254,
         n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264,
         n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274,
         n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284,
         n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294,
         n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304,
         n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314,
         n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324,
         n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334,
         n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344,
         n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354,
         n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364,
         n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374,
         n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384,
         n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394,
         n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404,
         n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414,
         n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424,
         n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434,
         n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444,
         n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454,
         n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464,
         n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474,
         n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484,
         n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494,
         n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504,
         n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514,
         n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524,
         n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534,
         n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544,
         n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554,
         n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564,
         n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574,
         n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584,
         n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594,
         n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604,
         n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614,
         n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624,
         n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634,
         n9635, n9636, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645,
         n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655,
         n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665,
         n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675,
         n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685,
         n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695,
         n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705,
         n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715,
         n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725,
         n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735,
         n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745,
         n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755,
         n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765,
         n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775,
         n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785,
         n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795,
         n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805,
         n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815,
         n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825,
         n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835,
         n9836, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846,
         n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856,
         n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866,
         n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876,
         n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886,
         n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896,
         n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906,
         n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916,
         n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926,
         n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936,
         n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946,
         n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956,
         n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966,
         n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976,
         n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986,
         n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996,
         n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005,
         n10006, n10007, n10008, n10009, n10010, n10011, n10012, n10013,
         n10014, n10015, n10016, n10017, n10018, n10019, n10020, n10021,
         n10022, n10023, n10024, n10025, n10026, n10027, n10028, n10029,
         n10030, n10031, n10032, n10033, n10034, n10035, n10036, n10037,
         n10038, n10039, n10040, n10041, n10042, n10043, n10044, n10045,
         n10046, n10047, n10048, n10049, n10050, n10051, n10052, n10053,
         n10054, n10055, n10056, n10057, n10058, n10059, n10060, n10061,
         n10062, n10063, n10064, n10065, n10066, n10067, n10068, n10069,
         n10070, n10071, n10072, n10073, n10074, n10075, n10076, n10077,
         n10078, n10079, n10080, n10081, n10082, n10083, n10084, n10085,
         n10086, n10087, n10088, n10089, n10090, n10091, n10092, n10093,
         n10094, n10095, n10096, n10097, n10098, n10099, n10100, n10101,
         n10102, n10103, n10104, n10105, n10106, n10107, n10108, n10109,
         n10110, n10111, n10112, n10113, n10114, n10115, n10116, n10117,
         n10118, n10119, n10120, n10121, n10122, n10123, n10124, n10125,
         n10126, n10127, n10128, n10129, n10130, n10131, n10132, n10133,
         n10134, n10135, n10136, n10137, n10138, n10139, n10140, n10141,
         n10142, n10143, n10144, n10145, n10146, n10147, n10148, n10149,
         n10150, n10151, n10152, n10153, n10154, n10155, n10156, n10157,
         n10158, n10159, n10160, n10161, n10162, n10163, n10164, n10165,
         n10166, n10167, n10168, n10169, n10170, n10171, n10172, n10173,
         n10174, n10175, n10176, n10177, n10178, n10179, n10180, n10181,
         n10182, n10183, n10184, n10185, n10186, n10187, n10188, n10189,
         n10190, n10191, n10192, n10196;

  AOI21_X1 U4850 ( .B1(n9229), .B2(n9821), .A(n9228), .ZN(n9391) );
  INV_X1 U4851 ( .A(n9861), .ZN(n8210) );
  NAND2_X1 U4852 ( .A1(n6075), .A2(n4349), .ZN(n8322) );
  CLKBUF_X2 U4853 ( .A(n6074), .Z(n4349) );
  INV_X1 U4854 ( .A(n6064), .ZN(n6749) );
  NAND2_X1 U4855 ( .A1(n5925), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5969) );
  INV_X1 U4856 ( .A(n6262), .ZN(n7282) );
  INV_X2 U4857 ( .A(n7941), .ZN(n7731) );
  CLKBUF_X2 U4858 ( .A(n5219), .Z(n8107) );
  NOR2_X1 U4859 ( .A1(n5508), .A2(P2_IR_REG_21__SCAN_IN), .ZN(n5561) );
  INV_X1 U4861 ( .A(n10196), .ZN(n4345) );
  INV_X1 U4862 ( .A(n7949), .ZN(n7922) );
  NOR2_X1 U4863 ( .A1(n7685), .A2(n7684), .ZN(n7692) );
  CLKBUF_X3 U4864 ( .A(n6204), .Z(n4347) );
  OAI211_X1 U4865 ( .C1(n8173), .C2(n9585), .A(n6181), .B(n6180), .ZN(n6615)
         );
  AND2_X1 U4866 ( .A1(n8559), .A2(n7816), .ZN(n7819) );
  NAND2_X1 U4867 ( .A1(n7576), .A2(n7482), .ZN(n5120) );
  NAND2_X1 U4868 ( .A1(n7576), .A2(n4917), .ZN(n5219) );
  INV_X1 U4869 ( .A(n4347), .ZN(n7714) );
  INV_X1 U4870 ( .A(n6642), .ZN(n6643) );
  INV_X1 U4871 ( .A(n6615), .ZN(n6626) );
  NAND2_X1 U4872 ( .A1(n5375), .A2(n5374), .ZN(n8852) );
  NOR2_X1 U4873 ( .A1(n5510), .A2(n5561), .ZN(n7979) );
  NAND2_X1 U4874 ( .A1(n7432), .A2(n7431), .ZN(n9454) );
  XNOR2_X1 U4875 ( .A(n5448), .B(n5447), .ZN(n7853) );
  XNOR2_X1 U4876 ( .A(n5969), .B(n5968), .ZN(n6075) );
  AND2_X1 U4877 ( .A1(n5069), .A2(n4962), .ZN(n5093) );
  NAND2_X1 U4878 ( .A1(n6158), .A2(n7949), .ZN(n4346) );
  NAND2_X2 U4879 ( .A1(n6158), .A2(n7949), .ZN(n6252) );
  NAND2_X1 U4880 ( .A1(n8173), .A2(n5052), .ZN(n6204) );
  XNOR2_X2 U4881 ( .A(n4935), .B(n4695), .ZN(n4934) );
  NAND2_X2 U4882 ( .A1(n4931), .A2(n4930), .ZN(n4935) );
  NOR2_X2 U4883 ( .A1(n7488), .A2(n8376), .ZN(n7641) );
  OAI22_X2 U4884 ( .A1(n9547), .A2(n4830), .B1(n4832), .B2(n8437), .ZN(n7488)
         );
  XNOR2_X2 U4885 ( .A(n4954), .B(SI_4_), .ZN(n5125) );
  XNOR2_X2 U4886 ( .A(n4687), .B(n4914), .ZN(n4918) );
  AOI21_X2 U4887 ( .B1(n8090), .B2(n8092), .A(n8093), .ZN(n8101) );
  OAI21_X1 U4888 ( .B1(n5606), .B2(n8134), .A(n5605), .ZN(n4348) );
  OAI21_X2 U4889 ( .B1(n5304), .B2(n4758), .A(n4756), .ZN(n5319) );
  INV_X4 U4890 ( .A(n5069), .ZN(n5127) );
  AOI21_X1 U4891 ( .B1(n4521), .B2(n4373), .A(n4519), .ZN(n8089) );
  INV_X1 U4892 ( .A(n8946), .ZN(n4544) );
  NAND2_X1 U4893 ( .A1(n5360), .A2(n5359), .ZN(n8928) );
  NAND2_X1 U4894 ( .A1(n5385), .A2(n5002), .ZN(n5010) );
  NAND2_X1 U4895 ( .A1(n6655), .A2(n6654), .ZN(n7141) );
  INV_X2 U4896 ( .A(n8322), .ZN(n8264) );
  NOR2_X1 U4897 ( .A1(n9081), .A2(n9830), .ZN(n9813) );
  INV_X4 U4898 ( .A(n7948), .ZN(n7709) );
  NAND4_X1 U4899 ( .A1(n5124), .A2(n5123), .A3(n5122), .A4(n5121), .ZN(n8600)
         );
  OR2_X1 U4900 ( .A1(n6204), .A2(n6179), .ZN(n6180) );
  CLKBUF_X1 U4901 ( .A(n6003), .Z(n6001) );
  NAND2_X2 U4902 ( .A1(n6484), .A2(n9567), .ZN(n8173) );
  NAND2_X1 U4903 ( .A1(n5997), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5991) );
  OR2_X1 U4904 ( .A1(n9389), .A2(n4477), .ZN(n4608) );
  AOI21_X1 U4905 ( .B1(n9239), .B2(n9821), .A(n9238), .ZN(n9398) );
  NAND2_X1 U4906 ( .A1(n7895), .A2(n7894), .ZN(n8935) );
  AND2_X1 U4907 ( .A1(n8093), .A2(n8092), .ZN(n8099) );
  OAI21_X1 U4908 ( .B1(n5681), .B2(n5680), .A(n8572), .ZN(n5706) );
  NOR3_X1 U4909 ( .A1(n8089), .A2(n8088), .A3(n8087), .ZN(n8093) );
  NAND2_X1 U4910 ( .A1(n4399), .A2(n4537), .ZN(n9026) );
  NAND2_X1 U4911 ( .A1(n4697), .A2(n4696), .ZN(n8728) );
  NAND2_X1 U4912 ( .A1(n8312), .A2(n8311), .ZN(n9390) );
  OR2_X1 U4913 ( .A1(n8887), .A2(n8732), .ZN(n7965) );
  NAND2_X1 U4914 ( .A1(n5054), .A2(n5053), .ZN(n8869) );
  NAND2_X1 U4915 ( .A1(n7937), .A2(n7936), .ZN(n9395) );
  NAND2_X1 U4916 ( .A1(n5466), .A2(n5465), .ZN(n8881) );
  OAI21_X1 U4917 ( .B1(n8571), .B2(n4842), .A(n4839), .ZN(n5657) );
  NAND2_X1 U4918 ( .A1(n5529), .A2(n8059), .ZN(n8774) );
  AND2_X1 U4919 ( .A1(n8275), .A2(n9210), .ZN(n9326) );
  AOI21_X1 U4920 ( .B1(n5656), .B2(n4841), .A(n4840), .ZN(n4839) );
  NAND2_X1 U4921 ( .A1(n7849), .A2(n7848), .ZN(n9416) );
  INV_X1 U4922 ( .A(n5656), .ZN(n4842) );
  NAND2_X1 U4923 ( .A1(n5436), .A2(n5435), .ZN(n7815) );
  OR2_X1 U4924 ( .A1(n8911), .A2(n8779), .ZN(n8063) );
  NAND2_X1 U4925 ( .A1(n5410), .A2(n5409), .ZN(n8905) );
  NAND2_X1 U4926 ( .A1(n7606), .A2(n5644), .ZN(n7672) );
  AOI21_X1 U4927 ( .B1(n7635), .B2(n7634), .A(n7633), .ZN(n9174) );
  NAND2_X1 U4928 ( .A1(n5402), .A2(n5401), .ZN(n8911) );
  OR2_X1 U4929 ( .A1(n9435), .A2(n9177), .ZN(n8356) );
  OR2_X1 U4930 ( .A1(n7605), .A2(n7604), .ZN(n7606) );
  XNOR2_X1 U4931 ( .A(n5424), .B(n5423), .ZN(n7778) );
  AOI21_X1 U4932 ( .B1(n7500), .B2(n8375), .A(n7499), .ZN(n7635) );
  NAND2_X1 U4933 ( .A1(n4745), .A2(n4412), .ZN(n5424) );
  OAI21_X1 U4934 ( .B1(n9729), .B2(n9735), .A(n8247), .ZN(n7276) );
  OR2_X1 U4935 ( .A1(n8852), .A2(n8576), .ZN(n8050) );
  AND2_X1 U4936 ( .A1(n7639), .A2(n7638), .ZN(n9173) );
  AND2_X1 U4937 ( .A1(n7716), .A2(n7715), .ZN(n8263) );
  NAND2_X1 U4938 ( .A1(n5525), .A2(n4594), .ZN(n10111) );
  NAND2_X1 U4939 ( .A1(n7330), .A2(n4550), .ZN(n4549) );
  OR2_X1 U4940 ( .A1(n5370), .A2(n5369), .ZN(n5385) );
  NAND2_X1 U4941 ( .A1(n6607), .A2(n4743), .ZN(n7072) );
  NAND2_X1 U4942 ( .A1(n5346), .A2(n5345), .ZN(n8544) );
  NAND2_X1 U4943 ( .A1(n7487), .A2(n7486), .ZN(n9449) );
  NAND2_X1 U4944 ( .A1(n5327), .A2(n5326), .ZN(n7679) );
  NAND2_X1 U4945 ( .A1(n5521), .A2(n7972), .ZN(n7077) );
  AND2_X1 U4946 ( .A1(n6777), .A2(n8229), .ZN(n8417) );
  AOI21_X1 U4947 ( .B1(n6799), .B2(n6798), .A(n4865), .ZN(n7172) );
  NAND2_X1 U4948 ( .A1(n5292), .A2(n5291), .ZN(n7407) );
  NAND2_X1 U4949 ( .A1(n7259), .A2(n7258), .ZN(n9918) );
  AND2_X1 U4950 ( .A1(n8422), .A2(n9745), .ZN(n8369) );
  OAI21_X1 U4951 ( .B1(n4620), .B2(n4619), .A(n6701), .ZN(n6799) );
  AOI22_X1 U4952 ( .A1(n6260), .A2(n6259), .B1(n6258), .B2(n6257), .ZN(n6442)
         );
  OR2_X1 U4953 ( .A1(n6523), .A2(n4562), .ZN(n4561) );
  AND2_X2 U4954 ( .A1(n5597), .A2(n10038), .ZN(n8797) );
  CLKBUF_X1 U4955 ( .A(n5226), .Z(n5245) );
  NOR2_X1 U4956 ( .A1(n5699), .A2(n5698), .ZN(n8580) );
  NAND2_X1 U4957 ( .A1(n6571), .A2(n6570), .ZN(n6642) );
  AND3_X1 U4958 ( .A1(n5166), .A2(n5165), .A3(n5164), .ZN(n6599) );
  OAI211_X2 U4960 ( .C1(n8173), .C2(n9620), .A(n6418), .B(n6417), .ZN(n6817)
         );
  NOR2_X1 U4961 ( .A1(n9978), .A2(n6406), .ZN(n9977) );
  AND3_X1 U4962 ( .A1(n5132), .A2(n5131), .A3(n5130), .ZN(n10070) );
  INV_X2 U4963 ( .A(n8500), .ZN(n6105) );
  AND3_X1 U4964 ( .A1(n6251), .A2(n6250), .A3(n6249), .ZN(n9849) );
  NAND2_X1 U4965 ( .A1(n6070), .A2(n6749), .ZN(n6166) );
  NAND4_X1 U4966 ( .A1(n6189), .A2(n6188), .A3(n6187), .A4(n6186), .ZN(n9080)
         );
  NAND4_X1 U4967 ( .A1(n6218), .A2(n6217), .A3(n6216), .A4(n6215), .ZN(n9079)
         );
  NAND2_X2 U4968 ( .A1(n6157), .A2(n6621), .ZN(n7948) );
  INV_X1 U4969 ( .A(n6130), .ZN(n4350) );
  CLKBUF_X1 U4970 ( .A(n7282), .Z(n7876) );
  AND3_X1 U4971 ( .A1(n5074), .A2(n5073), .A3(n5072), .ZN(n10054) );
  INV_X1 U4972 ( .A(n8496), .ZN(n7294) );
  NOR2_X1 U4973 ( .A1(n5339), .A2(P2_IR_REG_16__SCAN_IN), .ZN(n5343) );
  NAND2_X1 U4974 ( .A1(n5556), .A2(n5555), .ZN(n5572) );
  NAND2_X1 U4975 ( .A1(n5566), .A2(n5048), .ZN(n8496) );
  INV_X1 U4976 ( .A(n6003), .ZN(n7599) );
  NAND2_X1 U4977 ( .A1(n5324), .A2(n4872), .ZN(n5339) );
  XNOR2_X1 U4978 ( .A(n5558), .B(n5562), .ZN(n8497) );
  OR2_X1 U4979 ( .A1(n5551), .A2(n5563), .ZN(n5556) );
  XNOR2_X1 U4980 ( .A(n5047), .B(n5046), .ZN(n5538) );
  NAND2_X1 U4981 ( .A1(n5906), .A2(n4365), .ZN(n7306) );
  AND2_X1 U4982 ( .A1(n5557), .A2(n5554), .ZN(n5555) );
  XNOR2_X1 U4983 ( .A(n4916), .B(P2_IR_REG_29__SCAN_IN), .ZN(n7482) );
  NAND2_X1 U4984 ( .A1(n5050), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5047) );
  XNOR2_X1 U4985 ( .A(n5991), .B(n5995), .ZN(n9567) );
  MUX2_X1 U4986 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5049), .S(
        P2_IR_REG_27__SCAN_IN), .Z(n5051) );
  NOR2_X1 U4987 ( .A1(n6056), .A2(n5911), .ZN(n6061) );
  OR2_X1 U4988 ( .A1(n5997), .A2(n5996), .ZN(n7622) );
  AND4_X1 U4989 ( .A1(n4754), .A2(n4909), .A3(n5145), .A4(n4607), .ZN(n5045)
         );
  INV_X1 U4990 ( .A(n6200), .ZN(n5979) );
  NOR2_X1 U4991 ( .A1(n4389), .A2(n4755), .ZN(n4754) );
  NAND2_X1 U4992 ( .A1(n4926), .A2(n4925), .ZN(n4732) );
  NAND2_X1 U4993 ( .A1(n4928), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n4731) );
  NAND2_X1 U4994 ( .A1(n5974), .A2(n4611), .ZN(n4610) );
  NOR2_X1 U4995 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_4__SCAN_IN), .ZN(
        n5898) );
  NOR2_X2 U4996 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), .ZN(
        n5897) );
  INV_X2 U4997 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  INV_X4 U4998 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X1 U4999 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n4925) );
  NOR2_X1 U5000 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n4617) );
  NOR2_X1 U5001 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n4526) );
  NOR2_X1 U5002 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n4618) );
  NOR2_X1 U5003 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n4566) );
  INV_X1 U5004 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n6059) );
  NAND2_X2 U5005 ( .A1(n7482), .A2(n4918), .ZN(n5084) );
  INV_X4 U5006 ( .A(n5104), .ZN(n5540) );
  OAI22_X2 U5007 ( .A1(n5319), .A2(n4992), .B1(SI_16_), .B2(n5317), .ZN(n5337)
         );
  OR2_X4 U5008 ( .A1(n7601), .A2(n6003), .ZN(n7941) );
  NOR2_X2 U5009 ( .A1(n6443), .A2(n6444), .ZN(n6524) );
  OAI22_X2 U5010 ( .A1(n6442), .A2(n6441), .B1(n6440), .B2(n6439), .ZN(n6443)
         );
  AND3_X2 U5011 ( .A1(n6529), .A2(n6528), .A3(n6527), .ZN(n9861) );
  NOR2_X2 U5012 ( .A1(n7782), .A2(n7810), .ZN(n7800) );
  OR2_X2 U5013 ( .A1(n7766), .A2(n9032), .ZN(n7782) );
  XNOR2_X1 U5014 ( .A(n6060), .B(P1_IR_REG_19__SCAN_IN), .ZN(n6074) );
  XNOR2_X2 U5015 ( .A(n4612), .B(n5975), .ZN(n6484) );
  NOR2_X2 U5016 ( .A1(n7283), .A2(n9055), .ZN(n7436) );
  OR2_X2 U5017 ( .A1(n7263), .A2(n7262), .ZN(n7283) );
  XNOR2_X2 U5018 ( .A(n7943), .B(n7942), .ZN(n9244) );
  NOR2_X4 U5019 ( .A1(n5128), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n5145) );
  AND2_X1 U5020 ( .A1(n5420), .A2(n5423), .ZN(n5016) );
  INV_X1 U5021 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n5908) );
  INV_X1 U5022 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n4565) );
  NAND2_X1 U5023 ( .A1(n6749), .A2(n6151), .ZN(n6156) );
  NOR2_X1 U5024 ( .A1(n9252), .A2(n9395), .ZN(n9230) );
  OR2_X1 U5025 ( .A1(n9421), .A2(n9188), .ZN(n8379) );
  INV_X1 U5026 ( .A(SI_10_), .ZN(n4976) );
  INV_X1 U5027 ( .A(n8703), .ZN(n5873) );
  INV_X1 U5028 ( .A(n5120), .ZN(n5468) );
  OAI22_X1 U5029 ( .A1(n5219), .A2(n5066), .B1(n5084), .B2(n10121), .ZN(n4705)
         );
  AND2_X1 U5030 ( .A1(n6045), .A2(n5907), .ZN(n5924) );
  AOI21_X1 U5031 ( .B1(n8057), .B2(n8063), .A(n8085), .ZN(n4507) );
  NAND2_X1 U5032 ( .A1(n8058), .A2(n8063), .ZN(n4508) );
  NOR2_X1 U5033 ( .A1(n4588), .A2(n8118), .ZN(n4587) );
  INV_X1 U5034 ( .A(n4591), .ZN(n4588) );
  AND2_X1 U5035 ( .A1(n8668), .A2(n8169), .ZN(n5571) );
  NAND2_X1 U5036 ( .A1(n4961), .A2(n4960), .ZN(n4512) );
  NOR2_X2 U5037 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5896) );
  OAI21_X1 U5038 ( .B1(n4377), .B2(n4855), .A(n4856), .ZN(n4854) );
  OR2_X1 U5039 ( .A1(n7817), .A2(n8753), .ZN(n4856) );
  INV_X1 U5040 ( .A(n7482), .ZN(n4917) );
  NAND2_X1 U5041 ( .A1(n6356), .A2(n4460), .ZN(n5784) );
  OR2_X1 U5042 ( .A1(n6360), .A2(n5829), .ZN(n4460) );
  OR2_X1 U5043 ( .A1(n7679), .A2(n5335), .ZN(n8043) );
  INV_X1 U5044 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5560) );
  INV_X1 U5045 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5161) );
  INV_X1 U5046 ( .A(n4548), .ZN(n4546) );
  OR2_X1 U5047 ( .A1(n7549), .A2(n7548), .ZN(n7550) );
  INV_X1 U5048 ( .A(n4551), .ZN(n4550) );
  OAI21_X1 U5049 ( .B1(n4354), .B2(n7230), .A(n4552), .ZN(n4551) );
  INV_X1 U5050 ( .A(n7242), .ZN(n4552) );
  OR2_X1 U5051 ( .A1(n7871), .A2(n8970), .ZN(n7891) );
  AND2_X1 U5052 ( .A1(n7683), .A2(n4410), .ZN(n7684) );
  AND2_X1 U5053 ( .A1(n9380), .A2(n9163), .ZN(n8455) );
  NOR2_X1 U5054 ( .A1(n9643), .A2(n9642), .ZN(n9641) );
  OR2_X1 U5055 ( .A1(n9416), .A2(n9189), .ZN(n9213) );
  AOI21_X1 U5056 ( .B1(n4871), .B2(n9186), .A(n4396), .ZN(n4653) );
  INV_X1 U5057 ( .A(n6156), .ZN(n6621) );
  NAND2_X1 U5058 ( .A1(n7571), .A2(n7570), .ZN(n7617) );
  OR2_X1 U5059 ( .A1(n7569), .A2(n7568), .ZN(n7570) );
  AND2_X1 U5060 ( .A1(n5041), .A2(n5040), .ZN(n5056) );
  OR2_X1 U5061 ( .A1(n5039), .A2(n5038), .ZN(n5040) );
  NAND2_X1 U5062 ( .A1(n5669), .A2(n8474), .ZN(n5877) );
  NAND2_X1 U5063 ( .A1(n4875), .A2(n8668), .ZN(n4489) );
  NAND2_X1 U5064 ( .A1(n7482), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n4704) );
  NAND2_X1 U5065 ( .A1(n7314), .A2(n7315), .ZN(n7313) );
  XNOR2_X1 U5066 ( .A(n8689), .B(n8869), .ZN(n8482) );
  AOI21_X1 U5067 ( .B1(n4698), .B2(n4700), .A(n4395), .ZN(n4696) );
  NAND2_X1 U5068 ( .A1(n5418), .A2(n4698), .ZN(n4697) );
  OR2_X1 U5069 ( .A1(n8905), .A2(n7833), .ZN(n8068) );
  AOI21_X1 U5070 ( .B1(n4708), .B2(n4710), .A(n4419), .ZN(n4706) );
  OR2_X1 U5071 ( .A1(n8544), .A2(n7674), .ZN(n8802) );
  NOR2_X1 U5072 ( .A1(n4596), .A2(n7394), .ZN(n4595) );
  INV_X1 U5073 ( .A(n8039), .ZN(n4596) );
  AND2_X1 U5074 ( .A1(n5695), .A2(n8085), .ZN(n8807) );
  INV_X1 U5075 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n4914) );
  NAND2_X1 U5076 ( .A1(n7626), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4687) );
  NOR2_X2 U5077 ( .A1(n4908), .A2(n5253), .ZN(n4909) );
  NAND2_X1 U5078 ( .A1(n6155), .A2(n6152), .ZN(n6153) );
  NAND2_X1 U5079 ( .A1(n6166), .A2(n6156), .ZN(n6152) );
  AND2_X1 U5080 ( .A1(n7791), .A2(n7790), .ZN(n9188) );
  NAND2_X1 U5081 ( .A1(n9230), .A2(n9155), .ZN(n9231) );
  NAND2_X1 U5082 ( .A1(n4646), .A2(n4643), .ZN(n9278) );
  INV_X1 U5083 ( .A(n4644), .ZN(n4643) );
  OAI22_X1 U5084 ( .A1(n9191), .A2(n4645), .B1(n9190), .B2(n9416), .ZN(n4644)
         );
  NAND2_X1 U5085 ( .A1(n4809), .A2(n4359), .ZN(n4812) );
  NAND2_X1 U5086 ( .A1(n4641), .A2(n4388), .ZN(n9362) );
  NAND2_X1 U5087 ( .A1(n9174), .A2(n4870), .ZN(n4641) );
  NAND2_X1 U5088 ( .A1(n8173), .A2(n4962), .ZN(n7636) );
  NAND2_X1 U5089 ( .A1(n9812), .A2(n6617), .ZN(n6664) );
  OR2_X1 U5090 ( .A1(n6616), .A2(n6626), .ZN(n6617) );
  NAND2_X1 U5091 ( .A1(n9815), .A2(n9813), .ZN(n9812) );
  NOR2_X1 U5092 ( .A1(n4882), .A2(n5977), .ZN(n5978) );
  OR2_X1 U5093 ( .A1(n5976), .A2(P1_IR_REG_25__SCAN_IN), .ZN(n4882) );
  INV_X1 U5094 ( .A(n5977), .ZN(n5903) );
  NAND2_X1 U5095 ( .A1(n6062), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6063) );
  NAND2_X1 U5096 ( .A1(n4723), .A2(n4975), .ZN(n5212) );
  NAND2_X1 U5097 ( .A1(n4730), .A2(n4728), .ZN(n4723) );
  NAND2_X1 U5098 ( .A1(n5192), .A2(n4970), .ZN(n4730) );
  NAND2_X1 U5099 ( .A1(n4486), .A2(n4489), .ZN(n4484) );
  INV_X1 U5100 ( .A(n4487), .ZN(n4486) );
  AND2_X1 U5101 ( .A1(n8165), .A2(n7112), .ZN(n4449) );
  NAND2_X1 U5102 ( .A1(n5065), .A2(n5064), .ZN(n8703) );
  OAI21_X1 U5103 ( .B1(n8023), .B2(n8024), .A(n5265), .ZN(n4496) );
  INV_X1 U5104 ( .A(n8146), .ZN(n4497) );
  NAND2_X1 U5105 ( .A1(n4502), .A2(n4508), .ZN(n4501) );
  NOR2_X1 U5106 ( .A1(n4505), .A2(n4503), .ZN(n4502) );
  NAND2_X1 U5107 ( .A1(n4507), .A2(n4400), .ZN(n4503) );
  NAND2_X1 U5108 ( .A1(n5211), .A2(n4975), .ZN(n4726) );
  NOR2_X1 U5109 ( .A1(n4726), .A2(n4722), .ZN(n4721) );
  INV_X1 U5110 ( .A(n4970), .ZN(n4722) );
  OR2_X1 U5111 ( .A1(n5714), .A2(n8487), .ZN(n8123) );
  AND3_X1 U5112 ( .A1(n6596), .A2(n8006), .A3(n7991), .ZN(n4570) );
  INV_X1 U5113 ( .A(n8002), .ZN(n4572) );
  NOR2_X1 U5114 ( .A1(n4820), .A2(n9265), .ZN(n4814) );
  AND2_X1 U5115 ( .A1(n5487), .A2(n5486), .ZN(n7569) );
  OR2_X1 U5116 ( .A1(n5022), .A2(n5447), .ZN(n5035) );
  NOR2_X1 U5117 ( .A1(P1_IR_REG_23__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), .ZN(
        n5915) );
  AND2_X1 U5118 ( .A1(n8117), .A2(n4586), .ZN(n4585) );
  NAND2_X1 U5119 ( .A1(n9963), .A2(n9962), .ZN(n9961) );
  NAND2_X1 U5120 ( .A1(n9961), .A2(n4459), .ZN(n4458) );
  OR2_X1 U5121 ( .A1(n9965), .A2(n5775), .ZN(n4459) );
  NOR2_X1 U5122 ( .A1(n6313), .A2(n4776), .ZN(n5752) );
  NOR2_X1 U5123 ( .A1(n6323), .A2(n6610), .ZN(n4776) );
  NAND2_X1 U5124 ( .A1(n6737), .A2(n5786), .ZN(n5787) );
  NOR2_X1 U5125 ( .A1(n5467), .A2(n4897), .ZN(n4444) );
  NAND2_X1 U5126 ( .A1(n4480), .A2(n4479), .ZN(n7973) );
  INV_X1 U5127 ( .A(n4699), .ZN(n4698) );
  OAI21_X1 U5128 ( .B1(n8131), .B2(n4700), .A(n5432), .ZN(n4699) );
  OR2_X1 U5129 ( .A1(n7815), .A2(n8714), .ZN(n8130) );
  NAND2_X1 U5130 ( .A1(n4719), .A2(n4371), .ZN(n4718) );
  INV_X1 U5131 ( .A(n8790), .ZN(n4719) );
  OR2_X1 U5132 ( .A1(n8917), .A2(n8794), .ZN(n8060) );
  AND2_X1 U5133 ( .A1(n8132), .A2(n4577), .ZN(n4576) );
  NAND2_X1 U5134 ( .A1(n8049), .A2(n4578), .ZN(n4577) );
  INV_X1 U5135 ( .A(n8043), .ZN(n4578) );
  OR2_X1 U5136 ( .A1(n7603), .A2(n7584), .ZN(n8040) );
  AND2_X1 U5137 ( .A1(n5560), .A2(n5589), .ZN(n5552) );
  INV_X1 U5138 ( .A(n5320), .ZN(n5324) );
  NAND2_X1 U5139 ( .A1(n4543), .A2(n7775), .ZN(n4538) );
  AND2_X1 U5140 ( .A1(n4540), .A2(n7761), .ZN(n4539) );
  NAND2_X1 U5141 ( .A1(n7758), .A2(n7760), .ZN(n7761) );
  OR2_X1 U5142 ( .A1(n4541), .A2(n7739), .ZN(n4540) );
  INV_X1 U5143 ( .A(n7759), .ZN(n7760) );
  INV_X1 U5144 ( .A(n7757), .ZN(n4541) );
  INV_X1 U5145 ( .A(n6158), .ZN(n7924) );
  NOR2_X1 U5146 ( .A1(n9641), .A2(n4413), .ZN(n9494) );
  OR2_X1 U5147 ( .A1(n9494), .A2(n9495), .ZN(n4679) );
  NOR2_X1 U5148 ( .A1(n9481), .A2(n4682), .ZN(n9658) );
  AND2_X1 U5149 ( .A1(n9489), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n4682) );
  AOI21_X1 U5150 ( .B1(P1_REG2_REG_10__SCAN_IN), .B2(n9489), .A(n9484), .ZN(
        n9662) );
  OR2_X1 U5151 ( .A1(n9658), .A2(n9659), .ZN(n4681) );
  NOR2_X1 U5152 ( .A1(n9684), .A2(n4683), .ZN(n9101) );
  NOR2_X1 U5153 ( .A1(n9694), .A2(n7260), .ZN(n4683) );
  AOI21_X1 U5154 ( .B1(n4675), .B2(n4674), .A(n4673), .ZN(n4672) );
  INV_X1 U5155 ( .A(n9138), .ZN(n4673) );
  INV_X1 U5156 ( .A(n9135), .ZN(n4674) );
  NAND2_X1 U5157 ( .A1(n4672), .A2(n4670), .ZN(n4669) );
  NAND2_X1 U5158 ( .A1(n4676), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n4670) );
  INV_X1 U5159 ( .A(n9216), .ZN(n4823) );
  NOR2_X1 U5160 ( .A1(n9304), .A2(n9214), .ZN(n4827) );
  AND2_X1 U5161 ( .A1(n9213), .A2(n8334), .ZN(n9212) );
  OR2_X1 U5162 ( .A1(n8183), .A2(n9181), .ZN(n8355) );
  OR2_X1 U5163 ( .A1(n8184), .A2(n9176), .ZN(n8328) );
  INV_X1 U5164 ( .A(n9068), .ZN(n7362) );
  AND2_X1 U5165 ( .A1(n8252), .A2(n7269), .ZN(n8373) );
  OR2_X1 U5166 ( .A1(n9734), .A2(n7362), .ZN(n8247) );
  NAND2_X1 U5167 ( .A1(n9906), .A2(n7363), .ZN(n4661) );
  OR2_X1 U5168 ( .A1(n7173), .A2(n9070), .ZN(n8235) );
  NAND2_X1 U5169 ( .A1(n9873), .A2(n6758), .ZN(n8228) );
  XNOR2_X1 U5170 ( .A(n7569), .B(n7567), .ZN(n7566) );
  NAND2_X1 U5171 ( .A1(n5056), .A2(n5055), .ZN(n5482) );
  NOR2_X1 U5172 ( .A1(n5916), .A2(n5973), .ZN(n5917) );
  INV_X1 U5173 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5916) );
  NAND2_X1 U5174 ( .A1(n4746), .A2(n4863), .ZN(n5421) );
  INV_X1 U5175 ( .A(n5286), .ZN(n4988) );
  OR2_X1 U5176 ( .A1(n6090), .A2(P1_IR_REG_11__SCAN_IN), .ZN(n6091) );
  NOR2_X1 U5177 ( .A1(n5191), .A2(n4514), .ZN(n4513) );
  INV_X1 U5178 ( .A(n4965), .ZN(n4514) );
  NAND2_X1 U5179 ( .A1(n4511), .A2(n4518), .ZN(n4515) );
  AND2_X1 U5180 ( .A1(n4512), .A2(n4963), .ZN(n4518) );
  OR2_X1 U5181 ( .A1(n5945), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n5959) );
  INV_X1 U5182 ( .A(SI_1_), .ZN(n4695) );
  AND2_X1 U5183 ( .A1(n5876), .A2(n5875), .ZN(n8473) );
  INV_X1 U5184 ( .A(n4849), .ZN(n4848) );
  OAI21_X1 U5185 ( .B1(n4850), .B2(n7537), .A(n7536), .ZN(n4849) );
  NAND2_X1 U5186 ( .A1(n5664), .A2(n5663), .ZN(n8472) );
  OAI21_X1 U5187 ( .B1(n8513), .B2(n4855), .A(n4853), .ZN(n5664) );
  INV_X1 U5188 ( .A(n4854), .ZN(n4853) );
  OR2_X1 U5189 ( .A1(n5631), .A2(n5630), .ZN(n5632) );
  NAND2_X1 U5190 ( .A1(n5658), .A2(n8779), .ZN(n5659) );
  AND4_X1 U5191 ( .A1(n5333), .A2(n5332), .A3(n5331), .A4(n5330), .ZN(n5335)
         );
  NAND2_X1 U5192 ( .A1(n4357), .A2(n7576), .ZN(n4580) );
  XNOR2_X1 U5193 ( .A(n4458), .B(n6302), .ZN(n6294) );
  OR2_X1 U5194 ( .A1(n5741), .A2(n5932), .ZN(n5742) );
  NAND2_X1 U5195 ( .A1(n6357), .A2(n6358), .ZN(n6356) );
  NOR2_X1 U5196 ( .A1(n6350), .A2(n7058), .ZN(n4778) );
  XNOR2_X1 U5197 ( .A(n5784), .B(n7058), .ZN(n7056) );
  NAND2_X1 U5198 ( .A1(n6738), .A2(n6739), .ZN(n6737) );
  NAND2_X1 U5199 ( .A1(n4782), .A2(n4781), .ZN(n6348) );
  AND2_X1 U5200 ( .A1(n4779), .A2(n4784), .ZN(n7061) );
  AOI21_X1 U5201 ( .B1(n6351), .B2(n4787), .A(n4780), .ZN(n4779) );
  OAI21_X1 U5202 ( .B1(n4788), .B2(n4781), .A(n4783), .ZN(n4780) );
  AND2_X1 U5203 ( .A1(n4789), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n4783) );
  XNOR2_X1 U5204 ( .A(n5787), .B(n5839), .ZN(n7184) );
  NAND2_X1 U5205 ( .A1(n7313), .A2(n5789), .ZN(n5790) );
  INV_X1 U5206 ( .A(n4796), .ZN(n4793) );
  NOR2_X1 U5207 ( .A1(n8639), .A2(n5766), .ZN(n5767) );
  NAND2_X1 U5208 ( .A1(n4444), .A2(n6972), .ZN(n5598) );
  INV_X1 U5209 ( .A(n4444), .ZN(n5059) );
  OR2_X1 U5210 ( .A1(n4374), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n5437) );
  INV_X1 U5211 ( .A(n8593), .ZN(n7525) );
  NAND2_X1 U5212 ( .A1(n6693), .A2(n8102), .ZN(n4481) );
  INV_X1 U5213 ( .A(n8594), .ZN(n7477) );
  AND2_X1 U5214 ( .A1(n5208), .A2(n5197), .ZN(n4743) );
  AND2_X1 U5215 ( .A1(n7973), .A2(n7967), .ZN(n8143) );
  INV_X1 U5216 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n4885) );
  NOR2_X1 U5217 ( .A1(n10086), .A2(n7979), .ZN(n5709) );
  NAND2_X1 U5218 ( .A1(n4736), .A2(n4740), .ZN(n8688) );
  NAND2_X1 U5219 ( .A1(n8711), .A2(n4741), .ZN(n4736) );
  NAND2_X1 U5220 ( .A1(n8689), .A2(n8809), .ZN(n8691) );
  AND2_X1 U5221 ( .A1(n4400), .A2(n8068), .ZN(n4603) );
  NAND2_X1 U5222 ( .A1(n8747), .A2(n8069), .ZN(n4604) );
  NAND2_X1 U5223 ( .A1(n5418), .A2(n8131), .ZN(n8752) );
  NAND2_X1 U5224 ( .A1(n8765), .A2(n4371), .ZN(n4713) );
  INV_X1 U5225 ( .A(n4712), .ZN(n4711) );
  OAI21_X1 U5226 ( .B1(n4716), .B2(n4717), .A(n8762), .ZN(n4712) );
  INV_X1 U5227 ( .A(n5092), .ZN(n5357) );
  AND4_X1 U5228 ( .A1(n5352), .A2(n5351), .A3(n5350), .A4(n5349), .ZN(n7674)
         );
  NAND2_X1 U5229 ( .A1(n7509), .A2(n5334), .ZN(n7579) );
  NAND2_X1 U5230 ( .A1(n5697), .A2(n8085), .ZN(n10041) );
  AND2_X1 U5231 ( .A1(n8040), .A2(n8039), .ZN(n8149) );
  NOR2_X1 U5232 ( .A1(n8035), .A2(n4599), .ZN(n4598) );
  INV_X1 U5233 ( .A(n8031), .ZN(n4599) );
  INV_X1 U5234 ( .A(n10041), .ZN(n8809) );
  OR2_X1 U5235 ( .A1(n5535), .A2(n5603), .ZN(n6275) );
  NAND2_X1 U5236 ( .A1(n7070), .A2(n7101), .ZN(n10103) );
  INV_X1 U5237 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5589) );
  INV_X1 U5238 ( .A(n4902), .ZN(n4755) );
  INV_X1 U5239 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5228) );
  XNOR2_X1 U5240 ( .A(n5214), .B(P2_IR_REG_10__SCAN_IN), .ZN(n6360) );
  AND2_X1 U5241 ( .A1(n5179), .A2(n5205), .ZN(n10019) );
  AND2_X1 U5242 ( .A1(n4899), .A2(n4900), .ZN(n4852) );
  INV_X1 U5243 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n4900) );
  NAND2_X1 U5244 ( .A1(n4462), .A2(n4461), .ZN(n5095) );
  INV_X1 U5245 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n4462) );
  INV_X1 U5246 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n4461) );
  INV_X1 U5247 ( .A(n4555), .ZN(n4547) );
  AOI21_X1 U5248 ( .B1(n4546), .B2(n4555), .A(n4554), .ZN(n4545) );
  AND2_X1 U5249 ( .A1(n7357), .A2(n4556), .ZN(n4555) );
  INV_X1 U5250 ( .A(n9078), .ZN(n6639) );
  NAND2_X1 U5251 ( .A1(n8935), .A2(n4390), .ZN(n8939) );
  NAND2_X1 U5252 ( .A1(n4544), .A2(n4543), .ZN(n4542) );
  INV_X1 U5253 ( .A(n6524), .ZN(n4559) );
  NOR2_X1 U5254 ( .A1(n6523), .A2(n4564), .ZN(n4558) );
  NAND2_X1 U5255 ( .A1(n6695), .A2(n6694), .ZN(n7338) );
  NAND2_X1 U5256 ( .A1(n6252), .A2(n6614), .ZN(n6207) );
  NAND2_X1 U5257 ( .A1(n7872), .A2(n7891), .ZN(n8971) );
  AND2_X1 U5258 ( .A1(n7866), .A2(n7865), .ZN(n9193) );
  AOI21_X1 U5259 ( .B1(n9294), .B2(n7876), .A(n7807), .ZN(n9189) );
  AND3_X1 U5260 ( .A1(n7735), .A2(n7734), .A3(n7733), .ZN(n9177) );
  MUX2_X1 U5261 ( .A(n6489), .B(P1_REG1_REG_1__SCAN_IN), .S(n6491), .Z(n9577)
         );
  NOR2_X1 U5262 ( .A1(n9581), .A2(n9580), .ZN(n9579) );
  OR2_X1 U5263 ( .A1(n9595), .A2(n9594), .ZN(n4432) );
  NOR2_X1 U5264 ( .A1(n9614), .A2(n4411), .ZN(n9626) );
  NOR2_X1 U5265 ( .A1(n9626), .A2(n9627), .ZN(n9625) );
  NOR2_X1 U5266 ( .A1(n9523), .A2(n4433), .ZN(n9083) );
  AND2_X1 U5267 ( .A1(n6653), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n4433) );
  NAND2_X1 U5268 ( .A1(n9083), .A2(n9084), .ZN(n9082) );
  XNOR2_X1 U5269 ( .A(n9101), .B(n9115), .ZN(n9701) );
  NOR2_X1 U5270 ( .A1(n9701), .A2(n7279), .ZN(n9700) );
  XNOR2_X1 U5271 ( .A(n9114), .B(n9115), .ZN(n9705) );
  NOR2_X1 U5272 ( .A1(n9688), .A2(n4435), .ZN(n9114) );
  AND2_X1 U5273 ( .A1(n9113), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n4435) );
  NOR2_X1 U5274 ( .A1(n9705), .A2(n9704), .ZN(n9703) );
  NAND2_X1 U5275 ( .A1(n8321), .A2(n8320), .ZN(n9156) );
  NAND2_X1 U5276 ( .A1(n4637), .A2(n9195), .ZN(n4636) );
  NOR2_X1 U5277 ( .A1(n9297), .A2(n8278), .ZN(n4828) );
  AOI21_X1 U5278 ( .B1(n4653), .B2(n4650), .A(n4394), .ZN(n4649) );
  INV_X1 U5279 ( .A(n4871), .ZN(n4650) );
  INV_X1 U5280 ( .A(n4653), .ZN(n4651) );
  INV_X1 U5281 ( .A(n9212), .ZN(n9297) );
  NAND2_X1 U5282 ( .A1(n9310), .A2(n9311), .ZN(n9309) );
  OR2_X1 U5283 ( .A1(n9185), .A2(n9323), .ZN(n4871) );
  NAND2_X1 U5284 ( .A1(n8256), .A2(n8251), .ZN(n4830) );
  AND2_X1 U5285 ( .A1(n9454), .A2(n9065), .ZN(n7499) );
  NAND2_X1 U5286 ( .A1(n4831), .A2(n8251), .ZN(n4833) );
  INV_X1 U5287 ( .A(n9547), .ZN(n4831) );
  INV_X1 U5288 ( .A(n8373), .ZN(n7277) );
  NAND2_X1 U5289 ( .A1(n7162), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n7263) );
  OAI21_X1 U5290 ( .B1(n7253), .B2(n8372), .A(n4661), .ZN(n9736) );
  AOI22_X1 U5291 ( .A1(n9742), .A2(n9741), .B1(n9070), .B2(n9898), .ZN(n7253)
         );
  AND2_X1 U5292 ( .A1(n8235), .A2(n8236), .ZN(n9744) );
  INV_X1 U5293 ( .A(n4623), .ZN(n4619) );
  NAND2_X1 U5294 ( .A1(n9789), .A2(n9790), .ZN(n6839) );
  AND2_X1 U5295 ( .A1(n8412), .A2(n8420), .ZN(n9781) );
  NAND2_X1 U5296 ( .A1(n4476), .A2(n9844), .ZN(n9805) );
  INV_X1 U5297 ( .A(n9828), .ZN(n4476) );
  INV_X1 U5298 ( .A(n9821), .ZN(n9746) );
  INV_X1 U5299 ( .A(n9227), .ZN(n9228) );
  NAND2_X1 U5300 ( .A1(n7781), .A2(n7780), .ZN(n9421) );
  INV_X1 U5301 ( .A(n9173), .ZN(n9445) );
  AND2_X1 U5302 ( .A1(n6549), .A2(n6166), .ZN(n9919) );
  NAND2_X1 U5303 ( .A1(n6071), .A2(n8175), .ZN(n9821) );
  AND2_X1 U5304 ( .A1(n9382), .A2(n6065), .ZN(n6545) );
  OAI211_X1 U5305 ( .C1(n6042), .C2(n6044), .A(n6045), .B(n6043), .ZN(n9475)
         );
  INV_X1 U5306 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n5992) );
  INV_X1 U5307 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5995) );
  INV_X1 U5308 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5975) );
  XNOR2_X1 U5309 ( .A(n5389), .B(n5388), .ZN(n7723) );
  NAND2_X1 U5310 ( .A1(n5385), .A2(n5384), .ZN(n5389) );
  NAND2_X1 U5311 ( .A1(n4996), .A2(n4742), .ZN(n5356) );
  AND2_X1 U5312 ( .A1(n4998), .A2(n4995), .ZN(n4742) );
  INV_X1 U5313 ( .A(n5354), .ZN(n4998) );
  NOR2_X1 U5314 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n4805) );
  INV_X1 U5315 ( .A(n4615), .ZN(n4613) );
  XNOR2_X1 U5316 ( .A(n5252), .B(n5251), .ZN(n7149) );
  XNOR2_X1 U5317 ( .A(n4665), .B(P1_IR_REG_1__SCAN_IN), .ZN(n6491) );
  NAND2_X1 U5318 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n4665) );
  NAND2_X1 U5319 ( .A1(n5877), .A2(n5875), .ZN(n4838) );
  AND4_X1 U5320 ( .A1(n5417), .A2(n5416), .A3(n5415), .A4(n5414), .ZN(n7833)
         );
  INV_X1 U5321 ( .A(n7216), .ZN(n7389) );
  OR2_X1 U5322 ( .A1(n4875), .A2(n8668), .ZN(n4488) );
  XNOR2_X1 U5323 ( .A(n5507), .B(P2_IR_REG_22__SCAN_IN), .ZN(n8169) );
  INV_X1 U5324 ( .A(n8732), .ZN(n8702) );
  OAI211_X1 U5325 ( .C1(n8107), .C2(n5441), .A(n5440), .B(n5439), .ZN(n8741)
         );
  INV_X1 U5326 ( .A(n7833), .ZN(n8768) );
  INV_X1 U5327 ( .A(n4703), .ZN(n4701) );
  OAI22_X1 U5328 ( .A1(n5104), .A2(n5067), .B1(n4918), .B2(n4704), .ZN(n4703)
         );
  OR2_X1 U5329 ( .A1(n7182), .A2(n5280), .ZN(n4766) );
  XNOR2_X1 U5330 ( .A(n5790), .B(n5800), .ZN(n8606) );
  NAND2_X1 U5331 ( .A1(n8624), .A2(n8625), .ZN(n8623) );
  NOR2_X1 U5332 ( .A1(n8640), .A2(n7662), .ZN(n8639) );
  NAND2_X1 U5333 ( .A1(n5767), .A2(n5768), .ZN(n5769) );
  OAI211_X1 U5334 ( .C1(n8660), .C2(n5864), .A(n5863), .B(n5862), .ZN(n5865)
         );
  NAND2_X1 U5335 ( .A1(n5549), .A2(n4880), .ZN(n5708) );
  NOR2_X1 U5336 ( .A1(n8030), .A2(n8020), .ZN(n4594) );
  NAND2_X1 U5337 ( .A1(n4593), .A2(n8083), .ZN(n5891) );
  NAND2_X1 U5338 ( .A1(n5887), .A2(n5886), .ZN(n5888) );
  NAND2_X1 U5339 ( .A1(n8703), .A2(n8807), .ZN(n5886) );
  NAND2_X1 U5340 ( .A1(n5058), .A2(n5057), .ZN(n8875) );
  NAND2_X1 U5341 ( .A1(n10118), .A2(n10112), .ZN(n8892) );
  XNOR2_X1 U5342 ( .A(n5512), .B(n4860), .ZN(n8115) );
  XOR2_X1 U5343 ( .A(n7952), .B(n7951), .Z(n7953) );
  OAI22_X1 U5344 ( .A1(n7941), .A2(n6084), .B1(n6262), .B2(n6083), .ZN(n6085)
         );
  INV_X1 U5345 ( .A(n9151), .ZN(n9152) );
  OAI21_X1 U5346 ( .B1(n9150), .B2(n9699), .A(n9724), .ZN(n9151) );
  AND2_X1 U5347 ( .A1(n6483), .A2(n5981), .ZN(n9609) );
  NAND2_X1 U5348 ( .A1(n8174), .A2(n8173), .ZN(n9380) );
  OAI21_X1 U5349 ( .B1(n4631), .B2(n4629), .A(n4626), .ZN(n9201) );
  AOI21_X1 U5350 ( .B1(n4628), .B2(n4627), .A(n4393), .ZN(n4626) );
  AND2_X1 U5351 ( .A1(n9232), .A2(n9231), .ZN(n9389) );
  OR2_X1 U5352 ( .A1(n6171), .A2(n6170), .ZN(n9799) );
  NAND2_X1 U5353 ( .A1(n6775), .A2(n6774), .ZN(n7299) );
  AND2_X1 U5354 ( .A1(n7999), .A2(n7968), .ZN(n8010) );
  INV_X1 U5355 ( .A(n4496), .ZN(n4495) );
  NAND2_X1 U5356 ( .A1(n4492), .A2(n4497), .ZN(n4490) );
  INV_X1 U5357 ( .A(n4504), .ZN(n4500) );
  NAND2_X1 U5358 ( .A1(n4509), .A2(n4510), .ZN(n4506) );
  NAND2_X1 U5359 ( .A1(n4508), .A2(n4507), .ZN(n4510) );
  NAND2_X1 U5360 ( .A1(n8289), .A2(n8288), .ZN(n8308) );
  AOI21_X1 U5361 ( .B1(n4524), .B2(n8085), .A(n4522), .ZN(n4521) );
  OR2_X1 U5362 ( .A1(n8701), .A2(n4523), .ZN(n4522) );
  NAND2_X1 U5363 ( .A1(n8073), .A2(n8072), .ZN(n4524) );
  AND2_X1 U5364 ( .A1(n8074), .A2(n8098), .ZN(n4523) );
  NAND2_X1 U5365 ( .A1(n4520), .A2(n4590), .ZN(n4519) );
  INV_X1 U5366 ( .A(n8082), .ZN(n4520) );
  NAND2_X1 U5367 ( .A1(n4587), .A2(n4589), .ZN(n4586) );
  AOI21_X1 U5368 ( .B1(n8482), .B2(n4592), .A(n4360), .ZN(n4591) );
  NAND2_X1 U5369 ( .A1(n4590), .A2(n8482), .ZN(n4589) );
  INV_X1 U5370 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5322) );
  INV_X1 U5371 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5273) );
  AND2_X1 U5372 ( .A1(n4409), .A2(n7704), .ZN(n4527) );
  OR2_X1 U5373 ( .A1(n8990), .A2(n7705), .ZN(n7704) );
  AND2_X1 U5374 ( .A1(n5030), .A2(n5032), .ZN(n5031) );
  OR2_X1 U5375 ( .A1(n5037), .A2(n5036), .ZN(n5038) );
  INV_X1 U5376 ( .A(n4725), .ZN(n4724) );
  OAI21_X1 U5377 ( .B1(n4728), .B2(n4726), .A(n4978), .ZN(n4725) );
  INV_X1 U5378 ( .A(n7816), .ZN(n4855) );
  NOR2_X1 U5379 ( .A1(n8505), .A2(n4844), .ZN(n4843) );
  INV_X1 U5380 ( .A(n5652), .ZN(n4844) );
  AND2_X1 U5381 ( .A1(n7524), .A2(n5625), .ZN(n5626) );
  INV_X1 U5382 ( .A(n4843), .ZN(n4841) );
  INV_X1 U5383 ( .A(n5611), .ZN(n5628) );
  NAND2_X1 U5384 ( .A1(n8472), .A2(n8521), .ZN(n5669) );
  AND2_X1 U5385 ( .A1(n6330), .A2(n4760), .ZN(n4759) );
  INV_X1 U5386 ( .A(n8657), .ZN(n4801) );
  INV_X1 U5387 ( .A(n8663), .ZN(n4799) );
  NOR2_X1 U5388 ( .A1(n5392), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n4447) );
  NOR2_X1 U5389 ( .A1(n5328), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n4446) );
  NOR2_X1 U5390 ( .A1(n5235), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n4448) );
  INV_X1 U5391 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n6740) );
  NAND2_X1 U5392 ( .A1(n5516), .A2(n7981), .ZN(n6510) );
  NAND2_X1 U5393 ( .A1(n8123), .A2(n8121), .ZN(n8087) );
  OAI21_X1 U5394 ( .B1(n8709), .B2(n4735), .A(n4737), .ZN(n5884) );
  NAND2_X1 U5395 ( .A1(n4740), .A2(n8156), .ZN(n4735) );
  INV_X1 U5396 ( .A(n4738), .ZN(n4737) );
  OAI21_X1 U5397 ( .B1(n4741), .B2(n4739), .A(n5474), .ZN(n4738) );
  AND2_X1 U5398 ( .A1(n4358), .A2(n5458), .ZN(n4741) );
  NAND2_X1 U5399 ( .A1(n4603), .A2(n4601), .ZN(n4600) );
  INV_X1 U5400 ( .A(n8069), .ZN(n4601) );
  INV_X1 U5401 ( .A(n5419), .ZN(n4700) );
  NOR2_X1 U5402 ( .A1(n8775), .A2(n4714), .ZN(n4717) );
  INV_X1 U5403 ( .A(n5383), .ZN(n4714) );
  INV_X1 U5404 ( .A(n4709), .ZN(n4708) );
  OAI21_X1 U5405 ( .B1(n5334), .B2(n4710), .A(n7656), .ZN(n4709) );
  INV_X1 U5406 ( .A(n5336), .ZN(n4710) );
  NAND2_X1 U5407 ( .A1(n6391), .A2(n4570), .ZN(n4569) );
  INV_X1 U5408 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n4901) );
  INV_X1 U5409 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5323) );
  OR2_X1 U5410 ( .A1(n5205), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n5213) );
  INV_X1 U5411 ( .A(n7551), .ZN(n4556) );
  OR2_X1 U5412 ( .A1(n9380), .A2(n8342), .ZN(n4689) );
  NOR2_X1 U5413 ( .A1(n9589), .A2(n4376), .ZN(n9509) );
  NOR2_X1 U5414 ( .A1(n9509), .A2(n9510), .ZN(n9508) );
  OR2_X1 U5415 ( .A1(n9513), .A2(n9514), .ZN(n4430) );
  NAND2_X1 U5416 ( .A1(n6649), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n4678) );
  NAND2_X1 U5417 ( .A1(n4675), .A2(n9139), .ZN(n4671) );
  INV_X1 U5418 ( .A(n9197), .ZN(n4634) );
  AND2_X1 U5419 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(n7903), .ZN(n7957) );
  INV_X1 U5420 ( .A(n9062), .ZN(n8313) );
  OR2_X1 U5421 ( .A1(n7857), .A2(n8976), .ZN(n7875) );
  OR2_X1 U5422 ( .A1(n9411), .A2(n9193), .ZN(n8383) );
  NAND2_X1 U5423 ( .A1(n4649), .A2(n4651), .ZN(n4645) );
  NOR2_X1 U5424 ( .A1(n9191), .A2(n4648), .ZN(n4647) );
  INV_X1 U5425 ( .A(n4649), .ZN(n4648) );
  NOR2_X1 U5426 ( .A1(n4467), .A2(n8183), .ZN(n4466) );
  INV_X1 U5427 ( .A(n4468), .ZN(n4467) );
  NOR2_X1 U5428 ( .A1(n4811), .A2(n8325), .ZN(n4810) );
  INV_X1 U5429 ( .A(n9371), .ZN(n4811) );
  NOR2_X1 U5430 ( .A1(n9435), .A2(n8184), .ZN(n4468) );
  NOR2_X1 U5431 ( .A1(n4353), .A2(n4660), .ZN(n4659) );
  INV_X1 U5432 ( .A(n9735), .ZN(n4660) );
  INV_X1 U5433 ( .A(n4661), .ZN(n4656) );
  NOR2_X1 U5434 ( .A1(n9918), .A2(n9734), .ZN(n4474) );
  INV_X1 U5435 ( .A(n6702), .ZN(n4621) );
  OR2_X1 U5436 ( .A1(n7338), .A2(n7223), .ZN(n8233) );
  NOR2_X1 U5437 ( .A1(n6642), .A2(n8210), .ZN(n4471) );
  NAND2_X1 U5438 ( .A1(n6614), .A2(n6267), .ZN(n8197) );
  OR2_X2 U5439 ( .A1(n6075), .A2(n4349), .ZN(n6155) );
  AND2_X1 U5440 ( .A1(n8353), .A2(n6166), .ZN(n6163) );
  AOI21_X1 U5441 ( .B1(n4819), .B2(n4816), .A(n8339), .ZN(n4815) );
  NAND2_X1 U5442 ( .A1(n9257), .A2(n9198), .ZN(n4635) );
  NAND2_X1 U5443 ( .A1(n9217), .A2(n4633), .ZN(n4632) );
  INV_X1 U5444 ( .A(n4636), .ZN(n4633) );
  NOR2_X1 U5445 ( .A1(n9755), .A2(n7173), .ZN(n9756) );
  OR2_X1 U5446 ( .A1(n6801), .A2(n7299), .ZN(n9755) );
  INV_X1 U5447 ( .A(SI_23_), .ZN(n5018) );
  INV_X1 U5448 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5912) );
  INV_X1 U5449 ( .A(SI_20_), .ZN(n5386) );
  INV_X1 U5450 ( .A(SI_17_), .ZN(n6966) );
  NOR2_X1 U5451 ( .A1(n5302), .A2(SI_15_), .ZN(n4758) );
  OR2_X1 U5452 ( .A1(n4757), .A2(n5301), .ZN(n4756) );
  INV_X1 U5453 ( .A(n5302), .ZN(n4757) );
  AND2_X1 U5454 ( .A1(n4729), .A2(n4879), .ZN(n4728) );
  NAND2_X1 U5455 ( .A1(n5191), .A2(n4970), .ZN(n4729) );
  AND2_X1 U5456 ( .A1(n5897), .A2(n5896), .ZN(n5938) );
  NAND2_X1 U5457 ( .A1(n5052), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n4733) );
  OAI21_X1 U5458 ( .B1(n4962), .B2(n4945), .A(n4944), .ZN(n4946) );
  XNOR2_X1 U5459 ( .A(n4940), .B(SI_2_), .ZN(n5091) );
  NAND2_X1 U5460 ( .A1(n4927), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n4928) );
  INV_X1 U5461 ( .A(SI_24_), .ZN(n6907) );
  INV_X1 U5462 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n8539) );
  INV_X1 U5463 ( .A(SI_22_), .ZN(n6886) );
  INV_X1 U5464 ( .A(SI_12_), .ZN(n6898) );
  INV_X1 U5465 ( .A(SI_27_), .ZN(n6918) );
  INV_X1 U5466 ( .A(SI_16_), .ZN(n6964) );
  INV_X1 U5467 ( .A(SI_14_), .ZN(n6959) );
  INV_X1 U5468 ( .A(SI_26_), .ZN(n6973) );
  INV_X1 U5469 ( .A(SI_25_), .ZN(n6940) );
  INV_X1 U5470 ( .A(SI_19_), .ZN(n6936) );
  NAND2_X1 U5471 ( .A1(n6823), .A2(n6822), .ZN(n6821) );
  AND2_X1 U5472 ( .A1(n5670), .A2(n5667), .ZN(n8522) );
  INV_X1 U5473 ( .A(n8712), .ZN(n8529) );
  NAND2_X1 U5474 ( .A1(n5648), .A2(n4858), .ZN(n8536) );
  NOR2_X1 U5475 ( .A1(n8538), .A2(n4859), .ZN(n4858) );
  INV_X1 U5476 ( .A(n5647), .ZN(n4859) );
  NAND2_X1 U5477 ( .A1(n4890), .A2(n4889), .ZN(n5217) );
  INV_X1 U5478 ( .A(n5198), .ZN(n4890) );
  NAND2_X1 U5479 ( .A1(n8571), .A2(n4843), .ZN(n8503) );
  AND2_X1 U5480 ( .A1(n4851), .A2(n5636), .ZN(n4850) );
  INV_X1 U5481 ( .A(n7460), .ZN(n4851) );
  OR2_X1 U5482 ( .A1(n5217), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5235) );
  INV_X1 U5483 ( .A(n4448), .ZN(n5259) );
  OR2_X1 U5484 ( .A1(n5692), .A2(n5677), .ZN(n5699) );
  AOI21_X1 U5485 ( .B1(n4848), .B2(n7537), .A(n4420), .ZN(n4847) );
  INV_X1 U5486 ( .A(n9537), .ZN(n8547) );
  OR2_X1 U5487 ( .A1(n8107), .A2(n6406), .ZN(n5138) );
  OR2_X1 U5488 ( .A1(n5104), .A2(n4582), .ZN(n4581) );
  AOI21_X1 U5489 ( .B1(n6294), .B2(P2_REG1_REG_3__SCAN_IN), .A(n4397), .ZN(
        n6327) );
  NAND2_X1 U5490 ( .A1(n4762), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n6296) );
  OAI21_X1 U5491 ( .B1(n9977), .B2(n5746), .A(n9991), .ZN(n9994) );
  NOR2_X1 U5492 ( .A1(n10013), .A2(n5814), .ZN(n10012) );
  OAI21_X1 U5493 ( .B1(n10013), .B2(n4775), .A(n4774), .ZN(n6313) );
  NAND2_X1 U5494 ( .A1(n6312), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n4775) );
  NAND2_X1 U5495 ( .A1(n4777), .A2(n6312), .ZN(n4774) );
  NAND2_X1 U5496 ( .A1(n6368), .A2(n5783), .ZN(n6357) );
  OR2_X1 U5497 ( .A1(n5756), .A2(n7058), .ZN(n4789) );
  NAND2_X1 U5498 ( .A1(n7055), .A2(n5785), .ZN(n6738) );
  NAND2_X1 U5499 ( .A1(n7183), .A2(n5788), .ZN(n7314) );
  OR2_X1 U5500 ( .A1(n8603), .A2(n4771), .ZN(n4769) );
  NAND2_X1 U5501 ( .A1(n4772), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n4771) );
  INV_X1 U5502 ( .A(n8621), .ZN(n4772) );
  OR2_X1 U5503 ( .A1(n4366), .A2(n8621), .ZN(n4770) );
  OR2_X1 U5504 ( .A1(n8603), .A2(n8604), .ZN(n4773) );
  NAND2_X1 U5505 ( .A1(n8623), .A2(n4457), .ZN(n5792) );
  OR2_X1 U5506 ( .A1(n5798), .A2(n7590), .ZN(n4457) );
  AND3_X1 U5507 ( .A1(n4769), .A2(n4770), .A3(n5764), .ZN(n5765) );
  INV_X1 U5508 ( .A(n5537), .ZN(n8662) );
  NAND2_X1 U5509 ( .A1(n5857), .A2(n8660), .ZN(n5863) );
  NAND2_X1 U5510 ( .A1(n4798), .A2(n4797), .ZN(n4796) );
  NAND2_X1 U5511 ( .A1(n8663), .A2(n4801), .ZN(n4797) );
  NAND2_X1 U5512 ( .A1(n4800), .A2(n4799), .ZN(n4798) );
  NAND2_X1 U5513 ( .A1(n4801), .A2(n5768), .ZN(n4800) );
  NAND2_X1 U5514 ( .A1(n4803), .A2(n8663), .ZN(n4802) );
  INV_X1 U5515 ( .A(n5768), .ZN(n4803) );
  OR2_X1 U5516 ( .A1(n5451), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n5467) );
  NAND2_X1 U5517 ( .A1(n4447), .A2(n6888), .ZN(n5411) );
  INV_X1 U5518 ( .A(n4447), .ZN(n5403) );
  NAND2_X1 U5519 ( .A1(n4446), .A2(n8539), .ZN(n5361) );
  NAND2_X1 U5520 ( .A1(n4894), .A2(n4893), .ZN(n5328) );
  INV_X1 U5521 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n4893) );
  INV_X1 U5522 ( .A(n5310), .ZN(n4894) );
  INV_X1 U5523 ( .A(n4446), .ZN(n5347) );
  OR2_X1 U5524 ( .A1(n5294), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5310) );
  NAND2_X1 U5525 ( .A1(n4448), .A2(n6740), .ZN(n5278) );
  NAND2_X1 U5526 ( .A1(n4892), .A2(n4891), .ZN(n5294) );
  INV_X1 U5527 ( .A(n5278), .ZN(n4892) );
  AND2_X1 U5528 ( .A1(n8018), .A2(n8017), .ZN(n7121) );
  NAND2_X1 U5529 ( .A1(n4442), .A2(n4441), .ZN(n5198) );
  INV_X1 U5530 ( .A(n5185), .ZN(n4442) );
  AND3_X1 U5531 ( .A1(n5196), .A2(n5195), .A3(n5194), .ZN(n5620) );
  NAND2_X1 U5532 ( .A1(n4443), .A2(n4888), .ZN(n5185) );
  INV_X1 U5533 ( .A(n5169), .ZN(n4443) );
  OR2_X1 U5534 ( .A1(n5153), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5169) );
  NAND2_X1 U5535 ( .A1(n6515), .A2(n5516), .ZN(n10035) );
  CLKBUF_X1 U5536 ( .A(n6510), .Z(n8135) );
  NAND2_X1 U5537 ( .A1(n5576), .A2(n5575), .ZN(n5712) );
  OR2_X1 U5538 ( .A1(n5606), .A2(n5574), .ZN(n5575) );
  NAND2_X1 U5539 ( .A1(n8586), .A2(n8809), .ZN(n5887) );
  NAND2_X1 U5540 ( .A1(n4718), .A2(n5383), .ZN(n8776) );
  AOI21_X1 U5541 ( .B1(n4576), .B2(n4579), .A(n8048), .ZN(n4574) );
  INV_X1 U5542 ( .A(n8049), .ZN(n4579) );
  AND4_X1 U5543 ( .A1(n5315), .A2(n5314), .A3(n5313), .A4(n5312), .ZN(n7584)
         );
  AOI21_X1 U5544 ( .B1(n7393), .B2(n5300), .A(n4418), .ZN(n7510) );
  OR2_X1 U5545 ( .A1(n5596), .A2(n8169), .ZN(n10086) );
  OR2_X1 U5546 ( .A1(n5673), .A2(n8134), .ZN(n5720) );
  INV_X1 U5547 ( .A(n10103), .ZN(n10112) );
  XNOR2_X1 U5548 ( .A(n5590), .B(n5589), .ZN(n5734) );
  NAND2_X1 U5549 ( .A1(n5567), .A2(n7294), .ZN(n5983) );
  INV_X1 U5550 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n5562) );
  AND2_X1 U5551 ( .A1(n5552), .A2(n5563), .ZN(n5553) );
  AND2_X1 U5552 ( .A1(n5145), .A2(n4902), .ZN(n5255) );
  INV_X1 U5553 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n5342) );
  XNOR2_X1 U5554 ( .A(n5163), .B(P2_IR_REG_6__SCAN_IN), .ZN(n10000) );
  XNOR2_X1 U5555 ( .A(n5096), .B(P2_IR_REG_2__SCAN_IN), .ZN(n9965) );
  INV_X1 U5556 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n6580) );
  OR2_X1 U5557 ( .A1(n7642), .A2(n8955), .ZN(n7728) );
  INV_X1 U5558 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n6657) );
  NOR2_X1 U5559 ( .A1(n7728), .A2(n7727), .ZN(n7747) );
  AOI21_X1 U5560 ( .B1(n4550), .B2(n4354), .A(n4398), .ZN(n4548) );
  NAND2_X1 U5561 ( .A1(n4529), .A2(n8982), .ZN(n4528) );
  INV_X1 U5562 ( .A(n4876), .ZN(n4529) );
  NOR2_X1 U5563 ( .A1(n4532), .A2(n4533), .ZN(n4531) );
  INV_X1 U5564 ( .A(n9049), .ZN(n4533) );
  INV_X1 U5565 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n6673) );
  NAND2_X1 U5566 ( .A1(n6161), .A2(n6162), .ZN(n6177) );
  NAND2_X1 U5567 ( .A1(n7356), .A2(n7355), .ZN(n4557) );
  INV_X1 U5568 ( .A(n4534), .ZN(n9027) );
  NAND2_X1 U5569 ( .A1(n4544), .A2(n4536), .ZN(n4535) );
  NOR2_X1 U5570 ( .A1(n4541), .A2(n7740), .ZN(n4536) );
  AOI21_X1 U5571 ( .B1(n7330), .B2(n7230), .A(n4354), .ZN(n7371) );
  OR2_X1 U5572 ( .A1(n7898), .A2(n7897), .ZN(n8934) );
  INV_X1 U5573 ( .A(n9225), .ZN(n9017) );
  INV_X1 U5574 ( .A(n9162), .ZN(n9052) );
  AND2_X1 U5575 ( .A1(n7755), .A2(n7754), .ZN(n9181) );
  NAND2_X1 U5576 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n4664) );
  AOI21_X1 U5577 ( .B1(n6491), .B2(P1_REG1_REG_1__SCAN_IN), .A(n9575), .ZN(
        n9590) );
  NOR2_X1 U5578 ( .A1(n9590), .A2(n9591), .ZN(n9589) );
  AND2_X1 U5579 ( .A1(n4432), .A2(n4431), .ZN(n9513) );
  NAND2_X1 U5580 ( .A1(n6493), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n4431) );
  INV_X1 U5581 ( .A(n4430), .ZN(n9512) );
  NOR2_X1 U5582 ( .A1(n9508), .A2(n4684), .ZN(n9611) );
  AND2_X1 U5583 ( .A1(n6495), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n4684) );
  AND2_X1 U5584 ( .A1(n4430), .A2(n4429), .ZN(n9615) );
  NAND2_X1 U5585 ( .A1(n6495), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n4429) );
  NOR2_X1 U5586 ( .A1(n9625), .A2(n4408), .ZN(n9646) );
  NOR2_X1 U5587 ( .A1(n9646), .A2(n9647), .ZN(n9645) );
  INV_X1 U5588 ( .A(n4679), .ZN(n9493) );
  AOI21_X1 U5589 ( .B1(P1_REG2_REG_7__SCAN_IN), .B2(n6649), .A(n9497), .ZN(
        n9524) );
  NAND2_X1 U5590 ( .A1(n9082), .A2(n6478), .ZN(n9486) );
  NOR2_X1 U5591 ( .A1(n9486), .A2(n9485), .ZN(n9484) );
  INV_X1 U5592 ( .A(n4681), .ZN(n9657) );
  AND2_X1 U5593 ( .A1(n4681), .A2(n4680), .ZN(n6503) );
  NAND2_X1 U5594 ( .A1(n9656), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n4680) );
  NAND2_X1 U5595 ( .A1(n6503), .A2(n6502), .ZN(n9097) );
  NAND2_X1 U5596 ( .A1(n9111), .A2(n9110), .ZN(n9677) );
  NOR2_X1 U5597 ( .A1(n9677), .A2(n9676), .ZN(n9675) );
  AOI21_X1 U5598 ( .B1(P1_REG2_REG_13__SCAN_IN), .B2(n9680), .A(n9675), .ZN(
        n9689) );
  NOR2_X1 U5599 ( .A1(n9700), .A2(n9102), .ZN(n9103) );
  NAND3_X1 U5600 ( .A1(n4667), .A2(n4666), .A3(n4668), .ZN(n9150) );
  OAI21_X1 U5601 ( .B1(n4672), .B2(n9139), .A(n4669), .ZN(n4668) );
  OR2_X1 U5602 ( .A1(n9136), .A2(n4671), .ZN(n4667) );
  INV_X1 U5603 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n8955) );
  INV_X1 U5604 ( .A(n9266), .ZN(n4631) );
  INV_X1 U5605 ( .A(n4375), .ZN(n4627) );
  INV_X1 U5606 ( .A(n9230), .ZN(n9241) );
  NAND2_X1 U5607 ( .A1(n9217), .A2(n8385), .ZN(n4821) );
  NAND2_X1 U5608 ( .A1(n9265), .A2(n4822), .ZN(n4817) );
  NAND2_X1 U5609 ( .A1(n9291), .A2(n4392), .ZN(n9252) );
  NAND2_X1 U5610 ( .A1(n9291), .A2(n4356), .ZN(n9267) );
  NAND2_X1 U5611 ( .A1(n4826), .A2(n9213), .ZN(n4825) );
  INV_X1 U5612 ( .A(n4828), .ZN(n4826) );
  NAND2_X1 U5613 ( .A1(n9291), .A2(n9154), .ZN(n9292) );
  NAND2_X1 U5614 ( .A1(n9363), .A2(n4464), .ZN(n9319) );
  NOR2_X1 U5615 ( .A1(n9426), .A2(n4465), .ZN(n4464) );
  INV_X1 U5616 ( .A(n4466), .ZN(n4465) );
  AND2_X1 U5617 ( .A1(n8355), .A2(n9209), .ZN(n9340) );
  AOI21_X1 U5618 ( .B1(n9349), .B2(n9180), .A(n9179), .ZN(n9333) );
  AND2_X1 U5619 ( .A1(n9435), .A2(n9178), .ZN(n9179) );
  NAND2_X1 U5620 ( .A1(n9363), .A2(n4468), .ZN(n9350) );
  AND2_X1 U5621 ( .A1(n8356), .A2(n9206), .ZN(n9356) );
  INV_X1 U5622 ( .A(n4638), .ZN(n9349) );
  OAI21_X1 U5623 ( .B1(n9362), .B2(n4640), .A(n4639), .ZN(n4638) );
  NAND2_X1 U5624 ( .A1(n9370), .A2(n9176), .ZN(n4639) );
  AND2_X1 U5625 ( .A1(n8184), .A2(n9175), .ZN(n4640) );
  AND2_X1 U5626 ( .A1(n7648), .A2(n9173), .ZN(n9363) );
  NAND2_X1 U5627 ( .A1(n9363), .A2(n9370), .ZN(n9364) );
  NAND2_X1 U5628 ( .A1(n8992), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n7490) );
  NOR2_X1 U5629 ( .A1(n9558), .A2(n9454), .ZN(n7501) );
  OR2_X1 U5630 ( .A1(n7427), .A2(n9066), .ZN(n7426) );
  NAND2_X1 U5631 ( .A1(n9556), .A2(n7269), .ZN(n4829) );
  NAND2_X1 U5632 ( .A1(n7270), .A2(n4472), .ZN(n9558) );
  NOR2_X1 U5633 ( .A1(n7427), .A2(n4473), .ZN(n4472) );
  INV_X1 U5634 ( .A(n4474), .ZN(n4473) );
  INV_X1 U5635 ( .A(n4654), .ZN(n9557) );
  OAI21_X1 U5636 ( .B1(n7253), .B2(n4657), .A(n4655), .ZN(n4654) );
  AOI21_X1 U5637 ( .B1(n4659), .B2(n4656), .A(n4658), .ZN(n4655) );
  NAND2_X1 U5638 ( .A1(n4659), .A2(n7274), .ZN(n4657) );
  INV_X1 U5639 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n7262) );
  NAND2_X1 U5640 ( .A1(n7270), .A2(n9912), .ZN(n9737) );
  NOR2_X1 U5641 ( .A1(n7154), .A2(n7153), .ZN(n7162) );
  INV_X1 U5642 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n6787) );
  AND2_X1 U5643 ( .A1(n9744), .A2(n9745), .ZN(n7147) );
  OAI21_X1 U5644 ( .B1(n7172), .B2(n8369), .A(n7171), .ZN(n9742) );
  OR2_X1 U5645 ( .A1(n7299), .A2(n9072), .ZN(n7171) );
  INV_X1 U5646 ( .A(n9744), .ZN(n9741) );
  NOR2_X1 U5647 ( .A1(n6674), .A2(n6673), .ZN(n6708) );
  AND2_X1 U5648 ( .A1(n6714), .A2(n6713), .ZN(n7376) );
  AND2_X1 U5649 ( .A1(n9774), .A2(n9881), .ZN(n6704) );
  NAND2_X1 U5650 ( .A1(n6839), .A2(n4385), .ZN(n4622) );
  AND2_X1 U5651 ( .A1(n8190), .A2(n8222), .ZN(n6702) );
  INV_X1 U5652 ( .A(n8173), .ZN(n7713) );
  AND2_X1 U5653 ( .A1(n9792), .A2(n4470), .ZN(n9774) );
  AND2_X1 U5654 ( .A1(n9772), .A2(n4471), .ZN(n4470) );
  NAND2_X1 U5655 ( .A1(n9792), .A2(n9861), .ZN(n9791) );
  NAND2_X1 U5656 ( .A1(n9792), .A2(n4471), .ZN(n9776) );
  NAND2_X1 U5657 ( .A1(n6666), .A2(n8412), .ZN(n6833) );
  AND2_X1 U5658 ( .A1(n8416), .A2(n8192), .ZN(n8365) );
  OR2_X1 U5659 ( .A1(n9805), .A2(n6686), .ZN(n9806) );
  NOR2_X1 U5660 ( .A1(n9806), .A2(n6817), .ZN(n9792) );
  OR2_X1 U5661 ( .A1(n6627), .A2(n6064), .ZN(n9775) );
  OAI21_X1 U5662 ( .B1(n9815), .B2(n9816), .A(n6625), .ZN(n6634) );
  NAND2_X1 U5663 ( .A1(n8173), .A2(n4609), .ZN(n6181) );
  AND2_X1 U5664 ( .A1(n6178), .A2(n4962), .ZN(n4609) );
  OR2_X1 U5665 ( .A1(n9836), .A2(n6622), .ZN(n9754) );
  AND2_X1 U5666 ( .A1(n8464), .A2(n6151), .ZN(n8353) );
  OR2_X1 U5667 ( .A1(n6171), .A2(n6163), .ZN(n9381) );
  NAND2_X1 U5668 ( .A1(n4630), .A2(n4628), .ZN(n9393) );
  AND2_X1 U5669 ( .A1(n4624), .A2(n4625), .ZN(n9765) );
  NAND2_X1 U5670 ( .A1(n6839), .A2(n6647), .ZN(n4624) );
  OR2_X1 U5671 ( .A1(n4347), .A2(n4734), .ZN(n4475) );
  NOR2_X1 U5672 ( .A1(n8322), .A2(n6064), .ZN(n9903) );
  INV_X1 U5673 ( .A(n9919), .ZN(n9911) );
  INV_X1 U5674 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n5999) );
  XNOR2_X1 U5675 ( .A(n7621), .B(n7620), .ZN(n8172) );
  OAI21_X1 U5676 ( .B1(n7617), .B2(n7616), .A(n7615), .ZN(n7621) );
  XNOR2_X1 U5677 ( .A(n7617), .B(n7616), .ZN(n8318) );
  XNOR2_X1 U5678 ( .A(n7566), .B(n5488), .ZN(n8309) );
  XNOR2_X1 U5679 ( .A(n5044), .B(n5484), .ZN(n7934) );
  INV_X1 U5680 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n5974) );
  XNOR2_X1 U5681 ( .A(n5904), .B(P1_IR_REG_26__SCAN_IN), .ZN(n6045) );
  NAND2_X1 U5682 ( .A1(n4365), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5904) );
  XNOR2_X1 U5683 ( .A(n5464), .B(n5463), .ZN(n7838) );
  NOR2_X1 U5684 ( .A1(n5921), .A2(n5920), .ZN(n5922) );
  OAI21_X1 U5685 ( .B1(n5925), .B2(n5918), .A(n5917), .ZN(n5923) );
  NOR2_X1 U5686 ( .A1(P1_IR_REG_24__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n5920) );
  XNOR2_X1 U5687 ( .A(n5017), .B(n5018), .ZN(n5423) );
  NAND2_X1 U5688 ( .A1(n5008), .A2(n5007), .ZN(n5009) );
  NAND2_X1 U5689 ( .A1(n5004), .A2(n4862), .ZN(n5008) );
  AND2_X1 U5690 ( .A1(n5384), .A2(SI_20_), .ZN(n5002) );
  NOR2_X1 U5691 ( .A1(n4748), .A2(n4863), .ZN(n4747) );
  INV_X1 U5692 ( .A(n5420), .ZN(n4748) );
  INV_X1 U5693 ( .A(n5422), .ZN(n4744) );
  XNOR2_X1 U5694 ( .A(n5928), .B(n5927), .ZN(n5972) );
  INV_X1 U5695 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n5927) );
  INV_X1 U5696 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5968) );
  AND2_X1 U5697 ( .A1(n6095), .A2(n6100), .ZN(n9098) );
  XNOR2_X1 U5698 ( .A(n5204), .B(n4879), .ZN(n6693) );
  NAND2_X1 U5699 ( .A1(n4727), .A2(n4970), .ZN(n5204) );
  NAND2_X1 U5700 ( .A1(n4515), .A2(n4384), .ZN(n4727) );
  AND2_X1 U5701 ( .A1(n5963), .A2(n5987), .ZN(n6653) );
  AND2_X1 U5702 ( .A1(n5947), .A2(n5959), .ZN(n6568) );
  XNOR2_X1 U5703 ( .A(n4934), .B(n4694), .ZN(n6178) );
  INV_X1 U5704 ( .A(n5068), .ZN(n4694) );
  OR2_X1 U5705 ( .A1(n5637), .A2(n7537), .ZN(n4846) );
  NAND2_X1 U5706 ( .A1(n8571), .A2(n5652), .ZN(n8504) );
  AND2_X1 U5707 ( .A1(n8111), .A2(n5495), .ZN(n8487) );
  AND2_X1 U5708 ( .A1(n8479), .A2(n8478), .ZN(n8480) );
  NAND2_X1 U5709 ( .A1(n6821), .A2(n4834), .ZN(n7083) );
  NAND2_X1 U5710 ( .A1(n5619), .A2(n4835), .ZN(n4834) );
  NAND2_X1 U5711 ( .A1(n5648), .A2(n5647), .ZN(n8537) );
  AND2_X1 U5712 ( .A1(n5637), .A2(n4850), .ZN(n7538) );
  NAND2_X1 U5713 ( .A1(n5637), .A2(n5636), .ZN(n7461) );
  NAND2_X1 U5714 ( .A1(n8513), .A2(n5659), .ZN(n8558) );
  NAND2_X1 U5715 ( .A1(n6132), .A2(n5610), .ZN(n6193) );
  INV_X1 U5716 ( .A(n8810), .ZN(n8576) );
  NAND2_X1 U5717 ( .A1(n5682), .A2(n10038), .ZN(n9539) );
  INV_X1 U5718 ( .A(n8563), .ZN(n8577) );
  OAI211_X1 U5719 ( .C1(n8107), .C2(n8743), .A(n5431), .B(n5430), .ZN(n8753)
         );
  OR2_X1 U5720 ( .A1(n5219), .A2(n6395), .ZN(n5121) );
  NAND2_X1 U5721 ( .A1(n5540), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5089) );
  INV_X1 U5722 ( .A(n10020), .ZN(n9956) );
  NOR2_X1 U5723 ( .A1(P2_U3150), .A2(n5859), .ZN(n9946) );
  NOR2_X1 U5724 ( .A1(n5758), .A2(n7061), .ZN(n6730) );
  AND2_X1 U5725 ( .A1(n6348), .A2(n5756), .ZN(n5757) );
  AND2_X1 U5726 ( .A1(n4765), .A2(n4763), .ZN(n7311) );
  INV_X1 U5727 ( .A(n4764), .ZN(n4763) );
  OAI21_X1 U5728 ( .B1(n5761), .B2(P2_REG2_REG_13__SCAN_IN), .A(n4768), .ZN(
        n4764) );
  NAND2_X1 U5729 ( .A1(n8605), .A2(n5791), .ZN(n8624) );
  NAND2_X1 U5730 ( .A1(n4769), .A2(n4770), .ZN(n8620) );
  AND2_X1 U5731 ( .A1(n4773), .A2(n4366), .ZN(n8622) );
  XNOR2_X1 U5732 ( .A(n5792), .B(n5847), .ZN(n8642) );
  OAI21_X1 U5733 ( .B1(n5767), .B2(n4791), .A(n4452), .ZN(n4451) );
  NAND2_X1 U5734 ( .A1(n4804), .A2(n4794), .ZN(n4791) );
  INV_X1 U5735 ( .A(n8673), .ZN(n4452) );
  NAND2_X1 U5736 ( .A1(n4796), .A2(n4802), .ZN(n4794) );
  NOR2_X1 U5737 ( .A1(n10024), .A2(n4792), .ZN(n4790) );
  NOR2_X1 U5738 ( .A1(n4793), .A2(n4795), .ZN(n4792) );
  NOR2_X1 U5739 ( .A1(n8663), .A2(n8657), .ZN(n4795) );
  NAND2_X1 U5740 ( .A1(n8658), .A2(n4456), .ZN(n4455) );
  OR2_X1 U5741 ( .A1(n8660), .A2(n8855), .ZN(n4456) );
  NAND2_X1 U5742 ( .A1(n4898), .A2(n5598), .ZN(n8683) );
  NAND2_X1 U5743 ( .A1(n5525), .A2(n8017), .ZN(n7206) );
  NAND2_X1 U5744 ( .A1(n5258), .A2(n5257), .ZN(n10113) );
  NAND2_X1 U5745 ( .A1(n6607), .A2(n5197), .ZN(n7074) );
  AND3_X1 U5746 ( .A1(n5182), .A2(n5181), .A3(n5180), .ZN(n10085) );
  OR2_X1 U5747 ( .A1(n8797), .A2(n6390), .ZN(n8819) );
  OR2_X1 U5748 ( .A1(n5597), .A2(n10036), .ZN(n8681) );
  NAND2_X1 U5749 ( .A1(n5982), .A2(n5709), .ZN(n10038) );
  INV_X1 U5750 ( .A(n8819), .ZN(n7399) );
  INV_X1 U5751 ( .A(n10038), .ZN(n8815) );
  INV_X1 U5752 ( .A(n8681), .ZN(n8816) );
  AOI21_X1 U5753 ( .B1(n8693), .B2(n5513), .A(n8692), .ZN(n8873) );
  NAND2_X1 U5754 ( .A1(n8691), .A2(n8690), .ZN(n8692) );
  NAND2_X1 U5755 ( .A1(n8712), .A2(n8807), .ZN(n8690) );
  NAND2_X1 U5756 ( .A1(n8711), .A2(n5458), .ZN(n8700) );
  NAND2_X1 U5757 ( .A1(n4604), .A2(n4603), .ZN(n8726) );
  NAND2_X1 U5758 ( .A1(n8752), .A2(n5419), .ZN(n8740) );
  NAND2_X1 U5759 ( .A1(n4604), .A2(n8068), .ZN(n8738) );
  NAND2_X1 U5760 ( .A1(n5391), .A2(n5390), .ZN(n8917) );
  NAND2_X1 U5761 ( .A1(n7655), .A2(n8049), .ZN(n8803) );
  NAND2_X1 U5762 ( .A1(n7579), .A2(n5336), .ZN(n7657) );
  NAND2_X1 U5763 ( .A1(n5309), .A2(n5308), .ZN(n7603) );
  NAND2_X1 U5764 ( .A1(n4597), .A2(n8037), .ZN(n7508) );
  NAND2_X1 U5765 ( .A1(n5526), .A2(n8031), .ZN(n7398) );
  NAND2_X1 U5766 ( .A1(n5276), .A2(n5275), .ZN(n7467) );
  INV_X1 U5767 ( .A(n8892), .ZN(n8927) );
  AND2_X1 U5768 ( .A1(n5216), .A2(n5215), .ZN(n7216) );
  AND2_X1 U5769 ( .A1(n5734), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8495) );
  AND2_X1 U5770 ( .A1(n5046), .A2(n4913), .ZN(n4686) );
  INV_X1 U5771 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n4913) );
  NOR2_X1 U5772 ( .A1(P2_IR_REG_27__SCAN_IN), .A2(P2_IR_REG_28__SCAN_IN), .ZN(
        n4606) );
  INV_X1 U5773 ( .A(n5802), .ZN(n7320) );
  INV_X1 U5774 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6097) );
  INV_X1 U5775 ( .A(n6741), .ZN(n6099) );
  INV_X1 U5776 ( .A(n6360), .ZN(n6037) );
  INV_X1 U5777 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6010) );
  INV_X1 U5778 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n5957) );
  NAND2_X1 U5779 ( .A1(n5071), .A2(n5095), .ZN(n5738) );
  AND2_X1 U5780 ( .A1(n5972), .A2(P1_STATE_REG_SCAN_IN), .ZN(n5966) );
  NAND2_X1 U5781 ( .A1(n8939), .A2(n7933), .ZN(n7954) );
  NAND2_X1 U5782 ( .A1(n8959), .A2(n7757), .ZN(n8960) );
  NAND2_X1 U5783 ( .A1(n4542), .A2(n7739), .ZN(n8959) );
  NAND2_X1 U5784 ( .A1(n4549), .A2(n4548), .ZN(n7358) );
  INV_X1 U5785 ( .A(n8971), .ZN(n8972) );
  INV_X1 U5786 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n6540) );
  INV_X1 U5787 ( .A(n4560), .ZN(n6567) );
  OAI21_X1 U5788 ( .B1(n6524), .B2(n6523), .A(n4564), .ZN(n4560) );
  INV_X1 U5789 ( .A(n6817), .ZN(n9855) );
  AOI21_X1 U5790 ( .B1(n7358), .B2(n7357), .A(n4553), .ZN(n7552) );
  INV_X1 U5791 ( .A(n4557), .ZN(n4553) );
  NAND2_X1 U5792 ( .A1(n6172), .A2(n9799), .ZN(n9023) );
  INV_X1 U5793 ( .A(n9023), .ZN(n9061) );
  INV_X1 U5794 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n9055) );
  INV_X1 U5795 ( .A(n9018), .ZN(n9056) );
  INV_X1 U5796 ( .A(n9036), .ZN(n9050) );
  AND2_X1 U5797 ( .A1(n8353), .A2(n9603), .ZN(n9225) );
  NAND2_X1 U5798 ( .A1(n4750), .A2(n8459), .ZN(n4749) );
  NAND2_X1 U5799 ( .A1(n8460), .A2(n8461), .ZN(n4750) );
  INV_X1 U5800 ( .A(n4752), .ZN(n4751) );
  OAI21_X1 U5801 ( .B1(n8400), .B2(n4349), .A(n6064), .ZN(n4752) );
  INV_X1 U5802 ( .A(n6075), .ZN(n8464) );
  OR2_X1 U5803 ( .A1(n7947), .A2(n7946), .ZN(n9226) );
  OR2_X1 U5804 ( .A1(n7907), .A2(n7906), .ZN(n9063) );
  OR2_X1 U5805 ( .A1(n7496), .A2(n7495), .ZN(n9171) );
  OR2_X1 U5806 ( .A1(n7441), .A2(n7440), .ZN(n9065) );
  OR2_X1 U5807 ( .A1(n7167), .A2(n7166), .ZN(n9068) );
  AND2_X1 U5808 ( .A1(n6794), .A2(n6793), .ZN(n9070) );
  OR2_X1 U5809 ( .A1(n6680), .A2(n6679), .ZN(n9073) );
  OR2_X1 U5810 ( .A1(n6663), .A2(n6662), .ZN(n9074) );
  OR2_X1 U5811 ( .A1(n6586), .A2(n6585), .ZN(n9075) );
  OR2_X1 U5812 ( .A1(n6539), .A2(n6538), .ZN(n9076) );
  OR2_X1 U5813 ( .A1(n6427), .A2(n6426), .ZN(n9077) );
  OR2_X1 U5814 ( .A1(n6266), .A2(n6265), .ZN(n9078) );
  NAND4_X2 U5815 ( .A1(n6080), .A2(n6079), .A3(n6078), .A4(n6077), .ZN(n9081)
         );
  INV_X1 U5816 ( .A(n4432), .ZN(n9593) );
  NOR2_X1 U5817 ( .A1(n9661), .A2(n4434), .ZN(n6480) );
  AND2_X1 U5818 ( .A1(n9656), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n4434) );
  NAND2_X1 U5819 ( .A1(n6480), .A2(n6481), .ZN(n9111) );
  NOR2_X1 U5820 ( .A1(n9116), .A2(n9703), .ZN(n9119) );
  OR2_X1 U5821 ( .A1(n9573), .A2(n6485), .ZN(n9702) );
  NAND2_X1 U5822 ( .A1(n4677), .A2(n4675), .ZN(n9714) );
  AND2_X1 U5823 ( .A1(n4677), .A2(n4428), .ZN(n9716) );
  NAND2_X1 U5824 ( .A1(n9136), .A2(n9135), .ZN(n4677) );
  OR2_X1 U5825 ( .A1(n9573), .A2(n9603), .ZN(n9724) );
  INV_X1 U5826 ( .A(n9702), .ZN(n9718) );
  NAND2_X1 U5827 ( .A1(n9159), .A2(n9829), .ZN(n9379) );
  INV_X1 U5828 ( .A(n9380), .ZN(n9157) );
  INV_X1 U5829 ( .A(n9156), .ZN(n9387) );
  OAI21_X1 U5830 ( .B1(n9266), .B2(n9197), .A(n4636), .ZN(n9251) );
  NAND2_X1 U5831 ( .A1(n9309), .A2(n9211), .ZN(n9296) );
  NAND2_X1 U5832 ( .A1(n4642), .A2(n4649), .ZN(n9290) );
  OR2_X1 U5833 ( .A1(n9318), .A2(n4651), .ZN(n4642) );
  OR2_X1 U5834 ( .A1(n9318), .A2(n9186), .ZN(n4652) );
  AND2_X1 U5835 ( .A1(n4812), .A2(n8324), .ZN(n9372) );
  CLKBUF_X1 U5836 ( .A(n8263), .Z(n9370) );
  AND2_X1 U5837 ( .A1(n4833), .A2(n4832), .ZN(n7484) );
  AOI21_X1 U5838 ( .B1(n9736), .B2(n9735), .A(n4662), .ZN(n7422) );
  NAND2_X1 U5839 ( .A1(n6547), .A2(n9799), .ZN(n9335) );
  INV_X1 U5840 ( .A(n9799), .ZN(n9822) );
  OR2_X1 U5841 ( .A1(n9836), .A2(n6548), .ZN(n9825) );
  MUX2_X1 U5842 ( .A(n9570), .B(n9479), .S(n8173), .Z(n9830) );
  INV_X1 U5843 ( .A(n9248), .ZN(n9832) );
  INV_X1 U5844 ( .A(n9825), .ZN(n9753) );
  INV_X1 U5845 ( .A(n9945), .ZN(n9943) );
  NAND2_X1 U5846 ( .A1(n9390), .A2(n9919), .ZN(n4478) );
  OAI21_X1 U5847 ( .B1(n6000), .B2(n5994), .A(n5993), .ZN(n5998) );
  NAND2_X1 U5848 ( .A1(n5992), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5993) );
  INV_X1 U5849 ( .A(n6151), .ZN(n8405) );
  NAND2_X1 U5850 ( .A1(n4996), .A2(n4995), .ZN(n5353) );
  AND2_X1 U5851 ( .A1(n6019), .A2(n6090), .ZN(n9489) );
  INV_X1 U5852 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n5965) );
  INV_X1 U5853 ( .A(n6491), .ZN(n9585) );
  OAI21_X1 U5854 ( .B1(n8084), .B2(n8583), .A(n5881), .ZN(n5882) );
  OAI21_X1 U5855 ( .B1(n4485), .B2(n4487), .A(n4449), .ZN(n4482) );
  NAND2_X1 U5856 ( .A1(n4484), .A2(n7112), .ZN(n4483) );
  INV_X1 U5857 ( .A(n4766), .ZN(n7181) );
  NAND2_X1 U5858 ( .A1(n5797), .A2(n10017), .ZN(n5867) );
  OAI21_X1 U5859 ( .B1(n4453), .B2(n9981), .A(n4450), .ZN(P2_U3201) );
  XNOR2_X1 U5860 ( .A(n4455), .B(n4454), .ZN(n4453) );
  NOR2_X1 U5861 ( .A1(n4451), .A2(n4383), .ZN(n4450) );
  INV_X1 U5862 ( .A(n8664), .ZN(n4454) );
  NOR2_X1 U5863 ( .A1(n5717), .A2(n5716), .ZN(n5718) );
  NOR2_X1 U5864 ( .A1(n5728), .A2(n8836), .ZN(n5717) );
  OAI21_X1 U5865 ( .B1(n8872), .B2(n8859), .A(n5892), .ZN(n5893) );
  OAI22_X1 U5866 ( .A1(n5728), .A2(n8892), .B1(n10118), .B2(n5727), .ZN(n5729)
         );
  AOI21_X1 U5867 ( .B1(n9609), .B2(P1_ADDR_REG_19__SCAN_IN), .A(n9153), .ZN(
        n4685) );
  NAND2_X1 U5868 ( .A1(n4440), .A2(n6070), .ZN(n4439) );
  OR2_X1 U5869 ( .A1(n9380), .A2(n9163), .ZN(n4351) );
  INV_X1 U5870 ( .A(n9406), .ZN(n4637) );
  INV_X2 U5871 ( .A(n7636), .ZN(n7777) );
  AND2_X1 U5872 ( .A1(n8383), .A2(n9215), .ZN(n4352) );
  AND2_X1 U5873 ( .A1(n9918), .A2(n9067), .ZN(n4353) );
  OR2_X1 U5874 ( .A1(n7229), .A2(n7228), .ZN(n4354) );
  AND2_X1 U5875 ( .A1(n7446), .A2(n9066), .ZN(n8436) );
  AND2_X1 U5876 ( .A1(n9154), .A2(n9282), .ZN(n4355) );
  NAND2_X1 U5877 ( .A1(n4818), .A2(n4391), .ZN(n9237) );
  INV_X1 U5878 ( .A(n7427), .ZN(n7446) );
  AND2_X1 U5879 ( .A1(n4637), .A2(n4355), .ZN(n4356) );
  AND2_X1 U5880 ( .A1(n7482), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n4357) );
  OR2_X1 U5881 ( .A1(n8881), .A2(n8712), .ZN(n4358) );
  NOR2_X1 U5882 ( .A1(n9218), .A2(n4823), .ZN(n4822) );
  INV_X1 U5883 ( .A(n4822), .ZN(n4816) );
  AND2_X1 U5884 ( .A1(n8326), .A2(n8260), .ZN(n4359) );
  AND2_X1 U5885 ( .A1(n9918), .A2(n7556), .ZN(n9549) );
  NOR2_X1 U5886 ( .A1(n8869), .A2(n8095), .ZN(n4360) );
  INV_X1 U5887 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n4607) );
  INV_X1 U5888 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n6124) );
  NAND2_X1 U5889 ( .A1(n9772), .A2(n6758), .ZN(n4361) );
  AND2_X1 U5890 ( .A1(n4481), .A2(n5207), .ZN(n5209) );
  INV_X1 U5891 ( .A(n5209), .ZN(n4480) );
  OR2_X1 U5892 ( .A1(n4539), .A2(n4537), .ZN(n4362) );
  INV_X1 U5893 ( .A(n7058), .ZN(n4785) );
  NAND2_X1 U5894 ( .A1(n6123), .A2(n6124), .ZN(n6122) );
  AND2_X1 U5895 ( .A1(n4424), .A2(n5420), .ZN(n4363) );
  XNOR2_X1 U5896 ( .A(n6063), .B(P1_IR_REG_20__SCAN_IN), .ZN(n6064) );
  NAND2_X1 U5897 ( .A1(n9715), .A2(n4428), .ZN(n4676) );
  AND2_X1 U5898 ( .A1(n4672), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n4364) );
  OR2_X1 U5899 ( .A1(n5919), .A2(P1_IR_REG_25__SCAN_IN), .ZN(n4365) );
  INV_X1 U5900 ( .A(n8687), .ZN(n4590) );
  INV_X1 U5901 ( .A(n5084), .ZN(n8103) );
  NAND2_X1 U5902 ( .A1(n8199), .A2(n8197), .ZN(n8191) );
  OR2_X1 U5903 ( .A1(n5800), .A2(n5763), .ZN(n4366) );
  NAND3_X1 U5904 ( .A1(n5077), .A2(n5076), .A3(n4369), .ZN(n6130) );
  NAND2_X1 U5905 ( .A1(n8503), .A2(n5656), .ZN(n8509) );
  AND2_X1 U5906 ( .A1(n6596), .A2(n8006), .ZN(n4367) );
  NAND2_X1 U5907 ( .A1(n5924), .A2(n6042), .ZN(n6157) );
  OAI21_X1 U5908 ( .B1(n8790), .B2(n4713), .A(n4711), .ZN(n8748) );
  NAND2_X1 U5909 ( .A1(n4718), .A2(n4717), .ZN(n8764) );
  OR2_X1 U5910 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n4368) );
  AND2_X1 U5911 ( .A1(n4581), .A2(n4580), .ZN(n4369) );
  AND2_X1 U5912 ( .A1(n5087), .A2(n5086), .ZN(n4370) );
  OR2_X1 U5913 ( .A1(n8852), .A2(n8810), .ZN(n4371) );
  AND2_X1 U5914 ( .A1(n4632), .A2(n4635), .ZN(n4372) );
  AND3_X1 U5915 ( .A1(n4475), .A2(n6206), .A3(n6205), .ZN(n9844) );
  NAND2_X1 U5916 ( .A1(n4918), .A2(n4917), .ZN(n5104) );
  OR3_X1 U5917 ( .A1(n8077), .A2(n8085), .A3(n8156), .ZN(n4373) );
  OR2_X1 U5918 ( .A1(n5411), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n4374) );
  OAI21_X1 U5919 ( .B1(n8699), .B2(n8080), .A(n8079), .ZN(n8686) );
  AND2_X1 U5920 ( .A1(n4634), .A2(n9217), .ZN(n4375) );
  OAI21_X1 U5921 ( .B1(n5160), .B2(n4961), .A(n4960), .ZN(n5175) );
  NAND2_X1 U5922 ( .A1(n4584), .A2(n4591), .ZN(n8122) );
  NAND2_X1 U5923 ( .A1(n4652), .A2(n4871), .ZN(n9303) );
  AND2_X1 U5924 ( .A1(n6493), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n4376) );
  AND2_X1 U5925 ( .A1(n4857), .A2(n5659), .ZN(n4377) );
  NAND2_X1 U5926 ( .A1(n7919), .A2(n7918), .ZN(n9401) );
  NAND2_X1 U5927 ( .A1(n7856), .A2(n7855), .ZN(n9411) );
  INV_X1 U5928 ( .A(n9411), .ZN(n9282) );
  OR2_X1 U5929 ( .A1(n5767), .A2(n5768), .ZN(n4378) );
  NAND2_X1 U5930 ( .A1(n9421), .A2(n9188), .ZN(n9211) );
  NOR2_X1 U5931 ( .A1(n9319), .A2(n9421), .ZN(n9291) );
  NAND2_X1 U5932 ( .A1(n5255), .A2(n4909), .ZN(n5511) );
  AND2_X1 U5933 ( .A1(n4679), .A2(n4678), .ZN(n4379) );
  NOR3_X1 U5934 ( .A1(n8381), .A2(n9304), .A3(n8380), .ZN(n4380) );
  AND2_X1 U5935 ( .A1(n8881), .A2(n8712), .ZN(n4381) );
  NAND2_X1 U5936 ( .A1(n4852), .A2(n5094), .ZN(n5128) );
  NOR2_X1 U5937 ( .A1(n5208), .A2(n5523), .ZN(n4382) );
  AND2_X1 U5938 ( .A1(n5767), .A2(n4790), .ZN(n4383) );
  NAND2_X1 U5939 ( .A1(n5094), .A2(n4899), .ZN(n5112) );
  NAND2_X1 U5940 ( .A1(n7425), .A2(n7424), .ZN(n7427) );
  INV_X1 U5941 ( .A(n4918), .ZN(n7576) );
  AND2_X1 U5942 ( .A1(n8239), .A2(n8432), .ZN(n8372) );
  OR2_X1 U5943 ( .A1(n9079), .A2(n9849), .ZN(n8196) );
  AND2_X1 U5944 ( .A1(n4516), .A2(n4513), .ZN(n4384) );
  AND2_X1 U5945 ( .A1(n8002), .A2(n7995), .ZN(n7991) );
  INV_X1 U5946 ( .A(n9426), .ZN(n9323) );
  AND2_X1 U5947 ( .A1(n6647), .A2(n4361), .ZN(n4385) );
  NAND2_X1 U5948 ( .A1(n9291), .A2(n4355), .ZN(n4463) );
  AND2_X1 U5949 ( .A1(n4506), .A2(n8070), .ZN(n4386) );
  AND2_X1 U5950 ( .A1(n9309), .A2(n4828), .ZN(n4387) );
  OR2_X1 U5951 ( .A1(n9173), .A2(n9172), .ZN(n4388) );
  NAND4_X1 U5952 ( .A1(n4912), .A2(n4911), .A3(n4910), .A4(n5560), .ZN(n4389)
         );
  INV_X1 U5953 ( .A(n8034), .ZN(n4493) );
  AND2_X1 U5954 ( .A1(n8934), .A2(n4867), .ZN(n4390) );
  AND2_X1 U5955 ( .A1(n4821), .A2(n4817), .ZN(n4391) );
  AND2_X1 U5956 ( .A1(n4356), .A2(n9257), .ZN(n4392) );
  OR2_X1 U5957 ( .A1(n9395), .A2(n9199), .ZN(n8387) );
  NAND3_X1 U5958 ( .A1(n5089), .A2(n5088), .A3(n4370), .ZN(n5101) );
  NAND2_X1 U5959 ( .A1(n4702), .A2(n4701), .ZN(n5607) );
  INV_X1 U5960 ( .A(n5607), .ZN(n5609) );
  NOR2_X1 U5961 ( .A1(n9200), .A2(n9199), .ZN(n4393) );
  NOR2_X1 U5962 ( .A1(n9308), .A2(n9188), .ZN(n4394) );
  NOR2_X1 U5963 ( .A1(n8899), .A2(n8753), .ZN(n4395) );
  INV_X1 U5964 ( .A(n4820), .ZN(n4819) );
  NAND2_X1 U5965 ( .A1(n4821), .A2(n8387), .ZN(n4820) );
  INV_X1 U5966 ( .A(n9217), .ZN(n9258) );
  INV_X1 U5967 ( .A(n8762), .ZN(n4715) );
  NOR2_X1 U5968 ( .A1(n9421), .A2(n9187), .ZN(n4396) );
  INV_X1 U5969 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5046) );
  INV_X1 U5970 ( .A(n4629), .ZN(n4628) );
  NAND2_X1 U5971 ( .A1(n4372), .A2(n9242), .ZN(n4629) );
  AND2_X1 U5972 ( .A1(n4458), .A2(n5932), .ZN(n4397) );
  INV_X1 U5973 ( .A(n4663), .ZN(n4662) );
  NAND2_X1 U5974 ( .A1(n9912), .A2(n7362), .ZN(n4663) );
  OR2_X1 U5975 ( .A1(n9454), .A2(n7442), .ZN(n8256) );
  OAI21_X1 U5976 ( .B1(n4557), .B2(n7551), .A(n7550), .ZN(n4554) );
  OAI21_X1 U5977 ( .B1(n4353), .B2(n4663), .A(n7421), .ZN(n4658) );
  INV_X1 U5978 ( .A(n8083), .ZN(n4592) );
  OR2_X1 U5979 ( .A1(n7241), .A2(n4881), .ZN(n4398) );
  OAI21_X1 U5980 ( .B1(n8029), .B2(n4493), .A(n8033), .ZN(n4492) );
  INV_X1 U5981 ( .A(n8765), .ZN(n4716) );
  AND2_X1 U5982 ( .A1(n8251), .A2(n8187), .ZN(n9556) );
  INV_X1 U5983 ( .A(n4740), .ZN(n4739) );
  NAND2_X1 U5984 ( .A1(n4358), .A2(n4381), .ZN(n4740) );
  AND2_X1 U5985 ( .A1(n4535), .A2(n4539), .ZN(n4399) );
  NAND2_X1 U5986 ( .A1(n7841), .A2(n7840), .ZN(n9406) );
  NAND2_X1 U5987 ( .A1(n5532), .A2(n8753), .ZN(n4400) );
  AND2_X1 U5988 ( .A1(n8076), .A2(n4600), .ZN(n4401) );
  AND2_X1 U5989 ( .A1(n4516), .A2(n4965), .ZN(n4402) );
  AND2_X1 U5990 ( .A1(n8038), .A2(n8149), .ZN(n4403) );
  AND2_X1 U5991 ( .A1(n8935), .A2(n8934), .ZN(n4404) );
  INV_X1 U5992 ( .A(n4445), .ZN(n5376) );
  NOR2_X1 U5993 ( .A1(n5361), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n4445) );
  AND2_X1 U5994 ( .A1(n4497), .A2(n8034), .ZN(n4405) );
  OR2_X1 U5995 ( .A1(n4541), .A2(n4538), .ZN(n4406) );
  AND2_X1 U5996 ( .A1(n4630), .A2(n4372), .ZN(n4407) );
  INV_X1 U5997 ( .A(n7775), .ZN(n4537) );
  INV_X1 U5998 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n4734) );
  AND2_X1 U5999 ( .A1(n6499), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n4408) );
  NAND2_X1 U6000 ( .A1(n7698), .A2(n7697), .ZN(n4409) );
  NAND2_X1 U6001 ( .A1(n5528), .A2(n8043), .ZN(n7655) );
  NAND2_X1 U6002 ( .A1(n7072), .A2(n5210), .ZN(n7091) );
  NAND2_X1 U6003 ( .A1(n4575), .A2(n4574), .ZN(n8787) );
  XOR2_X1 U6004 ( .A(n7555), .B(n7949), .Z(n4410) );
  OAI21_X1 U6005 ( .B1(n7117), .B2(n5269), .A(n5268), .ZN(n7345) );
  NAND2_X1 U6006 ( .A1(n5285), .A2(n7346), .ZN(n7393) );
  AND2_X1 U6007 ( .A1(n6497), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n4411) );
  INV_X1 U6008 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n4860) );
  INV_X1 U6009 ( .A(n8510), .ZN(n4840) );
  AND2_X1 U6010 ( .A1(n7501), .A2(n7631), .ZN(n7648) );
  INV_X1 U6011 ( .A(n6350), .ZN(n4781) );
  INV_X1 U6012 ( .A(n9734), .ZN(n9912) );
  OR2_X1 U6013 ( .A1(n7159), .A2(n7158), .ZN(n9069) );
  NOR2_X1 U6014 ( .A1(n4747), .A2(n4744), .ZN(n4412) );
  NAND2_X1 U6015 ( .A1(n9363), .A2(n4466), .ZN(n4469) );
  AND2_X1 U6016 ( .A1(n6568), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n4413) );
  AND2_X1 U6017 ( .A1(n5624), .A2(n8595), .ZN(n4414) );
  AND2_X1 U6018 ( .A1(n4846), .A2(n4848), .ZN(n4415) );
  AND2_X1 U6019 ( .A1(n4766), .A2(n4767), .ZN(n4416) );
  AND2_X1 U6020 ( .A1(n4528), .A2(n4409), .ZN(n4417) );
  AND2_X1 U6021 ( .A1(n7407), .A2(n8590), .ZN(n4418) );
  AND2_X1 U6022 ( .A1(n8544), .A2(n8808), .ZN(n4419) );
  INV_X1 U6023 ( .A(n4788), .ZN(n4787) );
  NAND2_X1 U6024 ( .A1(n5756), .A2(n7058), .ZN(n4788) );
  AND2_X1 U6025 ( .A1(n5640), .A2(n7609), .ZN(n4420) );
  AND2_X1 U6026 ( .A1(n4530), .A2(n4417), .ZN(n4421) );
  INV_X1 U6027 ( .A(n9772), .ZN(n9873) );
  AND2_X1 U6028 ( .A1(n6651), .A2(n6650), .ZN(n9772) );
  OAI21_X1 U6029 ( .B1(n5983), .B2(P2_D_REG_0__SCAN_IN), .A(n5984), .ZN(n5606)
         );
  AND2_X1 U6030 ( .A1(n8363), .A2(n8228), .ZN(n4422) );
  INV_X1 U6031 ( .A(n6531), .ZN(n4564) );
  XNOR2_X1 U6032 ( .A(n5971), .B(P1_IR_REG_21__SCAN_IN), .ZN(n6151) );
  AND2_X1 U6033 ( .A1(n7270), .A2(n4474), .ZN(n4423) );
  AND2_X1 U6034 ( .A1(n5923), .A2(n5922), .ZN(n6042) );
  OR2_X1 U6035 ( .A1(n5012), .A2(n5011), .ZN(n4424) );
  AND2_X1 U6036 ( .A1(n9756), .A2(n9906), .ZN(n7270) );
  INV_X1 U6037 ( .A(n10024), .ZN(n4804) );
  NAND2_X1 U6038 ( .A1(n9952), .A2(n8662), .ZN(n10024) );
  AND2_X1 U6039 ( .A1(n4559), .A2(n4558), .ZN(n4425) );
  INV_X1 U6040 ( .A(n8595), .ZN(n4479) );
  NOR2_X1 U6041 ( .A1(n8668), .A2(n5603), .ZN(n4426) );
  INV_X1 U6042 ( .A(n9543), .ZN(n8572) );
  INV_X1 U6043 ( .A(n8597), .ZN(n4835) );
  NAND4_X1 U6044 ( .A1(n5141), .A2(n5140), .A3(n5139), .A4(n5138), .ZN(n8599)
         );
  INV_X1 U6045 ( .A(n8599), .ZN(n4571) );
  INV_X1 U6046 ( .A(n8668), .ZN(n5594) );
  AND2_X1 U6047 ( .A1(n9223), .A2(n9163), .ZN(n4427) );
  OR2_X1 U6048 ( .A1(n9140), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n4428) );
  INV_X1 U6049 ( .A(n4676), .ZN(n4675) );
  INV_X1 U6050 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n4441) );
  INV_X1 U6051 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n4884) );
  INV_X1 U6052 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n7049) );
  MUX2_X1 U6053 ( .A(n6084), .B(P1_REG2_REG_1__SCAN_IN), .S(n6491), .Z(n9581)
         );
  NAND3_X1 U6054 ( .A1(n4439), .A2(n4685), .A3(n4436), .ZN(P1_U3262) );
  NAND2_X1 U6055 ( .A1(n4437), .A2(n4349), .ZN(n4436) );
  NAND2_X1 U6056 ( .A1(n4438), .A2(n9152), .ZN(n4437) );
  NAND2_X1 U6057 ( .A1(n9149), .A2(n9718), .ZN(n4438) );
  OAI22_X1 U6058 ( .A1(n9149), .A2(n9702), .B1(n9148), .B2(n9699), .ZN(n4440)
         );
  INV_X2 U6059 ( .A(n5095), .ZN(n5094) );
  INV_X1 U6060 ( .A(n4463), .ZN(n9279) );
  INV_X1 U6061 ( .A(n4469), .ZN(n9334) );
  NAND3_X1 U6062 ( .A1(n9392), .A2(n9391), .A3(n4478), .ZN(n4477) );
  OAI211_X1 U6063 ( .C1(n8165), .C2(n4483), .A(n4482), .B(n8170), .ZN(P2_U3296) );
  AND2_X1 U6064 ( .A1(n8164), .A2(n5594), .ZN(n4485) );
  OAI21_X2 U6065 ( .B1(n8164), .B2(n4489), .A(n4488), .ZN(n4487) );
  NAND3_X1 U6066 ( .A1(n4491), .A2(n4403), .A3(n4490), .ZN(n8042) );
  NAND3_X1 U6067 ( .A1(n4495), .A2(n4405), .A3(n4494), .ZN(n4491) );
  OR2_X1 U6068 ( .A1(n8025), .A2(n8023), .ZN(n4494) );
  AOI21_X1 U6069 ( .B1(n8067), .B2(n8085), .A(n8131), .ZN(n4509) );
  OAI21_X1 U6070 ( .B1(n8131), .B2(n8085), .A(n4400), .ZN(n4504) );
  NAND4_X1 U6071 ( .A1(n4501), .A2(n8076), .A3(n4499), .A4(n4498), .ZN(n8071)
         );
  NAND3_X1 U6072 ( .A1(n8070), .A2(n8131), .A3(n4500), .ZN(n4498) );
  NAND3_X1 U6073 ( .A1(n8070), .A2(n8067), .A3(n4500), .ZN(n4499) );
  INV_X1 U6074 ( .A(n8070), .ZN(n4505) );
  INV_X1 U6075 ( .A(n5160), .ZN(n4511) );
  NAND2_X1 U6076 ( .A1(n4402), .A2(n4515), .ZN(n5192) );
  NAND3_X1 U6077 ( .A1(n4512), .A2(n4963), .A3(n4517), .ZN(n4516) );
  INV_X1 U6078 ( .A(n4960), .ZN(n4517) );
  INV_X1 U6079 ( .A(n4616), .ZN(n4614) );
  NAND4_X1 U6080 ( .A1(n5897), .A2(n4618), .A3(n4526), .A4(n4525), .ZN(n4616)
         );
  NOR2_X1 U6081 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n4525) );
  NAND2_X1 U6082 ( .A1(n9048), .A2(n4531), .ZN(n4530) );
  NAND3_X1 U6083 ( .A1(n4528), .A2(n4527), .A3(n4530), .ZN(n7707) );
  NAND2_X1 U6084 ( .A1(n9047), .A2(n4876), .ZN(n8981) );
  NAND2_X1 U6085 ( .A1(n9048), .A2(n9049), .ZN(n9047) );
  INV_X1 U6086 ( .A(n8982), .ZN(n4532) );
  OAI21_X1 U6087 ( .B1(n8946), .B2(n4406), .A(n4362), .ZN(n4534) );
  INV_X1 U6088 ( .A(n7740), .ZN(n4543) );
  OAI21_X2 U6089 ( .B1(n4549), .B2(n4547), .A(n4545), .ZN(n7683) );
  OAI22_X2 U6090 ( .A1(n6524), .A2(n4561), .B1(n6566), .B2(n4564), .ZN(n6757)
         );
  NOR2_X1 U6091 ( .A1(n6531), .A2(n4563), .ZN(n4562) );
  INV_X1 U6092 ( .A(n6566), .ZN(n4563) );
  NAND3_X1 U6093 ( .A1(n4907), .A2(n4566), .A3(n4565), .ZN(n5253) );
  NAND2_X1 U6094 ( .A1(n6391), .A2(n7991), .ZN(n4573) );
  NAND2_X1 U6095 ( .A1(n4569), .A2(n4567), .ZN(n5520) );
  AND2_X1 U6096 ( .A1(n8003), .A2(n4568), .ZN(n4567) );
  NAND3_X1 U6097 ( .A1(n6596), .A2(n8006), .A3(n4572), .ZN(n4568) );
  NAND2_X1 U6098 ( .A1(n4571), .A2(n6456), .ZN(n6596) );
  NAND2_X1 U6099 ( .A1(n6402), .A2(n4367), .ZN(n6597) );
  NAND2_X1 U6100 ( .A1(n4573), .A2(n8002), .ZN(n6402) );
  NAND2_X1 U6101 ( .A1(n5528), .A2(n4576), .ZN(n4575) );
  NAND2_X1 U6102 ( .A1(n4350), .A2(n9538), .ZN(n6516) );
  INV_X1 U6103 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n4582) );
  OR2_X1 U6104 ( .A1(n8686), .A2(n4589), .ZN(n4584) );
  NAND2_X1 U6105 ( .A1(n4583), .A2(n4585), .ZN(n8120) );
  NAND2_X1 U6106 ( .A1(n8686), .A2(n4587), .ZN(n4583) );
  OR2_X1 U6107 ( .A1(n8686), .A2(n8687), .ZN(n4593) );
  NAND2_X1 U6108 ( .A1(n10111), .A2(n8027), .ZN(n7349) );
  NAND2_X1 U6109 ( .A1(n5526), .A2(n4598), .ZN(n4597) );
  NAND2_X1 U6110 ( .A1(n4597), .A2(n4595), .ZN(n5527) );
  OAI21_X1 U6111 ( .B1(n8747), .B2(n4602), .A(n4401), .ZN(n5533) );
  INV_X1 U6112 ( .A(n4603), .ZN(n4602) );
  NAND2_X1 U6113 ( .A1(n4605), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4916) );
  NAND4_X1 U6114 ( .A1(n4754), .A2(n4909), .A3(n4606), .A4(n5145), .ZN(n4605)
         );
  NAND3_X1 U6115 ( .A1(n4754), .A2(n4909), .A3(n5145), .ZN(n5048) );
  AOI21_X2 U6116 ( .B1(n7132), .B2(n7131), .A(n7130), .ZN(n7330) );
  NAND2_X1 U6117 ( .A1(n7845), .A2(n7844), .ZN(n7895) );
  NOR2_X1 U6118 ( .A1(n7559), .A2(n7558), .ZN(n7685) );
  OAI22_X2 U6119 ( .A1(n6757), .A2(n6756), .B1(n6755), .B2(n6754), .ZN(n7132)
         );
  NAND2_X1 U6120 ( .A1(n5519), .A2(n7994), .ZN(n6391) );
  NAND2_X1 U6121 ( .A1(n5609), .A2(n6518), .ZN(n5516) );
  NOR3_X1 U6122 ( .A1(n8127), .A2(n8126), .A3(n8125), .ZN(n8163) );
  INV_X1 U6123 ( .A(n6516), .ZN(n7980) );
  MUX2_X1 U6124 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n4608), .S(n9945), .Z(
        P1_U3551) );
  MUX2_X1 U6125 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n4608), .S(n9927), .Z(
        P1_U3519) );
  XNOR2_X2 U6126 ( .A(n6616), .B(n6615), .ZN(n9815) );
  OAI21_X2 U6127 ( .B1(n5919), .B2(n4610), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n4612) );
  INV_X1 U6128 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n4611) );
  NAND3_X1 U6129 ( .A1(n4614), .A2(n4805), .A3(n4613), .ZN(n6200) );
  NAND3_X1 U6130 ( .A1(n5896), .A2(n5898), .A3(n4617), .ZN(n4615) );
  NOR2_X1 U6131 ( .A1(n4616), .A2(n4615), .ZN(n6123) );
  NAND3_X1 U6132 ( .A1(n5898), .A2(n5897), .A3(n5896), .ZN(n5945) );
  INV_X1 U6133 ( .A(n6646), .ZN(n4625) );
  OAI21_X1 U6134 ( .B1(n6646), .B2(n4422), .A(n4361), .ZN(n4623) );
  NAND2_X1 U6135 ( .A1(n4622), .A2(n4621), .ZN(n4620) );
  NAND2_X1 U6136 ( .A1(n4623), .A2(n4622), .ZN(n6703) );
  NAND2_X1 U6137 ( .A1(n4631), .A2(n4375), .ZN(n4630) );
  NAND2_X1 U6138 ( .A1(n9318), .A2(n4647), .ZN(n4646) );
  NOR2_X1 U6139 ( .A1(n9577), .A2(n4664), .ZN(n9575) );
  NAND2_X1 U6140 ( .A1(n9136), .A2(n4364), .ZN(n4666) );
  NAND2_X1 U6141 ( .A1(n5045), .A2(n4686), .ZN(n7626) );
  NOR2_X2 U6142 ( .A1(n4691), .A2(n4688), .ZN(n8323) );
  NOR2_X2 U6143 ( .A1(n4690), .A2(n4689), .ZN(n4688) );
  MUX2_X1 U6144 ( .A(n8264), .B(n4693), .S(n9156), .Z(n4690) );
  OAI21_X2 U6145 ( .B1(n4692), .B2(n4427), .A(n4351), .ZN(n4691) );
  MUX2_X1 U6146 ( .A(n4693), .B(n8322), .S(n9156), .Z(n4692) );
  AOI21_X2 U6147 ( .B1(n8317), .B2(n9221), .A(n8316), .ZN(n4693) );
  INV_X1 U6148 ( .A(n4705), .ZN(n4702) );
  NAND2_X1 U6149 ( .A1(n7509), .A2(n4708), .ZN(n4707) );
  NAND2_X2 U6150 ( .A1(n4707), .A2(n4706), .ZN(n8806) );
  NAND2_X1 U6151 ( .A1(n5192), .A2(n4721), .ZN(n4720) );
  NAND2_X1 U6152 ( .A1(n4720), .A2(n4724), .ZN(n5226) );
  NAND2_X4 U6153 ( .A1(n4732), .A2(n4731), .ZN(n5052) );
  OAI21_X1 U6154 ( .B1(n5052), .B2(n4734), .A(n4733), .ZN(n4940) );
  OR2_X1 U6155 ( .A1(n8709), .A2(n8721), .ZN(n8711) );
  NAND2_X1 U6156 ( .A1(n5356), .A2(n4999), .ZN(n5370) );
  NAND2_X1 U6157 ( .A1(n5010), .A2(n5009), .ZN(n5400) );
  NAND3_X1 U6158 ( .A1(n5010), .A2(n4363), .A3(n5009), .ZN(n4745) );
  NAND3_X1 U6159 ( .A1(n5010), .A2(n5009), .A3(n4424), .ZN(n4746) );
  AOI21_X2 U6160 ( .B1(n4753), .B2(n4751), .A(n4749), .ZN(n8467) );
  OR2_X2 U6161 ( .A1(n8399), .A2(n6070), .ZN(n4753) );
  NAND2_X1 U6162 ( .A1(n6295), .A2(n6329), .ZN(n4761) );
  NAND2_X1 U6163 ( .A1(n6329), .A2(n5105), .ZN(n4760) );
  INV_X1 U6164 ( .A(n6295), .ZN(n4762) );
  NAND2_X1 U6165 ( .A1(n4761), .A2(n4759), .ZN(n6332) );
  NAND2_X1 U6166 ( .A1(n4767), .A2(n7182), .ZN(n4765) );
  XNOR2_X1 U6167 ( .A(n5760), .B(n5839), .ZN(n7182) );
  INV_X1 U6168 ( .A(n5761), .ZN(n4767) );
  INV_X1 U6169 ( .A(n7312), .ZN(n4768) );
  INV_X1 U6170 ( .A(n4773), .ZN(n8602) );
  INV_X1 U6171 ( .A(n6314), .ZN(n4777) );
  NAND2_X1 U6172 ( .A1(n6348), .A2(n4787), .ZN(n4786) );
  NAND2_X1 U6173 ( .A1(n4782), .A2(n4778), .ZN(n4784) );
  INV_X1 U6174 ( .A(n6351), .ZN(n4782) );
  NAND3_X1 U6175 ( .A1(n4786), .A2(n4789), .A3(n4784), .ZN(n7062) );
  NAND3_X1 U6176 ( .A1(n4807), .A2(n8200), .A3(n4806), .ZN(n6665) );
  NAND2_X1 U6177 ( .A1(n9804), .A2(n8196), .ZN(n4806) );
  NAND3_X1 U6178 ( .A1(n8199), .A2(n8196), .A3(n8197), .ZN(n4807) );
  NAND2_X1 U6179 ( .A1(n4808), .A2(n8196), .ZN(n6807) );
  NAND2_X1 U6180 ( .A1(n8191), .A2(n9796), .ZN(n4808) );
  NAND2_X1 U6181 ( .A1(n4812), .A2(n4810), .ZN(n9205) );
  INV_X1 U6182 ( .A(n7641), .ZN(n4809) );
  NOR2_X1 U6183 ( .A1(n7641), .A2(n7640), .ZN(n8327) );
  INV_X1 U6184 ( .A(n9205), .ZN(n9208) );
  NAND2_X1 U6185 ( .A1(n9272), .A2(n8384), .ZN(n9271) );
  NAND2_X1 U6186 ( .A1(n4813), .A2(n4815), .ZN(n9222) );
  NAND2_X1 U6187 ( .A1(n9272), .A2(n4814), .ZN(n4813) );
  OR2_X1 U6188 ( .A1(n9272), .A2(n4816), .ZN(n4818) );
  NAND2_X1 U6189 ( .A1(n9271), .A2(n9216), .ZN(n9259) );
  NAND2_X1 U6190 ( .A1(n9310), .A2(n4827), .ZN(n4824) );
  NAND2_X1 U6191 ( .A1(n4824), .A2(n4825), .ZN(n9284) );
  INV_X1 U6192 ( .A(n8375), .ZN(n4832) );
  NOR2_X2 U6193 ( .A1(n9550), .A2(n4829), .ZN(n9547) );
  INV_X1 U6194 ( .A(n4833), .ZN(n7447) );
  AOI21_X2 U6195 ( .B1(n7103), .B2(n7102), .A(n4414), .ZN(n7470) );
  OAI22_X2 U6196 ( .A1(n7083), .A2(n5622), .B1(n7106), .B2(n5621), .ZN(n7103)
         );
  NAND2_X1 U6197 ( .A1(n4836), .A2(n5883), .ZN(P2_U3154) );
  NAND3_X1 U6198 ( .A1(n5878), .A2(n4837), .A3(n8572), .ZN(n4836) );
  NAND2_X1 U6199 ( .A1(n4838), .A2(n5874), .ZN(n4837) );
  NAND2_X1 U6200 ( .A1(n5637), .A2(n4848), .ZN(n4845) );
  NAND2_X1 U6201 ( .A1(n4845), .A2(n4847), .ZN(n7605) );
  NAND2_X1 U6202 ( .A1(n8513), .A2(n4377), .ZN(n8559) );
  INV_X1 U6203 ( .A(n8557), .ZN(n4857) );
  NAND2_X1 U6204 ( .A1(n8536), .A2(n8567), .ZN(n5650) );
  NAND4_X1 U6205 ( .A1(n4909), .A2(n5145), .A3(n4902), .A4(n4860), .ZN(n5508)
         );
  NAND2_X1 U6206 ( .A1(n8481), .A2(n8480), .ZN(n8484) );
  NAND2_X1 U6207 ( .A1(n7709), .A2(n9081), .ZN(n6159) );
  NAND2_X1 U6208 ( .A1(n5095), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5096) );
  XNOR2_X1 U6209 ( .A(n6184), .B(n7949), .ZN(n6210) );
  NAND2_X1 U6210 ( .A1(n4929), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n4931) );
  INV_X1 U6211 ( .A(n5052), .ZN(n4929) );
  XNOR2_X1 U6212 ( .A(n5370), .B(n5369), .ZN(n7712) );
  NAND2_X1 U6213 ( .A1(n5991), .A2(n5990), .ZN(n6000) );
  OR2_X1 U6214 ( .A1(n5607), .A2(n6518), .ZN(n5082) );
  NAND2_X1 U6215 ( .A1(n5434), .A2(n5433), .ZN(n5460) );
  AOI21_X1 U6216 ( .B1(n5421), .B2(n5016), .A(n4861), .ZN(n5434) );
  OAI21_X1 U6217 ( .B1(n5270), .B2(SI_13_), .A(n5271), .ZN(n4987) );
  XNOR2_X1 U6218 ( .A(n5270), .B(n5272), .ZN(n7254) );
  AND2_X1 U6219 ( .A1(n5255), .A2(n5254), .ZN(n5274) );
  OR3_X1 U6220 ( .A1(n8497), .A2(n5572), .A3(n8496), .ZN(n5732) );
  OR2_X1 U6221 ( .A1(n5983), .A2(n5587), .ZN(n5675) );
  OAI21_X2 U6222 ( .B1(n8806), .B2(n5368), .A(n5367), .ZN(n8790) );
  XNOR2_X1 U6223 ( .A(n5608), .B(n5607), .ZN(n6134) );
  NOR2_X2 U6224 ( .A1(n7276), .A2(n7277), .ZN(n9550) );
  INV_X1 U6225 ( .A(n5045), .ZN(n5050) );
  OR2_X1 U6226 ( .A1(n5598), .A2(n5120), .ZN(n8111) );
  NOR2_X1 U6227 ( .A1(n6720), .A2(n6721), .ZN(n6719) );
  INV_X2 U6228 ( .A(n10120), .ZN(n10118) );
  AND3_X2 U6229 ( .A1(n5713), .A2(n5712), .A3(n5711), .ZN(n10135) );
  INV_X1 U6230 ( .A(n10135), .ZN(n5719) );
  INV_X2 U6231 ( .A(n8797), .ZN(n10050) );
  NOR2_X1 U6232 ( .A1(n5015), .A2(n5422), .ZN(n4861) );
  NOR2_X1 U6233 ( .A1(n5369), .A2(n5006), .ZN(n4862) );
  OR2_X1 U6234 ( .A1(n5398), .A2(SI_21_), .ZN(n4863) );
  OR2_X1 U6235 ( .A1(n7706), .A2(n8989), .ZN(n4864) );
  AND2_X1 U6236 ( .A1(n9888), .A2(n7223), .ZN(n4865) );
  OR2_X1 U6237 ( .A1(n6176), .A2(n7949), .ZN(n4866) );
  AND2_X1 U6238 ( .A1(n7932), .A2(n7931), .ZN(n4867) );
  AND2_X1 U6239 ( .A1(n5707), .A2(n10052), .ZN(n4868) );
  INV_X1 U6240 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5563) );
  OR2_X1 U6241 ( .A1(n9181), .A2(n9337), .ZN(n4869) );
  OR2_X1 U6242 ( .A1(n9445), .A2(n9171), .ZN(n4870) );
  XNOR2_X1 U6243 ( .A(n6518), .B(n4348), .ZN(n5608) );
  AND3_X1 U6244 ( .A1(n5323), .A2(n5322), .A3(n5321), .ZN(n4872) );
  AND2_X1 U6245 ( .A1(n5612), .A2(n6229), .ZN(n4873) );
  OR2_X1 U6246 ( .A1(n6157), .A2(n6490), .ZN(n4874) );
  OR2_X1 U6247 ( .A1(n8678), .A2(n8675), .ZN(n4875) );
  INV_X1 U6248 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n4945) );
  OR2_X1 U6249 ( .A1(n7692), .A2(n7691), .ZN(n4876) );
  INV_X1 U6250 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n4891) );
  INV_X1 U6251 ( .A(n8779), .ZN(n8754) );
  AND4_X1 U6252 ( .A1(n5408), .A2(n5407), .A3(n5406), .A4(n5405), .ZN(n8779)
         );
  AND2_X1 U6253 ( .A1(n4956), .A2(n4953), .ZN(n4877) );
  NAND2_X1 U6254 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_29__SCAN_IN), 
        .ZN(n4878) );
  INV_X1 U6255 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n4889) );
  AND2_X1 U6256 ( .A1(n4975), .A2(n4974), .ZN(n4879) );
  INV_X1 U6257 ( .A(n5847), .ZN(n8646) );
  AND2_X1 U6258 ( .A1(n5344), .A2(n5371), .ZN(n5847) );
  INV_X1 U6259 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n4938) );
  AND2_X1 U6260 ( .A1(n5673), .A2(n8125), .ZN(n8792) );
  INV_X1 U6261 ( .A(n9416), .ZN(n9154) );
  AND2_X1 U6262 ( .A1(n5548), .A2(n5547), .ZN(n4880) );
  NAND2_X1 U6263 ( .A1(n4923), .A2(n4922), .ZN(n8689) );
  AND2_X1 U6264 ( .A1(n7240), .A2(n7372), .ZN(n4881) );
  AND2_X1 U6265 ( .A1(n8391), .A2(n8390), .ZN(n4883) );
  OR2_X1 U6266 ( .A1(n7453), .A2(n7452), .ZN(n9064) );
  NAND2_X1 U6267 ( .A1(n8014), .A2(n8013), .ZN(n8024) );
  NAND2_X1 U6268 ( .A1(n8404), .A2(n8264), .ZN(n8265) );
  INV_X1 U6269 ( .A(n8358), .ZN(n8359) );
  OAI21_X1 U6270 ( .B1(n8269), .B2(n8268), .A(n8267), .ZN(n8270) );
  OAI22_X1 U6271 ( .A1(n8279), .A2(n8278), .B1(n8264), .B2(n8277), .ZN(n8281)
         );
  AND2_X1 U6272 ( .A1(n8383), .A2(n8382), .ZN(n8284) );
  AND2_X1 U6273 ( .A1(n8386), .A2(n8264), .ZN(n8287) );
  AND2_X1 U6274 ( .A1(n8387), .A2(n8287), .ZN(n8288) );
  AND2_X1 U6275 ( .A1(n8305), .A2(n8304), .ZN(n8306) );
  INV_X1 U6276 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5899) );
  OAI211_X1 U6277 ( .C1(n8095), .C2(n5476), .A(n5475), .B(n5884), .ZN(n5477)
         );
  NOR2_X1 U6278 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n4907) );
  INV_X1 U6279 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n4899) );
  OR2_X1 U6280 ( .A1(n5027), .A2(n5461), .ZN(n5033) );
  OR2_X1 U6281 ( .A1(n7383), .A2(n7477), .ZN(n5625) );
  AOI211_X1 U6282 ( .C1(n8095), .C2(n8094), .A(n8159), .B(n8099), .ZN(n8114)
         );
  INV_X1 U6283 ( .A(n8149), .ZN(n5316) );
  INV_X1 U6284 ( .A(n8143), .ZN(n5208) );
  INV_X1 U6285 ( .A(n10058), .ZN(n5100) );
  AND2_X1 U6286 ( .A1(n4901), .A2(n5161), .ZN(n4902) );
  NOR2_X1 U6287 ( .A1(n8393), .A2(n8392), .ZN(n8397) );
  OR4_X1 U6288 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_5__SCAN_IN), .ZN(n6051) );
  INV_X1 U6289 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n6057) );
  INV_X1 U6290 ( .A(n5745), .ZN(n5746) );
  NAND2_X1 U6291 ( .A1(n5752), .A2(n6372), .ZN(n5753) );
  INV_X1 U6292 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n6958) );
  INV_X1 U6293 ( .A(n7843), .ZN(n7844) );
  INV_X1 U6294 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n7489) );
  INV_X1 U6295 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n7153) );
  INV_X1 U6296 ( .A(n9074), .ZN(n6700) );
  OR2_X1 U6297 ( .A1(n5485), .A2(n5484), .ZN(n5486) );
  AND2_X1 U6298 ( .A1(n5444), .A2(n5035), .ZN(n5459) );
  NOR2_X1 U6299 ( .A1(n4991), .A2(n6964), .ZN(n4992) );
  AND2_X1 U6300 ( .A1(n4983), .A2(n5249), .ZN(n4984) );
  INV_X1 U6301 ( .A(SI_9_), .ZN(n6921) );
  NAND2_X1 U6302 ( .A1(n5052), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n4930) );
  INV_X1 U6303 ( .A(n5437), .ZN(n4896) );
  AND2_X1 U6304 ( .A1(n5632), .A2(n7526), .ZN(n5633) );
  INV_X1 U6305 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n4886) );
  INV_X1 U6306 ( .A(n5861), .ZN(n5862) );
  NAND2_X1 U6307 ( .A1(n4445), .A2(n6958), .ZN(n5392) );
  OR2_X1 U6308 ( .A1(n5983), .A2(P2_D_REG_1__SCAN_IN), .ZN(n5569) );
  INV_X1 U6309 ( .A(n8792), .ZN(n5513) );
  INV_X1 U6310 ( .A(n5571), .ZN(n5535) );
  INV_X1 U6311 ( .A(n7957), .ZN(n7943) );
  INV_X1 U6312 ( .A(n6477), .ZN(n6478) );
  AOI22_X1 U6313 ( .A1(n9226), .A2(n9225), .B1(n9224), .B2(n9223), .ZN(n9227)
         );
  AND2_X1 U6314 ( .A1(n7875), .A2(n7858), .ZN(n9280) );
  NAND2_X1 U6315 ( .A1(n8206), .A2(n6642), .ZN(n8416) );
  OAI21_X1 U6316 ( .B1(n9208), .B2(n9207), .A(n9206), .ZN(n9339) );
  OR2_X1 U6317 ( .A1(n5026), .A2(n5025), .ZN(n5461) );
  INV_X1 U6318 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n4888) );
  INV_X1 U6319 ( .A(n8741), .ZN(n8714) );
  NAND2_X1 U6320 ( .A1(n4896), .A2(n4895), .ZN(n5451) );
  OR2_X1 U6321 ( .A1(n5635), .A2(n8026), .ZN(n5636) );
  NAND2_X1 U6322 ( .A1(n5608), .A2(n5609), .ZN(n5610) );
  INV_X1 U6323 ( .A(n8580), .ZN(n8530) );
  OR2_X1 U6324 ( .A1(n5120), .A2(n10037), .ZN(n5088) );
  AOI21_X1 U6325 ( .B1(P2_REG2_REG_12__SCAN_IN), .B2(n6099), .A(n6728), .ZN(
        n5760) );
  AOI21_X1 U6326 ( .B1(P2_REG2_REG_14__SCAN_IN), .B2(n7320), .A(n7311), .ZN(
        n5763) );
  INV_X1 U6327 ( .A(n8587), .ZN(n8793) );
  INV_X1 U6328 ( .A(n8590), .ZN(n7609) );
  AND2_X2 U6329 ( .A1(n7979), .A2(n8169), .ZN(n8085) );
  NAND2_X1 U6330 ( .A1(n5569), .A2(n5568), .ZN(n5676) );
  AND2_X1 U6331 ( .A1(n8050), .A2(n8059), .ZN(n8789) );
  INV_X1 U6332 ( .A(n8807), .ZN(n10043) );
  INV_X1 U6333 ( .A(n5699), .ZN(n5724) );
  OR2_X1 U6334 ( .A1(n5230), .A2(n4915), .ZN(n5231) );
  OR2_X1 U6335 ( .A1(n5178), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n5205) );
  OR2_X1 U6336 ( .A1(n4347), .A2(n7917), .ZN(n7918) );
  XNOR2_X1 U6337 ( .A(n6255), .B(n7949), .ZN(n6440) );
  AND2_X1 U6338 ( .A1(n7711), .A2(n7710), .ZN(n9040) );
  NAND2_X1 U6339 ( .A1(n8458), .A2(n6749), .ZN(n8459) );
  AOI21_X1 U6340 ( .B1(P1_REG2_REG_16__SCAN_IN), .B2(n9128), .A(n9127), .ZN(
        n9142) );
  INV_X1 U6341 ( .A(n9291), .ZN(n9305) );
  NOR2_X1 U6342 ( .A1(n9449), .A2(n9064), .ZN(n7633) );
  NAND2_X1 U6343 ( .A1(n7146), .A2(n7145), .ZN(n7173) );
  INV_X1 U6344 ( .A(n7338), .ZN(n9888) );
  NAND2_X1 U6345 ( .A1(n8197), .A2(n8407), .ZN(n8358) );
  NAND2_X1 U6346 ( .A1(n5966), .A2(n6157), .ZN(n6171) );
  OR2_X1 U6347 ( .A1(n6129), .A2(n7112), .ZN(n8563) );
  AND2_X1 U6348 ( .A1(n5457), .A2(n5456), .ZN(n8732) );
  AND4_X1 U6349 ( .A1(n5397), .A2(n5396), .A3(n5395), .A4(n5394), .ZN(n8794)
         );
  AND4_X1 U6350 ( .A1(n5264), .A2(n5263), .A3(n5262), .A4(n5261), .ZN(n8026)
         );
  NAND2_X1 U6351 ( .A1(n5854), .A2(n5853), .ZN(n10020) );
  INV_X1 U6352 ( .A(n6348), .ZN(n6349) );
  INV_X1 U6353 ( .A(n8671), .ZN(n10029) );
  AND2_X1 U6354 ( .A1(n7972), .A2(n7966), .ZN(n8141) );
  NOR2_X1 U6355 ( .A1(n10135), .A2(n5715), .ZN(n5716) );
  INV_X1 U6356 ( .A(n8836), .ZN(n8856) );
  OR2_X1 U6357 ( .A1(n5606), .A2(n5676), .ZN(n5711) );
  AND2_X1 U6358 ( .A1(n8675), .A2(n8674), .ZN(n8862) );
  XNOR2_X1 U6359 ( .A(n8875), .B(n5873), .ZN(n8687) );
  AND2_X1 U6360 ( .A1(n8060), .A2(n8760), .ZN(n8775) );
  INV_X1 U6361 ( .A(n7656), .ZN(n8046) );
  OR2_X1 U6362 ( .A1(n10079), .A2(n10052), .ZN(n10110) );
  AND3_X1 U6363 ( .A1(n6275), .A2(n10103), .A3(n5536), .ZN(n10079) );
  AND2_X1 U6364 ( .A1(n5732), .A2(n8495), .ZN(n5982) );
  INV_X1 U6365 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5372) );
  AND2_X1 U6366 ( .A1(n6270), .A2(n8466), .ZN(n9021) );
  INV_X1 U6367 ( .A(n7226), .ZN(n7225) );
  OR2_X1 U6368 ( .A1(n7637), .A2(n7636), .ZN(n7639) );
  AND2_X1 U6369 ( .A1(n6167), .A2(n8462), .ZN(n9018) );
  AND2_X1 U6370 ( .A1(n7884), .A2(n7883), .ZN(n9195) );
  AND3_X1 U6371 ( .A1(n7287), .A2(n7286), .A3(n7285), .ZN(n7686) );
  INV_X1 U6372 ( .A(n9699), .ZN(n9713) );
  INV_X1 U6373 ( .A(n9775), .ZN(n9829) );
  AND2_X1 U6374 ( .A1(n8328), .A2(n8445), .ZN(n9371) );
  INV_X1 U6375 ( .A(n9914), .ZN(n9457) );
  NAND2_X1 U6376 ( .A1(n9817), .A2(n9921), .ZN(n9914) );
  AND3_X1 U6377 ( .A1(n6147), .A2(n6145), .A3(n6170), .ZN(n9384) );
  INV_X1 U6378 ( .A(n6074), .ZN(n6070) );
  INV_X1 U6379 ( .A(n8495), .ZN(n6128) );
  INV_X1 U6380 ( .A(n7815), .ZN(n8893) );
  AND2_X1 U6381 ( .A1(n5679), .A2(n5678), .ZN(n9543) );
  INV_X1 U6382 ( .A(n9539), .ZN(n8583) );
  NAND2_X1 U6383 ( .A1(n5473), .A2(n5472), .ZN(n8712) );
  INV_X1 U6384 ( .A(n5335), .ZN(n8588) );
  INV_X1 U6385 ( .A(n9946), .ZN(n10033) );
  NAND2_X1 U6386 ( .A1(n5867), .A2(n5866), .ZN(n5868) );
  AND2_X1 U6387 ( .A1(n6597), .A2(n6403), .ZN(n10074) );
  NAND2_X1 U6388 ( .A1(n8827), .A2(n8826), .ZN(n8829) );
  NAND2_X1 U6389 ( .A1(n10135), .A2(n10110), .ZN(n8859) );
  INV_X1 U6390 ( .A(n5729), .ZN(n5730) );
  NAND2_X1 U6391 ( .A1(n10118), .A2(n10110), .ZN(n8931) );
  AND2_X1 U6392 ( .A1(n5726), .A2(n5725), .ZN(n10120) );
  NAND2_X1 U6393 ( .A1(n5983), .A2(n5982), .ZN(n8500) );
  INV_X1 U6394 ( .A(n8169), .ZN(n7101) );
  INV_X1 U6395 ( .A(n10019), .ZN(n5956) );
  INV_X1 U6396 ( .A(n8183), .ZN(n9337) );
  OR2_X1 U6397 ( .A1(n6169), .A2(n6150), .ZN(n9036) );
  OR2_X1 U6398 ( .A1(n7960), .A2(n7959), .ZN(n9062) );
  INV_X1 U6399 ( .A(n9181), .ZN(n9170) );
  OR2_X1 U6400 ( .A1(n7268), .A2(n7267), .ZN(n9067) );
  OR2_X1 U6401 ( .A1(n9573), .A2(n9569), .ZN(n9699) );
  OR2_X1 U6402 ( .A1(n9836), .A2(n4349), .ZN(n9248) );
  INV_X1 U6403 ( .A(n9809), .ZN(n9378) );
  INV_X1 U6404 ( .A(n9335), .ZN(n9823) );
  INV_X2 U6405 ( .A(n9335), .ZN(n9836) );
  AND2_X2 U6406 ( .A1(n9384), .A2(n9383), .ZN(n9945) );
  INV_X1 U6407 ( .A(n9927), .ZN(n9926) );
  AND2_X2 U6408 ( .A1(n9384), .A2(n6545), .ZN(n9927) );
  INV_X1 U6409 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n6096) );
  OR2_X1 U6410 ( .A1(n5869), .A2(n5868), .ZN(P2_U3200) );
  NAND2_X1 U6411 ( .A1(n5895), .A2(n5894), .ZN(P2_U3487) );
  AND2_X2 U6412 ( .A1(n6268), .A2(n5966), .ZN(P1_U3973) );
  NAND2_X1 U6413 ( .A1(n4885), .A2(n4884), .ZN(n5136) );
  INV_X1 U6414 ( .A(n5136), .ZN(n4887) );
  NAND2_X1 U6415 ( .A1(n4887), .A2(n4886), .ZN(n5153) );
  INV_X1 U6416 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n4895) );
  INV_X1 U6417 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n6976) );
  INV_X1 U6418 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n6942) );
  NAND2_X1 U6419 ( .A1(n6976), .A2(n6942), .ZN(n4897) );
  NAND2_X1 U6420 ( .A1(n5059), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n4898) );
  NOR2_X1 U6421 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n4906) );
  NOR2_X1 U6422 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_13__SCAN_IN), .ZN(
        n4905) );
  NOR2_X1 U6423 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n4904) );
  NOR2_X1 U6424 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n4903) );
  NAND4_X1 U6425 ( .A1(n4906), .A2(n4905), .A3(n4904), .A4(n4903), .ZN(n4908)
         );
  NOR2_X1 U6426 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), .ZN(
        n4912) );
  NOR2_X1 U6427 ( .A1(P2_IR_REG_25__SCAN_IN), .A2(P2_IR_REG_26__SCAN_IN), .ZN(
        n4911) );
  NOR2_X1 U6428 ( .A1(P2_IR_REG_24__SCAN_IN), .A2(P2_IR_REG_23__SCAN_IN), .ZN(
        n4910) );
  INV_X1 U6429 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n4915) );
  NAND2_X1 U6430 ( .A1(n8683), .A2(n5468), .ZN(n4923) );
  INV_X1 U6431 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n8682) );
  NAND2_X1 U6432 ( .A1(n8103), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n4920) );
  NAND2_X1 U6433 ( .A1(n5540), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n4919) );
  OAI211_X1 U6434 ( .C1(n8682), .C2(n8107), .A(n4920), .B(n4919), .ZN(n4921)
         );
  INV_X1 U6435 ( .A(n4921), .ZN(n4922) );
  INV_X1 U6436 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4924) );
  NAND2_X1 U6437 ( .A1(n7049), .A2(n4924), .ZN(n4926) );
  INV_X2 U6438 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4927) );
  AND2_X1 U6439 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n4932) );
  NAND2_X1 U6440 ( .A1(n4929), .A2(n4932), .ZN(n6068) );
  AND2_X1 U6441 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n4933) );
  NAND2_X1 U6442 ( .A1(n5052), .A2(n4933), .ZN(n5080) );
  NAND2_X1 U6443 ( .A1(n6068), .A2(n5080), .ZN(n5068) );
  NAND2_X1 U6444 ( .A1(n4934), .A2(n5068), .ZN(n4937) );
  NAND2_X1 U6445 ( .A1(n4935), .A2(SI_1_), .ZN(n4936) );
  NAND2_X1 U6446 ( .A1(n4937), .A2(n4936), .ZN(n5090) );
  INV_X1 U6447 ( .A(n5091), .ZN(n4939) );
  NAND2_X1 U6448 ( .A1(n5090), .A2(n4939), .ZN(n4942) );
  NAND2_X1 U6449 ( .A1(n4940), .A2(SI_2_), .ZN(n4941) );
  NAND2_X1 U6450 ( .A1(n4942), .A2(n4941), .ZN(n5110) );
  INV_X8 U6451 ( .A(n5052), .ZN(n4962) );
  INV_X1 U6452 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n4943) );
  OR2_X1 U6453 ( .A1(n5052), .A2(n4943), .ZN(n4944) );
  INV_X1 U6454 ( .A(SI_3_), .ZN(n6999) );
  XNOR2_X1 U6455 ( .A(n4946), .B(n6999), .ZN(n5111) );
  NAND2_X1 U6456 ( .A1(n5110), .A2(n5111), .ZN(n4948) );
  NAND2_X1 U6457 ( .A1(n4946), .A2(SI_3_), .ZN(n4947) );
  NAND2_X1 U6458 ( .A1(n4948), .A2(n4947), .ZN(n5126) );
  MUX2_X1 U6459 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .S(n4962), .Z(n4954) );
  INV_X1 U6460 ( .A(n5125), .ZN(n4949) );
  NAND2_X1 U6461 ( .A1(n5126), .A2(n4949), .ZN(n5143) );
  INV_X1 U6462 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n5943) );
  INV_X1 U6463 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6526) );
  MUX2_X1 U6464 ( .A(n5943), .B(n6526), .S(n4962), .Z(n4951) );
  INV_X1 U6465 ( .A(SI_5_), .ZN(n4950) );
  NAND2_X1 U6466 ( .A1(n4951), .A2(n4950), .ZN(n4956) );
  INV_X1 U6467 ( .A(n4951), .ZN(n4952) );
  NAND2_X1 U6468 ( .A1(n4952), .A2(SI_5_), .ZN(n4953) );
  NAND2_X1 U6469 ( .A1(n4954), .A2(SI_4_), .ZN(n5142) );
  AND2_X1 U6470 ( .A1(n4877), .A2(n5142), .ZN(n4955) );
  NAND2_X1 U6471 ( .A1(n5143), .A2(n4955), .ZN(n4957) );
  NAND2_X1 U6472 ( .A1(n4957), .A2(n4956), .ZN(n5160) );
  INV_X1 U6473 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n5949) );
  INV_X1 U6474 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n5948) );
  MUX2_X1 U6475 ( .A(n5949), .B(n5948), .S(n4962), .Z(n4958) );
  XNOR2_X1 U6476 ( .A(n4958), .B(SI_6_), .ZN(n5159) );
  INV_X1 U6477 ( .A(n5159), .ZN(n4961) );
  INV_X1 U6478 ( .A(n4958), .ZN(n4959) );
  NAND2_X1 U6479 ( .A1(n4959), .A2(SI_6_), .ZN(n4960) );
  MUX2_X1 U6480 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n4962), .Z(n4964) );
  XNOR2_X1 U6481 ( .A(n4964), .B(SI_7_), .ZN(n5176) );
  INV_X1 U6482 ( .A(n5176), .ZN(n4963) );
  NAND2_X1 U6483 ( .A1(n4964), .A2(SI_7_), .ZN(n4965) );
  MUX2_X1 U6484 ( .A(n5957), .B(n5965), .S(n4962), .Z(n4967) );
  INV_X1 U6485 ( .A(SI_8_), .ZN(n4966) );
  NAND2_X1 U6486 ( .A1(n4967), .A2(n4966), .ZN(n4970) );
  INV_X1 U6487 ( .A(n4967), .ZN(n4968) );
  NAND2_X1 U6488 ( .A1(n4968), .A2(SI_8_), .ZN(n4969) );
  NAND2_X1 U6489 ( .A1(n4970), .A2(n4969), .ZN(n5191) );
  INV_X1 U6490 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n4971) );
  MUX2_X1 U6491 ( .A(n6010), .B(n4971), .S(n4962), .Z(n4972) );
  NAND2_X1 U6492 ( .A1(n4972), .A2(n6921), .ZN(n4975) );
  INV_X1 U6493 ( .A(n4972), .ZN(n4973) );
  NAND2_X1 U6494 ( .A1(n4973), .A2(SI_9_), .ZN(n4974) );
  MUX2_X1 U6495 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .S(n4962), .Z(n4977) );
  XNOR2_X1 U6496 ( .A(n4977), .B(n4976), .ZN(n5211) );
  NAND2_X1 U6497 ( .A1(n4977), .A2(SI_10_), .ZN(n4978) );
  MUX2_X1 U6498 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .S(n4962), .Z(n5242) );
  MUX2_X1 U6499 ( .A(n6097), .B(n6096), .S(n4962), .Z(n4981) );
  NAND2_X1 U6500 ( .A1(n4981), .A2(n6898), .ZN(n5250) );
  OAI21_X1 U6501 ( .B1(SI_11_), .B2(n5242), .A(n5250), .ZN(n4979) );
  INV_X1 U6502 ( .A(n4979), .ZN(n4980) );
  NAND2_X1 U6503 ( .A1(n5226), .A2(n4980), .ZN(n4985) );
  NAND3_X1 U6504 ( .A1(n5250), .A2(n5242), .A3(SI_11_), .ZN(n4983) );
  INV_X1 U6505 ( .A(n4981), .ZN(n4982) );
  NAND2_X1 U6506 ( .A1(n4982), .A2(SI_12_), .ZN(n5249) );
  NAND2_X1 U6507 ( .A1(n4985), .A2(n4984), .ZN(n5270) );
  MUX2_X1 U6508 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n4962), .Z(n5271) );
  NAND2_X1 U6509 ( .A1(n5270), .A2(SI_13_), .ZN(n4986) );
  NAND2_X1 U6510 ( .A1(n4987), .A2(n4986), .ZN(n5288) );
  MUX2_X1 U6511 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n4962), .Z(n5286) );
  NOR2_X1 U6512 ( .A1(n4988), .A2(n6959), .ZN(n4990) );
  NAND2_X1 U6513 ( .A1(n4988), .A2(n6959), .ZN(n4989) );
  OAI21_X2 U6514 ( .B1(n5288), .B2(n4990), .A(n4989), .ZN(n5304) );
  INV_X1 U6515 ( .A(SI_15_), .ZN(n5301) );
  MUX2_X1 U6516 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .S(n4962), .Z(n5302) );
  MUX2_X1 U6517 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(P2_DATAO_REG_16__SCAN_IN), 
        .S(n4962), .Z(n5317) );
  INV_X1 U6518 ( .A(n5317), .ZN(n4991) );
  MUX2_X1 U6519 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(P2_DATAO_REG_17__SCAN_IN), 
        .S(n4962), .Z(n4993) );
  XNOR2_X1 U6520 ( .A(n4993), .B(n6966), .ZN(n5338) );
  NAND2_X1 U6521 ( .A1(n5337), .A2(n5338), .ZN(n4996) );
  INV_X1 U6522 ( .A(n4993), .ZN(n4994) );
  NAND2_X1 U6523 ( .A1(n4994), .A2(n6966), .ZN(n4995) );
  MUX2_X1 U6524 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n4962), .Z(n4997) );
  NAND2_X1 U6525 ( .A1(n4997), .A2(SI_18_), .ZN(n4999) );
  OAI21_X1 U6526 ( .B1(n4997), .B2(SI_18_), .A(n4999), .ZN(n5354) );
  MUX2_X1 U6527 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(P2_DATAO_REG_19__SCAN_IN), 
        .S(n4962), .Z(n5000) );
  XNOR2_X1 U6528 ( .A(n5000), .B(SI_19_), .ZN(n5369) );
  INV_X1 U6529 ( .A(n5000), .ZN(n5001) );
  NAND2_X1 U6530 ( .A1(n5001), .A2(n6936), .ZN(n5384) );
  INV_X1 U6531 ( .A(n5370), .ZN(n5004) );
  MUX2_X1 U6532 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(P2_DATAO_REG_20__SCAN_IN), 
        .S(n4962), .Z(n5387) );
  INV_X1 U6533 ( .A(n5387), .ZN(n5003) );
  NOR2_X1 U6534 ( .A1(n5003), .A2(n5386), .ZN(n5006) );
  AND2_X1 U6535 ( .A1(n5384), .A2(n5387), .ZN(n5005) );
  OR2_X1 U6536 ( .A1(n5006), .A2(n5005), .ZN(n5007) );
  MUX2_X1 U6537 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(P2_DATAO_REG_21__SCAN_IN), 
        .S(n4962), .Z(n5398) );
  INV_X1 U6538 ( .A(n5398), .ZN(n5012) );
  INV_X1 U6539 ( .A(SI_21_), .ZN(n5011) );
  MUX2_X1 U6540 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(P2_DATAO_REG_22__SCAN_IN), 
        .S(n4962), .Z(n5013) );
  XNOR2_X1 U6541 ( .A(n5013), .B(n6886), .ZN(n5420) );
  MUX2_X1 U6542 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(P2_DATAO_REG_23__SCAN_IN), 
        .S(n4962), .Z(n5017) );
  INV_X1 U6543 ( .A(n5423), .ZN(n5015) );
  INV_X1 U6544 ( .A(n5013), .ZN(n5014) );
  NAND2_X1 U6545 ( .A1(n5014), .A2(n6886), .ZN(n5422) );
  INV_X1 U6546 ( .A(n5017), .ZN(n5019) );
  NAND2_X1 U6547 ( .A1(n5019), .A2(n5018), .ZN(n5433) );
  MUX2_X1 U6548 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(P2_DATAO_REG_26__SCAN_IN), 
        .S(n4962), .Z(n5028) );
  XNOR2_X1 U6549 ( .A(n5028), .B(n6973), .ZN(n5463) );
  INV_X1 U6550 ( .A(n5463), .ZN(n5027) );
  MUX2_X1 U6551 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(P2_DATAO_REG_25__SCAN_IN), 
        .S(n4962), .Z(n5021) );
  INV_X1 U6552 ( .A(n5021), .ZN(n5020) );
  NAND2_X1 U6553 ( .A1(n5020), .A2(n6940), .ZN(n5024) );
  INV_X1 U6554 ( .A(n5024), .ZN(n5022) );
  XNOR2_X1 U6555 ( .A(n5021), .B(n6940), .ZN(n5447) );
  INV_X1 U6556 ( .A(n5035), .ZN(n5026) );
  MUX2_X1 U6557 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(P2_DATAO_REG_24__SCAN_IN), 
        .S(n4962), .Z(n5034) );
  INV_X1 U6558 ( .A(n5034), .ZN(n5023) );
  NAND2_X1 U6559 ( .A1(n5023), .A2(n6907), .ZN(n5445) );
  AND2_X1 U6560 ( .A1(n5445), .A2(n5024), .ZN(n5025) );
  AND2_X1 U6561 ( .A1(n5433), .A2(n5033), .ZN(n5030) );
  INV_X1 U6562 ( .A(n5028), .ZN(n5029) );
  NAND2_X1 U6563 ( .A1(n5029), .A2(n6973), .ZN(n5032) );
  NAND2_X1 U6564 ( .A1(n5434), .A2(n5031), .ZN(n5041) );
  INV_X1 U6565 ( .A(n5032), .ZN(n5039) );
  INV_X1 U6566 ( .A(n5033), .ZN(n5037) );
  XNOR2_X1 U6567 ( .A(n5034), .B(n6907), .ZN(n5444) );
  AND2_X1 U6568 ( .A1(n5459), .A2(n5463), .ZN(n5036) );
  MUX2_X1 U6569 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(P2_DATAO_REG_27__SCAN_IN), 
        .S(n4962), .Z(n5042) );
  XNOR2_X1 U6570 ( .A(n5042), .B(n6918), .ZN(n5055) );
  INV_X1 U6571 ( .A(n5042), .ZN(n5043) );
  NAND2_X1 U6572 ( .A1(n5043), .A2(n6918), .ZN(n5480) );
  NAND2_X1 U6573 ( .A1(n5482), .A2(n5480), .ZN(n5044) );
  MUX2_X1 U6574 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(P2_DATAO_REG_28__SCAN_IN), 
        .S(n4962), .Z(n5478) );
  INV_X1 U6575 ( .A(SI_28_), .ZN(n6938) );
  XNOR2_X1 U6576 ( .A(n5478), .B(n6938), .ZN(n5484) );
  NAND2_X1 U6577 ( .A1(n5048), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5049) );
  NAND2_X4 U6578 ( .A1(n5051), .A2(n5050), .ZN(n5537) );
  NAND2_X2 U6579 ( .A1(n5538), .A2(n5537), .ZN(n5069) );
  AND2_X2 U6580 ( .A1(n5069), .A2(n5052), .ZN(n5092) );
  NAND2_X1 U6581 ( .A1(n7934), .A2(n5092), .ZN(n5054) );
  NAND2_X1 U6582 ( .A1(n5489), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n5053) );
  INV_X1 U6583 ( .A(n8869), .ZN(n5476) );
  XNOR2_X1 U6584 ( .A(n5056), .B(n5055), .ZN(n7916) );
  NAND2_X1 U6585 ( .A1(n7916), .A2(n5092), .ZN(n5058) );
  NAND2_X1 U6586 ( .A1(n5489), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n5057) );
  OAI21_X1 U6587 ( .B1(n5467), .B2(P2_REG3_REG_26__SCAN_IN), .A(
        P2_REG3_REG_27__SCAN_IN), .ZN(n5060) );
  NAND2_X1 U6588 ( .A1(n5060), .A2(n5059), .ZN(n8695) );
  NAND2_X1 U6589 ( .A1(n8695), .A2(n5468), .ZN(n5065) );
  INV_X1 U6590 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n8694) );
  NAND2_X1 U6591 ( .A1(n8103), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n5062) );
  NAND2_X1 U6592 ( .A1(n5540), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n5061) );
  OAI211_X1 U6593 ( .C1(n8694), .C2(n8107), .A(n5062), .B(n5061), .ZN(n5063)
         );
  INV_X1 U6594 ( .A(n5063), .ZN(n5064) );
  AND2_X1 U6595 ( .A1(n8875), .A2(n8703), .ZN(n5499) );
  INV_X1 U6596 ( .A(n5499), .ZN(n5475) );
  INV_X1 U6597 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n5066) );
  INV_X1 U6598 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n5067) );
  INV_X1 U6599 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n6138) );
  NAND2_X1 U6600 ( .A1(n5092), .A2(n6178), .ZN(n5074) );
  NAND2_X1 U6601 ( .A1(n5093), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n5073) );
  NAND2_X1 U6602 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5070) );
  MUX2_X1 U6603 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5070), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n5071) );
  INV_X1 U6604 ( .A(n5738), .ZN(n6244) );
  NAND2_X1 U6605 ( .A1(n5127), .A2(n6244), .ZN(n5072) );
  INV_X1 U6606 ( .A(n10054), .ZN(n6518) );
  NAND2_X1 U6607 ( .A1(n5607), .A2(n10054), .ZN(n7981) );
  INV_X1 U6608 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n9947) );
  OR2_X1 U6609 ( .A1(n5084), .A2(n9947), .ZN(n5077) );
  INV_X1 U6610 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n9948) );
  OR2_X1 U6611 ( .A1(n5219), .A2(n9948), .ZN(n5076) );
  INV_X1 U6612 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n5075) );
  NAND2_X1 U6613 ( .A1(n5052), .A2(SI_0_), .ZN(n5079) );
  INV_X1 U6614 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5078) );
  NAND2_X1 U6615 ( .A1(n5079), .A2(n5078), .ZN(n5081) );
  AND2_X1 U6616 ( .A1(n5081), .A2(n5080), .ZN(n8933) );
  MUX2_X1 U6617 ( .A(P2_IR_REG_0__SCAN_IN), .B(n8933), .S(n5069), .Z(n9538) );
  NAND2_X1 U6618 ( .A1(n6130), .A2(n9538), .ZN(n6511) );
  NAND2_X1 U6619 ( .A1(n6510), .A2(n6511), .ZN(n5083) );
  NAND2_X1 U6620 ( .A1(n5083), .A2(n5082), .ZN(n10040) );
  INV_X1 U6621 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n10037) );
  INV_X1 U6622 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n5775) );
  OR2_X1 U6623 ( .A1(n5084), .A2(n5775), .ZN(n5087) );
  INV_X1 U6624 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n5085) );
  OR2_X1 U6625 ( .A1(n5219), .A2(n5085), .ZN(n5086) );
  XNOR2_X1 U6626 ( .A(n5090), .B(n5091), .ZN(n5930) );
  NAND2_X1 U6627 ( .A1(n5092), .A2(n5930), .ZN(n5099) );
  BUF_X4 U6628 ( .A(n5093), .Z(n5489) );
  NAND2_X1 U6629 ( .A1(n5489), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n5098) );
  NAND2_X1 U6630 ( .A1(n5127), .A2(n9965), .ZN(n5097) );
  AND3_X2 U6631 ( .A1(n5099), .A2(n5098), .A3(n5097), .ZN(n10058) );
  NAND2_X2 U6632 ( .A1(n6229), .A2(n5100), .ZN(n7987) );
  NAND2_X1 U6633 ( .A1(n5101), .A2(n10058), .ZN(n7988) );
  NAND2_X2 U6634 ( .A1(n7987), .A2(n7988), .ZN(n10039) );
  NAND2_X1 U6635 ( .A1(n10040), .A2(n10039), .ZN(n5103) );
  OR2_X1 U6636 ( .A1(n5101), .A2(n5100), .ZN(n5102) );
  NAND2_X1 U6637 ( .A1(n5103), .A2(n5102), .ZN(n6557) );
  NAND2_X1 U6638 ( .A1(n8103), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5109) );
  OR2_X1 U6639 ( .A1(n5104), .A2(n10067), .ZN(n5108) );
  INV_X1 U6640 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n5105) );
  OR2_X1 U6641 ( .A1(n5219), .A2(n5105), .ZN(n5107) );
  OR2_X1 U6642 ( .A1(n5120), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n5106) );
  NAND4_X1 U6643 ( .A1(n5109), .A2(n5108), .A3(n5107), .A4(n5106), .ZN(n8601)
         );
  XNOR2_X1 U6644 ( .A(n5110), .B(n5111), .ZN(n6248) );
  NAND2_X1 U6645 ( .A1(n5489), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n5115) );
  NAND2_X1 U6646 ( .A1(n5112), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5113) );
  XNOR2_X1 U6647 ( .A(n5113), .B(P2_IR_REG_3__SCAN_IN), .ZN(n6302) );
  NAND2_X1 U6648 ( .A1(n5127), .A2(n6302), .ZN(n5114) );
  OAI211_X1 U6649 ( .C1(n5357), .C2(n6248), .A(n5115), .B(n5114), .ZN(n6231)
         );
  NOR2_X1 U6650 ( .A1(n8601), .A2(n6231), .ZN(n5116) );
  INV_X1 U6651 ( .A(n8601), .ZN(n10042) );
  INV_X1 U6652 ( .A(n6231), .ZN(n10064) );
  OAI22_X1 U6653 ( .A1(n6557), .A2(n5116), .B1(n10042), .B2(n10064), .ZN(n5117) );
  INV_X1 U6654 ( .A(n5117), .ZN(n6393) );
  NAND2_X1 U6655 ( .A1(n8103), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5124) );
  INV_X1 U6656 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n5118) );
  OR2_X1 U6657 ( .A1(n5104), .A2(n5118), .ZN(n5123) );
  NAND2_X1 U6658 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n5119) );
  AND2_X1 U6659 ( .A1(n5136), .A2(n5119), .ZN(n6396) );
  OR2_X1 U6660 ( .A1(n5120), .A2(n6396), .ZN(n5122) );
  INV_X1 U6661 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n6395) );
  INV_X2 U6662 ( .A(n5357), .ZN(n8102) );
  XNOR2_X1 U6663 ( .A(n5126), .B(n5125), .ZN(n5936) );
  NAND2_X1 U6664 ( .A1(n8102), .A2(n5936), .ZN(n5132) );
  NAND2_X1 U6665 ( .A1(n5489), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n5131) );
  NAND2_X1 U6666 ( .A1(n5128), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5129) );
  XNOR2_X1 U6667 ( .A(n5129), .B(P2_IR_REG_4__SCAN_IN), .ZN(n6339) );
  NAND2_X1 U6668 ( .A1(n5127), .A2(n6339), .ZN(n5130) );
  OR2_X1 U6669 ( .A1(n8600), .A2(n10070), .ZN(n8002) );
  NAND2_X1 U6670 ( .A1(n8600), .A2(n10070), .ZN(n7995) );
  INV_X1 U6671 ( .A(n7991), .ZN(n5133) );
  NAND2_X1 U6672 ( .A1(n6393), .A2(n5133), .ZN(n6392) );
  INV_X1 U6673 ( .A(n10070), .ZN(n6398) );
  OR2_X1 U6674 ( .A1(n8600), .A2(n6398), .ZN(n5134) );
  NAND2_X1 U6675 ( .A1(n6392), .A2(n5134), .ZN(n6404) );
  NAND2_X1 U6676 ( .A1(n5540), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5141) );
  INV_X1 U6677 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n5135) );
  OR2_X1 U6678 ( .A1(n5084), .A2(n5135), .ZN(n5140) );
  NAND2_X1 U6679 ( .A1(n5136), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5137) );
  AND2_X1 U6680 ( .A1(n5153), .A2(n5137), .ZN(n6453) );
  OR2_X1 U6681 ( .A1(n5120), .A2(n6453), .ZN(n5139) );
  INV_X1 U6682 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n6406) );
  NAND2_X1 U6683 ( .A1(n5143), .A2(n5142), .ZN(n5144) );
  XNOR2_X1 U6684 ( .A(n5144), .B(n4877), .ZN(n6525) );
  NAND2_X1 U6685 ( .A1(n5489), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n5148) );
  OR2_X1 U6686 ( .A1(n5145), .A2(n4915), .ZN(n5146) );
  XNOR2_X1 U6687 ( .A(n5146), .B(P2_IR_REG_5__SCAN_IN), .ZN(n9984) );
  NAND2_X1 U6688 ( .A1(n5127), .A2(n9984), .ZN(n5147) );
  OAI211_X1 U6689 ( .C1(n5357), .C2(n6525), .A(n5148), .B(n5147), .ZN(n6456)
         );
  NAND2_X1 U6690 ( .A1(n8599), .A2(n6456), .ZN(n5149) );
  NAND2_X1 U6691 ( .A1(n6404), .A2(n5149), .ZN(n5151) );
  OR2_X1 U6692 ( .A1(n8599), .A2(n6456), .ZN(n5150) );
  NAND2_X1 U6693 ( .A1(n5151), .A2(n5150), .ZN(n6594) );
  NAND2_X1 U6694 ( .A1(n8103), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5158) );
  INV_X1 U6695 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n5152) );
  OR2_X1 U6696 ( .A1(n5104), .A2(n5152), .ZN(n5157) );
  NAND2_X1 U6697 ( .A1(n5153), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5154) );
  AND2_X1 U6698 ( .A1(n5169), .A2(n5154), .ZN(n6727) );
  OR2_X1 U6699 ( .A1(n5120), .A2(n6727), .ZN(n5156) );
  INV_X1 U6700 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n5747) );
  OR2_X1 U6701 ( .A1(n5219), .A2(n5747), .ZN(n5155) );
  NAND4_X1 U6702 ( .A1(n5158), .A2(n5157), .A3(n5156), .A4(n5155), .ZN(n8598)
         );
  XNOR2_X1 U6703 ( .A(n5160), .B(n5159), .ZN(n6569) );
  NAND2_X1 U6704 ( .A1(n8102), .A2(n6569), .ZN(n5166) );
  NAND2_X1 U6705 ( .A1(n5489), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n5165) );
  AND2_X1 U6706 ( .A1(n5145), .A2(n5161), .ZN(n5162) );
  OR2_X1 U6707 ( .A1(n5162), .A2(n4915), .ZN(n5163) );
  NAND2_X1 U6708 ( .A1(n5127), .A2(n10000), .ZN(n5164) );
  OR2_X1 U6709 ( .A1(n8598), .A2(n6599), .ZN(n8008) );
  NAND2_X1 U6710 ( .A1(n8598), .A2(n6599), .ZN(n7998) );
  NAND2_X1 U6711 ( .A1(n8008), .A2(n7998), .ZN(n8138) );
  NAND2_X1 U6712 ( .A1(n6594), .A2(n8138), .ZN(n5168) );
  INV_X1 U6713 ( .A(n6599), .ZN(n10081) );
  OR2_X1 U6714 ( .A1(n8598), .A2(n10081), .ZN(n5167) );
  NAND2_X1 U6715 ( .A1(n5168), .A2(n5167), .ZN(n6463) );
  NAND2_X1 U6716 ( .A1(n5540), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5174) );
  INV_X1 U6717 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n5813) );
  OR2_X1 U6718 ( .A1(n5084), .A2(n5813), .ZN(n5173) );
  NAND2_X1 U6719 ( .A1(n5169), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5170) );
  AND2_X1 U6720 ( .A1(n5185), .A2(n5170), .ZN(n6831) );
  OR2_X1 U6721 ( .A1(n5120), .A2(n6831), .ZN(n5172) );
  INV_X1 U6722 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n5814) );
  OR2_X1 U6723 ( .A1(n8107), .A2(n5814), .ZN(n5171) );
  NAND4_X1 U6724 ( .A1(n5174), .A2(n5173), .A3(n5172), .A4(n5171), .ZN(n8597)
         );
  XNOR2_X1 U6725 ( .A(n5175), .B(n5176), .ZN(n6648) );
  NAND2_X1 U6726 ( .A1(n8102), .A2(n6648), .ZN(n5182) );
  NAND2_X1 U6727 ( .A1(n5489), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n5181) );
  INV_X1 U6728 ( .A(n5255), .ZN(n5178) );
  NAND2_X1 U6729 ( .A1(n5178), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5177) );
  MUX2_X1 U6730 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5177), .S(
        P2_IR_REG_7__SCAN_IN), .Z(n5179) );
  NAND2_X1 U6731 ( .A1(n5127), .A2(n10019), .ZN(n5180) );
  OR2_X1 U6732 ( .A1(n8597), .A2(n10085), .ZN(n7971) );
  NAND2_X1 U6733 ( .A1(n8597), .A2(n10085), .ZN(n6603) );
  NAND2_X1 U6734 ( .A1(n7971), .A2(n6603), .ZN(n8139) );
  NAND2_X1 U6735 ( .A1(n6463), .A2(n8139), .ZN(n5184) );
  INV_X1 U6736 ( .A(n10085), .ZN(n6828) );
  OR2_X1 U6737 ( .A1(n8597), .A2(n6828), .ZN(n5183) );
  NAND2_X1 U6738 ( .A1(n5184), .A2(n5183), .ZN(n6605) );
  NAND2_X1 U6739 ( .A1(n5540), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n5190) );
  INV_X1 U6740 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n5818) );
  OR2_X1 U6741 ( .A1(n5084), .A2(n5818), .ZN(n5189) );
  NAND2_X1 U6742 ( .A1(n5185), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5186) );
  AND2_X1 U6743 ( .A1(n5198), .A2(n5186), .ZN(n7086) );
  OR2_X1 U6744 ( .A1(n5120), .A2(n7086), .ZN(n5188) );
  INV_X1 U6745 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n6610) );
  OR2_X1 U6746 ( .A1(n5219), .A2(n6610), .ZN(n5187) );
  NAND4_X1 U6747 ( .A1(n5190), .A2(n5189), .A3(n5188), .A4(n5187), .ZN(n8596)
         );
  XNOR2_X1 U6748 ( .A(n5192), .B(n5191), .ZN(n6652) );
  NAND2_X1 U6749 ( .A1(n8102), .A2(n6652), .ZN(n5196) );
  NAND2_X1 U6750 ( .A1(n5489), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n5195) );
  NAND2_X1 U6751 ( .A1(n5205), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5193) );
  XNOR2_X1 U6752 ( .A(n5193), .B(P2_IR_REG_8__SCAN_IN), .ZN(n6323) );
  NAND2_X1 U6753 ( .A1(n5127), .A2(n6323), .ZN(n5194) );
  OR2_X1 U6754 ( .A1(n8596), .A2(n5620), .ZN(n7972) );
  NAND2_X1 U6755 ( .A1(n8596), .A2(n5620), .ZN(n7966) );
  OR2_X2 U6756 ( .A1(n6605), .A2(n8141), .ZN(n6607) );
  INV_X1 U6757 ( .A(n5620), .ZN(n10093) );
  NAND2_X1 U6758 ( .A1(n8596), .A2(n10093), .ZN(n5197) );
  NAND2_X1 U6759 ( .A1(n5540), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5203) );
  INV_X1 U6760 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n5822) );
  OR2_X1 U6761 ( .A1(n5084), .A2(n5822), .ZN(n5202) );
  NAND2_X1 U6762 ( .A1(n5198), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n5199) );
  AND2_X1 U6763 ( .A1(n5217), .A2(n5199), .ZN(n7107) );
  OR2_X1 U6764 ( .A1(n5120), .A2(n7107), .ZN(n5201) );
  INV_X1 U6765 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n5823) );
  OR2_X1 U6766 ( .A1(n5219), .A2(n5823), .ZN(n5200) );
  NAND4_X1 U6767 ( .A1(n5203), .A2(n5202), .A3(n5201), .A4(n5200), .ZN(n8595)
         );
  NAND2_X1 U6768 ( .A1(n5213), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5206) );
  XNOR2_X1 U6769 ( .A(n5206), .B(P2_IR_REG_9__SCAN_IN), .ZN(n6372) );
  AOI22_X1 U6770 ( .A1(n5489), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n5127), .B2(
        n6372), .ZN(n5207) );
  NAND2_X1 U6771 ( .A1(n8595), .A2(n5209), .ZN(n7967) );
  OR2_X1 U6772 ( .A1(n8595), .A2(n4480), .ZN(n5210) );
  XNOR2_X1 U6773 ( .A(n5212), .B(n5211), .ZN(n6773) );
  NAND2_X1 U6774 ( .A1(n6773), .A2(n8102), .ZN(n5216) );
  NOR2_X1 U6775 ( .A1(n5213), .A2(P2_IR_REG_9__SCAN_IN), .ZN(n5229) );
  OR2_X1 U6776 ( .A1(n5229), .A2(n4915), .ZN(n5214) );
  AOI22_X1 U6777 ( .A1(n5489), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n5127), .B2(
        n6360), .ZN(n5215) );
  NAND2_X1 U6778 ( .A1(n5540), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5223) );
  INV_X1 U6779 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n5829) );
  OR2_X1 U6780 ( .A1(n5084), .A2(n5829), .ZN(n5222) );
  NAND2_X1 U6781 ( .A1(n5217), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5218) );
  AND2_X1 U6782 ( .A1(n5235), .A2(n5218), .ZN(n7392) );
  OR2_X1 U6783 ( .A1(n5120), .A2(n7392), .ZN(n5221) );
  INV_X1 U6784 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7095) );
  OR2_X1 U6785 ( .A1(n5219), .A2(n7095), .ZN(n5220) );
  NAND4_X1 U6786 ( .A1(n5223), .A2(n5222), .A3(n5221), .A4(n5220), .ZN(n8594)
         );
  NAND2_X1 U6787 ( .A1(n7216), .A2(n8594), .ZN(n8019) );
  NAND2_X1 U6788 ( .A1(n7477), .A2(n7389), .ZN(n8016) );
  NAND2_X1 U6789 ( .A1(n8019), .A2(n8016), .ZN(n7093) );
  NAND2_X1 U6790 ( .A1(n7091), .A2(n7093), .ZN(n5225) );
  OR2_X1 U6791 ( .A1(n8594), .A2(n7389), .ZN(n5224) );
  NAND2_X1 U6792 ( .A1(n5225), .A2(n5224), .ZN(n7117) );
  XNOR2_X1 U6793 ( .A(n5242), .B(SI_11_), .ZN(n5227) );
  XNOR2_X1 U6794 ( .A(n5245), .B(n5227), .ZN(n7144) );
  NAND2_X1 U6795 ( .A1(n7144), .A2(n8102), .ZN(n5233) );
  AND2_X1 U6796 ( .A1(n5229), .A2(n5228), .ZN(n5230) );
  XNOR2_X1 U6797 ( .A(n5231), .B(P2_IR_REG_11__SCAN_IN), .ZN(n7058) );
  AOI22_X1 U6798 ( .A1(n5489), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n5127), .B2(
        n7058), .ZN(n5232) );
  NAND2_X1 U6799 ( .A1(n5233), .A2(n5232), .ZN(n7123) );
  NAND2_X1 U6800 ( .A1(n5540), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5241) );
  INV_X1 U6801 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n5234) );
  OR2_X1 U6802 ( .A1(n8107), .A2(n5234), .ZN(n5240) );
  NAND2_X1 U6803 ( .A1(n5235), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5236) );
  AND2_X1 U6804 ( .A1(n5259), .A2(n5236), .ZN(n7474) );
  OR2_X1 U6805 ( .A1(n5120), .A2(n7474), .ZN(n5239) );
  INV_X1 U6806 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n5237) );
  OR2_X1 U6807 ( .A1(n5084), .A2(n5237), .ZN(n5238) );
  NAND4_X1 U6808 ( .A1(n5241), .A2(n5240), .A3(n5239), .A4(n5238), .ZN(n8593)
         );
  NOR2_X1 U6809 ( .A1(n7123), .A2(n8593), .ZN(n7197) );
  NAND2_X1 U6810 ( .A1(n5245), .A2(SI_11_), .ZN(n5244) );
  INV_X1 U6811 ( .A(n5242), .ZN(n5243) );
  NAND2_X1 U6812 ( .A1(n5244), .A2(n5243), .ZN(n5248) );
  INV_X1 U6813 ( .A(n5245), .ZN(n5246) );
  INV_X1 U6814 ( .A(SI_11_), .ZN(n6906) );
  NAND2_X1 U6815 ( .A1(n5246), .A2(n6906), .ZN(n5247) );
  NAND2_X1 U6816 ( .A1(n5248), .A2(n5247), .ZN(n5252) );
  AND2_X1 U6817 ( .A1(n5250), .A2(n5249), .ZN(n5251) );
  NAND2_X1 U6818 ( .A1(n7149), .A2(n8102), .ZN(n5258) );
  INV_X1 U6819 ( .A(n5253), .ZN(n5254) );
  OR2_X1 U6820 ( .A1(n5274), .A2(n4915), .ZN(n5256) );
  XNOR2_X1 U6821 ( .A(n5256), .B(P2_IR_REG_12__SCAN_IN), .ZN(n6741) );
  AOI22_X1 U6822 ( .A1(n5489), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n5127), .B2(
        n6741), .ZN(n5257) );
  NAND2_X1 U6823 ( .A1(n5540), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5264) );
  INV_X1 U6824 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n7204) );
  OR2_X1 U6825 ( .A1(n8107), .A2(n7204), .ZN(n5263) );
  NAND2_X1 U6826 ( .A1(n5259), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5260) );
  AND2_X1 U6827 ( .A1(n5278), .A2(n5260), .ZN(n7532) );
  OR2_X1 U6828 ( .A1(n5120), .A2(n7532), .ZN(n5262) );
  INV_X1 U6829 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n5837) );
  OR2_X1 U6830 ( .A1(n5084), .A2(n5837), .ZN(n5261) );
  XNOR2_X1 U6831 ( .A(n10113), .B(n8026), .ZN(n8030) );
  INV_X1 U6832 ( .A(n8030), .ZN(n5265) );
  OR2_X1 U6833 ( .A1(n7197), .A2(n5265), .ZN(n5269) );
  NAND2_X1 U6834 ( .A1(n7123), .A2(n8593), .ZN(n7198) );
  OR2_X1 U6835 ( .A1(n5265), .A2(n7198), .ZN(n5267) );
  INV_X1 U6836 ( .A(n8026), .ZN(n8592) );
  NAND2_X1 U6837 ( .A1(n10113), .A2(n8592), .ZN(n5266) );
  AND2_X1 U6838 ( .A1(n5267), .A2(n5266), .ZN(n5268) );
  XNOR2_X1 U6839 ( .A(n5271), .B(SI_13_), .ZN(n5272) );
  NAND2_X1 U6840 ( .A1(n7254), .A2(n8102), .ZN(n5276) );
  NAND2_X1 U6841 ( .A1(n5274), .A2(n5273), .ZN(n5320) );
  NAND2_X1 U6842 ( .A1(n5320), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5289) );
  XNOR2_X1 U6843 ( .A(n5289), .B(P2_IR_REG_13__SCAN_IN), .ZN(n5839) );
  AOI22_X1 U6844 ( .A1(n5489), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n5127), .B2(
        n5839), .ZN(n5275) );
  NAND2_X1 U6845 ( .A1(n5540), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5284) );
  INV_X1 U6846 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n5277) );
  OR2_X1 U6847 ( .A1(n5084), .A2(n5277), .ZN(n5283) );
  NAND2_X1 U6848 ( .A1(n5278), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n5279) );
  AND2_X1 U6849 ( .A1(n5294), .A2(n5279), .ZN(n7465) );
  OR2_X1 U6850 ( .A1(n5120), .A2(n7465), .ZN(n5282) );
  INV_X1 U6851 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n5280) );
  OR2_X1 U6852 ( .A1(n8107), .A2(n5280), .ZN(n5281) );
  NAND4_X1 U6853 ( .A1(n5284), .A2(n5283), .A3(n5282), .A4(n5281), .ZN(n8591)
         );
  OR2_X1 U6854 ( .A1(n7467), .A2(n8591), .ZN(n7347) );
  NAND2_X1 U6855 ( .A1(n7345), .A2(n7347), .ZN(n5285) );
  NAND2_X1 U6856 ( .A1(n7467), .A2(n8591), .ZN(n7346) );
  XNOR2_X1 U6857 ( .A(n5286), .B(SI_14_), .ZN(n5287) );
  XNOR2_X1 U6858 ( .A(n5288), .B(n5287), .ZN(n7257) );
  NAND2_X1 U6859 ( .A1(n7257), .A2(n8102), .ZN(n5292) );
  NAND2_X1 U6860 ( .A1(n5289), .A2(n5322), .ZN(n5290) );
  NAND2_X1 U6861 ( .A1(n5290), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5305) );
  XNOR2_X1 U6862 ( .A(n5305), .B(P2_IR_REG_14__SCAN_IN), .ZN(n5802) );
  AOI22_X1 U6863 ( .A1(n5489), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n5127), .B2(
        n5802), .ZN(n5291) );
  NAND2_X1 U6864 ( .A1(n5540), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5299) );
  INV_X1 U6865 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n5293) );
  OR2_X1 U6866 ( .A1(n8107), .A2(n5293), .ZN(n5298) );
  NAND2_X1 U6867 ( .A1(n5294), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5295) );
  AND2_X1 U6868 ( .A1(n5310), .A2(n5295), .ZN(n7540) );
  OR2_X1 U6869 ( .A1(n5120), .A2(n7540), .ZN(n5297) );
  INV_X1 U6870 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n7406) );
  OR2_X1 U6871 ( .A1(n5084), .A2(n7406), .ZN(n5296) );
  NAND4_X1 U6872 ( .A1(n5299), .A2(n5298), .A3(n5297), .A4(n5296), .ZN(n8590)
         );
  OR2_X1 U6873 ( .A1(n7407), .A2(n8590), .ZN(n5300) );
  XNOR2_X1 U6874 ( .A(n5302), .B(n5301), .ZN(n5303) );
  XNOR2_X1 U6875 ( .A(n5304), .B(n5303), .ZN(n7423) );
  NAND2_X1 U6876 ( .A1(n7423), .A2(n8102), .ZN(n5309) );
  NAND2_X1 U6877 ( .A1(n5305), .A2(n5323), .ZN(n5306) );
  NAND2_X1 U6878 ( .A1(n5306), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5307) );
  XNOR2_X1 U6879 ( .A(n5307), .B(P2_IR_REG_15__SCAN_IN), .ZN(n5800) );
  AOI22_X1 U6880 ( .A1(n5489), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n5127), .B2(
        n5800), .ZN(n5308) );
  NAND2_X1 U6881 ( .A1(n5540), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n5315) );
  INV_X1 U6882 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n7515) );
  OR2_X1 U6883 ( .A1(n5084), .A2(n7515), .ZN(n5314) );
  NAND2_X1 U6884 ( .A1(n5310), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n5311) );
  AND2_X1 U6885 ( .A1(n5328), .A2(n5311), .ZN(n7519) );
  OR2_X1 U6886 ( .A1(n5120), .A2(n7519), .ZN(n5313) );
  INV_X1 U6887 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n8604) );
  OR2_X1 U6888 ( .A1(n8107), .A2(n8604), .ZN(n5312) );
  NAND2_X1 U6889 ( .A1(n7603), .A2(n7584), .ZN(n8039) );
  NAND2_X1 U6890 ( .A1(n7510), .A2(n5316), .ZN(n7509) );
  XNOR2_X1 U6891 ( .A(n5317), .B(SI_16_), .ZN(n5318) );
  XNOR2_X1 U6892 ( .A(n5319), .B(n5318), .ZN(n7430) );
  NAND2_X1 U6893 ( .A1(n7430), .A2(n8102), .ZN(n5327) );
  INV_X1 U6894 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n5321) );
  NAND2_X1 U6895 ( .A1(n5339), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5325) );
  XNOR2_X1 U6896 ( .A(n5325), .B(P2_IR_REG_16__SCAN_IN), .ZN(n5798) );
  AOI22_X1 U6897 ( .A1(n5489), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n5127), .B2(
        n5798), .ZN(n5326) );
  NAND2_X1 U6898 ( .A1(n5540), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n5333) );
  INV_X1 U6899 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n7590) );
  OR2_X1 U6900 ( .A1(n5084), .A2(n7590), .ZN(n5332) );
  NAND2_X1 U6901 ( .A1(n5328), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5329) );
  AND2_X1 U6902 ( .A1(n5347), .A2(n5329), .ZN(n7677) );
  OR2_X1 U6903 ( .A1(n5120), .A2(n7677), .ZN(n5331) );
  INV_X1 U6904 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n7594) );
  OR2_X1 U6905 ( .A1(n8107), .A2(n7594), .ZN(n5330) );
  NAND2_X1 U6906 ( .A1(n7679), .A2(n5335), .ZN(n8044) );
  NAND2_X1 U6907 ( .A1(n8043), .A2(n8044), .ZN(n7580) );
  INV_X1 U6908 ( .A(n7584), .ZN(n8589) );
  OR2_X1 U6909 ( .A1(n7603), .A2(n8589), .ZN(n7581) );
  AND2_X1 U6910 ( .A1(n7580), .A2(n7581), .ZN(n5334) );
  NAND2_X1 U6911 ( .A1(n7679), .A2(n8588), .ZN(n5336) );
  XNOR2_X1 U6912 ( .A(n5337), .B(n5338), .ZN(n7485) );
  NAND2_X1 U6913 ( .A1(n7485), .A2(n8102), .ZN(n5346) );
  NOR2_X1 U6914 ( .A1(n5343), .A2(n4915), .ZN(n5340) );
  MUX2_X1 U6915 ( .A(n4915), .B(n5340), .S(P2_IR_REG_17__SCAN_IN), .Z(n5341)
         );
  INV_X1 U6916 ( .A(n5341), .ZN(n5344) );
  NAND2_X1 U6917 ( .A1(n5343), .A2(n5342), .ZN(n5371) );
  AOI22_X1 U6918 ( .A1(n5489), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n5847), .B2(
        n5127), .ZN(n5345) );
  NAND2_X1 U6919 ( .A1(n5540), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n5352) );
  INV_X1 U6920 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n7667) );
  OR2_X1 U6921 ( .A1(n5084), .A2(n7667), .ZN(n5351) );
  NAND2_X1 U6922 ( .A1(n5347), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n5348) );
  AND2_X1 U6923 ( .A1(n5361), .A2(n5348), .ZN(n8542) );
  OR2_X1 U6924 ( .A1(n5120), .A2(n8542), .ZN(n5350) );
  INV_X1 U6925 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n7662) );
  OR2_X1 U6926 ( .A1(n8107), .A2(n7662), .ZN(n5349) );
  NAND2_X1 U6927 ( .A1(n8544), .A2(n7674), .ZN(n8049) );
  NAND2_X1 U6928 ( .A1(n8802), .A2(n8049), .ZN(n7656) );
  INV_X1 U6929 ( .A(n7674), .ZN(n8808) );
  NAND2_X1 U6930 ( .A1(n5353), .A2(n5354), .ZN(n5355) );
  NAND2_X1 U6931 ( .A1(n5356), .A2(n5355), .ZN(n7637) );
  OR2_X1 U6932 ( .A1(n7637), .A2(n5357), .ZN(n5360) );
  NAND2_X1 U6933 ( .A1(n5371), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5358) );
  XNOR2_X1 U6934 ( .A(n5358), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8660) );
  AOI22_X1 U6935 ( .A1(n5489), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n5127), .B2(
        n8660), .ZN(n5359) );
  NAND2_X1 U6936 ( .A1(n5540), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n5366) );
  INV_X1 U6937 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8855) );
  OR2_X1 U6938 ( .A1(n5084), .A2(n8855), .ZN(n5365) );
  NAND2_X1 U6939 ( .A1(n5361), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5362) );
  AND2_X1 U6940 ( .A1(n5376), .A2(n5362), .ZN(n8813) );
  OR2_X1 U6941 ( .A1(n5120), .A2(n8813), .ZN(n5364) );
  INV_X1 U6942 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8812) );
  OR2_X1 U6943 ( .A1(n8107), .A2(n8812), .ZN(n5363) );
  NAND4_X1 U6944 ( .A1(n5366), .A2(n5365), .A3(n5364), .A4(n5363), .ZN(n8587)
         );
  AND2_X1 U6945 ( .A1(n8928), .A2(n8587), .ZN(n5368) );
  INV_X1 U6946 ( .A(n8928), .ZN(n8584) );
  NAND2_X1 U6947 ( .A1(n8584), .A2(n8793), .ZN(n5367) );
  NAND2_X1 U6948 ( .A1(n7712), .A2(n8102), .ZN(n5375) );
  OAI21_X2 U6949 ( .B1(n5371), .B2(P2_IR_REG_18__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5373) );
  XNOR2_X2 U6950 ( .A(n5373), .B(n5372), .ZN(n8668) );
  AOI22_X1 U6951 ( .A1(n5489), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n5594), .B2(
        n5127), .ZN(n5374) );
  NAND2_X1 U6952 ( .A1(n5540), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n5382) );
  INV_X1 U6953 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n8853) );
  OR2_X1 U6954 ( .A1(n5084), .A2(n8853), .ZN(n5381) );
  NAND2_X1 U6955 ( .A1(n5376), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n5377) );
  AND2_X1 U6956 ( .A1(n5392), .A2(n5377), .ZN(n8795) );
  OR2_X1 U6957 ( .A1(n5120), .A2(n8795), .ZN(n5380) );
  INV_X1 U6958 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n5378) );
  OR2_X1 U6959 ( .A1(n8107), .A2(n5378), .ZN(n5379) );
  NAND4_X1 U6960 ( .A1(n5382), .A2(n5381), .A3(n5380), .A4(n5379), .ZN(n8810)
         );
  NAND2_X1 U6961 ( .A1(n8852), .A2(n8810), .ZN(n5383) );
  XNOR2_X1 U6962 ( .A(n5387), .B(n5386), .ZN(n5388) );
  NAND2_X1 U6963 ( .A1(n7723), .A2(n8102), .ZN(n5391) );
  NAND2_X1 U6964 ( .A1(n5489), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n5390) );
  NAND2_X1 U6965 ( .A1(n8103), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n5397) );
  INV_X1 U6966 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n8915) );
  OR2_X1 U6967 ( .A1(n5104), .A2(n8915), .ZN(n5396) );
  NAND2_X1 U6968 ( .A1(n5392), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n5393) );
  AND2_X1 U6969 ( .A1(n5403), .A2(n5393), .ZN(n8783) );
  OR2_X1 U6970 ( .A1(n8783), .A2(n5120), .ZN(n5395) );
  INV_X1 U6971 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n8782) );
  OR2_X1 U6972 ( .A1(n8107), .A2(n8782), .ZN(n5394) );
  NAND2_X1 U6973 ( .A1(n8917), .A2(n8794), .ZN(n8760) );
  INV_X1 U6974 ( .A(n8794), .ZN(n8767) );
  OR2_X1 U6975 ( .A1(n8917), .A2(n8767), .ZN(n8765) );
  XNOR2_X1 U6976 ( .A(n5398), .B(SI_21_), .ZN(n5399) );
  XNOR2_X2 U6977 ( .A(n5400), .B(n5399), .ZN(n7743) );
  NAND2_X1 U6978 ( .A1(n7743), .A2(n8102), .ZN(n5402) );
  NAND2_X1 U6979 ( .A1(n5489), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n5401) );
  NAND2_X1 U6980 ( .A1(n5403), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n5404) );
  NAND2_X1 U6981 ( .A1(n5411), .A2(n5404), .ZN(n8771) );
  NAND2_X1 U6982 ( .A1(n5468), .A2(n8771), .ZN(n5408) );
  INV_X1 U6983 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n8845) );
  OR2_X1 U6984 ( .A1(n5084), .A2(n8845), .ZN(n5407) );
  INV_X1 U6985 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n8910) );
  OR2_X1 U6986 ( .A1(n5104), .A2(n8910), .ZN(n5406) );
  INV_X1 U6987 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n8770) );
  OR2_X1 U6988 ( .A1(n8107), .A2(n8770), .ZN(n5405) );
  NAND2_X1 U6989 ( .A1(n8911), .A2(n8779), .ZN(n5530) );
  NAND2_X1 U6990 ( .A1(n8063), .A2(n5530), .ZN(n8762) );
  OR2_X1 U6991 ( .A1(n8911), .A2(n8754), .ZN(n8749) );
  NAND2_X1 U6992 ( .A1(n8748), .A2(n8749), .ZN(n5418) );
  XNOR2_X1 U6993 ( .A(n5421), .B(n5420), .ZN(n7762) );
  NAND2_X1 U6994 ( .A1(n7762), .A2(n8102), .ZN(n5410) );
  NAND2_X1 U6995 ( .A1(n5489), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n5409) );
  NAND2_X1 U6996 ( .A1(n5411), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n5412) );
  NAND2_X1 U6997 ( .A1(n4374), .A2(n5412), .ZN(n8757) );
  NAND2_X1 U6998 ( .A1(n8757), .A2(n5468), .ZN(n5417) );
  NAND2_X1 U6999 ( .A1(n8103), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n5416) );
  NAND2_X1 U7000 ( .A1(n5540), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n5415) );
  INV_X1 U7001 ( .A(n8107), .ZN(n5413) );
  NAND2_X1 U7002 ( .A1(n5413), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n5414) );
  NAND2_X1 U7003 ( .A1(n8905), .A2(n7833), .ZN(n8069) );
  NAND2_X1 U7004 ( .A1(n8068), .A2(n8069), .ZN(n8131) );
  OR2_X1 U7005 ( .A1(n8905), .A2(n8768), .ZN(n5419) );
  NAND2_X1 U7006 ( .A1(n7778), .A2(n8102), .ZN(n5426) );
  NAND2_X1 U7007 ( .A1(n5489), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n5425) );
  NAND2_X2 U7008 ( .A1(n5426), .A2(n5425), .ZN(n8899) );
  INV_X1 U7009 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n8743) );
  NAND2_X1 U7010 ( .A1(n4374), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n5427) );
  NAND2_X1 U7011 ( .A1(n5437), .A2(n5427), .ZN(n8744) );
  NAND2_X1 U7012 ( .A1(n8744), .A2(n5468), .ZN(n5431) );
  NAND2_X1 U7013 ( .A1(n8103), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n5429) );
  NAND2_X1 U7014 ( .A1(n5540), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n5428) );
  AND2_X1 U7015 ( .A1(n5429), .A2(n5428), .ZN(n5430) );
  NAND2_X1 U7016 ( .A1(n8899), .A2(n8753), .ZN(n5432) );
  XNOR2_X1 U7017 ( .A(n5460), .B(n5444), .ZN(n7846) );
  NAND2_X1 U7018 ( .A1(n7846), .A2(n8102), .ZN(n5436) );
  NAND2_X1 U7019 ( .A1(n5489), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n5435) );
  INV_X1 U7020 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n5441) );
  NAND2_X1 U7021 ( .A1(n5437), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n5438) );
  NAND2_X1 U7022 ( .A1(n5451), .A2(n5438), .ZN(n8733) );
  NAND2_X1 U7023 ( .A1(n8733), .A2(n5468), .ZN(n5440) );
  AOI22_X1 U7024 ( .A1(n8103), .A2(P2_REG1_REG_24__SCAN_IN), .B1(n5540), .B2(
        P2_REG0_REG_24__SCAN_IN), .ZN(n5439) );
  NOR2_X1 U7025 ( .A1(n7815), .A2(n8741), .ZN(n5443) );
  NAND2_X1 U7026 ( .A1(n7815), .A2(n8741), .ZN(n5442) );
  OAI21_X2 U7027 ( .B1(n8728), .B2(n5443), .A(n5442), .ZN(n8709) );
  NAND2_X1 U7028 ( .A1(n5460), .A2(n5444), .ZN(n5446) );
  NAND2_X1 U7029 ( .A1(n5446), .A2(n5445), .ZN(n5448) );
  NAND2_X1 U7030 ( .A1(n7853), .A2(n8102), .ZN(n5450) );
  NAND2_X1 U7031 ( .A1(n5489), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n5449) );
  NAND2_X2 U7032 ( .A1(n5450), .A2(n5449), .ZN(n8887) );
  NAND2_X1 U7033 ( .A1(n5451), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n5452) );
  NAND2_X1 U7034 ( .A1(n5467), .A2(n5452), .ZN(n8717) );
  NAND2_X1 U7035 ( .A1(n8717), .A2(n5468), .ZN(n5457) );
  INV_X1 U7036 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n8722) );
  NAND2_X1 U7037 ( .A1(n5540), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n5454) );
  NAND2_X1 U7038 ( .A1(n8103), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n5453) );
  OAI211_X1 U7039 ( .C1(n8722), .C2(n8107), .A(n5454), .B(n5453), .ZN(n5455)
         );
  INV_X1 U7040 ( .A(n5455), .ZN(n5456) );
  NAND2_X1 U7041 ( .A1(n8887), .A2(n8732), .ZN(n8072) );
  AND2_X2 U7042 ( .A1(n7965), .A2(n8072), .ZN(n8721) );
  OR2_X1 U7043 ( .A1(n8887), .A2(n8702), .ZN(n5458) );
  NAND2_X1 U7044 ( .A1(n5460), .A2(n5459), .ZN(n5462) );
  NAND2_X1 U7045 ( .A1(n5462), .A2(n5461), .ZN(n5464) );
  NAND2_X1 U7046 ( .A1(n7838), .A2(n8102), .ZN(n5466) );
  NAND2_X1 U7047 ( .A1(n5489), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n5465) );
  XNOR2_X1 U7048 ( .A(n5467), .B(P2_REG3_REG_26__SCAN_IN), .ZN(n8706) );
  NAND2_X1 U7049 ( .A1(n8706), .A2(n5468), .ZN(n5473) );
  INV_X1 U7050 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n8705) );
  NAND2_X1 U7051 ( .A1(n8103), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n5470) );
  NAND2_X1 U7052 ( .A1(n5540), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n5469) );
  OAI211_X1 U7053 ( .C1(n8705), .C2(n8107), .A(n5470), .B(n5469), .ZN(n5471)
         );
  INV_X1 U7054 ( .A(n5471), .ZN(n5472) );
  OR2_X1 U7055 ( .A1(n8875), .A2(n8703), .ZN(n5474) );
  INV_X1 U7056 ( .A(n5477), .ZN(n5496) );
  INV_X1 U7057 ( .A(n5478), .ZN(n5479) );
  NAND2_X1 U7058 ( .A1(n5479), .A2(n6938), .ZN(n5483) );
  AND2_X1 U7059 ( .A1(n5480), .A2(n5483), .ZN(n5481) );
  NAND2_X1 U7060 ( .A1(n5482), .A2(n5481), .ZN(n5487) );
  INV_X1 U7061 ( .A(n5483), .ZN(n5485) );
  MUX2_X1 U7062 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .S(n4962), .Z(n7567) );
  INV_X1 U7063 ( .A(SI_29_), .ZN(n5488) );
  NAND2_X1 U7064 ( .A1(n8309), .A2(n5092), .ZN(n5491) );
  NAND2_X1 U7065 ( .A1(n5489), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n5490) );
  NAND2_X1 U7066 ( .A1(n5491), .A2(n5490), .ZN(n5714) );
  INV_X1 U7067 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n5599) );
  NAND2_X1 U7068 ( .A1(n5540), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n5493) );
  NAND2_X1 U7069 ( .A1(n8103), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n5492) );
  OAI211_X1 U7070 ( .C1(n8107), .C2(n5599), .A(n5493), .B(n5492), .ZN(n5494)
         );
  INV_X1 U7071 ( .A(n5494), .ZN(n5495) );
  NAND2_X1 U7072 ( .A1(n5714), .A2(n8487), .ZN(n8121) );
  NAND2_X1 U7073 ( .A1(n5496), .A2(n8087), .ZN(n5505) );
  NOR2_X1 U7074 ( .A1(n8869), .A2(n8689), .ZN(n5497) );
  NOR3_X1 U7075 ( .A1(n5884), .A2(n5497), .A3(n8087), .ZN(n5503) );
  INV_X1 U7076 ( .A(n5497), .ZN(n5501) );
  INV_X1 U7077 ( .A(n8689), .ZN(n8095) );
  AOI21_X1 U7078 ( .B1(n8095), .B2(n5475), .A(n5476), .ZN(n5498) );
  AOI211_X1 U7079 ( .C1(n5499), .C2(n8689), .A(n5498), .B(n8087), .ZN(n5500)
         );
  AOI21_X1 U7080 ( .B1(n8087), .B2(n5501), .A(n5500), .ZN(n5502) );
  NOR2_X1 U7081 ( .A1(n5503), .A2(n5502), .ZN(n5504) );
  NAND2_X1 U7082 ( .A1(n5505), .A2(n5504), .ZN(n5514) );
  INV_X1 U7083 ( .A(n5561), .ZN(n5506) );
  NAND2_X1 U7084 ( .A1(n5506), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5507) );
  NAND2_X1 U7085 ( .A1(n5594), .A2(n8169), .ZN(n5673) );
  AND2_X1 U7086 ( .A1(n5508), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5509) );
  MUX2_X1 U7087 ( .A(n4915), .B(n5509), .S(P2_IR_REG_21__SCAN_IN), .Z(n5510)
         );
  NAND2_X1 U7088 ( .A1(n5511), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5512) );
  INV_X1 U7089 ( .A(n8115), .ZN(n5570) );
  NAND2_X1 U7090 ( .A1(n7979), .A2(n5570), .ZN(n8125) );
  NAND2_X1 U7091 ( .A1(n5514), .A2(n5513), .ZN(n5549) );
  INV_X1 U7092 ( .A(n9538), .ZN(n6141) );
  INV_X1 U7093 ( .A(n6510), .ZN(n5515) );
  NAND2_X1 U7094 ( .A1(n7980), .A2(n5515), .ZN(n6515) );
  INV_X1 U7095 ( .A(n10039), .ZN(n5517) );
  NAND2_X1 U7096 ( .A1(n10035), .A2(n5517), .ZN(n5518) );
  NAND2_X1 U7097 ( .A1(n5518), .A2(n7987), .ZN(n6559) );
  XNOR2_X1 U7098 ( .A(n8601), .B(n6231), .ZN(n8136) );
  NAND2_X1 U7099 ( .A1(n6559), .A2(n8136), .ZN(n5519) );
  OR2_X1 U7100 ( .A1(n8601), .A2(n10064), .ZN(n7994) );
  INV_X1 U7101 ( .A(n6456), .ZN(n10073) );
  NAND2_X1 U7102 ( .A1(n8599), .A2(n10073), .ZN(n8006) );
  AND2_X1 U7103 ( .A1(n6596), .A2(n8008), .ZN(n8003) );
  NAND2_X1 U7104 ( .A1(n5520), .A2(n7998), .ZN(n6461) );
  INV_X1 U7105 ( .A(n8139), .ZN(n6460) );
  NAND2_X1 U7106 ( .A1(n6461), .A2(n6460), .ZN(n6459) );
  AND2_X1 U7107 ( .A1(n6603), .A2(n7966), .ZN(n7970) );
  NAND2_X1 U7108 ( .A1(n6459), .A2(n7970), .ZN(n5521) );
  INV_X1 U7109 ( .A(n7077), .ZN(n5522) );
  INV_X1 U7110 ( .A(n8016), .ZN(n5523) );
  NAND2_X1 U7111 ( .A1(n5522), .A2(n4382), .ZN(n7120) );
  OR2_X1 U7112 ( .A1(n7123), .A2(n7525), .ZN(n8018) );
  NAND2_X1 U7113 ( .A1(n7123), .A2(n7525), .ZN(n8017) );
  AND2_X1 U7114 ( .A1(n8019), .A2(n7967), .ZN(n7969) );
  OR2_X1 U7115 ( .A1(n5523), .A2(n7969), .ZN(n7119) );
  AND2_X1 U7116 ( .A1(n7121), .A2(n7119), .ZN(n5524) );
  NAND2_X1 U7117 ( .A1(n7120), .A2(n5524), .ZN(n5525) );
  OR2_X1 U7118 ( .A1(n10113), .A2(n8026), .ZN(n8027) );
  INV_X1 U7119 ( .A(n8591), .ZN(n7528) );
  NAND2_X1 U7120 ( .A1(n7467), .A2(n7528), .ZN(n8032) );
  NAND2_X1 U7121 ( .A1(n7349), .A2(n8032), .ZN(n5526) );
  OR2_X1 U7122 ( .A1(n7467), .A2(n7528), .ZN(n8031) );
  NOR2_X1 U7123 ( .A1(n7407), .A2(n7609), .ZN(n8035) );
  NAND2_X1 U7124 ( .A1(n7407), .A2(n7609), .ZN(n8037) );
  NAND2_X1 U7125 ( .A1(n5527), .A2(n8040), .ZN(n7578) );
  NAND2_X1 U7126 ( .A1(n7578), .A2(n8044), .ZN(n5528) );
  NAND2_X1 U7127 ( .A1(n8584), .A2(n8587), .ZN(n8801) );
  AND2_X1 U7128 ( .A1(n8801), .A2(n8802), .ZN(n8132) );
  NAND2_X1 U7129 ( .A1(n8928), .A2(n8793), .ZN(n8800) );
  NAND2_X1 U7130 ( .A1(n8852), .A2(n8576), .ZN(n8059) );
  NAND2_X1 U7131 ( .A1(n8787), .A2(n8789), .ZN(n5529) );
  NAND2_X1 U7132 ( .A1(n8774), .A2(n8060), .ZN(n8761) );
  AND2_X1 U7133 ( .A1(n5530), .A2(n8760), .ZN(n8065) );
  NAND2_X1 U7134 ( .A1(n8761), .A2(n8065), .ZN(n5531) );
  NAND2_X1 U7135 ( .A1(n5531), .A2(n8063), .ZN(n8747) );
  INV_X1 U7136 ( .A(n8899), .ZN(n5532) );
  NAND2_X1 U7137 ( .A1(n7815), .A2(n8714), .ZN(n8129) );
  INV_X1 U7138 ( .A(n8753), .ZN(n8731) );
  NAND2_X1 U7139 ( .A1(n8899), .A2(n8731), .ZN(n8725) );
  AND2_X1 U7140 ( .A1(n8129), .A2(n8725), .ZN(n8076) );
  NAND2_X1 U7141 ( .A1(n5533), .A2(n8130), .ZN(n8720) );
  NAND2_X1 U7142 ( .A1(n8720), .A2(n8072), .ZN(n5534) );
  NAND2_X1 U7143 ( .A1(n5534), .A2(n7965), .ZN(n8699) );
  NOR2_X1 U7144 ( .A1(n8881), .A2(n8529), .ZN(n8080) );
  NAND2_X1 U7145 ( .A1(n8881), .A2(n8529), .ZN(n8079) );
  OR2_X1 U7146 ( .A1(n8875), .A2(n5873), .ZN(n8083) );
  XNOR2_X1 U7147 ( .A(n8122), .B(n8087), .ZN(n5707) );
  NAND2_X1 U7148 ( .A1(n7979), .A2(n8115), .ZN(n5603) );
  INV_X1 U7149 ( .A(n7979), .ZN(n7070) );
  NAND2_X1 U7150 ( .A1(n8668), .A2(n8115), .ZN(n5604) );
  NAND2_X1 U7151 ( .A1(n5604), .A2(n5535), .ZN(n5536) );
  NAND2_X1 U7152 ( .A1(n5707), .A2(n10079), .ZN(n5548) );
  INV_X1 U7153 ( .A(n5538), .ZN(n8166) );
  NAND2_X1 U7154 ( .A1(n8662), .A2(n8166), .ZN(n5539) );
  NAND2_X1 U7155 ( .A1(n5069), .A2(n5539), .ZN(n5697) );
  INV_X1 U7156 ( .A(n5697), .ZN(n5695) );
  INV_X1 U7157 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n5543) );
  NAND2_X1 U7158 ( .A1(n8103), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n5542) );
  NAND2_X1 U7159 ( .A1(n5540), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n5541) );
  OAI211_X1 U7160 ( .C1(n5543), .C2(n8107), .A(n5542), .B(n5541), .ZN(n5544)
         );
  INV_X1 U7161 ( .A(n5544), .ZN(n5545) );
  NAND2_X1 U7162 ( .A1(n8111), .A2(n5545), .ZN(n8585) );
  AND2_X1 U7163 ( .A1(n5069), .A2(P2_B_REG_SCAN_IN), .ZN(n5546) );
  NOR2_X1 U7164 ( .A1(n10041), .A2(n5546), .ZN(n8674) );
  AOI22_X1 U7165 ( .A1(n8689), .A2(n8807), .B1(n8585), .B2(n8674), .ZN(n5547)
         );
  AND2_X1 U7166 ( .A1(n5707), .A2(n4426), .ZN(n5595) );
  NAND2_X1 U7167 ( .A1(n5561), .A2(n5552), .ZN(n5550) );
  NAND2_X1 U7168 ( .A1(n5550), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5551) );
  NAND2_X1 U7169 ( .A1(n5561), .A2(n5553), .ZN(n5557) );
  OR2_X1 U7170 ( .A1(P2_IR_REG_24__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n5554) );
  XNOR2_X1 U7171 ( .A(n5572), .B(P2_B_REG_SCAN_IN), .ZN(n5559) );
  NAND2_X1 U7172 ( .A1(n5557), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5558) );
  NAND2_X1 U7173 ( .A1(n5559), .A2(n8497), .ZN(n5567) );
  NAND2_X1 U7174 ( .A1(n5561), .A2(n5560), .ZN(n5588) );
  NAND3_X1 U7175 ( .A1(n5563), .A2(n5589), .A3(n5562), .ZN(n5564) );
  OAI21_X1 U7176 ( .B1(n5588), .B2(n5564), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n5565) );
  MUX2_X1 U7177 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5565), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n5566) );
  NAND2_X1 U7178 ( .A1(n8497), .A2(n8496), .ZN(n5568) );
  AOI21_X1 U7179 ( .B1(n5571), .B2(n5570), .A(n8085), .ZN(n5573) );
  OR2_X1 U7180 ( .A1(n5676), .A2(n5573), .ZN(n5576) );
  NAND2_X1 U7181 ( .A1(n5572), .A2(n8496), .ZN(n5984) );
  INV_X1 U7182 ( .A(n5573), .ZN(n5574) );
  INV_X1 U7183 ( .A(n5712), .ZN(n5593) );
  AND2_X1 U7184 ( .A1(n5606), .A2(n5676), .ZN(n5591) );
  NOR2_X1 U7185 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .ZN(
        n5580) );
  NOR4_X1 U7186 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_22__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n5579) );
  NOR4_X1 U7187 ( .A1(P2_D_REG_12__SCAN_IN), .A2(P2_D_REG_25__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_23__SCAN_IN), .ZN(n5578) );
  NOR4_X1 U7188 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_28__SCAN_IN), .A3(
        P2_D_REG_27__SCAN_IN), .A4(P2_D_REG_26__SCAN_IN), .ZN(n5577) );
  NAND4_X1 U7189 ( .A1(n5580), .A2(n5579), .A3(n5578), .A4(n5577), .ZN(n5586)
         );
  NOR4_X1 U7190 ( .A1(P2_D_REG_14__SCAN_IN), .A2(P2_D_REG_13__SCAN_IN), .A3(
        P2_D_REG_21__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n5584) );
  NOR4_X1 U7191 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_9__SCAN_IN), .A3(
        P2_D_REG_17__SCAN_IN), .A4(P2_D_REG_15__SCAN_IN), .ZN(n5583) );
  NOR4_X1 U7192 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n5582) );
  NOR4_X1 U7193 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_19__SCAN_IN), .ZN(n5581) );
  NAND4_X1 U7194 ( .A1(n5584), .A2(n5583), .A3(n5582), .A4(n5581), .ZN(n5585)
         );
  NOR2_X1 U7195 ( .A1(n5586), .A2(n5585), .ZN(n5587) );
  NAND2_X1 U7196 ( .A1(n5588), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5590) );
  NAND2_X1 U7197 ( .A1(n5604), .A2(n8085), .ZN(n5684) );
  NAND3_X1 U7198 ( .A1(n5675), .A2(n5982), .A3(n5684), .ZN(n5710) );
  NOR2_X1 U7199 ( .A1(n5591), .A2(n5710), .ZN(n5592) );
  NAND2_X1 U7200 ( .A1(n5593), .A2(n5592), .ZN(n5597) );
  NAND2_X1 U7201 ( .A1(n5594), .A2(n8115), .ZN(n5596) );
  OAI21_X1 U7202 ( .B1(n5708), .B2(n5595), .A(n10050), .ZN(n5602) );
  NAND2_X1 U7203 ( .A1(n5596), .A2(n10112), .ZN(n10036) );
  NOR2_X1 U7204 ( .A1(n5598), .A2(n10038), .ZN(n8676) );
  NOR2_X1 U7205 ( .A1(n10050), .A2(n5599), .ZN(n5600) );
  AOI211_X1 U7206 ( .C1(n5714), .C2(n8816), .A(n8676), .B(n5600), .ZN(n5601)
         );
  NAND2_X1 U7207 ( .A1(n5602), .A2(n5601), .ZN(P2_U3204) );
  OR2_X1 U7208 ( .A1(n7979), .A2(n8115), .ZN(n8134) );
  AND2_X1 U7209 ( .A1(n5604), .A2(n5603), .ZN(n5605) );
  OAI21_X2 U7210 ( .B1(n5606), .B2(n8134), .A(n5605), .ZN(n5611) );
  XNOR2_X1 U7211 ( .A(n8899), .B(n5628), .ZN(n7817) );
  XNOR2_X1 U7212 ( .A(n7407), .B(n5641), .ZN(n5640) );
  XNOR2_X1 U7213 ( .A(n5611), .B(n6828), .ZN(n5619) );
  INV_X2 U7214 ( .A(n5628), .ZN(n5641) );
  XNOR2_X1 U7215 ( .A(n5611), .B(n6599), .ZN(n5618) );
  INV_X1 U7216 ( .A(n8600), .ZN(n6452) );
  XNOR2_X1 U7217 ( .A(n5611), .B(n10070), .ZN(n5615) );
  INV_X1 U7218 ( .A(n5615), .ZN(n5616) );
  XNOR2_X1 U7219 ( .A(n5611), .B(n10064), .ZN(n5613) );
  INV_X1 U7220 ( .A(n5613), .ZN(n5614) );
  OAI21_X1 U7221 ( .B1(n5611), .B2(n9538), .A(n6516), .ZN(n6133) );
  NAND2_X1 U7222 ( .A1(n6134), .A2(n6133), .ZN(n6132) );
  XNOR2_X1 U7223 ( .A(n5611), .B(n5100), .ZN(n5612) );
  XNOR2_X1 U7224 ( .A(n5612), .B(n5101), .ZN(n6194) );
  INV_X1 U7225 ( .A(n5101), .ZN(n6229) );
  AOI21_X1 U7226 ( .B1(n6193), .B2(n6194), .A(n4873), .ZN(n6227) );
  XNOR2_X1 U7227 ( .A(n5613), .B(n10042), .ZN(n6226) );
  NAND2_X1 U7228 ( .A1(n6227), .A2(n6226), .ZN(n6225) );
  OAI21_X1 U7229 ( .B1(n10042), .B2(n5614), .A(n6225), .ZN(n6283) );
  XNOR2_X1 U7230 ( .A(n5615), .B(n8600), .ZN(n6284) );
  NOR2_X1 U7231 ( .A1(n6283), .A2(n6284), .ZN(n6282) );
  AOI21_X1 U7232 ( .B1(n6452), .B2(n5616), .A(n6282), .ZN(n6449) );
  XNOR2_X1 U7233 ( .A(n5611), .B(n10073), .ZN(n5617) );
  XNOR2_X1 U7234 ( .A(n5617), .B(n8599), .ZN(n6450) );
  OAI22_X1 U7235 ( .A1(n6449), .A2(n6450), .B1(n5617), .B2(n8599), .ZN(n6720)
         );
  XNOR2_X1 U7236 ( .A(n5618), .B(n8598), .ZN(n6721) );
  AOI21_X1 U7237 ( .B1(n5618), .B2(n8598), .A(n6719), .ZN(n6823) );
  XNOR2_X1 U7238 ( .A(n5619), .B(n8597), .ZN(n6822) );
  XNOR2_X1 U7239 ( .A(n5611), .B(n5620), .ZN(n7081) );
  NOR2_X1 U7240 ( .A1(n7081), .A2(n8596), .ZN(n5622) );
  INV_X1 U7241 ( .A(n8596), .ZN(n7106) );
  INV_X1 U7242 ( .A(n7081), .ZN(n5621) );
  XNOR2_X1 U7243 ( .A(n5641), .B(n4480), .ZN(n5623) );
  XNOR2_X1 U7244 ( .A(n5623), .B(n8595), .ZN(n7102) );
  INV_X1 U7245 ( .A(n5623), .ZN(n5624) );
  XNOR2_X1 U7246 ( .A(n7121), .B(n5641), .ZN(n7524) );
  XNOR2_X1 U7247 ( .A(n5641), .B(n7389), .ZN(n7383) );
  NAND2_X1 U7248 ( .A1(n7470), .A2(n5626), .ZN(n5634) );
  INV_X1 U7249 ( .A(n7121), .ZN(n8145) );
  NOR3_X1 U7250 ( .A1(n5628), .A2(n7216), .A3(n8594), .ZN(n5627) );
  AOI211_X1 U7251 ( .C1(n7525), .C2(n5628), .A(n8145), .B(n5627), .ZN(n5631)
         );
  NOR3_X1 U7252 ( .A1(n5641), .A2(n8594), .A3(n7389), .ZN(n5629) );
  AOI211_X1 U7253 ( .C1(n7525), .C2(n5641), .A(n7121), .B(n5629), .ZN(n5630)
         );
  XNOR2_X1 U7254 ( .A(n10113), .B(n5641), .ZN(n5635) );
  XNOR2_X1 U7255 ( .A(n5635), .B(n8592), .ZN(n7526) );
  NAND2_X1 U7256 ( .A1(n5634), .A2(n5633), .ZN(n5637) );
  XNOR2_X1 U7257 ( .A(n7467), .B(n5611), .ZN(n5638) );
  NAND2_X1 U7258 ( .A1(n5638), .A2(n7528), .ZN(n5639) );
  OAI21_X1 U7259 ( .B1(n5638), .B2(n7528), .A(n5639), .ZN(n7460) );
  INV_X1 U7260 ( .A(n5639), .ZN(n7537) );
  XNOR2_X1 U7261 ( .A(n5640), .B(n8590), .ZN(n7536) );
  XNOR2_X1 U7262 ( .A(n7603), .B(n5641), .ZN(n5642) );
  XNOR2_X1 U7263 ( .A(n5642), .B(n7584), .ZN(n7604) );
  INV_X1 U7264 ( .A(n5642), .ZN(n5643) );
  NAND2_X1 U7265 ( .A1(n5643), .A2(n8589), .ZN(n5644) );
  XNOR2_X1 U7266 ( .A(n7679), .B(n5641), .ZN(n5645) );
  XNOR2_X1 U7267 ( .A(n5645), .B(n8588), .ZN(n7671) );
  NAND2_X1 U7268 ( .A1(n7672), .A2(n7671), .ZN(n5648) );
  INV_X1 U7269 ( .A(n5645), .ZN(n5646) );
  NAND2_X1 U7270 ( .A1(n5646), .A2(n8588), .ZN(n5647) );
  XNOR2_X1 U7271 ( .A(n8544), .B(n5641), .ZN(n5649) );
  NAND2_X1 U7272 ( .A1(n5649), .A2(n7674), .ZN(n8567) );
  OAI21_X1 U7273 ( .B1(n5649), .B2(n7674), .A(n8567), .ZN(n8538) );
  XNOR2_X1 U7274 ( .A(n8928), .B(n5641), .ZN(n5651) );
  XNOR2_X1 U7275 ( .A(n5651), .B(n8587), .ZN(n8568) );
  NAND2_X1 U7276 ( .A1(n5650), .A2(n8568), .ZN(n8571) );
  NAND2_X1 U7277 ( .A1(n5651), .A2(n8793), .ZN(n5652) );
  XNOR2_X1 U7278 ( .A(n8852), .B(n5641), .ZN(n5654) );
  XNOR2_X1 U7279 ( .A(n5654), .B(n8576), .ZN(n8505) );
  XNOR2_X1 U7280 ( .A(n8917), .B(n5641), .ZN(n5653) );
  NAND2_X1 U7281 ( .A1(n5653), .A2(n8794), .ZN(n8510) );
  OAI21_X1 U7282 ( .B1(n5653), .B2(n8794), .A(n8510), .ZN(n8550) );
  INV_X1 U7283 ( .A(n5654), .ZN(n5655) );
  AND2_X1 U7284 ( .A1(n5655), .A2(n8810), .ZN(n8551) );
  NOR2_X1 U7285 ( .A1(n8550), .A2(n8551), .ZN(n5656) );
  XNOR2_X1 U7286 ( .A(n8911), .B(n5641), .ZN(n5658) );
  XNOR2_X1 U7287 ( .A(n5658), .B(n8754), .ZN(n8511) );
  NAND2_X1 U7288 ( .A1(n5657), .A2(n8511), .ZN(n8513) );
  XNOR2_X1 U7289 ( .A(n8905), .B(n5641), .ZN(n5660) );
  XNOR2_X1 U7290 ( .A(n5660), .B(n7833), .ZN(n8557) );
  INV_X1 U7291 ( .A(n5660), .ZN(n5661) );
  NAND2_X1 U7292 ( .A1(n5661), .A2(n8768), .ZN(n7816) );
  XNOR2_X1 U7293 ( .A(n7815), .B(n5641), .ZN(n5662) );
  NAND2_X1 U7294 ( .A1(n5662), .A2(n8714), .ZN(n8521) );
  OAI21_X1 U7295 ( .B1(n5662), .B2(n8714), .A(n8521), .ZN(n7820) );
  AOI21_X1 U7296 ( .B1(n7817), .B2(n8753), .A(n7820), .ZN(n5663) );
  XNOR2_X1 U7297 ( .A(n8887), .B(n5641), .ZN(n5665) );
  NAND2_X1 U7298 ( .A1(n5665), .A2(n8732), .ZN(n5670) );
  INV_X1 U7299 ( .A(n5665), .ZN(n5666) );
  NAND2_X1 U7300 ( .A1(n5666), .A2(n8702), .ZN(n5667) );
  NAND2_X1 U7301 ( .A1(n5669), .A2(n8522), .ZN(n8525) );
  XNOR2_X1 U7302 ( .A(n8881), .B(n5641), .ZN(n5870) );
  XNOR2_X1 U7303 ( .A(n5870), .B(n8712), .ZN(n5668) );
  INV_X1 U7304 ( .A(n5668), .ZN(n5671) );
  AND3_X1 U7305 ( .A1(n8525), .A2(n5670), .A3(n5671), .ZN(n5681) );
  AND2_X1 U7306 ( .A1(n8522), .A2(n5668), .ZN(n8474) );
  OR2_X1 U7307 ( .A1(n5671), .A2(n5670), .ZN(n5872) );
  NAND2_X1 U7308 ( .A1(n5877), .A2(n5872), .ZN(n5680) );
  INV_X1 U7309 ( .A(n5675), .ZN(n5672) );
  NOR2_X1 U7310 ( .A1(n5711), .A2(n5672), .ZN(n5689) );
  NAND2_X1 U7311 ( .A1(n5689), .A2(n5982), .ZN(n5722) );
  NOR2_X1 U7312 ( .A1(n8085), .A2(n10112), .ZN(n5674) );
  NAND2_X1 U7313 ( .A1(n5720), .A2(n5674), .ZN(n5683) );
  OR2_X1 U7314 ( .A1(n5722), .A2(n5683), .ZN(n5679) );
  NAND3_X1 U7315 ( .A1(n5606), .A2(n5676), .A3(n5675), .ZN(n5692) );
  INV_X1 U7316 ( .A(n5982), .ZN(n5677) );
  INV_X1 U7317 ( .A(n5720), .ZN(n5686) );
  NAND2_X1 U7318 ( .A1(n5724), .A2(n5686), .ZN(n5678) );
  INV_X1 U7319 ( .A(n8881), .ZN(n5703) );
  OR2_X1 U7320 ( .A1(n5722), .A2(n10103), .ZN(n5682) );
  NAND2_X1 U7321 ( .A1(n5683), .A2(n10036), .ZN(n5723) );
  INV_X1 U7322 ( .A(n5723), .ZN(n5688) );
  NAND2_X1 U7323 ( .A1(n5732), .A2(n5684), .ZN(n5685) );
  AOI21_X1 U7324 ( .B1(n5692), .B2(n5686), .A(n5685), .ZN(n5687) );
  OAI21_X1 U7325 ( .B1(n5689), .B2(n5688), .A(n5687), .ZN(n5690) );
  NAND2_X1 U7326 ( .A1(n5690), .A2(P2_STATE_REG_SCAN_IN), .ZN(n5694) );
  INV_X1 U7327 ( .A(n6275), .ZN(n5691) );
  AND2_X1 U7328 ( .A1(n5982), .A2(n5691), .ZN(n8167) );
  NAND2_X1 U7329 ( .A1(n5692), .A2(n8167), .ZN(n5693) );
  NAND2_X1 U7330 ( .A1(n5694), .A2(n5693), .ZN(n6129) );
  OR2_X1 U7331 ( .A1(n5734), .A2(P2_U3151), .ZN(n8171) );
  INV_X1 U7332 ( .A(n8171), .ZN(n7112) );
  NOR2_X1 U7333 ( .A1(n6275), .A2(n5695), .ZN(n5696) );
  NAND2_X1 U7334 ( .A1(n5724), .A2(n5696), .ZN(n9537) );
  OR2_X1 U7335 ( .A1(n6275), .A2(n5697), .ZN(n5698) );
  AOI22_X1 U7336 ( .A1(n8580), .A2(n8702), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3151), .ZN(n5700) );
  OAI21_X1 U7337 ( .B1(n5873), .B2(n9537), .A(n5700), .ZN(n5701) );
  AOI21_X1 U7338 ( .B1(n8706), .B2(n8563), .A(n5701), .ZN(n5702) );
  OAI21_X1 U7339 ( .B1(n5703), .B2(n8583), .A(n5702), .ZN(n5704) );
  INV_X1 U7340 ( .A(n5704), .ZN(n5705) );
  NAND2_X1 U7341 ( .A1(n5706), .A2(n5705), .ZN(P2_U3180) );
  INV_X1 U7342 ( .A(n10086), .ZN(n10052) );
  NOR2_X1 U7343 ( .A1(n5708), .A2(n4868), .ZN(n5731) );
  NOR2_X1 U7344 ( .A1(n5710), .A2(n5709), .ZN(n5713) );
  INV_X1 U7345 ( .A(n5714), .ZN(n5728) );
  NAND2_X1 U7346 ( .A1(n10135), .A2(n10112), .ZN(n8836) );
  INV_X1 U7347 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n5715) );
  OAI21_X1 U7348 ( .B1(n5731), .B2(n5719), .A(n5718), .ZN(P2_U3488) );
  AND2_X1 U7349 ( .A1(n5720), .A2(n6275), .ZN(n5721) );
  OR2_X1 U7350 ( .A1(n5722), .A2(n5721), .ZN(n5726) );
  NAND2_X1 U7351 ( .A1(n5724), .A2(n5723), .ZN(n5725) );
  INV_X1 U7352 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n5727) );
  OAI21_X1 U7353 ( .B1(n5731), .B2(n10120), .A(n5730), .ZN(P2_U3456) );
  NOR2_X4 U7354 ( .A1(n5732), .A2(n6128), .ZN(P2_U3893) );
  INV_X1 U7355 ( .A(n5732), .ZN(n5733) );
  NAND2_X1 U7356 ( .A1(n5733), .A2(n5734), .ZN(n5858) );
  NAND2_X1 U7357 ( .A1(n8085), .A2(n5734), .ZN(n5735) );
  NAND2_X1 U7358 ( .A1(n5858), .A2(n5735), .ZN(n5852) );
  OR2_X1 U7359 ( .A1(n5852), .A2(n5127), .ZN(n5736) );
  NAND2_X1 U7360 ( .A1(n5736), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3150) );
  INV_X1 U7361 ( .A(n6323), .ZN(n5958) );
  NOR2_X1 U7362 ( .A1(n9948), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n5737) );
  NAND2_X1 U7363 ( .A1(n5094), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5739) );
  OAI21_X1 U7364 ( .B1(n5738), .B2(n5737), .A(n5739), .ZN(n6240) );
  OR2_X1 U7365 ( .A1(n6240), .A2(n5066), .ZN(n6238) );
  NAND2_X1 U7366 ( .A1(n6238), .A2(n5739), .ZN(n9959) );
  XNOR2_X1 U7367 ( .A(n9965), .B(P2_REG2_REG_2__SCAN_IN), .ZN(n9957) );
  NAND2_X1 U7368 ( .A1(n9959), .A2(n9957), .ZN(n9958) );
  INV_X1 U7369 ( .A(n9965), .ZN(n5931) );
  NAND2_X1 U7370 ( .A1(n5931), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n5740) );
  NAND2_X1 U7371 ( .A1(n9958), .A2(n5740), .ZN(n5741) );
  INV_X1 U7372 ( .A(n6302), .ZN(n5932) );
  NAND2_X1 U7373 ( .A1(n5741), .A2(n5932), .ZN(n6329) );
  NAND2_X1 U7374 ( .A1(n6329), .A2(n5742), .ZN(n6295) );
  XNOR2_X1 U7375 ( .A(n6339), .B(P2_REG2_REG_4__SCAN_IN), .ZN(n6330) );
  OR2_X1 U7376 ( .A1(n6339), .A2(n6395), .ZN(n5743) );
  NAND2_X1 U7377 ( .A1(n6332), .A2(n5743), .ZN(n5744) );
  INV_X1 U7378 ( .A(n9984), .ZN(n5944) );
  NAND2_X1 U7379 ( .A1(n5744), .A2(n5944), .ZN(n5745) );
  OAI21_X1 U7380 ( .B1(n5744), .B2(n5944), .A(n5745), .ZN(n9978) );
  MUX2_X1 U7381 ( .A(n5747), .B(P2_REG2_REG_6__SCAN_IN), .S(n10000), .Z(n9991)
         );
  OR2_X1 U7382 ( .A1(n10000), .A2(n5747), .ZN(n5748) );
  NAND2_X1 U7383 ( .A1(n9994), .A2(n5748), .ZN(n5749) );
  NAND2_X1 U7384 ( .A1(n5749), .A2(n5956), .ZN(n6314) );
  INV_X1 U7385 ( .A(n5749), .ZN(n5750) );
  NAND2_X1 U7386 ( .A1(n5750), .A2(n10019), .ZN(n5751) );
  NAND2_X1 U7387 ( .A1(n6314), .A2(n5751), .ZN(n10013) );
  MUX2_X1 U7388 ( .A(n6610), .B(P2_REG2_REG_8__SCAN_IN), .S(n6323), .Z(n6312)
         );
  NOR2_X1 U7389 ( .A1(n5752), .A2(n6372), .ZN(n5755) );
  INV_X1 U7390 ( .A(n5755), .ZN(n5754) );
  NAND2_X1 U7391 ( .A1(n5754), .A2(n5753), .ZN(n6371) );
  NOR2_X1 U7392 ( .A1(n5823), .A2(n6371), .ZN(n6370) );
  NOR2_X1 U7393 ( .A1(n6370), .A2(n5755), .ZN(n6351) );
  AOI22_X1 U7394 ( .A1(n6360), .A2(P2_REG2_REG_10__SCAN_IN), .B1(n7095), .B2(
        n6037), .ZN(n6350) );
  NAND2_X1 U7395 ( .A1(n6037), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n5756) );
  NOR2_X1 U7396 ( .A1(n7058), .A2(n5757), .ZN(n5758) );
  NAND2_X1 U7397 ( .A1(P2_REG2_REG_12__SCAN_IN), .A2(n6099), .ZN(n5759) );
  OAI21_X1 U7398 ( .B1(P2_REG2_REG_12__SCAN_IN), .B2(n6099), .A(n5759), .ZN(
        n6729) );
  NOR2_X1 U7399 ( .A1(n6730), .A2(n6729), .ZN(n6728) );
  NOR2_X1 U7400 ( .A1(n5839), .A2(n5760), .ZN(n5761) );
  NAND2_X1 U7401 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n7320), .ZN(n5762) );
  OAI21_X1 U7402 ( .B1(P2_REG2_REG_14__SCAN_IN), .B2(n7320), .A(n5762), .ZN(
        n7312) );
  INV_X1 U7403 ( .A(n5800), .ZN(n8610) );
  XOR2_X1 U7404 ( .A(n8610), .B(n5763), .Z(n8603) );
  INV_X1 U7405 ( .A(n5798), .ZN(n8629) );
  NAND2_X1 U7406 ( .A1(P2_REG2_REG_16__SCAN_IN), .A2(n8629), .ZN(n5764) );
  OAI21_X1 U7407 ( .B1(P2_REG2_REG_16__SCAN_IN), .B2(n8629), .A(n5764), .ZN(
        n8621) );
  XNOR2_X1 U7408 ( .A(n5765), .B(n5847), .ZN(n8640) );
  NOR2_X1 U7409 ( .A1(n5847), .A2(n5765), .ZN(n5766) );
  INV_X1 U7410 ( .A(n8660), .ZN(n8656) );
  AOI22_X1 U7411 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n8660), .B1(n8656), .B2(
        n8812), .ZN(n5768) );
  OR2_X1 U7412 ( .A1(n5538), .A2(P2_U3151), .ZN(n7310) );
  OR2_X1 U7413 ( .A1(n5852), .A2(n7310), .ZN(n5796) );
  INV_X1 U7414 ( .A(n5796), .ZN(n9952) );
  AOI21_X1 U7415 ( .B1(n4378), .B2(n5769), .A(n10024), .ZN(n5869) );
  AOI22_X1 U7416 ( .A1(P2_REG1_REG_18__SCAN_IN), .A2(n8656), .B1(n8660), .B2(
        n8855), .ZN(n5795) );
  AOI22_X1 U7417 ( .A1(P2_REG1_REG_16__SCAN_IN), .A2(n8629), .B1(n5798), .B2(
        n7590), .ZN(n8625) );
  NAND2_X1 U7418 ( .A1(P2_REG1_REG_14__SCAN_IN), .A2(n7320), .ZN(n5789) );
  AOI22_X1 U7419 ( .A1(P2_REG1_REG_14__SCAN_IN), .A2(n7320), .B1(n5802), .B2(
        n7406), .ZN(n7315) );
  INV_X1 U7420 ( .A(n5839), .ZN(n7188) );
  NAND2_X1 U7421 ( .A1(P2_REG1_REG_12__SCAN_IN), .A2(n6099), .ZN(n5786) );
  AOI22_X1 U7422 ( .A1(P2_REG1_REG_12__SCAN_IN), .A2(n6099), .B1(n6741), .B2(
        n5837), .ZN(n6739) );
  AOI22_X1 U7423 ( .A1(n6360), .A2(n5829), .B1(P2_REG1_REG_10__SCAN_IN), .B2(
        n6037), .ZN(n6358) );
  MUX2_X1 U7424 ( .A(n5775), .B(P2_REG1_REG_2__SCAN_IN), .S(n9965), .Z(n9963)
         );
  NAND2_X1 U7425 ( .A1(n5094), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5773) );
  NAND2_X1 U7426 ( .A1(n5738), .A2(n5773), .ZN(n5772) );
  INV_X1 U7427 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n9955) );
  NAND2_X1 U7428 ( .A1(n9955), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5770) );
  OR2_X1 U7429 ( .A1(n5770), .A2(n5094), .ZN(n5771) );
  NAND2_X1 U7430 ( .A1(n5772), .A2(n5771), .ZN(n6237) );
  NAND2_X1 U7431 ( .A1(n6237), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5774) );
  NAND2_X1 U7432 ( .A1(n5774), .A2(n5773), .ZN(n9962) );
  INV_X1 U7433 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n10126) );
  MUX2_X1 U7434 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n10126), .S(n6339), .Z(n6328)
         );
  OAI22_X1 U7435 ( .A1(n6327), .A2(n6328), .B1(n6339), .B2(n10126), .ZN(n5776)
         );
  NAND2_X1 U7436 ( .A1(n5944), .A2(n5776), .ZN(n5778) );
  XNOR2_X1 U7437 ( .A(n9984), .B(n5776), .ZN(n9976) );
  NAND2_X1 U7438 ( .A1(P2_REG1_REG_5__SCAN_IN), .A2(n9976), .ZN(n5777) );
  NAND2_X1 U7439 ( .A1(n5778), .A2(n5777), .ZN(n9997) );
  INV_X1 U7440 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n5779) );
  MUX2_X1 U7441 ( .A(n5779), .B(P2_REG1_REG_6__SCAN_IN), .S(n10000), .Z(n9996)
         );
  NAND2_X1 U7442 ( .A1(n9997), .A2(n9996), .ZN(n9995) );
  OR2_X1 U7443 ( .A1(n10000), .A2(n5779), .ZN(n5780) );
  AND2_X1 U7444 ( .A1(n9995), .A2(n5780), .ZN(n5781) );
  XNOR2_X1 U7445 ( .A(n5781), .B(n5956), .ZN(n10015) );
  NAND2_X1 U7446 ( .A1(P2_REG1_REG_7__SCAN_IN), .A2(n10015), .ZN(n10014) );
  OAI21_X1 U7447 ( .B1(n5781), .B2(n10019), .A(n10014), .ZN(n6317) );
  MUX2_X1 U7448 ( .A(n5818), .B(P2_REG1_REG_8__SCAN_IN), .S(n6323), .Z(n6318)
         );
  NAND2_X1 U7449 ( .A1(n6317), .A2(n6318), .ZN(n6316) );
  OAI21_X1 U7450 ( .B1(n6323), .B2(n5818), .A(n6316), .ZN(n5782) );
  INV_X1 U7451 ( .A(n6372), .ZN(n6012) );
  NAND2_X1 U7452 ( .A1(n5782), .A2(n6012), .ZN(n5783) );
  XNOR2_X1 U7453 ( .A(n5782), .B(n6372), .ZN(n6369) );
  NAND2_X1 U7454 ( .A1(P2_REG1_REG_9__SCAN_IN), .A2(n6369), .ZN(n6368) );
  NAND2_X1 U7455 ( .A1(n4785), .A2(n5784), .ZN(n5785) );
  NAND2_X1 U7456 ( .A1(P2_REG1_REG_11__SCAN_IN), .A2(n7056), .ZN(n7055) );
  NAND2_X1 U7457 ( .A1(n7188), .A2(n5787), .ZN(n5788) );
  NAND2_X1 U7458 ( .A1(P2_REG1_REG_13__SCAN_IN), .A2(n7184), .ZN(n7183) );
  NAND2_X1 U7459 ( .A1(n8610), .A2(n5790), .ZN(n5791) );
  NAND2_X1 U7460 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n8606), .ZN(n8605) );
  NAND2_X1 U7461 ( .A1(n8646), .A2(n5792), .ZN(n5793) );
  NAND2_X1 U7462 ( .A1(P2_REG1_REG_17__SCAN_IN), .A2(n8642), .ZN(n8641) );
  NAND2_X1 U7463 ( .A1(n5793), .A2(n8641), .ZN(n5794) );
  NAND2_X1 U7464 ( .A1(n5795), .A2(n5794), .ZN(n8658) );
  OAI21_X1 U7465 ( .B1(n5795), .B2(n5794), .A(n8658), .ZN(n5797) );
  NOR2_X2 U7466 ( .A1(n5796), .A2(n8662), .ZN(n10017) );
  NAND2_X1 U7467 ( .A1(P2_U3893), .A2(n5538), .ZN(n8671) );
  MUX2_X1 U7468 ( .A(n7662), .B(n7667), .S(n5537), .Z(n5846) );
  XNOR2_X1 U7469 ( .A(n8646), .B(n5846), .ZN(n8645) );
  MUX2_X1 U7470 ( .A(P2_REG2_REG_16__SCAN_IN), .B(P2_REG1_REG_16__SCAN_IN), 
        .S(n5537), .Z(n5799) );
  OR2_X1 U7471 ( .A1(n5799), .A2(n8629), .ZN(n5844) );
  XNOR2_X1 U7472 ( .A(n5799), .B(n5798), .ZN(n8628) );
  MUX2_X1 U7473 ( .A(P2_REG2_REG_15__SCAN_IN), .B(P2_REG1_REG_15__SCAN_IN), 
        .S(n5537), .Z(n5801) );
  OR2_X1 U7474 ( .A1(n5801), .A2(n8610), .ZN(n5843) );
  XNOR2_X1 U7475 ( .A(n5801), .B(n5800), .ZN(n8609) );
  MUX2_X1 U7476 ( .A(P2_REG2_REG_14__SCAN_IN), .B(P2_REG1_REG_14__SCAN_IN), 
        .S(n5537), .Z(n5803) );
  OR2_X1 U7477 ( .A1(n5803), .A2(n7320), .ZN(n5842) );
  XNOR2_X1 U7478 ( .A(n5803), .B(n5802), .ZN(n7318) );
  MUX2_X1 U7479 ( .A(P2_REG2_REG_13__SCAN_IN), .B(P2_REG1_REG_13__SCAN_IN), 
        .S(n5537), .Z(n5840) );
  OR2_X1 U7480 ( .A1(n5840), .A2(n7188), .ZN(n5841) );
  MUX2_X1 U7481 ( .A(P2_REG2_REG_11__SCAN_IN), .B(P2_REG1_REG_11__SCAN_IN), 
        .S(n5537), .Z(n5835) );
  INV_X1 U7482 ( .A(n5835), .ZN(n5836) );
  MUX2_X1 U7483 ( .A(P2_REG2_REG_6__SCAN_IN), .B(P2_REG1_REG_6__SCAN_IN), .S(
        n5537), .Z(n5812) );
  INV_X1 U7484 ( .A(n10000), .ZN(n5951) );
  MUX2_X1 U7485 ( .A(P2_REG2_REG_4__SCAN_IN), .B(P2_REG1_REG_4__SCAN_IN), .S(
        n5537), .Z(n5809) );
  INV_X1 U7486 ( .A(n5809), .ZN(n5810) );
  INV_X1 U7487 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n10121) );
  MUX2_X1 U7488 ( .A(n5066), .B(n10121), .S(n5537), .Z(n5805) );
  XNOR2_X1 U7489 ( .A(n5805), .B(n6244), .ZN(n6236) );
  MUX2_X1 U7490 ( .A(P2_REG2_REG_0__SCAN_IN), .B(P2_REG1_REG_0__SCAN_IN), .S(
        n5537), .Z(n5804) );
  NOR2_X1 U7491 ( .A1(n5804), .A2(n9955), .ZN(n9951) );
  OAI22_X1 U7492 ( .A1(n6236), .A2(n9951), .B1(n6244), .B2(n5805), .ZN(n9971)
         );
  MUX2_X1 U7493 ( .A(P2_REG2_REG_2__SCAN_IN), .B(P2_REG1_REG_2__SCAN_IN), .S(
        n5537), .Z(n5806) );
  XNOR2_X1 U7494 ( .A(n5806), .B(n9965), .ZN(n9970) );
  AOI22_X1 U7495 ( .A1(n9971), .A2(n9970), .B1(n5806), .B2(n5931), .ZN(n6304)
         );
  MUX2_X1 U7496 ( .A(P2_REG2_REG_3__SCAN_IN), .B(P2_REG1_REG_3__SCAN_IN), .S(
        n5537), .Z(n5807) );
  XNOR2_X1 U7497 ( .A(n5807), .B(n6302), .ZN(n6303) );
  NAND2_X1 U7498 ( .A1(n6304), .A2(n6303), .ZN(n6341) );
  INV_X1 U7499 ( .A(n5807), .ZN(n5808) );
  NAND2_X1 U7500 ( .A1(n5808), .A2(n6302), .ZN(n6340) );
  XNOR2_X1 U7501 ( .A(n5809), .B(n6339), .ZN(n6343) );
  NAND3_X1 U7502 ( .A1(n6341), .A2(n6340), .A3(n6343), .ZN(n6342) );
  OAI21_X1 U7503 ( .B1(n6339), .B2(n5810), .A(n6342), .ZN(n9985) );
  MUX2_X1 U7504 ( .A(P2_REG2_REG_5__SCAN_IN), .B(P2_REG1_REG_5__SCAN_IN), .S(
        n5537), .Z(n5811) );
  XNOR2_X1 U7505 ( .A(n5811), .B(n9984), .ZN(n9986) );
  AOI22_X1 U7506 ( .A1(n9985), .A2(n9986), .B1(n5811), .B2(n5944), .ZN(n10007)
         );
  XNOR2_X1 U7507 ( .A(n5812), .B(n10000), .ZN(n10006) );
  NAND2_X1 U7508 ( .A1(n10007), .A2(n10006), .ZN(n10005) );
  OAI21_X1 U7509 ( .B1(n5812), .B2(n5951), .A(n10005), .ZN(n10027) );
  MUX2_X1 U7510 ( .A(n5814), .B(n5813), .S(n5537), .Z(n5815) );
  NAND2_X1 U7511 ( .A1(n5815), .A2(n10019), .ZN(n6310) );
  INV_X1 U7512 ( .A(n5815), .ZN(n5816) );
  NAND2_X1 U7513 ( .A1(n5816), .A2(n5956), .ZN(n5817) );
  AND2_X1 U7514 ( .A1(n6310), .A2(n5817), .ZN(n10028) );
  NAND2_X1 U7515 ( .A1(n10027), .A2(n10028), .ZN(n10026) );
  MUX2_X1 U7516 ( .A(n6610), .B(n5818), .S(n5537), .Z(n5819) );
  NAND2_X1 U7517 ( .A1(n5819), .A2(n6323), .ZN(n6378) );
  INV_X1 U7518 ( .A(n5819), .ZN(n5820) );
  NAND2_X1 U7519 ( .A1(n5820), .A2(n5958), .ZN(n5821) );
  NAND2_X1 U7520 ( .A1(n6378), .A2(n5821), .ZN(n6309) );
  AOI21_X1 U7521 ( .B1(n10026), .B2(n6310), .A(n6309), .ZN(n6376) );
  INV_X1 U7522 ( .A(n6378), .ZN(n5828) );
  MUX2_X1 U7523 ( .A(n5823), .B(n5822), .S(n5537), .Z(n5824) );
  NAND2_X1 U7524 ( .A1(n5824), .A2(n6372), .ZN(n6353) );
  INV_X1 U7525 ( .A(n5824), .ZN(n5825) );
  NAND2_X1 U7526 ( .A1(n5825), .A2(n6012), .ZN(n5826) );
  NAND2_X1 U7527 ( .A1(n6353), .A2(n5826), .ZN(n6377) );
  INV_X1 U7528 ( .A(n6377), .ZN(n5827) );
  OAI21_X1 U7529 ( .B1(n6376), .B2(n5828), .A(n5827), .ZN(n6381) );
  MUX2_X1 U7530 ( .A(n7095), .B(n5829), .S(n5537), .Z(n5830) );
  NAND2_X1 U7531 ( .A1(n5830), .A2(n6360), .ZN(n5833) );
  INV_X1 U7532 ( .A(n5830), .ZN(n5831) );
  NAND2_X1 U7533 ( .A1(n5831), .A2(n6037), .ZN(n5832) );
  NAND2_X1 U7534 ( .A1(n5833), .A2(n5832), .ZN(n6352) );
  AOI21_X1 U7535 ( .B1(n6381), .B2(n6353), .A(n6352), .ZN(n6355) );
  INV_X1 U7536 ( .A(n5833), .ZN(n5834) );
  NOR2_X1 U7537 ( .A1(n6355), .A2(n5834), .ZN(n7054) );
  XNOR2_X1 U7538 ( .A(n5835), .B(n4785), .ZN(n7053) );
  NOR2_X1 U7539 ( .A1(n7054), .A2(n7053), .ZN(n7052) );
  AOI21_X1 U7540 ( .B1(n7058), .B2(n5836), .A(n7052), .ZN(n6736) );
  MUX2_X1 U7541 ( .A(n7204), .B(n5837), .S(n5537), .Z(n5838) );
  NAND2_X1 U7542 ( .A1(n5838), .A2(n6741), .ZN(n6731) );
  NOR2_X1 U7543 ( .A1(n5838), .A2(n6741), .ZN(n6733) );
  AOI21_X1 U7544 ( .B1(n6736), .B2(n6731), .A(n6733), .ZN(n7186) );
  XNOR2_X1 U7545 ( .A(n5840), .B(n5839), .ZN(n7187) );
  NAND2_X1 U7546 ( .A1(n7186), .A2(n7187), .ZN(n7185) );
  NAND2_X1 U7547 ( .A1(n5841), .A2(n7185), .ZN(n7317) );
  NAND2_X1 U7548 ( .A1(n7318), .A2(n7317), .ZN(n7316) );
  NAND2_X1 U7549 ( .A1(n5842), .A2(n7316), .ZN(n8608) );
  NAND2_X1 U7550 ( .A1(n8609), .A2(n8608), .ZN(n8607) );
  NAND2_X1 U7551 ( .A1(n5843), .A2(n8607), .ZN(n8627) );
  NAND2_X1 U7552 ( .A1(n8628), .A2(n8627), .ZN(n8626) );
  NAND2_X1 U7553 ( .A1(n5844), .A2(n8626), .ZN(n8644) );
  NAND2_X1 U7554 ( .A1(n8645), .A2(n8644), .ZN(n8643) );
  INV_X1 U7555 ( .A(n8643), .ZN(n5845) );
  AOI21_X1 U7556 ( .B1(n5847), .B2(n5846), .A(n5845), .ZN(n5849) );
  MUX2_X1 U7557 ( .A(P2_REG2_REG_18__SCAN_IN), .B(P2_REG1_REG_18__SCAN_IN), 
        .S(n5537), .Z(n5848) );
  NOR2_X1 U7558 ( .A1(n5849), .A2(n5848), .ZN(n8661) );
  NAND2_X1 U7559 ( .A1(n5849), .A2(n5848), .ZN(n8659) );
  INV_X1 U7560 ( .A(n8659), .ZN(n5850) );
  NOR2_X1 U7561 ( .A1(n8661), .A2(n5850), .ZN(n5855) );
  OR2_X1 U7562 ( .A1(n8671), .A2(n5855), .ZN(n5864) );
  NOR2_X1 U7563 ( .A1(n5537), .A2(P2_U3151), .ZN(n7217) );
  NAND2_X1 U7564 ( .A1(n7217), .A2(n5538), .ZN(n5851) );
  OR2_X1 U7565 ( .A1(n5852), .A2(n5851), .ZN(n5854) );
  OR2_X1 U7566 ( .A1(n5858), .A2(n7310), .ZN(n5853) );
  AOI21_X1 U7567 ( .B1(P2_U3893), .B2(n5855), .A(n10020), .ZN(n5856) );
  INV_X1 U7568 ( .A(n5856), .ZN(n5857) );
  INV_X1 U7569 ( .A(n5858), .ZN(n5859) );
  INV_X1 U7570 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n5860) );
  NAND2_X1 U7571 ( .A1(P2_U3151), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8575) );
  OAI21_X1 U7572 ( .B1(n10033), .B2(n5860), .A(n8575), .ZN(n5861) );
  INV_X1 U7573 ( .A(n5865), .ZN(n5866) );
  NAND2_X1 U7574 ( .A1(n5870), .A2(n8529), .ZN(n5871) );
  AND2_X1 U7575 ( .A1(n5872), .A2(n5871), .ZN(n5875) );
  XNOR2_X1 U7576 ( .A(n8875), .B(n5641), .ZN(n8476) );
  XNOR2_X1 U7577 ( .A(n8476), .B(n5873), .ZN(n5874) );
  INV_X1 U7578 ( .A(n5874), .ZN(n5876) );
  NAND2_X1 U7579 ( .A1(n5877), .A2(n8473), .ZN(n5878) );
  INV_X1 U7580 ( .A(n8875), .ZN(n8084) );
  NOR2_X1 U7581 ( .A1(n8530), .A2(n8529), .ZN(n5880) );
  OAI22_X1 U7582 ( .A1(n8095), .A2(n9537), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6976), .ZN(n5879) );
  AOI211_X1 U7583 ( .C1(n8695), .C2(n8563), .A(n5880), .B(n5879), .ZN(n5881)
         );
  INV_X1 U7584 ( .A(n5882), .ZN(n5883) );
  INV_X1 U7585 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n5890) );
  NAND2_X1 U7586 ( .A1(n5884), .A2(n5475), .ZN(n5885) );
  XNOR2_X1 U7587 ( .A(n5885), .B(n8482), .ZN(n5889) );
  INV_X1 U7588 ( .A(n8487), .ZN(n8586) );
  AOI21_X1 U7589 ( .B1(n5889), .B2(n5513), .A(n5888), .ZN(n8867) );
  MUX2_X1 U7590 ( .A(n5890), .B(n8867), .S(n10135), .Z(n5895) );
  XNOR2_X1 U7591 ( .A(n5891), .B(n8482), .ZN(n8872) );
  NAND2_X1 U7592 ( .A1(n8869), .A2(n8856), .ZN(n5892) );
  INV_X1 U7593 ( .A(n5893), .ZN(n5894) );
  NAND2_X1 U7594 ( .A1(n6059), .A2(n5899), .ZN(n5909) );
  NOR2_X1 U7595 ( .A1(n5909), .A2(P1_IR_REG_24__SCAN_IN), .ZN(n5902) );
  NOR2_X1 U7596 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .ZN(
        n5901) );
  NOR2_X1 U7597 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_16__SCAN_IN), .ZN(
        n5900) );
  NAND4_X1 U7598 ( .A1(n5902), .A2(n5915), .A3(n5901), .A4(n5900), .ZN(n5977)
         );
  NAND2_X1 U7599 ( .A1(n5979), .A2(n5903), .ZN(n5919) );
  NAND2_X1 U7600 ( .A1(n5919), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5905) );
  MUX2_X1 U7601 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5905), .S(
        P1_IR_REG_25__SCAN_IN), .Z(n5906) );
  INV_X1 U7602 ( .A(n7306), .ZN(n5907) );
  NAND2_X1 U7603 ( .A1(n5979), .A2(n5908), .ZN(n6056) );
  INV_X1 U7604 ( .A(n5909), .ZN(n5910) );
  NAND2_X1 U7605 ( .A1(n5910), .A2(n6057), .ZN(n5911) );
  NAND2_X1 U7606 ( .A1(n6061), .A2(n5912), .ZN(n5970) );
  INV_X1 U7607 ( .A(n5970), .ZN(n5914) );
  INV_X1 U7608 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5913) );
  NAND2_X1 U7609 ( .A1(n5914), .A2(n5913), .ZN(n5925) );
  INV_X1 U7610 ( .A(n5915), .ZN(n5918) );
  INV_X1 U7611 ( .A(n5919), .ZN(n5921) );
  INV_X1 U7612 ( .A(n6157), .ZN(n6268) );
  NAND2_X1 U7613 ( .A1(n5969), .A2(n5968), .ZN(n5926) );
  NAND2_X1 U7614 ( .A1(n5926), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5928) );
  NAND2_X1 U7615 ( .A1(n5052), .A2(P2_U3151), .ZN(n8470) );
  INV_X1 U7616 ( .A(n6178), .ZN(n5935) );
  INV_X1 U7617 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n5929) );
  NOR2_X1 U7618 ( .A1(n5052), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7628) );
  INV_X1 U7619 ( .A(n7628), .ZN(n8491) );
  OAI222_X1 U7620 ( .A1(n5738), .A2(P2_U3151), .B1(n8470), .B2(n5935), .C1(
        n5929), .C2(n8491), .ZN(P2_U3294) );
  CLKBUF_X1 U7621 ( .A(n8470), .Z(n8494) );
  INV_X1 U7622 ( .A(n5930), .ZN(n6203) );
  OAI222_X1 U7623 ( .A1(n5931), .A2(P2_U3151), .B1(n8494), .B2(n6203), .C1(
        n4938), .C2(n8491), .ZN(P2_U3293) );
  OAI222_X1 U7624 ( .A1(n5932), .A2(P2_U3151), .B1(n8494), .B2(n6248), .C1(
        n4945), .C2(n8491), .ZN(P2_U3292) );
  NAND2_X2 U7625 ( .A1(n5052), .A2(P1_U3086), .ZN(n7913) );
  AND2_X1 U7626 ( .A1(n4962), .A2(P1_U3086), .ZN(n7115) );
  INV_X2 U7627 ( .A(n7115), .ZN(n7915) );
  NAND2_X1 U7628 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(n4368), .ZN(n5933) );
  XNOR2_X1 U7629 ( .A(n5933), .B(P1_IR_REG_2__SCAN_IN), .ZN(n6493) );
  INV_X1 U7630 ( .A(n6493), .ZN(n9599) );
  OAI222_X1 U7631 ( .A1(n7913), .A2(n4734), .B1(n7915), .B2(n6203), .C1(
        P1_U3086), .C2(n9599), .ZN(P1_U3353) );
  OAI21_X1 U7632 ( .B1(P1_IR_REG_2__SCAN_IN), .B2(n4368), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5934) );
  XNOR2_X1 U7633 ( .A(n5934), .B(P1_IR_REG_3__SCAN_IN), .ZN(n6495) );
  INV_X1 U7634 ( .A(n6495), .ZN(n9518) );
  OAI222_X1 U7635 ( .A1(n7913), .A2(n4943), .B1(n7915), .B2(n6248), .C1(
        P1_U3086), .C2(n9518), .ZN(P1_U3352) );
  INV_X1 U7636 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6179) );
  OAI222_X1 U7637 ( .A1(n7913), .A2(n6179), .B1(n7915), .B2(n5935), .C1(
        P1_U3086), .C2(n9585), .ZN(P1_U3354) );
  INV_X1 U7638 ( .A(n5936), .ZN(n6415) );
  AOI22_X1 U7639 ( .A1(n6339), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_4__SCAN_IN), .B2(n7628), .ZN(n5937) );
  OAI21_X1 U7640 ( .B1(n6415), .B2(n8494), .A(n5937), .ZN(P2_U3291) );
  INV_X1 U7641 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6416) );
  OR2_X1 U7642 ( .A1(n5938), .A2(n5973), .ZN(n5940) );
  XNOR2_X1 U7643 ( .A(n5940), .B(P1_IR_REG_4__SCAN_IN), .ZN(n6497) );
  INV_X1 U7644 ( .A(n6497), .ZN(n9620) );
  OAI222_X1 U7645 ( .A1(n7913), .A2(n6416), .B1(n7915), .B2(n6415), .C1(
        P1_U3086), .C2(n9620), .ZN(P1_U3351) );
  INV_X1 U7646 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n5939) );
  NAND2_X1 U7647 ( .A1(n5940), .A2(n5939), .ZN(n5941) );
  NAND2_X1 U7648 ( .A1(n5941), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5942) );
  XNOR2_X1 U7649 ( .A(n5942), .B(P1_IR_REG_5__SCAN_IN), .ZN(n6499) );
  INV_X1 U7650 ( .A(n6499), .ZN(n9635) );
  OAI222_X1 U7651 ( .A1(n7913), .A2(n6526), .B1(n7915), .B2(n6525), .C1(
        P1_U3086), .C2(n9635), .ZN(P1_U3350) );
  OAI222_X1 U7652 ( .A1(n5944), .A2(P2_U3151), .B1(n8494), .B2(n6525), .C1(
        n5943), .C2(n8491), .ZN(P2_U3290) );
  INV_X1 U7653 ( .A(n6569), .ZN(n5950) );
  NAND2_X1 U7654 ( .A1(n5945), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5946) );
  MUX2_X1 U7655 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5946), .S(
        P1_IR_REG_6__SCAN_IN), .Z(n5947) );
  INV_X1 U7656 ( .A(n6568), .ZN(n9651) );
  OAI222_X1 U7657 ( .A1(n7915), .A2(n5950), .B1(n9651), .B2(P1_U3086), .C1(
        n5948), .C2(n7913), .ZN(P1_U3349) );
  OAI222_X1 U7658 ( .A1(P2_U3151), .A2(n5951), .B1(n8470), .B2(n5950), .C1(
        n5949), .C2(n8491), .ZN(P2_U3289) );
  INV_X1 U7659 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n5953) );
  INV_X1 U7660 ( .A(n6648), .ZN(n5955) );
  NAND2_X1 U7661 ( .A1(n5959), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5952) );
  XNOR2_X1 U7662 ( .A(n5952), .B(P1_IR_REG_7__SCAN_IN), .ZN(n6649) );
  INV_X1 U7663 ( .A(n6649), .ZN(n9503) );
  OAI222_X1 U7664 ( .A1(n7913), .A2(n5953), .B1(n7915), .B2(n5955), .C1(
        P1_U3086), .C2(n9503), .ZN(P1_U3348) );
  INV_X1 U7665 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n5954) );
  OAI222_X1 U7666 ( .A1(n5956), .A2(P2_U3151), .B1(n8470), .B2(n5955), .C1(
        n5954), .C2(n8491), .ZN(P2_U3288) );
  INV_X1 U7667 ( .A(n6652), .ZN(n5964) );
  OAI222_X1 U7668 ( .A1(n5958), .A2(P2_U3151), .B1(n8470), .B2(n5964), .C1(
        n5957), .C2(n8491), .ZN(P2_U3287) );
  NOR2_X1 U7669 ( .A1(n5959), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n6014) );
  OR2_X1 U7670 ( .A1(n6014), .A2(n5973), .ZN(n5962) );
  INV_X1 U7671 ( .A(n5962), .ZN(n5960) );
  NAND2_X1 U7672 ( .A1(n5960), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n5963) );
  INV_X1 U7673 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n5961) );
  NAND2_X1 U7674 ( .A1(n5962), .A2(n5961), .ZN(n5987) );
  INV_X1 U7675 ( .A(n6653), .ZN(n9532) );
  OAI222_X1 U7676 ( .A1(n7913), .A2(n5965), .B1(n7915), .B2(n5964), .C1(
        P1_U3086), .C2(n9532), .ZN(P1_U3347) );
  INV_X1 U7677 ( .A(n5972), .ZN(n5967) );
  NAND2_X1 U7678 ( .A1(n5967), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8466) );
  NAND2_X1 U7679 ( .A1(n6171), .A2(n8466), .ZN(n6483) );
  NAND2_X1 U7680 ( .A1(n5970), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5971) );
  NAND2_X1 U7681 ( .A1(n8353), .A2(n5972), .ZN(n5980) );
  INV_X1 U7682 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n5973) );
  NAND2_X1 U7683 ( .A1(n5975), .A2(n5974), .ZN(n5976) );
  NAND2_X1 U7684 ( .A1(n5979), .A2(n5978), .ZN(n5997) );
  AND2_X1 U7685 ( .A1(n5980), .A2(n8173), .ZN(n6482) );
  INV_X1 U7686 ( .A(n6482), .ZN(n5981) );
  NOR2_X1 U7687 ( .A1(n9609), .A2(P1_U3973), .ZN(P1_U3085) );
  INV_X1 U7688 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n5986) );
  INV_X1 U7689 ( .A(n5984), .ZN(n5985) );
  AOI22_X1 U7690 ( .A1(n8500), .A2(n5986), .B1(n8495), .B2(n5985), .ZN(
        P2_U3376) );
  INV_X1 U7691 ( .A(n6693), .ZN(n6011) );
  NAND2_X1 U7692 ( .A1(n5987), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5988) );
  XNOR2_X1 U7693 ( .A(n5988), .B(P1_IR_REG_9__SCAN_IN), .ZN(n9091) );
  INV_X1 U7694 ( .A(n7913), .ZN(n7624) );
  AOI22_X1 U7695 ( .A1(n9091), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n7624), .ZN(n5989) );
  OAI21_X1 U7696 ( .B1(n6011), .B2(n7915), .A(n5989), .ZN(P1_U3346) );
  INV_X1 U7697 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n6009) );
  NAND2_X1 U7698 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_28__SCAN_IN), 
        .ZN(n5990) );
  NAND2_X1 U7699 ( .A1(n4878), .A2(P1_IR_REG_30__SCAN_IN), .ZN(n5994) );
  NAND3_X1 U7700 ( .A1(n5995), .A2(n5999), .A3(n5992), .ZN(n5996) );
  NAND2_X2 U7701 ( .A1(n5998), .A2(n7622), .ZN(n7601) );
  XNOR2_X2 U7702 ( .A(n6000), .B(n5999), .ZN(n6003) );
  INV_X1 U7703 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n6007) );
  NAND2_X4 U7704 ( .A1(n6001), .A2(n7601), .ZN(n8177) );
  INV_X1 U7705 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n6002) );
  OR2_X1 U7706 ( .A1(n8177), .A2(n6002), .ZN(n6006) );
  NAND2_X4 U7707 ( .A1(n7601), .A2(n7599), .ZN(n8179) );
  INV_X1 U7708 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n6004) );
  OR2_X1 U7709 ( .A1(n8179), .A2(n6004), .ZN(n6005) );
  OAI211_X1 U7710 ( .C1(n7941), .C2(n6007), .A(n6006), .B(n6005), .ZN(n9163)
         );
  NAND2_X1 U7711 ( .A1(n9163), .A2(P1_U3973), .ZN(n6008) );
  OAI21_X1 U7712 ( .B1(P1_U3973), .B2(n6009), .A(n6008), .ZN(P1_U3585) );
  OAI222_X1 U7713 ( .A1(P2_U3151), .A2(n6012), .B1(n8470), .B2(n6011), .C1(
        n6010), .C2(n8491), .ZN(P2_U3286) );
  INV_X1 U7714 ( .A(n6773), .ZN(n6036) );
  NOR2_X1 U7715 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n6013) );
  AND2_X1 U7716 ( .A1(n6014), .A2(n6013), .ZN(n6018) );
  NOR2_X1 U7717 ( .A1(n6018), .A2(n5973), .ZN(n6015) );
  MUX2_X1 U7718 ( .A(n5973), .B(n6015), .S(P1_IR_REG_10__SCAN_IN), .Z(n6016)
         );
  INV_X1 U7719 ( .A(n6016), .ZN(n6019) );
  INV_X1 U7720 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n6017) );
  NAND2_X1 U7721 ( .A1(n6018), .A2(n6017), .ZN(n6090) );
  AOI22_X1 U7722 ( .A1(n9489), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n7624), .ZN(n6020) );
  OAI21_X1 U7723 ( .B1(n6036), .B2(n7915), .A(n6020), .ZN(P1_U3345) );
  INV_X1 U7724 ( .A(P2_D_REG_11__SCAN_IN), .ZN(n6021) );
  NOR2_X1 U7725 ( .A1(n6105), .A2(n6021), .ZN(P2_U3254) );
  INV_X1 U7726 ( .A(P2_D_REG_17__SCAN_IN), .ZN(n6022) );
  NOR2_X1 U7727 ( .A1(n6105), .A2(n6022), .ZN(P2_U3248) );
  INV_X1 U7728 ( .A(P2_D_REG_12__SCAN_IN), .ZN(n6023) );
  NOR2_X1 U7729 ( .A1(n6105), .A2(n6023), .ZN(P2_U3253) );
  INV_X1 U7730 ( .A(P2_D_REG_19__SCAN_IN), .ZN(n6024) );
  NOR2_X1 U7731 ( .A1(n6105), .A2(n6024), .ZN(P2_U3246) );
  INV_X1 U7732 ( .A(P2_D_REG_13__SCAN_IN), .ZN(n6025) );
  NOR2_X1 U7733 ( .A1(n6105), .A2(n6025), .ZN(P2_U3252) );
  INV_X1 U7734 ( .A(P2_D_REG_15__SCAN_IN), .ZN(n6026) );
  NOR2_X1 U7735 ( .A1(n6105), .A2(n6026), .ZN(P2_U3250) );
  INV_X1 U7736 ( .A(P2_D_REG_16__SCAN_IN), .ZN(n6027) );
  NOR2_X1 U7737 ( .A1(n6105), .A2(n6027), .ZN(P2_U3249) );
  INV_X1 U7738 ( .A(P2_D_REG_14__SCAN_IN), .ZN(n6028) );
  NOR2_X1 U7739 ( .A1(n6105), .A2(n6028), .ZN(P2_U3251) );
  INV_X1 U7740 ( .A(P2_D_REG_18__SCAN_IN), .ZN(n6029) );
  NOR2_X1 U7741 ( .A1(n6105), .A2(n6029), .ZN(P2_U3247) );
  INV_X1 U7742 ( .A(P2_D_REG_25__SCAN_IN), .ZN(n6030) );
  NOR2_X1 U7743 ( .A1(n6105), .A2(n6030), .ZN(P2_U3240) );
  INV_X1 U7744 ( .A(P2_D_REG_23__SCAN_IN), .ZN(n6031) );
  NOR2_X1 U7745 ( .A1(n6105), .A2(n6031), .ZN(P2_U3242) );
  INV_X1 U7746 ( .A(P2_D_REG_21__SCAN_IN), .ZN(n6032) );
  NOR2_X1 U7747 ( .A1(n6105), .A2(n6032), .ZN(P2_U3244) );
  INV_X1 U7748 ( .A(P2_D_REG_24__SCAN_IN), .ZN(n6033) );
  NOR2_X1 U7749 ( .A1(n6105), .A2(n6033), .ZN(P2_U3241) );
  INV_X1 U7750 ( .A(P2_D_REG_20__SCAN_IN), .ZN(n6034) );
  NOR2_X1 U7751 ( .A1(n6105), .A2(n6034), .ZN(P2_U3245) );
  INV_X1 U7752 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6035) );
  OAI222_X1 U7753 ( .A1(P2_U3151), .A2(n6037), .B1(n8470), .B2(n6036), .C1(
        n6035), .C2(n8491), .ZN(P2_U3285) );
  INV_X1 U7754 ( .A(n7144), .ZN(n6041) );
  NAND2_X1 U7755 ( .A1(n6090), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6038) );
  XNOR2_X1 U7756 ( .A(n6038), .B(P1_IR_REG_11__SCAN_IN), .ZN(n9656) );
  AOI22_X1 U7757 ( .A1(n9656), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n7624), .ZN(n6039) );
  OAI21_X1 U7758 ( .B1(n6041), .B2(n7915), .A(n6039), .ZN(P1_U3344) );
  INV_X1 U7759 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6040) );
  OAI222_X1 U7760 ( .A1(n4785), .A2(P2_U3151), .B1(n8470), .B2(n6041), .C1(
        n6040), .C2(n8491), .ZN(P2_U3284) );
  NAND2_X1 U7761 ( .A1(n7306), .A2(P1_B_REG_SCAN_IN), .ZN(n6044) );
  INV_X1 U7762 ( .A(P1_B_REG_SCAN_IN), .ZN(n9160) );
  NAND2_X1 U7763 ( .A1(n6042), .A2(n9160), .ZN(n6043) );
  INV_X1 U7764 ( .A(n6045), .ZN(n7307) );
  NAND2_X1 U7765 ( .A1(n7307), .A2(n7306), .ZN(n9477) );
  OAI21_X1 U7766 ( .B1(n9475), .B2(P1_D_REG_1__SCAN_IN), .A(n9477), .ZN(n6147)
         );
  NOR4_X1 U7767 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n6054) );
  NOR4_X1 U7768 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n6053) );
  NOR4_X1 U7769 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n6049) );
  NOR4_X1 U7770 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_17__SCAN_IN), .ZN(n6048) );
  NOR4_X1 U7771 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n6047) );
  NOR4_X1 U7772 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n6046) );
  NAND4_X1 U7773 ( .A1(n6049), .A2(n6048), .A3(n6047), .A4(n6046), .ZN(n6050)
         );
  NOR4_X1 U7774 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        n6051), .A4(n6050), .ZN(n6052) );
  AND3_X1 U7775 ( .A1(n6054), .A2(n6053), .A3(n6052), .ZN(n6055) );
  OR2_X1 U7776 ( .A1(n9475), .A2(n6055), .ZN(n6145) );
  NAND2_X1 U7777 ( .A1(n6056), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6387) );
  NAND2_X1 U7778 ( .A1(n6387), .A2(n6057), .ZN(n6058) );
  NAND2_X1 U7779 ( .A1(n6058), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6410) );
  NAND2_X1 U7780 ( .A1(n6410), .A2(n6059), .ZN(n6413) );
  NAND2_X1 U7781 ( .A1(n6413), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6060) );
  INV_X1 U7782 ( .A(n6061), .ZN(n6062) );
  NAND2_X1 U7783 ( .A1(n9903), .A2(n8405), .ZN(n6170) );
  INV_X1 U7784 ( .A(n6042), .ZN(n7219) );
  NAND2_X1 U7785 ( .A1(n7219), .A2(n7307), .ZN(n9478) );
  OAI21_X1 U7786 ( .B1(n9475), .B2(P1_D_REG_0__SCAN_IN), .A(n9478), .ZN(n9382)
         );
  INV_X1 U7787 ( .A(n9381), .ZN(n6065) );
  INV_X1 U7788 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n6089) );
  NAND2_X1 U7789 ( .A1(n6075), .A2(n8405), .ZN(n6627) );
  INV_X1 U7790 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n9570) );
  INV_X1 U7791 ( .A(SI_0_), .ZN(n6067) );
  INV_X1 U7792 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n6066) );
  OAI21_X1 U7793 ( .B1(n5052), .B2(n6067), .A(n6066), .ZN(n6069) );
  NAND2_X1 U7794 ( .A1(n6069), .A2(n6068), .ZN(n9479) );
  OR2_X1 U7795 ( .A1(n6070), .A2(n6075), .ZN(n6071) );
  NAND2_X1 U7796 ( .A1(n6151), .A2(n6064), .ZN(n8175) );
  INV_X1 U7797 ( .A(n6166), .ZN(n6072) );
  NAND2_X1 U7798 ( .A1(n8353), .A2(n6072), .ZN(n6073) );
  AND2_X1 U7799 ( .A1(n6073), .A2(n6627), .ZN(n6553) );
  NAND2_X1 U7800 ( .A1(n6155), .A2(n6166), .ZN(n6076) );
  NAND2_X1 U7801 ( .A1(n6553), .A2(n6076), .ZN(n9817) );
  INV_X1 U7802 ( .A(n9903), .ZN(n9921) );
  OR2_X4 U7803 ( .A1(n7601), .A2(n7599), .ZN(n6262) );
  NAND2_X1 U7804 ( .A1(n7282), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n6080) );
  NAND2_X1 U7805 ( .A1(n7731), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n6079) );
  OR2_X1 U7806 ( .A1(n8179), .A2(n6089), .ZN(n6078) );
  INV_X1 U7807 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n6490) );
  OR2_X1 U7808 ( .A1(n8177), .A2(n6490), .ZN(n6077) );
  INV_X1 U7809 ( .A(n9813), .ZN(n6081) );
  NAND2_X1 U7810 ( .A1(n9081), .A2(n9830), .ZN(n8406) );
  NAND2_X1 U7811 ( .A1(n6081), .A2(n8406), .ZN(n8357) );
  OAI21_X1 U7812 ( .B1(n9821), .B2(n9914), .A(n8357), .ZN(n6087) );
  INV_X1 U7813 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n6489) );
  INV_X1 U7814 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n6082) );
  OAI22_X1 U7815 ( .A1(n8177), .A2(n6489), .B1(n8179), .B2(n6082), .ZN(n6086)
         );
  INV_X1 U7816 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n6084) );
  INV_X1 U7817 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n6083) );
  OR2_X2 U7818 ( .A1(n6086), .A2(n6085), .ZN(n6616) );
  NAND2_X1 U7819 ( .A1(n8353), .A2(n9567), .ZN(n9162) );
  NAND2_X1 U7820 ( .A1(n6616), .A2(n9052), .ZN(n6550) );
  OAI211_X1 U7821 ( .C1(n6627), .C2(n9830), .A(n6087), .B(n6550), .ZN(n9459)
         );
  NAND2_X1 U7822 ( .A1(n9459), .A2(n9927), .ZN(n6088) );
  OAI21_X1 U7823 ( .B1(n9927), .B2(n6089), .A(n6088), .ZN(P1_U3453) );
  INV_X1 U7824 ( .A(n7149), .ZN(n6098) );
  NAND2_X1 U7825 ( .A1(n6091), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6094) );
  INV_X1 U7826 ( .A(n6094), .ZN(n6092) );
  NAND2_X1 U7827 ( .A1(n6092), .A2(P1_IR_REG_12__SCAN_IN), .ZN(n6095) );
  INV_X1 U7828 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n6093) );
  NAND2_X1 U7829 ( .A1(n6094), .A2(n6093), .ZN(n6100) );
  INV_X1 U7830 ( .A(n9098), .ZN(n6505) );
  OAI222_X1 U7831 ( .A1(n7915), .A2(n6098), .B1(n6505), .B2(P1_U3086), .C1(
        n6096), .C2(n7913), .ZN(P1_U3343) );
  OAI222_X1 U7832 ( .A1(P2_U3151), .A2(n6099), .B1(n8470), .B2(n6098), .C1(
        n6097), .C2(n8491), .ZN(P2_U3283) );
  INV_X1 U7833 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n6102) );
  INV_X1 U7834 ( .A(n7254), .ZN(n6104) );
  NAND2_X1 U7835 ( .A1(n6100), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6101) );
  XNOR2_X1 U7836 ( .A(n6101), .B(P1_IR_REG_13__SCAN_IN), .ZN(n9680) );
  INV_X1 U7837 ( .A(n9680), .ZN(n9108) );
  OAI222_X1 U7838 ( .A1(n7913), .A2(n6102), .B1(n7915), .B2(n6104), .C1(
        P1_U3086), .C2(n9108), .ZN(P1_U3342) );
  INV_X1 U7839 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6103) );
  OAI222_X1 U7840 ( .A1(n7188), .A2(P2_U3151), .B1(n8470), .B2(n6104), .C1(
        n6103), .C2(n8491), .ZN(P2_U3282) );
  INV_X1 U7841 ( .A(P2_D_REG_3__SCAN_IN), .ZN(n6106) );
  NOR2_X1 U7842 ( .A1(n6105), .A2(n6106), .ZN(P2_U3262) );
  INV_X1 U7843 ( .A(P2_D_REG_22__SCAN_IN), .ZN(n6107) );
  NOR2_X1 U7844 ( .A1(n6105), .A2(n6107), .ZN(P2_U3243) );
  INV_X1 U7845 ( .A(P2_D_REG_2__SCAN_IN), .ZN(n6108) );
  NOR2_X1 U7846 ( .A1(n6105), .A2(n6108), .ZN(P2_U3263) );
  INV_X1 U7847 ( .A(P2_D_REG_6__SCAN_IN), .ZN(n6109) );
  NOR2_X1 U7848 ( .A1(n6105), .A2(n6109), .ZN(P2_U3259) );
  INV_X1 U7849 ( .A(P2_D_REG_31__SCAN_IN), .ZN(n6110) );
  NOR2_X1 U7850 ( .A1(n6105), .A2(n6110), .ZN(P2_U3234) );
  INV_X1 U7851 ( .A(P2_D_REG_29__SCAN_IN), .ZN(n6111) );
  NOR2_X1 U7852 ( .A1(n6105), .A2(n6111), .ZN(P2_U3236) );
  INV_X1 U7853 ( .A(P2_D_REG_4__SCAN_IN), .ZN(n6112) );
  NOR2_X1 U7854 ( .A1(n6105), .A2(n6112), .ZN(P2_U3261) );
  INV_X1 U7855 ( .A(P2_D_REG_28__SCAN_IN), .ZN(n6113) );
  NOR2_X1 U7856 ( .A1(n6105), .A2(n6113), .ZN(P2_U3237) );
  INV_X1 U7857 ( .A(P2_D_REG_5__SCAN_IN), .ZN(n6114) );
  NOR2_X1 U7858 ( .A1(n6105), .A2(n6114), .ZN(P2_U3260) );
  INV_X1 U7859 ( .A(P2_D_REG_27__SCAN_IN), .ZN(n6115) );
  NOR2_X1 U7860 ( .A1(n6105), .A2(n6115), .ZN(P2_U3238) );
  INV_X1 U7861 ( .A(P2_D_REG_9__SCAN_IN), .ZN(n6116) );
  NOR2_X1 U7862 ( .A1(n6105), .A2(n6116), .ZN(P2_U3256) );
  INV_X1 U7863 ( .A(P2_D_REG_7__SCAN_IN), .ZN(n6117) );
  NOR2_X1 U7864 ( .A1(n6105), .A2(n6117), .ZN(P2_U3258) );
  INV_X1 U7865 ( .A(P2_D_REG_30__SCAN_IN), .ZN(n6118) );
  NOR2_X1 U7866 ( .A1(n6105), .A2(n6118), .ZN(P2_U3235) );
  INV_X1 U7867 ( .A(P2_D_REG_10__SCAN_IN), .ZN(n6119) );
  NOR2_X1 U7868 ( .A1(n6105), .A2(n6119), .ZN(P2_U3255) );
  INV_X1 U7869 ( .A(P2_D_REG_26__SCAN_IN), .ZN(n6120) );
  NOR2_X1 U7870 ( .A1(n6105), .A2(n6120), .ZN(P2_U3239) );
  INV_X1 U7871 ( .A(P2_D_REG_8__SCAN_IN), .ZN(n6121) );
  NOR2_X1 U7872 ( .A1(n6105), .A2(n6121), .ZN(P2_U3257) );
  INV_X1 U7873 ( .A(n7257), .ZN(n6140) );
  OR2_X1 U7874 ( .A1(n6123), .A2(n5973), .ZN(n6125) );
  MUX2_X1 U7875 ( .A(n6125), .B(P1_IR_REG_31__SCAN_IN), .S(n6124), .Z(n6126)
         );
  AND2_X1 U7876 ( .A1(n6122), .A2(n6126), .ZN(n9113) );
  AOI22_X1 U7877 ( .A1(n9113), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n7624), .ZN(n6127) );
  OAI21_X1 U7878 ( .B1(n6140), .B2(n7915), .A(n6127), .ZN(P1_U3341) );
  NOR2_X1 U7879 ( .A1(n6129), .A2(n6128), .ZN(n9546) );
  OAI22_X1 U7880 ( .A1(n8530), .A2(n4350), .B1(n6229), .B2(n9537), .ZN(n6131)
         );
  AOI21_X1 U7881 ( .B1(n6518), .B2(n9539), .A(n6131), .ZN(n6137) );
  OAI21_X1 U7882 ( .B1(n6134), .B2(n6133), .A(n6132), .ZN(n6135) );
  NAND2_X1 U7883 ( .A1(n6135), .A2(n8572), .ZN(n6136) );
  OAI211_X1 U7884 ( .C1(n9546), .C2(n6138), .A(n6137), .B(n6136), .ZN(P2_U3162) );
  INV_X1 U7885 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6139) );
  OAI222_X1 U7886 ( .A1(n7320), .A2(P2_U3151), .B1(n8494), .B2(n6140), .C1(
        n6139), .C2(n8491), .ZN(P2_U3281) );
  AND2_X1 U7887 ( .A1(n6130), .A2(n6141), .ZN(n7982) );
  INV_X1 U7888 ( .A(n7982), .ZN(n7978) );
  AND2_X1 U7889 ( .A1(n6516), .A2(n7978), .ZN(n9542) );
  NOR2_X1 U7890 ( .A1(n10110), .A2(n5513), .ZN(n6143) );
  NAND2_X1 U7891 ( .A1(n9538), .A2(n10112), .ZN(n6142) );
  NAND2_X1 U7892 ( .A1(n5607), .A2(n8809), .ZN(n6276) );
  OAI211_X1 U7893 ( .C1(n9542), .C2(n6143), .A(n6142), .B(n6276), .ZN(n8860)
         );
  NAND2_X1 U7894 ( .A1(n10118), .A2(n8860), .ZN(n6144) );
  OAI21_X1 U7895 ( .B1(n10118), .B2(n4582), .A(n6144), .ZN(P2_U3390) );
  INV_X1 U7896 ( .A(n6145), .ZN(n6146) );
  NOR2_X1 U7897 ( .A1(n6147), .A2(n6146), .ZN(n6546) );
  INV_X1 U7898 ( .A(n9382), .ZN(n6148) );
  NAND2_X1 U7899 ( .A1(n6546), .A2(n6148), .ZN(n6169) );
  INV_X1 U7900 ( .A(n6171), .ZN(n9476) );
  INV_X1 U7901 ( .A(n8353), .ZN(n6149) );
  INV_X1 U7902 ( .A(n6627), .ZN(n6549) );
  NAND3_X1 U7903 ( .A1(n9476), .A2(n6149), .A3(n9911), .ZN(n6150) );
  NAND2_X2 U7904 ( .A1(n6157), .A2(n6153), .ZN(n6158) );
  INV_X1 U7905 ( .A(n9081), .ZN(n6154) );
  OAI222_X1 U7906 ( .A1(n7948), .A2(n9830), .B1(n6158), .B2(n6154), .C1(n6157), 
        .C2(n9570), .ZN(n6162) );
  NAND3_X4 U7907 ( .A1(n6157), .A2(n6156), .A3(n6155), .ZN(n7949) );
  INV_X1 U7908 ( .A(n9830), .ZN(n6623) );
  NAND2_X1 U7909 ( .A1(n6252), .A2(n6623), .ZN(n6160) );
  AND2_X1 U7910 ( .A1(n6160), .A2(n6159), .ZN(n6175) );
  NAND2_X1 U7911 ( .A1(n6175), .A2(n4874), .ZN(n6161) );
  OAI21_X1 U7912 ( .B1(n6162), .B2(n6161), .A(n6177), .ZN(n9601) );
  NAND2_X1 U7913 ( .A1(n6169), .A2(n6170), .ZN(n6165) );
  INV_X1 U7914 ( .A(n6163), .ZN(n6164) );
  NAND2_X1 U7915 ( .A1(n6165), .A2(n6164), .ZN(n6269) );
  NOR2_X1 U7916 ( .A1(n6269), .A2(n6171), .ZN(n8996) );
  INV_X1 U7917 ( .A(n8996), .ZN(n6221) );
  INV_X1 U7918 ( .A(n6169), .ZN(n6167) );
  NOR2_X1 U7919 ( .A1(n6171), .A2(n6166), .ZN(n8462) );
  OR2_X1 U7920 ( .A1(n6627), .A2(n6749), .ZN(n6548) );
  OR2_X1 U7921 ( .A1(n6171), .A2(n6548), .ZN(n6168) );
  OR2_X1 U7922 ( .A1(n6169), .A2(n6168), .ZN(n6172) );
  OAI22_X1 U7923 ( .A1(n9056), .A2(n6550), .B1(n9061), .B2(n9830), .ZN(n6173)
         );
  AOI21_X1 U7924 ( .B1(P1_REG3_REG_0__SCAN_IN), .B2(n6221), .A(n6173), .ZN(
        n6174) );
  OAI21_X1 U7925 ( .B1(n9036), .B2(n9601), .A(n6174), .ZN(P1_U3232) );
  INV_X1 U7926 ( .A(n6175), .ZN(n6176) );
  NAND2_X1 U7927 ( .A1(n6177), .A2(n4866), .ZN(n6213) );
  NAND2_X1 U7928 ( .A1(n4346), .A2(n6615), .ZN(n6183) );
  NAND2_X1 U7929 ( .A1(n6616), .A2(n7709), .ZN(n6182) );
  NAND2_X1 U7930 ( .A1(n6183), .A2(n6182), .ZN(n6184) );
  INV_X1 U7931 ( .A(n6616), .ZN(n6624) );
  OAI22_X1 U7932 ( .A1(n6624), .A2(n6158), .B1(n6626), .B2(n7948), .ZN(n6211)
         );
  XNOR2_X1 U7933 ( .A(n6210), .B(n6211), .ZN(n6212) );
  XOR2_X1 U7934 ( .A(n6213), .B(n6212), .Z(n6192) );
  INV_X1 U7935 ( .A(n9567), .ZN(n9603) );
  NAND2_X1 U7936 ( .A1(n7282), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n6189) );
  NAND2_X1 U7937 ( .A1(n7731), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6188) );
  INV_X1 U7938 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n6185) );
  OR2_X1 U7939 ( .A1(n8179), .A2(n6185), .ZN(n6187) );
  INV_X1 U7940 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n6492) );
  OR2_X1 U7941 ( .A1(n8177), .A2(n6492), .ZN(n6186) );
  AOI22_X1 U7942 ( .A1(n9225), .A2(n9081), .B1(n9080), .B2(n9052), .ZN(n9814)
         );
  OAI22_X1 U7943 ( .A1(n9814), .A2(n9056), .B1(n9061), .B2(n6626), .ZN(n6190)
         );
  AOI21_X1 U7944 ( .B1(P1_REG3_REG_1__SCAN_IN), .B2(n6221), .A(n6190), .ZN(
        n6191) );
  OAI21_X1 U7945 ( .B1(n6192), .B2(n9036), .A(n6191), .ZN(P1_U3222) );
  XOR2_X1 U7946 ( .A(n6194), .B(n6193), .Z(n6198) );
  OAI22_X1 U7947 ( .A1(n8530), .A2(n5609), .B1(n10042), .B2(n9537), .ZN(n6196)
         );
  NOR2_X1 U7948 ( .A1(n9546), .A2(n10037), .ZN(n6195) );
  AOI211_X1 U7949 ( .C1(n5100), .C2(n9539), .A(n6196), .B(n6195), .ZN(n6197)
         );
  OAI21_X1 U7950 ( .B1(n9543), .B2(n6198), .A(n6197), .ZN(P2_U3177) );
  INV_X1 U7951 ( .A(n7423), .ZN(n6235) );
  NAND2_X1 U7952 ( .A1(n6122), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6199) );
  MUX2_X1 U7953 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6199), .S(
        P1_IR_REG_15__SCAN_IN), .Z(n6201) );
  NAND2_X1 U7954 ( .A1(n6201), .A2(n6200), .ZN(n9115) );
  INV_X1 U7955 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n6202) );
  OAI222_X1 U7956 ( .A1(n7915), .A2(n6235), .B1(n9115), .B2(P1_U3086), .C1(
        n6202), .C2(n7913), .ZN(P1_U3340) );
  NAND2_X1 U7957 ( .A1(n9080), .A2(n7709), .ZN(n6208) );
  OR2_X1 U7958 ( .A1(n7636), .A2(n6203), .ZN(n6206) );
  OR2_X1 U7959 ( .A1(n8173), .A2(n9599), .ZN(n6205) );
  NAND2_X1 U7960 ( .A1(n6208), .A2(n6207), .ZN(n6209) );
  XNOR2_X1 U7961 ( .A(n6209), .B(n7949), .ZN(n6256) );
  AOI22_X1 U7962 ( .A1(n9080), .A2(n7924), .B1(n6614), .B2(n7709), .ZN(n6257)
         );
  XNOR2_X1 U7963 ( .A(n6256), .B(n6257), .ZN(n6259) );
  OAI22_X1 U7964 ( .A1(n6213), .A2(n6212), .B1(n6211), .B2(n6210), .ZN(n6260)
         );
  XOR2_X1 U7965 ( .A(n6259), .B(n6260), .Z(n6224) );
  NAND2_X1 U7966 ( .A1(n6616), .A2(n9225), .ZN(n6220) );
  INV_X1 U7967 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n6271) );
  NAND2_X1 U7968 ( .A1(n7282), .A2(n6271), .ZN(n6218) );
  NAND2_X1 U7969 ( .A1(n7731), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6217) );
  INV_X1 U7970 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n6214) );
  OR2_X1 U7971 ( .A1(n8179), .A2(n6214), .ZN(n6216) );
  INV_X1 U7972 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6494) );
  OR2_X1 U7973 ( .A1(n8177), .A2(n6494), .ZN(n6215) );
  NAND2_X1 U7974 ( .A1(n9079), .A2(n9052), .ZN(n6219) );
  NAND2_X1 U7975 ( .A1(n6220), .A2(n6219), .ZN(n6618) );
  AOI22_X1 U7976 ( .A1(n9018), .A2(n6618), .B1(n9023), .B2(n6614), .ZN(n6223)
         );
  NAND2_X1 U7977 ( .A1(n6221), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n6222) );
  OAI211_X1 U7978 ( .C1(n6224), .C2(n9036), .A(n6223), .B(n6222), .ZN(P1_U3237) );
  OAI211_X1 U7979 ( .C1(n6227), .C2(n6226), .A(n6225), .B(n8572), .ZN(n6233)
         );
  NOR2_X1 U7980 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n4884), .ZN(n6301) );
  AOI21_X1 U7981 ( .B1(n8547), .B2(n8600), .A(n6301), .ZN(n6228) );
  OAI21_X1 U7982 ( .B1(n6229), .B2(n8530), .A(n6228), .ZN(n6230) );
  AOI21_X1 U7983 ( .B1(n6231), .B2(n9539), .A(n6230), .ZN(n6232) );
  OAI211_X1 U7984 ( .C1(P2_REG3_REG_3__SCAN_IN), .C2(n8577), .A(n6233), .B(
        n6232), .ZN(P2_U3158) );
  INV_X1 U7985 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n6234) );
  OAI222_X1 U7986 ( .A1(P2_U3151), .A2(n8610), .B1(n8494), .B2(n6235), .C1(
        n6234), .C2(n8491), .ZN(P2_U3280) );
  XNOR2_X1 U7987 ( .A(n6236), .B(n9951), .ZN(n6247) );
  INV_X1 U7988 ( .A(n10017), .ZN(n9981) );
  XOR2_X1 U7989 ( .A(P2_REG1_REG_1__SCAN_IN), .B(n6237), .Z(n6242) );
  INV_X1 U7990 ( .A(n6238), .ZN(n6239) );
  AOI21_X1 U7991 ( .B1(n5066), .B2(n6240), .A(n6239), .ZN(n6241) );
  OAI22_X1 U7992 ( .A1(n9981), .A2(n6242), .B1(n6241), .B2(n10024), .ZN(n6243)
         );
  AOI21_X1 U7993 ( .B1(n9946), .B2(P2_ADDR_REG_1__SCAN_IN), .A(n6243), .ZN(
        n6246) );
  AOI22_X1 U7994 ( .A1(n10020), .A2(n6244), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        P2_U3151), .ZN(n6245) );
  OAI211_X1 U7995 ( .C1(n6247), .C2(n8671), .A(n6246), .B(n6245), .ZN(P2_U3183) );
  OR2_X1 U7996 ( .A1(n7636), .A2(n6248), .ZN(n6251) );
  OR2_X1 U7997 ( .A1(n4347), .A2(n4943), .ZN(n6250) );
  OR2_X1 U7998 ( .A1(n8173), .A2(n9518), .ZN(n6249) );
  INV_X1 U7999 ( .A(n9849), .ZN(n6686) );
  AOI22_X1 U8000 ( .A1(n9079), .A2(n7924), .B1(n6686), .B2(n7709), .ZN(n6438)
         );
  NAND2_X1 U8001 ( .A1(n9079), .A2(n7709), .ZN(n6254) );
  NAND2_X1 U8002 ( .A1(n6686), .A2(n6252), .ZN(n6253) );
  NAND2_X1 U8003 ( .A1(n6254), .A2(n6253), .ZN(n6255) );
  XOR2_X1 U8004 ( .A(n6438), .B(n6440), .Z(n6441) );
  INV_X1 U8005 ( .A(n6256), .ZN(n6258) );
  XOR2_X1 U8006 ( .A(n6441), .B(n6442), .Z(n6274) );
  INV_X1 U8007 ( .A(n9080), .ZN(n6267) );
  INV_X1 U8008 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6815) );
  INV_X1 U8009 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n6496) );
  OR2_X1 U8010 ( .A1(n8177), .A2(n6496), .ZN(n6261) );
  OAI21_X1 U8011 ( .B1(n7941), .B2(n6815), .A(n6261), .ZN(n6266) );
  NAND2_X1 U8012 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n6422) );
  OAI21_X1 U8013 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(n6422), .ZN(n6814) );
  INV_X1 U8014 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n6263) );
  OR2_X1 U8015 ( .A1(n8179), .A2(n6263), .ZN(n6264) );
  OAI21_X1 U8016 ( .B1(n6262), .B2(n6814), .A(n6264), .ZN(n6265) );
  OAI22_X1 U8017 ( .A1(n6267), .A2(n9017), .B1(n6639), .B2(n9162), .ZN(n9797)
         );
  AOI22_X1 U8018 ( .A1(n9018), .A2(n9797), .B1(n9023), .B2(n6686), .ZN(n6273)
         );
  OAI21_X1 U8019 ( .B1(n6269), .B2(n6268), .A(P1_STATE_REG_SCAN_IN), .ZN(n6270) );
  MUX2_X1 U8020 ( .A(P1_STATE_REG_SCAN_IN), .B(n9021), .S(n6271), .Z(n6272) );
  OAI211_X1 U8021 ( .C1(n6274), .C2(n9036), .A(n6273), .B(n6272), .ZN(P1_U3218) );
  NAND2_X1 U8022 ( .A1(n6275), .A2(n10103), .ZN(n6278) );
  NAND2_X1 U8023 ( .A1(n8815), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n6277) );
  OAI211_X1 U8024 ( .C1(n9542), .C2(n6278), .A(n6277), .B(n6276), .ZN(n6279)
         );
  MUX2_X1 U8025 ( .A(n6279), .B(P2_REG2_REG_0__SCAN_IN), .S(n8797), .Z(n6280)
         );
  AOI21_X1 U8026 ( .B1(n8816), .B2(n9538), .A(n6280), .ZN(n6281) );
  INV_X1 U8027 ( .A(n6281), .ZN(P2_U3233) );
  AOI21_X1 U8028 ( .B1(n6284), .B2(n6283), .A(n6282), .ZN(n6289) );
  AND2_X1 U8029 ( .A1(P2_U3151), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n6338) );
  AOI21_X1 U8030 ( .B1(n8547), .B2(n8599), .A(n6338), .ZN(n6285) );
  OAI21_X1 U8031 ( .B1(n10042), .B2(n8530), .A(n6285), .ZN(n6287) );
  NOR2_X1 U8032 ( .A1(n8577), .A2(n6396), .ZN(n6286) );
  AOI211_X1 U8033 ( .C1(n6398), .C2(n9539), .A(n6287), .B(n6286), .ZN(n6288)
         );
  OAI21_X1 U8034 ( .B1(n6289), .B2(n9543), .A(n6288), .ZN(P2_U3170) );
  INV_X1 U8035 ( .A(n7430), .ZN(n6292) );
  INV_X1 U8036 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n6290) );
  OAI222_X1 U8037 ( .A1(n8629), .A2(P2_U3151), .B1(n8494), .B2(n6292), .C1(
        n6290), .C2(n8491), .ZN(P2_U3279) );
  INV_X1 U8038 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n6293) );
  NAND2_X1 U8039 ( .A1(n6200), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6291) );
  XNOR2_X1 U8040 ( .A(n6291), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9128) );
  INV_X1 U8041 ( .A(n9128), .ZN(n9107) );
  OAI222_X1 U8042 ( .A1(n7913), .A2(n6293), .B1(n7915), .B2(n6292), .C1(
        P1_U3086), .C2(n9107), .ZN(P1_U3339) );
  INV_X1 U8043 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n6308) );
  XOR2_X1 U8044 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n6294), .Z(n6299) );
  INV_X1 U8045 ( .A(n6296), .ZN(n6297) );
  AOI21_X1 U8046 ( .B1(n5105), .B2(n6295), .A(n6297), .ZN(n6298) );
  OAI22_X1 U8047 ( .A1(n9981), .A2(n6299), .B1(n6298), .B2(n10024), .ZN(n6300)
         );
  AOI211_X1 U8048 ( .C1(n6302), .C2(n10020), .A(n6301), .B(n6300), .ZN(n6307)
         );
  OAI21_X1 U8049 ( .B1(n6304), .B2(n6303), .A(n6341), .ZN(n6305) );
  NAND2_X1 U8050 ( .A1(n6305), .A2(n10029), .ZN(n6306) );
  OAI211_X1 U8051 ( .C1(n6308), .C2(n10033), .A(n6307), .B(n6306), .ZN(
        P2_U3185) );
  INV_X1 U8052 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n6326) );
  AND3_X1 U8053 ( .A1(n10026), .A2(n6310), .A3(n6309), .ZN(n6311) );
  OAI21_X1 U8054 ( .B1(n6376), .B2(n6311), .A(n10029), .ZN(n6325) );
  NOR2_X1 U8055 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n4441), .ZN(n7084) );
  NOR2_X1 U8056 ( .A1(n6312), .A2(n10012), .ZN(n6315) );
  AOI21_X1 U8057 ( .B1(n6315), .B2(n6314), .A(n6313), .ZN(n6321) );
  OAI21_X1 U8058 ( .B1(n6318), .B2(n6317), .A(n6316), .ZN(n6319) );
  NAND2_X1 U8059 ( .A1(n10017), .A2(n6319), .ZN(n6320) );
  OAI21_X1 U8060 ( .B1(n6321), .B2(n10024), .A(n6320), .ZN(n6322) );
  AOI211_X1 U8061 ( .C1(n6323), .C2(n10020), .A(n7084), .B(n6322), .ZN(n6324)
         );
  OAI211_X1 U8062 ( .C1(n6326), .C2(n10033), .A(n6325), .B(n6324), .ZN(
        P2_U3190) );
  INV_X1 U8063 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n6347) );
  XOR2_X1 U8064 ( .A(n6328), .B(n6327), .Z(n6336) );
  INV_X1 U8065 ( .A(n6329), .ZN(n6331) );
  NOR2_X1 U8066 ( .A1(n6331), .A2(n6330), .ZN(n6334) );
  INV_X1 U8067 ( .A(n6332), .ZN(n6333) );
  AOI21_X1 U8068 ( .B1(n6334), .B2(n6296), .A(n6333), .ZN(n6335) );
  OAI22_X1 U8069 ( .A1(n9981), .A2(n6336), .B1(n6335), .B2(n10024), .ZN(n6337)
         );
  AOI211_X1 U8070 ( .C1(n6339), .C2(n10020), .A(n6338), .B(n6337), .ZN(n6346)
         );
  AND2_X1 U8071 ( .A1(n6341), .A2(n6340), .ZN(n6344) );
  OAI211_X1 U8072 ( .C1(n6344), .C2(n6343), .A(n10029), .B(n6342), .ZN(n6345)
         );
  OAI211_X1 U8073 ( .C1(n6347), .C2(n10033), .A(n6346), .B(n6345), .ZN(
        P2_U3186) );
  AOI21_X1 U8074 ( .B1(n6351), .B2(n6350), .A(n6349), .ZN(n6367) );
  AND3_X1 U8075 ( .A1(n6381), .A2(n6353), .A3(n6352), .ZN(n6354) );
  OAI21_X1 U8076 ( .B1(n6355), .B2(n6354), .A(n10029), .ZN(n6366) );
  OAI21_X1 U8077 ( .B1(n6358), .B2(n6357), .A(n6356), .ZN(n6364) );
  INV_X1 U8078 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n6362) );
  INV_X1 U8079 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n6359) );
  NOR2_X1 U8080 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6359), .ZN(n7386) );
  AOI21_X1 U8081 ( .B1(n10020), .B2(n6360), .A(n7386), .ZN(n6361) );
  OAI21_X1 U8082 ( .B1(n10033), .B2(n6362), .A(n6361), .ZN(n6363) );
  AOI21_X1 U8083 ( .B1(n6364), .B2(n10017), .A(n6363), .ZN(n6365) );
  OAI211_X1 U8084 ( .C1(n6367), .C2(n10024), .A(n6366), .B(n6365), .ZN(
        P2_U3192) );
  OAI21_X1 U8085 ( .B1(n6369), .B2(P2_REG1_REG_9__SCAN_IN), .A(n6368), .ZN(
        n6384) );
  AOI21_X1 U8086 ( .B1(n6371), .B2(n5823), .A(n6370), .ZN(n6375) );
  NAND2_X1 U8087 ( .A1(n9946), .A2(P2_ADDR_REG_9__SCAN_IN), .ZN(n6374) );
  NOR2_X1 U8088 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n4889), .ZN(n7104) );
  AOI21_X1 U8089 ( .B1(n10020), .B2(n6372), .A(n7104), .ZN(n6373) );
  OAI211_X1 U8090 ( .C1(n6375), .C2(n10024), .A(n6374), .B(n6373), .ZN(n6383)
         );
  INV_X1 U8091 ( .A(n6376), .ZN(n6379) );
  NAND3_X1 U8092 ( .A1(n6379), .A2(n6378), .A3(n6377), .ZN(n6380) );
  AOI21_X1 U8093 ( .B1(n6381), .B2(n6380), .A(n8671), .ZN(n6382) );
  AOI211_X1 U8094 ( .C1(n10017), .C2(n6384), .A(n6383), .B(n6382), .ZN(n6385)
         );
  INV_X1 U8095 ( .A(n6385), .ZN(P2_U3191) );
  INV_X1 U8096 ( .A(n7485), .ZN(n6388) );
  INV_X1 U8097 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n6386) );
  OAI222_X1 U8098 ( .A1(P2_U3151), .A2(n8646), .B1(n8494), .B2(n6388), .C1(
        n6386), .C2(n8491), .ZN(P2_U3278) );
  INV_X1 U8099 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n6389) );
  XNOR2_X1 U8100 ( .A(n6387), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9140) );
  INV_X1 U8101 ( .A(n9140), .ZN(n9130) );
  OAI222_X1 U8102 ( .A1(n7913), .A2(n6389), .B1(n9130), .B2(P1_U3086), .C1(
        n7915), .C2(n6388), .ZN(P1_U3338) );
  NOR2_X1 U8103 ( .A1(n10079), .A2(n4426), .ZN(n6390) );
  XNOR2_X1 U8104 ( .A(n6391), .B(n5133), .ZN(n10068) );
  OAI21_X1 U8105 ( .B1(n6393), .B2(n5133), .A(n6392), .ZN(n6394) );
  AOI222_X1 U8106 ( .A1(n5513), .A2(n6394), .B1(n8601), .B2(n8807), .C1(n8599), 
        .C2(n8809), .ZN(n10069) );
  MUX2_X1 U8107 ( .A(n6395), .B(n10069), .S(n10050), .Z(n6400) );
  INV_X1 U8108 ( .A(n6396), .ZN(n6397) );
  AOI22_X1 U8109 ( .A1(n8816), .A2(n6398), .B1(n8815), .B2(n6397), .ZN(n6399)
         );
  OAI211_X1 U8110 ( .C1(n8819), .C2(n10068), .A(n6400), .B(n6399), .ZN(
        P2_U3229) );
  INV_X1 U8111 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n6401) );
  OAI222_X1 U8112 ( .A1(P2_U3151), .A2(n8656), .B1(n8494), .B2(n7637), .C1(
        n6401), .C2(n8491), .ZN(P2_U3277) );
  OR2_X1 U8113 ( .A1(n6402), .A2(n4367), .ZN(n6403) );
  XOR2_X1 U8114 ( .A(n6404), .B(n4367), .Z(n6405) );
  AOI222_X1 U8115 ( .A1(n5513), .A2(n6405), .B1(n8598), .B2(n8809), .C1(n8600), 
        .C2(n8807), .ZN(n10075) );
  MUX2_X1 U8116 ( .A(n6406), .B(n10075), .S(n10050), .Z(n6409) );
  INV_X1 U8117 ( .A(n6453), .ZN(n6407) );
  AOI22_X1 U8118 ( .A1(n8816), .A2(n6456), .B1(n8815), .B2(n6407), .ZN(n6408)
         );
  OAI211_X1 U8119 ( .C1(n10074), .C2(n8819), .A(n6409), .B(n6408), .ZN(
        P2_U3228) );
  INV_X1 U8120 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n6414) );
  INV_X1 U8121 ( .A(n6410), .ZN(n6411) );
  NAND2_X1 U8122 ( .A1(n6411), .A2(P1_IR_REG_18__SCAN_IN), .ZN(n6412) );
  AND2_X1 U8123 ( .A1(n6413), .A2(n6412), .ZN(n9144) );
  INV_X1 U8124 ( .A(n9144), .ZN(n9723) );
  OAI222_X1 U8125 ( .A1(n7913), .A2(n6414), .B1(n9723), .B2(P1_U3086), .C1(
        n7915), .C2(n7637), .ZN(P1_U3337) );
  INV_X1 U8126 ( .A(n6814), .ZN(n6447) );
  INV_X1 U8127 ( .A(n9021), .ZN(n9058) );
  OR2_X1 U8128 ( .A1(n7636), .A2(n6415), .ZN(n6418) );
  OR2_X1 U8129 ( .A1(n4347), .A2(n6416), .ZN(n6417) );
  NAND2_X1 U8130 ( .A1(n9079), .A2(n9225), .ZN(n6429) );
  INV_X1 U8131 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n6421) );
  INV_X1 U8132 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n6419) );
  OR2_X1 U8133 ( .A1(n8177), .A2(n6419), .ZN(n6420) );
  OAI21_X1 U8134 ( .B1(n7941), .B2(n6421), .A(n6420), .ZN(n6427) );
  AND2_X1 U8135 ( .A1(n6422), .A2(n6540), .ZN(n6423) );
  NOR2_X1 U8136 ( .A1(n6422), .A2(n6540), .ZN(n6535) );
  OR2_X1 U8137 ( .A1(n6423), .A2(n6535), .ZN(n9785) );
  INV_X1 U8138 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n6424) );
  OR2_X1 U8139 ( .A1(n8179), .A2(n6424), .ZN(n6425) );
  OAI21_X1 U8140 ( .B1(n6262), .B2(n9785), .A(n6425), .ZN(n6426) );
  NAND2_X1 U8141 ( .A1(n9077), .A2(n9052), .ZN(n6428) );
  NAND2_X1 U8142 ( .A1(n6429), .A2(n6428), .ZN(n6809) );
  AOI22_X1 U8143 ( .A1(n9018), .A2(n6809), .B1(P1_REG3_REG_4__SCAN_IN), .B2(
        P1_U3086), .ZN(n6430) );
  OAI21_X1 U8144 ( .B1(n9855), .B2(n9061), .A(n6430), .ZN(n6446) );
  NAND2_X1 U8145 ( .A1(n9078), .A2(n7709), .ZN(n6432) );
  NAND2_X1 U8146 ( .A1(n6817), .A2(n4346), .ZN(n6431) );
  NAND2_X1 U8147 ( .A1(n6432), .A2(n6431), .ZN(n6433) );
  XNOR2_X1 U8148 ( .A(n6433), .B(n7949), .ZN(n6437) );
  NAND2_X1 U8149 ( .A1(n9078), .A2(n7924), .ZN(n6435) );
  NAND2_X1 U8150 ( .A1(n6817), .A2(n7709), .ZN(n6434) );
  NAND2_X1 U8151 ( .A1(n6435), .A2(n6434), .ZN(n6436) );
  NAND2_X1 U8152 ( .A1(n6437), .A2(n6436), .ZN(n6522) );
  OAI21_X1 U8153 ( .B1(n6437), .B2(n6436), .A(n6522), .ZN(n6444) );
  INV_X1 U8154 ( .A(n6438), .ZN(n6439) );
  AOI211_X1 U8155 ( .C1(n6444), .C2(n6443), .A(n9036), .B(n6524), .ZN(n6445)
         );
  AOI211_X1 U8156 ( .C1(n6447), .C2(n9058), .A(n6446), .B(n6445), .ZN(n6448)
         );
  INV_X1 U8157 ( .A(n6448), .ZN(P1_U3230) );
  XOR2_X1 U8158 ( .A(n6450), .B(n6449), .Z(n6458) );
  AND2_X1 U8159 ( .A1(P2_U3151), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n9983) );
  AOI21_X1 U8160 ( .B1(n8547), .B2(n8598), .A(n9983), .ZN(n6451) );
  OAI21_X1 U8161 ( .B1(n6452), .B2(n8530), .A(n6451), .ZN(n6455) );
  NOR2_X1 U8162 ( .A1(n8577), .A2(n6453), .ZN(n6454) );
  AOI211_X1 U8163 ( .C1(n6456), .C2(n9539), .A(n6455), .B(n6454), .ZN(n6457)
         );
  OAI21_X1 U8164 ( .B1(n6458), .B2(n9543), .A(n6457), .ZN(P2_U3167) );
  OR2_X1 U8165 ( .A1(n6461), .A2(n6460), .ZN(n6462) );
  NAND2_X1 U8166 ( .A1(n6459), .A2(n6462), .ZN(n10087) );
  INV_X1 U8167 ( .A(n10087), .ZN(n6467) );
  INV_X1 U8168 ( .A(n10079), .ZN(n10047) );
  XNOR2_X1 U8169 ( .A(n6463), .B(n8139), .ZN(n6464) );
  NAND2_X1 U8170 ( .A1(n6464), .A2(n5513), .ZN(n6466) );
  AOI22_X1 U8171 ( .A1(n8807), .A2(n8598), .B1(n8596), .B2(n8809), .ZN(n6465)
         );
  OAI211_X1 U8172 ( .C1(n10087), .C2(n10047), .A(n6466), .B(n6465), .ZN(n10089) );
  AOI21_X1 U8173 ( .B1(n4426), .B2(n6467), .A(n10089), .ZN(n6470) );
  OAI22_X1 U8174 ( .A1(n8681), .A2(n10085), .B1(n6831), .B2(n10038), .ZN(n6468) );
  AOI21_X1 U8175 ( .B1(n8797), .B2(P2_REG2_REG_7__SCAN_IN), .A(n6468), .ZN(
        n6469) );
  OAI21_X1 U8176 ( .B1(n6470), .B2(n8797), .A(n6469), .ZN(P2_U3226) );
  NOR2_X1 U8177 ( .A1(n9098), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n9109) );
  AOI21_X1 U8178 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(n9098), .A(n9109), .ZN(
        n6481) );
  NAND2_X1 U8179 ( .A1(n9489), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6471) );
  OAI21_X1 U8180 ( .B1(n9489), .B2(P1_REG2_REG_10__SCAN_IN), .A(n6471), .ZN(
        n9485) );
  INV_X1 U8181 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n9568) );
  NOR2_X1 U8182 ( .A1(n9570), .A2(n9568), .ZN(n9602) );
  INV_X1 U8183 ( .A(n9602), .ZN(n9580) );
  AOI21_X1 U8184 ( .B1(P1_REG2_REG_1__SCAN_IN), .B2(n6491), .A(n9579), .ZN(
        n9595) );
  INV_X1 U8185 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n6629) );
  AOI22_X1 U8186 ( .A1(n6493), .A2(n6629), .B1(P1_REG2_REG_2__SCAN_IN), .B2(
        n9599), .ZN(n9594) );
  INV_X1 U8187 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n6472) );
  AOI22_X1 U8188 ( .A1(n6495), .A2(n6472), .B1(P1_REG2_REG_3__SCAN_IN), .B2(
        n9518), .ZN(n9514) );
  AOI22_X1 U8189 ( .A1(n6497), .A2(n6815), .B1(P1_REG2_REG_4__SCAN_IN), .B2(
        n9620), .ZN(n9616) );
  NOR2_X1 U8190 ( .A1(n9615), .A2(n9616), .ZN(n9614) );
  NAND2_X1 U8191 ( .A1(n6499), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n6473) );
  OAI21_X1 U8192 ( .B1(n6499), .B2(P1_REG2_REG_5__SCAN_IN), .A(n6473), .ZN(
        n9627) );
  NAND2_X1 U8193 ( .A1(n6568), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6474) );
  OAI21_X1 U8194 ( .B1(n6568), .B2(P1_REG2_REG_6__SCAN_IN), .A(n6474), .ZN(
        n9647) );
  AOI21_X1 U8195 ( .B1(P1_REG2_REG_6__SCAN_IN), .B2(n6568), .A(n9645), .ZN(
        n9498) );
  INV_X1 U8196 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n6475) );
  AOI22_X1 U8197 ( .A1(n6649), .A2(n6475), .B1(P1_REG2_REG_7__SCAN_IN), .B2(
        n9503), .ZN(n9499) );
  NOR2_X1 U8198 ( .A1(n9498), .A2(n9499), .ZN(n9497) );
  NAND2_X1 U8199 ( .A1(n6653), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6476) );
  OAI21_X1 U8200 ( .B1(n6653), .B2(P1_REG2_REG_8__SCAN_IN), .A(n6476), .ZN(
        n9525) );
  NOR2_X1 U8201 ( .A1(n9524), .A2(n9525), .ZN(n9523) );
  NOR2_X1 U8202 ( .A1(n9091), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6477) );
  AOI21_X1 U8203 ( .B1(P1_REG2_REG_9__SCAN_IN), .B2(n9091), .A(n6477), .ZN(
        n9084) );
  NAND2_X1 U8204 ( .A1(n9656), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6479) );
  OAI21_X1 U8205 ( .B1(n9656), .B2(P1_REG2_REG_11__SCAN_IN), .A(n6479), .ZN(
        n9663) );
  NOR2_X1 U8206 ( .A1(n9662), .A2(n9663), .ZN(n9661) );
  OAI21_X1 U8207 ( .B1(n6481), .B2(n6480), .A(n9111), .ZN(n6486) );
  NAND2_X1 U8208 ( .A1(n6483), .A2(n6482), .ZN(n9573) );
  OR2_X1 U8209 ( .A1(n9567), .A2(n6484), .ZN(n6485) );
  NAND2_X1 U8210 ( .A1(n6486), .A2(n9718), .ZN(n6509) );
  NAND2_X1 U8211 ( .A1(n9489), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n6487) );
  OAI21_X1 U8212 ( .B1(n9489), .B2(P1_REG1_REG_10__SCAN_IN), .A(n6487), .ZN(
        n9482) );
  NOR2_X1 U8213 ( .A1(n9091), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6488) );
  AOI21_X1 U8214 ( .B1(P1_REG1_REG_9__SCAN_IN), .B2(n9091), .A(n6488), .ZN(
        n9089) );
  MUX2_X1 U8215 ( .A(n6492), .B(P1_REG1_REG_2__SCAN_IN), .S(n6493), .Z(n9591)
         );
  MUX2_X1 U8216 ( .A(n6494), .B(P1_REG1_REG_3__SCAN_IN), .S(n6495), .Z(n9510)
         );
  MUX2_X1 U8217 ( .A(n6496), .B(P1_REG1_REG_4__SCAN_IN), .S(n6497), .Z(n9612)
         );
  NOR2_X1 U8218 ( .A1(n9611), .A2(n9612), .ZN(n9610) );
  AOI21_X1 U8219 ( .B1(n6497), .B2(P1_REG1_REG_4__SCAN_IN), .A(n9610), .ZN(
        n9630) );
  NAND2_X1 U8220 ( .A1(n6499), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6498) );
  OAI21_X1 U8221 ( .B1(n6499), .B2(P1_REG1_REG_5__SCAN_IN), .A(n6498), .ZN(
        n9631) );
  NOR2_X1 U8222 ( .A1(n9630), .A2(n9631), .ZN(n9629) );
  AOI21_X1 U8223 ( .B1(n6499), .B2(P1_REG1_REG_5__SCAN_IN), .A(n9629), .ZN(
        n9643) );
  NAND2_X1 U8224 ( .A1(n6568), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6500) );
  OAI21_X1 U8225 ( .B1(n6568), .B2(P1_REG1_REG_6__SCAN_IN), .A(n6500), .ZN(
        n9642) );
  INV_X1 U8226 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n6578) );
  MUX2_X1 U8227 ( .A(n6578), .B(P1_REG1_REG_7__SCAN_IN), .S(n6649), .Z(n9495)
         );
  NAND2_X1 U8228 ( .A1(n6653), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6501) );
  OAI21_X1 U8229 ( .B1(n6653), .B2(P1_REG1_REG_8__SCAN_IN), .A(n6501), .ZN(
        n9528) );
  NOR2_X1 U8230 ( .A1(n4379), .A2(n9528), .ZN(n9527) );
  AOI21_X1 U8231 ( .B1(P1_REG1_REG_8__SCAN_IN), .B2(n6653), .A(n9527), .ZN(
        n9088) );
  NAND2_X1 U8232 ( .A1(n9089), .A2(n9088), .ZN(n9087) );
  OAI21_X1 U8233 ( .B1(n9091), .B2(P1_REG1_REG_9__SCAN_IN), .A(n9087), .ZN(
        n9483) );
  NOR2_X1 U8234 ( .A1(n9482), .A2(n9483), .ZN(n9481) );
  INV_X1 U8235 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n6783) );
  MUX2_X1 U8236 ( .A(n6783), .B(P1_REG1_REG_11__SCAN_IN), .S(n9656), .Z(n9659)
         );
  INV_X1 U8237 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n9940) );
  AOI22_X1 U8238 ( .A1(n9098), .A2(P1_REG1_REG_12__SCAN_IN), .B1(n9940), .B2(
        n6505), .ZN(n6502) );
  OAI21_X1 U8239 ( .B1(n6503), .B2(n6502), .A(n9097), .ZN(n6507) );
  INV_X1 U8240 ( .A(n6484), .ZN(n9569) );
  NAND2_X1 U8241 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n7248) );
  NAND2_X1 U8242 ( .A1(n9609), .A2(P1_ADDR_REG_12__SCAN_IN), .ZN(n6504) );
  OAI211_X1 U8243 ( .C1(n9724), .C2(n6505), .A(n7248), .B(n6504), .ZN(n6506)
         );
  AOI21_X1 U8244 ( .B1(n6507), .B2(n9713), .A(n6506), .ZN(n6508) );
  NAND2_X1 U8245 ( .A1(n6509), .A2(n6508), .ZN(P1_U3255) );
  XNOR2_X1 U8246 ( .A(n8135), .B(n6511), .ZN(n6512) );
  NAND2_X1 U8247 ( .A1(n6512), .A2(n5513), .ZN(n6514) );
  AOI22_X1 U8248 ( .A1(n8809), .A2(n5101), .B1(n6130), .B2(n8807), .ZN(n6513)
         );
  NAND2_X1 U8249 ( .A1(n6514), .A2(n6513), .ZN(n10056) );
  AOI21_X1 U8250 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(n8815), .A(n10056), .ZN(
        n6521) );
  NAND2_X1 U8251 ( .A1(n8135), .A2(n6516), .ZN(n6517) );
  NAND2_X1 U8252 ( .A1(n6515), .A2(n6517), .ZN(n10057) );
  NAND2_X1 U8253 ( .A1(n7399), .A2(n10057), .ZN(n6520) );
  AOI22_X1 U8254 ( .A1(n8816), .A2(n6518), .B1(n8797), .B2(
        P2_REG2_REG_1__SCAN_IN), .ZN(n6519) );
  OAI211_X1 U8255 ( .C1(n8797), .C2(n6521), .A(n6520), .B(n6519), .ZN(P2_U3232) );
  INV_X1 U8256 ( .A(n6522), .ZN(n6523) );
  OR2_X1 U8257 ( .A1(n7636), .A2(n6525), .ZN(n6529) );
  OR2_X1 U8258 ( .A1(n4347), .A2(n6526), .ZN(n6528) );
  OR2_X1 U8259 ( .A1(n8173), .A2(n9635), .ZN(n6527) );
  AOI22_X1 U8260 ( .A1(n9077), .A2(n7709), .B1(n8210), .B2(n6252), .ZN(n6530)
         );
  XNOR2_X1 U8261 ( .A(n6530), .B(n7949), .ZN(n6531) );
  NOR2_X1 U8262 ( .A1(n6567), .A2(n4425), .ZN(n6532) );
  INV_X1 U8263 ( .A(n9077), .ZN(n8203) );
  OAI22_X1 U8264 ( .A1(n8203), .A2(n6158), .B1(n9861), .B2(n7948), .ZN(n6566)
         );
  XNOR2_X1 U8265 ( .A(n6532), .B(n6566), .ZN(n6544) );
  INV_X1 U8266 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n6844) );
  INV_X1 U8267 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n6533) );
  OR2_X1 U8268 ( .A1(n8177), .A2(n6533), .ZN(n6534) );
  OAI21_X1 U8269 ( .B1(n7941), .B2(n6844), .A(n6534), .ZN(n6539) );
  NAND2_X1 U8270 ( .A1(n6535), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n6581) );
  OR2_X1 U8271 ( .A1(n6535), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n6536) );
  NAND2_X1 U8272 ( .A1(n6581), .A2(n6536), .ZN(n6843) );
  OR2_X1 U8273 ( .A1(n8179), .A2(n9871), .ZN(n6537) );
  OAI21_X1 U8274 ( .B1(n6262), .B2(n6843), .A(n6537), .ZN(n6538) );
  AOI22_X1 U8275 ( .A1(n9225), .A2(n9078), .B1(n9076), .B2(n9052), .ZN(n9782)
         );
  OAI22_X1 U8276 ( .A1(n9056), .A2(n9782), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n6540), .ZN(n6542) );
  NOR2_X1 U8277 ( .A1(n9021), .A2(n9785), .ZN(n6541) );
  AOI211_X1 U8278 ( .C1(n8210), .C2(n9023), .A(n6542), .B(n6541), .ZN(n6543)
         );
  OAI21_X1 U8279 ( .B1(n6544), .B2(n9036), .A(n6543), .ZN(P1_U3227) );
  NAND2_X1 U8280 ( .A1(n6546), .A2(n6545), .ZN(n6547) );
  AOI21_X1 U8281 ( .B1(n9832), .B2(n6549), .A(n9753), .ZN(n6556) );
  INV_X1 U8282 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n6551) );
  OAI21_X1 U8283 ( .B1(n9799), .B2(n6551), .A(n6550), .ZN(n6552) );
  AOI21_X1 U8284 ( .B1(n6553), .B2(n8357), .A(n6552), .ZN(n6554) );
  MUX2_X1 U8285 ( .A(n6554), .B(n9568), .S(n9836), .Z(n6555) );
  OAI21_X1 U8286 ( .B1(n6556), .B2(n9830), .A(n6555), .ZN(P1_U3293) );
  XOR2_X1 U8287 ( .A(n6557), .B(n8136), .Z(n6558) );
  AOI222_X1 U8288 ( .A1(n5513), .A2(n6558), .B1(n8600), .B2(n8809), .C1(n5101), 
        .C2(n8807), .ZN(n10063) );
  XNOR2_X1 U8289 ( .A(n6559), .B(n8136), .ZN(n10066) );
  OAI22_X1 U8290 ( .A1(n8681), .A2(n10064), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        n10038), .ZN(n6561) );
  AND2_X1 U8291 ( .A1(n8797), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n6560) );
  AOI211_X1 U8292 ( .C1(n7399), .C2(n10066), .A(n6561), .B(n6560), .ZN(n6562)
         );
  OAI21_X1 U8293 ( .B1(n10063), .B2(n8797), .A(n6562), .ZN(P2_U3230) );
  INV_X1 U8294 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n6563) );
  INV_X1 U8295 ( .A(n7712), .ZN(n6565) );
  OAI222_X1 U8296 ( .A1(n7913), .A2(n6563), .B1(n7915), .B2(n6565), .C1(n6070), 
        .C2(P1_U3086), .ZN(P1_U3336) );
  INV_X1 U8297 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n6564) );
  OAI222_X1 U8298 ( .A1(P2_U3151), .A2(n8668), .B1(n8470), .B2(n6565), .C1(
        n6564), .C2(n8491), .ZN(P2_U3276) );
  NAND2_X1 U8299 ( .A1(n9076), .A2(n7709), .ZN(n6573) );
  AOI22_X1 U8300 ( .A1(n7714), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n7713), .B2(
        n6568), .ZN(n6571) );
  NAND2_X1 U8301 ( .A1(n6569), .A2(n7777), .ZN(n6570) );
  INV_X1 U8302 ( .A(n6252), .ZN(n7717) );
  OR2_X1 U8303 ( .A1(n6643), .A2(n7717), .ZN(n6572) );
  NAND2_X1 U8304 ( .A1(n6573), .A2(n6572), .ZN(n6574) );
  XNOR2_X1 U8305 ( .A(n6574), .B(n7949), .ZN(n6753) );
  NAND2_X1 U8306 ( .A1(n9076), .A2(n7924), .ZN(n6576) );
  OR2_X1 U8307 ( .A1(n6643), .A2(n7948), .ZN(n6575) );
  NAND2_X1 U8308 ( .A1(n6576), .A2(n6575), .ZN(n6752) );
  INV_X1 U8309 ( .A(n6752), .ZN(n6754) );
  XNOR2_X1 U8310 ( .A(n6753), .B(n6754), .ZN(n6577) );
  XNOR2_X1 U8311 ( .A(n6757), .B(n6577), .ZN(n6592) );
  NAND2_X1 U8312 ( .A1(n9077), .A2(n9225), .ZN(n6588) );
  OR2_X1 U8313 ( .A1(n8177), .A2(n6578), .ZN(n6579) );
  OAI21_X1 U8314 ( .B1(n7941), .B2(n6475), .A(n6579), .ZN(n6586) );
  OR2_X2 U8315 ( .A1(n6581), .A2(n6580), .ZN(n6658) );
  NAND2_X1 U8316 ( .A1(n6581), .A2(n6580), .ZN(n6582) );
  NAND2_X1 U8317 ( .A1(n6658), .A2(n6582), .ZN(n9769) );
  INV_X1 U8318 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n6583) );
  OR2_X1 U8319 ( .A1(n8179), .A2(n6583), .ZN(n6584) );
  OAI21_X1 U8320 ( .B1(n6262), .B2(n9769), .A(n6584), .ZN(n6585) );
  NAND2_X1 U8321 ( .A1(n9075), .A2(n9052), .ZN(n6587) );
  NAND2_X1 U8322 ( .A1(n6588), .A2(n6587), .ZN(n6835) );
  AOI22_X1 U8323 ( .A1(n9018), .A2(n6835), .B1(P1_REG3_REG_6__SCAN_IN), .B2(
        P1_U3086), .ZN(n6590) );
  NAND2_X1 U8324 ( .A1(n9023), .A2(n6642), .ZN(n6589) );
  OAI211_X1 U8325 ( .C1(n9021), .C2(n6843), .A(n6590), .B(n6589), .ZN(n6591)
         );
  AOI21_X1 U8326 ( .B1(n6592), .B2(n9050), .A(n6591), .ZN(n6593) );
  INV_X1 U8327 ( .A(n6593), .ZN(P1_U3239) );
  XNOR2_X1 U8328 ( .A(n6594), .B(n8138), .ZN(n6595) );
  AOI222_X1 U8329 ( .A1(n5513), .A2(n6595), .B1(n8597), .B2(n8809), .C1(n8599), 
        .C2(n8807), .ZN(n10084) );
  NAND2_X1 U8330 ( .A1(n6597), .A2(n6596), .ZN(n6598) );
  XOR2_X1 U8331 ( .A(n8138), .B(n6598), .Z(n10082) );
  NOR2_X1 U8332 ( .A1(n10050), .A2(n5747), .ZN(n6601) );
  OAI22_X1 U8333 ( .A1(n8681), .A2(n6599), .B1(n6727), .B2(n10038), .ZN(n6600)
         );
  AOI211_X1 U8334 ( .C1(n10082), .C2(n7399), .A(n6601), .B(n6600), .ZN(n6602)
         );
  OAI21_X1 U8335 ( .B1(n10084), .B2(n8797), .A(n6602), .ZN(P2_U3227) );
  NAND2_X1 U8336 ( .A1(n6459), .A2(n6603), .ZN(n6604) );
  XNOR2_X1 U8337 ( .A(n6604), .B(n8141), .ZN(n10092) );
  NAND2_X1 U8338 ( .A1(n6605), .A2(n8141), .ZN(n6606) );
  NAND3_X1 U8339 ( .A1(n6607), .A2(n5513), .A3(n6606), .ZN(n6609) );
  AOI22_X1 U8340 ( .A1(n8809), .A2(n8595), .B1(n8597), .B2(n8807), .ZN(n6608)
         );
  AND2_X1 U8341 ( .A1(n6609), .A2(n6608), .ZN(n10096) );
  MUX2_X1 U8342 ( .A(n10096), .B(n6610), .S(n8797), .Z(n6613) );
  INV_X1 U8343 ( .A(n7086), .ZN(n6611) );
  AOI22_X1 U8344 ( .A1(n8816), .A2(n10093), .B1(n8815), .B2(n6611), .ZN(n6612)
         );
  OAI211_X1 U8345 ( .C1(n10092), .C2(n8819), .A(n6613), .B(n6612), .ZN(
        P2_U3225) );
  INV_X1 U8346 ( .A(n9844), .ZN(n6614) );
  NAND2_X1 U8347 ( .A1(n9080), .A2(n9844), .ZN(n8407) );
  XNOR2_X1 U8348 ( .A(n8358), .B(n6664), .ZN(n6620) );
  INV_X1 U8349 ( .A(n6618), .ZN(n6619) );
  OAI21_X1 U8350 ( .B1(n6620), .B2(n9746), .A(n6619), .ZN(n9845) );
  AOI21_X1 U8351 ( .B1(P1_REG3_REG_2__SCAN_IN), .B2(n9822), .A(n9845), .ZN(
        n6633) );
  NAND2_X1 U8352 ( .A1(n6621), .A2(n4349), .ZN(n6622) );
  OAI21_X2 U8353 ( .B1(n9836), .B2(n9817), .A(n9754), .ZN(n9809) );
  AND2_X1 U8354 ( .A1(n9081), .A2(n6623), .ZN(n9816) );
  NAND2_X1 U8355 ( .A1(n6624), .A2(n6626), .ZN(n6625) );
  XNOR2_X1 U8356 ( .A(n6634), .B(n8358), .ZN(n9847) );
  NAND2_X1 U8357 ( .A1(n6626), .A2(n9830), .ZN(n9828) );
  AOI21_X1 U8358 ( .B1(n9828), .B2(n6614), .A(n9775), .ZN(n6628) );
  NAND2_X1 U8359 ( .A1(n6628), .A2(n9805), .ZN(n9843) );
  NOR2_X1 U8360 ( .A1(n9248), .A2(n9843), .ZN(n6631) );
  OAI22_X1 U8361 ( .A1(n9844), .A2(n9825), .B1(n9335), .B2(n6629), .ZN(n6630)
         );
  AOI211_X1 U8362 ( .C1(n9809), .C2(n9847), .A(n6631), .B(n6630), .ZN(n6632)
         );
  OAI21_X1 U8363 ( .B1(n6633), .B2(n9823), .A(n6632), .ZN(P1_U3291) );
  NAND2_X1 U8364 ( .A1(n6634), .A2(n8358), .ZN(n6636) );
  OR2_X1 U8365 ( .A1(n9080), .A2(n6614), .ZN(n6635) );
  NAND2_X1 U8366 ( .A1(n6636), .A2(n6635), .ZN(n9803) );
  NAND2_X1 U8367 ( .A1(n9079), .A2(n9849), .ZN(n8201) );
  AND2_X1 U8368 ( .A1(n8196), .A2(n8201), .ZN(n9796) );
  INV_X1 U8369 ( .A(n9796), .ZN(n9804) );
  NAND2_X1 U8370 ( .A1(n9803), .A2(n9804), .ZN(n6638) );
  OR2_X1 U8371 ( .A1(n9079), .A2(n6686), .ZN(n6637) );
  NAND2_X1 U8372 ( .A1(n6638), .A2(n6637), .ZN(n6811) );
  NAND2_X1 U8373 ( .A1(n6639), .A2(n6817), .ZN(n8413) );
  NAND2_X1 U8374 ( .A1(n9078), .A2(n9855), .ZN(n8200) );
  NAND2_X1 U8375 ( .A1(n8413), .A2(n8200), .ZN(n8361) );
  NAND2_X1 U8376 ( .A1(n6811), .A2(n8361), .ZN(n6641) );
  NAND2_X1 U8377 ( .A1(n6639), .A2(n9855), .ZN(n6640) );
  NAND2_X1 U8378 ( .A1(n6641), .A2(n6640), .ZN(n9789) );
  NAND2_X1 U8379 ( .A1(n8203), .A2(n8210), .ZN(n8412) );
  NAND2_X1 U8380 ( .A1(n9077), .A2(n9861), .ZN(n8420) );
  INV_X1 U8381 ( .A(n9781), .ZN(n9790) );
  NAND2_X1 U8382 ( .A1(n8203), .A2(n9861), .ZN(n6838) );
  INV_X1 U8383 ( .A(n9076), .ZN(n8206) );
  NAND2_X1 U8384 ( .A1(n8206), .A2(n6643), .ZN(n6644) );
  AND2_X1 U8385 ( .A1(n6838), .A2(n6644), .ZN(n6647) );
  NAND2_X1 U8386 ( .A1(n9076), .A2(n6643), .ZN(n8192) );
  INV_X1 U8387 ( .A(n8365), .ZN(n6840) );
  INV_X1 U8388 ( .A(n6644), .ZN(n6645) );
  NOR2_X1 U8389 ( .A1(n6840), .A2(n6645), .ZN(n6646) );
  NAND2_X1 U8390 ( .A1(n6648), .A2(n7777), .ZN(n6651) );
  AOI22_X1 U8391 ( .A1(n7714), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n7713), .B2(
        n6649), .ZN(n6650) );
  NAND2_X1 U8392 ( .A1(n9772), .A2(n9075), .ZN(n8363) );
  INV_X1 U8393 ( .A(n9075), .ZN(n6758) );
  NAND2_X1 U8394 ( .A1(n6652), .A2(n7777), .ZN(n6655) );
  AOI22_X1 U8395 ( .A1(n7714), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n7713), .B2(
        n6653), .ZN(n6654) );
  INV_X1 U8396 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n6685) );
  OR2_X1 U8397 ( .A1(n8177), .A2(n9935), .ZN(n6656) );
  OAI21_X1 U8398 ( .B1(n7941), .B2(n6685), .A(n6656), .ZN(n6663) );
  OR2_X2 U8399 ( .A1(n6658), .A2(n6657), .ZN(n6674) );
  NAND2_X1 U8400 ( .A1(n6658), .A2(n6657), .ZN(n6659) );
  NAND2_X1 U8401 ( .A1(n6674), .A2(n6659), .ZN(n7139) );
  INV_X1 U8402 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n6660) );
  OR2_X1 U8403 ( .A1(n8179), .A2(n6660), .ZN(n6661) );
  OAI21_X1 U8404 ( .B1(n6262), .B2(n7139), .A(n6661), .ZN(n6662) );
  OR2_X1 U8405 ( .A1(n7141), .A2(n6700), .ZN(n8190) );
  NAND2_X1 U8406 ( .A1(n7141), .A2(n6700), .ZN(n8222) );
  XNOR2_X1 U8407 ( .A(n6703), .B(n6702), .ZN(n9878) );
  INV_X1 U8408 ( .A(n9878), .ZN(n6692) );
  NAND2_X1 U8409 ( .A1(n6664), .A2(n8407), .ZN(n8199) );
  NAND2_X1 U8410 ( .A1(n6665), .A2(n8413), .ZN(n9780) );
  NAND2_X1 U8411 ( .A1(n9780), .A2(n9781), .ZN(n6666) );
  NAND2_X1 U8412 ( .A1(n6833), .A2(n8365), .ZN(n6832) );
  NAND2_X1 U8413 ( .A1(n6832), .A2(n8416), .ZN(n9764) );
  AND2_X1 U8414 ( .A1(n9764), .A2(n4422), .ZN(n9762) );
  INV_X1 U8415 ( .A(n8228), .ZN(n6667) );
  OR2_X1 U8416 ( .A1(n9762), .A2(n6667), .ZN(n6668) );
  XNOR2_X1 U8417 ( .A(n6668), .B(n6702), .ZN(n6669) );
  NAND2_X1 U8418 ( .A1(n6669), .A2(n9821), .ZN(n6684) );
  NAND2_X1 U8419 ( .A1(n9075), .A2(n9225), .ZN(n6682) );
  INV_X1 U8420 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n6672) );
  INV_X1 U8421 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n6670) );
  OR2_X1 U8422 ( .A1(n8177), .A2(n6670), .ZN(n6671) );
  OAI21_X1 U8423 ( .B1(n7941), .B2(n6672), .A(n6671), .ZN(n6680) );
  INV_X1 U8424 ( .A(n6708), .ZN(n6676) );
  NAND2_X1 U8425 ( .A1(n6674), .A2(n6673), .ZN(n6675) );
  NAND2_X1 U8426 ( .A1(n6676), .A2(n6675), .ZN(n7341) );
  INV_X1 U8427 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n6677) );
  OR2_X1 U8428 ( .A1(n8179), .A2(n6677), .ZN(n6678) );
  OAI21_X1 U8429 ( .B1(n6262), .B2(n7341), .A(n6678), .ZN(n6679) );
  NAND2_X1 U8430 ( .A1(n9073), .A2(n9052), .ZN(n6681) );
  NAND2_X1 U8431 ( .A1(n6682), .A2(n6681), .ZN(n7137) );
  INV_X1 U8432 ( .A(n7137), .ZN(n6683) );
  NAND2_X1 U8433 ( .A1(n6684), .A2(n6683), .ZN(n9884) );
  NAND2_X1 U8434 ( .A1(n9884), .A2(n9335), .ZN(n6691) );
  OAI22_X1 U8435 ( .A1(n9335), .A2(n6685), .B1(n7139), .B2(n9799), .ZN(n6689)
         );
  INV_X1 U8436 ( .A(n7141), .ZN(n9881) );
  OAI21_X1 U8437 ( .B1(n9774), .B2(n9881), .A(n9829), .ZN(n6687) );
  OR2_X1 U8438 ( .A1(n6687), .A2(n6704), .ZN(n9879) );
  NOR2_X1 U8439 ( .A1(n9879), .A2(n9248), .ZN(n6688) );
  AOI211_X1 U8440 ( .C1(n9753), .C2(n7141), .A(n6689), .B(n6688), .ZN(n6690)
         );
  OAI211_X1 U8441 ( .C1(n9378), .C2(n6692), .A(n6691), .B(n6690), .ZN(P1_U3285) );
  INV_X1 U8442 ( .A(n7341), .ZN(n6699) );
  NAND2_X1 U8443 ( .A1(n9074), .A2(n9225), .ZN(n7336) );
  INV_X1 U8444 ( .A(n7336), .ZN(n6698) );
  NAND2_X1 U8445 ( .A1(n6693), .A2(n7777), .ZN(n6695) );
  AOI22_X1 U8446 ( .A1(n7714), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n7713), .B2(
        n9091), .ZN(n6694) );
  INV_X1 U8447 ( .A(n9073), .ZN(n7223) );
  NAND2_X1 U8448 ( .A1(n7338), .A2(n7223), .ZN(n8229) );
  NAND2_X1 U8449 ( .A1(n8233), .A2(n8229), .ZN(n6798) );
  NAND2_X1 U8450 ( .A1(n8222), .A2(n8228), .ZN(n8219) );
  OAI21_X1 U8451 ( .B1(n9762), .B2(n8219), .A(n8190), .ZN(n6696) );
  XOR2_X1 U8452 ( .A(n6798), .B(n6696), .Z(n6697) );
  NOR2_X1 U8453 ( .A1(n6697), .A2(n9746), .ZN(n9889) );
  AOI211_X1 U8454 ( .C1(n9822), .C2(n6699), .A(n6698), .B(n9889), .ZN(n6718)
         );
  NAND2_X1 U8455 ( .A1(n9881), .A2(n6700), .ZN(n6701) );
  XNOR2_X1 U8456 ( .A(n6799), .B(n6798), .ZN(n9891) );
  NAND2_X1 U8457 ( .A1(n6704), .A2(n9888), .ZN(n6801) );
  OAI211_X1 U8458 ( .C1(n6704), .C2(n9888), .A(n9829), .B(n6801), .ZN(n9887)
         );
  INV_X1 U8459 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n6800) );
  INV_X1 U8460 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n6705) );
  OR2_X1 U8461 ( .A1(n8179), .A2(n6705), .ZN(n6706) );
  OAI21_X1 U8462 ( .B1(n7941), .B2(n6800), .A(n6706), .ZN(n6707) );
  INV_X1 U8463 ( .A(n6707), .ZN(n6714) );
  NAND2_X1 U8464 ( .A1(n6708), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n6788) );
  OR2_X1 U8465 ( .A1(n6708), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n6709) );
  NAND2_X1 U8466 ( .A1(n6788), .A2(n6709), .ZN(n7302) );
  INV_X1 U8467 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n6710) );
  OR2_X1 U8468 ( .A1(n8177), .A2(n6710), .ZN(n6711) );
  OAI21_X1 U8469 ( .B1(n6262), .B2(n7302), .A(n6711), .ZN(n6712) );
  INV_X1 U8470 ( .A(n6712), .ZN(n6713) );
  OR2_X1 U8471 ( .A1(n7376), .A2(n9162), .ZN(n7337) );
  AOI21_X1 U8472 ( .B1(n9887), .B2(n7337), .A(n9248), .ZN(n6716) );
  OAI22_X1 U8473 ( .A1(n9888), .A2(n9825), .B1(n6672), .B2(n9335), .ZN(n6715)
         );
  AOI211_X1 U8474 ( .C1(n9891), .C2(n9809), .A(n6716), .B(n6715), .ZN(n6717)
         );
  OAI21_X1 U8475 ( .B1(n6718), .B2(n9823), .A(n6717), .ZN(P1_U3284) );
  AOI211_X1 U8476 ( .C1(n6721), .C2(n6720), .A(n9543), .B(n6719), .ZN(n6722)
         );
  INV_X1 U8477 ( .A(n6722), .ZN(n6726) );
  INV_X1 U8478 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n6948) );
  NOR2_X1 U8479 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6948), .ZN(n9999) );
  AOI21_X1 U8480 ( .B1(n8547), .B2(n8597), .A(n9999), .ZN(n6723) );
  OAI21_X1 U8481 ( .B1(n4571), .B2(n8530), .A(n6723), .ZN(n6724) );
  AOI21_X1 U8482 ( .B1(n10081), .B2(n9539), .A(n6724), .ZN(n6725) );
  OAI211_X1 U8483 ( .C1(n6727), .C2(n8577), .A(n6726), .B(n6725), .ZN(P2_U3179) );
  AOI21_X1 U8484 ( .B1(n6730), .B2(n6729), .A(n6728), .ZN(n6748) );
  INV_X1 U8485 ( .A(n6731), .ZN(n6732) );
  NOR2_X1 U8486 ( .A1(n6733), .A2(n6732), .ZN(n6735) );
  NAND2_X1 U8487 ( .A1(n6736), .A2(n6735), .ZN(n6734) );
  OAI211_X1 U8488 ( .C1(n6736), .C2(n6735), .A(n10029), .B(n6734), .ZN(n6747)
         );
  OAI21_X1 U8489 ( .B1(n6739), .B2(n6738), .A(n6737), .ZN(n6745) );
  INV_X1 U8490 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n6743) );
  NOR2_X1 U8491 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6740), .ZN(n7530) );
  AOI21_X1 U8492 ( .B1(n10020), .B2(n6741), .A(n7530), .ZN(n6742) );
  OAI21_X1 U8493 ( .B1(n10033), .B2(n6743), .A(n6742), .ZN(n6744) );
  AOI21_X1 U8494 ( .B1(n6745), .B2(n10017), .A(n6744), .ZN(n6746) );
  OAI211_X1 U8495 ( .C1(n6748), .C2(n10024), .A(n6747), .B(n6746), .ZN(
        P2_U3194) );
  INV_X1 U8496 ( .A(n7723), .ZN(n6751) );
  INV_X1 U8497 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7724) );
  OAI222_X1 U8498 ( .A1(n7915), .A2(n6751), .B1(P1_U3086), .B2(n6749), .C1(
        n7724), .C2(n7913), .ZN(P1_U3335) );
  INV_X1 U8499 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n6750) );
  OAI222_X1 U8500 ( .A1(n8115), .A2(P2_U3151), .B1(n8494), .B2(n6751), .C1(
        n6750), .C2(n8491), .ZN(P2_U3275) );
  NOR2_X1 U8501 ( .A1(n6753), .A2(n6752), .ZN(n6756) );
  INV_X1 U8502 ( .A(n6753), .ZN(n6755) );
  OAI22_X1 U8503 ( .A1(n9772), .A2(n7717), .B1(n6758), .B2(n7948), .ZN(n6759)
         );
  XNOR2_X1 U8504 ( .A(n6759), .B(n7922), .ZN(n6763) );
  OR2_X1 U8505 ( .A1(n9772), .A2(n7948), .ZN(n6761) );
  NAND2_X1 U8506 ( .A1(n9075), .A2(n7924), .ZN(n6760) );
  AND2_X1 U8507 ( .A1(n6761), .A2(n6760), .ZN(n6762) );
  NOR2_X1 U8508 ( .A1(n6763), .A2(n6762), .ZN(n7130) );
  INV_X1 U8509 ( .A(n7130), .ZN(n6764) );
  NAND2_X1 U8510 ( .A1(n6763), .A2(n6762), .ZN(n7131) );
  NAND2_X1 U8511 ( .A1(n6764), .A2(n7131), .ZN(n6765) );
  XNOR2_X1 U8512 ( .A(n7132), .B(n6765), .ZN(n6771) );
  NAND2_X1 U8513 ( .A1(n9076), .A2(n9225), .ZN(n6767) );
  NAND2_X1 U8514 ( .A1(n9074), .A2(n9052), .ZN(n6766) );
  NAND2_X1 U8515 ( .A1(n6767), .A2(n6766), .ZN(n9767) );
  AOI22_X1 U8516 ( .A1(n9018), .A2(n9767), .B1(P1_REG3_REG_7__SCAN_IN), .B2(
        P1_U3086), .ZN(n6769) );
  NAND2_X1 U8517 ( .A1(n9023), .A2(n9873), .ZN(n6768) );
  OAI211_X1 U8518 ( .C1(n9021), .C2(n9769), .A(n6769), .B(n6768), .ZN(n6770)
         );
  AOI21_X1 U8519 ( .B1(n6771), .B2(n9050), .A(n6770), .ZN(n6772) );
  INV_X1 U8520 ( .A(n6772), .ZN(P1_U3213) );
  NAND2_X1 U8521 ( .A1(n6773), .A2(n7777), .ZN(n6775) );
  AOI22_X1 U8522 ( .A1(n7714), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n7713), .B2(
        n9489), .ZN(n6774) );
  OR2_X1 U8523 ( .A1(n7299), .A2(n7376), .ZN(n8422) );
  AND2_X1 U8524 ( .A1(n7299), .A2(n7376), .ZN(n8232) );
  INV_X1 U8525 ( .A(n8232), .ZN(n9745) );
  NAND2_X1 U8526 ( .A1(n8233), .A2(n8190), .ZN(n8366) );
  INV_X1 U8527 ( .A(n8366), .ZN(n6776) );
  NAND2_X1 U8528 ( .A1(n6776), .A2(n8219), .ZN(n6777) );
  INV_X1 U8529 ( .A(n6833), .ZN(n6778) );
  NAND3_X1 U8530 ( .A1(n8417), .A2(n6778), .A3(n8416), .ZN(n6781) );
  NAND2_X1 U8531 ( .A1(n8363), .A2(n8192), .ZN(n6779) );
  OR2_X1 U8532 ( .A1(n8366), .A2(n6779), .ZN(n6780) );
  NAND2_X1 U8533 ( .A1(n8417), .A2(n6780), .ZN(n8423) );
  AND2_X1 U8534 ( .A1(n6781), .A2(n8423), .ZN(n6782) );
  NAND2_X1 U8535 ( .A1(n6782), .A2(n8369), .ZN(n7148) );
  OAI21_X1 U8536 ( .B1(n8369), .B2(n6782), .A(n7148), .ZN(n6797) );
  INV_X1 U8537 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n6785) );
  OR2_X1 U8538 ( .A1(n8177), .A2(n6783), .ZN(n6784) );
  OAI21_X1 U8539 ( .B1(n7941), .B2(n6785), .A(n6784), .ZN(n6786) );
  INV_X1 U8540 ( .A(n6786), .ZN(n6794) );
  OR2_X2 U8541 ( .A1(n6788), .A2(n6787), .ZN(n7154) );
  NAND2_X1 U8542 ( .A1(n6788), .A2(n6787), .ZN(n6789) );
  NAND2_X1 U8543 ( .A1(n7154), .A2(n6789), .ZN(n9751) );
  INV_X1 U8544 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n6790) );
  OR2_X1 U8545 ( .A1(n8179), .A2(n6790), .ZN(n6791) );
  OAI21_X1 U8546 ( .B1(n6262), .B2(n9751), .A(n6791), .ZN(n6792) );
  INV_X1 U8547 ( .A(n6792), .ZN(n6793) );
  OR2_X1 U8548 ( .A1(n9070), .A2(n9162), .ZN(n6796) );
  NAND2_X1 U8549 ( .A1(n9073), .A2(n9225), .ZN(n6795) );
  NAND2_X1 U8550 ( .A1(n6796), .A2(n6795), .ZN(n7298) );
  AOI21_X1 U8551 ( .B1(n6797), .B2(n9821), .A(n7298), .ZN(n9893) );
  XNOR2_X1 U8552 ( .A(n7172), .B(n8369), .ZN(n9896) );
  NAND2_X1 U8553 ( .A1(n9896), .A2(n9809), .ZN(n6806) );
  OAI22_X1 U8554 ( .A1(n9335), .A2(n6800), .B1(n7302), .B2(n9799), .ZN(n6804)
         );
  INV_X1 U8555 ( .A(n6801), .ZN(n6802) );
  INV_X1 U8556 ( .A(n7299), .ZN(n9894) );
  OAI211_X1 U8557 ( .C1(n6802), .C2(n9894), .A(n9829), .B(n9755), .ZN(n9892)
         );
  NOR2_X1 U8558 ( .A1(n9892), .A2(n9248), .ZN(n6803) );
  AOI211_X1 U8559 ( .C1(n9753), .C2(n7299), .A(n6804), .B(n6803), .ZN(n6805)
         );
  OAI211_X1 U8560 ( .C1(n9836), .C2(n9893), .A(n6806), .B(n6805), .ZN(P1_U3283) );
  INV_X1 U8561 ( .A(n8361), .ZN(n6808) );
  XNOR2_X1 U8562 ( .A(n6807), .B(n6808), .ZN(n6810) );
  AOI21_X1 U8563 ( .B1(n6810), .B2(n9821), .A(n6809), .ZN(n9859) );
  XNOR2_X1 U8564 ( .A(n6811), .B(n8361), .ZN(n9857) );
  NAND2_X1 U8565 ( .A1(n9806), .A2(n6817), .ZN(n6812) );
  NAND2_X1 U8566 ( .A1(n6812), .A2(n9829), .ZN(n6813) );
  OR2_X1 U8567 ( .A1(n6813), .A2(n9792), .ZN(n9854) );
  OAI22_X1 U8568 ( .A1(n9335), .A2(n6815), .B1(n6814), .B2(n9799), .ZN(n6816)
         );
  AOI21_X1 U8569 ( .B1(n9753), .B2(n6817), .A(n6816), .ZN(n6818) );
  OAI21_X1 U8570 ( .B1(n9248), .B2(n9854), .A(n6818), .ZN(n6819) );
  AOI21_X1 U8571 ( .B1(n9857), .B2(n9809), .A(n6819), .ZN(n6820) );
  OAI21_X1 U8572 ( .B1(n9859), .B2(n9823), .A(n6820), .ZN(P1_U3289) );
  OAI21_X1 U8573 ( .B1(n6823), .B2(n6822), .A(n6821), .ZN(n6824) );
  NAND2_X1 U8574 ( .A1(n6824), .A2(n8572), .ZN(n6830) );
  INV_X1 U8575 ( .A(n8598), .ZN(n6826) );
  NOR2_X1 U8576 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n4888), .ZN(n10018) );
  AOI21_X1 U8577 ( .B1(n8547), .B2(n8596), .A(n10018), .ZN(n6825) );
  OAI21_X1 U8578 ( .B1(n6826), .B2(n8530), .A(n6825), .ZN(n6827) );
  AOI21_X1 U8579 ( .B1(n6828), .B2(n9539), .A(n6827), .ZN(n6829) );
  OAI211_X1 U8580 ( .C1(n6831), .C2(n8577), .A(n6830), .B(n6829), .ZN(P2_U3153) );
  OAI21_X1 U8581 ( .B1(n8365), .B2(n6833), .A(n6832), .ZN(n6834) );
  NAND2_X1 U8582 ( .A1(n6834), .A2(n9821), .ZN(n6837) );
  INV_X1 U8583 ( .A(n6835), .ZN(n6836) );
  NAND2_X1 U8584 ( .A1(n6837), .A2(n6836), .ZN(n9869) );
  INV_X1 U8585 ( .A(n9869), .ZN(n6849) );
  NAND2_X1 U8586 ( .A1(n6839), .A2(n6838), .ZN(n6841) );
  XNOR2_X1 U8587 ( .A(n6841), .B(n6840), .ZN(n9866) );
  AOI21_X1 U8588 ( .B1(n9791), .B2(n6642), .A(n9775), .ZN(n6842) );
  NAND2_X1 U8589 ( .A1(n6842), .A2(n9776), .ZN(n9867) );
  OAI22_X1 U8590 ( .A1(n9335), .A2(n6844), .B1(n6843), .B2(n9799), .ZN(n6845)
         );
  AOI21_X1 U8591 ( .B1(n9753), .B2(n6642), .A(n6845), .ZN(n6846) );
  OAI21_X1 U8592 ( .B1(n9867), .B2(n9248), .A(n6846), .ZN(n6847) );
  AOI21_X1 U8593 ( .B1(n9866), .B2(n9809), .A(n6847), .ZN(n6848) );
  OAI21_X1 U8594 ( .B1(n6849), .B2(n9823), .A(n6848), .ZN(P1_U3287) );
  INV_X1 U8595 ( .A(SI_6_), .ZN(n7028) );
  AOI22_X1 U8596 ( .A1(SI_2_), .A2(keyinput_f30), .B1(P2_REG3_REG_10__SCAN_IN), 
        .B2(keyinput_f39), .ZN(n6850) );
  OAI221_X1 U8597 ( .B1(SI_2_), .B2(keyinput_f30), .C1(P2_REG3_REG_10__SCAN_IN), .C2(keyinput_f39), .A(n6850), .ZN(n6857) );
  AOI22_X1 U8598 ( .A1(SI_0_), .A2(keyinput_f32), .B1(P2_REG3_REG_23__SCAN_IN), 
        .B2(keyinput_f38), .ZN(n6851) );
  OAI221_X1 U8599 ( .B1(SI_0_), .B2(keyinput_f32), .C1(P2_REG3_REG_23__SCAN_IN), .C2(keyinput_f38), .A(n6851), .ZN(n6856) );
  AOI22_X1 U8600 ( .A1(keyinput_f0), .A2(P2_WR_REG_SCAN_IN), .B1(
        P2_REG3_REG_11__SCAN_IN), .B2(keyinput_f58), .ZN(n6852) );
  OAI221_X1 U8601 ( .B1(keyinput_f0), .B2(P2_WR_REG_SCAN_IN), .C1(
        P2_REG3_REG_11__SCAN_IN), .C2(keyinput_f58), .A(n6852), .ZN(n6855) );
  AOI22_X1 U8602 ( .A1(SI_7_), .A2(keyinput_f25), .B1(SI_20_), .B2(
        keyinput_f12), .ZN(n6853) );
  OAI221_X1 U8603 ( .B1(SI_7_), .B2(keyinput_f25), .C1(SI_20_), .C2(
        keyinput_f12), .A(n6853), .ZN(n6854) );
  NOR4_X1 U8604 ( .A1(n6857), .A2(n6856), .A3(n6855), .A4(n6854), .ZN(n6884)
         );
  XNOR2_X1 U8605 ( .A(n5075), .B(keyinput_f54), .ZN(n6864) );
  AOI22_X1 U8606 ( .A1(SI_8_), .A2(keyinput_f24), .B1(SI_26_), .B2(keyinput_f6), .ZN(n6858) );
  OAI221_X1 U8607 ( .B1(SI_8_), .B2(keyinput_f24), .C1(SI_26_), .C2(
        keyinput_f6), .A(n6858), .ZN(n6863) );
  AOI22_X1 U8608 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(keyinput_f40), .B1(
        P2_REG3_REG_22__SCAN_IN), .B2(keyinput_f57), .ZN(n6859) );
  OAI221_X1 U8609 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(keyinput_f40), .C1(
        P2_REG3_REG_22__SCAN_IN), .C2(keyinput_f57), .A(n6859), .ZN(n6862) );
  AOI22_X1 U8610 ( .A1(SI_23_), .A2(keyinput_f9), .B1(P2_REG3_REG_9__SCAN_IN), 
        .B2(keyinput_f53), .ZN(n6860) );
  OAI221_X1 U8611 ( .B1(SI_23_), .B2(keyinput_f9), .C1(P2_REG3_REG_9__SCAN_IN), 
        .C2(keyinput_f53), .A(n6860), .ZN(n6861) );
  NOR4_X1 U8612 ( .A1(n6864), .A2(n6863), .A3(n6862), .A4(n6861), .ZN(n6883)
         );
  AOI22_X1 U8613 ( .A1(SI_21_), .A2(keyinput_f11), .B1(P2_REG3_REG_4__SCAN_IN), 
        .B2(keyinput_f52), .ZN(n6865) );
  OAI221_X1 U8614 ( .B1(SI_21_), .B2(keyinput_f11), .C1(P2_REG3_REG_4__SCAN_IN), .C2(keyinput_f52), .A(n6865), .ZN(n6872) );
  AOI22_X1 U8615 ( .A1(SI_5_), .A2(keyinput_f27), .B1(SI_10_), .B2(
        keyinput_f22), .ZN(n6866) );
  OAI221_X1 U8616 ( .B1(SI_5_), .B2(keyinput_f27), .C1(SI_10_), .C2(
        keyinput_f22), .A(n6866), .ZN(n6871) );
  AOI22_X1 U8617 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(keyinput_f46), .B1(
        P2_REG3_REG_15__SCAN_IN), .B2(keyinput_f63), .ZN(n6867) );
  OAI221_X1 U8618 ( .B1(P2_REG3_REG_12__SCAN_IN), .B2(keyinput_f46), .C1(
        P2_REG3_REG_15__SCAN_IN), .C2(keyinput_f63), .A(n6867), .ZN(n6870) );
  AOI22_X1 U8619 ( .A1(SI_30_), .A2(keyinput_f2), .B1(SI_17_), .B2(
        keyinput_f15), .ZN(n6868) );
  OAI221_X1 U8620 ( .B1(SI_30_), .B2(keyinput_f2), .C1(SI_17_), .C2(
        keyinput_f15), .A(n6868), .ZN(n6869) );
  NOR4_X1 U8621 ( .A1(n6872), .A2(n6871), .A3(n6870), .A4(n6869), .ZN(n6882)
         );
  AOI22_X1 U8622 ( .A1(SI_14_), .A2(keyinput_f18), .B1(SI_25_), .B2(
        keyinput_f7), .ZN(n6873) );
  OAI221_X1 U8623 ( .B1(SI_14_), .B2(keyinput_f18), .C1(SI_25_), .C2(
        keyinput_f7), .A(n6873), .ZN(n6880) );
  AOI22_X1 U8624 ( .A1(P2_REG3_REG_1__SCAN_IN), .A2(keyinput_f44), .B1(
        P2_REG3_REG_27__SCAN_IN), .B2(keyinput_f36), .ZN(n6874) );
  OAI221_X1 U8625 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(keyinput_f44), .C1(
        P2_REG3_REG_27__SCAN_IN), .C2(keyinput_f36), .A(n6874), .ZN(n6879) );
  AOI22_X1 U8626 ( .A1(SI_31_), .A2(keyinput_f1), .B1(P2_REG3_REG_18__SCAN_IN), 
        .B2(keyinput_f60), .ZN(n6875) );
  OAI221_X1 U8627 ( .B1(SI_31_), .B2(keyinput_f1), .C1(P2_REG3_REG_18__SCAN_IN), .C2(keyinput_f60), .A(n6875), .ZN(n6878) );
  AOI22_X1 U8628 ( .A1(SI_29_), .A2(keyinput_f3), .B1(P2_REG3_REG_24__SCAN_IN), 
        .B2(keyinput_f51), .ZN(n6876) );
  OAI221_X1 U8629 ( .B1(SI_29_), .B2(keyinput_f3), .C1(P2_REG3_REG_24__SCAN_IN), .C2(keyinput_f51), .A(n6876), .ZN(n6877) );
  NOR4_X1 U8630 ( .A1(n6880), .A2(n6879), .A3(n6878), .A4(n6877), .ZN(n6881)
         );
  NAND4_X1 U8631 ( .A1(n6884), .A2(n6883), .A3(n6882), .A4(n6881), .ZN(n6933)
         );
  AOI22_X1 U8632 ( .A1(n6886), .A2(keyinput_f10), .B1(n4888), .B2(keyinput_f35), .ZN(n6885) );
  OAI221_X1 U8633 ( .B1(n6886), .B2(keyinput_f10), .C1(n4888), .C2(
        keyinput_f35), .A(n6885), .ZN(n6894) );
  INV_X1 U8634 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n6888) );
  AOI22_X1 U8635 ( .A1(n8539), .A2(keyinput_f50), .B1(n6888), .B2(keyinput_f45), .ZN(n6887) );
  OAI221_X1 U8636 ( .B1(n8539), .B2(keyinput_f50), .C1(n6888), .C2(
        keyinput_f45), .A(n6887), .ZN(n6893) );
  AOI22_X1 U8637 ( .A1(n6948), .A2(keyinput_f61), .B1(keyinput_f16), .B2(n6964), .ZN(n6889) );
  OAI221_X1 U8638 ( .B1(n6948), .B2(keyinput_f61), .C1(n6964), .C2(
        keyinput_f16), .A(n6889), .ZN(n6892) );
  INV_X1 U8639 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n7319) );
  AOI22_X1 U8640 ( .A1(n7319), .A2(keyinput_f37), .B1(keyinput_f17), .B2(n5301), .ZN(n6890) );
  OAI221_X1 U8641 ( .B1(n7319), .B2(keyinput_f37), .C1(n5301), .C2(
        keyinput_f17), .A(n6890), .ZN(n6891) );
  NOR4_X1 U8642 ( .A1(n6894), .A2(n6893), .A3(n6892), .A4(n6891), .ZN(n6931)
         );
  AOI22_X1 U8643 ( .A1(SI_28_), .A2(keyinput_f4), .B1(P2_REG3_REG_20__SCAN_IN), 
        .B2(keyinput_f55), .ZN(n6895) );
  OAI221_X1 U8644 ( .B1(SI_28_), .B2(keyinput_f4), .C1(P2_REG3_REG_20__SCAN_IN), .C2(keyinput_f55), .A(n6895), .ZN(n6903) );
  AOI22_X1 U8645 ( .A1(SI_19_), .A2(keyinput_f13), .B1(P2_REG3_REG_5__SCAN_IN), 
        .B2(keyinput_f49), .ZN(n6896) );
  OAI221_X1 U8646 ( .B1(SI_19_), .B2(keyinput_f13), .C1(P2_REG3_REG_5__SCAN_IN), .C2(keyinput_f49), .A(n6896), .ZN(n6902) );
  AOI22_X1 U8647 ( .A1(n6942), .A2(keyinput_f62), .B1(keyinput_f20), .B2(n6898), .ZN(n6897) );
  OAI221_X1 U8648 ( .B1(n6942), .B2(keyinput_f62), .C1(n6898), .C2(
        keyinput_f20), .A(n6897), .ZN(n6901) );
  INV_X1 U8649 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n6972) );
  AOI22_X1 U8650 ( .A1(n4441), .A2(keyinput_f43), .B1(n6972), .B2(keyinput_f42), .ZN(n6899) );
  OAI221_X1 U8651 ( .B1(n4441), .B2(keyinput_f43), .C1(n6972), .C2(
        keyinput_f42), .A(n6899), .ZN(n6900) );
  NOR4_X1 U8652 ( .A1(n6903), .A2(n6902), .A3(n6901), .A4(n6900), .ZN(n6930)
         );
  AOI22_X1 U8653 ( .A1(P2_U3151), .A2(keyinput_f34), .B1(keyinput_f33), .B2(
        n4927), .ZN(n6904) );
  OAI221_X1 U8654 ( .B1(P2_U3151), .B2(keyinput_f34), .C1(n4927), .C2(
        keyinput_f33), .A(n6904), .ZN(n6914) );
  AOI22_X1 U8655 ( .A1(n6907), .A2(keyinput_f8), .B1(keyinput_f21), .B2(n6906), 
        .ZN(n6905) );
  OAI221_X1 U8656 ( .B1(n6907), .B2(keyinput_f8), .C1(n6906), .C2(keyinput_f21), .A(n6905), .ZN(n6913) );
  XOR2_X1 U8657 ( .A(n4891), .B(keyinput_f56), .Z(n6911) );
  XNOR2_X1 U8658 ( .A(SI_4_), .B(keyinput_f28), .ZN(n6910) );
  XNOR2_X1 U8659 ( .A(SI_3_), .B(keyinput_f29), .ZN(n6909) );
  XNOR2_X1 U8660 ( .A(SI_1_), .B(keyinput_f31), .ZN(n6908) );
  NAND4_X1 U8661 ( .A1(n6911), .A2(n6910), .A3(n6909), .A4(n6908), .ZN(n6912)
         );
  NOR3_X1 U8662 ( .A1(n6914), .A2(n6913), .A3(n6912), .ZN(n6929) );
  INV_X1 U8663 ( .A(SI_13_), .ZN(n6916) );
  AOI22_X1 U8664 ( .A1(n6958), .A2(keyinput_f41), .B1(keyinput_f19), .B2(n6916), .ZN(n6915) );
  OAI221_X1 U8665 ( .B1(n6958), .B2(keyinput_f41), .C1(n6916), .C2(
        keyinput_f19), .A(n6915), .ZN(n6927) );
  INV_X1 U8666 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n8528) );
  AOI22_X1 U8667 ( .A1(n8528), .A2(keyinput_f47), .B1(keyinput_f5), .B2(n6918), 
        .ZN(n6917) );
  OAI221_X1 U8668 ( .B1(n8528), .B2(keyinput_f47), .C1(n6918), .C2(keyinput_f5), .A(n6917), .ZN(n6926) );
  INV_X1 U8669 ( .A(SI_18_), .ZN(n6920) );
  AOI22_X1 U8670 ( .A1(n6921), .A2(keyinput_f23), .B1(n6920), .B2(keyinput_f14), .ZN(n6919) );
  OAI221_X1 U8671 ( .B1(n6921), .B2(keyinput_f23), .C1(n6920), .C2(
        keyinput_f14), .A(n6919), .ZN(n6925) );
  XNOR2_X1 U8672 ( .A(P2_REG3_REG_2__SCAN_IN), .B(keyinput_f59), .ZN(n6923) );
  XNOR2_X1 U8673 ( .A(P2_REG3_REG_16__SCAN_IN), .B(keyinput_f48), .ZN(n6922)
         );
  NAND2_X1 U8674 ( .A1(n6923), .A2(n6922), .ZN(n6924) );
  NOR4_X1 U8675 ( .A1(n6927), .A2(n6926), .A3(n6925), .A4(n6924), .ZN(n6928)
         );
  NAND4_X1 U8676 ( .A1(n6931), .A2(n6930), .A3(n6929), .A4(n6928), .ZN(n6932)
         );
  OAI22_X1 U8677 ( .A1(keyinput_f26), .A2(n7028), .B1(n6933), .B2(n6932), .ZN(
        n6934) );
  AOI21_X1 U8678 ( .B1(keyinput_f26), .B2(n7028), .A(n6934), .ZN(n7027) );
  INV_X1 U8679 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n7673) );
  AOI22_X1 U8680 ( .A1(n6936), .A2(keyinput_g13), .B1(n7673), .B2(keyinput_g48), .ZN(n6935) );
  OAI221_X1 U8681 ( .B1(n6936), .B2(keyinput_g13), .C1(n7673), .C2(
        keyinput_g48), .A(n6935), .ZN(n6946) );
  AOI22_X1 U8682 ( .A1(n5301), .A2(keyinput_g17), .B1(n6938), .B2(keyinput_g4), 
        .ZN(n6937) );
  OAI221_X1 U8683 ( .B1(n5301), .B2(keyinput_g17), .C1(n6938), .C2(keyinput_g4), .A(n6937), .ZN(n6945) );
  AOI22_X1 U8684 ( .A1(n6940), .A2(keyinput_g7), .B1(n4927), .B2(keyinput_g33), 
        .ZN(n6939) );
  OAI221_X1 U8685 ( .B1(n6940), .B2(keyinput_g7), .C1(n4927), .C2(keyinput_g33), .A(n6939), .ZN(n6944) );
  INV_X1 U8686 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n7057) );
  AOI22_X1 U8687 ( .A1(n6942), .A2(keyinput_g62), .B1(keyinput_g58), .B2(n7057), .ZN(n6941) );
  OAI221_X1 U8688 ( .B1(n6942), .B2(keyinput_g62), .C1(n7057), .C2(
        keyinput_g58), .A(n6941), .ZN(n6943) );
  NOR4_X1 U8689 ( .A1(n6946), .A2(n6945), .A3(n6944), .A4(n6943), .ZN(n6987)
         );
  AOI22_X1 U8690 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(keyinput_g50), .B1(n6948), 
        .B2(keyinput_g61), .ZN(n6947) );
  OAI221_X1 U8691 ( .B1(P2_REG3_REG_17__SCAN_IN), .B2(keyinput_g50), .C1(n6948), .C2(keyinput_g61), .A(n6947), .ZN(n6956) );
  AOI22_X1 U8692 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(keyinput_g52), .B1(
        P2_STATE_REG_SCAN_IN), .B2(keyinput_g34), .ZN(n6949) );
  OAI221_X1 U8693 ( .B1(P2_REG3_REG_4__SCAN_IN), .B2(keyinput_g52), .C1(
        P2_STATE_REG_SCAN_IN), .C2(keyinput_g34), .A(n6949), .ZN(n6955) );
  AOI22_X1 U8694 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(keyinput_g49), .B1(
        P2_REG3_REG_12__SCAN_IN), .B2(keyinput_g46), .ZN(n6950) );
  OAI221_X1 U8695 ( .B1(P2_REG3_REG_5__SCAN_IN), .B2(keyinput_g49), .C1(
        P2_REG3_REG_12__SCAN_IN), .C2(keyinput_g46), .A(n6950), .ZN(n6954) );
  XNOR2_X1 U8696 ( .A(P2_REG3_REG_2__SCAN_IN), .B(keyinput_g59), .ZN(n6952) );
  XNOR2_X1 U8697 ( .A(P2_REG3_REG_24__SCAN_IN), .B(keyinput_g51), .ZN(n6951)
         );
  NAND2_X1 U8698 ( .A1(n6952), .A2(n6951), .ZN(n6953) );
  NOR4_X1 U8699 ( .A1(n6956), .A2(n6955), .A3(n6954), .A4(n6953), .ZN(n6986)
         );
  AOI22_X1 U8700 ( .A1(n6959), .A2(keyinput_g18), .B1(n6958), .B2(keyinput_g41), .ZN(n6957) );
  OAI221_X1 U8701 ( .B1(n6959), .B2(keyinput_g18), .C1(n6958), .C2(
        keyinput_g41), .A(n6957), .ZN(n6970) );
  INV_X1 U8702 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n6962) );
  INV_X1 U8703 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n6961) );
  AOI22_X1 U8704 ( .A1(n6962), .A2(keyinput_g57), .B1(n6961), .B2(keyinput_g38), .ZN(n6960) );
  OAI221_X1 U8705 ( .B1(n6962), .B2(keyinput_g57), .C1(n6961), .C2(
        keyinput_g38), .A(n6960), .ZN(n6969) );
  AOI22_X1 U8706 ( .A1(n6964), .A2(keyinput_g16), .B1(n4888), .B2(keyinput_g35), .ZN(n6963) );
  OAI221_X1 U8707 ( .B1(n6964), .B2(keyinput_g16), .C1(n4888), .C2(
        keyinput_g35), .A(n6963), .ZN(n6968) );
  AOI22_X1 U8708 ( .A1(n4889), .A2(keyinput_g53), .B1(keyinput_g15), .B2(n6966), .ZN(n6965) );
  OAI221_X1 U8709 ( .B1(n4889), .B2(keyinput_g53), .C1(n6966), .C2(
        keyinput_g15), .A(n6965), .ZN(n6967) );
  NOR4_X1 U8710 ( .A1(n6970), .A2(n6969), .A3(n6968), .A4(n6967), .ZN(n6985)
         );
  AOI22_X1 U8711 ( .A1(n6973), .A2(keyinput_g6), .B1(n6972), .B2(keyinput_g42), 
        .ZN(n6971) );
  OAI221_X1 U8712 ( .B1(n6973), .B2(keyinput_g6), .C1(n6972), .C2(keyinput_g42), .A(n6971), .ZN(n6983) );
  INV_X1 U8713 ( .A(SI_30_), .ZN(n6975) );
  AOI22_X1 U8714 ( .A1(n6976), .A2(keyinput_g36), .B1(keyinput_g2), .B2(n6975), 
        .ZN(n6974) );
  OAI221_X1 U8715 ( .B1(n6976), .B2(keyinput_g36), .C1(n6975), .C2(keyinput_g2), .A(n6974), .ZN(n6982) );
  INV_X1 U8716 ( .A(SI_31_), .ZN(n7618) );
  AOI22_X1 U8717 ( .A1(n4884), .A2(keyinput_g40), .B1(keyinput_g1), .B2(n7618), 
        .ZN(n6977) );
  OAI221_X1 U8718 ( .B1(n4884), .B2(keyinput_g40), .C1(n7618), .C2(keyinput_g1), .A(n6977), .ZN(n6981) );
  XNOR2_X1 U8719 ( .A(P2_REG3_REG_10__SCAN_IN), .B(keyinput_g39), .ZN(n6979)
         );
  XNOR2_X1 U8720 ( .A(SI_2_), .B(keyinput_g30), .ZN(n6978) );
  NAND2_X1 U8721 ( .A1(n6979), .A2(n6978), .ZN(n6980) );
  NOR4_X1 U8722 ( .A1(n6983), .A2(n6982), .A3(n6981), .A4(n6980), .ZN(n6984)
         );
  NAND4_X1 U8723 ( .A1(n6987), .A2(n6986), .A3(n6985), .A4(n6984), .ZN(n7025)
         );
  AOI22_X1 U8724 ( .A1(SI_0_), .A2(keyinput_g32), .B1(SI_21_), .B2(
        keyinput_g11), .ZN(n6988) );
  OAI221_X1 U8725 ( .B1(SI_0_), .B2(keyinput_g32), .C1(SI_21_), .C2(
        keyinput_g11), .A(n6988), .ZN(n6995) );
  AOI22_X1 U8726 ( .A1(SI_20_), .A2(keyinput_g12), .B1(SI_29_), .B2(
        keyinput_g3), .ZN(n6989) );
  OAI221_X1 U8727 ( .B1(SI_20_), .B2(keyinput_g12), .C1(SI_29_), .C2(
        keyinput_g3), .A(n6989), .ZN(n6994) );
  AOI22_X1 U8728 ( .A1(SI_8_), .A2(keyinput_g24), .B1(SI_23_), .B2(keyinput_g9), .ZN(n6990) );
  OAI221_X1 U8729 ( .B1(SI_8_), .B2(keyinput_g24), .C1(SI_23_), .C2(
        keyinput_g9), .A(n6990), .ZN(n6993) );
  AOI22_X1 U8730 ( .A1(SI_5_), .A2(keyinput_g27), .B1(SI_18_), .B2(
        keyinput_g14), .ZN(n6991) );
  OAI221_X1 U8731 ( .B1(SI_5_), .B2(keyinput_g27), .C1(SI_18_), .C2(
        keyinput_g14), .A(n6991), .ZN(n6992) );
  NOR4_X1 U8732 ( .A1(n6995), .A2(n6994), .A3(n6993), .A4(n6992), .ZN(n7023)
         );
  AOI22_X1 U8733 ( .A1(P2_REG3_REG_1__SCAN_IN), .A2(keyinput_g44), .B1(SI_9_), 
        .B2(keyinput_g23), .ZN(n6996) );
  OAI221_X1 U8734 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(keyinput_g44), .C1(SI_9_), 
        .C2(keyinput_g23), .A(n6996), .ZN(n7003) );
  AOI22_X1 U8735 ( .A1(SI_4_), .A2(keyinput_g28), .B1(P2_REG3_REG_14__SCAN_IN), 
        .B2(keyinput_g37), .ZN(n6997) );
  OAI221_X1 U8736 ( .B1(SI_4_), .B2(keyinput_g28), .C1(P2_REG3_REG_14__SCAN_IN), .C2(keyinput_g37), .A(n6997), .ZN(n7002) );
  AOI22_X1 U8737 ( .A1(SI_11_), .A2(keyinput_g21), .B1(P2_REG3_REG_13__SCAN_IN), .B2(keyinput_g56), .ZN(n6998) );
  OAI221_X1 U8738 ( .B1(SI_11_), .B2(keyinput_g21), .C1(
        P2_REG3_REG_13__SCAN_IN), .C2(keyinput_g56), .A(n6998), .ZN(n7001) );
  XNOR2_X1 U8739 ( .A(n6999), .B(keyinput_g29), .ZN(n7000) );
  NOR4_X1 U8740 ( .A1(n7003), .A2(n7002), .A3(n7001), .A4(n7000), .ZN(n7022)
         );
  AOI22_X1 U8741 ( .A1(P2_WR_REG_SCAN_IN), .A2(keyinput_g0), .B1(SI_27_), .B2(
        keyinput_g5), .ZN(n7004) );
  OAI221_X1 U8742 ( .B1(P2_WR_REG_SCAN_IN), .B2(keyinput_g0), .C1(SI_27_), 
        .C2(keyinput_g5), .A(n7004), .ZN(n7011) );
  AOI22_X1 U8743 ( .A1(SI_12_), .A2(keyinput_g20), .B1(SI_13_), .B2(
        keyinput_g19), .ZN(n7005) );
  OAI221_X1 U8744 ( .B1(SI_12_), .B2(keyinput_g20), .C1(SI_13_), .C2(
        keyinput_g19), .A(n7005), .ZN(n7010) );
  AOI22_X1 U8745 ( .A1(P2_REG3_REG_15__SCAN_IN), .A2(keyinput_g63), .B1(
        P2_REG3_REG_18__SCAN_IN), .B2(keyinput_g60), .ZN(n7006) );
  OAI221_X1 U8746 ( .B1(P2_REG3_REG_15__SCAN_IN), .B2(keyinput_g63), .C1(
        P2_REG3_REG_18__SCAN_IN), .C2(keyinput_g60), .A(n7006), .ZN(n7009) );
  AOI22_X1 U8747 ( .A1(SI_7_), .A2(keyinput_g25), .B1(P2_REG3_REG_21__SCAN_IN), 
        .B2(keyinput_g45), .ZN(n7007) );
  OAI221_X1 U8748 ( .B1(SI_7_), .B2(keyinput_g25), .C1(P2_REG3_REG_21__SCAN_IN), .C2(keyinput_g45), .A(n7007), .ZN(n7008) );
  NOR4_X1 U8749 ( .A1(n7011), .A2(n7010), .A3(n7009), .A4(n7008), .ZN(n7021)
         );
  AOI22_X1 U8750 ( .A1(SI_10_), .A2(keyinput_g22), .B1(SI_22_), .B2(
        keyinput_g10), .ZN(n7012) );
  OAI221_X1 U8751 ( .B1(SI_10_), .B2(keyinput_g22), .C1(SI_22_), .C2(
        keyinput_g10), .A(n7012), .ZN(n7019) );
  AOI22_X1 U8752 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(keyinput_g43), .B1(
        P2_REG3_REG_25__SCAN_IN), .B2(keyinput_g47), .ZN(n7013) );
  OAI221_X1 U8753 ( .B1(P2_REG3_REG_8__SCAN_IN), .B2(keyinput_g43), .C1(
        P2_REG3_REG_25__SCAN_IN), .C2(keyinput_g47), .A(n7013), .ZN(n7018) );
  AOI22_X1 U8754 ( .A1(SI_1_), .A2(keyinput_g31), .B1(SI_24_), .B2(keyinput_g8), .ZN(n7014) );
  OAI221_X1 U8755 ( .B1(SI_1_), .B2(keyinput_g31), .C1(SI_24_), .C2(
        keyinput_g8), .A(n7014), .ZN(n7017) );
  AOI22_X1 U8756 ( .A1(P2_REG3_REG_0__SCAN_IN), .A2(keyinput_g54), .B1(
        P2_REG3_REG_20__SCAN_IN), .B2(keyinput_g55), .ZN(n7015) );
  OAI221_X1 U8757 ( .B1(P2_REG3_REG_0__SCAN_IN), .B2(keyinput_g54), .C1(
        P2_REG3_REG_20__SCAN_IN), .C2(keyinput_g55), .A(n7015), .ZN(n7016) );
  NOR4_X1 U8758 ( .A1(n7019), .A2(n7018), .A3(n7017), .A4(n7016), .ZN(n7020)
         );
  NAND4_X1 U8759 ( .A1(n7023), .A2(n7022), .A3(n7021), .A4(n7020), .ZN(n7024)
         );
  OAI22_X1 U8760 ( .A1(keyinput_g26), .A2(n7028), .B1(n7025), .B2(n7024), .ZN(
        n7026) );
  AOI211_X1 U8761 ( .C1(keyinput_g26), .C2(n7028), .A(n7027), .B(n7026), .ZN(
        n7048) );
  INV_X1 U8762 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n10142) );
  NOR2_X1 U8763 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n7029) );
  AOI21_X1 U8764 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n7029), .ZN(n10147) );
  NOR2_X1 U8765 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n7030) );
  AOI21_X1 U8766 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n7030), .ZN(n10150) );
  NOR2_X1 U8767 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n7031) );
  AOI21_X1 U8768 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n7031), .ZN(n10153) );
  NOR2_X1 U8769 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n7032) );
  AOI21_X1 U8770 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n7032), .ZN(n10156) );
  NOR2_X1 U8771 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n7033) );
  AOI21_X1 U8772 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n7033), .ZN(n10159) );
  NOR2_X1 U8773 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n7034) );
  AOI21_X1 U8774 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n7034), .ZN(n10162) );
  NOR2_X1 U8775 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n7035) );
  AOI21_X1 U8776 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n7035), .ZN(n10165) );
  NOR2_X1 U8777 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n7036) );
  AOI21_X1 U8778 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n7036), .ZN(n10168) );
  NOR2_X1 U8779 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n7037) );
  AOI21_X1 U8780 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(P2_ADDR_REG_9__SCAN_IN), 
        .A(n7037), .ZN(n10174) );
  NOR2_X1 U8781 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n7038) );
  AOI21_X1 U8782 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(P2_ADDR_REG_8__SCAN_IN), 
        .A(n7038), .ZN(n10177) );
  NOR2_X1 U8783 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n7039) );
  AOI21_X1 U8784 ( .B1(P1_ADDR_REG_7__SCAN_IN), .B2(P2_ADDR_REG_7__SCAN_IN), 
        .A(n7039), .ZN(n10180) );
  NOR2_X1 U8785 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(P1_ADDR_REG_6__SCAN_IN), 
        .ZN(n7040) );
  AOI21_X1 U8786 ( .B1(P1_ADDR_REG_6__SCAN_IN), .B2(P2_ADDR_REG_6__SCAN_IN), 
        .A(n7040), .ZN(n10183) );
  NOR2_X1 U8787 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(P2_ADDR_REG_5__SCAN_IN), 
        .ZN(n7041) );
  AOI21_X1 U8788 ( .B1(P2_ADDR_REG_5__SCAN_IN), .B2(P1_ADDR_REG_5__SCAN_IN), 
        .A(n7041), .ZN(n10186) );
  AND2_X1 U8789 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .ZN(n7042) );
  NOR2_X1 U8790 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(n7042), .ZN(n10137) );
  INV_X1 U8791 ( .A(n10137), .ZN(n10138) );
  INV_X1 U8792 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10140) );
  NAND3_X1 U8793 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(P1_ADDR_REG_0__SCAN_IN), 
        .A3(P2_ADDR_REG_0__SCAN_IN), .ZN(n10139) );
  NAND2_X1 U8794 ( .A1(n10140), .A2(n10139), .ZN(n10136) );
  NAND2_X1 U8795 ( .A1(n10138), .A2(n10136), .ZN(n10171) );
  NAND2_X1 U8796 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n7043) );
  OAI21_X1 U8797 ( .B1(P1_ADDR_REG_2__SCAN_IN), .B2(P2_ADDR_REG_2__SCAN_IN), 
        .A(n7043), .ZN(n10170) );
  NOR2_X1 U8798 ( .A1(n10171), .A2(n10170), .ZN(n10169) );
  AOI21_X1 U8799 ( .B1(P2_ADDR_REG_2__SCAN_IN), .B2(P1_ADDR_REG_2__SCAN_IN), 
        .A(n10169), .ZN(n10189) );
  NAND2_X1 U8800 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n7044) );
  OAI21_X1 U8801 ( .B1(P1_ADDR_REG_3__SCAN_IN), .B2(P2_ADDR_REG_3__SCAN_IN), 
        .A(n7044), .ZN(n10188) );
  NOR2_X1 U8802 ( .A1(n10189), .A2(n10188), .ZN(n10187) );
  AOI21_X1 U8803 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(P1_ADDR_REG_3__SCAN_IN), 
        .A(n10187), .ZN(n10192) );
  NOR2_X1 U8804 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n7045) );
  AOI21_X1 U8805 ( .B1(P2_ADDR_REG_4__SCAN_IN), .B2(P1_ADDR_REG_4__SCAN_IN), 
        .A(n7045), .ZN(n10191) );
  NAND2_X1 U8806 ( .A1(n10192), .A2(n10191), .ZN(n10190) );
  OAI21_X1 U8807 ( .B1(P1_ADDR_REG_4__SCAN_IN), .B2(P2_ADDR_REG_4__SCAN_IN), 
        .A(n10190), .ZN(n10185) );
  NAND2_X1 U8808 ( .A1(n10186), .A2(n10185), .ZN(n10184) );
  OAI21_X1 U8809 ( .B1(P1_ADDR_REG_5__SCAN_IN), .B2(P2_ADDR_REG_5__SCAN_IN), 
        .A(n10184), .ZN(n10182) );
  NAND2_X1 U8810 ( .A1(n10183), .A2(n10182), .ZN(n10181) );
  OAI21_X1 U8811 ( .B1(P2_ADDR_REG_6__SCAN_IN), .B2(P1_ADDR_REG_6__SCAN_IN), 
        .A(n10181), .ZN(n10179) );
  NAND2_X1 U8812 ( .A1(n10180), .A2(n10179), .ZN(n10178) );
  OAI21_X1 U8813 ( .B1(P2_ADDR_REG_7__SCAN_IN), .B2(P1_ADDR_REG_7__SCAN_IN), 
        .A(n10178), .ZN(n10176) );
  NAND2_X1 U8814 ( .A1(n10177), .A2(n10176), .ZN(n10175) );
  OAI21_X1 U8815 ( .B1(P2_ADDR_REG_8__SCAN_IN), .B2(P1_ADDR_REG_8__SCAN_IN), 
        .A(n10175), .ZN(n10173) );
  NAND2_X1 U8816 ( .A1(n10174), .A2(n10173), .ZN(n10172) );
  OAI21_X1 U8817 ( .B1(P2_ADDR_REG_9__SCAN_IN), .B2(P1_ADDR_REG_9__SCAN_IN), 
        .A(n10172), .ZN(n10167) );
  NAND2_X1 U8818 ( .A1(n10168), .A2(n10167), .ZN(n10166) );
  OAI21_X1 U8819 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n10166), .ZN(n10164) );
  NAND2_X1 U8820 ( .A1(n10165), .A2(n10164), .ZN(n10163) );
  OAI21_X1 U8821 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n10163), .ZN(n10161) );
  NAND2_X1 U8822 ( .A1(n10162), .A2(n10161), .ZN(n10160) );
  OAI21_X1 U8823 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10160), .ZN(n10158) );
  NAND2_X1 U8824 ( .A1(n10159), .A2(n10158), .ZN(n10157) );
  OAI21_X1 U8825 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n10157), .ZN(n10155) );
  NAND2_X1 U8826 ( .A1(n10156), .A2(n10155), .ZN(n10154) );
  OAI21_X1 U8827 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10154), .ZN(n10152) );
  NAND2_X1 U8828 ( .A1(n10153), .A2(n10152), .ZN(n10151) );
  OAI21_X1 U8829 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n10151), .ZN(n10149) );
  NAND2_X1 U8830 ( .A1(n10150), .A2(n10149), .ZN(n10148) );
  OAI21_X1 U8831 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n10148), .ZN(n10146) );
  NAND2_X1 U8832 ( .A1(n10147), .A2(n10146), .ZN(n10145) );
  OAI21_X1 U8833 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10145), .ZN(n10143) );
  NAND2_X1 U8834 ( .A1(n10142), .A2(n10143), .ZN(n7046) );
  NOR2_X1 U8835 ( .A1(n10142), .A2(n10143), .ZN(n10141) );
  AOI21_X1 U8836 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(n7046), .A(n10141), .ZN(
        n7047) );
  XOR2_X1 U8837 ( .A(n7048), .B(n7047), .Z(n7051) );
  XNOR2_X1 U8838 ( .A(n7049), .B(P1_ADDR_REG_19__SCAN_IN), .ZN(n7050) );
  XNOR2_X1 U8839 ( .A(n7051), .B(n7050), .ZN(ADD_1068_U4) );
  AOI21_X1 U8840 ( .B1(n7054), .B2(n7053), .A(n7052), .ZN(n7068) );
  OAI21_X1 U8841 ( .B1(P2_REG1_REG_11__SCAN_IN), .B2(n7056), .A(n7055), .ZN(
        n7066) );
  INV_X1 U8842 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n7060) );
  NOR2_X1 U8843 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7057), .ZN(n7475) );
  AOI21_X1 U8844 ( .B1(n10020), .B2(n7058), .A(n7475), .ZN(n7059) );
  OAI21_X1 U8845 ( .B1(n10033), .B2(n7060), .A(n7059), .ZN(n7065) );
  AOI21_X1 U8846 ( .B1(n5234), .B2(n7062), .A(n7061), .ZN(n7063) );
  NOR2_X1 U8847 ( .A1(n7063), .A2(n10024), .ZN(n7064) );
  AOI211_X1 U8848 ( .C1(n10017), .C2(n7066), .A(n7065), .B(n7064), .ZN(n7067)
         );
  OAI21_X1 U8849 ( .B1(n7068), .B2(n8671), .A(n7067), .ZN(P2_U3193) );
  INV_X1 U8850 ( .A(n7743), .ZN(n7071) );
  INV_X1 U8851 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7069) );
  OAI222_X1 U8852 ( .A1(P2_U3151), .A2(n7070), .B1(n8470), .B2(n7071), .C1(
        n7069), .C2(n8491), .ZN(P2_U3274) );
  INV_X1 U8853 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7744) );
  OAI222_X1 U8854 ( .A1(n7913), .A2(n7744), .B1(n7915), .B2(n7071), .C1(
        P1_U3086), .C2(n8405), .ZN(P1_U3334) );
  INV_X1 U8855 ( .A(n7072), .ZN(n7073) );
  AOI21_X1 U8856 ( .B1(n8143), .B2(n7074), .A(n7073), .ZN(n7075) );
  OAI222_X1 U8857 ( .A1(n10043), .A2(n7106), .B1(n10041), .B2(n7477), .C1(
        n8792), .C2(n7075), .ZN(n10100) );
  INV_X1 U8858 ( .A(n10100), .ZN(n7080) );
  OAI22_X1 U8859 ( .A1(n10050), .A2(n5823), .B1(n7107), .B2(n10038), .ZN(n7076) );
  AOI21_X1 U8860 ( .B1(n8816), .B2(n4480), .A(n7076), .ZN(n7079) );
  OR2_X1 U8861 ( .A1(n7077), .A2(n5208), .ZN(n10099) );
  NAND2_X1 U8862 ( .A1(n7077), .A2(n5208), .ZN(n10098) );
  NAND3_X1 U8863 ( .A1(n10099), .A2(n7399), .A3(n10098), .ZN(n7078) );
  OAI211_X1 U8864 ( .C1(n7080), .C2(n8797), .A(n7079), .B(n7078), .ZN(P2_U3224) );
  XNOR2_X1 U8865 ( .A(n7081), .B(n8596), .ZN(n7082) );
  XNOR2_X1 U8866 ( .A(n7083), .B(n7082), .ZN(n7090) );
  AOI21_X1 U8867 ( .B1(n8547), .B2(n8595), .A(n7084), .ZN(n7085) );
  OAI21_X1 U8868 ( .B1(n4835), .B2(n8530), .A(n7085), .ZN(n7088) );
  NOR2_X1 U8869 ( .A1(n8577), .A2(n7086), .ZN(n7087) );
  AOI211_X1 U8870 ( .C1(n10093), .C2(n9539), .A(n7088), .B(n7087), .ZN(n7089)
         );
  OAI21_X1 U8871 ( .B1(n7090), .B2(n9543), .A(n7089), .ZN(P2_U3161) );
  INV_X1 U8872 ( .A(n7093), .ZN(n8142) );
  XNOR2_X1 U8873 ( .A(n7091), .B(n8142), .ZN(n7092) );
  OAI222_X1 U8874 ( .A1(n10043), .A2(n4479), .B1(n10041), .B2(n7525), .C1(
        n8792), .C2(n7092), .ZN(n7210) );
  INV_X1 U8875 ( .A(n7210), .ZN(n7099) );
  NAND2_X1 U8876 ( .A1(n10099), .A2(n7967), .ZN(n7094) );
  XNOR2_X1 U8877 ( .A(n7094), .B(n7093), .ZN(n7211) );
  NOR2_X1 U8878 ( .A1(n8681), .A2(n7216), .ZN(n7097) );
  OAI22_X1 U8879 ( .A1(n10050), .A2(n7095), .B1(n7392), .B2(n10038), .ZN(n7096) );
  AOI211_X1 U8880 ( .C1(n7211), .C2(n7399), .A(n7097), .B(n7096), .ZN(n7098)
         );
  OAI21_X1 U8881 ( .B1(n7099), .B2(n8797), .A(n7098), .ZN(P2_U3223) );
  INV_X1 U8882 ( .A(n7762), .ZN(n7682) );
  INV_X1 U8883 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7100) );
  OAI222_X1 U8884 ( .A1(n7101), .A2(P2_U3151), .B1(n8494), .B2(n7682), .C1(
        n7100), .C2(n8491), .ZN(P2_U3273) );
  XNOR2_X1 U8885 ( .A(n7103), .B(n7102), .ZN(n7111) );
  AOI21_X1 U8886 ( .B1(n8547), .B2(n8594), .A(n7104), .ZN(n7105) );
  OAI21_X1 U8887 ( .B1(n7106), .B2(n8530), .A(n7105), .ZN(n7109) );
  NOR2_X1 U8888 ( .A1(n8577), .A2(n7107), .ZN(n7108) );
  AOI211_X1 U8889 ( .C1(n4480), .C2(n9539), .A(n7109), .B(n7108), .ZN(n7110)
         );
  OAI21_X1 U8890 ( .B1(n7111), .B2(n9543), .A(n7110), .ZN(P2_U3171) );
  INV_X1 U8891 ( .A(n7778), .ZN(n7114) );
  AOI21_X1 U8892 ( .B1(P1_DATAO_REG_23__SCAN_IN), .B2(n7628), .A(n7112), .ZN(
        n7113) );
  OAI21_X1 U8893 ( .B1(n7114), .B2(n8494), .A(n7113), .ZN(P2_U3272) );
  INV_X1 U8894 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n7779) );
  NAND2_X1 U8895 ( .A1(n7778), .A2(n7115), .ZN(n7116) );
  OAI211_X1 U8896 ( .C1(n7779), .C2(n7913), .A(n7116), .B(n8466), .ZN(P1_U3332) );
  XNOR2_X1 U8897 ( .A(n7117), .B(n7121), .ZN(n7118) );
  OAI222_X1 U8898 ( .A1(n10043), .A2(n7477), .B1(n10041), .B2(n8026), .C1(
        n8792), .C2(n7118), .ZN(n10105) );
  INV_X1 U8899 ( .A(n10105), .ZN(n7127) );
  AND2_X1 U8900 ( .A1(n7120), .A2(n7119), .ZN(n7122) );
  XNOR2_X1 U8901 ( .A(n7122), .B(n7121), .ZN(n10107) );
  INV_X1 U8902 ( .A(n7123), .ZN(n10104) );
  NOR2_X1 U8903 ( .A1(n8681), .A2(n10104), .ZN(n7125) );
  OAI22_X1 U8904 ( .A1(n10050), .A2(n5234), .B1(n7474), .B2(n10038), .ZN(n7124) );
  AOI211_X1 U8905 ( .C1(n10107), .C2(n7399), .A(n7125), .B(n7124), .ZN(n7126)
         );
  OAI21_X1 U8906 ( .B1(n7127), .B2(n8797), .A(n7126), .ZN(P2_U3222) );
  NAND2_X1 U8907 ( .A1(n7141), .A2(n7709), .ZN(n7129) );
  NAND2_X1 U8908 ( .A1(n9074), .A2(n7924), .ZN(n7128) );
  AND2_X1 U8909 ( .A1(n7129), .A2(n7128), .ZN(n7226) );
  NAND2_X1 U8910 ( .A1(n7141), .A2(n6252), .ZN(n7134) );
  NAND2_X1 U8911 ( .A1(n9074), .A2(n7709), .ZN(n7133) );
  NAND2_X1 U8912 ( .A1(n7134), .A2(n7133), .ZN(n7135) );
  XNOR2_X1 U8913 ( .A(n7135), .B(n7922), .ZN(n7331) );
  XNOR2_X1 U8914 ( .A(n7330), .B(n7331), .ZN(n7136) );
  NOR2_X1 U8915 ( .A1(n7136), .A2(n7225), .ZN(n7329) );
  AOI21_X1 U8916 ( .B1(n7225), .B2(n7136), .A(n7329), .ZN(n7143) );
  AOI22_X1 U8917 ( .A1(n9018), .A2(n7137), .B1(P1_REG3_REG_8__SCAN_IN), .B2(
        P1_U3086), .ZN(n7138) );
  OAI21_X1 U8918 ( .B1(n9021), .B2(n7139), .A(n7138), .ZN(n7140) );
  AOI21_X1 U8919 ( .B1(n7141), .B2(n9023), .A(n7140), .ZN(n7142) );
  OAI21_X1 U8920 ( .B1(n7143), .B2(n9036), .A(n7142), .ZN(P1_U3221) );
  NAND2_X1 U8921 ( .A1(n7144), .A2(n7777), .ZN(n7146) );
  AOI22_X1 U8922 ( .A1(n7714), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n7713), .B2(
        n9656), .ZN(n7145) );
  NAND2_X1 U8923 ( .A1(n7173), .A2(n9070), .ZN(n8236) );
  NAND2_X1 U8924 ( .A1(n7148), .A2(n7147), .ZN(n9743) );
  NAND2_X1 U8925 ( .A1(n9743), .A2(n8235), .ZN(n7275) );
  NAND2_X1 U8926 ( .A1(n7149), .A2(n7777), .ZN(n7151) );
  AOI22_X1 U8927 ( .A1(n7714), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n7713), .B2(
        n9098), .ZN(n7150) );
  NAND2_X1 U8928 ( .A1(n7151), .A2(n7150), .ZN(n7174) );
  INV_X1 U8929 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n7175) );
  OR2_X1 U8930 ( .A1(n8177), .A2(n9940), .ZN(n7152) );
  OAI21_X1 U8931 ( .B1(n7941), .B2(n7175), .A(n7152), .ZN(n7159) );
  AND2_X1 U8932 ( .A1(n7154), .A2(n7153), .ZN(n7155) );
  OR2_X1 U8933 ( .A1(n7155), .A2(n7162), .ZN(n7249) );
  INV_X1 U8934 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n7156) );
  OR2_X1 U8935 ( .A1(n8179), .A2(n7156), .ZN(n7157) );
  OAI21_X1 U8936 ( .B1(n6262), .B2(n7249), .A(n7157), .ZN(n7158) );
  INV_X1 U8937 ( .A(n9069), .ZN(n7363) );
  OR2_X1 U8938 ( .A1(n7174), .A2(n7363), .ZN(n8239) );
  NAND2_X1 U8939 ( .A1(n7174), .A2(n7363), .ZN(n8432) );
  INV_X1 U8940 ( .A(n8372), .ZN(n7274) );
  XNOR2_X1 U8941 ( .A(n7275), .B(n7274), .ZN(n7170) );
  OR2_X1 U8942 ( .A1(n9070), .A2(n9017), .ZN(n7169) );
  INV_X1 U8943 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n7161) );
  INV_X1 U8944 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n9096) );
  OR2_X1 U8945 ( .A1(n8177), .A2(n9096), .ZN(n7160) );
  OAI21_X1 U8946 ( .B1(n7941), .B2(n7161), .A(n7160), .ZN(n7167) );
  OR2_X1 U8947 ( .A1(n7162), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n7163) );
  NAND2_X1 U8948 ( .A1(n7263), .A2(n7163), .ZN(n9732) );
  INV_X1 U8949 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n7164) );
  OR2_X1 U8950 ( .A1(n8179), .A2(n7164), .ZN(n7165) );
  OAI21_X1 U8951 ( .B1(n6262), .B2(n9732), .A(n7165), .ZN(n7166) );
  NAND2_X1 U8952 ( .A1(n9068), .A2(n9052), .ZN(n7168) );
  NAND2_X1 U8953 ( .A1(n7169), .A2(n7168), .ZN(n7246) );
  AOI21_X1 U8954 ( .B1(n7170), .B2(n9821), .A(n7246), .ZN(n9905) );
  INV_X1 U8955 ( .A(n7376), .ZN(n9072) );
  INV_X1 U8956 ( .A(n7173), .ZN(n9898) );
  XNOR2_X1 U8957 ( .A(n7253), .B(n8372), .ZN(n9908) );
  NAND2_X1 U8958 ( .A1(n9908), .A2(n9809), .ZN(n7180) );
  OAI22_X1 U8959 ( .A1(n9335), .A2(n7175), .B1(n7249), .B2(n9799), .ZN(n7178)
         );
  INV_X1 U8960 ( .A(n7174), .ZN(n9906) );
  INV_X1 U8961 ( .A(n7270), .ZN(n7176) );
  OAI211_X1 U8962 ( .C1(n9906), .C2(n9756), .A(n7176), .B(n9829), .ZN(n9904)
         );
  NOR2_X1 U8963 ( .A1(n9904), .A2(n9248), .ZN(n7177) );
  AOI211_X1 U8964 ( .C1(n9753), .C2(n7174), .A(n7178), .B(n7177), .ZN(n7179)
         );
  OAI211_X1 U8965 ( .C1(n9836), .C2(n9905), .A(n7180), .B(n7179), .ZN(P1_U3281) );
  AOI21_X1 U8966 ( .B1(n5280), .B2(n7182), .A(n7181), .ZN(n7196) );
  OAI21_X1 U8967 ( .B1(P2_REG1_REG_13__SCAN_IN), .B2(n7184), .A(n7183), .ZN(
        n7194) );
  INV_X1 U8968 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n7192) );
  OAI21_X1 U8969 ( .B1(n7187), .B2(n7186), .A(n7185), .ZN(n7190) );
  NOR2_X1 U8970 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n4891), .ZN(n7463) );
  NOR2_X1 U8971 ( .A1(n9956), .A2(n7188), .ZN(n7189) );
  AOI211_X1 U8972 ( .C1(n10029), .C2(n7190), .A(n7463), .B(n7189), .ZN(n7191)
         );
  OAI21_X1 U8973 ( .B1(n10033), .B2(n7192), .A(n7191), .ZN(n7193) );
  AOI21_X1 U8974 ( .B1(n7194), .B2(n10017), .A(n7193), .ZN(n7195) );
  OAI21_X1 U8975 ( .B1(n7196), .B2(n10024), .A(n7195), .ZN(P2_U3195) );
  OR2_X1 U8976 ( .A1(n7117), .A2(n7197), .ZN(n7199) );
  NAND2_X1 U8977 ( .A1(n7199), .A2(n7198), .ZN(n7200) );
  XNOR2_X1 U8978 ( .A(n7200), .B(n5265), .ZN(n7201) );
  NAND2_X1 U8979 ( .A1(n7201), .A2(n5513), .ZN(n7203) );
  AOI22_X1 U8980 ( .A1(n8807), .A2(n8593), .B1(n8591), .B2(n8809), .ZN(n7202)
         );
  NAND2_X1 U8981 ( .A1(n7203), .A2(n7202), .ZN(n10117) );
  INV_X1 U8982 ( .A(n10117), .ZN(n7209) );
  OAI22_X1 U8983 ( .A1(n10050), .A2(n7204), .B1(n7532), .B2(n10038), .ZN(n7205) );
  AOI21_X1 U8984 ( .B1(n8816), .B2(n10113), .A(n7205), .ZN(n7208) );
  NAND2_X1 U8985 ( .A1(n7206), .A2(n8030), .ZN(n10109) );
  NAND3_X1 U8986 ( .A1(n10111), .A2(n10109), .A3(n7399), .ZN(n7207) );
  OAI211_X1 U8987 ( .C1(n7209), .C2(n8797), .A(n7208), .B(n7207), .ZN(P2_U3221) );
  AOI21_X1 U8988 ( .B1(n10110), .B2(n7211), .A(n7210), .ZN(n7213) );
  MUX2_X1 U8989 ( .A(n5829), .B(n7213), .S(n10135), .Z(n7212) );
  OAI21_X1 U8990 ( .B1(n7216), .B2(n8836), .A(n7212), .ZN(P2_U3469) );
  INV_X1 U8991 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n7214) );
  MUX2_X1 U8992 ( .A(n7214), .B(n7213), .S(n10118), .Z(n7215) );
  OAI21_X1 U8993 ( .B1(n7216), .B2(n8892), .A(n7215), .ZN(P2_U3420) );
  INV_X1 U8994 ( .A(n7916), .ZN(n7837) );
  AOI21_X1 U8995 ( .B1(n7628), .B2(P1_DATAO_REG_27__SCAN_IN), .A(n7217), .ZN(
        n7218) );
  OAI21_X1 U8996 ( .B1(n7837), .B2(n8494), .A(n7218), .ZN(P2_U3268) );
  INV_X1 U8997 ( .A(n7846), .ZN(n8469) );
  INV_X1 U8998 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7847) );
  OAI222_X1 U8999 ( .A1(n7915), .A2(n8469), .B1(P1_U3086), .B2(n7219), .C1(
        n7847), .C2(n7913), .ZN(P1_U3331) );
  NAND2_X1 U9000 ( .A1(n7338), .A2(n6252), .ZN(n7221) );
  NAND2_X1 U9001 ( .A1(n9073), .A2(n7709), .ZN(n7220) );
  NAND2_X1 U9002 ( .A1(n7221), .A2(n7220), .ZN(n7222) );
  XNOR2_X1 U9003 ( .A(n7222), .B(n7949), .ZN(n7333) );
  OAI22_X1 U9004 ( .A1(n9888), .A2(n7948), .B1(n7223), .B2(n6158), .ZN(n7332)
         );
  INV_X1 U9005 ( .A(n7331), .ZN(n7224) );
  AOI22_X1 U9006 ( .A1(n7333), .A2(n7332), .B1(n7225), .B2(n7224), .ZN(n7230)
         );
  NOR3_X1 U9007 ( .A1(n7332), .A2(n7225), .A3(n7224), .ZN(n7229) );
  NAND2_X1 U9008 ( .A1(n7331), .A2(n7226), .ZN(n7227) );
  AOI21_X1 U9009 ( .B1(n7332), .B2(n7227), .A(n7333), .ZN(n7228) );
  NAND2_X1 U9010 ( .A1(n7173), .A2(n4346), .ZN(n7232) );
  OR2_X1 U9011 ( .A1(n9070), .A2(n7948), .ZN(n7231) );
  NAND2_X1 U9012 ( .A1(n7232), .A2(n7231), .ZN(n7233) );
  XNOR2_X1 U9013 ( .A(n7233), .B(n7922), .ZN(n7373) );
  NOR2_X1 U9014 ( .A1(n9070), .A2(n6158), .ZN(n7234) );
  AOI21_X1 U9015 ( .B1(n7173), .B2(n7709), .A(n7234), .ZN(n7372) );
  NOR2_X1 U9016 ( .A1(n7376), .A2(n6158), .ZN(n7235) );
  AOI21_X1 U9017 ( .B1(n7299), .B2(n7709), .A(n7235), .ZN(n7297) );
  NAND2_X1 U9018 ( .A1(n7299), .A2(n6252), .ZN(n7237) );
  OR2_X1 U9019 ( .A1(n7376), .A2(n7948), .ZN(n7236) );
  NAND2_X1 U9020 ( .A1(n7237), .A2(n7236), .ZN(n7238) );
  XNOR2_X1 U9021 ( .A(n7238), .B(n7922), .ZN(n7368) );
  OAI22_X1 U9022 ( .A1(n7373), .A2(n7372), .B1(n7297), .B2(n7368), .ZN(n7242)
         );
  AND2_X1 U9023 ( .A1(n7368), .A2(n7297), .ZN(n7240) );
  OAI21_X1 U9024 ( .B1(n7240), .B2(n7372), .A(n7373), .ZN(n7239) );
  INV_X1 U9025 ( .A(n7239), .ZN(n7241) );
  OAI22_X1 U9026 ( .A1(n9906), .A2(n7948), .B1(n7363), .B2(n6158), .ZN(n7354)
         );
  NAND2_X1 U9027 ( .A1(n7174), .A2(n6252), .ZN(n7244) );
  NAND2_X1 U9028 ( .A1(n9069), .A2(n7709), .ZN(n7243) );
  NAND2_X1 U9029 ( .A1(n7244), .A2(n7243), .ZN(n7245) );
  XNOR2_X1 U9030 ( .A(n7245), .B(n7949), .ZN(n7353) );
  XOR2_X1 U9031 ( .A(n7354), .B(n7353), .Z(n7357) );
  XOR2_X1 U9032 ( .A(n7358), .B(n7357), .Z(n7252) );
  NAND2_X1 U9033 ( .A1(n9018), .A2(n7246), .ZN(n7247) );
  OAI211_X1 U9034 ( .C1(n9021), .C2(n7249), .A(n7248), .B(n7247), .ZN(n7250)
         );
  AOI21_X1 U9035 ( .B1(n7174), .B2(n9023), .A(n7250), .ZN(n7251) );
  OAI21_X1 U9036 ( .B1(n7252), .B2(n9036), .A(n7251), .ZN(P1_U3224) );
  NAND2_X1 U9037 ( .A1(n7254), .A2(n7777), .ZN(n7256) );
  AOI22_X1 U9038 ( .A1(n7714), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n7713), .B2(
        n9680), .ZN(n7255) );
  NAND2_X1 U9039 ( .A1(n7256), .A2(n7255), .ZN(n9734) );
  NAND2_X1 U9040 ( .A1(n9734), .A2(n7362), .ZN(n8248) );
  NAND2_X1 U9041 ( .A1(n8247), .A2(n8248), .ZN(n9735) );
  NAND2_X1 U9042 ( .A1(n7257), .A2(n7777), .ZN(n7259) );
  AOI22_X1 U9043 ( .A1(n7714), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n7713), .B2(
        n9113), .ZN(n7258) );
  INV_X1 U9044 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n7271) );
  INV_X1 U9045 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n7260) );
  OR2_X1 U9046 ( .A1(n8177), .A2(n7260), .ZN(n7261) );
  OAI21_X1 U9047 ( .B1(n7941), .B2(n7271), .A(n7261), .ZN(n7268) );
  NAND2_X1 U9048 ( .A1(n7263), .A2(n7262), .ZN(n7264) );
  NAND2_X1 U9049 ( .A1(n7283), .A2(n7264), .ZN(n7562) );
  INV_X1 U9050 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n7265) );
  OR2_X1 U9051 ( .A1(n8179), .A2(n7265), .ZN(n7266) );
  OAI21_X1 U9052 ( .B1(n6262), .B2(n7562), .A(n7266), .ZN(n7267) );
  INV_X1 U9053 ( .A(n9067), .ZN(n7556) );
  OR2_X1 U9054 ( .A1(n9918), .A2(n7556), .ZN(n8252) );
  INV_X1 U9055 ( .A(n9549), .ZN(n7269) );
  XNOR2_X1 U9056 ( .A(n7422), .B(n7277), .ZN(n9922) );
  AOI211_X1 U9057 ( .C1(n9918), .C2(n9737), .A(n9775), .B(n4423), .ZN(n9917)
         );
  INV_X1 U9058 ( .A(n9918), .ZN(n7557) );
  NOR2_X1 U9059 ( .A1(n7557), .A2(n9825), .ZN(n7273) );
  OAI22_X1 U9060 ( .A1(n9335), .A2(n7271), .B1(n7562), .B2(n9799), .ZN(n7272)
         );
  AOI211_X1 U9061 ( .C1(n9917), .C2(n9832), .A(n7273), .B(n7272), .ZN(n7293)
         );
  OAI21_X2 U9062 ( .B1(n7275), .B2(n7274), .A(n8432), .ZN(n9729) );
  AOI21_X1 U9063 ( .B1(n7277), .B2(n7276), .A(n9550), .ZN(n7291) );
  INV_X1 U9064 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n7278) );
  OR2_X1 U9065 ( .A1(n8179), .A2(n7278), .ZN(n7281) );
  INV_X1 U9066 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n7279) );
  OR2_X1 U9067 ( .A1(n8177), .A2(n7279), .ZN(n7280) );
  AND2_X1 U9068 ( .A1(n7281), .A2(n7280), .ZN(n7287) );
  AND2_X1 U9069 ( .A1(n7283), .A2(n9055), .ZN(n7284) );
  NOR2_X1 U9070 ( .A1(n7436), .A2(n7284), .ZN(n9555) );
  NAND2_X1 U9071 ( .A1(n7876), .A2(n9555), .ZN(n7286) );
  NAND2_X1 U9072 ( .A1(n7731), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n7285) );
  OR2_X1 U9073 ( .A1(n7686), .A2(n9162), .ZN(n7289) );
  NAND2_X1 U9074 ( .A1(n9068), .A2(n9225), .ZN(n7288) );
  NAND2_X1 U9075 ( .A1(n7289), .A2(n7288), .ZN(n7560) );
  INV_X1 U9076 ( .A(n7560), .ZN(n7290) );
  OAI21_X1 U9077 ( .B1(n7291), .B2(n9746), .A(n7290), .ZN(n9916) );
  NAND2_X1 U9078 ( .A1(n9916), .A2(n9335), .ZN(n7292) );
  OAI211_X1 U9079 ( .C1(n9922), .C2(n9378), .A(n7293), .B(n7292), .ZN(P1_U3279) );
  INV_X1 U9080 ( .A(n7838), .ZN(n7308) );
  AOI22_X1 U9081 ( .A1(n7294), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_26__SCAN_IN), .B2(n7628), .ZN(n7295) );
  OAI21_X1 U9082 ( .B1(n7308), .B2(n8494), .A(n7295), .ZN(P2_U3269) );
  XNOR2_X1 U9083 ( .A(n7371), .B(n7368), .ZN(n7296) );
  NAND2_X1 U9084 ( .A1(n7296), .A2(n7297), .ZN(n7369) );
  OAI21_X1 U9085 ( .B1(n7297), .B2(n7296), .A(n7369), .ZN(n7304) );
  AOI22_X1 U9086 ( .A1(n9018), .A2(n7298), .B1(P1_REG3_REG_10__SCAN_IN), .B2(
        P1_U3086), .ZN(n7301) );
  NAND2_X1 U9087 ( .A1(n7299), .A2(n9023), .ZN(n7300) );
  OAI211_X1 U9088 ( .C1(n9021), .C2(n7302), .A(n7301), .B(n7300), .ZN(n7303)
         );
  AOI21_X1 U9089 ( .B1(n7304), .B2(n9050), .A(n7303), .ZN(n7305) );
  INV_X1 U9090 ( .A(n7305), .ZN(P1_U3217) );
  INV_X1 U9091 ( .A(n7853), .ZN(n8493) );
  INV_X1 U9092 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7854) );
  OAI222_X1 U9093 ( .A1(n7915), .A2(n8493), .B1(P1_U3086), .B2(n7306), .C1(
        n7854), .C2(n7913), .ZN(P1_U3330) );
  INV_X1 U9094 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n7839) );
  OAI222_X1 U9095 ( .A1(n7915), .A2(n7308), .B1(P1_U3086), .B2(n7307), .C1(
        n7839), .C2(n7913), .ZN(P1_U3329) );
  INV_X1 U9096 ( .A(n7934), .ZN(n7914) );
  NAND2_X1 U9097 ( .A1(n7628), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n7309) );
  OAI211_X1 U9098 ( .C1(n7914), .C2(n8494), .A(n7310), .B(n7309), .ZN(P2_U3267) );
  AOI21_X1 U9099 ( .B1(n4416), .B2(n7312), .A(n7311), .ZN(n7328) );
  OAI21_X1 U9100 ( .B1(n7315), .B2(n7314), .A(n7313), .ZN(n7326) );
  INV_X1 U9101 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n7324) );
  OAI21_X1 U9102 ( .B1(n7318), .B2(n7317), .A(n7316), .ZN(n7322) );
  NOR2_X1 U9103 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7319), .ZN(n7541) );
  NOR2_X1 U9104 ( .A1(n9956), .A2(n7320), .ZN(n7321) );
  AOI211_X1 U9105 ( .C1(n10029), .C2(n7322), .A(n7541), .B(n7321), .ZN(n7323)
         );
  OAI21_X1 U9106 ( .B1(n10033), .B2(n7324), .A(n7323), .ZN(n7325) );
  AOI21_X1 U9107 ( .B1(n7326), .B2(n10017), .A(n7325), .ZN(n7327) );
  OAI21_X1 U9108 ( .B1(n7328), .B2(n10024), .A(n7327), .ZN(P2_U3196) );
  AOI21_X1 U9109 ( .B1(n7331), .B2(n7330), .A(n7329), .ZN(n7335) );
  XNOR2_X1 U9110 ( .A(n7333), .B(n7332), .ZN(n7334) );
  XNOR2_X1 U9111 ( .A(n7335), .B(n7334), .ZN(n7343) );
  NAND2_X1 U9112 ( .A1(n7337), .A2(n7336), .ZN(n9885) );
  AND2_X1 U9113 ( .A1(P1_U3086), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n9086) );
  AOI21_X1 U9114 ( .B1(n9018), .B2(n9885), .A(n9086), .ZN(n7340) );
  NAND2_X1 U9115 ( .A1(n7338), .A2(n9023), .ZN(n7339) );
  OAI211_X1 U9116 ( .C1(n9021), .C2(n7341), .A(n7340), .B(n7339), .ZN(n7342)
         );
  AOI21_X1 U9117 ( .B1(n7343), .B2(n9050), .A(n7342), .ZN(n7344) );
  INV_X1 U9118 ( .A(n7344), .ZN(P1_U3231) );
  INV_X1 U9119 ( .A(n10036), .ZN(n8718) );
  NAND2_X1 U9120 ( .A1(n7347), .A2(n7346), .ZN(n8034) );
  XNOR2_X1 U9121 ( .A(n7345), .B(n4493), .ZN(n7348) );
  OAI222_X1 U9122 ( .A1(n10041), .A2(n7609), .B1(n10043), .B2(n8026), .C1(
        n8792), .C2(n7348), .ZN(n7411) );
  AOI21_X1 U9123 ( .B1(n8718), .B2(n7467), .A(n7411), .ZN(n7352) );
  XNOR2_X1 U9124 ( .A(n7349), .B(n4493), .ZN(n7418) );
  OAI22_X1 U9125 ( .A1(n10050), .A2(n5280), .B1(n7465), .B2(n10038), .ZN(n7350) );
  AOI21_X1 U9126 ( .B1(n7418), .B2(n7399), .A(n7350), .ZN(n7351) );
  OAI21_X1 U9127 ( .B1(n7352), .B2(n8797), .A(n7351), .ZN(P2_U3220) );
  INV_X1 U9128 ( .A(n7353), .ZN(n7356) );
  INV_X1 U9129 ( .A(n7354), .ZN(n7355) );
  NAND2_X1 U9130 ( .A1(n9734), .A2(n6252), .ZN(n7360) );
  NAND2_X1 U9131 ( .A1(n9068), .A2(n7709), .ZN(n7359) );
  NAND2_X1 U9132 ( .A1(n7360), .A2(n7359), .ZN(n7361) );
  XNOR2_X1 U9133 ( .A(n7361), .B(n7949), .ZN(n7549) );
  OAI22_X1 U9134 ( .A1(n9912), .A2(n7948), .B1(n7362), .B2(n6158), .ZN(n7548)
         );
  XNOR2_X1 U9135 ( .A(n7549), .B(n7548), .ZN(n7551) );
  XOR2_X1 U9136 ( .A(n7552), .B(n7551), .Z(n7367) );
  OAI22_X1 U9137 ( .A1(n7363), .A2(n9017), .B1(n7556), .B2(n9162), .ZN(n9730)
         );
  AOI22_X1 U9138 ( .A1(n9018), .A2(n9730), .B1(P1_REG3_REG_13__SCAN_IN), .B2(
        P1_U3086), .ZN(n7364) );
  OAI21_X1 U9139 ( .B1(n9021), .B2(n9732), .A(n7364), .ZN(n7365) );
  AOI21_X1 U9140 ( .B1(n9734), .B2(n9023), .A(n7365), .ZN(n7366) );
  OAI21_X1 U9141 ( .B1(n7367), .B2(n9036), .A(n7366), .ZN(P1_U3234) );
  INV_X1 U9142 ( .A(n7368), .ZN(n7370) );
  OAI21_X1 U9143 ( .B1(n7371), .B2(n7370), .A(n7369), .ZN(n7375) );
  XNOR2_X1 U9144 ( .A(n7373), .B(n7372), .ZN(n7374) );
  XNOR2_X1 U9145 ( .A(n7375), .B(n7374), .ZN(n7382) );
  OR2_X1 U9146 ( .A1(n7376), .A2(n9017), .ZN(n7378) );
  NAND2_X1 U9147 ( .A1(n9069), .A2(n9052), .ZN(n7377) );
  NAND2_X1 U9148 ( .A1(n7378), .A2(n7377), .ZN(n9749) );
  AOI22_X1 U9149 ( .A1(n9018), .A2(n9749), .B1(P1_REG3_REG_11__SCAN_IN), .B2(
        P1_U3086), .ZN(n7379) );
  OAI21_X1 U9150 ( .B1(n9021), .B2(n9751), .A(n7379), .ZN(n7380) );
  AOI21_X1 U9151 ( .B1(n7173), .B2(n9023), .A(n7380), .ZN(n7381) );
  OAI21_X1 U9152 ( .B1(n7382), .B2(n9036), .A(n7381), .ZN(P1_U3236) );
  XNOR2_X1 U9153 ( .A(n7470), .B(n8594), .ZN(n7384) );
  NAND2_X1 U9154 ( .A1(n7384), .A2(n7383), .ZN(n7472) );
  OAI21_X1 U9155 ( .B1(n7384), .B2(n7383), .A(n7472), .ZN(n7385) );
  NAND2_X1 U9156 ( .A1(n7385), .A2(n8572), .ZN(n7391) );
  AOI21_X1 U9157 ( .B1(n8547), .B2(n8593), .A(n7386), .ZN(n7387) );
  OAI21_X1 U9158 ( .B1(n4479), .B2(n8530), .A(n7387), .ZN(n7388) );
  AOI21_X1 U9159 ( .B1(n7389), .B2(n9539), .A(n7388), .ZN(n7390) );
  OAI211_X1 U9160 ( .C1(n7392), .C2(n8577), .A(n7391), .B(n7390), .ZN(P2_U3157) );
  INV_X1 U9161 ( .A(n8037), .ZN(n7394) );
  OR2_X1 U9162 ( .A1(n8035), .A2(n7394), .ZN(n8146) );
  XOR2_X1 U9163 ( .A(n7393), .B(n8146), .Z(n7395) );
  AOI222_X1 U9164 ( .A1(n5513), .A2(n7395), .B1(n8589), .B2(n8809), .C1(n8591), 
        .C2(n8807), .ZN(n7405) );
  INV_X1 U9165 ( .A(n7405), .ZN(n7397) );
  INV_X1 U9166 ( .A(n7407), .ZN(n7547) );
  OAI22_X1 U9167 ( .A1(n7547), .A2(n10036), .B1(n7540), .B2(n10038), .ZN(n7396) );
  OAI21_X1 U9168 ( .B1(n7397), .B2(n7396), .A(n10050), .ZN(n7401) );
  XNOR2_X1 U9169 ( .A(n7398), .B(n8146), .ZN(n7408) );
  AOI22_X1 U9170 ( .A1(n7408), .A2(n7399), .B1(P2_REG2_REG_14__SCAN_IN), .B2(
        n8797), .ZN(n7400) );
  NAND2_X1 U9171 ( .A1(n7401), .A2(n7400), .ZN(P2_U3219) );
  INV_X1 U9172 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n7402) );
  MUX2_X1 U9173 ( .A(n7402), .B(n7405), .S(n10118), .Z(n7404) );
  INV_X1 U9174 ( .A(n8931), .ZN(n7417) );
  AOI22_X1 U9175 ( .A1(n7408), .A2(n7417), .B1(n8927), .B2(n7407), .ZN(n7403)
         );
  NAND2_X1 U9176 ( .A1(n7404), .A2(n7403), .ZN(P2_U3432) );
  MUX2_X1 U9177 ( .A(n7406), .B(n7405), .S(n10135), .Z(n7410) );
  INV_X1 U9178 ( .A(n8859), .ZN(n7412) );
  AOI22_X1 U9179 ( .A1(n7408), .A2(n7412), .B1(n8856), .B2(n7407), .ZN(n7409)
         );
  NAND2_X1 U9180 ( .A1(n7410), .A2(n7409), .ZN(P2_U3473) );
  INV_X1 U9181 ( .A(n7411), .ZN(n7415) );
  MUX2_X1 U9182 ( .A(n5277), .B(n7415), .S(n10135), .Z(n7414) );
  AOI22_X1 U9183 ( .A1(n7418), .A2(n7412), .B1(n8856), .B2(n7467), .ZN(n7413)
         );
  NAND2_X1 U9184 ( .A1(n7414), .A2(n7413), .ZN(P2_U3472) );
  INV_X1 U9185 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n7416) );
  MUX2_X1 U9186 ( .A(n7416), .B(n7415), .S(n10118), .Z(n7420) );
  AOI22_X1 U9187 ( .A1(n7418), .A2(n7417), .B1(n8927), .B2(n7467), .ZN(n7419)
         );
  NAND2_X1 U9188 ( .A1(n7420), .A2(n7419), .ZN(P2_U3429) );
  NAND2_X1 U9189 ( .A1(n7557), .A2(n7556), .ZN(n7421) );
  NAND2_X1 U9190 ( .A1(n7423), .A2(n7777), .ZN(n7425) );
  INV_X1 U9191 ( .A(n9115), .ZN(n9708) );
  AOI22_X1 U9192 ( .A1(n7714), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n7713), .B2(
        n9708), .ZN(n7424) );
  INV_X1 U9193 ( .A(n7686), .ZN(n9066) );
  NAND2_X1 U9194 ( .A1(n9557), .A2(n7426), .ZN(n7429) );
  OR2_X1 U9195 ( .A1(n7446), .A2(n7686), .ZN(n7428) );
  NAND2_X1 U9196 ( .A1(n7429), .A2(n7428), .ZN(n7500) );
  NAND2_X1 U9197 ( .A1(n7430), .A2(n7777), .ZN(n7432) );
  AOI22_X1 U9198 ( .A1(n7714), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n7713), .B2(
        n9128), .ZN(n7431) );
  INV_X1 U9199 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n7435) );
  INV_X1 U9200 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n7433) );
  OR2_X1 U9201 ( .A1(n8177), .A2(n7433), .ZN(n7434) );
  OAI21_X1 U9202 ( .B1(n7941), .B2(n7435), .A(n7434), .ZN(n7441) );
  AND2_X2 U9203 ( .A1(n7436), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n8992) );
  NOR2_X1 U9204 ( .A1(n7436), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n7437) );
  OR2_X1 U9205 ( .A1(n8992), .A2(n7437), .ZN(n8985) );
  INV_X1 U9206 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n7438) );
  OR2_X1 U9207 ( .A1(n8179), .A2(n7438), .ZN(n7439) );
  OAI21_X1 U9208 ( .B1(n6262), .B2(n8985), .A(n7439), .ZN(n7440) );
  INV_X1 U9209 ( .A(n9065), .ZN(n7442) );
  NAND2_X1 U9210 ( .A1(n9454), .A2(n7442), .ZN(n8435) );
  NAND2_X1 U9211 ( .A1(n8256), .A2(n8435), .ZN(n8375) );
  XNOR2_X1 U9212 ( .A(n7500), .B(n8375), .ZN(n9458) );
  AOI211_X1 U9213 ( .C1(n9454), .C2(n9558), .A(n9775), .B(n7501), .ZN(n9453)
         );
  INV_X1 U9214 ( .A(n9454), .ZN(n7445) );
  INV_X1 U9215 ( .A(n8985), .ZN(n7443) );
  AOI22_X1 U9216 ( .A1(n9823), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n7443), .B2(
        n9822), .ZN(n7444) );
  OAI21_X1 U9217 ( .B1(n7445), .B2(n9825), .A(n7444), .ZN(n7458) );
  INV_X1 U9218 ( .A(n8436), .ZN(n8251) );
  NAND2_X1 U9219 ( .A1(n7427), .A2(n7686), .ZN(n8187) );
  INV_X1 U9220 ( .A(n9556), .ZN(n9548) );
  AOI211_X1 U9221 ( .C1(n7447), .C2(n8375), .A(n9746), .B(n7484), .ZN(n7456)
         );
  OR2_X1 U9222 ( .A1(n7686), .A2(n9017), .ZN(n7455) );
  INV_X1 U9223 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n9126) );
  INV_X1 U9224 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n9124) );
  OR2_X1 U9225 ( .A1(n8177), .A2(n9124), .ZN(n7448) );
  OAI21_X1 U9226 ( .B1(n7941), .B2(n9126), .A(n7448), .ZN(n7453) );
  OR2_X1 U9227 ( .A1(n8992), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n7449) );
  NAND2_X1 U9228 ( .A1(n7490), .A2(n7449), .ZN(n7503) );
  INV_X1 U9229 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n7450) );
  OR2_X1 U9230 ( .A1(n8179), .A2(n7450), .ZN(n7451) );
  OAI21_X1 U9231 ( .B1(n6262), .B2(n7503), .A(n7451), .ZN(n7452) );
  NAND2_X1 U9232 ( .A1(n9064), .A2(n9052), .ZN(n7454) );
  NAND2_X1 U9233 ( .A1(n7455), .A2(n7454), .ZN(n8983) );
  NOR2_X1 U9234 ( .A1(n7456), .A2(n8983), .ZN(n9456) );
  NOR2_X1 U9235 ( .A1(n9456), .A2(n9823), .ZN(n7457) );
  AOI211_X1 U9236 ( .C1(n9453), .C2(n9832), .A(n7458), .B(n7457), .ZN(n7459)
         );
  OAI21_X1 U9237 ( .B1(n9378), .B2(n9458), .A(n7459), .ZN(P1_U3277) );
  AOI21_X1 U9238 ( .B1(n7461), .B2(n7460), .A(n7538), .ZN(n7469) );
  NOR2_X1 U9239 ( .A1(n9537), .A2(n7609), .ZN(n7462) );
  AOI211_X1 U9240 ( .C1(n8580), .C2(n8592), .A(n7463), .B(n7462), .ZN(n7464)
         );
  OAI21_X1 U9241 ( .B1(n7465), .B2(n8577), .A(n7464), .ZN(n7466) );
  AOI21_X1 U9242 ( .B1(n7467), .B2(n9539), .A(n7466), .ZN(n7468) );
  OAI21_X1 U9243 ( .B1(n7469), .B2(n9543), .A(n7468), .ZN(P2_U3174) );
  NAND2_X1 U9244 ( .A1(n7470), .A2(n7477), .ZN(n7471) );
  AND2_X1 U9245 ( .A1(n7472), .A2(n7471), .ZN(n7473) );
  NAND3_X1 U9246 ( .A1(n7472), .A2(n7524), .A3(n7471), .ZN(n7523) );
  OAI211_X1 U9247 ( .C1(n7473), .C2(n7524), .A(n8572), .B(n7523), .ZN(n7481)
         );
  INV_X1 U9248 ( .A(n7474), .ZN(n7479) );
  AOI21_X1 U9249 ( .B1(n8547), .B2(n8592), .A(n7475), .ZN(n7476) );
  OAI21_X1 U9250 ( .B1(n7477), .B2(n8530), .A(n7476), .ZN(n7478) );
  AOI21_X1 U9251 ( .B1(n7479), .B2(n8563), .A(n7478), .ZN(n7480) );
  OAI211_X1 U9252 ( .C1(n10104), .C2(n8583), .A(n7481), .B(n7480), .ZN(
        P2_U3176) );
  INV_X1 U9253 ( .A(n8309), .ZN(n7600) );
  AOI22_X1 U9254 ( .A1(n7482), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_29__SCAN_IN), .B2(n7628), .ZN(n7483) );
  OAI21_X1 U9255 ( .B1(n7600), .B2(n8494), .A(n7483), .ZN(P2_U3266) );
  INV_X1 U9256 ( .A(n8256), .ZN(n8437) );
  NAND2_X1 U9257 ( .A1(n7485), .A2(n7777), .ZN(n7487) );
  AOI22_X1 U9258 ( .A1(n7714), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n7713), .B2(
        n9140), .ZN(n7486) );
  INV_X1 U9259 ( .A(n9064), .ZN(n7632) );
  OR2_X1 U9260 ( .A1(n9449), .A2(n7632), .ZN(n8260) );
  NAND2_X1 U9261 ( .A1(n9449), .A2(n7632), .ZN(n8443) );
  NAND2_X1 U9262 ( .A1(n8260), .A2(n8443), .ZN(n8376) );
  AOI211_X1 U9263 ( .C1(n7488), .C2(n8376), .A(n9746), .B(n7641), .ZN(n7498)
         );
  OR2_X2 U9264 ( .A1(n7490), .A2(n7489), .ZN(n7642) );
  NAND2_X1 U9265 ( .A1(n7490), .A2(n7489), .ZN(n7491) );
  NAND2_X1 U9266 ( .A1(n7642), .A2(n7491), .ZN(n7650) );
  INV_X1 U9267 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n7492) );
  OAI22_X1 U9268 ( .A1(n7650), .A2(n6262), .B1(n8177), .B2(n7492), .ZN(n7496)
         );
  INV_X1 U9269 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n7494) );
  INV_X1 U9270 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n7493) );
  OAI22_X1 U9271 ( .A1(n7941), .A2(n7494), .B1(n8179), .B2(n7493), .ZN(n7495)
         );
  AOI22_X1 U9272 ( .A1(n9171), .A2(n9052), .B1(n9065), .B2(n9225), .ZN(n8994)
         );
  INV_X1 U9273 ( .A(n8994), .ZN(n7497) );
  NOR2_X1 U9274 ( .A1(n7498), .A2(n7497), .ZN(n9451) );
  XOR2_X1 U9275 ( .A(n7635), .B(n8376), .Z(n9452) );
  OR2_X1 U9276 ( .A1(n9452), .A2(n9378), .ZN(n7507) );
  INV_X1 U9277 ( .A(n7501), .ZN(n7502) );
  INV_X1 U9278 ( .A(n9449), .ZN(n7631) );
  AOI211_X1 U9279 ( .C1(n9449), .C2(n7502), .A(n9775), .B(n7648), .ZN(n9448)
         );
  NOR2_X1 U9280 ( .A1(n7631), .A2(n9825), .ZN(n7505) );
  OAI22_X1 U9281 ( .A1(n9335), .A2(n9126), .B1(n7503), .B2(n9799), .ZN(n7504)
         );
  AOI211_X1 U9282 ( .C1(n9448), .C2(n9832), .A(n7505), .B(n7504), .ZN(n7506)
         );
  OAI211_X1 U9283 ( .C1(n9836), .C2(n9451), .A(n7507), .B(n7506), .ZN(P1_U3276) );
  XOR2_X1 U9284 ( .A(n7508), .B(n8149), .Z(n7522) );
  INV_X1 U9285 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n7512) );
  OAI21_X1 U9286 ( .B1(n7510), .B2(n5316), .A(n7509), .ZN(n7511) );
  AOI222_X1 U9287 ( .A1(n5513), .A2(n7511), .B1(n8590), .B2(n8807), .C1(n8588), 
        .C2(n8809), .ZN(n7518) );
  MUX2_X1 U9288 ( .A(n7512), .B(n7518), .S(n10118), .Z(n7514) );
  NAND2_X1 U9289 ( .A1(n8927), .A2(n7603), .ZN(n7513) );
  OAI211_X1 U9290 ( .C1(n7522), .C2(n8931), .A(n7514), .B(n7513), .ZN(P2_U3435) );
  MUX2_X1 U9291 ( .A(n7515), .B(n7518), .S(n10135), .Z(n7517) );
  NAND2_X1 U9292 ( .A1(n7603), .A2(n8856), .ZN(n7516) );
  OAI211_X1 U9293 ( .C1(n8859), .C2(n7522), .A(n7517), .B(n7516), .ZN(P2_U3474) );
  MUX2_X1 U9294 ( .A(n8604), .B(n7518), .S(n10050), .Z(n7521) );
  INV_X1 U9295 ( .A(n7519), .ZN(n7611) );
  AOI22_X1 U9296 ( .A1(n7603), .A2(n8816), .B1(n8815), .B2(n7611), .ZN(n7520)
         );
  OAI211_X1 U9297 ( .C1(n7522), .C2(n8819), .A(n7521), .B(n7520), .ZN(P2_U3218) );
  OAI21_X1 U9298 ( .B1(n7525), .B2(n7524), .A(n7523), .ZN(n7527) );
  XNOR2_X1 U9299 ( .A(n7527), .B(n7526), .ZN(n7535) );
  NOR2_X1 U9300 ( .A1(n9537), .A2(n7528), .ZN(n7529) );
  AOI211_X1 U9301 ( .C1(n8580), .C2(n8593), .A(n7530), .B(n7529), .ZN(n7531)
         );
  OAI21_X1 U9302 ( .B1(n7532), .B2(n8577), .A(n7531), .ZN(n7533) );
  AOI21_X1 U9303 ( .B1(n10113), .B2(n9539), .A(n7533), .ZN(n7534) );
  OAI21_X1 U9304 ( .B1(n7535), .B2(n9543), .A(n7534), .ZN(P2_U3164) );
  NOR3_X1 U9305 ( .A1(n7538), .A2(n7537), .A3(n7536), .ZN(n7539) );
  OAI21_X1 U9306 ( .B1(n4415), .B2(n7539), .A(n8572), .ZN(n7546) );
  INV_X1 U9307 ( .A(n7540), .ZN(n7544) );
  AOI21_X1 U9308 ( .B1(n8580), .B2(n8591), .A(n7541), .ZN(n7542) );
  OAI21_X1 U9309 ( .B1(n7584), .B2(n9537), .A(n7542), .ZN(n7543) );
  AOI21_X1 U9310 ( .B1(n7544), .B2(n8563), .A(n7543), .ZN(n7545) );
  OAI211_X1 U9311 ( .C1(n7547), .C2(n8583), .A(n7546), .B(n7545), .ZN(P2_U3155) );
  NAND2_X1 U9312 ( .A1(n9918), .A2(n6252), .ZN(n7554) );
  NAND2_X1 U9313 ( .A1(n9067), .A2(n7709), .ZN(n7553) );
  NAND2_X1 U9314 ( .A1(n7554), .A2(n7553), .ZN(n7555) );
  XNOR2_X1 U9315 ( .A(n7683), .B(n4410), .ZN(n7559) );
  OAI22_X1 U9316 ( .A1(n7557), .A2(n7948), .B1(n7556), .B2(n6158), .ZN(n7558)
         );
  AOI21_X1 U9317 ( .B1(n7559), .B2(n7558), .A(n7685), .ZN(n7565) );
  AOI22_X1 U9318 ( .A1(n9018), .A2(n7560), .B1(P1_REG3_REG_14__SCAN_IN), .B2(
        P1_U3086), .ZN(n7561) );
  OAI21_X1 U9319 ( .B1(n9021), .B2(n7562), .A(n7561), .ZN(n7563) );
  AOI21_X1 U9320 ( .B1(n9918), .B2(n9023), .A(n7563), .ZN(n7564) );
  OAI21_X1 U9321 ( .B1(n7565), .B2(n9036), .A(n7564), .ZN(P1_U3215) );
  NAND2_X1 U9322 ( .A1(n7566), .A2(SI_29_), .ZN(n7571) );
  INV_X1 U9323 ( .A(n7567), .ZN(n7568) );
  INV_X1 U9324 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n8319) );
  INV_X1 U9325 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n7572) );
  MUX2_X1 U9326 ( .A(n8319), .B(n7572), .S(n5052), .Z(n7573) );
  NAND2_X1 U9327 ( .A1(n7573), .A2(n6975), .ZN(n7615) );
  INV_X1 U9328 ( .A(n7573), .ZN(n7574) );
  NAND2_X1 U9329 ( .A1(n7574), .A2(SI_30_), .ZN(n7575) );
  NAND2_X1 U9330 ( .A1(n7615), .A2(n7575), .ZN(n7616) );
  INV_X1 U9331 ( .A(n8318), .ZN(n7602) );
  AOI22_X1 U9332 ( .A1(n7576), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n7628), .ZN(n7577) );
  OAI21_X1 U9333 ( .B1(n7602), .B2(n8494), .A(n7577), .ZN(P2_U3265) );
  INV_X1 U9334 ( .A(n7580), .ZN(n8150) );
  XNOR2_X1 U9335 ( .A(n7578), .B(n8150), .ZN(n7598) );
  INV_X1 U9336 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n7587) );
  INV_X1 U9337 ( .A(n7579), .ZN(n7583) );
  AOI21_X1 U9338 ( .B1(n7509), .B2(n7581), .A(n7580), .ZN(n7582) );
  NOR3_X1 U9339 ( .A1(n7583), .A2(n7582), .A3(n8792), .ZN(n7586) );
  OAI22_X1 U9340 ( .A1(n7584), .A2(n10043), .B1(n7674), .B2(n10041), .ZN(n7585) );
  NOR2_X1 U9341 ( .A1(n7586), .A2(n7585), .ZN(n7593) );
  MUX2_X1 U9342 ( .A(n7587), .B(n7593), .S(n10118), .Z(n7589) );
  NAND2_X1 U9343 ( .A1(n8927), .A2(n7679), .ZN(n7588) );
  OAI211_X1 U9344 ( .C1(n7598), .C2(n8931), .A(n7589), .B(n7588), .ZN(P2_U3438) );
  MUX2_X1 U9345 ( .A(n7590), .B(n7593), .S(n10135), .Z(n7592) );
  NAND2_X1 U9346 ( .A1(n7679), .A2(n8856), .ZN(n7591) );
  OAI211_X1 U9347 ( .C1(n7598), .C2(n8859), .A(n7592), .B(n7591), .ZN(P2_U3475) );
  MUX2_X1 U9348 ( .A(n7594), .B(n7593), .S(n10050), .Z(n7597) );
  INV_X1 U9349 ( .A(n7677), .ZN(n7595) );
  AOI22_X1 U9350 ( .A1(n7679), .A2(n8816), .B1(n8815), .B2(n7595), .ZN(n7596)
         );
  OAI211_X1 U9351 ( .C1(n7598), .C2(n8819), .A(n7597), .B(n7596), .ZN(P2_U3217) );
  INV_X1 U9352 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n8310) );
  OAI222_X1 U9353 ( .A1(n7915), .A2(n7600), .B1(P1_U3086), .B2(n7599), .C1(
        n8310), .C2(n7913), .ZN(P1_U3326) );
  OAI222_X1 U9354 ( .A1(n7913), .A2(n8319), .B1(n7915), .B2(n7602), .C1(
        P1_U3086), .C2(n7601), .ZN(P1_U3325) );
  INV_X1 U9355 ( .A(n7603), .ZN(n7614) );
  AOI21_X1 U9356 ( .B1(n7605), .B2(n7604), .A(n9543), .ZN(n7607) );
  NAND2_X1 U9357 ( .A1(n7607), .A2(n7606), .ZN(n7613) );
  AND2_X1 U9358 ( .A1(P2_U3151), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8612) );
  AOI21_X1 U9359 ( .B1(n8547), .B2(n8588), .A(n8612), .ZN(n7608) );
  OAI21_X1 U9360 ( .B1(n7609), .B2(n8530), .A(n7608), .ZN(n7610) );
  AOI21_X1 U9361 ( .B1(n7611), .B2(n8563), .A(n7610), .ZN(n7612) );
  OAI211_X1 U9362 ( .C1(n7614), .C2(n8583), .A(n7613), .B(n7612), .ZN(P2_U3181) );
  MUX2_X1 U9363 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n5052), .Z(n7619) );
  XNOR2_X1 U9364 ( .A(n7619), .B(n7618), .ZN(n7620) );
  INV_X1 U9365 ( .A(n8172), .ZN(n7630) );
  NOR3_X1 U9366 ( .A1(n7622), .A2(n5973), .A3(P1_U3086), .ZN(n7623) );
  AOI21_X1 U9367 ( .B1(n7624), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n7623), .ZN(
        n7625) );
  OAI21_X1 U9368 ( .B1(n7630), .B2(n7915), .A(n7625), .ZN(P1_U3324) );
  NOR4_X1 U9369 ( .A1(n7626), .A2(P2_IR_REG_30__SCAN_IN), .A3(P2_U3151), .A4(
        n4915), .ZN(n7627) );
  AOI21_X1 U9370 ( .B1(n7628), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n7627), .ZN(
        n7629) );
  OAI21_X1 U9371 ( .B1(n7630), .B2(n8494), .A(n7629), .ZN(P2_U3264) );
  NAND2_X1 U9372 ( .A1(n9449), .A2(n9064), .ZN(n7634) );
  AOI22_X1 U9373 ( .A1(n7714), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n7713), .B2(
        n9144), .ZN(n7638) );
  NAND2_X1 U9374 ( .A1(n9173), .A2(n9171), .ZN(n8262) );
  INV_X1 U9375 ( .A(n9171), .ZN(n9172) );
  NAND2_X1 U9376 ( .A1(n9445), .A2(n9172), .ZN(n8324) );
  NAND2_X1 U9377 ( .A1(n8262), .A2(n8324), .ZN(n8377) );
  XNOR2_X1 U9378 ( .A(n9174), .B(n8377), .ZN(n9447) );
  INV_X1 U9379 ( .A(n8260), .ZN(n7640) );
  XNOR2_X1 U9380 ( .A(n8327), .B(n8377), .ZN(n7647) );
  NAND2_X1 U9381 ( .A1(n7642), .A2(n8955), .ZN(n7643) );
  NAND2_X1 U9382 ( .A1(n7728), .A2(n7643), .ZN(n9367) );
  INV_X1 U9383 ( .A(n8179), .ZN(n7644) );
  AOI22_X1 U9384 ( .A1(n7731), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n7644), .B2(
        P1_REG0_REG_19__SCAN_IN), .ZN(n7646) );
  INV_X1 U9385 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n9139) );
  OR2_X1 U9386 ( .A1(n8177), .A2(n9139), .ZN(n7645) );
  OAI211_X1 U9387 ( .C1(n9367), .C2(n6262), .A(n7646), .B(n7645), .ZN(n9175)
         );
  AOI22_X1 U9388 ( .A1(n9175), .A2(n9052), .B1(n9225), .B2(n9064), .ZN(n9042)
         );
  OAI21_X1 U9389 ( .B1(n7647), .B2(n9746), .A(n9042), .ZN(n9443) );
  INV_X1 U9390 ( .A(n7648), .ZN(n7649) );
  AOI211_X1 U9391 ( .C1(n9445), .C2(n7649), .A(n9775), .B(n9363), .ZN(n9444)
         );
  NAND2_X1 U9392 ( .A1(n9444), .A2(n9832), .ZN(n7652) );
  INV_X1 U9393 ( .A(n7650), .ZN(n9044) );
  AOI22_X1 U9394 ( .A1(n9823), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9044), .B2(
        n9822), .ZN(n7651) );
  OAI211_X1 U9395 ( .C1(n9173), .C2(n9825), .A(n7652), .B(n7651), .ZN(n7653)
         );
  AOI21_X1 U9396 ( .B1(n9443), .B2(n9335), .A(n7653), .ZN(n7654) );
  OAI21_X1 U9397 ( .B1(n9447), .B2(n9378), .A(n7654), .ZN(P1_U3275) );
  XNOR2_X1 U9398 ( .A(n7655), .B(n8046), .ZN(n7670) );
  INV_X1 U9399 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n7659) );
  XNOR2_X1 U9400 ( .A(n7657), .B(n8046), .ZN(n7658) );
  AOI222_X1 U9401 ( .A1(n5513), .A2(n7658), .B1(n8587), .B2(n8809), .C1(n8588), 
        .C2(n8807), .ZN(n7666) );
  MUX2_X1 U9402 ( .A(n7659), .B(n7666), .S(n10118), .Z(n7661) );
  NAND2_X1 U9403 ( .A1(n8544), .A2(n8927), .ZN(n7660) );
  OAI211_X1 U9404 ( .C1(n7670), .C2(n8931), .A(n7661), .B(n7660), .ZN(P2_U3441) );
  MUX2_X1 U9405 ( .A(n7662), .B(n7666), .S(n10050), .Z(n7665) );
  INV_X1 U9406 ( .A(n8542), .ZN(n7663) );
  AOI22_X1 U9407 ( .A1(n8544), .A2(n8816), .B1(n8815), .B2(n7663), .ZN(n7664)
         );
  OAI211_X1 U9408 ( .C1(n7670), .C2(n8819), .A(n7665), .B(n7664), .ZN(P2_U3216) );
  MUX2_X1 U9409 ( .A(n7667), .B(n7666), .S(n10135), .Z(n7669) );
  NAND2_X1 U9410 ( .A1(n8544), .A2(n8856), .ZN(n7668) );
  OAI211_X1 U9411 ( .C1(n7670), .C2(n8859), .A(n7669), .B(n7668), .ZN(P2_U3476) );
  XNOR2_X1 U9412 ( .A(n7672), .B(n7671), .ZN(n7681) );
  NOR2_X1 U9413 ( .A1(n7673), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8631) );
  NOR2_X1 U9414 ( .A1(n9537), .A2(n7674), .ZN(n7675) );
  AOI211_X1 U9415 ( .C1(n8580), .C2(n8589), .A(n8631), .B(n7675), .ZN(n7676)
         );
  OAI21_X1 U9416 ( .B1(n7677), .B2(n8577), .A(n7676), .ZN(n7678) );
  AOI21_X1 U9417 ( .B1(n7679), .B2(n9539), .A(n7678), .ZN(n7680) );
  OAI21_X1 U9418 ( .B1(n7681), .B2(n9543), .A(n7680), .ZN(P2_U3166) );
  INV_X1 U9419 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7763) );
  OAI222_X1 U9420 ( .A1(n7915), .A2(n7682), .B1(n6075), .B2(P1_U3086), .C1(
        n7763), .C2(n7913), .ZN(P1_U3333) );
  NAND2_X1 U9421 ( .A1(n7427), .A2(n6252), .ZN(n7688) );
  OR2_X1 U9422 ( .A1(n7686), .A2(n7948), .ZN(n7687) );
  NAND2_X1 U9423 ( .A1(n7688), .A2(n7687), .ZN(n7689) );
  XNOR2_X1 U9424 ( .A(n7689), .B(n7922), .ZN(n7690) );
  XNOR2_X1 U9425 ( .A(n7692), .B(n7690), .ZN(n9048) );
  AOI22_X1 U9426 ( .A1(n7427), .A2(n7709), .B1(n7924), .B2(n9066), .ZN(n9049)
         );
  INV_X1 U9427 ( .A(n7690), .ZN(n7691) );
  NAND2_X1 U9428 ( .A1(n9454), .A2(n4346), .ZN(n7694) );
  NAND2_X1 U9429 ( .A1(n9065), .A2(n7709), .ZN(n7693) );
  NAND2_X1 U9430 ( .A1(n7694), .A2(n7693), .ZN(n7695) );
  XNOR2_X1 U9431 ( .A(n7695), .B(n7949), .ZN(n7696) );
  AOI22_X1 U9432 ( .A1(n9454), .A2(n7709), .B1(n7924), .B2(n9065), .ZN(n7697)
         );
  XNOR2_X1 U9433 ( .A(n7696), .B(n7697), .ZN(n8982) );
  INV_X1 U9434 ( .A(n7696), .ZN(n7698) );
  NAND2_X1 U9435 ( .A1(n9449), .A2(n4346), .ZN(n7700) );
  NAND2_X1 U9436 ( .A1(n9064), .A2(n7709), .ZN(n7699) );
  NAND2_X1 U9437 ( .A1(n7700), .A2(n7699), .ZN(n7701) );
  XNOR2_X1 U9438 ( .A(n7701), .B(n7949), .ZN(n8990) );
  NAND2_X1 U9439 ( .A1(n9449), .A2(n7709), .ZN(n7703) );
  NAND2_X1 U9440 ( .A1(n9064), .A2(n7924), .ZN(n7702) );
  NAND2_X1 U9441 ( .A1(n7703), .A2(n7702), .ZN(n7705) );
  INV_X1 U9442 ( .A(n8990), .ZN(n7706) );
  INV_X1 U9443 ( .A(n7705), .ZN(n8989) );
  NAND2_X1 U9444 ( .A1(n7707), .A2(n4864), .ZN(n8946) );
  OAI22_X1 U9445 ( .A1(n9173), .A2(n7717), .B1(n9172), .B2(n7948), .ZN(n7708)
         );
  XNOR2_X1 U9446 ( .A(n7708), .B(n7922), .ZN(n8947) );
  NAND2_X1 U9447 ( .A1(n9445), .A2(n7709), .ZN(n7711) );
  NAND2_X1 U9448 ( .A1(n9171), .A2(n7924), .ZN(n7710) );
  NAND2_X1 U9449 ( .A1(n7712), .A2(n7777), .ZN(n7716) );
  AOI22_X1 U9450 ( .A1(n7714), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n4349), .B2(
        n7713), .ZN(n7715) );
  INV_X1 U9451 ( .A(n9175), .ZN(n9176) );
  OAI22_X1 U9452 ( .A1(n9370), .A2(n7717), .B1(n9176), .B2(n7948), .ZN(n7718)
         );
  XNOR2_X1 U9453 ( .A(n7718), .B(n7949), .ZN(n8949) );
  OR2_X1 U9454 ( .A1(n9370), .A2(n7948), .ZN(n7720) );
  NAND2_X1 U9455 ( .A1(n9175), .A2(n7924), .ZN(n7719) );
  NAND2_X1 U9456 ( .A1(n7720), .A2(n7719), .ZN(n7722) );
  NAND2_X1 U9457 ( .A1(n8949), .A2(n7722), .ZN(n9010) );
  OAI21_X1 U9458 ( .B1(n8947), .B2(n9040), .A(n9010), .ZN(n7740) );
  INV_X1 U9459 ( .A(n7722), .ZN(n8948) );
  NAND2_X1 U9460 ( .A1(n8947), .A2(n9040), .ZN(n7721) );
  INV_X1 U9461 ( .A(n7721), .ZN(n7738) );
  AOI21_X1 U9462 ( .B1(n7722), .B2(n7721), .A(n8949), .ZN(n7737) );
  NAND2_X1 U9463 ( .A1(n7723), .A2(n7777), .ZN(n7726) );
  OR2_X1 U9464 ( .A1(n4347), .A2(n7724), .ZN(n7725) );
  NAND2_X2 U9465 ( .A1(n7726), .A2(n7725), .ZN(n9435) );
  INV_X1 U9466 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n7727) );
  AND2_X1 U9467 ( .A1(n7728), .A2(n7727), .ZN(n7729) );
  NOR2_X1 U9468 ( .A1(n7747), .A2(n7729), .ZN(n9352) );
  NAND2_X1 U9469 ( .A1(n9352), .A2(n7876), .ZN(n7735) );
  INV_X1 U9470 ( .A(n8177), .ZN(n7730) );
  AOI22_X1 U9471 ( .A1(n7731), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n7730), .B2(
        P1_REG1_REG_20__SCAN_IN), .ZN(n7734) );
  INV_X1 U9472 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n7732) );
  OR2_X1 U9473 ( .A1(n8179), .A2(n7732), .ZN(n7733) );
  INV_X1 U9474 ( .A(n9177), .ZN(n9178) );
  AOI22_X1 U9475 ( .A1(n9435), .A2(n6252), .B1(n7709), .B2(n9178), .ZN(n7736)
         );
  XOR2_X1 U9476 ( .A(n7949), .B(n7736), .Z(n7742) );
  INV_X1 U9477 ( .A(n9435), .ZN(n9354) );
  OAI22_X1 U9478 ( .A1(n9354), .A2(n7948), .B1(n9177), .B2(n6158), .ZN(n7741)
         );
  NOR2_X1 U9479 ( .A1(n7742), .A2(n7741), .ZN(n9014) );
  AOI211_X1 U9480 ( .C1(n8948), .C2(n7738), .A(n7737), .B(n9014), .ZN(n7739)
         );
  NAND2_X1 U9481 ( .A1(n7742), .A2(n7741), .ZN(n9012) );
  NAND2_X1 U9482 ( .A1(n7743), .A2(n7777), .ZN(n7746) );
  OR2_X1 U9483 ( .A1(n4347), .A2(n7744), .ZN(n7745) );
  NAND2_X2 U9484 ( .A1(n7746), .A2(n7745), .ZN(n8183) );
  OR2_X1 U9485 ( .A1(n7747), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n7748) );
  NAND2_X1 U9486 ( .A1(n7747), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n7766) );
  AND2_X1 U9487 ( .A1(n7748), .A2(n7766), .ZN(n9344) );
  NAND2_X1 U9488 ( .A1(n9344), .A2(n7876), .ZN(n7755) );
  INV_X1 U9489 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n9336) );
  INV_X1 U9490 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n7749) );
  OR2_X1 U9491 ( .A1(n8177), .A2(n7749), .ZN(n7752) );
  INV_X1 U9492 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n7750) );
  OR2_X1 U9493 ( .A1(n8179), .A2(n7750), .ZN(n7751) );
  OAI211_X1 U9494 ( .C1(n7941), .C2(n9336), .A(n7752), .B(n7751), .ZN(n7753)
         );
  INV_X1 U9495 ( .A(n7753), .ZN(n7754) );
  AOI22_X1 U9496 ( .A1(n8183), .A2(n4346), .B1(n7709), .B2(n9170), .ZN(n7756)
         );
  XNOR2_X1 U9497 ( .A(n7756), .B(n7949), .ZN(n7758) );
  OAI22_X1 U9498 ( .A1(n9337), .A2(n7948), .B1(n9181), .B2(n6158), .ZN(n7759)
         );
  XNOR2_X1 U9499 ( .A(n7758), .B(n7759), .ZN(n8962) );
  AND2_X1 U9500 ( .A1(n9012), .A2(n8962), .ZN(n7757) );
  NAND2_X1 U9501 ( .A1(n7762), .A2(n7777), .ZN(n7765) );
  OR2_X1 U9502 ( .A1(n4347), .A2(n7763), .ZN(n7764) );
  NAND2_X2 U9503 ( .A1(n7765), .A2(n7764), .ZN(n9426) );
  INV_X1 U9504 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n9032) );
  NAND2_X1 U9505 ( .A1(n7766), .A2(n9032), .ZN(n7767) );
  AND2_X1 U9506 ( .A1(n7782), .A2(n7767), .ZN(n9321) );
  INV_X1 U9507 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n7772) );
  INV_X1 U9508 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n7768) );
  OR2_X1 U9509 ( .A1(n8177), .A2(n7768), .ZN(n7771) );
  INV_X1 U9510 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n7769) );
  OR2_X1 U9511 ( .A1(n8179), .A2(n7769), .ZN(n7770) );
  OAI211_X1 U9512 ( .C1(n7941), .C2(n7772), .A(n7771), .B(n7770), .ZN(n7773)
         );
  AOI21_X1 U9513 ( .B1(n9321), .B2(n7876), .A(n7773), .ZN(n9185) );
  INV_X1 U9514 ( .A(n9185), .ZN(n9184) );
  AOI22_X1 U9515 ( .A1(n9426), .A2(n4346), .B1(n7709), .B2(n9184), .ZN(n7774)
         );
  XNOR2_X1 U9516 ( .A(n7774), .B(n7949), .ZN(n7775) );
  OAI22_X1 U9517 ( .A1(n9323), .A2(n7948), .B1(n9185), .B2(n6158), .ZN(n9029)
         );
  NAND2_X1 U9518 ( .A1(n9027), .A2(n9029), .ZN(n7776) );
  NAND2_X1 U9519 ( .A1(n7776), .A2(n9026), .ZN(n7842) );
  NAND2_X1 U9520 ( .A1(n7778), .A2(n7777), .ZN(n7781) );
  OR2_X1 U9521 ( .A1(n4347), .A2(n7779), .ZN(n7780) );
  NAND2_X1 U9522 ( .A1(n9421), .A2(n4346), .ZN(n7793) );
  INV_X1 U9523 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n7810) );
  AND2_X1 U9524 ( .A1(n7782), .A2(n7810), .ZN(n7783) );
  NOR2_X1 U9525 ( .A1(n7800), .A2(n7783), .ZN(n9306) );
  NAND2_X1 U9526 ( .A1(n9306), .A2(n7876), .ZN(n7791) );
  INV_X1 U9527 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n7788) );
  INV_X1 U9528 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n7784) );
  OR2_X1 U9529 ( .A1(n8177), .A2(n7784), .ZN(n7787) );
  INV_X1 U9530 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n7785) );
  OR2_X1 U9531 ( .A1(n8179), .A2(n7785), .ZN(n7786) );
  OAI211_X1 U9532 ( .C1(n7941), .C2(n7788), .A(n7787), .B(n7786), .ZN(n7789)
         );
  INV_X1 U9533 ( .A(n7789), .ZN(n7790) );
  OR2_X1 U9534 ( .A1(n9188), .A2(n7948), .ZN(n7792) );
  NAND2_X1 U9535 ( .A1(n7793), .A2(n7792), .ZN(n7794) );
  XNOR2_X1 U9536 ( .A(n7794), .B(n7922), .ZN(n7797) );
  NOR2_X1 U9537 ( .A1(n9188), .A2(n6158), .ZN(n7795) );
  AOI21_X1 U9538 ( .B1(n9421), .B2(n7709), .A(n7795), .ZN(n7796) );
  NOR2_X1 U9539 ( .A1(n7797), .A2(n7796), .ZN(n7843) );
  NAND2_X1 U9540 ( .A1(n7797), .A2(n7796), .ZN(n7893) );
  INV_X1 U9541 ( .A(n7893), .ZN(n7798) );
  NOR2_X1 U9542 ( .A1(n7843), .A2(n7798), .ZN(n7799) );
  XNOR2_X1 U9543 ( .A(n7842), .B(n7799), .ZN(n7814) );
  NAND2_X1 U9544 ( .A1(n7800), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n7857) );
  OR2_X1 U9545 ( .A1(n7800), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n7801) );
  AND2_X1 U9546 ( .A1(n7857), .A2(n7801), .ZN(n9294) );
  INV_X1 U9547 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n7806) );
  INV_X1 U9548 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n7802) );
  OR2_X1 U9549 ( .A1(n8177), .A2(n7802), .ZN(n7805) );
  INV_X1 U9550 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n7803) );
  OR2_X1 U9551 ( .A1(n8179), .A2(n7803), .ZN(n7804) );
  OAI211_X1 U9552 ( .C1(n7941), .C2(n7806), .A(n7805), .B(n7804), .ZN(n7807)
         );
  OR2_X1 U9553 ( .A1(n9189), .A2(n9162), .ZN(n7809) );
  OR2_X1 U9554 ( .A1(n9185), .A2(n9017), .ZN(n7808) );
  AND2_X1 U9555 ( .A1(n7809), .A2(n7808), .ZN(n9312) );
  OAI22_X1 U9556 ( .A1(n9312), .A2(n9056), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n7810), .ZN(n7812) );
  INV_X1 U9557 ( .A(n9421), .ZN(n9308) );
  NOR2_X1 U9558 ( .A1(n9308), .A2(n9061), .ZN(n7811) );
  AOI211_X1 U9559 ( .C1(n9306), .C2(n9058), .A(n7812), .B(n7811), .ZN(n7813)
         );
  OAI21_X1 U9560 ( .B1(n7814), .B2(n9036), .A(n7813), .ZN(P1_U3216) );
  INV_X1 U9561 ( .A(n7817), .ZN(n7818) );
  NAND2_X1 U9562 ( .A1(n7819), .A2(n7818), .ZN(n7821) );
  OAI21_X1 U9563 ( .B1(n7819), .B2(n7818), .A(n7821), .ZN(n7829) );
  NOR2_X1 U9564 ( .A1(n7829), .A2(n8753), .ZN(n7830) );
  INV_X1 U9565 ( .A(n7820), .ZN(n7823) );
  INV_X1 U9566 ( .A(n7821), .ZN(n7822) );
  NOR3_X1 U9567 ( .A1(n7830), .A2(n7823), .A3(n7822), .ZN(n7824) );
  INV_X1 U9568 ( .A(n8472), .ZN(n8524) );
  OAI21_X1 U9569 ( .B1(n7824), .B2(n8524), .A(n8572), .ZN(n7828) );
  AOI22_X1 U9570 ( .A1(n8547), .A2(n8702), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3151), .ZN(n7825) );
  OAI21_X1 U9571 ( .B1(n8731), .B2(n8530), .A(n7825), .ZN(n7826) );
  AOI21_X1 U9572 ( .B1(n8733), .B2(n8563), .A(n7826), .ZN(n7827) );
  OAI211_X1 U9573 ( .C1(n8893), .C2(n8583), .A(n7828), .B(n7827), .ZN(P2_U3169) );
  AOI21_X1 U9574 ( .B1(n8753), .B2(n7829), .A(n7830), .ZN(n7836) );
  NAND2_X1 U9575 ( .A1(n8563), .A2(n8744), .ZN(n7832) );
  AOI22_X1 U9576 ( .A1(n8547), .A2(n8741), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3151), .ZN(n7831) );
  OAI211_X1 U9577 ( .C1(n7833), .C2(n8530), .A(n7832), .B(n7831), .ZN(n7834)
         );
  AOI21_X1 U9578 ( .B1(n8899), .B2(n9539), .A(n7834), .ZN(n7835) );
  OAI21_X1 U9579 ( .B1(n7836), .B2(n9543), .A(n7835), .ZN(P2_U3156) );
  INV_X1 U9580 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n7917) );
  OAI222_X1 U9581 ( .A1(n7915), .A2(n7837), .B1(n6484), .B2(P1_U3086), .C1(
        n7917), .C2(n7913), .ZN(P1_U3328) );
  NAND2_X1 U9582 ( .A1(n7838), .A2(n7777), .ZN(n7841) );
  OR2_X1 U9583 ( .A1(n4347), .A2(n7839), .ZN(n7840) );
  INV_X1 U9584 ( .A(n7842), .ZN(n7845) );
  NAND2_X1 U9585 ( .A1(n7895), .A2(n7893), .ZN(n9002) );
  NAND2_X1 U9586 ( .A1(n7846), .A2(n7777), .ZN(n7849) );
  OR2_X1 U9587 ( .A1(n4347), .A2(n7847), .ZN(n7848) );
  INV_X1 U9588 ( .A(n9189), .ZN(n9190) );
  AOI22_X1 U9589 ( .A1(n9416), .A2(n6252), .B1(n7709), .B2(n9190), .ZN(n7850)
         );
  XOR2_X1 U9590 ( .A(n7949), .B(n7850), .Z(n7852) );
  OAI22_X1 U9591 ( .A1(n9154), .A2(n7948), .B1(n9189), .B2(n6158), .ZN(n7851)
         );
  NOR2_X1 U9592 ( .A1(n7852), .A2(n7851), .ZN(n7870) );
  AOI21_X1 U9593 ( .B1(n7852), .B2(n7851), .A(n7870), .ZN(n9003) );
  NAND2_X1 U9594 ( .A1(n7853), .A2(n7777), .ZN(n7856) );
  OR2_X1 U9595 ( .A1(n4347), .A2(n7854), .ZN(n7855) );
  INV_X1 U9596 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n8976) );
  NAND2_X1 U9597 ( .A1(n7857), .A2(n8976), .ZN(n7858) );
  NAND2_X1 U9598 ( .A1(n9280), .A2(n7876), .ZN(n7866) );
  INV_X1 U9599 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n7863) );
  INV_X1 U9600 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n7859) );
  OR2_X1 U9601 ( .A1(n8177), .A2(n7859), .ZN(n7862) );
  INV_X1 U9602 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n7860) );
  OR2_X1 U9603 ( .A1(n8179), .A2(n7860), .ZN(n7861) );
  OAI211_X1 U9604 ( .C1(n7941), .C2(n7863), .A(n7862), .B(n7861), .ZN(n7864)
         );
  INV_X1 U9605 ( .A(n7864), .ZN(n7865) );
  OAI22_X1 U9606 ( .A1(n9282), .A2(n7948), .B1(n9193), .B2(n6158), .ZN(n7873)
         );
  NAND2_X1 U9607 ( .A1(n9411), .A2(n6252), .ZN(n7868) );
  INV_X1 U9608 ( .A(n9193), .ZN(n9192) );
  NAND2_X1 U9609 ( .A1(n9192), .A2(n7709), .ZN(n7867) );
  NAND2_X1 U9610 ( .A1(n7868), .A2(n7867), .ZN(n7869) );
  XNOR2_X1 U9611 ( .A(n7869), .B(n7949), .ZN(n7874) );
  XOR2_X1 U9612 ( .A(n7873), .B(n7874), .Z(n8974) );
  AND2_X1 U9613 ( .A1(n9003), .A2(n8974), .ZN(n7897) );
  NAND2_X1 U9614 ( .A1(n9002), .A2(n7897), .ZN(n7872) );
  INV_X1 U9615 ( .A(n8974), .ZN(n7871) );
  INV_X1 U9616 ( .A(n7870), .ZN(n8970) );
  NOR2_X1 U9617 ( .A1(n7874), .A2(n7873), .ZN(n7889) );
  NAND2_X1 U9618 ( .A1(n9406), .A2(n4346), .ZN(n7886) );
  INV_X1 U9619 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n7908) );
  NOR2_X2 U9620 ( .A1(n7875), .A2(n7908), .ZN(n7903) );
  AOI21_X1 U9621 ( .B1(n7875), .B2(n7908), .A(n7903), .ZN(n9269) );
  NAND2_X1 U9622 ( .A1(n9269), .A2(n7876), .ZN(n7884) );
  INV_X1 U9623 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n7881) );
  INV_X1 U9624 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n7877) );
  OR2_X1 U9625 ( .A1(n8177), .A2(n7877), .ZN(n7880) );
  INV_X1 U9626 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n7878) );
  OR2_X1 U9627 ( .A1(n8179), .A2(n7878), .ZN(n7879) );
  OAI211_X1 U9628 ( .C1(n7941), .C2(n7881), .A(n7880), .B(n7879), .ZN(n7882)
         );
  INV_X1 U9629 ( .A(n7882), .ZN(n7883) );
  OR2_X1 U9630 ( .A1(n9195), .A2(n7948), .ZN(n7885) );
  NAND2_X1 U9631 ( .A1(n7886), .A2(n7885), .ZN(n7887) );
  XNOR2_X1 U9632 ( .A(n7887), .B(n7922), .ZN(n7927) );
  NOR2_X1 U9633 ( .A1(n9195), .A2(n6158), .ZN(n7888) );
  AOI21_X1 U9634 ( .B1(n9406), .B2(n7709), .A(n7888), .ZN(n7928) );
  XNOR2_X1 U9635 ( .A(n7927), .B(n7928), .ZN(n7890) );
  OAI21_X1 U9636 ( .B1(n8971), .B2(n7889), .A(n7890), .ZN(n7899) );
  NOR2_X1 U9637 ( .A1(n7890), .A2(n7889), .ZN(n7892) );
  AND2_X1 U9638 ( .A1(n7892), .A2(n7891), .ZN(n7896) );
  AND2_X1 U9639 ( .A1(n7893), .A2(n7896), .ZN(n7894) );
  INV_X1 U9640 ( .A(n7896), .ZN(n7898) );
  NAND3_X1 U9641 ( .A1(n7899), .A2(n4404), .A3(n9050), .ZN(n7912) );
  INV_X1 U9642 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n7902) );
  INV_X1 U9643 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n7900) );
  OR2_X1 U9644 ( .A1(n8177), .A2(n7900), .ZN(n7901) );
  OAI21_X1 U9645 ( .B1(n7941), .B2(n7902), .A(n7901), .ZN(n7907) );
  OAI21_X1 U9646 ( .B1(P1_REG3_REG_27__SCAN_IN), .B2(n7903), .A(n7943), .ZN(
        n9254) );
  INV_X1 U9647 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n7904) );
  OR2_X1 U9648 ( .A1(n8179), .A2(n7904), .ZN(n7905) );
  OAI21_X1 U9649 ( .B1(n6262), .B2(n9254), .A(n7905), .ZN(n7906) );
  INV_X2 U9650 ( .A(n9063), .ZN(n9198) );
  OAI22_X1 U9651 ( .A1(n9193), .A2(n9017), .B1(n9198), .B2(n9162), .ZN(n9273)
         );
  INV_X1 U9652 ( .A(n9269), .ZN(n7909) );
  OAI22_X1 U9653 ( .A1(n7909), .A2(n9021), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n7908), .ZN(n7910) );
  AOI21_X1 U9654 ( .B1(n9273), .B2(n9018), .A(n7910), .ZN(n7911) );
  OAI211_X1 U9655 ( .C1(n4637), .C2(n9061), .A(n7912), .B(n7911), .ZN(P1_U3240) );
  INV_X1 U9656 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n7935) );
  OAI222_X1 U9657 ( .A1(n7915), .A2(n7914), .B1(n9567), .B2(P1_U3086), .C1(
        n7935), .C2(n7913), .ZN(P1_U3327) );
  NAND2_X1 U9658 ( .A1(n7916), .A2(n7777), .ZN(n7919) );
  NAND2_X1 U9659 ( .A1(n9401), .A2(n6252), .ZN(n7921) );
  NAND2_X1 U9660 ( .A1(n9063), .A2(n7709), .ZN(n7920) );
  NAND2_X1 U9661 ( .A1(n7921), .A2(n7920), .ZN(n7923) );
  XNOR2_X1 U9662 ( .A(n7923), .B(n7922), .ZN(n7926) );
  AOI22_X1 U9663 ( .A1(n9401), .A2(n7709), .B1(n7924), .B2(n9063), .ZN(n7925)
         );
  NAND2_X1 U9664 ( .A1(n7926), .A2(n7925), .ZN(n7933) );
  OAI21_X1 U9665 ( .B1(n7926), .B2(n7925), .A(n7933), .ZN(n8936) );
  INV_X1 U9666 ( .A(n8936), .ZN(n7932) );
  INV_X1 U9667 ( .A(n7927), .ZN(n7930) );
  INV_X1 U9668 ( .A(n7928), .ZN(n7929) );
  AND2_X1 U9669 ( .A1(n7930), .A2(n7929), .ZN(n8937) );
  INV_X1 U9670 ( .A(n8937), .ZN(n7931) );
  NAND2_X1 U9671 ( .A1(n7934), .A2(n7777), .ZN(n7937) );
  OR2_X1 U9672 ( .A1(n4347), .A2(n7935), .ZN(n7936) );
  INV_X1 U9673 ( .A(n9395), .ZN(n9200) );
  INV_X1 U9674 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n7940) );
  INV_X1 U9675 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n7938) );
  OR2_X1 U9676 ( .A1(n8177), .A2(n7938), .ZN(n7939) );
  OAI21_X1 U9677 ( .B1(n7941), .B2(n7940), .A(n7939), .ZN(n7947) );
  INV_X1 U9678 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n7942) );
  INV_X1 U9679 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n7944) );
  OR2_X1 U9680 ( .A1(n8179), .A2(n7944), .ZN(n7945) );
  OAI21_X1 U9681 ( .B1(n6262), .B2(n9244), .A(n7945), .ZN(n7946) );
  INV_X2 U9682 ( .A(n9226), .ZN(n9199) );
  OAI22_X1 U9683 ( .A1(n9200), .A2(n7948), .B1(n9199), .B2(n6158), .ZN(n7952)
         );
  AOI22_X1 U9684 ( .A1(n9395), .A2(n6252), .B1(n7709), .B2(n9226), .ZN(n7950)
         );
  XNOR2_X1 U9685 ( .A(n7950), .B(n7949), .ZN(n7951) );
  XNOR2_X1 U9686 ( .A(n7954), .B(n7953), .ZN(n7964) );
  INV_X1 U9687 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n7956) );
  INV_X1 U9688 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n7955) );
  OAI22_X1 U9689 ( .A1(n7941), .A2(n7956), .B1(n8177), .B2(n7955), .ZN(n7960)
         );
  NAND2_X1 U9690 ( .A1(n7957), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n9203) );
  INV_X1 U9691 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n7958) );
  OAI22_X1 U9692 ( .A1(n6262), .A2(n9203), .B1(n8179), .B2(n7958), .ZN(n7959)
         );
  OAI22_X1 U9693 ( .A1(n8313), .A2(n9162), .B1(n9198), .B2(n9017), .ZN(n9238)
         );
  AOI22_X1 U9694 ( .A1(n9018), .A2(n9238), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3086), .ZN(n7961) );
  OAI21_X1 U9695 ( .B1(n9021), .B2(n9244), .A(n7961), .ZN(n7962) );
  AOI21_X1 U9696 ( .B1(n9395), .B2(n9023), .A(n7962), .ZN(n7963) );
  OAI21_X1 U9697 ( .B1(n7964), .B2(n9036), .A(n7963), .ZN(P1_U3220) );
  INV_X1 U9698 ( .A(n8087), .ZN(n8090) );
  MUX2_X1 U9699 ( .A(n8869), .B(n8689), .S(n8085), .Z(n8092) );
  INV_X1 U9700 ( .A(n7965), .ZN(n8074) );
  INV_X1 U9701 ( .A(n8085), .ZN(n8098) );
  NAND3_X1 U9702 ( .A1(n7972), .A2(n7973), .A3(n8098), .ZN(n7999) );
  NAND3_X1 U9703 ( .A1(n7967), .A2(n7966), .A3(n8085), .ZN(n7968) );
  OAI21_X1 U9704 ( .B1(n8010), .B2(n7970), .A(n7969), .ZN(n7976) );
  AND2_X1 U9705 ( .A1(n7972), .A2(n7971), .ZN(n7974) );
  OAI211_X1 U9706 ( .C1(n8010), .C2(n7974), .A(n7973), .B(n8016), .ZN(n7975)
         );
  MUX2_X1 U9707 ( .A(n7976), .B(n7975), .S(n8085), .Z(n7977) );
  NOR2_X1 U9708 ( .A1(n7977), .A2(n8145), .ZN(n8025) );
  OAI22_X1 U9709 ( .A1(n7980), .A2(n7979), .B1(n8169), .B2(n7978), .ZN(n7986)
         );
  INV_X1 U9710 ( .A(n7981), .ZN(n7984) );
  OAI21_X1 U9711 ( .B1(n8135), .B2(n7982), .A(n5516), .ZN(n7983) );
  MUX2_X1 U9712 ( .A(n7984), .B(n7983), .S(n8085), .Z(n7985) );
  AOI211_X1 U9713 ( .C1(n5516), .C2(n7986), .A(n10039), .B(n7985), .ZN(n7993)
         );
  NAND2_X1 U9714 ( .A1(n7994), .A2(n7987), .ZN(n7990) );
  NAND2_X1 U9715 ( .A1(n8601), .A2(n10064), .ZN(n8001) );
  NAND2_X1 U9716 ( .A1(n7988), .A2(n8001), .ZN(n7989) );
  MUX2_X1 U9717 ( .A(n7990), .B(n7989), .S(n8085), .Z(n7992) );
  OAI21_X1 U9718 ( .B1(n7993), .B2(n7992), .A(n7991), .ZN(n8005) );
  INV_X1 U9719 ( .A(n7994), .ZN(n7996) );
  OAI211_X1 U9720 ( .C1(n8005), .C2(n7996), .A(n8006), .B(n7995), .ZN(n7997)
         );
  AND2_X1 U9721 ( .A1(n7997), .A2(n8003), .ZN(n8000) );
  INV_X1 U9722 ( .A(n7998), .ZN(n8007) );
  OAI21_X1 U9723 ( .B1(n8000), .B2(n8007), .A(n7999), .ZN(n8014) );
  INV_X1 U9724 ( .A(n8001), .ZN(n8004) );
  OAI211_X1 U9725 ( .C1(n8005), .C2(n8004), .A(n8003), .B(n8002), .ZN(n8012)
         );
  INV_X1 U9726 ( .A(n8006), .ZN(n8009) );
  AOI211_X1 U9727 ( .C1(n8009), .C2(n8008), .A(n8085), .B(n8007), .ZN(n8011)
         );
  AOI211_X1 U9728 ( .C1(n8012), .C2(n8011), .A(n8010), .B(n8139), .ZN(n8013)
         );
  INV_X1 U9729 ( .A(n8018), .ZN(n8015) );
  AOI21_X1 U9730 ( .B1(n8017), .B2(n8016), .A(n8015), .ZN(n8022) );
  INV_X1 U9731 ( .A(n8017), .ZN(n8020) );
  OAI21_X1 U9732 ( .B1(n8020), .B2(n8019), .A(n8018), .ZN(n8021) );
  MUX2_X1 U9733 ( .A(n8022), .B(n8021), .S(n8085), .Z(n8023) );
  NAND2_X1 U9734 ( .A1(n10113), .A2(n8026), .ZN(n8028) );
  MUX2_X1 U9735 ( .A(n8028), .B(n8027), .S(n8085), .Z(n8029) );
  MUX2_X1 U9736 ( .A(n8032), .B(n8031), .S(n8085), .Z(n8033) );
  INV_X1 U9737 ( .A(n8035), .ZN(n8036) );
  MUX2_X1 U9738 ( .A(n8037), .B(n8036), .S(n8085), .Z(n8038) );
  MUX2_X1 U9739 ( .A(n8040), .B(n8039), .S(n8085), .Z(n8041) );
  NAND3_X1 U9740 ( .A1(n8042), .A2(n8150), .A3(n8041), .ZN(n8047) );
  MUX2_X1 U9741 ( .A(n8044), .B(n8043), .S(n8085), .Z(n8045) );
  NAND3_X1 U9742 ( .A1(n8047), .A2(n8046), .A3(n8045), .ZN(n8052) );
  INV_X1 U9743 ( .A(n8800), .ZN(n8048) );
  AOI21_X1 U9744 ( .B1(n8052), .B2(n8132), .A(n8048), .ZN(n8054) );
  AND2_X1 U9745 ( .A1(n8800), .A2(n8049), .ZN(n8133) );
  INV_X1 U9746 ( .A(n8801), .ZN(n8051) );
  INV_X1 U9747 ( .A(n8050), .ZN(n8055) );
  AOI211_X1 U9748 ( .C1(n8052), .C2(n8133), .A(n8051), .B(n8055), .ZN(n8053)
         );
  MUX2_X1 U9749 ( .A(n8054), .B(n8053), .S(n8085), .Z(n8062) );
  INV_X1 U9750 ( .A(n8060), .ZN(n8056) );
  AOI211_X1 U9751 ( .C1(n8062), .C2(n8059), .A(n8056), .B(n8055), .ZN(n8058)
         );
  INV_X1 U9752 ( .A(n8065), .ZN(n8057) );
  INV_X1 U9753 ( .A(n8059), .ZN(n8061) );
  OAI21_X1 U9754 ( .B1(n8062), .B2(n8061), .A(n8060), .ZN(n8066) );
  INV_X1 U9755 ( .A(n8063), .ZN(n8064) );
  AOI21_X1 U9756 ( .B1(n8066), .B2(n8065), .A(n8064), .ZN(n8067) );
  MUX2_X1 U9757 ( .A(n8069), .B(n8068), .S(n8085), .Z(n8070) );
  NAND3_X1 U9758 ( .A1(n8071), .A2(n8721), .A3(n8130), .ZN(n8073) );
  NAND2_X1 U9759 ( .A1(n4400), .A2(n8130), .ZN(n8075) );
  AOI22_X1 U9760 ( .A1(n4386), .A2(n8076), .B1(n8129), .B2(n8075), .ZN(n8077)
         );
  INV_X1 U9761 ( .A(n8721), .ZN(n8156) );
  INV_X1 U9762 ( .A(n8080), .ZN(n8078) );
  NAND2_X1 U9763 ( .A1(n8078), .A2(n8079), .ZN(n8701) );
  INV_X1 U9764 ( .A(n8079), .ZN(n8081) );
  MUX2_X1 U9765 ( .A(n8081), .B(n8080), .S(n8085), .Z(n8082) );
  NOR2_X1 U9766 ( .A1(n8084), .A2(n8703), .ZN(n8086) );
  MUX2_X1 U9767 ( .A(n4592), .B(n8086), .S(n8085), .Z(n8088) );
  INV_X1 U9768 ( .A(n8101), .ZN(n8094) );
  AOI22_X1 U9769 ( .A1(n8318), .A2(n8102), .B1(P1_DATAO_REG_30__SCAN_IN), .B2(
        n5489), .ZN(n8866) );
  INV_X1 U9770 ( .A(n8866), .ZN(n8822) );
  INV_X1 U9771 ( .A(n8585), .ZN(n8091) );
  NAND2_X1 U9772 ( .A1(n8822), .A2(n8091), .ZN(n8096) );
  NAND2_X1 U9773 ( .A1(n8096), .A2(n8121), .ZN(n8159) );
  INV_X1 U9774 ( .A(n8096), .ZN(n8097) );
  NAND2_X1 U9775 ( .A1(n8866), .A2(n8585), .ZN(n8119) );
  OAI21_X1 U9776 ( .B1(n8097), .B2(n8098), .A(n8119), .ZN(n8113) );
  NAND2_X1 U9777 ( .A1(n8119), .A2(n8123), .ZN(n8160) );
  NOR3_X1 U9778 ( .A1(n8099), .A2(n8098), .A3(n8160), .ZN(n8100) );
  OAI21_X1 U9779 ( .B1(n8101), .B2(n8869), .A(n8100), .ZN(n8112) );
  AOI22_X1 U9780 ( .A1(n8172), .A2(n8102), .B1(n5489), .B2(
        P1_DATAO_REG_31__SCAN_IN), .ZN(n8678) );
  INV_X1 U9781 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n8108) );
  NAND2_X1 U9782 ( .A1(n8103), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n8106) );
  INV_X1 U9783 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n8104) );
  OR2_X1 U9784 ( .A1(n5104), .A2(n8104), .ZN(n8105) );
  OAI211_X1 U9785 ( .C1(n8108), .C2(n8107), .A(n8106), .B(n8105), .ZN(n8109)
         );
  INV_X1 U9786 ( .A(n8109), .ZN(n8110) );
  NAND2_X1 U9787 ( .A1(n8111), .A2(n8110), .ZN(n8675) );
  NAND2_X1 U9788 ( .A1(n8678), .A2(n8675), .ZN(n8128) );
  OAI211_X1 U9789 ( .C1(n8114), .C2(n8113), .A(n8112), .B(n8128), .ZN(n8116)
         );
  NAND2_X1 U9790 ( .A1(n8116), .A2(n8115), .ZN(n8165) );
  INV_X1 U9791 ( .A(n8123), .ZN(n8118) );
  INV_X1 U9792 ( .A(n8159), .ZN(n8117) );
  AOI21_X1 U9793 ( .B1(n8120), .B2(n8119), .A(n8678), .ZN(n8127) );
  NAND2_X1 U9794 ( .A1(n8122), .A2(n8121), .ZN(n8124) );
  AOI211_X1 U9795 ( .C1(n8124), .C2(n8123), .A(n8822), .B(n8675), .ZN(n8126)
         );
  INV_X1 U9796 ( .A(n8128), .ZN(n8161) );
  INV_X1 U9797 ( .A(n8701), .ZN(n8698) );
  NAND2_X1 U9798 ( .A1(n8130), .A2(n8129), .ZN(n8729) );
  NAND2_X1 U9799 ( .A1(n4400), .A2(n8725), .ZN(n8739) );
  INV_X1 U9800 ( .A(n8131), .ZN(n8750) );
  INV_X1 U9801 ( .A(n8789), .ZN(n8788) );
  INV_X1 U9802 ( .A(n8132), .ZN(n8153) );
  INV_X1 U9803 ( .A(n8133), .ZN(n8152) );
  NOR4_X1 U9804 ( .A1(n5133), .A2(n8135), .A3(n10039), .A4(n8134), .ZN(n8137)
         );
  NAND4_X1 U9805 ( .A1(n8137), .A2(n4367), .A3(n9542), .A4(n8136), .ZN(n8140)
         );
  NOR3_X1 U9806 ( .A1(n8140), .A2(n8139), .A3(n8138), .ZN(n8144) );
  NAND4_X1 U9807 ( .A1(n8144), .A2(n8143), .A3(n8142), .A4(n8141), .ZN(n8147)
         );
  NOR4_X1 U9808 ( .A1(n8147), .A2(n8146), .A3(n4493), .A4(n8145), .ZN(n8148)
         );
  NAND4_X1 U9809 ( .A1(n8150), .A2(n8149), .A3(n8148), .A4(n5265), .ZN(n8151)
         );
  NOR4_X1 U9810 ( .A1(n8788), .A2(n8153), .A3(n8152), .A4(n8151), .ZN(n8154)
         );
  NAND4_X1 U9811 ( .A1(n8750), .A2(n4715), .A3(n8775), .A4(n8154), .ZN(n8155)
         );
  NOR4_X1 U9812 ( .A1(n8156), .A2(n8729), .A3(n8739), .A4(n8155), .ZN(n8157)
         );
  NAND4_X1 U9813 ( .A1(n8482), .A2(n8698), .A3(n8157), .A4(n4590), .ZN(n8158)
         );
  NOR4_X1 U9814 ( .A1(n8161), .A2(n8160), .A3(n8159), .A4(n8158), .ZN(n8162)
         );
  NOR2_X1 U9815 ( .A1(n8163), .A2(n8162), .ZN(n8164) );
  INV_X1 U9816 ( .A(n8678), .ZN(n8861) );
  NAND3_X1 U9817 ( .A1(n8167), .A2(n8166), .A3(n5537), .ZN(n8168) );
  OAI211_X1 U9818 ( .C1(n8169), .C2(n8171), .A(n8168), .B(P2_B_REG_SCAN_IN), 
        .ZN(n8170) );
  MUX2_X1 U9819 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n8172), .S(n4962), .Z(n8174) );
  AOI211_X1 U9820 ( .C1(n8455), .C2(n4349), .A(n8464), .B(n8175), .ZN(n8461)
         );
  INV_X1 U9821 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n8182) );
  INV_X1 U9822 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n8176) );
  OR2_X1 U9823 ( .A1(n8177), .A2(n8176), .ZN(n8181) );
  INV_X1 U9824 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n8178) );
  OR2_X1 U9825 ( .A1(n8179), .A2(n8178), .ZN(n8180) );
  OAI211_X1 U9826 ( .C1(n7941), .C2(n8182), .A(n8181), .B(n8180), .ZN(n9223)
         );
  OR2_X1 U9827 ( .A1(n9426), .A2(n9185), .ZN(n8275) );
  NAND2_X1 U9828 ( .A1(n8379), .A2(n8275), .ZN(n8329) );
  NAND2_X1 U9829 ( .A1(n8355), .A2(n8356), .ZN(n8403) );
  NAND2_X1 U9830 ( .A1(n8183), .A2(n9181), .ZN(n9209) );
  NAND2_X1 U9831 ( .A1(n9435), .A2(n9177), .ZN(n9206) );
  NAND2_X1 U9832 ( .A1(n9209), .A2(n9206), .ZN(n8337) );
  MUX2_X1 U9833 ( .A(n8403), .B(n8337), .S(n8264), .Z(n8274) );
  AOI21_X1 U9834 ( .B1(n9206), .B2(n9370), .A(n8264), .ZN(n8186) );
  INV_X1 U9835 ( .A(n8263), .ZN(n8184) );
  NAND2_X1 U9836 ( .A1(n8356), .A2(n8328), .ZN(n9207) );
  NAND3_X1 U9837 ( .A1(n9206), .A2(n8322), .A3(n9175), .ZN(n8185) );
  OAI21_X1 U9838 ( .B1(n8186), .B2(n9207), .A(n8185), .ZN(n8271) );
  NAND2_X1 U9839 ( .A1(n8435), .A2(n8187), .ZN(n8257) );
  NAND2_X1 U9840 ( .A1(n8252), .A2(n8247), .ZN(n8431) );
  NOR2_X1 U9841 ( .A1(n8431), .A2(n8248), .ZN(n8188) );
  OR3_X1 U9842 ( .A1(n8257), .A2(n9549), .A3(n8188), .ZN(n8440) );
  AND2_X1 U9843 ( .A1(n8363), .A2(n8264), .ZN(n8189) );
  NAND2_X1 U9844 ( .A1(n8190), .A2(n8189), .ZN(n8227) );
  NAND2_X1 U9845 ( .A1(n8191), .A2(n8201), .ZN(n8195) );
  AND2_X1 U9846 ( .A1(n8196), .A2(n8413), .ZN(n8194) );
  NAND4_X1 U9847 ( .A1(n8200), .A2(n8420), .A3(n8192), .A4(n8264), .ZN(n8193)
         );
  AOI21_X1 U9848 ( .B1(n8195), .B2(n8194), .A(n8193), .ZN(n8218) );
  AND2_X1 U9849 ( .A1(n8197), .A2(n8196), .ZN(n8198) );
  NAND2_X1 U9850 ( .A1(n8199), .A2(n8198), .ZN(n8408) );
  AND2_X1 U9851 ( .A1(n8201), .A2(n8200), .ZN(n8411) );
  NAND4_X1 U9852 ( .A1(n8413), .A2(n8416), .A3(n8412), .A4(n8322), .ZN(n8202)
         );
  AOI21_X1 U9853 ( .B1(n8408), .B2(n8411), .A(n8202), .ZN(n8217) );
  NAND2_X1 U9854 ( .A1(n8203), .A2(n8264), .ZN(n8205) );
  OAI22_X1 U9855 ( .A1(n8205), .A2(n9861), .B1(n8322), .B2(n9076), .ZN(n8204)
         );
  NAND2_X1 U9856 ( .A1(n8204), .A2(n6642), .ZN(n8215) );
  OAI21_X1 U9857 ( .B1(n8205), .B2(n9076), .A(n8210), .ZN(n8208) );
  NAND2_X1 U9858 ( .A1(n9077), .A2(n8322), .ZN(n8211) );
  OAI21_X1 U9859 ( .B1(n8211), .B2(n8206), .A(n9861), .ZN(n8207) );
  NAND2_X1 U9860 ( .A1(n8208), .A2(n8207), .ZN(n8214) );
  NAND2_X1 U9861 ( .A1(n9076), .A2(n8322), .ZN(n8209) );
  OAI21_X1 U9862 ( .B1(n8211), .B2(n8210), .A(n8209), .ZN(n8212) );
  NAND2_X1 U9863 ( .A1(n8212), .A2(n6643), .ZN(n8213) );
  NAND4_X1 U9864 ( .A1(n8215), .A2(n8214), .A3(n8363), .A4(n8213), .ZN(n8216)
         );
  OR3_X1 U9865 ( .A1(n8218), .A2(n8217), .A3(n8216), .ZN(n8221) );
  OAI21_X1 U9866 ( .B1(n8219), .B2(n8264), .A(n8227), .ZN(n8220) );
  NAND2_X1 U9867 ( .A1(n8221), .A2(n8220), .ZN(n8226) );
  NAND2_X1 U9868 ( .A1(n8229), .A2(n8222), .ZN(n8223) );
  MUX2_X1 U9869 ( .A(n8223), .B(n8366), .S(n8322), .Z(n8224) );
  INV_X1 U9870 ( .A(n8224), .ZN(n8225) );
  OAI211_X1 U9871 ( .C1(n8228), .C2(n8227), .A(n8226), .B(n8225), .ZN(n8234)
         );
  NAND2_X1 U9872 ( .A1(n8234), .A2(n8229), .ZN(n8230) );
  NAND2_X1 U9873 ( .A1(n8236), .A2(n9745), .ZN(n8429) );
  AOI21_X1 U9874 ( .B1(n8230), .B2(n8422), .A(n8429), .ZN(n8231) );
  NAND2_X1 U9875 ( .A1(n8239), .A2(n8235), .ZN(n8427) );
  OAI21_X1 U9876 ( .B1(n8231), .B2(n8427), .A(n8432), .ZN(n8242) );
  AOI21_X1 U9877 ( .B1(n8234), .B2(n8233), .A(n8232), .ZN(n8238) );
  NAND2_X1 U9878 ( .A1(n8235), .A2(n8422), .ZN(n8237) );
  OAI211_X1 U9879 ( .C1(n8238), .C2(n8237), .A(n8432), .B(n8236), .ZN(n8240)
         );
  NAND2_X1 U9880 ( .A1(n8240), .A2(n8239), .ZN(n8241) );
  MUX2_X1 U9881 ( .A(n8242), .B(n8241), .S(n8264), .Z(n8246) );
  NOR2_X1 U9882 ( .A1(n8246), .A2(n8431), .ZN(n8244) );
  NAND2_X1 U9883 ( .A1(n8435), .A2(n8436), .ZN(n8243) );
  OAI211_X1 U9884 ( .C1(n8440), .C2(n8244), .A(n8256), .B(n8243), .ZN(n8245)
         );
  INV_X1 U9885 ( .A(n8245), .ZN(n8255) );
  INV_X1 U9886 ( .A(n8246), .ZN(n8250) );
  INV_X1 U9887 ( .A(n8247), .ZN(n8249) );
  OAI211_X1 U9888 ( .C1(n8250), .C2(n8249), .A(n8373), .B(n8248), .ZN(n8253)
         );
  NAND4_X1 U9889 ( .A1(n8253), .A2(n8256), .A3(n8252), .A4(n8251), .ZN(n8254)
         );
  MUX2_X1 U9890 ( .A(n8255), .B(n8254), .S(n8322), .Z(n8259) );
  NAND3_X1 U9891 ( .A1(n8257), .A2(n8322), .A3(n8256), .ZN(n8258) );
  AOI21_X1 U9892 ( .B1(n8259), .B2(n8258), .A(n8376), .ZN(n8269) );
  NAND2_X1 U9893 ( .A1(n8262), .A2(n8260), .ZN(n8434) );
  NAND2_X1 U9894 ( .A1(n8324), .A2(n8443), .ZN(n8261) );
  MUX2_X1 U9895 ( .A(n8434), .B(n8261), .S(n8322), .Z(n8268) );
  NAND2_X1 U9896 ( .A1(n8328), .A2(n8262), .ZN(n8446) );
  NAND2_X1 U9897 ( .A1(n8446), .A2(n8322), .ZN(n8266) );
  NAND2_X1 U9898 ( .A1(n8184), .A2(n9176), .ZN(n8445) );
  NAND2_X1 U9899 ( .A1(n8445), .A2(n8324), .ZN(n8404) );
  AND2_X1 U9900 ( .A1(n8266), .A2(n8265), .ZN(n8267) );
  AND2_X1 U9901 ( .A1(n8271), .A2(n8270), .ZN(n8273) );
  MUX2_X1 U9902 ( .A(n8355), .B(n9209), .S(n8322), .Z(n8272) );
  OAI21_X1 U9903 ( .B1(n8274), .B2(n8273), .A(n8272), .ZN(n8276) );
  NAND2_X1 U9904 ( .A1(n9426), .A2(n9185), .ZN(n9210) );
  AOI22_X1 U9905 ( .A1(n8329), .A2(n8264), .B1(n8276), .B2(n9326), .ZN(n8279)
         );
  INV_X1 U9906 ( .A(n9211), .ZN(n8278) );
  AND2_X1 U9907 ( .A1(n9211), .A2(n9210), .ZN(n8277) );
  NAND2_X1 U9908 ( .A1(n9416), .A2(n9189), .ZN(n8334) );
  OR3_X1 U9909 ( .A1(n9421), .A2(n8264), .A3(n9188), .ZN(n8280) );
  NAND3_X1 U9910 ( .A1(n8281), .A2(n9212), .A3(n8280), .ZN(n8283) );
  MUX2_X1 U9911 ( .A(n8334), .B(n9213), .S(n8264), .Z(n8282) );
  NAND2_X1 U9912 ( .A1(n8283), .A2(n8282), .ZN(n8290) );
  NAND2_X1 U9913 ( .A1(n9411), .A2(n9193), .ZN(n9215) );
  NAND2_X1 U9914 ( .A1(n8290), .A2(n9215), .ZN(n8285) );
  OR2_X1 U9915 ( .A1(n9406), .A2(n9195), .ZN(n8382) );
  NAND2_X1 U9916 ( .A1(n8285), .A2(n8284), .ZN(n8286) );
  NAND2_X1 U9917 ( .A1(n9406), .A2(n9195), .ZN(n9216) );
  NAND2_X1 U9918 ( .A1(n8286), .A2(n9216), .ZN(n8289) );
  OR2_X1 U9919 ( .A1(n9401), .A2(n9198), .ZN(n8386) );
  NAND2_X1 U9920 ( .A1(n8290), .A2(n8383), .ZN(n8291) );
  NAND3_X1 U9921 ( .A1(n8291), .A2(n9216), .A3(n9215), .ZN(n8292) );
  NAND2_X1 U9922 ( .A1(n8292), .A2(n8382), .ZN(n8294) );
  NAND2_X1 U9923 ( .A1(n9395), .A2(n9199), .ZN(n9219) );
  NAND2_X1 U9924 ( .A1(n9401), .A2(n9198), .ZN(n8385) );
  AND3_X1 U9925 ( .A1(n9219), .A2(n8322), .A3(n8385), .ZN(n8293) );
  NAND2_X1 U9926 ( .A1(n8294), .A2(n8293), .ZN(n8307) );
  NAND2_X1 U9927 ( .A1(n9063), .A2(n8322), .ZN(n8295) );
  OAI22_X1 U9928 ( .A1(n9401), .A2(n8295), .B1(n8264), .B2(n9199), .ZN(n8299)
         );
  NAND2_X1 U9929 ( .A1(n9198), .A2(n8264), .ZN(n8300) );
  OAI21_X1 U9930 ( .B1(n9226), .B2(n8300), .A(n9401), .ZN(n8298) );
  NOR2_X1 U9931 ( .A1(n8295), .A2(n9199), .ZN(n8296) );
  OR2_X1 U9932 ( .A1(n9401), .A2(n8296), .ZN(n8297) );
  AOI22_X1 U9933 ( .A1(n9200), .A2(n8299), .B1(n8298), .B2(n8297), .ZN(n8305)
         );
  INV_X1 U9934 ( .A(n8300), .ZN(n8301) );
  NAND2_X1 U9935 ( .A1(n9401), .A2(n8301), .ZN(n8302) );
  OAI21_X1 U9936 ( .B1(n9226), .B2(n8322), .A(n8302), .ZN(n8303) );
  NAND2_X1 U9937 ( .A1(n8303), .A2(n9395), .ZN(n8304) );
  NAND3_X1 U9938 ( .A1(n8308), .A2(n8307), .A3(n8306), .ZN(n8317) );
  NAND2_X1 U9939 ( .A1(n8309), .A2(n7777), .ZN(n8312) );
  OR2_X1 U9940 ( .A1(n4347), .A2(n8310), .ZN(n8311) );
  NOR2_X1 U9941 ( .A1(n9390), .A2(n8313), .ZN(n8344) );
  INV_X1 U9942 ( .A(n8344), .ZN(n8314) );
  AND2_X1 U9943 ( .A1(n9390), .A2(n8313), .ZN(n8315) );
  INV_X1 U9944 ( .A(n8315), .ZN(n8333) );
  AND2_X2 U9945 ( .A1(n8314), .A2(n8333), .ZN(n9221) );
  MUX2_X1 U9946 ( .A(n8315), .B(n8344), .S(n8322), .Z(n8316) );
  NAND2_X1 U9947 ( .A1(n8318), .A2(n7777), .ZN(n8321) );
  OR2_X1 U9948 ( .A1(n4347), .A2(n8319), .ZN(n8320) );
  INV_X1 U9949 ( .A(n9223), .ZN(n8342) );
  NOR2_X1 U9950 ( .A1(n8323), .A2(n8455), .ZN(n8396) );
  OAI21_X1 U9951 ( .B1(n6070), .B2(n4351), .A(n8396), .ZN(n8460) );
  INV_X1 U9952 ( .A(n8377), .ZN(n8326) );
  INV_X1 U9953 ( .A(n8324), .ZN(n8325) );
  NAND2_X1 U9954 ( .A1(n9205), .A2(n8328), .ZN(n9355) );
  NAND2_X1 U9955 ( .A1(n8329), .A2(n9211), .ZN(n8330) );
  NAND2_X1 U9956 ( .A1(n9213), .A2(n8330), .ZN(n8331) );
  NAND2_X1 U9957 ( .A1(n8331), .A2(n8334), .ZN(n8332) );
  NAND2_X1 U9958 ( .A1(n8383), .A2(n8332), .ZN(n8402) );
  NOR3_X1 U9959 ( .A1(n9355), .A2(n8403), .A3(n8402), .ZN(n8350) );
  NAND2_X1 U9960 ( .A1(n9156), .A2(n8342), .ZN(n8390) );
  NAND2_X1 U9961 ( .A1(n8390), .A2(n8333), .ZN(n8347) );
  INV_X1 U9962 ( .A(n8347), .ZN(n8341) );
  AND2_X1 U9963 ( .A1(n8386), .A2(n8382), .ZN(n8343) );
  NAND2_X1 U9964 ( .A1(n9211), .A2(n9210), .ZN(n8336) );
  INV_X1 U9965 ( .A(n8334), .ZN(n8335) );
  AOI211_X1 U9966 ( .C1(n8355), .C2(n8337), .A(n8336), .B(n8335), .ZN(n8338)
         );
  OAI21_X1 U9967 ( .B1(n8338), .B2(n8402), .A(n9215), .ZN(n8340) );
  INV_X1 U9968 ( .A(n8385), .ZN(n9218) );
  INV_X1 U9969 ( .A(n9219), .ZN(n8339) );
  AOI211_X1 U9970 ( .C1(n8343), .C2(n8340), .A(n9218), .B(n8339), .ZN(n8346)
         );
  NAND3_X1 U9971 ( .A1(n8341), .A2(n8346), .A3(n9216), .ZN(n8401) );
  OR2_X1 U9972 ( .A1(n9156), .A2(n8342), .ZN(n8391) );
  INV_X1 U9973 ( .A(n8391), .ZN(n8452) );
  INV_X1 U9974 ( .A(n8343), .ZN(n8345) );
  INV_X1 U9975 ( .A(n8387), .ZN(n9220) );
  AOI211_X1 U9976 ( .C1(n8346), .C2(n8345), .A(n9220), .B(n8344), .ZN(n8348)
         );
  NOR2_X1 U9977 ( .A1(n8348), .A2(n8347), .ZN(n8451) );
  AOI21_X1 U9978 ( .B1(n8452), .B2(n9163), .A(n8451), .ZN(n8349) );
  OAI21_X1 U9979 ( .B1(n8350), .B2(n8401), .A(n8349), .ZN(n8352) );
  INV_X1 U9980 ( .A(n8455), .ZN(n8351) );
  OAI211_X1 U9981 ( .C1(n9387), .C2(n9163), .A(n8352), .B(n8351), .ZN(n8354)
         );
  NAND3_X1 U9982 ( .A1(n8354), .A2(n8353), .A3(n4351), .ZN(n8395) );
  INV_X1 U9983 ( .A(n9221), .ZN(n8389) );
  NOR2_X1 U9984 ( .A1(n8357), .A2(n6151), .ZN(n8360) );
  NAND4_X1 U9985 ( .A1(n8360), .A2(n9796), .A3(n8359), .A4(n9815), .ZN(n8362)
         );
  NOR2_X1 U9986 ( .A1(n8362), .A2(n8361), .ZN(n8364) );
  NAND4_X1 U9987 ( .A1(n8365), .A2(n8364), .A3(n9781), .A4(n8363), .ZN(n8367)
         );
  NOR2_X1 U9988 ( .A1(n8367), .A2(n8366), .ZN(n8368) );
  NAND4_X1 U9989 ( .A1(n9744), .A2(n8417), .A3(n8369), .A4(n8368), .ZN(n8370)
         );
  NOR2_X1 U9990 ( .A1(n9735), .A2(n8370), .ZN(n8371) );
  NAND4_X1 U9991 ( .A1(n9556), .A2(n8373), .A3(n8372), .A4(n8371), .ZN(n8374)
         );
  NOR4_X1 U9992 ( .A1(n8377), .A2(n8376), .A3(n8375), .A4(n8374), .ZN(n8378)
         );
  NAND4_X1 U9993 ( .A1(n9340), .A2(n9356), .A3(n9371), .A4(n8378), .ZN(n8381)
         );
  NAND2_X1 U9994 ( .A1(n8379), .A2(n9211), .ZN(n9304) );
  INV_X1 U9995 ( .A(n9326), .ZN(n8380) );
  NAND2_X1 U9996 ( .A1(n8382), .A2(n9216), .ZN(n9265) );
  INV_X1 U9997 ( .A(n9265), .ZN(n8384) );
  NAND4_X1 U9998 ( .A1(n4380), .A2(n8384), .A3(n4352), .A4(n9212), .ZN(n8388)
         );
  NAND2_X1 U9999 ( .A1(n8386), .A2(n8385), .ZN(n9217) );
  NAND2_X1 U10000 ( .A1(n8387), .A2(n9219), .ZN(n9242) );
  OR4_X1 U10001 ( .A1(n8389), .A2(n8388), .A3(n9217), .A4(n9242), .ZN(n8393)
         );
  NAND3_X1 U10002 ( .A1(n8351), .A2(n4351), .A3(n4883), .ZN(n8392) );
  INV_X1 U10003 ( .A(n8397), .ZN(n8394) );
  NAND2_X1 U10004 ( .A1(n8395), .A2(n8394), .ZN(n8400) );
  NAND2_X1 U10005 ( .A1(n8396), .A2(n8464), .ZN(n8398) );
  AOI21_X1 U10006 ( .B1(n8398), .B2(n6151), .A(n8397), .ZN(n8399) );
  INV_X1 U10007 ( .A(n8401), .ZN(n8454) );
  INV_X1 U10008 ( .A(n8402), .ZN(n8450) );
  INV_X1 U10009 ( .A(n8403), .ZN(n8449) );
  INV_X1 U10010 ( .A(n8404), .ZN(n8444) );
  AOI21_X1 U10011 ( .B1(n6616), .B2(n6626), .A(n8405), .ZN(n8410) );
  AND2_X1 U10012 ( .A1(n8407), .A2(n8406), .ZN(n8409) );
  AOI21_X1 U10013 ( .B1(n8410), .B2(n8409), .A(n8408), .ZN(n8415) );
  INV_X1 U10014 ( .A(n8411), .ZN(n8414) );
  OAI211_X1 U10015 ( .C1(n8415), .C2(n8414), .A(n8413), .B(n8412), .ZN(n8421)
         );
  INV_X1 U10016 ( .A(n8416), .ZN(n8419) );
  INV_X1 U10017 ( .A(n8417), .ZN(n8418) );
  AOI211_X1 U10018 ( .C1(n8421), .C2(n8420), .A(n8419), .B(n8418), .ZN(n8426)
         );
  INV_X1 U10019 ( .A(n8422), .ZN(n8425) );
  INV_X1 U10020 ( .A(n8423), .ZN(n8424) );
  NOR3_X1 U10021 ( .A1(n8426), .A2(n8425), .A3(n8424), .ZN(n8430) );
  INV_X1 U10022 ( .A(n8427), .ZN(n8428) );
  OAI21_X1 U10023 ( .B1(n8430), .B2(n8429), .A(n8428), .ZN(n8433) );
  AOI21_X1 U10024 ( .B1(n8433), .B2(n8432), .A(n8431), .ZN(n8441) );
  INV_X1 U10025 ( .A(n8434), .ZN(n8439) );
  OAI21_X1 U10026 ( .B1(n8437), .B2(n8436), .A(n8435), .ZN(n8438) );
  OAI211_X1 U10027 ( .C1(n8441), .C2(n8440), .A(n8439), .B(n8438), .ZN(n8442)
         );
  NAND3_X1 U10028 ( .A1(n8444), .A2(n8443), .A3(n8442), .ZN(n8448) );
  NAND2_X1 U10029 ( .A1(n8446), .A2(n8445), .ZN(n8447) );
  NAND4_X1 U10030 ( .A1(n8450), .A2(n8449), .A3(n8448), .A4(n8447), .ZN(n8453)
         );
  AOI211_X1 U10031 ( .C1(n8454), .C2(n8453), .A(n8452), .B(n8451), .ZN(n8456)
         );
  OAI21_X1 U10032 ( .B1(n8456), .B2(n8455), .A(n4351), .ZN(n8457) );
  XNOR2_X1 U10033 ( .A(n8457), .B(n4349), .ZN(n8458) );
  NAND3_X1 U10034 ( .A1(n8462), .A2(n9569), .A3(n9225), .ZN(n8463) );
  OAI211_X1 U10035 ( .C1(n8464), .C2(n8466), .A(n8463), .B(P1_B_REG_SCAN_IN), 
        .ZN(n8465) );
  OAI21_X1 U10036 ( .B1(n8467), .B2(n8466), .A(n8465), .ZN(P1_U3242) );
  INV_X1 U10037 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n8468) );
  OAI222_X1 U10038 ( .A1(n5572), .A2(P2_U3151), .B1(n8470), .B2(n8469), .C1(
        n8468), .C2(n8491), .ZN(P2_U3271) );
  AND2_X1 U10039 ( .A1(n8521), .A2(n8473), .ZN(n8471) );
  NAND2_X1 U10040 ( .A1(n8472), .A2(n8471), .ZN(n8481) );
  INV_X1 U10041 ( .A(n8473), .ZN(n8475) );
  OR2_X1 U10042 ( .A1(n8475), .A2(n8474), .ZN(n8479) );
  INV_X1 U10043 ( .A(n8476), .ZN(n8477) );
  NAND2_X1 U10044 ( .A1(n8477), .A2(n8703), .ZN(n8478) );
  XNOR2_X1 U10045 ( .A(n8482), .B(n5641), .ZN(n8483) );
  XNOR2_X1 U10046 ( .A(n8484), .B(n8483), .ZN(n8490) );
  NAND2_X1 U10047 ( .A1(n8563), .A2(n8683), .ZN(n8486) );
  AOI22_X1 U10048 ( .A1(n8580), .A2(n8703), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3151), .ZN(n8485) );
  OAI211_X1 U10049 ( .C1(n8487), .C2(n9537), .A(n8486), .B(n8485), .ZN(n8488)
         );
  AOI21_X1 U10050 ( .B1(n8869), .B2(n9539), .A(n8488), .ZN(n8489) );
  OAI21_X1 U10051 ( .B1(n8490), .B2(n9543), .A(n8489), .ZN(P2_U3160) );
  INV_X1 U10052 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n8492) );
  OAI222_X1 U10053 ( .A1(n8497), .A2(P2_U3151), .B1(n8494), .B2(n8493), .C1(
        n8492), .C2(n8491), .ZN(P2_U3270) );
  INV_X1 U10054 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n8499) );
  AND2_X1 U10055 ( .A1(n8496), .A2(n8495), .ZN(n8498) );
  AOI22_X1 U10056 ( .A1(n8500), .A2(n8499), .B1(n8498), .B2(n8497), .ZN(
        P2_U3377) );
  NAND2_X1 U10057 ( .A1(P2_U3151), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8667) );
  OAI21_X1 U10058 ( .B1(n9537), .B2(n8794), .A(n8667), .ZN(n8501) );
  AOI21_X1 U10059 ( .B1(n8580), .B2(n8587), .A(n8501), .ZN(n8502) );
  OAI21_X1 U10060 ( .B1(n8577), .B2(n8795), .A(n8502), .ZN(n8507) );
  INV_X1 U10061 ( .A(n8503), .ZN(n8552) );
  AOI211_X1 U10062 ( .C1(n8505), .C2(n8504), .A(n9543), .B(n8552), .ZN(n8506)
         );
  AOI211_X1 U10063 ( .C1(n8852), .C2(n9539), .A(n8507), .B(n8506), .ZN(n8508)
         );
  INV_X1 U10064 ( .A(n8508), .ZN(P2_U3159) );
  INV_X1 U10065 ( .A(n8911), .ZN(n8520) );
  INV_X1 U10066 ( .A(n8509), .ZN(n8512) );
  NOR3_X1 U10067 ( .A1(n8512), .A2(n4840), .A3(n8511), .ZN(n8515) );
  INV_X1 U10068 ( .A(n8513), .ZN(n8514) );
  OAI21_X1 U10069 ( .B1(n8515), .B2(n8514), .A(n8572), .ZN(n8519) );
  AOI22_X1 U10070 ( .A1(n8547), .A2(n8768), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3151), .ZN(n8516) );
  OAI21_X1 U10071 ( .B1(n8794), .B2(n8530), .A(n8516), .ZN(n8517) );
  AOI21_X1 U10072 ( .B1(n8771), .B2(n8563), .A(n8517), .ZN(n8518) );
  OAI211_X1 U10073 ( .C1(n8520), .C2(n8583), .A(n8519), .B(n8518), .ZN(
        P2_U3163) );
  INV_X1 U10074 ( .A(n8887), .ZN(n8535) );
  INV_X1 U10075 ( .A(n8521), .ZN(n8523) );
  NOR3_X1 U10076 ( .A1(n8524), .A2(n8523), .A3(n8522), .ZN(n8527) );
  INV_X1 U10077 ( .A(n8525), .ZN(n8526) );
  OAI21_X1 U10078 ( .B1(n8527), .B2(n8526), .A(n8572), .ZN(n8534) );
  OAI22_X1 U10079 ( .A1(n9537), .A2(n8529), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8528), .ZN(n8532) );
  NOR2_X1 U10080 ( .A1(n8530), .A2(n8714), .ZN(n8531) );
  AOI211_X1 U10081 ( .C1(n8717), .C2(n8563), .A(n8532), .B(n8531), .ZN(n8533)
         );
  OAI211_X1 U10082 ( .C1(n8535), .C2(n8583), .A(n8534), .B(n8533), .ZN(
        P2_U3165) );
  INV_X1 U10083 ( .A(n8536), .ZN(n8570) );
  AOI21_X1 U10084 ( .B1(n8538), .B2(n8537), .A(n8570), .ZN(n8546) );
  NOR2_X1 U10085 ( .A1(n8539), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8648) );
  NOR2_X1 U10086 ( .A1(n9537), .A2(n8793), .ZN(n8540) );
  AOI211_X1 U10087 ( .C1(n8580), .C2(n8588), .A(n8648), .B(n8540), .ZN(n8541)
         );
  OAI21_X1 U10088 ( .B1(n8542), .B2(n8577), .A(n8541), .ZN(n8543) );
  AOI21_X1 U10089 ( .B1(n8544), .B2(n9539), .A(n8543), .ZN(n8545) );
  OAI21_X1 U10090 ( .B1(n8546), .B2(n9543), .A(n8545), .ZN(P2_U3168) );
  AOI22_X1 U10091 ( .A1(n8547), .A2(n8754), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3151), .ZN(n8549) );
  NAND2_X1 U10092 ( .A1(n8580), .A2(n8810), .ZN(n8548) );
  OAI211_X1 U10093 ( .C1(n8577), .C2(n8783), .A(n8549), .B(n8548), .ZN(n8555)
         );
  OAI21_X1 U10094 ( .B1(n8552), .B2(n8551), .A(n8550), .ZN(n8553) );
  AOI21_X1 U10095 ( .B1(n8553), .B2(n8509), .A(n9543), .ZN(n8554) );
  AOI211_X1 U10096 ( .C1(n8917), .C2(n9539), .A(n8555), .B(n8554), .ZN(n8556)
         );
  INV_X1 U10097 ( .A(n8556), .ZN(P2_U3173) );
  INV_X1 U10098 ( .A(n8905), .ZN(n8566) );
  AOI21_X1 U10099 ( .B1(n8558), .B2(n8557), .A(n9543), .ZN(n8560) );
  NAND2_X1 U10100 ( .A1(n8560), .A2(n8559), .ZN(n8565) );
  AOI22_X1 U10101 ( .A1(n8580), .A2(n8754), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3151), .ZN(n8561) );
  OAI21_X1 U10102 ( .B1(n8731), .B2(n9537), .A(n8561), .ZN(n8562) );
  AOI21_X1 U10103 ( .B1(n8757), .B2(n8563), .A(n8562), .ZN(n8564) );
  OAI211_X1 U10104 ( .C1(n8566), .C2(n8583), .A(n8565), .B(n8564), .ZN(
        P2_U3175) );
  INV_X1 U10105 ( .A(n8567), .ZN(n8569) );
  NOR3_X1 U10106 ( .A1(n8570), .A2(n8569), .A3(n8568), .ZN(n8574) );
  INV_X1 U10107 ( .A(n8571), .ZN(n8573) );
  OAI21_X1 U10108 ( .B1(n8574), .B2(n8573), .A(n8572), .ZN(n8582) );
  OAI21_X1 U10109 ( .B1(n9537), .B2(n8576), .A(n8575), .ZN(n8579) );
  NOR2_X1 U10110 ( .A1(n8577), .A2(n8813), .ZN(n8578) );
  AOI211_X1 U10111 ( .C1(n8580), .C2(n8808), .A(n8579), .B(n8578), .ZN(n8581)
         );
  OAI211_X1 U10112 ( .C1(n8584), .C2(n8583), .A(n8582), .B(n8581), .ZN(
        P2_U3178) );
  MUX2_X1 U10113 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n8675), .S(P2_U3893), .Z(
        P2_U3522) );
  MUX2_X1 U10114 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n8585), .S(P2_U3893), .Z(
        P2_U3521) );
  MUX2_X1 U10115 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n8586), .S(P2_U3893), .Z(
        P2_U3520) );
  MUX2_X1 U10116 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n8689), .S(P2_U3893), .Z(
        P2_U3519) );
  MUX2_X1 U10117 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8703), .S(P2_U3893), .Z(
        P2_U3518) );
  MUX2_X1 U10118 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n8712), .S(P2_U3893), .Z(
        P2_U3517) );
  MUX2_X1 U10119 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n8702), .S(P2_U3893), .Z(
        P2_U3516) );
  MUX2_X1 U10120 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n8741), .S(P2_U3893), .Z(
        P2_U3515) );
  MUX2_X1 U10121 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(n8753), .S(P2_U3893), .Z(
        P2_U3514) );
  MUX2_X1 U10122 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8768), .S(P2_U3893), .Z(
        P2_U3513) );
  MUX2_X1 U10123 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n8754), .S(P2_U3893), .Z(
        P2_U3512) );
  MUX2_X1 U10124 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8767), .S(P2_U3893), .Z(
        P2_U3511) );
  MUX2_X1 U10125 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n8810), .S(P2_U3893), .Z(
        P2_U3510) );
  MUX2_X1 U10126 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n8587), .S(P2_U3893), .Z(
        P2_U3509) );
  MUX2_X1 U10127 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8808), .S(P2_U3893), .Z(
        P2_U3508) );
  MUX2_X1 U10128 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n8588), .S(P2_U3893), .Z(
        P2_U3507) );
  MUX2_X1 U10129 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n8589), .S(P2_U3893), .Z(
        P2_U3506) );
  MUX2_X1 U10130 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n8590), .S(P2_U3893), .Z(
        P2_U3505) );
  MUX2_X1 U10131 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n8591), .S(P2_U3893), .Z(
        P2_U3504) );
  MUX2_X1 U10132 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n8592), .S(P2_U3893), .Z(
        P2_U3503) );
  MUX2_X1 U10133 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n8593), .S(P2_U3893), .Z(
        P2_U3502) );
  MUX2_X1 U10134 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n8594), .S(P2_U3893), .Z(
        P2_U3501) );
  MUX2_X1 U10135 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n8595), .S(P2_U3893), .Z(
        P2_U3500) );
  MUX2_X1 U10136 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n8596), .S(P2_U3893), .Z(
        P2_U3499) );
  MUX2_X1 U10137 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n8597), .S(P2_U3893), .Z(
        P2_U3498) );
  MUX2_X1 U10138 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n8598), .S(P2_U3893), .Z(
        P2_U3497) );
  MUX2_X1 U10139 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(n8599), .S(P2_U3893), .Z(
        P2_U3496) );
  MUX2_X1 U10140 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n8600), .S(P2_U3893), .Z(
        P2_U3495) );
  MUX2_X1 U10141 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(n8601), .S(P2_U3893), .Z(
        P2_U3494) );
  MUX2_X1 U10142 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(n5101), .S(P2_U3893), .Z(
        P2_U3493) );
  MUX2_X1 U10143 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n5607), .S(P2_U3893), .Z(
        P2_U3492) );
  MUX2_X1 U10144 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(n6130), .S(P2_U3893), .Z(
        P2_U3491) );
  AOI21_X1 U10145 ( .B1(n8604), .B2(n8603), .A(n8602), .ZN(n8619) );
  OAI21_X1 U10146 ( .B1(P2_REG1_REG_15__SCAN_IN), .B2(n8606), .A(n8605), .ZN(
        n8617) );
  INV_X1 U10147 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n8615) );
  OAI21_X1 U10148 ( .B1(n8609), .B2(n8608), .A(n8607), .ZN(n8613) );
  NOR2_X1 U10149 ( .A1(n9956), .A2(n8610), .ZN(n8611) );
  AOI211_X1 U10150 ( .C1(n10029), .C2(n8613), .A(n8612), .B(n8611), .ZN(n8614)
         );
  OAI21_X1 U10151 ( .B1(n10033), .B2(n8615), .A(n8614), .ZN(n8616) );
  AOI21_X1 U10152 ( .B1(n8617), .B2(n10017), .A(n8616), .ZN(n8618) );
  OAI21_X1 U10153 ( .B1(n8619), .B2(n10024), .A(n8618), .ZN(P2_U3197) );
  AOI21_X1 U10154 ( .B1(n8622), .B2(n8621), .A(n8620), .ZN(n8638) );
  OAI21_X1 U10155 ( .B1(n8625), .B2(n8624), .A(n8623), .ZN(n8636) );
  INV_X1 U10156 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n8634) );
  OAI21_X1 U10157 ( .B1(n8628), .B2(n8627), .A(n8626), .ZN(n8632) );
  NOR2_X1 U10158 ( .A1(n9956), .A2(n8629), .ZN(n8630) );
  AOI211_X1 U10159 ( .C1(n10029), .C2(n8632), .A(n8631), .B(n8630), .ZN(n8633)
         );
  OAI21_X1 U10160 ( .B1(n10033), .B2(n8634), .A(n8633), .ZN(n8635) );
  AOI21_X1 U10161 ( .B1(n8636), .B2(n10017), .A(n8635), .ZN(n8637) );
  OAI21_X1 U10162 ( .B1(n8638), .B2(n10024), .A(n8637), .ZN(P2_U3198) );
  AOI21_X1 U10163 ( .B1(n7662), .B2(n8640), .A(n8639), .ZN(n8655) );
  OAI21_X1 U10164 ( .B1(P2_REG1_REG_17__SCAN_IN), .B2(n8642), .A(n8641), .ZN(
        n8653) );
  INV_X1 U10165 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n8651) );
  OAI21_X1 U10166 ( .B1(n8645), .B2(n8644), .A(n8643), .ZN(n8649) );
  NOR2_X1 U10167 ( .A1(n9956), .A2(n8646), .ZN(n8647) );
  AOI211_X1 U10168 ( .C1(n10029), .C2(n8649), .A(n8648), .B(n8647), .ZN(n8650)
         );
  OAI21_X1 U10169 ( .B1(n10033), .B2(n8651), .A(n8650), .ZN(n8652) );
  AOI21_X1 U10170 ( .B1(n8653), .B2(n10017), .A(n8652), .ZN(n8654) );
  OAI21_X1 U10171 ( .B1(n8655), .B2(n10024), .A(n8654), .ZN(P2_U3199) );
  NOR2_X1 U10172 ( .A1(n8660), .A2(n8812), .ZN(n8657) );
  MUX2_X1 U10173 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n5378), .S(n8668), .Z(n8663) );
  XNOR2_X1 U10174 ( .A(n8668), .B(n8853), .ZN(n8664) );
  OAI21_X1 U10175 ( .B1(n8661), .B2(n8660), .A(n8659), .ZN(n8666) );
  MUX2_X1 U10176 ( .A(n8664), .B(n8663), .S(n8662), .Z(n8665) );
  XNOR2_X1 U10177 ( .A(n8666), .B(n8665), .ZN(n8672) );
  OAI21_X1 U10178 ( .B1(n9956), .B2(n8668), .A(n8667), .ZN(n8669) );
  AOI21_X1 U10179 ( .B1(P2_ADDR_REG_19__SCAN_IN), .B2(n9946), .A(n8669), .ZN(
        n8670) );
  OAI21_X1 U10180 ( .B1(n8672), .B2(n8671), .A(n8670), .ZN(n8673) );
  AOI21_X1 U10181 ( .B1(n10050), .B2(n8862), .A(n8676), .ZN(n8680) );
  NAND2_X1 U10182 ( .A1(n8797), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n8677) );
  OAI211_X1 U10183 ( .C1(n8678), .C2(n8681), .A(n8680), .B(n8677), .ZN(
        P2_U3202) );
  NAND2_X1 U10184 ( .A1(n8797), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n8679) );
  OAI211_X1 U10185 ( .C1(n8866), .C2(n8681), .A(n8680), .B(n8679), .ZN(
        P2_U3203) );
  MUX2_X1 U10186 ( .A(n8682), .B(n8867), .S(n10050), .Z(n8685) );
  AOI22_X1 U10187 ( .A1(n8869), .A2(n8816), .B1(n8815), .B2(n8683), .ZN(n8684)
         );
  OAI211_X1 U10188 ( .C1(n8872), .C2(n8819), .A(n8685), .B(n8684), .ZN(
        P2_U3205) );
  XNOR2_X1 U10189 ( .A(n8686), .B(n8687), .ZN(n8878) );
  XOR2_X1 U10190 ( .A(n8688), .B(n8687), .Z(n8693) );
  MUX2_X1 U10191 ( .A(n8694), .B(n8873), .S(n10050), .Z(n8697) );
  AOI22_X1 U10192 ( .A1(n8875), .A2(n8816), .B1(n8815), .B2(n8695), .ZN(n8696)
         );
  OAI211_X1 U10193 ( .C1(n8878), .C2(n8819), .A(n8697), .B(n8696), .ZN(
        P2_U3206) );
  XNOR2_X1 U10194 ( .A(n8699), .B(n8698), .ZN(n8884) );
  XNOR2_X1 U10195 ( .A(n8700), .B(n8701), .ZN(n8704) );
  AOI222_X1 U10196 ( .A1(n5513), .A2(n8704), .B1(n8703), .B2(n8809), .C1(n8702), .C2(n8807), .ZN(n8879) );
  MUX2_X1 U10197 ( .A(n8705), .B(n8879), .S(n10050), .Z(n8708) );
  AOI22_X1 U10198 ( .A1(n8881), .A2(n8816), .B1(n8706), .B2(n8815), .ZN(n8707)
         );
  OAI211_X1 U10199 ( .C1(n8884), .C2(n8819), .A(n8708), .B(n8707), .ZN(
        P2_U3207) );
  NAND2_X1 U10200 ( .A1(n8709), .A2(n8721), .ZN(n8710) );
  NAND2_X1 U10201 ( .A1(n8711), .A2(n8710), .ZN(n8716) );
  NAND2_X1 U10202 ( .A1(n8712), .A2(n8809), .ZN(n8713) );
  OAI21_X1 U10203 ( .B1(n8714), .B2(n10043), .A(n8713), .ZN(n8715) );
  AOI21_X1 U10204 ( .B1(n8716), .B2(n5513), .A(n8715), .ZN(n8886) );
  AOI22_X1 U10205 ( .A1(n8887), .A2(n8718), .B1(n8815), .B2(n8717), .ZN(n8719)
         );
  AOI21_X1 U10206 ( .B1(n8886), .B2(n8719), .A(n8797), .ZN(n8724) );
  XNOR2_X1 U10207 ( .A(n8720), .B(n8721), .ZN(n8890) );
  OAI22_X1 U10208 ( .A1(n8890), .A2(n8819), .B1(n8722), .B2(n10050), .ZN(n8723) );
  OR2_X1 U10209 ( .A1(n8724), .A2(n8723), .ZN(P2_U3208) );
  NAND2_X1 U10210 ( .A1(n8726), .A2(n8725), .ZN(n8727) );
  XNOR2_X1 U10211 ( .A(n8727), .B(n8729), .ZN(n8894) );
  XOR2_X1 U10212 ( .A(n8729), .B(n8728), .Z(n8730) );
  OAI222_X1 U10213 ( .A1(n10041), .A2(n8732), .B1(n10043), .B2(n8731), .C1(
        n8792), .C2(n8730), .ZN(n8891) );
  INV_X1 U10214 ( .A(n8733), .ZN(n8734) );
  OAI22_X1 U10215 ( .A1(n8893), .A2(n10036), .B1(n8734), .B2(n10038), .ZN(
        n8735) );
  OAI21_X1 U10216 ( .B1(n8891), .B2(n8735), .A(n10050), .ZN(n8737) );
  NAND2_X1 U10217 ( .A1(n8797), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n8736) );
  OAI211_X1 U10218 ( .C1(n8894), .C2(n8819), .A(n8737), .B(n8736), .ZN(
        P2_U3209) );
  XOR2_X1 U10219 ( .A(n8739), .B(n8738), .Z(n8902) );
  XNOR2_X1 U10220 ( .A(n8740), .B(n8739), .ZN(n8742) );
  AOI222_X1 U10221 ( .A1(n5513), .A2(n8742), .B1(n8741), .B2(n8809), .C1(n8768), .C2(n8807), .ZN(n8897) );
  MUX2_X1 U10222 ( .A(n8743), .B(n8897), .S(n10050), .Z(n8746) );
  AOI22_X1 U10223 ( .A1(n8899), .A2(n8816), .B1(n8815), .B2(n8744), .ZN(n8745)
         );
  OAI211_X1 U10224 ( .C1(n8902), .C2(n8819), .A(n8746), .B(n8745), .ZN(
        P2_U3210) );
  XNOR2_X1 U10225 ( .A(n8747), .B(n8750), .ZN(n8908) );
  INV_X1 U10226 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n8756) );
  NAND3_X1 U10227 ( .A1(n8748), .A2(n8750), .A3(n8749), .ZN(n8751) );
  NAND2_X1 U10228 ( .A1(n8752), .A2(n8751), .ZN(n8755) );
  AOI222_X1 U10229 ( .A1(n5513), .A2(n8755), .B1(n8754), .B2(n8807), .C1(n8753), .C2(n8809), .ZN(n8903) );
  MUX2_X1 U10230 ( .A(n8756), .B(n8903), .S(n10050), .Z(n8759) );
  AOI22_X1 U10231 ( .A1(n8905), .A2(n8816), .B1(n8815), .B2(n8757), .ZN(n8758)
         );
  OAI211_X1 U10232 ( .C1(n8908), .C2(n8819), .A(n8759), .B(n8758), .ZN(
        P2_U3211) );
  NAND2_X1 U10233 ( .A1(n8761), .A2(n8760), .ZN(n8763) );
  XNOR2_X1 U10234 ( .A(n8763), .B(n8762), .ZN(n8914) );
  NAND3_X1 U10235 ( .A1(n8764), .A2(n4715), .A3(n8765), .ZN(n8766) );
  NAND2_X1 U10236 ( .A1(n8748), .A2(n8766), .ZN(n8769) );
  AOI222_X1 U10237 ( .A1(n5513), .A2(n8769), .B1(n8768), .B2(n8809), .C1(n8767), .C2(n8807), .ZN(n8909) );
  MUX2_X1 U10238 ( .A(n8770), .B(n8909), .S(n10050), .Z(n8773) );
  AOI22_X1 U10239 ( .A1(n8911), .A2(n8816), .B1(n8815), .B2(n8771), .ZN(n8772)
         );
  OAI211_X1 U10240 ( .C1(n8914), .C2(n8819), .A(n8773), .B(n8772), .ZN(
        P2_U3212) );
  XOR2_X1 U10241 ( .A(n8774), .B(n8775), .Z(n8920) );
  NAND2_X1 U10242 ( .A1(n8776), .A2(n8775), .ZN(n8777) );
  NAND2_X1 U10243 ( .A1(n8764), .A2(n8777), .ZN(n8781) );
  NAND2_X1 U10244 ( .A1(n8810), .A2(n8807), .ZN(n8778) );
  OAI21_X1 U10245 ( .B1(n8779), .B2(n10041), .A(n8778), .ZN(n8780) );
  AOI21_X1 U10246 ( .B1(n8781), .B2(n5513), .A(n8780), .ZN(n8916) );
  MUX2_X1 U10247 ( .A(n8916), .B(n8782), .S(n8797), .Z(n8786) );
  INV_X1 U10248 ( .A(n8783), .ZN(n8784) );
  AOI22_X1 U10249 ( .A1(n8917), .A2(n8816), .B1(n8815), .B2(n8784), .ZN(n8785)
         );
  OAI211_X1 U10250 ( .C1(n8920), .C2(n8819), .A(n8786), .B(n8785), .ZN(
        P2_U3213) );
  XNOR2_X1 U10251 ( .A(n8787), .B(n8788), .ZN(n8924) );
  XNOR2_X1 U10252 ( .A(n8790), .B(n8789), .ZN(n8791) );
  OAI222_X1 U10253 ( .A1(n10041), .A2(n8794), .B1(n10043), .B2(n8793), .C1(
        n8792), .C2(n8791), .ZN(n8851) );
  NOR2_X1 U10254 ( .A1(n10038), .A2(n8795), .ZN(n8796) );
  OAI21_X1 U10255 ( .B1(n8851), .B2(n8796), .A(n10050), .ZN(n8799) );
  AOI22_X1 U10256 ( .A1(n8852), .A2(n8816), .B1(P2_REG2_REG_19__SCAN_IN), .B2(
        n8797), .ZN(n8798) );
  OAI211_X1 U10257 ( .C1(n8924), .C2(n8819), .A(n8799), .B(n8798), .ZN(
        P2_U3214) );
  NAND2_X1 U10258 ( .A1(n8801), .A2(n8800), .ZN(n8805) );
  NAND2_X1 U10259 ( .A1(n8803), .A2(n8802), .ZN(n8804) );
  XOR2_X1 U10260 ( .A(n8805), .B(n8804), .Z(n8932) );
  XOR2_X1 U10261 ( .A(n8806), .B(n8805), .Z(n8811) );
  AOI222_X1 U10262 ( .A1(n5513), .A2(n8811), .B1(n8810), .B2(n8809), .C1(n8808), .C2(n8807), .ZN(n8925) );
  MUX2_X1 U10263 ( .A(n8812), .B(n8925), .S(n10050), .Z(n8818) );
  INV_X1 U10264 ( .A(n8813), .ZN(n8814) );
  AOI22_X1 U10265 ( .A1(n8928), .A2(n8816), .B1(n8815), .B2(n8814), .ZN(n8817)
         );
  OAI211_X1 U10266 ( .C1(n8932), .C2(n8819), .A(n8818), .B(n8817), .ZN(
        P2_U3215) );
  INV_X1 U10267 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n8821) );
  NAND2_X1 U10268 ( .A1(n8861), .A2(n8856), .ZN(n8820) );
  NAND2_X1 U10269 ( .A1(n8862), .A2(n10135), .ZN(n8823) );
  OAI211_X1 U10270 ( .C1(n10135), .C2(n8821), .A(n8820), .B(n8823), .ZN(
        P2_U3490) );
  INV_X1 U10271 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n8825) );
  NAND2_X1 U10272 ( .A1(n8822), .A2(n8856), .ZN(n8824) );
  OAI211_X1 U10273 ( .C1(n10135), .C2(n8825), .A(n8824), .B(n8823), .ZN(
        P2_U3489) );
  NAND2_X1 U10274 ( .A1(n8873), .A2(n10135), .ZN(n8827) );
  OR2_X1 U10275 ( .A1(n10135), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n8826) );
  NAND2_X1 U10276 ( .A1(n8875), .A2(n8856), .ZN(n8828) );
  OAI211_X1 U10277 ( .C1(n8878), .C2(n8859), .A(n8829), .B(n8828), .ZN(
        P2_U3486) );
  INV_X1 U10278 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n8830) );
  MUX2_X1 U10279 ( .A(n8830), .B(n8879), .S(n10135), .Z(n8832) );
  NAND2_X1 U10280 ( .A1(n8881), .A2(n8856), .ZN(n8831) );
  OAI211_X1 U10281 ( .C1(n8884), .C2(n8859), .A(n8832), .B(n8831), .ZN(
        P2_U3485) );
  INV_X1 U10282 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n8833) );
  MUX2_X1 U10283 ( .A(n8886), .B(n8833), .S(n5719), .Z(n8835) );
  NAND2_X1 U10284 ( .A1(n8887), .A2(n8856), .ZN(n8834) );
  OAI211_X1 U10285 ( .C1(n8890), .C2(n8859), .A(n8835), .B(n8834), .ZN(
        P2_U3484) );
  MUX2_X1 U10286 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n8891), .S(n10135), .Z(
        n8838) );
  OAI22_X1 U10287 ( .A1(n8894), .A2(n8859), .B1(n8893), .B2(n8836), .ZN(n8837)
         );
  OR2_X1 U10288 ( .A1(n8838), .A2(n8837), .ZN(P2_U3483) );
  INV_X1 U10289 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n8839) );
  MUX2_X1 U10290 ( .A(n8839), .B(n8897), .S(n10135), .Z(n8841) );
  NAND2_X1 U10291 ( .A1(n8899), .A2(n8856), .ZN(n8840) );
  OAI211_X1 U10292 ( .C1(n8902), .C2(n8859), .A(n8841), .B(n8840), .ZN(
        P2_U3482) );
  INV_X1 U10293 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n8842) );
  MUX2_X1 U10294 ( .A(n8842), .B(n8903), .S(n10135), .Z(n8844) );
  NAND2_X1 U10295 ( .A1(n8905), .A2(n8856), .ZN(n8843) );
  OAI211_X1 U10296 ( .C1(n8908), .C2(n8859), .A(n8844), .B(n8843), .ZN(
        P2_U3481) );
  MUX2_X1 U10297 ( .A(n8845), .B(n8909), .S(n10135), .Z(n8847) );
  NAND2_X1 U10298 ( .A1(n8911), .A2(n8856), .ZN(n8846) );
  OAI211_X1 U10299 ( .C1(n8859), .C2(n8914), .A(n8847), .B(n8846), .ZN(
        P2_U3480) );
  INV_X1 U10300 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n8848) );
  MUX2_X1 U10301 ( .A(n8848), .B(n8916), .S(n10135), .Z(n8850) );
  NAND2_X1 U10302 ( .A1(n8917), .A2(n8856), .ZN(n8849) );
  OAI211_X1 U10303 ( .C1(n8859), .C2(n8920), .A(n8850), .B(n8849), .ZN(
        P2_U3479) );
  AOI21_X1 U10304 ( .B1(n10112), .B2(n8852), .A(n8851), .ZN(n8921) );
  MUX2_X1 U10305 ( .A(n8853), .B(n8921), .S(n10135), .Z(n8854) );
  OAI21_X1 U10306 ( .B1(n8859), .B2(n8924), .A(n8854), .ZN(P2_U3478) );
  MUX2_X1 U10307 ( .A(n8855), .B(n8925), .S(n10135), .Z(n8858) );
  NAND2_X1 U10308 ( .A1(n8928), .A2(n8856), .ZN(n8857) );
  OAI211_X1 U10309 ( .C1(n8932), .C2(n8859), .A(n8858), .B(n8857), .ZN(
        P2_U3477) );
  MUX2_X1 U10310 ( .A(P2_REG1_REG_0__SCAN_IN), .B(n8860), .S(n10135), .Z(
        P2_U3459) );
  NAND2_X1 U10311 ( .A1(n8861), .A2(n8927), .ZN(n8863) );
  NAND2_X1 U10312 ( .A1(n10118), .A2(n8862), .ZN(n8864) );
  OAI211_X1 U10313 ( .C1(n8104), .C2(n10118), .A(n8863), .B(n8864), .ZN(
        P2_U3458) );
  NAND2_X1 U10314 ( .A1(n10120), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n8865) );
  OAI211_X1 U10315 ( .C1(n8866), .C2(n8892), .A(n8865), .B(n8864), .ZN(
        P2_U3457) );
  INV_X1 U10316 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n8868) );
  MUX2_X1 U10317 ( .A(n8868), .B(n8867), .S(n10118), .Z(n8871) );
  NAND2_X1 U10318 ( .A1(n8869), .A2(n8927), .ZN(n8870) );
  OAI211_X1 U10319 ( .C1(n8872), .C2(n8931), .A(n8871), .B(n8870), .ZN(
        P2_U3455) );
  INV_X1 U10320 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n8874) );
  MUX2_X1 U10321 ( .A(n8874), .B(n8873), .S(n10118), .Z(n8877) );
  NAND2_X1 U10322 ( .A1(n8875), .A2(n8927), .ZN(n8876) );
  OAI211_X1 U10323 ( .C1(n8878), .C2(n8931), .A(n8877), .B(n8876), .ZN(
        P2_U3454) );
  INV_X1 U10324 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n8880) );
  MUX2_X1 U10325 ( .A(n8880), .B(n8879), .S(n10118), .Z(n8883) );
  NAND2_X1 U10326 ( .A1(n8881), .A2(n8927), .ZN(n8882) );
  OAI211_X1 U10327 ( .C1(n8884), .C2(n8931), .A(n8883), .B(n8882), .ZN(
        P2_U3453) );
  INV_X1 U10328 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n8885) );
  MUX2_X1 U10329 ( .A(n8886), .B(n8885), .S(n10120), .Z(n8889) );
  NAND2_X1 U10330 ( .A1(n8887), .A2(n8927), .ZN(n8888) );
  OAI211_X1 U10331 ( .C1(n8890), .C2(n8931), .A(n8889), .B(n8888), .ZN(
        P2_U3452) );
  MUX2_X1 U10332 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n8891), .S(n10118), .Z(
        n8896) );
  OAI22_X1 U10333 ( .A1(n8894), .A2(n8931), .B1(n8893), .B2(n8892), .ZN(n8895)
         );
  OR2_X1 U10334 ( .A1(n8896), .A2(n8895), .ZN(P2_U3451) );
  INV_X1 U10335 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n8898) );
  MUX2_X1 U10336 ( .A(n8898), .B(n8897), .S(n10118), .Z(n8901) );
  NAND2_X1 U10337 ( .A1(n8899), .A2(n8927), .ZN(n8900) );
  OAI211_X1 U10338 ( .C1(n8902), .C2(n8931), .A(n8901), .B(n8900), .ZN(
        P2_U3450) );
  INV_X1 U10339 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n8904) );
  MUX2_X1 U10340 ( .A(n8904), .B(n8903), .S(n10118), .Z(n8907) );
  NAND2_X1 U10341 ( .A1(n8905), .A2(n8927), .ZN(n8906) );
  OAI211_X1 U10342 ( .C1(n8908), .C2(n8931), .A(n8907), .B(n8906), .ZN(
        P2_U3449) );
  MUX2_X1 U10343 ( .A(n8910), .B(n8909), .S(n10118), .Z(n8913) );
  NAND2_X1 U10344 ( .A1(n8911), .A2(n8927), .ZN(n8912) );
  OAI211_X1 U10345 ( .C1(n8914), .C2(n8931), .A(n8913), .B(n8912), .ZN(
        P2_U3448) );
  MUX2_X1 U10346 ( .A(n8916), .B(n8915), .S(n10120), .Z(n8919) );
  NAND2_X1 U10347 ( .A1(n8917), .A2(n8927), .ZN(n8918) );
  OAI211_X1 U10348 ( .C1(n8920), .C2(n8931), .A(n8919), .B(n8918), .ZN(
        P2_U3447) );
  INV_X1 U10349 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n8922) );
  MUX2_X1 U10350 ( .A(n8922), .B(n8921), .S(n10118), .Z(n8923) );
  OAI21_X1 U10351 ( .B1(n8924), .B2(n8931), .A(n8923), .ZN(P2_U3446) );
  INV_X1 U10352 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n8926) );
  MUX2_X1 U10353 ( .A(n8926), .B(n8925), .S(n10118), .Z(n8930) );
  NAND2_X1 U10354 ( .A1(n8928), .A2(n8927), .ZN(n8929) );
  OAI211_X1 U10355 ( .C1(n8932), .C2(n8931), .A(n8930), .B(n8929), .ZN(
        P2_U3444) );
  MUX2_X1 U10356 ( .A(n8933), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  INV_X1 U10357 ( .A(n9401), .ZN(n9257) );
  NAND2_X1 U10358 ( .A1(n8935), .A2(n8934), .ZN(n8938) );
  OAI21_X1 U10359 ( .B1(n8938), .B2(n8937), .A(n8936), .ZN(n8940) );
  AOI21_X1 U10360 ( .B1(n8940), .B2(n8939), .A(n9036), .ZN(n8941) );
  INV_X1 U10361 ( .A(n8941), .ZN(n8945) );
  OAI22_X1 U10362 ( .A1(n9195), .A2(n9017), .B1(n9199), .B2(n9162), .ZN(n9260)
         );
  INV_X1 U10363 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n8942) );
  OAI22_X1 U10364 ( .A1(n9021), .A2(n9254), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8942), .ZN(n8943) );
  AOI21_X1 U10365 ( .B1(n9260), .B2(n9018), .A(n8943), .ZN(n8944) );
  OAI211_X1 U10366 ( .C1(n9257), .C2(n9061), .A(n8945), .B(n8944), .ZN(
        P1_U3214) );
  XNOR2_X1 U10367 ( .A(n8946), .B(n8947), .ZN(n9039) );
  NAND2_X1 U10368 ( .A1(n9039), .A2(n9040), .ZN(n9038) );
  NAND2_X1 U10369 ( .A1(n4544), .A2(n8947), .ZN(n8950) );
  AND2_X1 U10370 ( .A1(n9038), .A2(n8950), .ZN(n8952) );
  XNOR2_X1 U10371 ( .A(n8949), .B(n8948), .ZN(n8951) );
  NAND3_X1 U10372 ( .A1(n9038), .A2(n8951), .A3(n8950), .ZN(n9011) );
  OAI211_X1 U10373 ( .C1(n8952), .C2(n8951), .A(n9050), .B(n9011), .ZN(n8958)
         );
  OR2_X1 U10374 ( .A1(n9177), .A2(n9162), .ZN(n8954) );
  NAND2_X1 U10375 ( .A1(n9171), .A2(n9225), .ZN(n8953) );
  NAND2_X1 U10376 ( .A1(n8954), .A2(n8953), .ZN(n9373) );
  NOR2_X1 U10377 ( .A1(n8955), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9153) );
  NOR2_X1 U10378 ( .A1(n9021), .A2(n9367), .ZN(n8956) );
  AOI211_X1 U10379 ( .C1(n9018), .C2(n9373), .A(n9153), .B(n8956), .ZN(n8957)
         );
  OAI211_X1 U10380 ( .C1(n9370), .C2(n9061), .A(n8958), .B(n8957), .ZN(
        P1_U3219) );
  AND2_X1 U10381 ( .A1(n8959), .A2(n9012), .ZN(n8961) );
  OAI21_X1 U10382 ( .B1(n8962), .B2(n8961), .A(n8960), .ZN(n8963) );
  NAND2_X1 U10383 ( .A1(n8963), .A2(n9050), .ZN(n8969) );
  OR2_X1 U10384 ( .A1(n9185), .A2(n9162), .ZN(n8965) );
  OR2_X1 U10385 ( .A1(n9177), .A2(n9017), .ZN(n8964) );
  AND2_X1 U10386 ( .A1(n8965), .A2(n8964), .ZN(n9341) );
  INV_X1 U10387 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n8966) );
  OAI22_X1 U10388 ( .A1(n9341), .A2(n9056), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8966), .ZN(n8967) );
  AOI21_X1 U10389 ( .B1(n9344), .B2(n9058), .A(n8967), .ZN(n8968) );
  OAI211_X1 U10390 ( .C1(n9337), .C2(n9061), .A(n8969), .B(n8968), .ZN(
        P1_U3223) );
  NAND2_X1 U10391 ( .A1(n9002), .A2(n9003), .ZN(n9001) );
  NAND2_X1 U10392 ( .A1(n9001), .A2(n8970), .ZN(n8973) );
  OAI21_X1 U10393 ( .B1(n8974), .B2(n8973), .A(n8972), .ZN(n8975) );
  NAND2_X1 U10394 ( .A1(n8975), .A2(n9050), .ZN(n8980) );
  OAI22_X1 U10395 ( .A1(n9195), .A2(n9162), .B1(n9189), .B2(n9017), .ZN(n9285)
         );
  INV_X1 U10396 ( .A(n9280), .ZN(n8977) );
  OAI22_X1 U10397 ( .A1(n8977), .A2(n9021), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8976), .ZN(n8978) );
  AOI21_X1 U10398 ( .B1(n9285), .B2(n9018), .A(n8978), .ZN(n8979) );
  OAI211_X1 U10399 ( .C1(n9282), .C2(n9061), .A(n8980), .B(n8979), .ZN(
        P1_U3225) );
  XOR2_X1 U10400 ( .A(n8982), .B(n8981), .Z(n8988) );
  NAND2_X1 U10401 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9106) );
  NAND2_X1 U10402 ( .A1(n9018), .A2(n8983), .ZN(n8984) );
  OAI211_X1 U10403 ( .C1(n9021), .C2(n8985), .A(n9106), .B(n8984), .ZN(n8986)
         );
  AOI21_X1 U10404 ( .B1(n9454), .B2(n9023), .A(n8986), .ZN(n8987) );
  OAI21_X1 U10405 ( .B1(n8988), .B2(n9036), .A(n8987), .ZN(P1_U3226) );
  XNOR2_X1 U10406 ( .A(n8990), .B(n8989), .ZN(n8991) );
  XNOR2_X1 U10407 ( .A(n4421), .B(n8991), .ZN(n9000) );
  INV_X1 U10408 ( .A(n8992), .ZN(n8993) );
  NOR3_X1 U10409 ( .A1(n9021), .A2(P1_REG3_REG_17__SCAN_IN), .A3(n8993), .ZN(
        n8998) );
  OAI21_X1 U10410 ( .B1(n8993), .B2(P1_U3086), .A(P1_REG3_REG_17__SCAN_IN), 
        .ZN(n8995) );
  OAI22_X1 U10411 ( .A1(n8996), .A2(n8995), .B1(n9056), .B2(n8994), .ZN(n8997)
         );
  AOI211_X1 U10412 ( .C1(n9449), .C2(n9023), .A(n8998), .B(n8997), .ZN(n8999)
         );
  OAI21_X1 U10413 ( .B1(n9000), .B2(n9036), .A(n8999), .ZN(P1_U3228) );
  OAI21_X1 U10414 ( .B1(n9003), .B2(n9002), .A(n9001), .ZN(n9004) );
  NAND2_X1 U10415 ( .A1(n9004), .A2(n9050), .ZN(n9009) );
  OAI22_X1 U10416 ( .A1(n9193), .A2(n9162), .B1(n9188), .B2(n9017), .ZN(n9298)
         );
  INV_X1 U10417 ( .A(n9294), .ZN(n9006) );
  INV_X1 U10418 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n9005) );
  OAI22_X1 U10419 ( .A1(n9006), .A2(n9021), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9005), .ZN(n9007) );
  AOI21_X1 U10420 ( .B1(n9298), .B2(n9018), .A(n9007), .ZN(n9008) );
  OAI211_X1 U10421 ( .C1(n9154), .C2(n9061), .A(n9009), .B(n9008), .ZN(
        P1_U3229) );
  NAND2_X1 U10422 ( .A1(n9011), .A2(n9010), .ZN(n9016) );
  INV_X1 U10423 ( .A(n9012), .ZN(n9013) );
  NOR2_X1 U10424 ( .A1(n9014), .A2(n9013), .ZN(n9015) );
  XNOR2_X1 U10425 ( .A(n9016), .B(n9015), .ZN(n9025) );
  INV_X1 U10426 ( .A(n9352), .ZN(n9020) );
  OAI22_X1 U10427 ( .A1(n9181), .A2(n9162), .B1(n9176), .B2(n9017), .ZN(n9357)
         );
  AOI22_X1 U10428 ( .A1(n9357), .A2(n9018), .B1(P1_REG3_REG_20__SCAN_IN), .B2(
        P1_U3086), .ZN(n9019) );
  OAI21_X1 U10429 ( .B1(n9021), .B2(n9020), .A(n9019), .ZN(n9022) );
  AOI21_X1 U10430 ( .B1(n9435), .B2(n9023), .A(n9022), .ZN(n9024) );
  OAI21_X1 U10431 ( .B1(n9025), .B2(n9036), .A(n9024), .ZN(P1_U3233) );
  NAND2_X1 U10432 ( .A1(n9027), .A2(n9026), .ZN(n9028) );
  XOR2_X1 U10433 ( .A(n9029), .B(n9028), .Z(n9037) );
  OR2_X1 U10434 ( .A1(n9188), .A2(n9162), .ZN(n9031) );
  NAND2_X1 U10435 ( .A1(n9170), .A2(n9225), .ZN(n9030) );
  AND2_X1 U10436 ( .A1(n9031), .A2(n9030), .ZN(n9327) );
  OAI22_X1 U10437 ( .A1(n9327), .A2(n9056), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9032), .ZN(n9034) );
  NOR2_X1 U10438 ( .A1(n9323), .A2(n9061), .ZN(n9033) );
  AOI211_X1 U10439 ( .C1(n9321), .C2(n9058), .A(n9034), .B(n9033), .ZN(n9035)
         );
  OAI21_X1 U10440 ( .B1(n9037), .B2(n9036), .A(n9035), .ZN(P1_U3235) );
  OAI21_X1 U10441 ( .B1(n9040), .B2(n9039), .A(n9038), .ZN(n9041) );
  NAND2_X1 U10442 ( .A1(n9041), .A2(n9050), .ZN(n9046) );
  NAND2_X1 U10443 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9726) );
  OAI21_X1 U10444 ( .B1(n9056), .B2(n9042), .A(n9726), .ZN(n9043) );
  AOI21_X1 U10445 ( .B1(n9058), .B2(n9044), .A(n9043), .ZN(n9045) );
  OAI211_X1 U10446 ( .C1(n9173), .C2(n9061), .A(n9046), .B(n9045), .ZN(
        P1_U3238) );
  OAI21_X1 U10447 ( .B1(n9049), .B2(n9048), .A(n9047), .ZN(n9051) );
  NAND2_X1 U10448 ( .A1(n9051), .A2(n9050), .ZN(n9060) );
  NAND2_X1 U10449 ( .A1(n9067), .A2(n9225), .ZN(n9054) );
  NAND2_X1 U10450 ( .A1(n9065), .A2(n9052), .ZN(n9053) );
  AND2_X1 U10451 ( .A1(n9054), .A2(n9053), .ZN(n9551) );
  OAI22_X1 U10452 ( .A1(n9056), .A2(n9551), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9055), .ZN(n9057) );
  AOI21_X1 U10453 ( .B1(n9058), .B2(n9555), .A(n9057), .ZN(n9059) );
  OAI211_X1 U10454 ( .C1(n7446), .C2(n9061), .A(n9060), .B(n9059), .ZN(
        P1_U3241) );
  MUX2_X1 U10455 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9223), .S(P1_U3973), .Z(
        P1_U3584) );
  MUX2_X1 U10456 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n9062), .S(P1_U3973), .Z(
        P1_U3583) );
  MUX2_X1 U10457 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9226), .S(P1_U3973), .Z(
        P1_U3582) );
  MUX2_X1 U10458 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9063), .S(P1_U3973), .Z(
        P1_U3581) );
  INV_X1 U10459 ( .A(n9195), .ZN(n9196) );
  MUX2_X1 U10460 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9196), .S(P1_U3973), .Z(
        P1_U3580) );
  MUX2_X1 U10461 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9192), .S(P1_U3973), .Z(
        P1_U3579) );
  MUX2_X1 U10462 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9190), .S(P1_U3973), .Z(
        P1_U3578) );
  INV_X1 U10463 ( .A(n9188), .ZN(n9187) );
  MUX2_X1 U10464 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9187), .S(P1_U3973), .Z(
        P1_U3577) );
  MUX2_X1 U10465 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9184), .S(P1_U3973), .Z(
        P1_U3576) );
  MUX2_X1 U10466 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9170), .S(P1_U3973), .Z(
        P1_U3575) );
  MUX2_X1 U10467 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9178), .S(P1_U3973), .Z(
        P1_U3574) );
  MUX2_X1 U10468 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9175), .S(P1_U3973), .Z(
        P1_U3573) );
  MUX2_X1 U10469 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9171), .S(P1_U3973), .Z(
        P1_U3572) );
  MUX2_X1 U10470 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9064), .S(P1_U3973), .Z(
        P1_U3571) );
  MUX2_X1 U10471 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9065), .S(P1_U3973), .Z(
        P1_U3570) );
  MUX2_X1 U10472 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n9066), .S(P1_U3973), .Z(
        P1_U3569) );
  MUX2_X1 U10473 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n9067), .S(P1_U3973), .Z(
        P1_U3568) );
  MUX2_X1 U10474 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9068), .S(P1_U3973), .Z(
        P1_U3567) );
  MUX2_X1 U10475 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n9069), .S(P1_U3973), .Z(
        P1_U3566) );
  INV_X1 U10476 ( .A(n9070), .ZN(n9071) );
  MUX2_X1 U10477 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n9071), .S(P1_U3973), .Z(
        P1_U3565) );
  MUX2_X1 U10478 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n9072), .S(P1_U3973), .Z(
        P1_U3564) );
  MUX2_X1 U10479 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n9073), .S(P1_U3973), .Z(
        P1_U3563) );
  MUX2_X1 U10480 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n9074), .S(P1_U3973), .Z(
        P1_U3562) );
  MUX2_X1 U10481 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n9075), .S(P1_U3973), .Z(
        P1_U3561) );
  MUX2_X1 U10482 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n9076), .S(P1_U3973), .Z(
        P1_U3560) );
  MUX2_X1 U10483 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n9077), .S(P1_U3973), .Z(
        P1_U3559) );
  MUX2_X1 U10484 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n9078), .S(P1_U3973), .Z(
        P1_U3558) );
  MUX2_X1 U10485 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n9079), .S(P1_U3973), .Z(
        P1_U3557) );
  MUX2_X1 U10486 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n9080), .S(P1_U3973), .Z(
        P1_U3556) );
  MUX2_X1 U10487 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n6616), .S(P1_U3973), .Z(
        P1_U3555) );
  MUX2_X1 U10488 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n9081), .S(P1_U3973), .Z(
        P1_U3554) );
  OAI21_X1 U10489 ( .B1(n9084), .B2(n9083), .A(n9082), .ZN(n9085) );
  NAND2_X1 U10490 ( .A1(n9085), .A2(n9718), .ZN(n9095) );
  AOI21_X1 U10491 ( .B1(n9609), .B2(P1_ADDR_REG_9__SCAN_IN), .A(n9086), .ZN(
        n9094) );
  OAI21_X1 U10492 ( .B1(n9089), .B2(n9088), .A(n9087), .ZN(n9090) );
  NAND2_X1 U10493 ( .A1(n9090), .A2(n9713), .ZN(n9093) );
  INV_X1 U10494 ( .A(n9724), .ZN(n9709) );
  NAND2_X1 U10495 ( .A1(n9709), .A2(n9091), .ZN(n9092) );
  NAND4_X1 U10496 ( .A1(n9095), .A2(n9094), .A3(n9093), .A4(n9092), .ZN(
        P1_U3252) );
  AOI22_X1 U10497 ( .A1(n9128), .A2(P1_REG1_REG_16__SCAN_IN), .B1(n7433), .B2(
        n9107), .ZN(n9104) );
  MUX2_X1 U10498 ( .A(n9096), .B(P1_REG1_REG_13__SCAN_IN), .S(n9680), .Z(n9673) );
  OAI21_X1 U10499 ( .B1(P1_REG1_REG_12__SCAN_IN), .B2(n9098), .A(n9097), .ZN(
        n9674) );
  NOR2_X1 U10500 ( .A1(n9673), .A2(n9674), .ZN(n9672) );
  AOI21_X1 U10501 ( .B1(n9680), .B2(P1_REG1_REG_13__SCAN_IN), .A(n9672), .ZN(
        n9686) );
  INV_X1 U10502 ( .A(n9113), .ZN(n9694) );
  NAND2_X1 U10503 ( .A1(n9694), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n9100) );
  NAND2_X1 U10504 ( .A1(n9113), .A2(n7260), .ZN(n9099) );
  AND2_X1 U10505 ( .A1(n9100), .A2(n9099), .ZN(n9685) );
  NOR2_X1 U10506 ( .A1(n9686), .A2(n9685), .ZN(n9684) );
  NOR2_X1 U10507 ( .A1(n9101), .A2(n9115), .ZN(n9102) );
  NAND2_X1 U10508 ( .A1(n9104), .A2(n9103), .ZN(n9125) );
  OAI21_X1 U10509 ( .B1(n9104), .B2(n9103), .A(n9125), .ZN(n9122) );
  NAND2_X1 U10510 ( .A1(n9609), .A2(P1_ADDR_REG_16__SCAN_IN), .ZN(n9105) );
  OAI211_X1 U10511 ( .C1(n9724), .C2(n9107), .A(n9106), .B(n9105), .ZN(n9121)
         );
  AOI22_X1 U10512 ( .A1(n9680), .A2(n7161), .B1(P1_REG2_REG_13__SCAN_IN), .B2(
        n9108), .ZN(n9676) );
  INV_X1 U10513 ( .A(n9109), .ZN(n9110) );
  NAND2_X1 U10514 ( .A1(n9113), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n9112) );
  OAI21_X1 U10515 ( .B1(n9113), .B2(P1_REG2_REG_14__SCAN_IN), .A(n9112), .ZN(
        n9690) );
  NOR2_X1 U10516 ( .A1(n9689), .A2(n9690), .ZN(n9688) );
  NOR2_X1 U10517 ( .A1(n9114), .A2(n9115), .ZN(n9116) );
  INV_X1 U10518 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n9704) );
  NAND2_X1 U10519 ( .A1(n9128), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n9117) );
  OAI21_X1 U10520 ( .B1(n9128), .B2(P1_REG2_REG_16__SCAN_IN), .A(n9117), .ZN(
        n9118) );
  NOR2_X1 U10521 ( .A1(n9119), .A2(n9118), .ZN(n9127) );
  AOI211_X1 U10522 ( .C1(n9119), .C2(n9118), .A(n9127), .B(n9702), .ZN(n9120)
         );
  AOI211_X1 U10523 ( .C1(n9713), .C2(n9122), .A(n9121), .B(n9120), .ZN(n9123)
         );
  INV_X1 U10524 ( .A(n9123), .ZN(P1_U3259) );
  XNOR2_X1 U10525 ( .A(n9140), .B(n9124), .ZN(n9135) );
  OAI21_X1 U10526 ( .B1(n9128), .B2(P1_REG1_REG_16__SCAN_IN), .A(n9125), .ZN(
        n9136) );
  XOR2_X1 U10527 ( .A(n9135), .B(n9136), .Z(n9134) );
  XNOR2_X1 U10528 ( .A(n9140), .B(n9126), .ZN(n9143) );
  XNOR2_X1 U10529 ( .A(n9143), .B(n9142), .ZN(n9132) );
  AOI22_X1 U10530 ( .A1(n9609), .A2(P1_ADDR_REG_17__SCAN_IN), .B1(
        P1_REG3_REG_17__SCAN_IN), .B2(P1_U3086), .ZN(n9129) );
  OAI21_X1 U10531 ( .B1(n9130), .B2(n9724), .A(n9129), .ZN(n9131) );
  AOI21_X1 U10532 ( .B1(n9718), .B2(n9132), .A(n9131), .ZN(n9133) );
  OAI21_X1 U10533 ( .B1(n9134), .B2(n9699), .A(n9133), .ZN(P1_U3260) );
  NAND2_X1 U10534 ( .A1(n9144), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n9138) );
  OR2_X1 U10535 ( .A1(n9144), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n9137) );
  AND2_X1 U10536 ( .A1(n9138), .A2(n9137), .ZN(n9715) );
  INV_X1 U10537 ( .A(n9150), .ZN(n9148) );
  NOR2_X1 U10538 ( .A1(n9140), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n9141) );
  AOI21_X1 U10539 ( .B1(n9143), .B2(n9142), .A(n9141), .ZN(n9719) );
  NAND2_X1 U10540 ( .A1(n9144), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9146) );
  OR2_X1 U10541 ( .A1(n9144), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9145) );
  AND2_X1 U10542 ( .A1(n9146), .A2(n9145), .ZN(n9720) );
  NAND2_X1 U10543 ( .A1(n9719), .A2(n9720), .ZN(n9717) );
  NAND2_X1 U10544 ( .A1(n9717), .A2(n9146), .ZN(n9147) );
  XNOR2_X1 U10545 ( .A(n9147), .B(P1_REG2_REG_19__SCAN_IN), .ZN(n9149) );
  INV_X1 U10546 ( .A(n9390), .ZN(n9155) );
  NOR2_X1 U10547 ( .A1(n9156), .A2(n9231), .ZN(n9158) );
  XNOR2_X1 U10548 ( .A(n9158), .B(n9157), .ZN(n9159) );
  NOR2_X1 U10549 ( .A1(n6484), .A2(n9160), .ZN(n9161) );
  NOR2_X1 U10550 ( .A1(n9162), .A2(n9161), .ZN(n9224) );
  NAND2_X1 U10551 ( .A1(n9163), .A2(n9224), .ZN(n9385) );
  NOR2_X1 U10552 ( .A1(n9836), .A2(n9385), .ZN(n9168) );
  NOR2_X1 U10553 ( .A1(n9380), .A2(n9825), .ZN(n9164) );
  AOI211_X1 U10554 ( .C1(n9836), .C2(P1_REG2_REG_31__SCAN_IN), .A(n9168), .B(
        n9164), .ZN(n9165) );
  OAI21_X1 U10555 ( .B1(n9379), .B2(n9248), .A(n9165), .ZN(P1_U3263) );
  XNOR2_X1 U10556 ( .A(n9231), .B(n9387), .ZN(n9166) );
  NAND2_X1 U10557 ( .A1(n9166), .A2(n9829), .ZN(n9386) );
  NOR2_X1 U10558 ( .A1(n9387), .A2(n9825), .ZN(n9167) );
  AOI211_X1 U10559 ( .C1(n9836), .C2(P1_REG2_REG_30__SCAN_IN), .A(n9168), .B(
        n9167), .ZN(n9169) );
  OAI21_X1 U10560 ( .B1(n9248), .B2(n9386), .A(n9169), .ZN(P1_U3264) );
  OR2_X1 U10561 ( .A1(n8183), .A2(n9170), .ZN(n9183) );
  NAND2_X1 U10562 ( .A1(n9354), .A2(n9177), .ZN(n9180) );
  NAND2_X1 U10563 ( .A1(n9333), .A2(n4869), .ZN(n9182) );
  NAND2_X1 U10564 ( .A1(n9183), .A2(n9182), .ZN(n9318) );
  NOR2_X1 U10565 ( .A1(n9426), .A2(n9184), .ZN(n9186) );
  NOR2_X1 U10566 ( .A1(n9154), .A2(n9189), .ZN(n9191) );
  NOR2_X1 U10567 ( .A1(n9411), .A2(n9192), .ZN(n9194) );
  OAI22_X1 U10568 ( .A1(n9278), .A2(n9194), .B1(n9282), .B2(n9193), .ZN(n9266)
         );
  NOR2_X1 U10569 ( .A1(n4637), .A2(n9195), .ZN(n9197) );
  XNOR2_X1 U10570 ( .A(n9201), .B(n9221), .ZN(n9388) );
  NAND2_X1 U10571 ( .A1(n9388), .A2(n9809), .ZN(n9236) );
  NAND2_X1 U10572 ( .A1(n9836), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n9202) );
  OAI21_X1 U10573 ( .B1(n9799), .B2(n9203), .A(n9202), .ZN(n9204) );
  AOI21_X1 U10574 ( .B1(n9390), .B2(n9753), .A(n9204), .ZN(n9235) );
  NAND2_X1 U10575 ( .A1(n9339), .A2(n9340), .ZN(n9338) );
  NAND2_X1 U10576 ( .A1(n9338), .A2(n9209), .ZN(n9325) );
  NAND2_X1 U10577 ( .A1(n9325), .A2(n9326), .ZN(n9324) );
  NAND2_X1 U10578 ( .A1(n9324), .A2(n9210), .ZN(n9310) );
  INV_X1 U10579 ( .A(n9304), .ZN(n9311) );
  INV_X1 U10580 ( .A(n9213), .ZN(n9214) );
  NAND2_X1 U10581 ( .A1(n9284), .A2(n4352), .ZN(n9283) );
  NAND2_X1 U10582 ( .A1(n9283), .A2(n9215), .ZN(n9272) );
  XNOR2_X1 U10583 ( .A(n9222), .B(n9221), .ZN(n9229) );
  OR2_X1 U10584 ( .A1(n9391), .A2(n9836), .ZN(n9234) );
  AOI21_X1 U10585 ( .B1(n9390), .B2(n9241), .A(n9775), .ZN(n9232) );
  NAND2_X1 U10586 ( .A1(n9389), .A2(n9832), .ZN(n9233) );
  NAND4_X1 U10587 ( .A1(n9236), .A2(n9235), .A3(n9234), .A4(n9233), .ZN(
        P1_U3356) );
  XNOR2_X1 U10588 ( .A(n9237), .B(n9242), .ZN(n9239) );
  NAND2_X1 U10589 ( .A1(n9395), .A2(n9252), .ZN(n9240) );
  NAND3_X1 U10590 ( .A1(n9241), .A2(n9829), .A3(n9240), .ZN(n9397) );
  OR2_X1 U10591 ( .A1(n4407), .A2(n9242), .ZN(n9394) );
  NAND3_X1 U10592 ( .A1(n9394), .A2(n9393), .A3(n9809), .ZN(n9247) );
  NAND2_X1 U10593 ( .A1(n9836), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n9243) );
  OAI21_X1 U10594 ( .B1(n9799), .B2(n9244), .A(n9243), .ZN(n9245) );
  AOI21_X1 U10595 ( .B1(n9395), .B2(n9753), .A(n9245), .ZN(n9246) );
  OAI211_X1 U10596 ( .C1(n9397), .C2(n9248), .A(n9247), .B(n9246), .ZN(n9249)
         );
  INV_X1 U10597 ( .A(n9249), .ZN(n9250) );
  OAI21_X1 U10598 ( .B1(n9836), .B2(n9398), .A(n9250), .ZN(P1_U3265) );
  XNOR2_X1 U10599 ( .A(n9251), .B(n9258), .ZN(n9404) );
  INV_X1 U10600 ( .A(n9252), .ZN(n9253) );
  AOI211_X1 U10601 ( .C1(n9401), .C2(n9267), .A(n9775), .B(n9253), .ZN(n9400)
         );
  INV_X1 U10602 ( .A(n9254), .ZN(n9255) );
  AOI22_X1 U10603 ( .A1(n9823), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n9255), .B2(
        n9822), .ZN(n9256) );
  OAI21_X1 U10604 ( .B1(n9257), .B2(n9825), .A(n9256), .ZN(n9263) );
  XNOR2_X1 U10605 ( .A(n9259), .B(n9258), .ZN(n9261) );
  AOI21_X1 U10606 ( .B1(n9261), .B2(n9821), .A(n9260), .ZN(n9403) );
  NOR2_X1 U10607 ( .A1(n9403), .A2(n9823), .ZN(n9262) );
  AOI211_X1 U10608 ( .C1(n9400), .C2(n9832), .A(n9263), .B(n9262), .ZN(n9264)
         );
  OAI21_X1 U10609 ( .B1(n9404), .B2(n9378), .A(n9264), .ZN(P1_U3266) );
  XNOR2_X1 U10610 ( .A(n9266), .B(n9265), .ZN(n9409) );
  INV_X1 U10611 ( .A(n9267), .ZN(n9268) );
  AOI211_X1 U10612 ( .C1(n9406), .C2(n4463), .A(n9775), .B(n9268), .ZN(n9405)
         );
  AOI22_X1 U10613 ( .A1(n9269), .A2(n9822), .B1(P1_REG2_REG_26__SCAN_IN), .B2(
        n9823), .ZN(n9270) );
  OAI21_X1 U10614 ( .B1(n4637), .B2(n9825), .A(n9270), .ZN(n9276) );
  OAI21_X1 U10615 ( .B1(n8384), .B2(n9272), .A(n9271), .ZN(n9274) );
  AOI21_X1 U10616 ( .B1(n9274), .B2(n9821), .A(n9273), .ZN(n9408) );
  NOR2_X1 U10617 ( .A1(n9408), .A2(n9823), .ZN(n9275) );
  AOI211_X1 U10618 ( .C1(n9405), .C2(n9832), .A(n9276), .B(n9275), .ZN(n9277)
         );
  OAI21_X1 U10619 ( .B1(n9409), .B2(n9378), .A(n9277), .ZN(P1_U3267) );
  XNOR2_X1 U10620 ( .A(n9278), .B(n4352), .ZN(n9414) );
  AOI211_X1 U10621 ( .C1(n9411), .C2(n9292), .A(n9775), .B(n9279), .ZN(n9410)
         );
  AOI22_X1 U10622 ( .A1(n9280), .A2(n9822), .B1(P1_REG2_REG_25__SCAN_IN), .B2(
        n9823), .ZN(n9281) );
  OAI21_X1 U10623 ( .B1(n9282), .B2(n9825), .A(n9281), .ZN(n9288) );
  OAI21_X1 U10624 ( .B1(n4352), .B2(n9284), .A(n9283), .ZN(n9286) );
  AOI21_X1 U10625 ( .B1(n9286), .B2(n9821), .A(n9285), .ZN(n9413) );
  NOR2_X1 U10626 ( .A1(n9413), .A2(n9836), .ZN(n9287) );
  AOI211_X1 U10627 ( .C1(n9410), .C2(n9832), .A(n9288), .B(n9287), .ZN(n9289)
         );
  OAI21_X1 U10628 ( .B1(n9414), .B2(n9378), .A(n9289), .ZN(P1_U3268) );
  XNOR2_X1 U10629 ( .A(n9290), .B(n9297), .ZN(n9419) );
  INV_X1 U10630 ( .A(n9292), .ZN(n9293) );
  AOI211_X1 U10631 ( .C1(n9416), .C2(n9305), .A(n9775), .B(n9293), .ZN(n9415)
         );
  AOI22_X1 U10632 ( .A1(n9294), .A2(n9822), .B1(P1_REG2_REG_24__SCAN_IN), .B2(
        n9823), .ZN(n9295) );
  OAI21_X1 U10633 ( .B1(n9154), .B2(n9825), .A(n9295), .ZN(n9301) );
  AOI211_X1 U10634 ( .C1(n9297), .C2(n9296), .A(n9746), .B(n4387), .ZN(n9299)
         );
  NOR2_X1 U10635 ( .A1(n9299), .A2(n9298), .ZN(n9418) );
  NOR2_X1 U10636 ( .A1(n9418), .A2(n9823), .ZN(n9300) );
  AOI211_X1 U10637 ( .C1(n9415), .C2(n9832), .A(n9301), .B(n9300), .ZN(n9302)
         );
  OAI21_X1 U10638 ( .B1(n9378), .B2(n9419), .A(n9302), .ZN(P1_U3269) );
  XNOR2_X1 U10639 ( .A(n9303), .B(n9304), .ZN(n9424) );
  AOI211_X1 U10640 ( .C1(n9421), .C2(n9319), .A(n9775), .B(n9291), .ZN(n9420)
         );
  AOI22_X1 U10641 ( .A1(n9306), .A2(n9822), .B1(P1_REG2_REG_23__SCAN_IN), .B2(
        n9823), .ZN(n9307) );
  OAI21_X1 U10642 ( .B1(n9308), .B2(n9825), .A(n9307), .ZN(n9316) );
  OAI21_X1 U10643 ( .B1(n9311), .B2(n9310), .A(n9309), .ZN(n9314) );
  INV_X1 U10644 ( .A(n9312), .ZN(n9313) );
  AOI21_X1 U10645 ( .B1(n9314), .B2(n9821), .A(n9313), .ZN(n9423) );
  NOR2_X1 U10646 ( .A1(n9423), .A2(n9823), .ZN(n9315) );
  AOI211_X1 U10647 ( .C1(n9420), .C2(n9832), .A(n9316), .B(n9315), .ZN(n9317)
         );
  OAI21_X1 U10648 ( .B1(n9424), .B2(n9378), .A(n9317), .ZN(P1_U3270) );
  XNOR2_X1 U10649 ( .A(n9318), .B(n9326), .ZN(n9429) );
  INV_X1 U10650 ( .A(n9319), .ZN(n9320) );
  AOI211_X1 U10651 ( .C1(n9426), .C2(n4469), .A(n9775), .B(n9320), .ZN(n9425)
         );
  AOI22_X1 U10652 ( .A1(n9321), .A2(n9822), .B1(n9823), .B2(
        P1_REG2_REG_22__SCAN_IN), .ZN(n9322) );
  OAI21_X1 U10653 ( .B1(n9323), .B2(n9825), .A(n9322), .ZN(n9331) );
  OAI21_X1 U10654 ( .B1(n9326), .B2(n9325), .A(n9324), .ZN(n9329) );
  INV_X1 U10655 ( .A(n9327), .ZN(n9328) );
  AOI21_X1 U10656 ( .B1(n9329), .B2(n9821), .A(n9328), .ZN(n9428) );
  NOR2_X1 U10657 ( .A1(n9428), .A2(n9836), .ZN(n9330) );
  AOI211_X1 U10658 ( .C1(n9425), .C2(n9832), .A(n9331), .B(n9330), .ZN(n9332)
         );
  OAI21_X1 U10659 ( .B1(n9429), .B2(n9378), .A(n9332), .ZN(P1_U3271) );
  XNOR2_X1 U10660 ( .A(n9333), .B(n9340), .ZN(n9433) );
  AOI211_X1 U10661 ( .C1(n8183), .C2(n9350), .A(n9775), .B(n9334), .ZN(n9430)
         );
  OAI22_X1 U10662 ( .A1(n9337), .A2(n9825), .B1(n9336), .B2(n9335), .ZN(n9347)
         );
  OAI21_X1 U10663 ( .B1(n9340), .B2(n9339), .A(n9338), .ZN(n9343) );
  INV_X1 U10664 ( .A(n9341), .ZN(n9342) );
  AOI21_X1 U10665 ( .B1(n9343), .B2(n9821), .A(n9342), .ZN(n9432) );
  NAND2_X1 U10666 ( .A1(n9344), .A2(n9822), .ZN(n9345) );
  AOI21_X1 U10667 ( .B1(n9432), .B2(n9345), .A(n9836), .ZN(n9346) );
  AOI211_X1 U10668 ( .C1(n9430), .C2(n9832), .A(n9347), .B(n9346), .ZN(n9348)
         );
  OAI21_X1 U10669 ( .B1(n9433), .B2(n9378), .A(n9348), .ZN(P1_U3272) );
  XOR2_X1 U10670 ( .A(n9356), .B(n9349), .Z(n9438) );
  INV_X1 U10671 ( .A(n9350), .ZN(n9351) );
  AOI211_X1 U10672 ( .C1(n9435), .C2(n9364), .A(n9775), .B(n9351), .ZN(n9434)
         );
  AOI22_X1 U10673 ( .A1(n9823), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9352), .B2(
        n9822), .ZN(n9353) );
  OAI21_X1 U10674 ( .B1(n9354), .B2(n9825), .A(n9353), .ZN(n9360) );
  XOR2_X1 U10675 ( .A(n9356), .B(n9355), .Z(n9358) );
  AOI21_X1 U10676 ( .B1(n9358), .B2(n9821), .A(n9357), .ZN(n9437) );
  NOR2_X1 U10677 ( .A1(n9437), .A2(n9836), .ZN(n9359) );
  AOI211_X1 U10678 ( .C1(n9434), .C2(n9832), .A(n9360), .B(n9359), .ZN(n9361)
         );
  OAI21_X1 U10679 ( .B1(n9438), .B2(n9378), .A(n9361), .ZN(P1_U3273) );
  XOR2_X1 U10680 ( .A(n9362), .B(n9371), .Z(n9442) );
  INV_X1 U10681 ( .A(n9363), .ZN(n9366) );
  INV_X1 U10682 ( .A(n9364), .ZN(n9365) );
  AOI211_X1 U10683 ( .C1(n8184), .C2(n9366), .A(n9775), .B(n9365), .ZN(n9439)
         );
  INV_X1 U10684 ( .A(n9367), .ZN(n9368) );
  AOI22_X1 U10685 ( .A1(n9823), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9368), .B2(
        n9822), .ZN(n9369) );
  OAI21_X1 U10686 ( .B1(n9370), .B2(n9825), .A(n9369), .ZN(n9376) );
  XOR2_X1 U10687 ( .A(n9372), .B(n9371), .Z(n9374) );
  AOI21_X1 U10688 ( .B1(n9374), .B2(n9821), .A(n9373), .ZN(n9441) );
  NOR2_X1 U10689 ( .A1(n9441), .A2(n9823), .ZN(n9375) );
  AOI211_X1 U10690 ( .C1(n9439), .C2(n9832), .A(n9376), .B(n9375), .ZN(n9377)
         );
  OAI21_X1 U10691 ( .B1(n9378), .B2(n9442), .A(n9377), .ZN(P1_U3274) );
  OAI211_X1 U10692 ( .C1(n9380), .C2(n9911), .A(n9379), .B(n9385), .ZN(n9460)
         );
  NOR2_X1 U10693 ( .A1(n9382), .A2(n9381), .ZN(n9383) );
  MUX2_X1 U10694 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n9460), .S(n9945), .Z(
        P1_U3553) );
  OAI211_X1 U10695 ( .C1(n9387), .C2(n9911), .A(n9386), .B(n9385), .ZN(n9461)
         );
  MUX2_X1 U10696 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n9461), .S(n9945), .Z(
        P1_U3552) );
  NAND2_X1 U10697 ( .A1(n9388), .A2(n9914), .ZN(n9392) );
  NAND3_X1 U10698 ( .A1(n9394), .A2(n9393), .A3(n9914), .ZN(n9399) );
  NAND2_X1 U10699 ( .A1(n9395), .A2(n9919), .ZN(n9396) );
  NAND4_X1 U10700 ( .A1(n9399), .A2(n9398), .A3(n9397), .A4(n9396), .ZN(n9462)
         );
  MUX2_X1 U10701 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n9462), .S(n9945), .Z(
        P1_U3550) );
  AOI21_X1 U10702 ( .B1(n9919), .B2(n9401), .A(n9400), .ZN(n9402) );
  OAI211_X1 U10703 ( .C1(n9404), .C2(n9457), .A(n9403), .B(n9402), .ZN(n9463)
         );
  MUX2_X1 U10704 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9463), .S(n9945), .Z(
        P1_U3549) );
  AOI21_X1 U10705 ( .B1(n9919), .B2(n9406), .A(n9405), .ZN(n9407) );
  OAI211_X1 U10706 ( .C1(n9409), .C2(n9457), .A(n9408), .B(n9407), .ZN(n9464)
         );
  MUX2_X1 U10707 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9464), .S(n9945), .Z(
        P1_U3548) );
  AOI21_X1 U10708 ( .B1(n9919), .B2(n9411), .A(n9410), .ZN(n9412) );
  OAI211_X1 U10709 ( .C1(n9414), .C2(n9457), .A(n9413), .B(n9412), .ZN(n9465)
         );
  MUX2_X1 U10710 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9465), .S(n9945), .Z(
        P1_U3547) );
  AOI21_X1 U10711 ( .B1(n9919), .B2(n9416), .A(n9415), .ZN(n9417) );
  OAI211_X1 U10712 ( .C1(n9419), .C2(n9457), .A(n9418), .B(n9417), .ZN(n9466)
         );
  MUX2_X1 U10713 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9466), .S(n9945), .Z(
        P1_U3546) );
  AOI21_X1 U10714 ( .B1(n9919), .B2(n9421), .A(n9420), .ZN(n9422) );
  OAI211_X1 U10715 ( .C1(n9424), .C2(n9457), .A(n9423), .B(n9422), .ZN(n9467)
         );
  MUX2_X1 U10716 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9467), .S(n9945), .Z(
        P1_U3545) );
  AOI21_X1 U10717 ( .B1(n9919), .B2(n9426), .A(n9425), .ZN(n9427) );
  OAI211_X1 U10718 ( .C1(n9429), .C2(n9457), .A(n9428), .B(n9427), .ZN(n9468)
         );
  MUX2_X1 U10719 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9468), .S(n9945), .Z(
        P1_U3544) );
  AOI21_X1 U10720 ( .B1(n9919), .B2(n8183), .A(n9430), .ZN(n9431) );
  OAI211_X1 U10721 ( .C1(n9433), .C2(n9457), .A(n9432), .B(n9431), .ZN(n9469)
         );
  MUX2_X1 U10722 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9469), .S(n9945), .Z(
        P1_U3543) );
  AOI21_X1 U10723 ( .B1(n9919), .B2(n9435), .A(n9434), .ZN(n9436) );
  OAI211_X1 U10724 ( .C1(n9438), .C2(n9457), .A(n9437), .B(n9436), .ZN(n9470)
         );
  MUX2_X1 U10725 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9470), .S(n9945), .Z(
        P1_U3542) );
  AOI21_X1 U10726 ( .B1(n9919), .B2(n8184), .A(n9439), .ZN(n9440) );
  OAI211_X1 U10727 ( .C1(n9442), .C2(n9457), .A(n9441), .B(n9440), .ZN(n9471)
         );
  MUX2_X1 U10728 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9471), .S(n9945), .Z(
        P1_U3541) );
  AOI211_X1 U10729 ( .C1(n9919), .C2(n9445), .A(n9444), .B(n9443), .ZN(n9446)
         );
  OAI21_X1 U10730 ( .B1(n9457), .B2(n9447), .A(n9446), .ZN(n9472) );
  MUX2_X1 U10731 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9472), .S(n9945), .Z(
        P1_U3540) );
  AOI21_X1 U10732 ( .B1(n9919), .B2(n9449), .A(n9448), .ZN(n9450) );
  OAI211_X1 U10733 ( .C1(n9452), .C2(n9457), .A(n9451), .B(n9450), .ZN(n9473)
         );
  MUX2_X1 U10734 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9473), .S(n9945), .Z(
        P1_U3539) );
  AOI21_X1 U10735 ( .B1(n9919), .B2(n9454), .A(n9453), .ZN(n9455) );
  OAI211_X1 U10736 ( .C1(n9458), .C2(n9457), .A(n9456), .B(n9455), .ZN(n9474)
         );
  MUX2_X1 U10737 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9474), .S(n9945), .Z(
        P1_U3538) );
  MUX2_X1 U10738 ( .A(n9459), .B(P1_REG1_REG_0__SCAN_IN), .S(n9943), .Z(
        P1_U3522) );
  MUX2_X1 U10739 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n9460), .S(n9927), .Z(
        P1_U3521) );
  MUX2_X1 U10740 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n9461), .S(n9927), .Z(
        P1_U3520) );
  MUX2_X1 U10741 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n9462), .S(n9927), .Z(
        P1_U3518) );
  MUX2_X1 U10742 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9463), .S(n9927), .Z(
        P1_U3517) );
  MUX2_X1 U10743 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9464), .S(n9927), .Z(
        P1_U3516) );
  MUX2_X1 U10744 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9465), .S(n9927), .Z(
        P1_U3515) );
  MUX2_X1 U10745 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9466), .S(n9927), .Z(
        P1_U3514) );
  MUX2_X1 U10746 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9467), .S(n9927), .Z(
        P1_U3513) );
  MUX2_X1 U10747 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9468), .S(n9927), .Z(
        P1_U3512) );
  MUX2_X1 U10748 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9469), .S(n9927), .Z(
        P1_U3511) );
  MUX2_X1 U10749 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9470), .S(n9927), .Z(
        P1_U3510) );
  MUX2_X1 U10750 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9471), .S(n9927), .Z(
        P1_U3509) );
  MUX2_X1 U10751 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9472), .S(n9927), .Z(
        P1_U3507) );
  MUX2_X1 U10752 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9473), .S(n9927), .Z(
        P1_U3504) );
  MUX2_X1 U10753 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n9474), .S(n9927), .Z(
        P1_U3501) );
  MUX2_X1 U10754 ( .A(n9477), .B(P1_D_REG_1__SCAN_IN), .S(n4345), .Z(P1_U3440)
         );
  MUX2_X1 U10755 ( .A(n9478), .B(P1_D_REG_0__SCAN_IN), .S(n4345), .Z(P1_U3439)
         );
  INV_X1 U10756 ( .A(n9479), .ZN(n9480) );
  MUX2_X1 U10757 ( .A(n9480), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  INV_X1 U10758 ( .A(n9609), .ZN(n9728) );
  INV_X1 U10759 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n9492) );
  AOI211_X1 U10760 ( .C1(n9483), .C2(n9482), .A(n9481), .B(n9699), .ZN(n9488)
         );
  AOI211_X1 U10761 ( .C1(n9486), .C2(n9485), .A(n9484), .B(n9702), .ZN(n9487)
         );
  AOI211_X1 U10762 ( .C1(n9709), .C2(n9489), .A(n9488), .B(n9487), .ZN(n9491)
         );
  NAND2_X1 U10763 ( .A1(P1_REG3_REG_10__SCAN_IN), .A2(P1_U3086), .ZN(n9490) );
  OAI211_X1 U10764 ( .C1(n9728), .C2(n9492), .A(n9491), .B(n9490), .ZN(
        P1_U3253) );
  INV_X1 U10765 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n9507) );
  AOI21_X1 U10766 ( .B1(n9495), .B2(n9494), .A(n9493), .ZN(n9496) );
  NAND2_X1 U10767 ( .A1(n9713), .A2(n9496), .ZN(n9502) );
  AOI21_X1 U10768 ( .B1(n9499), .B2(n9498), .A(n9497), .ZN(n9500) );
  NAND2_X1 U10769 ( .A1(n9718), .A2(n9500), .ZN(n9501) );
  OAI211_X1 U10770 ( .C1(n9724), .C2(n9503), .A(n9502), .B(n9501), .ZN(n9504)
         );
  INV_X1 U10771 ( .A(n9504), .ZN(n9506) );
  NAND2_X1 U10772 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3086), .ZN(n9505) );
  OAI211_X1 U10773 ( .C1(n9728), .C2(n9507), .A(n9506), .B(n9505), .ZN(
        P1_U3250) );
  INV_X1 U10774 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n9522) );
  AOI21_X1 U10775 ( .B1(n9510), .B2(n9509), .A(n9508), .ZN(n9511) );
  NAND2_X1 U10776 ( .A1(n9713), .A2(n9511), .ZN(n9517) );
  AOI21_X1 U10777 ( .B1(n9514), .B2(n9513), .A(n9512), .ZN(n9515) );
  NAND2_X1 U10778 ( .A1(n9718), .A2(n9515), .ZN(n9516) );
  OAI211_X1 U10779 ( .C1(n9724), .C2(n9518), .A(n9517), .B(n9516), .ZN(n9519)
         );
  INV_X1 U10780 ( .A(n9519), .ZN(n9521) );
  NAND2_X1 U10781 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_U3086), .ZN(n9520) );
  OAI211_X1 U10782 ( .C1(n9522), .C2(n9728), .A(n9521), .B(n9520), .ZN(
        P1_U3246) );
  INV_X1 U10783 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n9536) );
  AOI21_X1 U10784 ( .B1(n9525), .B2(n9524), .A(n9523), .ZN(n9526) );
  NAND2_X1 U10785 ( .A1(n9718), .A2(n9526), .ZN(n9531) );
  AOI21_X1 U10786 ( .B1(n9528), .B2(n4379), .A(n9527), .ZN(n9529) );
  NAND2_X1 U10787 ( .A1(n9713), .A2(n9529), .ZN(n9530) );
  OAI211_X1 U10788 ( .C1(n9724), .C2(n9532), .A(n9531), .B(n9530), .ZN(n9533)
         );
  INV_X1 U10789 ( .A(n9533), .ZN(n9535) );
  NAND2_X1 U10790 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_U3086), .ZN(n9534) );
  OAI211_X1 U10791 ( .C1(n9728), .C2(n9536), .A(n9535), .B(n9534), .ZN(
        P1_U3251) );
  OR2_X1 U10792 ( .A1(n9537), .A2(n5609), .ZN(n9541) );
  NAND2_X1 U10793 ( .A1(n9539), .A2(n9538), .ZN(n9540) );
  OAI211_X1 U10794 ( .C1(n9543), .C2(n9542), .A(n9541), .B(n9540), .ZN(n9544)
         );
  INV_X1 U10795 ( .A(n9544), .ZN(n9545) );
  OAI21_X1 U10796 ( .B1(n9546), .B2(n5075), .A(n9545), .ZN(P2_U3172) );
  NOR2_X1 U10797 ( .A1(n9547), .A2(n9746), .ZN(n9554) );
  OAI21_X1 U10798 ( .B1(n9550), .B2(n9549), .A(n9548), .ZN(n9553) );
  INV_X1 U10799 ( .A(n9551), .ZN(n9552) );
  AOI21_X1 U10800 ( .B1(n9554), .B2(n9553), .A(n9552), .ZN(n9563) );
  AOI222_X1 U10801 ( .A1(n7427), .A2(n9753), .B1(P1_REG2_REG_15__SCAN_IN), 
        .B2(n9836), .C1(n9822), .C2(n9555), .ZN(n9561) );
  XNOR2_X1 U10802 ( .A(n9557), .B(n9556), .ZN(n9565) );
  OAI211_X1 U10803 ( .C1(n4423), .C2(n7446), .A(n9829), .B(n9558), .ZN(n9562)
         );
  INV_X1 U10804 ( .A(n9562), .ZN(n9559) );
  AOI22_X1 U10805 ( .A1(n9565), .A2(n9809), .B1(n9832), .B2(n9559), .ZN(n9560)
         );
  OAI211_X1 U10806 ( .C1(n9836), .C2(n9563), .A(n9561), .B(n9560), .ZN(
        P1_U3278) );
  OAI211_X1 U10807 ( .C1(n7446), .C2(n9911), .A(n9563), .B(n9562), .ZN(n9564)
         );
  AOI21_X1 U10808 ( .B1(n9565), .B2(n9914), .A(n9564), .ZN(n9566) );
  AOI22_X1 U10809 ( .A1(n9945), .A2(n9566), .B1(n7279), .B2(n9943), .ZN(
        P1_U3537) );
  AOI22_X1 U10810 ( .A1(n9927), .A2(n9566), .B1(n7278), .B2(n9926), .ZN(
        P1_U3498) );
  XNOR2_X1 U10811 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XOR2_X1 U10812 ( .A(n4927), .B(P1_RD_REG_SCAN_IN), .Z(U126) );
  AOI21_X1 U10813 ( .B1(n9569), .B2(n9568), .A(n9567), .ZN(n9606) );
  OAI21_X1 U10814 ( .B1(n9569), .B2(P1_REG1_REG_0__SCAN_IN), .A(n9606), .ZN(
        n9571) );
  XNOR2_X1 U10815 ( .A(n9571), .B(n9570), .ZN(n9574) );
  AOI22_X1 U10816 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(n9609), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n9572) );
  OAI21_X1 U10817 ( .B1(n9574), .B2(n9573), .A(n9572), .ZN(P1_U3243) );
  AOI22_X1 U10818 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(n9609), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n9588) );
  NAND2_X1 U10819 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n9576) );
  AOI21_X1 U10820 ( .B1(n9577), .B2(n9576), .A(n9575), .ZN(n9578) );
  NAND2_X1 U10821 ( .A1(n9713), .A2(n9578), .ZN(n9584) );
  AOI21_X1 U10822 ( .B1(n9581), .B2(n9580), .A(n9579), .ZN(n9582) );
  NAND2_X1 U10823 ( .A1(n9718), .A2(n9582), .ZN(n9583) );
  OAI211_X1 U10824 ( .C1(n9724), .C2(n9585), .A(n9584), .B(n9583), .ZN(n9586)
         );
  INV_X1 U10825 ( .A(n9586), .ZN(n9587) );
  NAND2_X1 U10826 ( .A1(n9588), .A2(n9587), .ZN(P1_U3244) );
  AOI22_X1 U10827 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(n9609), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n9608) );
  AOI21_X1 U10828 ( .B1(n9591), .B2(n9590), .A(n9589), .ZN(n9592) );
  NAND2_X1 U10829 ( .A1(n9713), .A2(n9592), .ZN(n9598) );
  AOI21_X1 U10830 ( .B1(n9595), .B2(n9594), .A(n9593), .ZN(n9596) );
  NAND2_X1 U10831 ( .A1(n9718), .A2(n9596), .ZN(n9597) );
  OAI211_X1 U10832 ( .C1(n9724), .C2(n9599), .A(n9598), .B(n9597), .ZN(n9600)
         );
  INV_X1 U10833 ( .A(n9600), .ZN(n9607) );
  MUX2_X1 U10834 ( .A(n9602), .B(n9601), .S(n6484), .Z(n9604) );
  NAND2_X1 U10835 ( .A1(n9604), .A2(n9603), .ZN(n9605) );
  OAI211_X1 U10836 ( .C1(P1_IR_REG_0__SCAN_IN), .C2(n9606), .A(n9605), .B(
        P1_U3973), .ZN(n9622) );
  NAND3_X1 U10837 ( .A1(n9608), .A2(n9607), .A3(n9622), .ZN(P1_U3245) );
  AOI22_X1 U10838 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(n9609), .B1(
        P1_REG3_REG_4__SCAN_IN), .B2(P1_U3086), .ZN(n9624) );
  AOI21_X1 U10839 ( .B1(n9612), .B2(n9611), .A(n9610), .ZN(n9613) );
  NAND2_X1 U10840 ( .A1(n9713), .A2(n9613), .ZN(n9619) );
  AOI21_X1 U10841 ( .B1(n9616), .B2(n9615), .A(n9614), .ZN(n9617) );
  NAND2_X1 U10842 ( .A1(n9718), .A2(n9617), .ZN(n9618) );
  OAI211_X1 U10843 ( .C1(n9724), .C2(n9620), .A(n9619), .B(n9618), .ZN(n9621)
         );
  INV_X1 U10844 ( .A(n9621), .ZN(n9623) );
  NAND3_X1 U10845 ( .A1(n9624), .A2(n9623), .A3(n9622), .ZN(P1_U3247) );
  INV_X1 U10846 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n9640) );
  AOI21_X1 U10847 ( .B1(n9627), .B2(n9626), .A(n9625), .ZN(n9628) );
  NAND2_X1 U10848 ( .A1(n9718), .A2(n9628), .ZN(n9634) );
  AOI21_X1 U10849 ( .B1(n9631), .B2(n9630), .A(n9629), .ZN(n9632) );
  NAND2_X1 U10850 ( .A1(n9713), .A2(n9632), .ZN(n9633) );
  OAI211_X1 U10851 ( .C1(n9724), .C2(n9635), .A(n9634), .B(n9633), .ZN(n9636)
         );
  INV_X1 U10852 ( .A(n9636), .ZN(n9639) );
  NAND2_X1 U10853 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n9638) );
  OAI211_X1 U10854 ( .C1(n9728), .C2(n9640), .A(n9639), .B(n9638), .ZN(
        P1_U3248) );
  INV_X1 U10855 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n9655) );
  AOI21_X1 U10856 ( .B1(n9643), .B2(n9642), .A(n9641), .ZN(n9644) );
  NAND2_X1 U10857 ( .A1(n9713), .A2(n9644), .ZN(n9650) );
  AOI21_X1 U10858 ( .B1(n9647), .B2(n9646), .A(n9645), .ZN(n9648) );
  NAND2_X1 U10859 ( .A1(n9718), .A2(n9648), .ZN(n9649) );
  OAI211_X1 U10860 ( .C1(n9724), .C2(n9651), .A(n9650), .B(n9649), .ZN(n9652)
         );
  INV_X1 U10861 ( .A(n9652), .ZN(n9654) );
  NAND2_X1 U10862 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_U3086), .ZN(n9653) );
  OAI211_X1 U10863 ( .C1(n9728), .C2(n9655), .A(n9654), .B(n9653), .ZN(
        P1_U3249) );
  INV_X1 U10864 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n9671) );
  INV_X1 U10865 ( .A(n9656), .ZN(n9667) );
  AOI21_X1 U10866 ( .B1(n9659), .B2(n9658), .A(n9657), .ZN(n9660) );
  NAND2_X1 U10867 ( .A1(n9713), .A2(n9660), .ZN(n9666) );
  AOI21_X1 U10868 ( .B1(n9663), .B2(n9662), .A(n9661), .ZN(n9664) );
  NAND2_X1 U10869 ( .A1(n9718), .A2(n9664), .ZN(n9665) );
  OAI211_X1 U10870 ( .C1(n9724), .C2(n9667), .A(n9666), .B(n9665), .ZN(n9668)
         );
  INV_X1 U10871 ( .A(n9668), .ZN(n9670) );
  NAND2_X1 U10872 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n9669) );
  OAI211_X1 U10873 ( .C1(n9728), .C2(n9671), .A(n9670), .B(n9669), .ZN(
        P1_U3254) );
  INV_X1 U10874 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n9683) );
  AOI211_X1 U10875 ( .C1(n9674), .C2(n9673), .A(n9672), .B(n9699), .ZN(n9679)
         );
  AOI211_X1 U10876 ( .C1(n9677), .C2(n9676), .A(n9675), .B(n9702), .ZN(n9678)
         );
  AOI211_X1 U10877 ( .C1(n9709), .C2(n9680), .A(n9679), .B(n9678), .ZN(n9682)
         );
  NAND2_X1 U10878 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3086), .ZN(n9681) );
  OAI211_X1 U10879 ( .C1(n9728), .C2(n9683), .A(n9682), .B(n9681), .ZN(
        P1_U3256) );
  INV_X1 U10880 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n9698) );
  AOI21_X1 U10881 ( .B1(n9686), .B2(n9685), .A(n9684), .ZN(n9687) );
  NAND2_X1 U10882 ( .A1(n9713), .A2(n9687), .ZN(n9693) );
  AOI21_X1 U10883 ( .B1(n9690), .B2(n9689), .A(n9688), .ZN(n9691) );
  NAND2_X1 U10884 ( .A1(n9718), .A2(n9691), .ZN(n9692) );
  OAI211_X1 U10885 ( .C1(n9724), .C2(n9694), .A(n9693), .B(n9692), .ZN(n9695)
         );
  INV_X1 U10886 ( .A(n9695), .ZN(n9697) );
  NAND2_X1 U10887 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n9696) );
  OAI211_X1 U10888 ( .C1(n9728), .C2(n9698), .A(n9697), .B(n9696), .ZN(
        P1_U3257) );
  INV_X1 U10889 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n9712) );
  AOI211_X1 U10890 ( .C1(n9701), .C2(n7279), .A(n9700), .B(n9699), .ZN(n9707)
         );
  AOI211_X1 U10891 ( .C1(n9705), .C2(n9704), .A(n9703), .B(n9702), .ZN(n9706)
         );
  AOI211_X1 U10892 ( .C1(n9709), .C2(n9708), .A(n9707), .B(n9706), .ZN(n9711)
         );
  NAND2_X1 U10893 ( .A1(P1_REG3_REG_15__SCAN_IN), .A2(P1_U3086), .ZN(n9710) );
  OAI211_X1 U10894 ( .C1(n9728), .C2(n9712), .A(n9711), .B(n9710), .ZN(
        P1_U3258) );
  OAI211_X1 U10895 ( .C1(n9716), .C2(n9715), .A(n9714), .B(n9713), .ZN(n9722)
         );
  OAI211_X1 U10896 ( .C1(n9720), .C2(n9719), .A(n9718), .B(n9717), .ZN(n9721)
         );
  OAI211_X1 U10897 ( .C1(n9724), .C2(n9723), .A(n9722), .B(n9721), .ZN(n9725)
         );
  INV_X1 U10898 ( .A(n9725), .ZN(n9727) );
  OAI211_X1 U10899 ( .C1(n9728), .C2(n10142), .A(n9727), .B(n9726), .ZN(
        P1_U3261) );
  XOR2_X1 U10900 ( .A(n9729), .B(n9735), .Z(n9731) );
  AOI21_X1 U10901 ( .B1(n9731), .B2(n9821), .A(n9730), .ZN(n9910) );
  INV_X1 U10902 ( .A(n9732), .ZN(n9733) );
  AOI222_X1 U10903 ( .A1(n9734), .A2(n9753), .B1(n9733), .B2(n9822), .C1(
        P1_REG2_REG_13__SCAN_IN), .C2(n9836), .ZN(n9740) );
  XNOR2_X1 U10904 ( .A(n9736), .B(n9735), .ZN(n9915) );
  OAI211_X1 U10905 ( .C1(n7270), .C2(n9912), .A(n9829), .B(n9737), .ZN(n9909)
         );
  INV_X1 U10906 ( .A(n9909), .ZN(n9738) );
  AOI22_X1 U10907 ( .A1(n9915), .A2(n9809), .B1(n9832), .B2(n9738), .ZN(n9739)
         );
  OAI211_X1 U10908 ( .C1(n9836), .C2(n9910), .A(n9740), .B(n9739), .ZN(
        P1_U3280) );
  XNOR2_X1 U10909 ( .A(n9742), .B(n9741), .ZN(n9902) );
  INV_X1 U10910 ( .A(n9817), .ZN(n9925) );
  INV_X1 U10911 ( .A(n9743), .ZN(n9748) );
  AOI21_X1 U10912 ( .B1(n7148), .B2(n9745), .A(n9744), .ZN(n9747) );
  NOR3_X1 U10913 ( .A1(n9748), .A2(n9747), .A3(n9746), .ZN(n9750) );
  AOI211_X1 U10914 ( .C1(n9902), .C2(n9925), .A(n9750), .B(n9749), .ZN(n9899)
         );
  INV_X1 U10915 ( .A(n9751), .ZN(n9752) );
  AOI222_X1 U10916 ( .A1(n7173), .A2(n9753), .B1(n9752), .B2(n9822), .C1(
        P1_REG2_REG_11__SCAN_IN), .C2(n9836), .ZN(n9761) );
  INV_X1 U10917 ( .A(n9754), .ZN(n9833) );
  INV_X1 U10918 ( .A(n9755), .ZN(n9758) );
  INV_X1 U10919 ( .A(n9756), .ZN(n9757) );
  OAI211_X1 U10920 ( .C1(n9898), .C2(n9758), .A(n9757), .B(n9829), .ZN(n9897)
         );
  INV_X1 U10921 ( .A(n9897), .ZN(n9759) );
  AOI22_X1 U10922 ( .A1(n9902), .A2(n9833), .B1(n9832), .B2(n9759), .ZN(n9760)
         );
  OAI211_X1 U10923 ( .C1(n9836), .C2(n9899), .A(n9761), .B(n9760), .ZN(
        P1_U3282) );
  INV_X1 U10924 ( .A(n9762), .ZN(n9763) );
  OAI21_X1 U10925 ( .B1(n4422), .B2(n9764), .A(n9763), .ZN(n9768) );
  XNOR2_X1 U10926 ( .A(n9765), .B(n4422), .ZN(n9876) );
  NOR2_X1 U10927 ( .A1(n9876), .A2(n9817), .ZN(n9766) );
  AOI211_X1 U10928 ( .C1(n9821), .C2(n9768), .A(n9767), .B(n9766), .ZN(n9875)
         );
  NOR2_X1 U10929 ( .A1(n9799), .A2(n9769), .ZN(n9770) );
  AOI21_X1 U10930 ( .B1(n9836), .B2(P1_REG2_REG_7__SCAN_IN), .A(n9770), .ZN(
        n9771) );
  OAI21_X1 U10931 ( .B1(n9825), .B2(n9772), .A(n9771), .ZN(n9773) );
  INV_X1 U10932 ( .A(n9773), .ZN(n9779) );
  INV_X1 U10933 ( .A(n9876), .ZN(n9777) );
  AOI211_X1 U10934 ( .C1(n9873), .C2(n9776), .A(n9775), .B(n9774), .ZN(n9872)
         );
  AOI22_X1 U10935 ( .A1(n9777), .A2(n9833), .B1(n9832), .B2(n9872), .ZN(n9778)
         );
  OAI211_X1 U10936 ( .C1(n9836), .C2(n9875), .A(n9779), .B(n9778), .ZN(
        P1_U3286) );
  XNOR2_X1 U10937 ( .A(n9780), .B(n9781), .ZN(n9784) );
  INV_X1 U10938 ( .A(n9782), .ZN(n9783) );
  AOI21_X1 U10939 ( .B1(n9784), .B2(n9821), .A(n9783), .ZN(n9862) );
  NOR2_X1 U10940 ( .A1(n9799), .A2(n9785), .ZN(n9786) );
  AOI21_X1 U10941 ( .B1(n9836), .B2(P1_REG2_REG_5__SCAN_IN), .A(n9786), .ZN(
        n9787) );
  OAI21_X1 U10942 ( .B1(n9825), .B2(n9861), .A(n9787), .ZN(n9788) );
  INV_X1 U10943 ( .A(n9788), .ZN(n9795) );
  XNOR2_X1 U10944 ( .A(n9789), .B(n9790), .ZN(n9865) );
  OAI211_X1 U10945 ( .C1(n9792), .C2(n9861), .A(n9791), .B(n9829), .ZN(n9860)
         );
  INV_X1 U10946 ( .A(n9860), .ZN(n9793) );
  AOI22_X1 U10947 ( .A1(n9865), .A2(n9809), .B1(n9832), .B2(n9793), .ZN(n9794)
         );
  OAI211_X1 U10948 ( .C1(n9836), .C2(n9862), .A(n9795), .B(n9794), .ZN(
        P1_U3288) );
  XNOR2_X1 U10949 ( .A(n8191), .B(n9796), .ZN(n9798) );
  AOI21_X1 U10950 ( .B1(n9798), .B2(n9821), .A(n9797), .ZN(n9850) );
  NOR2_X1 U10951 ( .A1(n9799), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n9800) );
  AOI21_X1 U10952 ( .B1(n9836), .B2(P1_REG2_REG_3__SCAN_IN), .A(n9800), .ZN(
        n9801) );
  OAI21_X1 U10953 ( .B1(n9825), .B2(n9849), .A(n9801), .ZN(n9802) );
  INV_X1 U10954 ( .A(n9802), .ZN(n9811) );
  XNOR2_X1 U10955 ( .A(n9803), .B(n9804), .ZN(n9853) );
  INV_X1 U10956 ( .A(n9805), .ZN(n9807) );
  OAI211_X1 U10957 ( .C1(n9807), .C2(n9849), .A(n9829), .B(n9806), .ZN(n9848)
         );
  INV_X1 U10958 ( .A(n9848), .ZN(n9808) );
  AOI22_X1 U10959 ( .A1(n9853), .A2(n9809), .B1(n9832), .B2(n9808), .ZN(n9810)
         );
  OAI211_X1 U10960 ( .C1(n9836), .C2(n9850), .A(n9811), .B(n9810), .ZN(
        P1_U3290) );
  OAI21_X1 U10961 ( .B1(n9813), .B2(n9815), .A(n9812), .ZN(n9820) );
  INV_X1 U10962 ( .A(n9814), .ZN(n9819) );
  XOR2_X1 U10963 ( .A(n9816), .B(n9815), .Z(n9827) );
  NOR2_X1 U10964 ( .A1(n9827), .A2(n9817), .ZN(n9818) );
  AOI211_X1 U10965 ( .C1(n9821), .C2(n9820), .A(n9819), .B(n9818), .ZN(n9839)
         );
  AOI22_X1 U10966 ( .A1(n9823), .A2(P1_REG2_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(n9822), .ZN(n9824) );
  OAI21_X1 U10967 ( .B1(n9825), .B2(n6626), .A(n9824), .ZN(n9826) );
  INV_X1 U10968 ( .A(n9826), .ZN(n9835) );
  INV_X1 U10969 ( .A(n9827), .ZN(n9842) );
  OAI211_X1 U10970 ( .C1(n6626), .C2(n9830), .A(n9829), .B(n9828), .ZN(n9838)
         );
  INV_X1 U10971 ( .A(n9838), .ZN(n9831) );
  AOI22_X1 U10972 ( .A1(n9842), .A2(n9833), .B1(n9832), .B2(n9831), .ZN(n9834)
         );
  OAI211_X1 U10973 ( .C1(n9836), .C2(n9839), .A(n9835), .B(n9834), .ZN(
        P1_U3292) );
  AND2_X1 U10974 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n4345), .ZN(P1_U3294) );
  AND2_X1 U10975 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n4345), .ZN(P1_U3295) );
  AND2_X1 U10976 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n4345), .ZN(P1_U3296) );
  AND2_X1 U10977 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n4345), .ZN(P1_U3297) );
  AND2_X1 U10978 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n4345), .ZN(P1_U3298) );
  AND2_X1 U10979 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n4345), .ZN(P1_U3299) );
  AND2_X1 U10980 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n4345), .ZN(P1_U3300) );
  AND2_X1 U10981 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n4345), .ZN(P1_U3301) );
  AND2_X1 U10982 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n4345), .ZN(P1_U3302) );
  AND2_X1 U10983 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n4345), .ZN(P1_U3303) );
  AND2_X1 U10984 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n4345), .ZN(P1_U3304) );
  AND2_X1 U10985 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n4345), .ZN(P1_U3305) );
  AND2_X1 U10986 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n4345), .ZN(P1_U3306) );
  AND2_X1 U10987 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n4345), .ZN(P1_U3307) );
  AND2_X1 U10988 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n4345), .ZN(P1_U3308) );
  AND2_X1 U10989 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n4345), .ZN(P1_U3309) );
  AND2_X1 U10990 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n4345), .ZN(P1_U3310) );
  AND2_X1 U10991 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n4345), .ZN(P1_U3311) );
  AND2_X1 U10992 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n4345), .ZN(P1_U3312) );
  AND2_X1 U10993 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n4345), .ZN(P1_U3313) );
  AND2_X1 U10994 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n4345), .ZN(P1_U3314) );
  AND2_X1 U10995 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n4345), .ZN(P1_U3315) );
  AND2_X1 U10996 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n4345), .ZN(P1_U3316) );
  AND2_X1 U10997 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n4345), .ZN(P1_U3317) );
  AND2_X1 U10998 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n4345), .ZN(P1_U3318) );
  AND2_X1 U10999 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n4345), .ZN(P1_U3319) );
  AND2_X1 U11000 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n4345), .ZN(P1_U3320) );
  AND2_X1 U11001 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n4345), .ZN(P1_U3321) );
  AND2_X1 U11002 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n4345), .ZN(P1_U3322) );
  AND2_X1 U11003 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n4345), .ZN(P1_U3323) );
  OAI21_X1 U11004 ( .B1(n6626), .B2(n9911), .A(n9838), .ZN(n9841) );
  INV_X1 U11005 ( .A(n9839), .ZN(n9840) );
  AOI211_X1 U11006 ( .C1(n9903), .C2(n9842), .A(n9841), .B(n9840), .ZN(n9928)
         );
  AOI22_X1 U11007 ( .A1(n9927), .A2(n9928), .B1(n6082), .B2(n9926), .ZN(
        P1_U3456) );
  OAI21_X1 U11008 ( .B1(n9844), .B2(n9911), .A(n9843), .ZN(n9846) );
  AOI211_X1 U11009 ( .C1(n9914), .C2(n9847), .A(n9846), .B(n9845), .ZN(n9929)
         );
  AOI22_X1 U11010 ( .A1(n9927), .A2(n9929), .B1(n6185), .B2(n9926), .ZN(
        P1_U3459) );
  OAI21_X1 U11011 ( .B1(n9849), .B2(n9911), .A(n9848), .ZN(n9852) );
  INV_X1 U11012 ( .A(n9850), .ZN(n9851) );
  AOI211_X1 U11013 ( .C1(n9914), .C2(n9853), .A(n9852), .B(n9851), .ZN(n9930)
         );
  AOI22_X1 U11014 ( .A1(n9927), .A2(n9930), .B1(n6214), .B2(n9926), .ZN(
        P1_U3462) );
  OAI21_X1 U11015 ( .B1(n9855), .B2(n9911), .A(n9854), .ZN(n9856) );
  AOI21_X1 U11016 ( .B1(n9857), .B2(n9914), .A(n9856), .ZN(n9858) );
  AND2_X1 U11017 ( .A1(n9859), .A2(n9858), .ZN(n9931) );
  AOI22_X1 U11018 ( .A1(n9927), .A2(n9931), .B1(n6263), .B2(n9926), .ZN(
        P1_U3465) );
  OAI21_X1 U11019 ( .B1(n9861), .B2(n9911), .A(n9860), .ZN(n9864) );
  INV_X1 U11020 ( .A(n9862), .ZN(n9863) );
  AOI211_X1 U11021 ( .C1(n9914), .C2(n9865), .A(n9864), .B(n9863), .ZN(n9932)
         );
  AOI22_X1 U11022 ( .A1(n9927), .A2(n9932), .B1(n6424), .B2(n9926), .ZN(
        P1_U3468) );
  AND2_X1 U11023 ( .A1(n9866), .A2(n9914), .ZN(n9870) );
  OAI21_X1 U11024 ( .B1(n6643), .B2(n9911), .A(n9867), .ZN(n9868) );
  NOR3_X1 U11025 ( .A1(n9870), .A2(n9869), .A3(n9868), .ZN(n9933) );
  INV_X1 U11026 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n9871) );
  AOI22_X1 U11027 ( .A1(n9927), .A2(n9933), .B1(n9871), .B2(n9926), .ZN(
        P1_U3471) );
  AOI21_X1 U11028 ( .B1(n9919), .B2(n9873), .A(n9872), .ZN(n9874) );
  OAI211_X1 U11029 ( .C1(n9876), .C2(n9921), .A(n9875), .B(n9874), .ZN(n9877)
         );
  INV_X1 U11030 ( .A(n9877), .ZN(n9934) );
  AOI22_X1 U11031 ( .A1(n9927), .A2(n9934), .B1(n6583), .B2(n9926), .ZN(
        P1_U3474) );
  AND2_X1 U11032 ( .A1(n9878), .A2(n9925), .ZN(n9883) );
  NAND2_X1 U11033 ( .A1(n9878), .A2(n9903), .ZN(n9880) );
  OAI211_X1 U11034 ( .C1(n9881), .C2(n9911), .A(n9880), .B(n9879), .ZN(n9882)
         );
  NOR3_X1 U11035 ( .A1(n9884), .A2(n9883), .A3(n9882), .ZN(n9936) );
  AOI22_X1 U11036 ( .A1(n9927), .A2(n9936), .B1(n6660), .B2(n9926), .ZN(
        P1_U3477) );
  INV_X1 U11037 ( .A(n9885), .ZN(n9886) );
  OAI211_X1 U11038 ( .C1(n9888), .C2(n9911), .A(n9887), .B(n9886), .ZN(n9890)
         );
  AOI211_X1 U11039 ( .C1(n9914), .C2(n9891), .A(n9890), .B(n9889), .ZN(n9937)
         );
  AOI22_X1 U11040 ( .A1(n9927), .A2(n9937), .B1(n6677), .B2(n9926), .ZN(
        P1_U3480) );
  OAI211_X1 U11041 ( .C1(n9894), .C2(n9911), .A(n9893), .B(n9892), .ZN(n9895)
         );
  AOI21_X1 U11042 ( .B1(n9896), .B2(n9914), .A(n9895), .ZN(n9938) );
  AOI22_X1 U11043 ( .A1(n9927), .A2(n9938), .B1(n6705), .B2(n9926), .ZN(
        P1_U3483) );
  OAI21_X1 U11044 ( .B1(n9898), .B2(n9911), .A(n9897), .ZN(n9901) );
  INV_X1 U11045 ( .A(n9899), .ZN(n9900) );
  AOI211_X1 U11046 ( .C1(n9903), .C2(n9902), .A(n9901), .B(n9900), .ZN(n9939)
         );
  AOI22_X1 U11047 ( .A1(n9927), .A2(n9939), .B1(n6790), .B2(n9926), .ZN(
        P1_U3486) );
  OAI211_X1 U11048 ( .C1(n9906), .C2(n9911), .A(n9905), .B(n9904), .ZN(n9907)
         );
  AOI21_X1 U11049 ( .B1(n9908), .B2(n9914), .A(n9907), .ZN(n9941) );
  AOI22_X1 U11050 ( .A1(n9927), .A2(n9941), .B1(n7156), .B2(n9926), .ZN(
        P1_U3489) );
  OAI211_X1 U11051 ( .C1(n9912), .C2(n9911), .A(n9910), .B(n9909), .ZN(n9913)
         );
  AOI21_X1 U11052 ( .B1(n9915), .B2(n9914), .A(n9913), .ZN(n9942) );
  AOI22_X1 U11053 ( .A1(n9927), .A2(n9942), .B1(n7164), .B2(n9926), .ZN(
        P1_U3492) );
  INV_X1 U11054 ( .A(n9922), .ZN(n9924) );
  AOI211_X1 U11055 ( .C1(n9919), .C2(n9918), .A(n9917), .B(n9916), .ZN(n9920)
         );
  OAI21_X1 U11056 ( .B1(n9922), .B2(n9921), .A(n9920), .ZN(n9923) );
  AOI21_X1 U11057 ( .B1(n9925), .B2(n9924), .A(n9923), .ZN(n9944) );
  AOI22_X1 U11058 ( .A1(n9927), .A2(n9944), .B1(n7265), .B2(n9926), .ZN(
        P1_U3495) );
  AOI22_X1 U11059 ( .A1(n9945), .A2(n9928), .B1(n6489), .B2(n9943), .ZN(
        P1_U3523) );
  AOI22_X1 U11060 ( .A1(n9945), .A2(n9929), .B1(n6492), .B2(n9943), .ZN(
        P1_U3524) );
  AOI22_X1 U11061 ( .A1(n9945), .A2(n9930), .B1(n6494), .B2(n9943), .ZN(
        P1_U3525) );
  AOI22_X1 U11062 ( .A1(n9945), .A2(n9931), .B1(n6496), .B2(n9943), .ZN(
        P1_U3526) );
  AOI22_X1 U11063 ( .A1(n9945), .A2(n9932), .B1(n6419), .B2(n9943), .ZN(
        P1_U3527) );
  AOI22_X1 U11064 ( .A1(n9945), .A2(n9933), .B1(n6533), .B2(n9943), .ZN(
        P1_U3528) );
  AOI22_X1 U11065 ( .A1(n9945), .A2(n9934), .B1(n6578), .B2(n9943), .ZN(
        P1_U3529) );
  INV_X1 U11066 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n9935) );
  AOI22_X1 U11067 ( .A1(n9945), .A2(n9936), .B1(n9935), .B2(n9943), .ZN(
        P1_U3530) );
  AOI22_X1 U11068 ( .A1(n9945), .A2(n9937), .B1(n6670), .B2(n9943), .ZN(
        P1_U3531) );
  AOI22_X1 U11069 ( .A1(n9945), .A2(n9938), .B1(n6710), .B2(n9943), .ZN(
        P1_U3532) );
  AOI22_X1 U11070 ( .A1(n9945), .A2(n9939), .B1(n6783), .B2(n9943), .ZN(
        P1_U3533) );
  AOI22_X1 U11071 ( .A1(n9945), .A2(n9941), .B1(n9940), .B2(n9943), .ZN(
        P1_U3534) );
  AOI22_X1 U11072 ( .A1(n9945), .A2(n9942), .B1(n9096), .B2(n9943), .ZN(
        P1_U3535) );
  AOI22_X1 U11073 ( .A1(n9945), .A2(n9944), .B1(n7260), .B2(n9943), .ZN(
        P1_U3536) );
  AOI22_X1 U11074 ( .A1(P2_ADDR_REG_0__SCAN_IN), .A2(n9946), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3151), .ZN(n9954) );
  MUX2_X1 U11075 ( .A(n9948), .B(n9947), .S(n5537), .Z(n9949) );
  NOR2_X1 U11076 ( .A1(n9949), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n9950) );
  OAI22_X1 U11077 ( .A1(n9952), .A2(n10029), .B1(n9951), .B2(n9950), .ZN(n9953) );
  OAI211_X1 U11078 ( .C1(n9956), .C2(n9955), .A(n9954), .B(n9953), .ZN(
        P2_U3182) );
  INV_X1 U11079 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n9975) );
  OAI21_X1 U11080 ( .B1(n9957), .B2(n9959), .A(n9958), .ZN(n9960) );
  INV_X1 U11081 ( .A(n9960), .ZN(n9968) );
  OAI21_X1 U11082 ( .B1(n9963), .B2(n9962), .A(n9961), .ZN(n9964) );
  NAND2_X1 U11083 ( .A1(n10017), .A2(n9964), .ZN(n9967) );
  AOI22_X1 U11084 ( .A1(n10020), .A2(n9965), .B1(P2_REG3_REG_2__SCAN_IN), .B2(
        P2_U3151), .ZN(n9966) );
  OAI211_X1 U11085 ( .C1(n10024), .C2(n9968), .A(n9967), .B(n9966), .ZN(n9969)
         );
  INV_X1 U11086 ( .A(n9969), .ZN(n9974) );
  XOR2_X1 U11087 ( .A(n9971), .B(n9970), .Z(n9972) );
  NAND2_X1 U11088 ( .A1(n9972), .A2(n10029), .ZN(n9973) );
  OAI211_X1 U11089 ( .C1(n9975), .C2(n10033), .A(n9974), .B(n9973), .ZN(
        P2_U3184) );
  INV_X1 U11090 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n9990) );
  XOR2_X1 U11091 ( .A(n9976), .B(P2_REG1_REG_5__SCAN_IN), .Z(n9980) );
  AOI21_X1 U11092 ( .B1(n9978), .B2(n6406), .A(n9977), .ZN(n9979) );
  OAI22_X1 U11093 ( .A1(n9981), .A2(n9980), .B1(n9979), .B2(n10024), .ZN(n9982) );
  AOI211_X1 U11094 ( .C1(n9984), .C2(n10020), .A(n9983), .B(n9982), .ZN(n9989)
         );
  XOR2_X1 U11095 ( .A(n9986), .B(n9985), .Z(n9987) );
  NAND2_X1 U11096 ( .A1(n9987), .A2(n10029), .ZN(n9988) );
  OAI211_X1 U11097 ( .C1(n9990), .C2(n10033), .A(n9989), .B(n9988), .ZN(
        P2_U3187) );
  INV_X1 U11098 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n10011) );
  NOR2_X1 U11099 ( .A1(n9991), .A2(n9977), .ZN(n9992) );
  NAND2_X1 U11100 ( .A1(n5745), .A2(n9992), .ZN(n9993) );
  AND2_X1 U11101 ( .A1(n9994), .A2(n9993), .ZN(n10003) );
  OAI21_X1 U11102 ( .B1(n9997), .B2(n9996), .A(n9995), .ZN(n9998) );
  NAND2_X1 U11103 ( .A1(n10017), .A2(n9998), .ZN(n10002) );
  AOI21_X1 U11104 ( .B1(n10020), .B2(n10000), .A(n9999), .ZN(n10001) );
  OAI211_X1 U11105 ( .C1(n10024), .C2(n10003), .A(n10002), .B(n10001), .ZN(
        n10004) );
  INV_X1 U11106 ( .A(n10004), .ZN(n10010) );
  OAI21_X1 U11107 ( .B1(n10007), .B2(n10006), .A(n10005), .ZN(n10008) );
  NAND2_X1 U11108 ( .A1(n10008), .A2(n10029), .ZN(n10009) );
  OAI211_X1 U11109 ( .C1(n10011), .C2(n10033), .A(n10010), .B(n10009), .ZN(
        P2_U3188) );
  INV_X1 U11110 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n10034) );
  AOI21_X1 U11111 ( .B1(n10013), .B2(n5814), .A(n10012), .ZN(n10023) );
  OAI21_X1 U11112 ( .B1(n10015), .B2(P2_REG1_REG_7__SCAN_IN), .A(n10014), .ZN(
        n10016) );
  NAND2_X1 U11113 ( .A1(n10017), .A2(n10016), .ZN(n10022) );
  AOI21_X1 U11114 ( .B1(n10020), .B2(n10019), .A(n10018), .ZN(n10021) );
  OAI211_X1 U11115 ( .C1(n10024), .C2(n10023), .A(n10022), .B(n10021), .ZN(
        n10025) );
  INV_X1 U11116 ( .A(n10025), .ZN(n10032) );
  OAI21_X1 U11117 ( .B1(n10028), .B2(n10027), .A(n10026), .ZN(n10030) );
  NAND2_X1 U11118 ( .A1(n10030), .A2(n10029), .ZN(n10031) );
  OAI211_X1 U11119 ( .C1(n10034), .C2(n10033), .A(n10032), .B(n10031), .ZN(
        P2_U3189) );
  XNOR2_X1 U11120 ( .A(n10035), .B(n10039), .ZN(n10059) );
  INV_X1 U11121 ( .A(n10059), .ZN(n10049) );
  OAI22_X1 U11122 ( .A1(n10038), .A2(n10037), .B1(n10058), .B2(n10036), .ZN(
        n10048) );
  XNOR2_X1 U11123 ( .A(n10040), .B(n10039), .ZN(n10045) );
  OAI22_X1 U11124 ( .A1(n5609), .A2(n10043), .B1(n10042), .B2(n10041), .ZN(
        n10044) );
  AOI21_X1 U11125 ( .B1(n10045), .B2(n5513), .A(n10044), .ZN(n10046) );
  OAI21_X1 U11126 ( .B1(n10059), .B2(n10047), .A(n10046), .ZN(n10061) );
  AOI211_X1 U11127 ( .C1(n4426), .C2(n10049), .A(n10048), .B(n10061), .ZN(
        n10051) );
  AOI22_X1 U11128 ( .A1(n8797), .A2(n5085), .B1(n10051), .B2(n10050), .ZN(
        P2_U3231) );
  NAND2_X1 U11129 ( .A1(n10057), .A2(n10052), .ZN(n10053) );
  OAI21_X1 U11130 ( .B1(n10054), .B2(n10103), .A(n10053), .ZN(n10055) );
  AOI211_X1 U11131 ( .C1(n10079), .C2(n10057), .A(n10056), .B(n10055), .ZN(
        n10122) );
  AOI22_X1 U11132 ( .A1(n10120), .A2(n5067), .B1(n10122), .B2(n10118), .ZN(
        P2_U3393) );
  INV_X1 U11133 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n10062) );
  OAI22_X1 U11134 ( .A1(n10059), .A2(n10086), .B1(n10058), .B2(n10103), .ZN(
        n10060) );
  NOR2_X1 U11135 ( .A1(n10061), .A2(n10060), .ZN(n10123) );
  AOI22_X1 U11136 ( .A1(n10120), .A2(n10062), .B1(n10123), .B2(n10118), .ZN(
        P2_U3396) );
  INV_X1 U11137 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n10067) );
  OAI21_X1 U11138 ( .B1(n10064), .B2(n10103), .A(n10063), .ZN(n10065) );
  AOI21_X1 U11139 ( .B1(n10110), .B2(n10066), .A(n10065), .ZN(n10125) );
  AOI22_X1 U11140 ( .A1(n10120), .A2(n10067), .B1(n10125), .B2(n10118), .ZN(
        P2_U3399) );
  INV_X1 U11141 ( .A(n10068), .ZN(n10072) );
  OAI21_X1 U11142 ( .B1(n10070), .B2(n10103), .A(n10069), .ZN(n10071) );
  AOI21_X1 U11143 ( .B1(n10072), .B2(n10110), .A(n10071), .ZN(n10127) );
  AOI22_X1 U11144 ( .A1(n10120), .A2(n5118), .B1(n10127), .B2(n10118), .ZN(
        P2_U3402) );
  INV_X1 U11145 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n10080) );
  INV_X1 U11146 ( .A(n10074), .ZN(n10078) );
  OAI22_X1 U11147 ( .A1(n10074), .A2(n10086), .B1(n10073), .B2(n10103), .ZN(
        n10077) );
  INV_X1 U11148 ( .A(n10075), .ZN(n10076) );
  AOI211_X1 U11149 ( .C1(n10079), .C2(n10078), .A(n10077), .B(n10076), .ZN(
        n10128) );
  AOI22_X1 U11150 ( .A1(n10120), .A2(n10080), .B1(n10128), .B2(n10118), .ZN(
        P2_U3405) );
  AOI22_X1 U11151 ( .A1(n10082), .A2(n10110), .B1(n10112), .B2(n10081), .ZN(
        n10083) );
  AND2_X1 U11152 ( .A1(n10084), .A2(n10083), .ZN(n10129) );
  AOI22_X1 U11153 ( .A1(n10120), .A2(n5152), .B1(n10129), .B2(n10118), .ZN(
        P2_U3408) );
  INV_X1 U11154 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n10090) );
  OAI22_X1 U11155 ( .A1(n10087), .A2(n10086), .B1(n10085), .B2(n10103), .ZN(
        n10088) );
  NOR2_X1 U11156 ( .A1(n10089), .A2(n10088), .ZN(n10130) );
  AOI22_X1 U11157 ( .A1(n10120), .A2(n10090), .B1(n10130), .B2(n10118), .ZN(
        P2_U3411) );
  INV_X1 U11158 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n10097) );
  INV_X1 U11159 ( .A(n10110), .ZN(n10091) );
  OR2_X1 U11160 ( .A1(n10092), .A2(n10091), .ZN(n10095) );
  NAND2_X1 U11161 ( .A1(n10093), .A2(n10112), .ZN(n10094) );
  AND3_X1 U11162 ( .A1(n10096), .A2(n10095), .A3(n10094), .ZN(n10131) );
  AOI22_X1 U11163 ( .A1(n10120), .A2(n10097), .B1(n10131), .B2(n10118), .ZN(
        P2_U3414) );
  INV_X1 U11164 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n10102) );
  AND3_X1 U11165 ( .A1(n10099), .A2(n10110), .A3(n10098), .ZN(n10101) );
  AOI211_X1 U11166 ( .C1(n10112), .C2(n4480), .A(n10101), .B(n10100), .ZN(
        n10132) );
  AOI22_X1 U11167 ( .A1(n10120), .A2(n10102), .B1(n10132), .B2(n10118), .ZN(
        P2_U3417) );
  INV_X1 U11168 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n10108) );
  NOR2_X1 U11169 ( .A1(n10104), .A2(n10103), .ZN(n10106) );
  AOI211_X1 U11170 ( .C1(n10107), .C2(n10110), .A(n10106), .B(n10105), .ZN(
        n10133) );
  AOI22_X1 U11171 ( .A1(n10120), .A2(n10108), .B1(n10133), .B2(n10118), .ZN(
        P2_U3423) );
  INV_X1 U11172 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n10119) );
  NAND3_X1 U11173 ( .A1(n10111), .A2(n10110), .A3(n10109), .ZN(n10115) );
  NAND2_X1 U11174 ( .A1(n10113), .A2(n10112), .ZN(n10114) );
  NAND2_X1 U11175 ( .A1(n10115), .A2(n10114), .ZN(n10116) );
  NOR2_X1 U11176 ( .A1(n10117), .A2(n10116), .ZN(n10134) );
  AOI22_X1 U11177 ( .A1(n10120), .A2(n10119), .B1(n10134), .B2(n10118), .ZN(
        P2_U3426) );
  AOI22_X1 U11178 ( .A1(n10135), .A2(n10122), .B1(n10121), .B2(n5719), .ZN(
        P2_U3460) );
  AOI22_X1 U11179 ( .A1(n10135), .A2(n10123), .B1(n5775), .B2(n5719), .ZN(
        P2_U3461) );
  INV_X1 U11180 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n10124) );
  AOI22_X1 U11181 ( .A1(n10135), .A2(n10125), .B1(n10124), .B2(n5719), .ZN(
        P2_U3462) );
  AOI22_X1 U11182 ( .A1(n10135), .A2(n10127), .B1(n10126), .B2(n5719), .ZN(
        P2_U3463) );
  AOI22_X1 U11183 ( .A1(n10135), .A2(n10128), .B1(n5135), .B2(n5719), .ZN(
        P2_U3464) );
  AOI22_X1 U11184 ( .A1(n10135), .A2(n10129), .B1(n5779), .B2(n5719), .ZN(
        P2_U3465) );
  AOI22_X1 U11185 ( .A1(n10135), .A2(n10130), .B1(n5813), .B2(n5719), .ZN(
        P2_U3466) );
  AOI22_X1 U11186 ( .A1(n10135), .A2(n10131), .B1(n5818), .B2(n5719), .ZN(
        P2_U3467) );
  AOI22_X1 U11187 ( .A1(n10135), .A2(n10132), .B1(n5822), .B2(n5719), .ZN(
        P2_U3468) );
  AOI22_X1 U11188 ( .A1(n10135), .A2(n10133), .B1(n5237), .B2(n5719), .ZN(
        P2_U3470) );
  AOI22_X1 U11189 ( .A1(n10135), .A2(n10134), .B1(n5837), .B2(n5719), .ZN(
        P2_U3471) );
  OAI222_X1 U11190 ( .A1(n10140), .A2(n10139), .B1(n10140), .B2(n10138), .C1(
        n10137), .C2(n10136), .ZN(ADD_1068_U5) );
  XOR2_X1 U11191 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1068_U46) );
  AOI21_X1 U11192 ( .B1(n10143), .B2(n10142), .A(n10141), .ZN(n10144) );
  XOR2_X1 U11193 ( .A(n10144), .B(P2_ADDR_REG_18__SCAN_IN), .Z(ADD_1068_U55)
         );
  OAI21_X1 U11194 ( .B1(n10147), .B2(n10146), .A(n10145), .ZN(ADD_1068_U56) );
  OAI21_X1 U11195 ( .B1(n10150), .B2(n10149), .A(n10148), .ZN(ADD_1068_U57) );
  OAI21_X1 U11196 ( .B1(n10153), .B2(n10152), .A(n10151), .ZN(ADD_1068_U58) );
  OAI21_X1 U11197 ( .B1(n10156), .B2(n10155), .A(n10154), .ZN(ADD_1068_U59) );
  OAI21_X1 U11198 ( .B1(n10159), .B2(n10158), .A(n10157), .ZN(ADD_1068_U60) );
  OAI21_X1 U11199 ( .B1(n10162), .B2(n10161), .A(n10160), .ZN(ADD_1068_U61) );
  OAI21_X1 U11200 ( .B1(n10165), .B2(n10164), .A(n10163), .ZN(ADD_1068_U62) );
  OAI21_X1 U11201 ( .B1(n10168), .B2(n10167), .A(n10166), .ZN(ADD_1068_U63) );
  AOI21_X1 U11202 ( .B1(n10171), .B2(n10170), .A(n10169), .ZN(ADD_1068_U54) );
  OAI21_X1 U11203 ( .B1(n10174), .B2(n10173), .A(n10172), .ZN(ADD_1068_U47) );
  OAI21_X1 U11204 ( .B1(n10177), .B2(n10176), .A(n10175), .ZN(ADD_1068_U48) );
  OAI21_X1 U11205 ( .B1(n10180), .B2(n10179), .A(n10178), .ZN(ADD_1068_U49) );
  OAI21_X1 U11206 ( .B1(n10183), .B2(n10182), .A(n10181), .ZN(ADD_1068_U50) );
  OAI21_X1 U11207 ( .B1(n10186), .B2(n10185), .A(n10184), .ZN(ADD_1068_U51) );
  AOI21_X1 U11208 ( .B1(n10189), .B2(n10188), .A(n10187), .ZN(ADD_1068_U53) );
  OAI21_X1 U11209 ( .B1(n10192), .B2(n10191), .A(n10190), .ZN(ADD_1068_U52) );
  AND2_X1 U4860 ( .A1(n9476), .A2(n9475), .ZN(n10196) );
endmodule

