

module b14_C_AntiSAT_k_256_10 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, 
        REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, 
        REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, 
        REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, 
        REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, 
        REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, 
        REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, 
        REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, 
        IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, 
        IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, 
        IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, 
        IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, 
        IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, 
        IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, 
        IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, 
        IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, 
        IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, 
        IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, 
        IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, 
        D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, 
        D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, 
        D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, 
        D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, 
        D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, 
        D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, 
        D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, 
        D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, 
        D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, 
        D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, 
        REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, 
        REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, 
        REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, 
        REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, 
        REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, 
        REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, 
        REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, 
        REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, 
        REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, 
        REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, 
        REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, 
        REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, 
        REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, 
        REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, 
        REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, 
        REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, 
        REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, 
        REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, 
        REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, 
        REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, 
        REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, 
        REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, 
        REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, 
        REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, 
        REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, 
        REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, 
        REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, 
        REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, 
        REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, 
        REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, 
        REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, 
        REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, 
        ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, 
        ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, 
        ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, 
        ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, 
        ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, 
        ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, 
        ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, 
        REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, 
        REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, 
        keyinput128, keyinput129, keyinput130, keyinput131, keyinput132, 
        keyinput133, keyinput134, keyinput135, keyinput136, keyinput137, 
        keyinput138, keyinput139, keyinput140, keyinput141, keyinput142, 
        keyinput143, keyinput144, keyinput145, keyinput146, keyinput147, 
        keyinput148, keyinput149, keyinput150, keyinput151, keyinput152, 
        keyinput153, keyinput154, keyinput155, keyinput156, keyinput157, 
        keyinput158, keyinput159, keyinput160, keyinput161, keyinput162, 
        keyinput163, keyinput164, keyinput165, keyinput166, keyinput167, 
        keyinput168, keyinput169, keyinput170, keyinput171, keyinput172, 
        keyinput173, keyinput174, keyinput175, keyinput176, keyinput177, 
        keyinput178, keyinput179, keyinput180, keyinput181, keyinput182, 
        keyinput183, keyinput184, keyinput185, keyinput186, keyinput187, 
        keyinput188, keyinput189, keyinput190, keyinput191, keyinput192, 
        keyinput193, keyinput194, keyinput195, keyinput196, keyinput197, 
        keyinput198, keyinput199, keyinput200, keyinput201, keyinput202, 
        keyinput203, keyinput204, keyinput205, keyinput206, keyinput207, 
        keyinput208, keyinput209, keyinput210, keyinput211, keyinput212, 
        keyinput213, keyinput214, keyinput215, keyinput216, keyinput217, 
        keyinput218, keyinput219, keyinput220, keyinput221, keyinput222, 
        keyinput223, keyinput224, keyinput225, keyinput226, keyinput227, 
        keyinput228, keyinput229, keyinput230, keyinput231, keyinput232, 
        keyinput233, keyinput234, keyinput235, keyinput236, keyinput237, 
        keyinput238, keyinput239, keyinput240, keyinput241, keyinput242, 
        keyinput243, keyinput244, keyinput245, keyinput246, keyinput247, 
        keyinput248, keyinput249, keyinput250, keyinput251, keyinput252, 
        keyinput253, keyinput254, keyinput255, U3352, U3351, U3350, U3349, 
        U3348, U3347, U3346, U3345, U3344, U3343, U3342, U3341, U3340, U3339, 
        U3338, U3337, U3336, U3335, U3334, U3333, U3332, U3331, U3330, U3329, 
        U3328, U3327, U3326, U3325, U3324, U3323, U3322, U3321, U3458, U3459, 
        U3320, U3319, U3318, U3317, U3316, U3315, U3314, U3313, U3312, U3311, 
        U3310, U3309, U3308, U3307, U3306, U3305, U3304, U3303, U3302, U3301, 
        U3300, U3299, U3298, U3297, U3296, U3295, U3294, U3293, U3292, U3291, 
        U3467, U3469, U3471, U3473, U3475, U3477, U3479, U3481, U3483, U3485, 
        U3487, U3489, U3491, U3493, U3495, U3497, U3499, U3501, U3503, U3505, 
        U3506, U3507, U3508, U3509, U3510, U3511, U3512, U3513, U3514, U3515, 
        U3516, U3517, U3518, U3519, U3520, U3521, U3522, U3523, U3524, U3525, 
        U3526, U3527, U3528, U3529, U3530, U3531, U3532, U3533, U3534, U3535, 
        U3536, U3537, U3538, U3539, U3540, U3541, U3542, U3543, U3544, U3545, 
        U3546, U3547, U3548, U3549, U3290, U3289, U3288, U3287, U3286, U3285, 
        U3284, U3283, U3282, U3281, U3280, U3279, U3278, U3277, U3276, U3275, 
        U3274, U3273, U3272, U3271, U3270, U3269, U3268, U3267, U3266, U3265, 
        U3264, U3263, U3262, U3354, U3261, U3260, U3259, U3258, U3257, U3256, 
        U3255, U3254, U3253, U3252, U3251, U3250, U3249, U3248, U3247, U3246, 
        U3245, U3244, U3243, U3242, U3241, U3240, U3550, U3551, U3552, U3553, 
        U3554, U3555, U3556, U3557, U3558, U3559, U3560, U3561, U3562, U3563, 
        U3564, U3565, U3566, U3567, U3568, U3569, U3570, U3571, U3572, U3573, 
        U3574, U3575, U3576, U3577, U3578, U3579, U3580, U3581, U3239, U3238, 
        U3237, U3236, U3235, U3234, U3233, U3232, U3231, U3230, U3229, U3228, 
        U3227, U3226, U3225, U3224, U3223, U3222, U3221, U3220, U3219, U3218, 
        U3217, U3216, U3215, U3214, U3213, U3212, U3211, U3210, U3149, U3148, 
        U4043 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
         REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
         REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
         REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
         REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
         REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
         REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
         REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
         IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
         IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
         IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
         IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
         IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
         IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
         IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
         IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
         IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
         IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
         IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
         D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
         D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN,
         D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
         D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
         D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
         D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
         D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
         D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
         D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
         D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
         D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
         REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
         REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
         REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
         REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
         REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
         REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
         REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
         REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
         REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
         REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
         REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
         REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
         REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
         REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
         REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
         REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
         REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
         REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
         REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
         REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
         REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
         REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
         REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
         REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
         REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
         REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
         REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
         REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
         REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
         REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
         REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
         REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
         ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
         ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
         ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
         ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
         ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
         ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
         DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
         DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
         DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
         DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
         DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
         DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
         DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
         DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
         DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
         DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
         DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
         REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
         REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
         REG3_REG_22__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127, keyinput128, keyinput129,
         keyinput130, keyinput131, keyinput132, keyinput133, keyinput134,
         keyinput135, keyinput136, keyinput137, keyinput138, keyinput139,
         keyinput140, keyinput141, keyinput142, keyinput143, keyinput144,
         keyinput145, keyinput146, keyinput147, keyinput148, keyinput149,
         keyinput150, keyinput151, keyinput152, keyinput153, keyinput154,
         keyinput155, keyinput156, keyinput157, keyinput158, keyinput159,
         keyinput160, keyinput161, keyinput162, keyinput163, keyinput164,
         keyinput165, keyinput166, keyinput167, keyinput168, keyinput169,
         keyinput170, keyinput171, keyinput172, keyinput173, keyinput174,
         keyinput175, keyinput176, keyinput177, keyinput178, keyinput179,
         keyinput180, keyinput181, keyinput182, keyinput183, keyinput184,
         keyinput185, keyinput186, keyinput187, keyinput188, keyinput189,
         keyinput190, keyinput191, keyinput192, keyinput193, keyinput194,
         keyinput195, keyinput196, keyinput197, keyinput198, keyinput199,
         keyinput200, keyinput201, keyinput202, keyinput203, keyinput204,
         keyinput205, keyinput206, keyinput207, keyinput208, keyinput209,
         keyinput210, keyinput211, keyinput212, keyinput213, keyinput214,
         keyinput215, keyinput216, keyinput217, keyinput218, keyinput219,
         keyinput220, keyinput221, keyinput222, keyinput223, keyinput224,
         keyinput225, keyinput226, keyinput227, keyinput228, keyinput229,
         keyinput230, keyinput231, keyinput232, keyinput233, keyinput234,
         keyinput235, keyinput236, keyinput237, keyinput238, keyinput239,
         keyinput240, keyinput241, keyinput242, keyinput243, keyinput244,
         keyinput245, keyinput246, keyinput247, keyinput248, keyinput249,
         keyinput250, keyinput251, keyinput252, keyinput253, keyinput254,
         keyinput255;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244,
         n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254,
         n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264,
         n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274,
         n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284,
         n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294,
         n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304,
         n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314,
         n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324,
         n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334,
         n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344,
         n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354,
         n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364,
         n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374,
         n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384,
         n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394,
         n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404,
         n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414,
         n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424,
         n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434,
         n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444,
         n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454,
         n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464,
         n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474,
         n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484,
         n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494,
         n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504,
         n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514,
         n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524,
         n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534,
         n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544,
         n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554,
         n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564,
         n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574,
         n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584,
         n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594,
         n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604,
         n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614,
         n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624,
         n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634,
         n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644,
         n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654,
         n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664,
         n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674,
         n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684,
         n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694,
         n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704,
         n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714,
         n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724,
         n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734,
         n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744,
         n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754,
         n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764,
         n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774,
         n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784,
         n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794,
         n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804,
         n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814,
         n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824,
         n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834,
         n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844,
         n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854,
         n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864,
         n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874,
         n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884,
         n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894,
         n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904,
         n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914,
         n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924,
         n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934,
         n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944,
         n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954,
         n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964,
         n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974,
         n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984,
         n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994,
         n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004,
         n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014,
         n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024,
         n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034,
         n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044,
         n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054,
         n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064,
         n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074,
         n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084,
         n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094,
         n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104,
         n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114,
         n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124,
         n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134,
         n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144,
         n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154,
         n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164,
         n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174,
         n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184,
         n3185, n3186, n3187, n3188, n3189, n3191, n3192, n3193, n3194, n3195,
         n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205,
         n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215,
         n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225,
         n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235,
         n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245,
         n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255,
         n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265,
         n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275,
         n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285,
         n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295,
         n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305,
         n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315,
         n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325,
         n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335,
         n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345,
         n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355,
         n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365,
         n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375,
         n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385,
         n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395,
         n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405,
         n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415,
         n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425,
         n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435,
         n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445,
         n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455,
         n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465,
         n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475,
         n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485,
         n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495,
         n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505,
         n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515,
         n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525,
         n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535,
         n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545,
         n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555,
         n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565,
         n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575,
         n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585,
         n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595,
         n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605,
         n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615,
         n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625,
         n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635,
         n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645,
         n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655,
         n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665,
         n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675,
         n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685,
         n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695,
         n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705,
         n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715,
         n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725,
         n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735,
         n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745,
         n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755,
         n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765,
         n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775,
         n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785,
         n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795,
         n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805,
         n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815,
         n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825,
         n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835,
         n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845,
         n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855,
         n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865,
         n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875,
         n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885,
         n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895,
         n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905,
         n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915,
         n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925,
         n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935,
         n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945,
         n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955,
         n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965,
         n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975,
         n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985,
         n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995,
         n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005,
         n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015,
         n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025,
         n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035,
         n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045,
         n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055,
         n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065,
         n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075,
         n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085,
         n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095,
         n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105,
         n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115,
         n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125,
         n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135,
         n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145,
         n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155,
         n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165,
         n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175,
         n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185,
         n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195,
         n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205,
         n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215,
         n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226,
         n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236,
         n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246,
         n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256,
         n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266,
         n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276,
         n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286,
         n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296,
         n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306,
         n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316,
         n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326,
         n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336,
         n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346,
         n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356,
         n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366,
         n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376,
         n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386,
         n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396,
         n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406,
         n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416,
         n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426,
         n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436,
         n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446,
         n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456,
         n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466,
         n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476,
         n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486,
         n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496,
         n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506,
         n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516,
         n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526,
         n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536,
         n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546,
         n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556,
         n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566,
         n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576,
         n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586,
         n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596,
         n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606,
         n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616,
         n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626,
         n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636,
         n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646,
         n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656,
         n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666,
         n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676,
         n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686,
         n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696,
         n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706,
         n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716,
         n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726,
         n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736,
         n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746,
         n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756,
         n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766,
         n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776,
         n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786,
         n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796,
         n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806,
         n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816,
         n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826,
         n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836,
         n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846,
         n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856,
         n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866,
         n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876,
         n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886,
         n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896,
         n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906,
         n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916,
         n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926,
         n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936,
         n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946,
         n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956,
         n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966,
         n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976,
         n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986,
         n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996,
         n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006,
         n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016,
         n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026,
         n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036,
         n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046,
         n5047, n5048, n5049, n5050, n5051, n5052;

  BUF_X4 U2477 ( .A(n2571), .Z(n2951) );
  INV_X4 U2478 ( .A(n2947), .ZN(n2920) );
  INV_X1 U2479 ( .A(n2944), .ZN(n2571) );
  INV_X1 U2481 ( .A(n2601), .ZN(n2563) );
  XNOR2_X1 U2482 ( .A(n2486), .B(n3108), .ZN(n2488) );
  NOR2_X2 U2483 ( .A1(IR_REG_1__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n2590)
         );
  INV_X1 U2484 ( .A(n2684), .ZN(n3230) );
  XNOR2_X1 U2485 ( .A(n2325), .B(n2324), .ZN(n2490) );
  XNOR2_X1 U2486 ( .A(n2554), .B(IR_REG_1__SCAN_IN), .ZN(n3143) );
  AOI21_X2 U2487 ( .B1(n3391), .B2(n2455), .A(n2453), .ZN(n3486) );
  OR2_X2 U2488 ( .A1(n4306), .A2(n3094), .ZN(n4172) );
  OAI22_X2 U2489 ( .A1(n3213), .A2(n3021), .B1(n3266), .B2(n3173), .ZN(n3192)
         );
  NAND2_X1 U2490 ( .A1(n2544), .A2(n3051), .ZN(n2944) );
  NAND2_X1 U2491 ( .A1(n2360), .A2(n2358), .ZN(n3965) );
  AND2_X1 U2492 ( .A1(n3728), .A2(n4403), .ZN(n2796) );
  AOI21_X1 U2493 ( .B1(n4086), .B2(n3044), .A(n2468), .ZN(n4070) );
  NAND2_X1 U2494 ( .A1(n2354), .A2(n2353), .ZN(n4165) );
  AOI21_X1 U2495 ( .B1(n3447), .B2(n3446), .A(n2465), .ZN(n3476) );
  AND2_X1 U2496 ( .A1(n3757), .A2(n2332), .ZN(n2331) );
  NOR2_X1 U2497 ( .A1(n2581), .A2(n2466), .ZN(n3162) );
  NAND2_X1 U2498 ( .A1(n4225), .A2(n4224), .ZN(n2326) );
  INV_X2 U2499 ( .A(n4577), .ZN(n4213) );
  NAND2_X1 U2500 ( .A1(n2972), .A2(n3848), .ZN(n4638) );
  OR2_X1 U2501 ( .A1(n2542), .A2(n3762), .ZN(n2535) );
  NOR2_X1 U2502 ( .A1(n2258), .A2(n2239), .ZN(n3136) );
  NAND2_X1 U2503 ( .A1(n2531), .A2(n2534), .ZN(n3959) );
  NAND2_X1 U2504 ( .A1(n2531), .A2(IR_REG_31__SCAN_IN), .ZN(n2515) );
  NAND2_X1 U2505 ( .A1(n2248), .A2(n2526), .ZN(n3137) );
  XNOR2_X1 U2506 ( .A(n2530), .B(n2529), .ZN(n3897) );
  NAND2_X1 U2507 ( .A1(n2533), .A2(n2532), .ZN(n2531) );
  OR2_X1 U2508 ( .A1(n2999), .A2(n2743), .ZN(n2325) );
  NAND2_X1 U2509 ( .A1(n2247), .A2(IR_REG_31__SCAN_IN), .ZN(n2533) );
  INV_X1 U2510 ( .A(n2508), .ZN(n2483) );
  AND2_X1 U2511 ( .A1(n2481), .A2(n2480), .ZN(n2482) );
  AND2_X1 U2512 ( .A1(n2474), .A2(n2475), .ZN(n2460) );
  AND4_X1 U2513 ( .A1(n2478), .A2(n2970), .A3(n2529), .A4(n2477), .ZN(n2481)
         );
  NOR2_X1 U2514 ( .A1(IR_REG_3__SCAN_IN), .A2(IR_REG_2__SCAN_IN), .ZN(n2470)
         );
  INV_X1 U2515 ( .A(IR_REG_4__SCAN_IN), .ZN(n4896) );
  INV_X1 U2516 ( .A(IR_REG_15__SCAN_IN), .ZN(n2786) );
  NOR2_X1 U2517 ( .A1(IR_REG_12__SCAN_IN), .A2(IR_REG_11__SCAN_IN), .ZN(n2474)
         );
  INV_X1 U2518 ( .A(IR_REG_23__SCAN_IN), .ZN(n2970) );
  NOR2_X1 U2519 ( .A1(IR_REG_26__SCAN_IN), .A2(IR_REG_25__SCAN_IN), .ZN(n2499)
         );
  INV_X1 U2520 ( .A(IR_REG_8__SCAN_IN), .ZN(n2695) );
  AOI21_X2 U2521 ( .B1(n2263), .B2(n2736), .A(n2735), .ZN(n3552) );
  NAND2_X4 U2522 ( .A1(n2488), .A2(n4376), .ZN(n2601) );
  AOI21_X1 U2523 ( .B1(n2366), .B2(n2364), .A(n2266), .ZN(n2363) );
  INV_X1 U2524 ( .A(n2261), .ZN(n2364) );
  NAND2_X1 U2525 ( .A1(n3136), .A2(IR_REG_28__SCAN_IN), .ZN(n2370) );
  NAND2_X1 U2526 ( .A1(n3137), .A2(n2527), .ZN(n2371) );
  AND2_X1 U2527 ( .A1(n3605), .A2(n3754), .ZN(n3878) );
  NAND2_X1 U2528 ( .A1(n3336), .A2(n3277), .ZN(n2351) );
  NAND2_X1 U2529 ( .A1(n2394), .A2(n2393), .ZN(n2392) );
  NAND2_X1 U2530 ( .A1(n2401), .A2(n4432), .ZN(n2393) );
  NAND2_X1 U2531 ( .A1(n2402), .A2(n3134), .ZN(n2394) );
  NAND2_X1 U2532 ( .A1(n4488), .A2(n2464), .ZN(n3944) );
  OR2_X1 U2533 ( .A1(n4494), .A2(n3932), .ZN(n3934) );
  INV_X1 U2534 ( .A(n3048), .ZN(n2367) );
  NOR2_X1 U2535 ( .A1(n3534), .A2(n3533), .ZN(n3568) );
  INV_X1 U2536 ( .A(IR_REG_21__SCAN_IN), .ZN(n2518) );
  NOR2_X1 U2537 ( .A1(n2508), .A2(n2509), .ZN(n2519) );
  OR2_X1 U2538 ( .A1(IR_REG_18__SCAN_IN), .A2(n2252), .ZN(n2509) );
  INV_X1 U2539 ( .A(IR_REG_13__SCAN_IN), .ZN(n2475) );
  INV_X1 U2540 ( .A(IR_REG_9__SCAN_IN), .ZN(n2471) );
  INV_X1 U2541 ( .A(IR_REG_5__SCAN_IN), .ZN(n2472) );
  NAND2_X1 U2542 ( .A1(n2434), .A2(n2432), .ZN(n3635) );
  AOI21_X1 U2543 ( .B1(n2235), .B2(n2244), .A(n2433), .ZN(n2432) );
  INV_X1 U2544 ( .A(n3707), .ZN(n2433) );
  AOI21_X1 U2545 ( .B1(n3018), .B2(n2795), .A(n2555), .ZN(n2560) );
  INV_X1 U2546 ( .A(n2566), .ZN(n2991) );
  INV_X1 U2547 ( .A(n2564), .ZN(n2684) );
  NAND2_X1 U2548 ( .A1(n3107), .A2(IR_REG_31__SCAN_IN), .ZN(n2486) );
  INV_X1 U2549 ( .A(n2363), .ZN(n2362) );
  NAND2_X1 U2550 ( .A1(n2302), .A2(n2305), .ZN(n2301) );
  INV_X1 U2551 ( .A(n3874), .ZN(n2302) );
  AND2_X1 U2552 ( .A1(n2715), .A2(n3455), .ZN(n2455) );
  XNOR2_X1 U2553 ( .A(n2597), .B(n2947), .ZN(n2598) );
  OAI21_X1 U2554 ( .B1(n2719), .B2(n2454), .A(n2278), .ZN(n2453) );
  INV_X1 U2555 ( .A(n3455), .ZN(n2454) );
  INV_X1 U2556 ( .A(n3484), .ZN(n2452) );
  NAND2_X1 U2557 ( .A1(n3391), .A2(n2451), .ZN(n2450) );
  AND2_X1 U2558 ( .A1(n2455), .A2(n2452), .ZN(n2451) );
  INV_X1 U2559 ( .A(n2420), .ZN(n3132) );
  NOR2_X1 U2560 ( .A1(n3600), .A2(n2362), .ZN(n2361) );
  NOR3_X1 U2561 ( .A1(n3600), .A2(n2362), .A3(n2366), .ZN(n2359) );
  AND2_X1 U2562 ( .A1(n2306), .A2(n3781), .ZN(n2305) );
  NAND2_X1 U2563 ( .A1(n4030), .A2(n3874), .ZN(n2307) );
  NAND2_X1 U2564 ( .A1(n2311), .A2(n2309), .ZN(n4106) );
  NOR2_X1 U2565 ( .A1(n3862), .A2(n2310), .ZN(n2309) );
  INV_X1 U2566 ( .A(n2313), .ZN(n2310) );
  NAND2_X1 U2567 ( .A1(n2295), .A2(n3828), .ZN(n4205) );
  NAND2_X1 U2568 ( .A1(n3471), .A2(n3826), .ZN(n2295) );
  INV_X1 U2569 ( .A(n2341), .ZN(n2339) );
  NAND2_X1 U2570 ( .A1(n2262), .A2(n2338), .ZN(n2337) );
  INV_X1 U2571 ( .A(n3026), .ZN(n2338) );
  OR2_X1 U2572 ( .A1(n3905), .A2(n3420), .ZN(n3822) );
  NAND2_X1 U2573 ( .A1(n2255), .A2(n2351), .ZN(n2346) );
  AND2_X1 U2574 ( .A1(n3193), .A2(n2351), .ZN(n2348) );
  NOR2_X1 U2575 ( .A1(n2542), .A2(n3762), .ZN(n3051) );
  OR2_X1 U2576 ( .A1(n2576), .A2(n4232), .ZN(n3788) );
  OR2_X1 U2577 ( .A1(n3018), .A2(n3253), .ZN(n3787) );
  INV_X1 U2578 ( .A(n3036), .ZN(n2356) );
  AND2_X1 U2579 ( .A1(n3762), .A2(n3897), .ZN(n2972) );
  OR2_X1 U2580 ( .A1(n2484), .A2(IR_REG_27__SCAN_IN), .ZN(n2485) );
  AND3_X1 U2581 ( .A1(n2532), .A2(n2479), .A3(n2518), .ZN(n2480) );
  AND2_X1 U2582 ( .A1(n3410), .A2(n3408), .ZN(n2715) );
  INV_X1 U2583 ( .A(n3715), .ZN(n2444) );
  NAND2_X1 U2584 ( .A1(n2425), .A2(n2424), .ZN(n3354) );
  AOI21_X1 U2585 ( .B1(n2426), .B2(n2429), .A(n2249), .ZN(n2424) );
  INV_X1 U2586 ( .A(n2572), .ZN(n3741) );
  NAND2_X1 U2587 ( .A1(n2800), .A2(n2799), .ZN(n2801) );
  INV_X1 U2588 ( .A(n2798), .ZN(n2800) );
  NAND2_X1 U2589 ( .A1(n3627), .A2(n2898), .ZN(n3674) );
  AND2_X1 U2590 ( .A1(n2897), .A2(n2896), .ZN(n2898) );
  NAND2_X1 U2591 ( .A1(n2842), .A2(n2841), .ZN(n2843) );
  INV_X1 U2592 ( .A(n2840), .ZN(n2842) );
  NAND2_X1 U2593 ( .A1(n3686), .A2(n2457), .ZN(n2456) );
  NOR2_X1 U2594 ( .A1(n3642), .A2(n2458), .ZN(n2457) );
  NAND2_X1 U2595 ( .A1(n2716), .A2(n2718), .ZN(n2719) );
  INV_X1 U2596 ( .A(n2717), .ZN(n2718) );
  XNOR2_X1 U2597 ( .A(n2575), .B(n2947), .ZN(n2580) );
  OR2_X1 U2598 ( .A1(n2797), .A2(n2235), .ZN(n2435) );
  NAND2_X1 U2599 ( .A1(n2264), .A2(n2443), .ZN(n2445) );
  INV_X1 U2600 ( .A(n2584), .ZN(n2996) );
  NOR2_X1 U2601 ( .A1(n2507), .A2(n3106), .ZN(n2514) );
  NAND2_X1 U2602 ( .A1(n5041), .A2(n3131), .ZN(n3912) );
  NAND2_X1 U2603 ( .A1(n3913), .A2(n3912), .ZN(n3911) );
  NAND2_X1 U2604 ( .A1(n2283), .A2(n2282), .ZN(n3510) );
  NAND2_X1 U2605 ( .A1(n4382), .A2(REG2_REG_5__SCAN_IN), .ZN(n2282) );
  NAND2_X1 U2606 ( .A1(n3508), .A2(n2284), .ZN(n2283) );
  NAND2_X1 U2607 ( .A1(n3509), .A2(n3129), .ZN(n2284) );
  OAI211_X1 U2608 ( .C1(n3147), .C2(n2396), .A(n2395), .B(n2391), .ZN(n3496)
         );
  NAND2_X1 U2609 ( .A1(n4382), .A2(REG1_REG_5__SCAN_IN), .ZN(n2395) );
  NAND2_X1 U2610 ( .A1(n2402), .A2(n4432), .ZN(n2396) );
  NAND2_X1 U2611 ( .A1(n4451), .A2(n3512), .ZN(n3514) );
  OAI22_X1 U2612 ( .A1(n4447), .A2(n3498), .B1(REG1_REG_7__SCAN_IN), .B2(n4445), .ZN(n3500) );
  AND2_X1 U2613 ( .A1(n4445), .A2(REG1_REG_7__SCAN_IN), .ZN(n3498) );
  NOR2_X1 U2614 ( .A1(n4464), .A2(n2412), .ZN(n3503) );
  AND2_X1 U2615 ( .A1(n3507), .A2(REG1_REG_9__SCAN_IN), .ZN(n2412) );
  OR2_X1 U2616 ( .A1(n4475), .A2(n4476), .ZN(n2410) );
  NAND2_X1 U2617 ( .A1(n2291), .A2(n3947), .ZN(n3948) );
  OR2_X1 U2618 ( .A1(n4509), .A2(n2407), .ZN(n2405) );
  NAND2_X1 U2619 ( .A1(n2409), .A2(REG1_REG_14__SCAN_IN), .ZN(n2407) );
  NAND2_X1 U2620 ( .A1(n3935), .A2(n2409), .ZN(n2406) );
  OR2_X1 U2621 ( .A1(n4509), .A2(n4508), .ZN(n2408) );
  NAND2_X1 U2622 ( .A1(n4537), .A2(n2385), .ZN(n4550) );
  NAND2_X1 U2623 ( .A1(n4586), .A2(n4304), .ZN(n2385) );
  NAND2_X1 U2624 ( .A1(n4540), .A2(n2290), .ZN(n4553) );
  OR2_X1 U2625 ( .A1(n3954), .A2(REG2_REG_17__SCAN_IN), .ZN(n2290) );
  OR2_X1 U2626 ( .A1(n2902), .A2(n2901), .ZN(n2914) );
  NAND2_X1 U2627 ( .A1(n2357), .A2(n2363), .ZN(n4011) );
  OR2_X1 U2628 ( .A1(n4045), .A2(n2365), .ZN(n2357) );
  OR2_X1 U2629 ( .A1(n4146), .A2(n4138), .ZN(n3040) );
  AOI22_X1 U2630 ( .A1(n3476), .A2(n3030), .B1(n3029), .B2(n3543), .ZN(n3534)
         );
  OR2_X1 U2631 ( .A1(n3905), .A2(n3425), .ZN(n3027) );
  NAND2_X1 U2632 ( .A1(n3424), .A2(n2265), .ZN(n3028) );
  OR2_X1 U2633 ( .A1(n2701), .A2(n3412), .ZN(n2721) );
  NAND2_X1 U2634 ( .A1(n3394), .A2(n3367), .ZN(n2341) );
  OAI21_X1 U2635 ( .B1(n3194), .B2(n3056), .A(n3798), .ZN(n3319) );
  NAND2_X1 U2636 ( .A1(n2326), .A2(n3020), .ZN(n3213) );
  AND2_X1 U2637 ( .A1(n3240), .A2(n3019), .ZN(n4225) );
  AND2_X1 U2638 ( .A1(n3750), .A2(n3236), .ZN(n3241) );
  NOR2_X1 U2639 ( .A1(n4060), .A2(n2376), .ZN(n4019) );
  AND2_X1 U2640 ( .A1(n4226), .A2(n4614), .ZN(n4605) );
  NAND2_X1 U2641 ( .A1(n4378), .A2(n2956), .ZN(n3113) );
  NOR2_X1 U2642 ( .A1(IR_REG_26__SCAN_IN), .A2(IR_REG_31__SCAN_IN), .ZN(n2500)
         );
  NAND2_X1 U2643 ( .A1(n2511), .A2(IR_REG_31__SCAN_IN), .ZN(n2971) );
  AND2_X1 U2644 ( .A1(n2518), .A2(n2529), .ZN(n2510) );
  XNOR2_X1 U2645 ( .A(n2971), .B(n2970), .ZN(n3120) );
  NOR2_X1 U2646 ( .A1(IR_REG_10__SCAN_IN), .A2(IR_REG_17__SCAN_IN), .ZN(n2297)
         );
  NOR3_X1 U2647 ( .A1(n2473), .A2(n2624), .A3(IR_REG_10__SCAN_IN), .ZN(n2521)
         );
  INV_X1 U2648 ( .A(IR_REG_3__SCAN_IN), .ZN(n2592) );
  NAND2_X1 U2649 ( .A1(n3391), .A2(n2715), .ZN(n3409) );
  INV_X1 U2650 ( .A(n4112), .ZN(n4146) );
  OR3_X1 U2651 ( .A1(n2879), .A2(n2878), .A3(n2877), .ZN(n4072) );
  NAND4_X1 U2652 ( .A1(n2605), .A2(n2604), .A3(n2603), .A4(n2602), .ZN(n3909)
         );
  OR2_X1 U2653 ( .A1(n2584), .A2(n3273), .ZN(n2603) );
  XNOR2_X1 U2654 ( .A(n3510), .B(n4598), .ZN(n4439) );
  NAND2_X1 U2655 ( .A1(n4439), .A2(REG2_REG_6__SCAN_IN), .ZN(n4438) );
  NAND2_X1 U2656 ( .A1(n4452), .A2(n4453), .ZN(n4451) );
  XNOR2_X1 U2657 ( .A(n3514), .B(n3499), .ZN(n4461) );
  XNOR2_X1 U2658 ( .A(n3503), .B(n2411), .ZN(n4475) );
  OAI21_X1 U2659 ( .B1(n4560), .B2(n4950), .A(n4559), .ZN(n2414) );
  NAND2_X1 U2660 ( .A1(n2384), .A2(n2383), .ZN(n4558) );
  INV_X1 U2661 ( .A(n4549), .ZN(n2383) );
  INV_X1 U2662 ( .A(n4550), .ZN(n2384) );
  AOI21_X1 U2663 ( .B1(n4553), .B2(n4552), .A(n4551), .ZN(n2415) );
  OAI21_X1 U2664 ( .B1(n2319), .B2(n4236), .A(n2318), .ZN(n4259) );
  AND2_X1 U2665 ( .A1(n3608), .A2(n3609), .ZN(n2318) );
  XNOR2_X1 U2666 ( .A(n3607), .B(n3778), .ZN(n2319) );
  OR2_X1 U2667 ( .A1(n3071), .A2(n4125), .ZN(n3862) );
  INV_X1 U2668 ( .A(IR_REG_24__SCAN_IN), .ZN(n2477) );
  INV_X1 U2669 ( .A(IR_REG_20__SCAN_IN), .ZN(n2478) );
  NAND2_X1 U2670 ( .A1(n2237), .A2(n3284), .ZN(n2429) );
  NOR2_X1 U2671 ( .A1(n3148), .A2(n2403), .ZN(n2402) );
  OR2_X1 U2672 ( .A1(n2294), .A2(n3519), .ZN(n2293) );
  INV_X1 U2673 ( .A(n4522), .ZN(n2409) );
  OAI21_X1 U2674 ( .B1(n4030), .B2(n2300), .A(n2299), .ZN(n3992) );
  NAND2_X1 U2675 ( .A1(n2308), .A2(n3872), .ZN(n2300) );
  NAND2_X1 U2676 ( .A1(n2256), .A2(n2308), .ZN(n2299) );
  NOR2_X1 U2677 ( .A1(n2334), .A2(n2329), .ZN(n2328) );
  INV_X1 U2678 ( .A(n3039), .ZN(n2329) );
  INV_X1 U2679 ( .A(n3041), .ZN(n2334) );
  NAND2_X1 U2680 ( .A1(n2333), .A2(n3041), .ZN(n2332) );
  INV_X1 U2681 ( .A(n3040), .ZN(n2333) );
  AND2_X1 U2682 ( .A1(n4105), .A2(n3075), .ZN(n3867) );
  AOI21_X1 U2683 ( .B1(n4182), .B2(n2315), .A(n2314), .ZN(n2313) );
  INV_X1 U2684 ( .A(n3812), .ZN(n2315) );
  NAND2_X1 U2685 ( .A1(n2312), .A2(n4182), .ZN(n2311) );
  OR2_X1 U2686 ( .A1(n3904), .A2(n4201), .ZN(n3830) );
  NAND2_X1 U2687 ( .A1(n4205), .A2(n4206), .ZN(n4204) );
  NAND2_X1 U2688 ( .A1(n3362), .A2(n3806), .ZN(n2322) );
  INV_X1 U2689 ( .A(n3082), .ZN(n3121) );
  NAND2_X1 U2690 ( .A1(n2375), .A2(n3721), .ZN(n2374) );
  INV_X1 U2691 ( .A(n2376), .ZN(n2375) );
  NAND2_X1 U2692 ( .A1(n3679), .A2(n4021), .ZN(n2376) );
  NAND2_X1 U2693 ( .A1(n2379), .A2(n4114), .ZN(n2378) );
  INV_X1 U2694 ( .A(n2380), .ZN(n2379) );
  NAND2_X1 U2695 ( .A1(n4145), .A2(n4138), .ZN(n2380) );
  INV_X1 U2696 ( .A(IR_REG_7__SCAN_IN), .ZN(n2659) );
  INV_X1 U2697 ( .A(n3285), .ZN(n2431) );
  AND2_X1 U2698 ( .A1(n2431), .A2(n3308), .ZN(n2426) );
  NAND2_X1 U2699 ( .A1(n2430), .A2(n2428), .ZN(n2427) );
  INV_X1 U2700 ( .A(n2429), .ZN(n2428) );
  INV_X1 U2701 ( .A(DATAI_1_), .ZN(n2373) );
  INV_X1 U2702 ( .A(n3143), .ZN(n2372) );
  AND2_X1 U2703 ( .A1(n2864), .A2(n2863), .ZN(n3642) );
  XNOR2_X1 U2704 ( .A(n2610), .B(n2920), .ZN(n2614) );
  INV_X1 U2705 ( .A(n3352), .ZN(n2682) );
  NAND2_X1 U2706 ( .A1(n2678), .A2(n3351), .ZN(n2683) );
  OR2_X1 U2707 ( .A1(n2855), .A2(n2854), .ZN(n3688) );
  NAND2_X1 U2708 ( .A1(n2450), .A2(n2449), .ZN(n2735) );
  OAI21_X1 U2709 ( .B1(n2453), .B2(n2263), .A(n2452), .ZN(n2449) );
  INV_X1 U2710 ( .A(n2778), .ZN(n2774) );
  INV_X1 U2711 ( .A(n2989), .ZN(n3008) );
  INV_X1 U2712 ( .A(n2542), .ZN(n3848) );
  NAND2_X1 U2713 ( .A1(n4379), .A2(n3959), .ZN(n2986) );
  AND2_X1 U2714 ( .A1(n5039), .A2(n2390), .ZN(n5036) );
  NOR2_X1 U2715 ( .A1(n5035), .A2(n5034), .ZN(n2390) );
  NAND2_X1 U2716 ( .A1(n2287), .A2(n2286), .ZN(n5043) );
  NAND2_X1 U2717 ( .A1(n3143), .A2(n3247), .ZN(n2286) );
  OR2_X1 U2718 ( .A1(n3143), .A2(n3247), .ZN(n2287) );
  NAND2_X1 U2719 ( .A1(n5043), .A2(n5044), .ZN(n5041) );
  NOR2_X1 U2720 ( .A1(n3917), .A2(n3916), .ZN(n3915) );
  NOR2_X1 U2721 ( .A1(n3915), .A2(n3145), .ZN(n3146) );
  AND2_X1 U2722 ( .A1(n3144), .A2(REG1_REG_2__SCAN_IN), .ZN(n3145) );
  NAND2_X1 U2723 ( .A1(n3911), .A2(n2254), .ZN(n2420) );
  NAND2_X1 U2724 ( .A1(n3133), .A2(n4432), .ZN(n2285) );
  INV_X1 U2725 ( .A(n3148), .ZN(n2401) );
  AND2_X1 U2726 ( .A1(n3147), .A2(n4432), .ZN(n2404) );
  NAND2_X1 U2727 ( .A1(n4469), .A2(n3516), .ZN(n3517) );
  NOR2_X1 U2728 ( .A1(n4483), .A2(n3504), .ZN(n2388) );
  NAND2_X1 U2729 ( .A1(n2387), .A2(n4381), .ZN(n3929) );
  INV_X1 U2730 ( .A(n2388), .ZN(n2387) );
  XNOR2_X1 U2731 ( .A(n3944), .B(n2417), .ZN(n3519) );
  NAND2_X1 U2732 ( .A1(n3519), .A2(REG2_REG_12__SCAN_IN), .ZN(n3945) );
  AND2_X1 U2733 ( .A1(n3948), .A2(n4512), .ZN(n3949) );
  XNOR2_X1 U2734 ( .A(n3937), .B(n4587), .ZN(n4529) );
  NOR2_X1 U2735 ( .A1(n4516), .A2(n2421), .ZN(n3952) );
  AND2_X1 U2736 ( .A1(n3951), .A2(REG2_REG_15__SCAN_IN), .ZN(n2421) );
  NAND2_X1 U2737 ( .A1(n4538), .A2(n4539), .ZN(n4537) );
  INV_X1 U2738 ( .A(IR_REG_19__SCAN_IN), .ZN(n2532) );
  AND2_X1 U2739 ( .A1(n3876), .A2(n3845), .ZN(n3964) );
  NOR2_X1 U2740 ( .A1(n2253), .A2(n2359), .ZN(n2358) );
  NAND2_X1 U2741 ( .A1(n4045), .A2(n2361), .ZN(n2360) );
  INV_X1 U2742 ( .A(n3964), .ZN(n3966) );
  INV_X1 U2743 ( .A(n3616), .ZN(n3995) );
  NAND2_X1 U2744 ( .A1(n2307), .A2(n2305), .ZN(n3606) );
  NOR2_X1 U2745 ( .A1(n2304), .A2(n3780), .ZN(n4012) );
  INV_X1 U2746 ( .A(n2307), .ZN(n2304) );
  NAND2_X1 U2747 ( .A1(n2867), .A2(n2866), .ZN(n2875) );
  INV_X1 U2748 ( .A(n2865), .ZN(n2867) );
  AND2_X1 U2749 ( .A1(n3741), .A2(DATAI_23_), .ZN(n4054) );
  NAND2_X1 U2750 ( .A1(n4073), .A2(n2382), .ZN(n3044) );
  AOI21_X1 U2751 ( .B1(n4106), .B2(n3867), .A(n3866), .ZN(n4087) );
  INV_X1 U2752 ( .A(n2831), .ZN(n2829) );
  NAND2_X1 U2753 ( .A1(n2802), .A2(REG3_REG_17__SCAN_IN), .ZN(n2815) );
  INV_X1 U2754 ( .A(n2804), .ZN(n2802) );
  AOI21_X1 U2755 ( .B1(n2242), .B2(n2236), .A(n2268), .ZN(n2353) );
  NAND2_X1 U2756 ( .A1(n3568), .A2(n2242), .ZN(n2354) );
  NAND2_X1 U2757 ( .A1(n2311), .A2(n2313), .ZN(n4166) );
  AND2_X1 U2758 ( .A1(n3477), .A2(n2271), .ZN(n3575) );
  INV_X1 U2759 ( .A(REG3_REG_16__SCAN_IN), .ZN(n4396) );
  NAND2_X1 U2760 ( .A1(n3069), .A2(n3812), .ZN(n4183) );
  NAND2_X1 U2761 ( .A1(n2766), .A2(n2765), .ZN(n2780) );
  AND2_X1 U2762 ( .A1(REG3_REG_14__SCAN_IN), .A2(REG3_REG_15__SCAN_IN), .ZN(
        n2765) );
  AND2_X1 U2763 ( .A1(n2737), .A2(REG3_REG_13__SCAN_IN), .ZN(n2766) );
  NAND2_X1 U2764 ( .A1(n3060), .A2(n3822), .ZN(n3471) );
  INV_X1 U2765 ( .A(REG3_REG_10__SCAN_IN), .ZN(n3412) );
  INV_X1 U2766 ( .A(n3425), .ZN(n3420) );
  NAND2_X1 U2767 ( .A1(n2323), .A2(n3807), .ZN(n3419) );
  NAND2_X1 U2768 ( .A1(n2322), .A2(n2320), .ZN(n2323) );
  NOR2_X1 U2769 ( .A1(n3823), .A2(n2321), .ZN(n2320) );
  INV_X1 U2770 ( .A(n3804), .ZN(n2321) );
  NOR2_X1 U2771 ( .A1(n3083), .A2(n3082), .ZN(n4188) );
  NAND2_X1 U2772 ( .A1(n2241), .A2(n2262), .ZN(n2335) );
  OR2_X1 U2773 ( .A1(n3372), .A2(n2337), .ZN(n2336) );
  INV_X1 U2774 ( .A(REG3_REG_9__SCAN_IN), .ZN(n2687) );
  OR2_X1 U2775 ( .A1(n2688), .A2(n2687), .ZN(n2701) );
  NAND2_X1 U2776 ( .A1(n2322), .A2(n3804), .ZN(n3379) );
  NAND2_X1 U2777 ( .A1(n2670), .A2(REG3_REG_8__SCAN_IN), .ZN(n2688) );
  CLKBUF_X1 U2778 ( .A(n4188), .Z(n4227) );
  NAND2_X1 U2779 ( .A1(n2342), .A2(n2343), .ZN(n3301) );
  INV_X1 U2780 ( .A(n2344), .ZN(n2343) );
  OAI21_X1 U2781 ( .B1(n2346), .B2(n2345), .A(n2463), .ZN(n2344) );
  OR2_X1 U2782 ( .A1(n3319), .A2(n3318), .ZN(n3057) );
  NAND2_X1 U2783 ( .A1(n3192), .A2(n2348), .ZN(n2347) );
  INV_X1 U2784 ( .A(n3195), .ZN(n3267) );
  NAND2_X1 U2785 ( .A1(n3219), .A2(n3267), .ZN(n3326) );
  NAND2_X1 U2786 ( .A1(n3055), .A2(n3793), .ZN(n3194) );
  AND2_X1 U2787 ( .A1(n3793), .A2(n3790), .ZN(n3769) );
  NOR2_X1 U2788 ( .A1(n4609), .A2(n3220), .ZN(n3219) );
  INV_X1 U2789 ( .A(n4255), .ZN(n4055) );
  INV_X1 U2790 ( .A(n4236), .ZN(n4571) );
  NAND2_X1 U2791 ( .A1(n3121), .A2(n3083), .ZN(n4574) );
  AND2_X1 U2792 ( .A1(n3089), .A2(n3116), .ZN(n3205) );
  AND2_X1 U2793 ( .A1(n2969), .A2(n3114), .ZN(n3098) );
  NAND2_X1 U2794 ( .A1(n2972), .A2(n2542), .ZN(n4255) );
  NOR2_X1 U2795 ( .A1(n4060), .A2(n4037), .ZN(n4038) );
  OR2_X1 U2796 ( .A1(n4281), .A2(n4054), .ZN(n4060) );
  NAND2_X1 U2797 ( .A1(n4096), .A2(n4081), .ZN(n4281) );
  NOR3_X1 U2798 ( .A1(n4172), .A2(n2378), .A3(n2382), .ZN(n4096) );
  NOR2_X1 U2799 ( .A1(n4172), .A2(n2378), .ZN(n4116) );
  NOR2_X1 U2800 ( .A1(n4172), .A2(n2380), .ZN(n4136) );
  INV_X1 U2801 ( .A(n3094), .ZN(n4173) );
  NAND2_X1 U2802 ( .A1(n2355), .A2(n2242), .ZN(n4189) );
  OR2_X1 U2803 ( .A1(n3568), .A2(n2236), .ZN(n2355) );
  NAND2_X1 U2804 ( .A1(n3477), .A2(n2243), .ZN(n4211) );
  NAND2_X1 U2805 ( .A1(n3477), .A2(n3488), .ZN(n3545) );
  INV_X1 U2806 ( .A(n3029), .ZN(n3488) );
  AND2_X1 U2807 ( .A1(n3449), .A2(n3459), .ZN(n3477) );
  OR2_X1 U2808 ( .A1(n3385), .A2(n3384), .ZN(n3426) );
  NOR2_X1 U2809 ( .A1(n3426), .A2(n3425), .ZN(n3449) );
  NOR2_X1 U2810 ( .A1(n3342), .A2(n3302), .ZN(n3368) );
  OR2_X1 U2811 ( .A1(n3326), .A2(n3325), .ZN(n3344) );
  NAND2_X1 U2812 ( .A1(n2369), .A2(n3289), .ZN(n3342) );
  INV_X1 U2813 ( .A(n3344), .ZN(n2369) );
  INV_X1 U2814 ( .A(n4605), .ZN(n4642) );
  AND3_X1 U2815 ( .A1(n3091), .A2(n3090), .A3(n3089), .ZN(n3099) );
  AND2_X1 U2816 ( .A1(n2544), .A2(n3117), .ZN(n3202) );
  NOR2_X1 U2817 ( .A1(n2485), .A2(IR_REG_28__SCAN_IN), .ZN(n2461) );
  INV_X1 U2818 ( .A(IR_REG_27__SCAN_IN), .ZN(n2525) );
  NAND2_X1 U2819 ( .A1(n2520), .A2(n2528), .ZN(n3762) );
  MUX2_X1 U2820 ( .A(IR_REG_31__SCAN_IN), .B(n2517), .S(IR_REG_21__SCAN_IN), 
        .Z(n2520) );
  INV_X1 U2821 ( .A(IR_REG_14__SCAN_IN), .ZN(n2476) );
  AND2_X1 U2822 ( .A1(n2521), .A2(n2474), .ZN(n2744) );
  AND2_X1 U2823 ( .A1(n2427), .A2(n2431), .ZN(n3309) );
  NAND2_X1 U2824 ( .A1(n2427), .A2(n2426), .ZN(n3307) );
  NAND2_X1 U2825 ( .A1(n2440), .A2(n2439), .ZN(n3615) );
  NAND2_X1 U2826 ( .A1(n2444), .A2(n2448), .ZN(n2439) );
  NAND2_X1 U2827 ( .A1(n3656), .A2(n2441), .ZN(n2440) );
  NOR2_X1 U2828 ( .A1(n3715), .A2(n2443), .ZN(n2441) );
  NAND2_X1 U2829 ( .A1(n2447), .A2(n2443), .ZN(n2442) );
  NAND2_X1 U2830 ( .A1(n2456), .A2(n3643), .ZN(n3696) );
  NAND2_X1 U2831 ( .A1(n3409), .A2(n2719), .ZN(n3457) );
  OR2_X1 U2832 ( .A1(n2796), .A2(n2235), .ZN(n2436) );
  NAND2_X1 U2833 ( .A1(n2446), .A2(n2445), .ZN(n3718) );
  AND2_X2 U2834 ( .A1(n2990), .A2(n3152), .ZN(n4410) );
  OR3_X1 U2835 ( .A1(n2987), .A2(n4584), .A3(n2986), .ZN(n3900) );
  INV_X1 U2836 ( .A(n3779), .ZN(n3971) );
  OAI211_X1 U2837 ( .C1(n3230), .C2(n2906), .A(n2905), .B(n2904), .ZN(n3232)
         );
  NAND2_X1 U2838 ( .A1(n2892), .A2(n2891), .ZN(n4016) );
  NAND4_X1 U2839 ( .A1(n2836), .A2(n2835), .A3(n2834), .A4(n2833), .ZN(n4112)
         );
  NAND4_X1 U2840 ( .A1(n2494), .A2(n2493), .A3(n2492), .A4(n2491), .ZN(n3543)
         );
  NAND4_X1 U2841 ( .A1(n2706), .A2(n2705), .A3(n2704), .A4(n2703), .ZN(n3905)
         );
  NAND4_X1 U2842 ( .A1(n2623), .A2(n2622), .A3(n2621), .A4(n2620), .ZN(n3196)
         );
  OR2_X1 U2843 ( .A1(n2584), .A2(n3328), .ZN(n2621) );
  NAND2_X1 U2844 ( .A1(n2589), .A2(n2588), .ZN(n4229) );
  NOR2_X1 U2845 ( .A1(n2462), .A2(n2587), .ZN(n2589) );
  OR2_X1 U2846 ( .A1(n2564), .A2(n3130), .ZN(n2568) );
  OR2_X1 U2847 ( .A1(n2584), .A2(n3168), .ZN(n2569) );
  OR2_X1 U2848 ( .A1(n2566), .A2(n2549), .ZN(n2550) );
  OR2_X1 U2849 ( .A1(n2564), .A2(n3247), .ZN(n2553) );
  OR2_X1 U2850 ( .A1(n2584), .A2(n3260), .ZN(n2552) );
  NAND4_X1 U2851 ( .A1(n2541), .A2(n2540), .A3(n2539), .A4(n2538), .ZN(n3750)
         );
  OR2_X1 U2852 ( .A1(n2566), .A2(n2537), .ZN(n2538) );
  INV_X1 U2853 ( .A(IR_REG_0__SCAN_IN), .ZN(n5035) );
  XNOR2_X1 U2854 ( .A(n2420), .B(n2419), .ZN(n4390) );
  OR2_X1 U2855 ( .A1(n2400), .A2(n2399), .ZN(n3495) );
  OAI21_X1 U2856 ( .B1(n2404), .B2(REG1_REG_4__SCAN_IN), .A(n2401), .ZN(n2399)
         );
  NOR2_X1 U2857 ( .A1(n4426), .A2(n2404), .ZN(n2400) );
  INV_X1 U2858 ( .A(n2404), .ZN(n2398) );
  NAND2_X1 U2859 ( .A1(n4426), .A2(REG1_REG_4__SCAN_IN), .ZN(n2397) );
  NAND2_X1 U2860 ( .A1(n4438), .A2(n3511), .ZN(n4452) );
  NAND2_X1 U2861 ( .A1(n4436), .A2(n3497), .ZN(n4447) );
  NAND2_X1 U2862 ( .A1(n4460), .A2(n3515), .ZN(n4470) );
  NAND2_X1 U2863 ( .A1(n4470), .A2(n4471), .ZN(n4469) );
  XNOR2_X1 U2864 ( .A(n3517), .B(n2411), .ZN(n4480) );
  INV_X1 U2865 ( .A(n2410), .ZN(n4474) );
  AND2_X1 U2866 ( .A1(n2410), .A2(n2257), .ZN(n4485) );
  NOR2_X1 U2867 ( .A1(n3505), .A2(n2487), .ZN(n3930) );
  NAND2_X1 U2868 ( .A1(n3929), .A2(n2386), .ZN(n3505) );
  NAND2_X1 U2869 ( .A1(n2388), .A2(n2417), .ZN(n2386) );
  NAND2_X1 U2870 ( .A1(n3945), .A2(n3946), .ZN(n4501) );
  NOR2_X1 U2871 ( .A1(n4506), .A2(n4215), .ZN(n4505) );
  OR2_X1 U2872 ( .A1(n3949), .A2(n2418), .ZN(n4506) );
  NOR2_X1 U2873 ( .A1(n3948), .A2(n4512), .ZN(n2418) );
  INV_X1 U2874 ( .A(n2408), .ZN(n4507) );
  OR2_X1 U2875 ( .A1(n4422), .A2(n3922), .ZN(n4551) );
  NAND2_X1 U2876 ( .A1(n2405), .A2(n2406), .ZN(n4521) );
  XNOR2_X1 U2877 ( .A(n3952), .B(n2791), .ZN(n4531) );
  NAND2_X1 U2878 ( .A1(n4541), .A2(n4542), .ZN(n4540) );
  INV_X1 U2879 ( .A(n4551), .ZN(n5042) );
  OR2_X1 U2880 ( .A1(n4422), .A2(n4419), .ZN(n4548) );
  NAND2_X1 U2881 ( .A1(n4558), .A2(n3940), .ZN(n3942) );
  AND2_X1 U2882 ( .A1(n2289), .A2(n2288), .ZN(n3956) );
  NAND2_X1 U2883 ( .A1(n4554), .A2(REG2_REG_18__SCAN_IN), .ZN(n2288) );
  OR2_X1 U2884 ( .A1(n2937), .A2(n3003), .ZN(n3610) );
  INV_X1 U2885 ( .A(n3984), .ZN(n3985) );
  NAND2_X1 U2886 ( .A1(n2368), .A2(n3048), .ZN(n4027) );
  NAND2_X1 U2887 ( .A1(n4045), .A2(n2261), .ZN(n2368) );
  NAND2_X1 U2888 ( .A1(n4123), .A2(n3040), .ZN(n2330) );
  NAND2_X1 U2889 ( .A1(n3575), .A2(n4395), .ZN(n4306) );
  NAND2_X1 U2890 ( .A1(n2340), .A2(n2341), .ZN(n3383) );
  OR2_X1 U2891 ( .A1(n3372), .A2(n3026), .ZN(n2340) );
  AND2_X1 U2892 ( .A1(n3576), .A2(n3959), .ZN(n4158) );
  NAND2_X1 U2893 ( .A1(n3192), .A2(n3193), .ZN(n2349) );
  INV_X1 U2894 ( .A(n4180), .ZN(n4196) );
  AND2_X1 U2895 ( .A1(n3202), .A2(n3087), .ZN(n4577) );
  INV_X1 U2896 ( .A(REG1_REG_2__SCAN_IN), .ZN(n4879) );
  INV_X1 U2897 ( .A(REG1_REG_0__SCAN_IN), .ZN(n5034) );
  AND2_X2 U2898 ( .A1(n3099), .A2(n3098), .ZN(n4658) );
  INV_X1 U2899 ( .A(n4658), .ZN(n4656) );
  AOI21_X1 U2900 ( .B1(n4253), .B2(n4252), .A(n4251), .ZN(n4415) );
  OAI21_X1 U2901 ( .B1(n4261), .B2(n4605), .A(n2317), .ZN(n2316) );
  NAND2_X1 U2902 ( .A1(n4260), .A2(n4619), .ZN(n2317) );
  AND2_X2 U2903 ( .A1(n3099), .A2(n3206), .ZN(n4645) );
  INV_X1 U2904 ( .A(n4584), .ZN(n3117) );
  NAND2_X1 U2905 ( .A1(n3113), .A2(n3202), .ZN(n4583) );
  INV_X1 U2906 ( .A(IR_REG_30__SCAN_IN), .ZN(n3108) );
  INV_X1 U2907 ( .A(n2490), .ZN(n4376) );
  INV_X1 U2908 ( .A(IR_REG_26__SCAN_IN), .ZN(n2496) );
  NAND2_X1 U2909 ( .A1(n2506), .A2(n2505), .ZN(n3106) );
  NAND2_X1 U2910 ( .A1(n2512), .A2(IR_REG_31__SCAN_IN), .ZN(n2513) );
  INV_X1 U2911 ( .A(n3762), .ZN(n3785) );
  XNOR2_X1 U2912 ( .A(n2607), .B(IR_REG_4__SCAN_IN), .ZN(n4432) );
  XNOR2_X1 U2913 ( .A(n2423), .B(n2422), .ZN(n3144) );
  NOR2_X1 U2914 ( .A1(n2590), .A2(n2743), .ZN(n2423) );
  NAND2_X1 U2915 ( .A1(n2416), .A2(n2413), .ZN(U3258) );
  AOI21_X1 U2916 ( .B1(n2289), .B2(n2415), .A(n2279), .ZN(n2413) );
  NAND2_X1 U2917 ( .A1(n4558), .A2(n4557), .ZN(n2416) );
  OR2_X1 U2918 ( .A1(n4003), .A2(n4323), .ZN(n3096) );
  INV_X1 U2919 ( .A(IR_REG_31__SCAN_IN), .ZN(n2743) );
  NAND2_X1 U2920 ( .A1(n2269), .A2(n2801), .ZN(n2235) );
  OR2_X1 U2921 ( .A1(n3033), .A2(n3035), .ZN(n2236) );
  AND2_X1 U2922 ( .A1(n2606), .A2(n2594), .ZN(n4383) );
  INV_X1 U2923 ( .A(n4383), .ZN(n2419) );
  NAND2_X1 U2924 ( .A1(n2632), .A2(n2631), .ZN(n2237) );
  AND2_X1 U2925 ( .A1(n2408), .A2(n3933), .ZN(n2238) );
  INV_X1 U2926 ( .A(IR_REG_2__SCAN_IN), .ZN(n2422) );
  NAND2_X1 U2927 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_27__SCAN_IN), .ZN(n2239) );
  OR2_X1 U2928 ( .A1(n4553), .A2(n4552), .ZN(n2289) );
  AND2_X1 U2929 ( .A1(n2482), .A2(n2461), .ZN(n2240) );
  OR2_X1 U2930 ( .A1(n2251), .A2(n2339), .ZN(n2241) );
  AND2_X1 U2931 ( .A1(n2356), .A2(n4190), .ZN(n2242) );
  AND2_X1 U2932 ( .A1(n3488), .A2(n3558), .ZN(n2243) );
  AND2_X1 U2933 ( .A1(n2274), .A2(n2813), .ZN(n2244) );
  INV_X1 U2934 ( .A(n3654), .ZN(n2443) );
  OR2_X1 U2935 ( .A1(n4060), .A2(n2374), .ZN(n2245) );
  AND2_X1 U2936 ( .A1(n2243), .A2(n4201), .ZN(n2246) );
  AND2_X1 U2937 ( .A1(n2349), .A2(n2352), .ZN(n3324) );
  NAND2_X1 U2938 ( .A1(n3111), .A2(n2490), .ZN(n2564) );
  XNOR2_X1 U2939 ( .A(n2515), .B(IR_REG_20__SCAN_IN), .ZN(n2542) );
  NAND2_X1 U2940 ( .A1(n2514), .A2(n2954), .ZN(n2544) );
  NAND2_X1 U2941 ( .A1(n2490), .A2(n2488), .ZN(n2566) );
  OR2_X1 U2942 ( .A1(n2508), .A2(IR_REG_18__SCAN_IN), .ZN(n2247) );
  OR2_X1 U2943 ( .A1(n2503), .A2(n2485), .ZN(n2248) );
  AND2_X1 U2944 ( .A1(n2666), .A2(n2668), .ZN(n2249) );
  AND2_X1 U2945 ( .A1(n3196), .A2(n3325), .ZN(n2250) );
  AND2_X1 U2946 ( .A1(n3414), .A2(n3395), .ZN(n2251) );
  OR2_X1 U2947 ( .A1(IR_REG_19__SCAN_IN), .A2(IR_REG_20__SCAN_IN), .ZN(n2252)
         );
  NAND2_X1 U2948 ( .A1(n3599), .A2(n3598), .ZN(n2253) );
  NAND2_X1 U2949 ( .A1(n3144), .A2(REG2_REG_2__SCAN_IN), .ZN(n2254) );
  OR2_X1 U2950 ( .A1(n2250), .A2(n2350), .ZN(n2255) );
  NAND2_X1 U2951 ( .A1(n3878), .A2(n2301), .ZN(n2256) );
  OR2_X1 U2952 ( .A1(n3503), .A2(n2411), .ZN(n2257) );
  AND2_X1 U2953 ( .A1(n2499), .A2(n2498), .ZN(n2258) );
  AND3_X1 U2954 ( .A1(n2476), .A2(n2789), .A3(n2786), .ZN(n2259) );
  OR2_X1 U2955 ( .A1(n4259), .A2(n2316), .ZN(n2260) );
  INV_X1 U2956 ( .A(n3022), .ZN(n2345) );
  OR2_X1 U2957 ( .A1(n4072), .A2(n4054), .ZN(n2261) );
  NAND2_X1 U2958 ( .A1(n3714), .A2(n2264), .ZN(n2448) );
  NAND2_X1 U2959 ( .A1(n3906), .A2(n3384), .ZN(n2262) );
  NAND3_X1 U2960 ( .A1(n2590), .A2(n2470), .A3(n4896), .ZN(n2624) );
  INV_X1 U2961 ( .A(n2624), .ZN(n2298) );
  NAND2_X1 U2962 ( .A1(n2521), .A2(n2460), .ZN(n2758) );
  XOR2_X1 U2963 ( .A(n2536), .B(n2947), .Z(n2263) );
  NAND2_X1 U2964 ( .A1(n4152), .A2(n3039), .ZN(n4123) );
  NAND2_X1 U2965 ( .A1(n2330), .A2(n3041), .ZN(n4102) );
  NAND2_X1 U2966 ( .A1(n2437), .A2(n2801), .ZN(n3664) );
  OR2_X1 U2967 ( .A1(n2912), .A2(n2911), .ZN(n2264) );
  INV_X1 U2968 ( .A(n4210), .ZN(n4201) );
  INV_X1 U2969 ( .A(n3025), .ZN(n3367) );
  INV_X1 U2970 ( .A(IR_REG_22__SCAN_IN), .ZN(n2529) );
  NAND2_X1 U2971 ( .A1(n2298), .A2(n2296), .ZN(n2707) );
  NOR3_X1 U2972 ( .A1(n4060), .A2(n2374), .A3(n3995), .ZN(n2377) );
  OR2_X1 U2973 ( .A1(n3462), .A2(n3420), .ZN(n2265) );
  INV_X1 U2974 ( .A(n2381), .ZN(n4156) );
  NOR2_X1 U2975 ( .A1(n4172), .A2(n4155), .ZN(n2381) );
  INV_X1 U2976 ( .A(n2366), .ZN(n2365) );
  NOR2_X1 U2977 ( .A1(n3049), .A2(n2367), .ZN(n2366) );
  AND2_X1 U2978 ( .A1(n4059), .A2(n3679), .ZN(n2266) );
  INV_X1 U2979 ( .A(n2305), .ZN(n2303) );
  INV_X1 U2980 ( .A(IR_REG_28__SCAN_IN), .ZN(n2527) );
  NOR2_X1 U2981 ( .A1(IR_REG_6__SCAN_IN), .A2(IR_REG_7__SCAN_IN), .ZN(n2694)
         );
  AND3_X1 U2982 ( .A1(n3614), .A2(n2444), .A3(n2442), .ZN(n2267) );
  INV_X1 U2983 ( .A(n3780), .ZN(n2306) );
  INV_X1 U2984 ( .A(IR_REG_29__SCAN_IN), .ZN(n2324) );
  AND2_X1 U2985 ( .A1(n4169), .A2(n4191), .ZN(n2268) );
  OR2_X1 U2986 ( .A1(n3665), .A2(n3666), .ZN(n2269) );
  AND2_X1 U2987 ( .A1(n2874), .A2(n3643), .ZN(n2270) );
  AND2_X1 U2988 ( .A1(n2246), .A2(n3732), .ZN(n2271) );
  AND2_X1 U2989 ( .A1(n2355), .A2(n2356), .ZN(n2272) );
  INV_X1 U2990 ( .A(n2448), .ZN(n2447) );
  AND2_X1 U2991 ( .A1(n3207), .A2(n4213), .ZN(n4581) );
  INV_X1 U2992 ( .A(REG1_REG_4__SCAN_IN), .ZN(n2403) );
  NAND2_X1 U2993 ( .A1(n3274), .A2(n3275), .ZN(n2430) );
  INV_X1 U2994 ( .A(n4593), .ZN(n2411) );
  INV_X1 U2995 ( .A(n4094), .ZN(n2382) );
  INV_X1 U2996 ( .A(n3687), .ZN(n2458) );
  INV_X1 U2997 ( .A(n3832), .ZN(n2314) );
  AND2_X1 U2998 ( .A1(n2502), .A2(n2501), .ZN(n4378) );
  AND2_X1 U2999 ( .A1(n3477), .A2(n2246), .ZN(n2273) );
  NAND2_X1 U3000 ( .A1(n2336), .A2(n2335), .ZN(n3424) );
  NAND2_X1 U3001 ( .A1(n2347), .A2(n2346), .ZN(n3332) );
  XNOR2_X1 U3002 ( .A(n2513), .B(IR_REG_24__SCAN_IN), .ZN(n2954) );
  OR2_X1 U3003 ( .A1(n2828), .A2(n2827), .ZN(n2274) );
  INV_X1 U3004 ( .A(n3095), .ZN(n4138) );
  NAND2_X1 U3005 ( .A1(n2521), .A2(n2459), .ZN(n2275) );
  INV_X1 U3006 ( .A(n3679), .ZN(n4037) );
  NAND2_X1 U3007 ( .A1(n3741), .A2(DATAI_24_), .ZN(n3679) );
  AND2_X1 U3008 ( .A1(n2430), .A2(n2237), .ZN(n2276) );
  AND2_X1 U3009 ( .A1(n3547), .A2(n4590), .ZN(n2277) );
  XNOR2_X1 U3010 ( .A(n3147), .B(n3134), .ZN(n4426) );
  NAND4_X1 U3011 ( .A1(n2551), .A2(n2553), .A3(n2552), .A4(n2550), .ZN(n3018)
         );
  OAI21_X1 U3012 ( .B1(n4427), .B2(n3135), .A(n2285), .ZN(n3508) );
  OR2_X1 U3013 ( .A1(n2734), .A2(n2733), .ZN(n2278) );
  OR2_X1 U3014 ( .A1(n4556), .A2(n2414), .ZN(n2279) );
  NAND2_X1 U3015 ( .A1(n2398), .A2(n2397), .ZN(n2280) );
  NAND2_X1 U3016 ( .A1(n3951), .A2(REG1_REG_15__SCAN_IN), .ZN(n2281) );
  INV_X1 U3017 ( .A(n2352), .ZN(n2350) );
  INV_X1 U3018 ( .A(n4381), .ZN(n2417) );
  INV_X1 U3019 ( .A(IR_REG_16__SCAN_IN), .ZN(n2789) );
  INV_X1 U3020 ( .A(n2488), .ZN(n3111) );
  NAND3_X1 U3021 ( .A1(n2483), .A2(n2324), .A3(n2240), .ZN(n3107) );
  NAND2_X1 U3022 ( .A1(n2293), .A2(n2292), .ZN(n2291) );
  AOI21_X1 U3023 ( .B1(n3946), .B2(n3479), .A(n2277), .ZN(n2292) );
  INV_X1 U3024 ( .A(n3946), .ZN(n2294) );
  NAND2_X1 U3025 ( .A1(n4531), .A2(n4193), .ZN(n4530) );
  NOR2_X1 U3026 ( .A1(n4518), .A2(n4517), .ZN(n4516) );
  NAND4_X2 U3027 ( .A1(n2296), .A2(n2297), .A3(n2459), .A4(n2298), .ZN(n2508)
         );
  INV_X1 U3028 ( .A(n2473), .ZN(n2296) );
  AND2_X2 U3029 ( .A1(n2460), .A2(n2259), .ZN(n2459) );
  NAND2_X1 U3030 ( .A1(n3992), .A2(n3993), .ZN(n3991) );
  INV_X1 U3031 ( .A(n3881), .ZN(n2308) );
  INV_X1 U3032 ( .A(n3069), .ZN(n2312) );
  OAI21_X1 U3033 ( .B1(n4224), .B2(n4225), .A(n2326), .ZN(n4613) );
  NAND2_X1 U3034 ( .A1(n2571), .A2(n3018), .ZN(n2557) );
  AND2_X1 U3035 ( .A1(n2483), .A2(n2240), .ZN(n2999) );
  NAND2_X1 U3036 ( .A1(n2327), .A2(n2331), .ZN(n3043) );
  NAND2_X1 U3037 ( .A1(n4152), .A2(n2328), .ZN(n2327) );
  NAND3_X1 U3038 ( .A1(n3192), .A2(n2348), .A3(n3022), .ZN(n2342) );
  NAND2_X1 U3039 ( .A1(n3909), .A2(n3195), .ZN(n2352) );
  INV_X1 U3040 ( .A(n3253), .ZN(n3243) );
  MUX2_X1 U3041 ( .A(n2373), .B(n2372), .S(n2572), .Z(n3253) );
  NAND2_X2 U3042 ( .A1(n2371), .A2(n2370), .ZN(n2572) );
  INV_X1 U3043 ( .A(n2377), .ZN(n3986) );
  OAI21_X1 U3044 ( .B1(n3143), .B2(n4647), .A(n2389), .ZN(n5039) );
  NAND2_X1 U3045 ( .A1(n3143), .A2(n4647), .ZN(n2389) );
  NAND2_X1 U3046 ( .A1(n3147), .A2(n2392), .ZN(n2391) );
  NAND3_X1 U3047 ( .A1(n2405), .A2(n2406), .A3(n2281), .ZN(n3937) );
  NAND3_X1 U3048 ( .A1(n2426), .A2(n3274), .A3(n3275), .ZN(n2425) );
  NAND3_X1 U3049 ( .A1(n2797), .A2(n2796), .A3(n2244), .ZN(n2434) );
  NAND3_X1 U3050 ( .A1(n2436), .A2(n2435), .A3(n2813), .ZN(n3706) );
  NAND2_X1 U3051 ( .A1(n2797), .A2(n2796), .ZN(n2437) );
  NAND2_X1 U3052 ( .A1(n2900), .A2(n3675), .ZN(n3656) );
  NAND2_X1 U3053 ( .A1(n2438), .A2(n2267), .ZN(n3017) );
  NAND3_X1 U3054 ( .A1(n2900), .A2(n2447), .A3(n3675), .ZN(n2438) );
  NAND3_X1 U3055 ( .A1(n2900), .A2(n2264), .A3(n3675), .ZN(n2446) );
  NAND2_X1 U3056 ( .A1(n2456), .A2(n2270), .ZN(n3624) );
  NAND2_X1 U3057 ( .A1(n3686), .A2(n3687), .ZN(n3648) );
  NAND2_X1 U3058 ( .A1(n2483), .A2(n2482), .ZN(n2503) );
  INV_X1 U3059 ( .A(n3372), .ZN(n3373) );
  NOR2_X1 U3060 ( .A1(n2561), .A2(n2560), .ZN(n2562) );
  XNOR2_X1 U3061 ( .A(n2559), .B(n2561), .ZN(n3250) );
  INV_X1 U3062 ( .A(n2880), .ZN(n2949) );
  NAND2_X1 U3063 ( .A1(n3195), .A2(n2880), .ZN(n2608) );
  NAND2_X1 U3064 ( .A1(n2519), .A2(n2510), .ZN(n2511) );
  AND2_X1 U3065 ( .A1(n3354), .A2(n2680), .ZN(n2681) );
  OAI21_X1 U3066 ( .B1(n4011), .B2(n3983), .A(n3982), .ZN(n3984) );
  OAI21_X1 U3067 ( .B1(n4011), .B2(n3592), .A(n3593), .ZN(n3050) );
  AOI22_X1 U3068 ( .A1(n3196), .A2(n2951), .B1(n2880), .B2(n3325), .ZN(n2628)
         );
  NAND2_X1 U3069 ( .A1(n3909), .A2(n2951), .ZN(n2609) );
  AND2_X1 U3070 ( .A1(n2563), .A2(REG1_REG_3__SCAN_IN), .ZN(n2462) );
  INV_X1 U3071 ( .A(n3733), .ZN(n3165) );
  INV_X1 U3072 ( .A(REG2_REG_1__SCAN_IN), .ZN(n3247) );
  OR2_X1 U3073 ( .A1(n3312), .A2(n3289), .ZN(n2463) );
  OR2_X1 U3074 ( .A1(n4493), .A2(n3450), .ZN(n2464) );
  AND2_X1 U3075 ( .A1(n3489), .A2(n3459), .ZN(n2465) );
  AND2_X1 U3076 ( .A1(n2580), .A2(n2579), .ZN(n2466) );
  INV_X1 U3077 ( .A(n4547), .ZN(n5046) );
  NAND4_X1 U3078 ( .A1(n2820), .A2(n2819), .A3(n2818), .A4(n2817), .ZN(n4133)
         );
  INV_X1 U3079 ( .A(n4133), .ZN(n3038) );
  INV_X1 U3080 ( .A(n4049), .ZN(n3045) );
  OR2_X1 U3081 ( .A1(n3146), .A2(n2419), .ZN(n2467) );
  AND2_X1 U3082 ( .A1(n4104), .A2(n4094), .ZN(n2468) );
  NAND2_X1 U3083 ( .A1(n3741), .A2(DATAI_21_), .ZN(n4094) );
  INV_X1 U3084 ( .A(n4073), .ZN(n4104) );
  AND3_X1 U3085 ( .A1(n2979), .A2(n4405), .A3(n2978), .ZN(n2469) );
  INV_X1 U3086 ( .A(IR_REG_18__SCAN_IN), .ZN(n2479) );
  NAND2_X1 U3087 ( .A1(n2880), .A2(n3243), .ZN(n2556) );
  INV_X1 U3088 ( .A(n4206), .ZN(n3031) );
  NAND2_X1 U3089 ( .A1(n4229), .A2(n2951), .ZN(n2596) );
  NAND2_X1 U3090 ( .A1(n3032), .A2(n3031), .ZN(n3033) );
  NAND2_X1 U3091 ( .A1(n2596), .A2(n2595), .ZN(n2597) );
  INV_X1 U3092 ( .A(REG2_REG_2__SCAN_IN), .ZN(n3130) );
  NAND2_X1 U3093 ( .A1(n3038), .A2(n4145), .ZN(n3039) );
  INV_X1 U3094 ( .A(n3697), .ZN(n2874) );
  AOI21_X1 U3095 ( .B1(n3251), .B2(n3250), .A(n2562), .ZN(n3160) );
  INV_X1 U3096 ( .A(n3513), .ZN(n3499) );
  OR2_X1 U3097 ( .A1(n3596), .A2(n3595), .ZN(n3982) );
  OR2_X1 U3098 ( .A1(n4133), .A2(n4145), .ZN(n4126) );
  AND2_X1 U3099 ( .A1(n3830), .A2(n3811), .ZN(n4206) );
  INV_X1 U3100 ( .A(n4586), .ZN(n3954) );
  NOR2_X1 U3101 ( .A1(n3394), .A2(n3367), .ZN(n3026) );
  OR2_X1 U3102 ( .A1(n3113), .A2(D_REG_1__SCAN_IN), .ZN(n3203) );
  INV_X1 U3103 ( .A(REG3_REG_7__SCAN_IN), .ZN(n2651) );
  AND3_X1 U3104 ( .A1(REG3_REG_4__SCAN_IN), .A2(REG3_REG_3__SCAN_IN), .A3(
        REG3_REG_5__SCAN_IN), .ZN(n2616) );
  INV_X1 U3105 ( .A(n2613), .ZN(n2612) );
  INV_X1 U3106 ( .A(n3442), .ZN(n3459) );
  INV_X1 U3107 ( .A(REG3_REG_18__SCAN_IN), .ZN(n4967) );
  INV_X1 U3108 ( .A(n4169), .ZN(n3735) );
  AND2_X1 U3109 ( .A1(n3610), .A2(n2938), .ZN(n3976) );
  NAND4_X1 U3110 ( .A1(n2570), .A2(n2569), .A3(n2568), .A4(n2567), .ZN(n2576)
         );
  INV_X1 U3111 ( .A(REG3_REG_11__SCAN_IN), .ZN(n3460) );
  NOR2_X1 U3112 ( .A1(n4555), .A2(n4547), .ZN(n4556) );
  INV_X1 U3113 ( .A(n4016), .ZN(n4059) );
  AND2_X1 U3114 ( .A1(n3077), .A2(n4050), .ZN(n4049) );
  INV_X1 U3115 ( .A(n4191), .ZN(n4395) );
  INV_X1 U3116 ( .A(n4239), .ZN(n4232) );
  OR2_X1 U3117 ( .A1(n3113), .A2(D_REG_0__SCAN_IN), .ZN(n2969) );
  NAND2_X1 U3118 ( .A1(n3741), .A2(DATAI_20_), .ZN(n4114) );
  AND2_X1 U3119 ( .A1(n3888), .A2(n3080), .ZN(n4236) );
  OR2_X1 U3120 ( .A1(n3113), .A2(n2967), .ZN(n3089) );
  NOR2_X1 U3121 ( .A1(n2652), .A2(n2651), .ZN(n2670) );
  OR2_X1 U3122 ( .A1(n2875), .A2(n3629), .ZN(n2902) );
  NAND2_X1 U3123 ( .A1(n2829), .A2(REG3_REG_19__SCAN_IN), .ZN(n2844) );
  AND2_X1 U3124 ( .A1(n2722), .A2(REG3_REG_12__SCAN_IN), .ZN(n2737) );
  OR2_X1 U3125 ( .A1(n2780), .A2(n4396), .ZN(n2804) );
  AND2_X1 U3126 ( .A1(n3008), .A2(n3002), .ZN(n3618) );
  OR2_X1 U3127 ( .A1(n2844), .A2(n4867), .ZN(n2865) );
  NOR2_X1 U3128 ( .A1(n2721), .A2(n3460), .ZN(n2722) );
  OR2_X1 U3129 ( .A1(n2815), .A2(n4967), .ZN(n2831) );
  AND2_X2 U3130 ( .A1(n3008), .A2(n2974), .ZN(n4405) );
  AND2_X1 U3131 ( .A1(n2934), .A2(n2933), .ZN(n3779) );
  AND4_X1 U3132 ( .A1(n2872), .A2(n2871), .A3(n2870), .A4(n2869), .ZN(n4089)
         );
  NAND4_X1 U3133 ( .A1(n2742), .A2(n2741), .A3(n2740), .A4(n2739), .ZN(n4203)
         );
  NAND2_X1 U3134 ( .A1(n4489), .A2(n4490), .ZN(n4488) );
  INV_X1 U3135 ( .A(n4548), .ZN(n5038) );
  AOI22_X1 U3136 ( .A1(n3965), .A2(n3966), .B1(n3975), .B2(n3990), .ZN(n3601)
         );
  AND2_X1 U3137 ( .A1(n4158), .A2(n4619), .ZN(n4563) );
  AND2_X1 U3138 ( .A1(n4658), .A2(n4619), .ZN(n4264) );
  INV_X1 U3139 ( .A(n3034), .ZN(n3732) );
  AND2_X1 U3140 ( .A1(n4645), .A2(n4619), .ZN(n4329) );
  INV_X1 U3141 ( .A(n4638), .ZN(n4619) );
  INV_X1 U3142 ( .A(n3098), .ZN(n3206) );
  NAND2_X1 U3143 ( .A1(n3120), .A2(STATE_REG_SCAN_IN), .ZN(n4584) );
  AND2_X1 U3144 ( .A1(n2676), .A2(n2661), .ZN(n4445) );
  AND2_X1 U3145 ( .A1(n3128), .A2(n3122), .ZN(n5045) );
  AND2_X1 U3146 ( .A1(n3013), .A2(n3012), .ZN(n3014) );
  NAND2_X1 U3147 ( .A1(n2943), .A2(n2942), .ZN(n3990) );
  NAND4_X1 U31480 ( .A1(n2785), .A2(n2784), .A3(n2783), .A4(n2782), .ZN(n4169)
         );
  OR2_X1 U31490 ( .A1(n2544), .A2(n4584), .ZN(n3910) );
  INV_X1 U3150 ( .A(n4382), .ZN(n3509) );
  OR2_X1 U3151 ( .A1(n4422), .A2(n4377), .ZN(n4547) );
  NAND2_X1 U3152 ( .A1(n3576), .A2(n3239), .ZN(n4180) );
  INV_X1 U3153 ( .A(n4563), .ZN(n4175) );
  INV_X1 U3154 ( .A(n4264), .ZN(n4323) );
  OR2_X1 U3155 ( .A1(n4003), .A2(n4374), .ZN(n3102) );
  INV_X1 U3156 ( .A(n4329), .ZN(n4374) );
  INV_X1 U3157 ( .A(n4645), .ZN(n4644) );
  INV_X1 U3158 ( .A(n4583), .ZN(n4582) );
  INV_X1 U3159 ( .A(n3897), .ZN(n4379) );
  AND2_X1 U3160 ( .A1(n2626), .A2(n2697), .ZN(n4382) );
  NAND4_X1 U3161 ( .A1(n2694), .A2(n2472), .A3(n2471), .A4(n2695), .ZN(n2473)
         );
  INV_X1 U3162 ( .A(n2499), .ZN(n2484) );
  NAND2_X1 U3163 ( .A1(n2991), .A2(REG0_REG_12__SCAN_IN), .ZN(n2494) );
  INV_X1 U3164 ( .A(REG1_REG_12__SCAN_IN), .ZN(n2487) );
  OR2_X1 U3165 ( .A1(n2601), .A2(n2487), .ZN(n2493) );
  NAND2_X2 U3166 ( .A1(n3111), .A2(n4376), .ZN(n2584) );
  NAND2_X1 U3167 ( .A1(n2616), .A2(REG3_REG_6__SCAN_IN), .ZN(n2652) );
  NOR2_X1 U3168 ( .A1(n2722), .A2(REG3_REG_12__SCAN_IN), .ZN(n2489) );
  OR2_X1 U3169 ( .A1(n2737), .A2(n2489), .ZN(n3494) );
  OR2_X1 U3170 ( .A1(n2584), .A2(n3494), .ZN(n2492) );
  INV_X1 U3171 ( .A(REG2_REG_12__SCAN_IN), .ZN(n3479) );
  OR2_X1 U3172 ( .A1(n3230), .A2(n3479), .ZN(n2491) );
  INV_X1 U3173 ( .A(n2503), .ZN(n2498) );
  INV_X1 U3174 ( .A(IR_REG_25__SCAN_IN), .ZN(n2495) );
  NAND2_X1 U3175 ( .A1(n2498), .A2(n2495), .ZN(n2505) );
  NAND2_X1 U3176 ( .A1(n2505), .A2(IR_REG_31__SCAN_IN), .ZN(n2497) );
  OR2_X1 U3177 ( .A1(n2497), .A2(n2496), .ZN(n2502) );
  NOR2_X1 U3178 ( .A1(n2258), .A2(n2500), .ZN(n2501) );
  INV_X1 U3179 ( .A(n4378), .ZN(n2507) );
  NAND2_X1 U3180 ( .A1(n2503), .A2(IR_REG_31__SCAN_IN), .ZN(n2504) );
  MUX2_X1 U3181 ( .A(IR_REG_31__SCAN_IN), .B(n2504), .S(IR_REG_25__SCAN_IN), 
        .Z(n2506) );
  NAND2_X1 U3182 ( .A1(n2971), .A2(n2970), .ZN(n2512) );
  INV_X1 U3183 ( .A(n2519), .ZN(n2516) );
  NAND2_X1 U3184 ( .A1(n2516), .A2(IR_REG_31__SCAN_IN), .ZN(n2517) );
  NAND2_X1 U3185 ( .A1(n2519), .A2(n2518), .ZN(n2528) );
  AND2_X4 U3186 ( .A1(n2535), .A2(n2544), .ZN(n2880) );
  OR2_X1 U3187 ( .A1(n2521), .A2(n2743), .ZN(n2728) );
  INV_X1 U3188 ( .A(IR_REG_11__SCAN_IN), .ZN(n2522) );
  NAND2_X1 U3189 ( .A1(n2728), .A2(n2522), .ZN(n2523) );
  NAND2_X1 U3190 ( .A1(n2523), .A2(IR_REG_31__SCAN_IN), .ZN(n2524) );
  XNOR2_X1 U3191 ( .A(n2524), .B(IR_REG_12__SCAN_IN), .ZN(n4381) );
  NAND2_X1 U3192 ( .A1(n2743), .A2(n2525), .ZN(n2526) );
  MUX2_X1 U3193 ( .A(DATAI_12_), .B(n4381), .S(n2572), .Z(n3029) );
  AOI22_X1 U3194 ( .A1(n3543), .A2(n2951), .B1(n2880), .B2(n3029), .ZN(n2536)
         );
  NAND2_X1 U3195 ( .A1(n2528), .A2(IR_REG_31__SCAN_IN), .ZN(n2530) );
  OR2_X1 U3196 ( .A1(n2533), .A2(n2532), .ZN(n2534) );
  NAND2_X4 U3197 ( .A1(n2535), .A2(n2986), .ZN(n2947) );
  NAND2_X1 U3198 ( .A1(n2684), .A2(REG2_REG_0__SCAN_IN), .ZN(n2541) );
  INV_X1 U3199 ( .A(REG3_REG_0__SCAN_IN), .ZN(n3159) );
  OR2_X1 U3200 ( .A1(n2584), .A2(n3159), .ZN(n2540) );
  OR2_X1 U3201 ( .A1(n2601), .A2(n5034), .ZN(n2539) );
  INV_X1 U3202 ( .A(REG0_REG_0__SCAN_IN), .ZN(n2537) );
  AND2_X4 U3203 ( .A1(n2880), .A2(n4638), .ZN(n2795) );
  INV_X1 U3204 ( .A(DATAI_0_), .ZN(n2543) );
  MUX2_X1 U3205 ( .A(n2543), .B(n5035), .S(n2572), .Z(n4569) );
  OAI22_X1 U3206 ( .A1(n4569), .A2(n2944), .B1(n2544), .B2(n5035), .ZN(n2545)
         );
  AOI21_X1 U3207 ( .B1(n3750), .B2(n2795), .A(n2545), .ZN(n3155) );
  INV_X1 U3208 ( .A(n4569), .ZN(n3236) );
  NAND2_X1 U3209 ( .A1(n2880), .A2(n3236), .ZN(n2547) );
  OAI21_X1 U32100 ( .B1(n2544), .B2(n5034), .A(n2547), .ZN(n2546) );
  AOI21_X1 U32110 ( .B1(n3750), .B2(n2571), .A(n2546), .ZN(n3156) );
  INV_X1 U32120 ( .A(n2547), .ZN(n2548) );
  OAI22_X1 U32130 ( .A1(n3155), .A2(n3156), .B1(n2548), .B2(n2947), .ZN(n3251)
         );
  INV_X1 U32140 ( .A(REG3_REG_1__SCAN_IN), .ZN(n3260) );
  NAND2_X1 U32150 ( .A1(n2563), .A2(REG1_REG_1__SCAN_IN), .ZN(n2551) );
  INV_X1 U32160 ( .A(REG0_REG_1__SCAN_IN), .ZN(n2549) );
  NAND2_X1 U32170 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n2554) );
  NOR2_X1 U32180 ( .A1(n3253), .A2(n2944), .ZN(n2555) );
  INV_X1 U32190 ( .A(n2560), .ZN(n2559) );
  NAND2_X1 U32200 ( .A1(n2557), .A2(n2556), .ZN(n2558) );
  XNOR2_X1 U32210 ( .A(n2558), .B(n2920), .ZN(n2561) );
  NAND2_X1 U32220 ( .A1(n2563), .A2(REG1_REG_2__SCAN_IN), .ZN(n2570) );
  INV_X1 U32230 ( .A(REG3_REG_2__SCAN_IN), .ZN(n3168) );
  INV_X1 U32240 ( .A(REG0_REG_2__SCAN_IN), .ZN(n2565) );
  OR2_X1 U32250 ( .A1(n2566), .A2(n2565), .ZN(n2567) );
  NAND2_X1 U32260 ( .A1(n2576), .A2(n2571), .ZN(n2574) );
  MUX2_X1 U32270 ( .A(DATAI_2_), .B(n3144), .S(n2572), .Z(n4239) );
  NAND2_X1 U32280 ( .A1(n2880), .A2(n4239), .ZN(n2573) );
  NAND2_X1 U32290 ( .A1(n2574), .A2(n2573), .ZN(n2575) );
  NAND2_X1 U32300 ( .A1(n2576), .A2(n2795), .ZN(n2578) );
  NAND2_X1 U32310 ( .A1(n2571), .A2(n4239), .ZN(n2577) );
  NAND2_X1 U32320 ( .A1(n2578), .A2(n2577), .ZN(n2579) );
  NOR2_X1 U32330 ( .A1(n2580), .A2(n2579), .ZN(n2581) );
  NAND2_X1 U32340 ( .A1(n3160), .A2(n3162), .ZN(n3161) );
  INV_X1 U32350 ( .A(n2581), .ZN(n2582) );
  NAND2_X1 U32360 ( .A1(n3161), .A2(n2582), .ZN(n3170) );
  INV_X1 U32370 ( .A(REG0_REG_3__SCAN_IN), .ZN(n2583) );
  OR2_X1 U32380 ( .A1(n2566), .A2(n2583), .ZN(n2586) );
  OR2_X1 U32390 ( .A1(n2584), .A2(REG3_REG_3__SCAN_IN), .ZN(n2585) );
  NAND2_X1 U32400 ( .A1(n2586), .A2(n2585), .ZN(n2587) );
  INV_X1 U32410 ( .A(REG2_REG_3__SCAN_IN), .ZN(n3221) );
  OR2_X1 U32420 ( .A1(n3230), .A2(n3221), .ZN(n2588) );
  NAND2_X1 U32430 ( .A1(n2590), .A2(n2422), .ZN(n2591) );
  NAND2_X1 U32440 ( .A1(n2591), .A2(IR_REG_31__SCAN_IN), .ZN(n2593) );
  NAND2_X1 U32450 ( .A1(n2593), .A2(n2592), .ZN(n2606) );
  OR2_X1 U32460 ( .A1(n2593), .A2(n2592), .ZN(n2594) );
  MUX2_X1 U32470 ( .A(DATAI_3_), .B(n4383), .S(n2572), .Z(n3220) );
  NAND2_X1 U32480 ( .A1(n2880), .A2(n3220), .ZN(n2595) );
  AOI22_X1 U32490 ( .A1(n4229), .A2(n2795), .B1(n2951), .B2(n3220), .ZN(n2599)
         );
  XNOR2_X1 U32500 ( .A(n2598), .B(n2599), .ZN(n3171) );
  NAND2_X1 U32510 ( .A1(n3170), .A2(n3171), .ZN(n3169) );
  INV_X1 U32520 ( .A(n2598), .ZN(n2600) );
  NAND2_X1 U32530 ( .A1(n2600), .A2(n2599), .ZN(n3262) );
  NAND2_X1 U32540 ( .A1(n2991), .A2(REG0_REG_4__SCAN_IN), .ZN(n2605) );
  OR2_X1 U32550 ( .A1(n2601), .A2(n2403), .ZN(n2604) );
  XNOR2_X1 U32560 ( .A(REG3_REG_4__SCAN_IN), .B(REG3_REG_3__SCAN_IN), .ZN(
        n3273) );
  INV_X1 U32570 ( .A(REG2_REG_4__SCAN_IN), .ZN(n3135) );
  OR2_X1 U32580 ( .A1(n3230), .A2(n3135), .ZN(n2602) );
  NAND2_X1 U32590 ( .A1(n2606), .A2(IR_REG_31__SCAN_IN), .ZN(n2607) );
  MUX2_X1 U32600 ( .A(DATAI_4_), .B(n4432), .S(n2572), .Z(n3195) );
  NAND2_X1 U32610 ( .A1(n2609), .A2(n2608), .ZN(n2610) );
  NOR2_X1 U32620 ( .A1(n3267), .A2(n2987), .ZN(n2611) );
  AOI21_X1 U32630 ( .B1(n3909), .B2(n2795), .A(n2611), .ZN(n2613) );
  XNOR2_X1 U32640 ( .A(n2614), .B(n2612), .ZN(n3264) );
  NAND3_X1 U32650 ( .A1(n3169), .A2(n3262), .A3(n3264), .ZN(n3263) );
  OR2_X1 U32660 ( .A1(n2614), .A2(n2613), .ZN(n2615) );
  NAND2_X1 U32670 ( .A1(n3263), .A2(n2615), .ZN(n3274) );
  NAND2_X1 U32680 ( .A1(n2991), .A2(REG0_REG_5__SCAN_IN), .ZN(n2623) );
  INV_X1 U32690 ( .A(REG1_REG_5__SCAN_IN), .ZN(n3142) );
  OR2_X1 U32700 ( .A1(n2601), .A2(n3142), .ZN(n2622) );
  INV_X1 U32710 ( .A(n2616), .ZN(n2633) );
  INV_X1 U32720 ( .A(REG3_REG_5__SCAN_IN), .ZN(n2618) );
  NAND2_X1 U32730 ( .A1(REG3_REG_4__SCAN_IN), .A2(REG3_REG_3__SCAN_IN), .ZN(
        n2617) );
  NAND2_X1 U32740 ( .A1(n2618), .A2(n2617), .ZN(n2619) );
  NAND2_X1 U32750 ( .A1(n2633), .A2(n2619), .ZN(n3328) );
  INV_X1 U32760 ( .A(REG2_REG_5__SCAN_IN), .ZN(n3129) );
  OR2_X1 U32770 ( .A1(n3230), .A2(n3129), .ZN(n2620) );
  NAND2_X1 U32780 ( .A1(n2624), .A2(IR_REG_31__SCAN_IN), .ZN(n2625) );
  MUX2_X1 U32790 ( .A(IR_REG_31__SCAN_IN), .B(n2625), .S(IR_REG_5__SCAN_IN), 
        .Z(n2626) );
  OR2_X1 U32800 ( .A1(n2624), .A2(IR_REG_5__SCAN_IN), .ZN(n2697) );
  MUX2_X1 U32810 ( .A(DATAI_5_), .B(n4382), .S(n2572), .Z(n3325) );
  INV_X1 U32820 ( .A(n3325), .ZN(n3277) );
  NOR2_X1 U32830 ( .A1(n3277), .A2(n2987), .ZN(n2627) );
  AOI21_X1 U32840 ( .B1(n3196), .B2(n2795), .A(n2627), .ZN(n2630) );
  XNOR2_X1 U32850 ( .A(n2628), .B(n2947), .ZN(n2629) );
  XOR2_X1 U32860 ( .A(n2630), .B(n2629), .Z(n3275) );
  INV_X1 U32870 ( .A(n2629), .ZN(n2632) );
  INV_X1 U32880 ( .A(n2630), .ZN(n2631) );
  NAND2_X1 U32890 ( .A1(n2991), .A2(REG0_REG_6__SCAN_IN), .ZN(n2640) );
  INV_X1 U32900 ( .A(REG3_REG_6__SCAN_IN), .ZN(n4963) );
  NAND2_X1 U32910 ( .A1(n2633), .A2(n4963), .ZN(n2634) );
  AND2_X1 U32920 ( .A1(n2634), .A2(n2652), .ZN(n4561) );
  INV_X1 U32930 ( .A(n4561), .ZN(n3295) );
  OR2_X1 U32940 ( .A1(n2584), .A2(n3295), .ZN(n2639) );
  INV_X1 U32950 ( .A(REG1_REG_6__SCAN_IN), .ZN(n2635) );
  OR2_X1 U32960 ( .A1(n2601), .A2(n2635), .ZN(n2638) );
  INV_X1 U32970 ( .A(REG2_REG_6__SCAN_IN), .ZN(n2636) );
  OR2_X1 U32980 ( .A1(n3230), .A2(n2636), .ZN(n2637) );
  NAND4_X1 U32990 ( .A1(n2640), .A2(n2639), .A3(n2638), .A4(n2637), .ZN(n3908)
         );
  NAND2_X1 U33000 ( .A1(n3908), .A2(n2951), .ZN(n2643) );
  NAND2_X1 U33010 ( .A1(n2697), .A2(IR_REG_31__SCAN_IN), .ZN(n2641) );
  XNOR2_X1 U33020 ( .A(n2641), .B(IR_REG_6__SCAN_IN), .ZN(n4440) );
  MUX2_X1 U33030 ( .A(DATAI_6_), .B(n4440), .S(n2572), .Z(n3345) );
  NAND2_X1 U33040 ( .A1(n2880), .A2(n3345), .ZN(n2642) );
  NAND2_X1 U33050 ( .A1(n2643), .A2(n2642), .ZN(n2644) );
  XNOR2_X1 U33060 ( .A(n2644), .B(n2920), .ZN(n2649) );
  INV_X1 U33070 ( .A(n2649), .ZN(n2647) );
  INV_X1 U33080 ( .A(n3345), .ZN(n3289) );
  NOR2_X1 U33090 ( .A1(n3289), .A2(n2987), .ZN(n2645) );
  AOI21_X1 U33100 ( .B1(n3908), .B2(n2795), .A(n2645), .ZN(n2648) );
  INV_X1 U33110 ( .A(n2648), .ZN(n2646) );
  NAND2_X1 U33120 ( .A1(n2647), .A2(n2646), .ZN(n3284) );
  AND2_X1 U33130 ( .A1(n2649), .A2(n2648), .ZN(n3285) );
  NAND2_X1 U33140 ( .A1(n2991), .A2(REG0_REG_7__SCAN_IN), .ZN(n2658) );
  INV_X1 U33150 ( .A(REG1_REG_7__SCAN_IN), .ZN(n2650) );
  OR2_X1 U33160 ( .A1(n2601), .A2(n2650), .ZN(n2657) );
  AND2_X1 U33170 ( .A1(n2652), .A2(n2651), .ZN(n2653) );
  OR2_X1 U33180 ( .A1(n2653), .A2(n2670), .ZN(n3317) );
  OR2_X1 U33190 ( .A1(n2584), .A2(n3317), .ZN(n2656) );
  INV_X1 U33200 ( .A(REG2_REG_7__SCAN_IN), .ZN(n2654) );
  OR2_X1 U33210 ( .A1(n3230), .A2(n2654), .ZN(n2655) );
  NAND4_X1 U33220 ( .A1(n2658), .A2(n2657), .A3(n2656), .A4(n2655), .ZN(n3366)
         );
  NAND2_X1 U33230 ( .A1(n3366), .A2(n2951), .ZN(n2663) );
  OAI21_X1 U33240 ( .B1(n2697), .B2(IR_REG_6__SCAN_IN), .A(IR_REG_31__SCAN_IN), 
        .ZN(n2660) );
  NAND2_X1 U33250 ( .A1(n2660), .A2(n2659), .ZN(n2676) );
  OR2_X1 U33260 ( .A1(n2660), .A2(n2659), .ZN(n2661) );
  MUX2_X1 U33270 ( .A(DATAI_7_), .B(n4445), .S(n2572), .Z(n3302) );
  NAND2_X1 U33280 ( .A1(n2880), .A2(n3302), .ZN(n2662) );
  NAND2_X1 U33290 ( .A1(n2663), .A2(n2662), .ZN(n2664) );
  XNOR2_X1 U33300 ( .A(n2664), .B(n2947), .ZN(n2666) );
  INV_X1 U33310 ( .A(n3302), .ZN(n3310) );
  NOR2_X1 U33320 ( .A1(n3310), .A2(n2987), .ZN(n2665) );
  AOI21_X1 U33330 ( .B1(n3366), .B2(n2795), .A(n2665), .ZN(n2667) );
  XNOR2_X1 U33340 ( .A(n2666), .B(n2667), .ZN(n3308) );
  INV_X1 U33350 ( .A(n2667), .ZN(n2668) );
  INV_X1 U33360 ( .A(n3354), .ZN(n2678) );
  NAND2_X1 U33370 ( .A1(n2991), .A2(REG0_REG_8__SCAN_IN), .ZN(n2675) );
  INV_X1 U33380 ( .A(REG1_REG_8__SCAN_IN), .ZN(n2669) );
  OR2_X1 U33390 ( .A1(n2601), .A2(n2669), .ZN(n2674) );
  OR2_X1 U33400 ( .A1(n2670), .A2(REG3_REG_8__SCAN_IN), .ZN(n2671) );
  NAND2_X1 U33410 ( .A1(n2688), .A2(n2671), .ZN(n3370) );
  OR2_X1 U33420 ( .A1(n2584), .A2(n3370), .ZN(n2673) );
  INV_X1 U33430 ( .A(REG2_REG_8__SCAN_IN), .ZN(n3371) );
  OR2_X1 U33440 ( .A1(n3230), .A2(n3371), .ZN(n2672) );
  NAND4_X1 U33450 ( .A1(n2675), .A2(n2674), .A3(n2673), .A4(n2672), .ZN(n3907)
         );
  NAND2_X1 U33460 ( .A1(n2676), .A2(IR_REG_31__SCAN_IN), .ZN(n2677) );
  XNOR2_X1 U33470 ( .A(n2677), .B(IR_REG_8__SCAN_IN), .ZN(n3513) );
  MUX2_X1 U33480 ( .A(DATAI_8_), .B(n3513), .S(n2572), .Z(n3025) );
  AOI22_X1 U33490 ( .A1(n3907), .A2(n2795), .B1(n2951), .B2(n3025), .ZN(n3351)
         );
  AOI22_X1 U33500 ( .A1(n3907), .A2(n2951), .B1(n2880), .B2(n3025), .ZN(n2679)
         );
  XNOR2_X1 U33510 ( .A(n2679), .B(n2947), .ZN(n3352) );
  INV_X1 U33520 ( .A(n3351), .ZN(n2680) );
  AOI21_X2 U3353 ( .B1(n2683), .B2(n2682), .A(n2681), .ZN(n3390) );
  NAND2_X1 U33540 ( .A1(n2684), .A2(REG2_REG_9__SCAN_IN), .ZN(n2693) );
  INV_X1 U3355 ( .A(REG1_REG_9__SCAN_IN), .ZN(n2685) );
  OR2_X1 U3356 ( .A1(n2601), .A2(n2685), .ZN(n2692) );
  INV_X1 U3357 ( .A(REG0_REG_9__SCAN_IN), .ZN(n2686) );
  OR2_X1 U3358 ( .A1(n2566), .A2(n2686), .ZN(n2691) );
  NAND2_X1 U3359 ( .A1(n2688), .A2(n2687), .ZN(n2689) );
  NAND2_X1 U3360 ( .A1(n2701), .A2(n2689), .ZN(n3399) );
  OR2_X1 U3361 ( .A1(n2584), .A2(n3399), .ZN(n2690) );
  NAND4_X1 U3362 ( .A1(n2693), .A2(n2692), .A3(n2691), .A4(n2690), .ZN(n3906)
         );
  NAND2_X1 U3363 ( .A1(n2694), .A2(n2695), .ZN(n2696) );
  OAI21_X1 U3364 ( .B1(n2697), .B2(n2696), .A(IR_REG_31__SCAN_IN), .ZN(n2698)
         );
  XNOR2_X1 U3365 ( .A(n2698), .B(IR_REG_9__SCAN_IN), .ZN(n3507) );
  MUX2_X1 U3366 ( .A(DATAI_9_), .B(n3507), .S(n2572), .Z(n3384) );
  AOI22_X1 U3367 ( .A1(n3906), .A2(n2795), .B1(n2951), .B2(n3384), .ZN(n2713)
         );
  AOI22_X1 U3368 ( .A1(n3906), .A2(n2951), .B1(n2880), .B2(n3384), .ZN(n2699)
         );
  XNOR2_X1 U3369 ( .A(n2699), .B(n2947), .ZN(n2714) );
  XOR2_X1 U3370 ( .A(n2713), .B(n2714), .Z(n3392) );
  NAND2_X1 U3371 ( .A1(n3390), .A2(n3392), .ZN(n3391) );
  NAND2_X1 U3372 ( .A1(n2563), .A2(REG1_REG_10__SCAN_IN), .ZN(n2706) );
  INV_X1 U3373 ( .A(REG0_REG_10__SCAN_IN), .ZN(n2700) );
  OR2_X1 U3374 ( .A1(n2566), .A2(n2700), .ZN(n2705) );
  NAND2_X1 U3375 ( .A1(n2701), .A2(n3412), .ZN(n2702) );
  NAND2_X1 U3376 ( .A1(n2721), .A2(n2702), .ZN(n3429) );
  OR2_X1 U3377 ( .A1(n2584), .A2(n3429), .ZN(n2704) );
  INV_X1 U3378 ( .A(REG2_REG_10__SCAN_IN), .ZN(n3430) );
  OR2_X1 U3379 ( .A1(n3230), .A2(n3430), .ZN(n2703) );
  NAND2_X1 U3380 ( .A1(n3905), .A2(n2951), .ZN(n2710) );
  NAND2_X1 U3381 ( .A1(n2707), .A2(IR_REG_31__SCAN_IN), .ZN(n2708) );
  XNOR2_X1 U3382 ( .A(n2708), .B(IR_REG_10__SCAN_IN), .ZN(n4593) );
  MUX2_X1 U3383 ( .A(DATAI_10_), .B(n4593), .S(n2572), .Z(n3425) );
  NAND2_X1 U3384 ( .A1(n2880), .A2(n3425), .ZN(n2709) );
  NAND2_X1 U3385 ( .A1(n2710), .A2(n2709), .ZN(n2711) );
  XNOR2_X1 U3386 ( .A(n2711), .B(n2947), .ZN(n2716) );
  NOR2_X1 U3387 ( .A1(n3420), .A2(n2987), .ZN(n2712) );
  AOI21_X1 U3388 ( .B1(n3905), .B2(n2795), .A(n2712), .ZN(n2717) );
  XNOR2_X1 U3389 ( .A(n2716), .B(n2717), .ZN(n3410) );
  NAND2_X1 U3390 ( .A1(n2714), .A2(n2713), .ZN(n3408) );
  NAND2_X1 U3391 ( .A1(n2563), .A2(REG1_REG_11__SCAN_IN), .ZN(n2727) );
  INV_X1 U3392 ( .A(REG0_REG_11__SCAN_IN), .ZN(n2720) );
  OR2_X1 U3393 ( .A1(n2566), .A2(n2720), .ZN(n2726) );
  AND2_X1 U3394 ( .A1(n2721), .A2(n3460), .ZN(n2723) );
  OR2_X1 U3395 ( .A1(n2723), .A2(n2722), .ZN(n3467) );
  OR2_X1 U3396 ( .A1(n2584), .A2(n3467), .ZN(n2725) );
  INV_X1 U3397 ( .A(REG2_REG_11__SCAN_IN), .ZN(n3450) );
  OR2_X1 U3398 ( .A1(n3230), .A2(n3450), .ZN(n2724) );
  NAND4_X1 U3399 ( .A1(n2727), .A2(n2726), .A3(n2725), .A4(n2724), .ZN(n3473)
         );
  NAND2_X1 U3400 ( .A1(n3473), .A2(n2951), .ZN(n2730) );
  XNOR2_X1 U3401 ( .A(n2728), .B(IR_REG_11__SCAN_IN), .ZN(n4591) );
  MUX2_X1 U3402 ( .A(DATAI_11_), .B(n4591), .S(n2572), .Z(n3442) );
  NAND2_X1 U3403 ( .A1(n2880), .A2(n3442), .ZN(n2729) );
  NAND2_X1 U3404 ( .A1(n2730), .A2(n2729), .ZN(n2731) );
  XNOR2_X1 U3405 ( .A(n2731), .B(n2920), .ZN(n2734) );
  NOR2_X1 U3406 ( .A1(n3459), .A2(n2987), .ZN(n2732) );
  AOI21_X1 U3407 ( .B1(n3473), .B2(n2795), .A(n2732), .ZN(n2733) );
  NAND2_X1 U3408 ( .A1(n2734), .A2(n2733), .ZN(n3455) );
  INV_X1 U3409 ( .A(n3486), .ZN(n2736) );
  AOI22_X1 U3410 ( .A1(n3543), .A2(n2795), .B1(n2951), .B2(n3029), .ZN(n3484)
         );
  NAND2_X1 U3411 ( .A1(n2684), .A2(REG2_REG_13__SCAN_IN), .ZN(n2742) );
  INV_X1 U3412 ( .A(REG0_REG_13__SCAN_IN), .ZN(n4372) );
  OR2_X1 U3413 ( .A1(n2566), .A2(n4372), .ZN(n2741) );
  INV_X1 U3414 ( .A(REG1_REG_13__SCAN_IN), .ZN(n4321) );
  OR2_X1 U3415 ( .A1(n2601), .A2(n4321), .ZN(n2740) );
  NOR2_X1 U3416 ( .A1(n2737), .A2(REG3_REG_13__SCAN_IN), .ZN(n2738) );
  OR2_X1 U3417 ( .A1(n2766), .A2(n2738), .ZN(n3566) );
  OR2_X1 U3418 ( .A1(n2584), .A2(n3566), .ZN(n2739) );
  NAND2_X1 U3419 ( .A1(n4203), .A2(n2951), .ZN(n2747) );
  OR2_X1 U3420 ( .A1(n2744), .A2(n2743), .ZN(n2745) );
  XNOR2_X1 U3421 ( .A(n2745), .B(IR_REG_13__SCAN_IN), .ZN(n4499) );
  MUX2_X1 U3422 ( .A(DATAI_13_), .B(n4499), .S(n2572), .Z(n3093) );
  NAND2_X1 U3423 ( .A1(n2880), .A2(n3093), .ZN(n2746) );
  NAND2_X1 U3424 ( .A1(n2747), .A2(n2746), .ZN(n2748) );
  XNOR2_X1 U3425 ( .A(n2748), .B(n2920), .ZN(n2753) );
  INV_X1 U3426 ( .A(n2753), .ZN(n2751) );
  INV_X1 U3427 ( .A(n3093), .ZN(n3558) );
  NOR2_X1 U3428 ( .A1(n3558), .A2(n2987), .ZN(n2749) );
  AOI21_X1 U3429 ( .B1(n4203), .B2(n2795), .A(n2749), .ZN(n2752) );
  INV_X1 U3430 ( .A(n2752), .ZN(n2750) );
  NAND2_X1 U3431 ( .A1(n2751), .A2(n2750), .ZN(n3553) );
  AND2_X1 U3432 ( .A1(n2753), .A2(n2752), .ZN(n3554) );
  AOI21_X1 U3433 ( .B1(n3552), .B2(n3553), .A(n3554), .ZN(n3584) );
  NAND2_X1 U3434 ( .A1(n2991), .A2(REG0_REG_14__SCAN_IN), .ZN(n2757) );
  INV_X1 U3435 ( .A(REG1_REG_14__SCAN_IN), .ZN(n4508) );
  OR2_X1 U3436 ( .A1(n2601), .A2(n4508), .ZN(n2756) );
  XNOR2_X1 U3437 ( .A(n2766), .B(REG3_REG_14__SCAN_IN), .ZN(n4214) );
  OR2_X1 U3438 ( .A1(n2584), .A2(n4214), .ZN(n2755) );
  INV_X1 U3439 ( .A(REG2_REG_14__SCAN_IN), .ZN(n4215) );
  OR2_X1 U3440 ( .A1(n3230), .A2(n4215), .ZN(n2754) );
  NAND4_X1 U3441 ( .A1(n2757), .A2(n2756), .A3(n2755), .A4(n2754), .ZN(n3904)
         );
  NAND2_X1 U3442 ( .A1(n2758), .A2(IR_REG_31__SCAN_IN), .ZN(n2759) );
  XNOR2_X1 U3443 ( .A(n2759), .B(IR_REG_14__SCAN_IN), .ZN(n4512) );
  MUX2_X1 U3444 ( .A(DATAI_14_), .B(n4512), .S(n2572), .Z(n4210) );
  AOI22_X1 U3445 ( .A1(n3904), .A2(n2951), .B1(n2880), .B2(n4210), .ZN(n2760)
         );
  XOR2_X1 U3446 ( .A(n2947), .B(n2760), .Z(n3582) );
  INV_X1 U3447 ( .A(n3904), .ZN(n3731) );
  INV_X1 U3448 ( .A(n2795), .ZN(n2935) );
  OAI22_X1 U3449 ( .A1(n3731), .A2(n2935), .B1(n2987), .B2(n4201), .ZN(n3581)
         );
  OAI21_X1 U3450 ( .B1(n3584), .B2(n3582), .A(n3581), .ZN(n2762) );
  NAND2_X1 U3451 ( .A1(n3584), .A2(n3582), .ZN(n2761) );
  NAND2_X1 U3452 ( .A1(n2762), .A2(n2761), .ZN(n2779) );
  INV_X1 U3453 ( .A(n2779), .ZN(n2775) );
  INV_X1 U3454 ( .A(REG0_REG_15__SCAN_IN), .ZN(n4892) );
  OR2_X1 U3455 ( .A1(n2566), .A2(n4892), .ZN(n2771) );
  INV_X1 U3456 ( .A(REG1_REG_15__SCAN_IN), .ZN(n4313) );
  OR2_X1 U3457 ( .A1(n2601), .A2(n4313), .ZN(n2770) );
  NAND2_X1 U34580 ( .A1(n2766), .A2(REG3_REG_14__SCAN_IN), .ZN(n2764) );
  INV_X1 U34590 ( .A(REG3_REG_15__SCAN_IN), .ZN(n2763) );
  NAND2_X1 U3460 ( .A1(n2764), .A2(n2763), .ZN(n2767) );
  NAND2_X1 U3461 ( .A1(n2767), .A2(n2780), .ZN(n3740) );
  OR2_X1 U3462 ( .A1(n2584), .A2(n3740), .ZN(n2769) );
  INV_X1 U3463 ( .A(REG2_REG_15__SCAN_IN), .ZN(n3950) );
  OR2_X1 U3464 ( .A1(n3230), .A2(n3950), .ZN(n2768) );
  NAND4_X1 U3465 ( .A1(n2771), .A2(n2770), .A3(n2769), .A4(n2768), .ZN(n4187)
         );
  OR2_X1 U3466 ( .A1(n2758), .A2(IR_REG_14__SCAN_IN), .ZN(n2772) );
  NAND2_X1 U34670 ( .A1(n2772), .A2(IR_REG_31__SCAN_IN), .ZN(n2787) );
  XNOR2_X1 U3468 ( .A(n2787), .B(IR_REG_15__SCAN_IN), .ZN(n3951) );
  MUX2_X1 U34690 ( .A(DATAI_15_), .B(n3951), .S(n2572), .Z(n3034) );
  AOI22_X1 U3470 ( .A1(n4187), .A2(n2951), .B1(n2880), .B2(n3034), .ZN(n2773)
         );
  XOR2_X1 U34710 ( .A(n2947), .B(n2773), .Z(n2778) );
  NAND2_X1 U3472 ( .A1(n2775), .A2(n2774), .ZN(n3727) );
  NAND2_X1 U34730 ( .A1(n4187), .A2(n2795), .ZN(n2777) );
  NAND2_X1 U3474 ( .A1(n2951), .A2(n3034), .ZN(n2776) );
  NAND2_X1 U34750 ( .A1(n2777), .A2(n2776), .ZN(n4401) );
  NAND2_X1 U3476 ( .A1(n3727), .A2(n4401), .ZN(n2797) );
  NAND2_X1 U34770 ( .A1(n2779), .A2(n2778), .ZN(n3728) );
  NAND2_X1 U3478 ( .A1(n2780), .A2(n4396), .ZN(n2781) );
  NAND2_X1 U34790 ( .A1(n2804), .A2(n2781), .ZN(n4409) );
  OR2_X1 U3480 ( .A1(n2584), .A2(n4409), .ZN(n2785) );
  INV_X1 U34810 ( .A(REG1_REG_16__SCAN_IN), .ZN(n4528) );
  OR2_X1 U3482 ( .A1(n2601), .A2(n4528), .ZN(n2784) );
  INV_X1 U34830 ( .A(REG2_REG_16__SCAN_IN), .ZN(n4193) );
  OR2_X1 U3484 ( .A1(n3230), .A2(n4193), .ZN(n2783) );
  INV_X1 U34850 ( .A(REG0_REG_16__SCAN_IN), .ZN(n4807) );
  OR2_X1 U3486 ( .A1(n2566), .A2(n4807), .ZN(n2782) );
  NAND2_X1 U34870 ( .A1(n4169), .A2(n2951), .ZN(n2793) );
  NAND2_X1 U3488 ( .A1(n2787), .A2(n2786), .ZN(n2788) );
  NAND2_X1 U34890 ( .A1(n2788), .A2(IR_REG_31__SCAN_IN), .ZN(n2790) );
  XNOR2_X1 U3490 ( .A(n2790), .B(n2789), .ZN(n4587) );
  INV_X1 U34910 ( .A(n4587), .ZN(n2791) );
  MUX2_X1 U3492 ( .A(DATAI_16_), .B(n2791), .S(n2572), .Z(n4191) );
  NAND2_X1 U34930 ( .A1(n2880), .A2(n4191), .ZN(n2792) );
  NAND2_X1 U3494 ( .A1(n2793), .A2(n2792), .ZN(n2794) );
  XNOR2_X1 U34950 ( .A(n2794), .B(n2947), .ZN(n2798) );
  AOI22_X1 U3496 ( .A1(n4169), .A2(n2795), .B1(n2951), .B2(n4191), .ZN(n2799)
         );
  XNOR2_X1 U34970 ( .A(n2798), .B(n2799), .ZN(n4403) );
  INV_X1 U3498 ( .A(REG3_REG_17__SCAN_IN), .ZN(n2803) );
  NAND2_X1 U34990 ( .A1(n2804), .A2(n2803), .ZN(n2805) );
  NAND2_X1 U3500 ( .A1(n2815), .A2(n2805), .ZN(n4176) );
  OR2_X1 U35010 ( .A1(n2584), .A2(n4176), .ZN(n2809) );
  INV_X1 U3502 ( .A(REG1_REG_17__SCAN_IN), .ZN(n4304) );
  OR2_X1 U35030 ( .A1(n2601), .A2(n4304), .ZN(n2808) );
  INV_X1 U3504 ( .A(REG2_REG_17__SCAN_IN), .ZN(n4829) );
  OR2_X1 U35050 ( .A1(n3230), .A2(n4829), .ZN(n2807) );
  INV_X1 U35060 ( .A(REG0_REG_17__SCAN_IN), .ZN(n4932) );
  OR2_X1 U35070 ( .A1(n2566), .A2(n4932), .ZN(n2806) );
  NAND4_X1 U35080 ( .A1(n2809), .A2(n2808), .A3(n2807), .A4(n2806), .ZN(n4151)
         );
  NAND2_X1 U35090 ( .A1(n2275), .A2(IR_REG_31__SCAN_IN), .ZN(n2810) );
  MUX2_X1 U35100 ( .A(IR_REG_31__SCAN_IN), .B(n2810), .S(IR_REG_17__SCAN_IN), 
        .Z(n2811) );
  NAND2_X1 U35110 ( .A1(n2811), .A2(n2508), .ZN(n4586) );
  MUX2_X1 U35120 ( .A(DATAI_17_), .B(n3954), .S(n2572), .Z(n3094) );
  AOI22_X1 U35130 ( .A1(n4151), .A2(n2951), .B1(n2880), .B2(n3094), .ZN(n2812)
         );
  XOR2_X1 U35140 ( .A(n2947), .B(n2812), .Z(n3665) );
  INV_X1 U35150 ( .A(n4151), .ZN(n4398) );
  OAI22_X1 U35160 ( .A1(n4398), .A2(n2935), .B1(n2987), .B2(n4173), .ZN(n3666)
         );
  NAND2_X1 U35170 ( .A1(n3665), .A2(n3666), .ZN(n2813) );
  NAND2_X1 U35180 ( .A1(n2991), .A2(REG0_REG_18__SCAN_IN), .ZN(n2820) );
  INV_X1 U35190 ( .A(REG1_REG_18__SCAN_IN), .ZN(n2814) );
  OR2_X1 U35200 ( .A1(n2601), .A2(n2814), .ZN(n2819) );
  NAND2_X1 U35210 ( .A1(n2815), .A2(n4967), .ZN(n2816) );
  NAND2_X1 U35220 ( .A1(n2831), .A2(n2816), .ZN(n4160) );
  OR2_X1 U35230 ( .A1(n2584), .A2(n4160), .ZN(n2818) );
  INV_X1 U35240 ( .A(REG2_REG_18__SCAN_IN), .ZN(n4161) );
  OR2_X1 U35250 ( .A1(n3230), .A2(n4161), .ZN(n2817) );
  NAND2_X1 U35260 ( .A1(n4133), .A2(n2951), .ZN(n2824) );
  NAND2_X1 U35270 ( .A1(n2508), .A2(IR_REG_31__SCAN_IN), .ZN(n2821) );
  MUX2_X1 U35280 ( .A(IR_REG_31__SCAN_IN), .B(n2821), .S(IR_REG_18__SCAN_IN), 
        .Z(n2822) );
  AND2_X1 U35290 ( .A1(n2822), .A2(n2247), .ZN(n4554) );
  MUX2_X1 U35300 ( .A(DATAI_18_), .B(n4554), .S(n2572), .Z(n4155) );
  NAND2_X1 U35310 ( .A1(n2880), .A2(n4155), .ZN(n2823) );
  NAND2_X1 U35320 ( .A1(n2824), .A2(n2823), .ZN(n2825) );
  XNOR2_X1 U35330 ( .A(n2825), .B(n2920), .ZN(n2828) );
  INV_X1 U35340 ( .A(n4155), .ZN(n4145) );
  NOR2_X1 U35350 ( .A1(n4145), .A2(n2987), .ZN(n2826) );
  AOI21_X1 U35360 ( .B1(n4133), .B2(n2795), .A(n2826), .ZN(n2827) );
  NAND2_X1 U35370 ( .A1(n2828), .A2(n2827), .ZN(n3707) );
  NAND2_X1 U35380 ( .A1(n2991), .A2(REG0_REG_19__SCAN_IN), .ZN(n2836) );
  INV_X1 U35390 ( .A(REG1_REG_19__SCAN_IN), .ZN(n4296) );
  OR2_X1 U35400 ( .A1(n2601), .A2(n4296), .ZN(n2835) );
  INV_X1 U35410 ( .A(REG3_REG_19__SCAN_IN), .ZN(n2830) );
  NAND2_X1 U35420 ( .A1(n2831), .A2(n2830), .ZN(n2832) );
  NAND2_X1 U35430 ( .A1(n2844), .A2(n2832), .ZN(n4139) );
  OR2_X1 U35440 ( .A1(n2584), .A2(n4139), .ZN(n2834) );
  INV_X1 U35450 ( .A(REG2_REG_19__SCAN_IN), .ZN(n4140) );
  OR2_X1 U35460 ( .A1(n3230), .A2(n4140), .ZN(n2833) );
  NAND2_X1 U35470 ( .A1(n4112), .A2(n2951), .ZN(n2838) );
  INV_X1 U35480 ( .A(n3959), .ZN(n4380) );
  MUX2_X1 U35490 ( .A(DATAI_19_), .B(n4380), .S(n2572), .Z(n3095) );
  NAND2_X1 U35500 ( .A1(n2880), .A2(n3095), .ZN(n2837) );
  NAND2_X1 U35510 ( .A1(n2838), .A2(n2837), .ZN(n2839) );
  XNOR2_X1 U35520 ( .A(n2839), .B(n2947), .ZN(n2840) );
  AOI22_X1 U35530 ( .A1(n4112), .A2(n2795), .B1(n2951), .B2(n3095), .ZN(n2841)
         );
  XNOR2_X1 U35540 ( .A(n2840), .B(n2841), .ZN(n3636) );
  NAND2_X1 U35550 ( .A1(n3635), .A2(n3636), .ZN(n3634) );
  NAND2_X1 U35560 ( .A1(n3634), .A2(n2843), .ZN(n3645) );
  NAND2_X1 U35570 ( .A1(n2991), .A2(REG0_REG_20__SCAN_IN), .ZN(n2849) );
  INV_X1 U35580 ( .A(REG1_REG_20__SCAN_IN), .ZN(n4935) );
  OR2_X1 U35590 ( .A1(n2601), .A2(n4935), .ZN(n2848) );
  INV_X1 U35600 ( .A(REG3_REG_20__SCAN_IN), .ZN(n4867) );
  NAND2_X1 U35610 ( .A1(n2844), .A2(n4867), .ZN(n2845) );
  NAND2_X1 U35620 ( .A1(n2865), .A2(n2845), .ZN(n4117) );
  OR2_X1 U35630 ( .A1(n2584), .A2(n4117), .ZN(n2847) );
  INV_X1 U35640 ( .A(REG2_REG_20__SCAN_IN), .ZN(n4118) );
  OR2_X1 U35650 ( .A1(n3230), .A2(n4118), .ZN(n2846) );
  NAND4_X1 U35660 ( .A1(n2849), .A2(n2848), .A3(n2847), .A4(n2846), .ZN(n4091)
         );
  NAND2_X1 U35670 ( .A1(n4091), .A2(n2571), .ZN(n2851) );
  OR2_X1 U35680 ( .A1(n2949), .A2(n4114), .ZN(n2850) );
  NAND2_X1 U35690 ( .A1(n2851), .A2(n2850), .ZN(n2852) );
  XNOR2_X1 U35700 ( .A(n2852), .B(n2920), .ZN(n2855) );
  NOR2_X1 U35710 ( .A1(n2987), .A2(n4114), .ZN(n2853) );
  AOI21_X1 U35720 ( .B1(n4091), .B2(n2795), .A(n2853), .ZN(n2854) );
  NAND2_X1 U35730 ( .A1(n3645), .A2(n3688), .ZN(n3686) );
  NAND2_X1 U35740 ( .A1(n2855), .A2(n2854), .ZN(n3687) );
  INV_X1 U35750 ( .A(REG3_REG_21__SCAN_IN), .ZN(n3649) );
  XNOR2_X1 U35760 ( .A(n2865), .B(n3649), .ZN(n4097) );
  OR2_X1 U35770 ( .A1(n4097), .A2(n2584), .ZN(n2859) );
  INV_X1 U35780 ( .A(REG0_REG_21__SCAN_IN), .ZN(n4348) );
  OR2_X1 U35790 ( .A1(n2566), .A2(n4348), .ZN(n2858) );
  INV_X1 U35800 ( .A(REG1_REG_21__SCAN_IN), .ZN(n4288) );
  OR2_X1 U35810 ( .A1(n2601), .A2(n4288), .ZN(n2857) );
  INV_X1 U3582 ( .A(REG2_REG_21__SCAN_IN), .ZN(n4831) );
  OR2_X1 U3583 ( .A1(n3230), .A2(n4831), .ZN(n2856) );
  NAND4_X1 U3584 ( .A1(n2859), .A2(n2858), .A3(n2857), .A4(n2856), .ZN(n4073)
         );
  NOR2_X1 U3585 ( .A1(n2949), .A2(n4094), .ZN(n2860) );
  AOI21_X1 U3586 ( .B1(n4073), .B2(n2571), .A(n2860), .ZN(n2861) );
  XNOR2_X1 U3587 ( .A(n2861), .B(n2947), .ZN(n2864) );
  NOR2_X1 U3588 ( .A1(n2987), .A2(n4094), .ZN(n2862) );
  AOI21_X1 U3589 ( .B1(n4073), .B2(n2795), .A(n2862), .ZN(n2863) );
  OR2_X1 U3590 ( .A1(n2864), .A2(n2863), .ZN(n3643) );
  NAND2_X1 U3591 ( .A1(n2563), .A2(REG1_REG_22__SCAN_IN), .ZN(n2872) );
  INV_X1 U3592 ( .A(REG0_REG_22__SCAN_IN), .ZN(n4934) );
  OR2_X1 U3593 ( .A1(n2566), .A2(n4934), .ZN(n2871) );
  INV_X1 U3594 ( .A(REG3_REG_22__SCAN_IN), .ZN(n3698) );
  OAI21_X1 U3595 ( .B1(n2865), .B2(n3649), .A(n3698), .ZN(n2868) );
  AND2_X1 U3596 ( .A1(REG3_REG_21__SCAN_IN), .A2(REG3_REG_22__SCAN_IN), .ZN(
        n2866) );
  NAND2_X1 U3597 ( .A1(n2868), .A2(n2875), .ZN(n4078) );
  OR2_X1 U3598 ( .A1(n2584), .A2(n4078), .ZN(n2870) );
  INV_X1 U3599 ( .A(REG2_REG_22__SCAN_IN), .ZN(n4079) );
  OR2_X1 U3600 ( .A1(n3230), .A2(n4079), .ZN(n2869) );
  NAND2_X1 U3601 ( .A1(n3741), .A2(DATAI_22_), .ZN(n4081) );
  OAI22_X1 U3602 ( .A1(n4089), .A2(n2987), .B1(n2949), .B2(n4081), .ZN(n2873)
         );
  XNOR2_X1 U3603 ( .A(n2873), .B(n2947), .ZN(n2884) );
  OAI22_X1 U3604 ( .A1(n4089), .A2(n2935), .B1(n2987), .B2(n4081), .ZN(n2883)
         );
  XNOR2_X1 U3605 ( .A(n2884), .B(n2883), .ZN(n3697) );
  INV_X1 U3606 ( .A(REG3_REG_23__SCAN_IN), .ZN(n3629) );
  NAND2_X1 U3607 ( .A1(n2875), .A2(n3629), .ZN(n2876) );
  NAND2_X1 U3608 ( .A1(n2902), .A2(n2876), .ZN(n4063) );
  NOR2_X1 U3609 ( .A1(n4063), .A2(n2584), .ZN(n2879) );
  INV_X1 U3610 ( .A(REG1_REG_23__SCAN_IN), .ZN(n4942) );
  INV_X1 U3611 ( .A(REG0_REG_23__SCAN_IN), .ZN(n4343) );
  OAI22_X1 U3612 ( .A1(n2601), .A2(n4942), .B1(n2566), .B2(n4343), .ZN(n2878)
         );
  INV_X1 U3613 ( .A(REG2_REG_23__SCAN_IN), .ZN(n4064) );
  NOR2_X1 U3614 ( .A1(n3230), .A2(n4064), .ZN(n2877) );
  AOI22_X1 U3615 ( .A1(n4072), .A2(n2951), .B1(n2880), .B2(n4054), .ZN(n2881)
         );
  XNOR2_X1 U3616 ( .A(n2881), .B(n2947), .ZN(n2887) );
  INV_X1 U3617 ( .A(n4054), .ZN(n4061) );
  NOR2_X1 U3618 ( .A1(n2987), .A2(n4061), .ZN(n2882) );
  AOI21_X1 U3619 ( .B1(n4072), .B2(n2795), .A(n2882), .ZN(n2886) );
  XNOR2_X1 U3620 ( .A(n2887), .B(n2886), .ZN(n3625) );
  NOR2_X1 U3621 ( .A1(n2884), .A2(n2883), .ZN(n3626) );
  NOR2_X1 U3622 ( .A1(n3625), .A2(n3626), .ZN(n2885) );
  NAND2_X2 U3623 ( .A1(n3624), .A2(n2885), .ZN(n3627) );
  OR2_X1 U3624 ( .A1(n2887), .A2(n2886), .ZN(n2897) );
  NAND2_X1 U3625 ( .A1(n3627), .A2(n2897), .ZN(n2895) );
  INV_X1 U3626 ( .A(REG1_REG_24__SCAN_IN), .ZN(n4941) );
  NAND2_X1 U3627 ( .A1(n2991), .A2(REG0_REG_24__SCAN_IN), .ZN(n2889) );
  NAND2_X1 U3628 ( .A1(n2684), .A2(REG2_REG_24__SCAN_IN), .ZN(n2888) );
  OAI211_X1 U3629 ( .C1(n2601), .C2(n4941), .A(n2889), .B(n2888), .ZN(n2890)
         );
  INV_X1 U3630 ( .A(n2890), .ZN(n2892) );
  XNOR2_X1 U3631 ( .A(n2902), .B(REG3_REG_24__SCAN_IN), .ZN(n4040) );
  NAND2_X1 U3632 ( .A1(n4040), .A2(n2996), .ZN(n2891) );
  NOR2_X1 U3633 ( .A1(n2944), .A2(n3679), .ZN(n2893) );
  AOI21_X1 U3634 ( .B1(n4016), .B2(n2795), .A(n2893), .ZN(n2896) );
  INV_X1 U3635 ( .A(n2896), .ZN(n2894) );
  NAND2_X1 U3636 ( .A1(n2895), .A2(n2894), .ZN(n3675) );
  OAI22_X1 U3637 ( .A1(n4059), .A2(n2987), .B1(n2949), .B2(n3679), .ZN(n2899)
         );
  XNOR2_X1 U3638 ( .A(n2899), .B(n2947), .ZN(n3676) );
  NAND2_X1 U3639 ( .A1(n3674), .A2(n3676), .ZN(n2900) );
  INV_X1 U3640 ( .A(REG2_REG_25__SCAN_IN), .ZN(n2906) );
  NAND2_X1 U3641 ( .A1(REG3_REG_24__SCAN_IN), .A2(REG3_REG_25__SCAN_IN), .ZN(
        n2901) );
  INV_X1 U3642 ( .A(REG3_REG_24__SCAN_IN), .ZN(n3680) );
  INV_X1 U3643 ( .A(REG3_REG_25__SCAN_IN), .ZN(n3658) );
  OAI21_X1 U3644 ( .B1(n2902), .B2(n3680), .A(n3658), .ZN(n2903) );
  AND2_X1 U3645 ( .A1(n2914), .A2(n2903), .ZN(n4022) );
  NAND2_X1 U3646 ( .A1(n4022), .A2(n2996), .ZN(n2905) );
  AOI22_X1 U3647 ( .A1(n2563), .A2(REG1_REG_25__SCAN_IN), .B1(n2991), .B2(
        REG0_REG_25__SCAN_IN), .ZN(n2904) );
  NAND2_X1 U3648 ( .A1(n3232), .A2(n2951), .ZN(n2908) );
  NAND2_X1 U3649 ( .A1(n3741), .A2(DATAI_25_), .ZN(n4021) );
  OR2_X1 U3650 ( .A1(n2949), .A2(n4021), .ZN(n2907) );
  NAND2_X1 U3651 ( .A1(n2908), .A2(n2907), .ZN(n2909) );
  XNOR2_X1 U3652 ( .A(n2909), .B(n2920), .ZN(n2912) );
  NOR2_X1 U3653 ( .A1(n2987), .A2(n4021), .ZN(n2910) );
  AOI21_X1 U3654 ( .B1(n3232), .B2(n2795), .A(n2910), .ZN(n2911) );
  NAND2_X1 U3655 ( .A1(n2912), .A2(n2911), .ZN(n3654) );
  INV_X1 U3656 ( .A(REG2_REG_26__SCAN_IN), .ZN(n4005) );
  INV_X1 U3657 ( .A(n2914), .ZN(n2913) );
  NAND2_X1 U3658 ( .A1(n2913), .A2(REG3_REG_26__SCAN_IN), .ZN(n2927) );
  INV_X1 U3659 ( .A(REG3_REG_26__SCAN_IN), .ZN(n4852) );
  NAND2_X1 U3660 ( .A1(n2914), .A2(n4852), .ZN(n2915) );
  NAND2_X1 U3661 ( .A1(n2927), .A2(n2915), .ZN(n4004) );
  OR2_X1 U3662 ( .A1(n4004), .A2(n2584), .ZN(n2917) );
  AOI22_X1 U3663 ( .A1(n2563), .A2(REG1_REG_26__SCAN_IN), .B1(n2991), .B2(
        REG0_REG_26__SCAN_IN), .ZN(n2916) );
  OAI211_X1 U3664 ( .C1(n3230), .C2(n4005), .A(n2917), .B(n2916), .ZN(n3996)
         );
  NAND2_X1 U3665 ( .A1(n3996), .A2(n2571), .ZN(n2919) );
  NAND2_X1 U3666 ( .A1(n3741), .A2(DATAI_26_), .ZN(n3721) );
  OR2_X1 U3667 ( .A1(n2949), .A2(n3721), .ZN(n2918) );
  NAND2_X1 U3668 ( .A1(n2919), .A2(n2918), .ZN(n2921) );
  XNOR2_X1 U3669 ( .A(n2921), .B(n2920), .ZN(n2924) );
  NOR2_X1 U3670 ( .A1(n2987), .A2(n3721), .ZN(n2922) );
  AOI21_X1 U3671 ( .B1(n3996), .B2(n2795), .A(n2922), .ZN(n2923) );
  OR2_X1 U3672 ( .A1(n2924), .A2(n2923), .ZN(n3714) );
  AND2_X1 U3673 ( .A1(n2924), .A2(n2923), .ZN(n3715) );
  INV_X1 U3674 ( .A(n2927), .ZN(n2925) );
  NAND2_X1 U3675 ( .A1(n2925), .A2(REG3_REG_27__SCAN_IN), .ZN(n2937) );
  INV_X1 U3676 ( .A(REG3_REG_27__SCAN_IN), .ZN(n2926) );
  NAND2_X1 U3677 ( .A1(n2927), .A2(n2926), .ZN(n2928) );
  NAND2_X1 U3678 ( .A1(n2937), .A2(n2928), .ZN(n3987) );
  OR2_X1 U3679 ( .A1(n3987), .A2(n2584), .ZN(n2934) );
  INV_X1 U3680 ( .A(REG0_REG_27__SCAN_IN), .ZN(n2931) );
  NAND2_X1 U3681 ( .A1(n2684), .A2(REG2_REG_27__SCAN_IN), .ZN(n2930) );
  NAND2_X1 U3682 ( .A1(n2563), .A2(REG1_REG_27__SCAN_IN), .ZN(n2929) );
  OAI211_X1 U3683 ( .C1(n2566), .C2(n2931), .A(n2930), .B(n2929), .ZN(n2932)
         );
  INV_X1 U3684 ( .A(n2932), .ZN(n2933) );
  NAND2_X1 U3685 ( .A1(n3741), .A2(DATAI_27_), .ZN(n3616) );
  OAI22_X1 U3686 ( .A1(n3779), .A2(n2935), .B1(n2987), .B2(n3616), .ZN(n2976)
         );
  OAI22_X1 U3687 ( .A1(n3779), .A2(n2987), .B1(n3616), .B2(n2949), .ZN(n2936)
         );
  XNOR2_X1 U3688 ( .A(n2936), .B(n2947), .ZN(n2977) );
  XOR2_X1 U3689 ( .A(n2976), .B(n2977), .Z(n3614) );
  INV_X1 U3690 ( .A(REG3_REG_28__SCAN_IN), .ZN(n3003) );
  NAND2_X1 U3691 ( .A1(n2937), .A2(n3003), .ZN(n2938) );
  NAND2_X1 U3692 ( .A1(n3976), .A2(n2996), .ZN(n2943) );
  INV_X1 U3693 ( .A(REG1_REG_28__SCAN_IN), .ZN(n4819) );
  NAND2_X1 U3694 ( .A1(n2684), .A2(REG2_REG_28__SCAN_IN), .ZN(n2940) );
  INV_X1 U3695 ( .A(REG0_REG_28__SCAN_IN), .ZN(n4945) );
  OR2_X1 U3696 ( .A1(n2566), .A2(n4945), .ZN(n2939) );
  OAI211_X1 U3697 ( .C1(n2601), .C2(n4819), .A(n2940), .B(n2939), .ZN(n2941)
         );
  INV_X1 U3698 ( .A(n2941), .ZN(n2942) );
  NAND2_X1 U3699 ( .A1(n3990), .A2(n2795), .ZN(n2946) );
  NAND2_X1 U3700 ( .A1(n3741), .A2(DATAI_28_), .ZN(n3968) );
  OR2_X1 U3701 ( .A1(n2944), .A2(n3968), .ZN(n2945) );
  NAND2_X1 U3702 ( .A1(n2946), .A2(n2945), .ZN(n2948) );
  XNOR2_X1 U3703 ( .A(n2948), .B(n2947), .ZN(n2953) );
  NOR2_X1 U3704 ( .A1(n2949), .A2(n3968), .ZN(n2950) );
  AOI21_X1 U3705 ( .B1(n3990), .B2(n2951), .A(n2950), .ZN(n2952) );
  XNOR2_X1 U3706 ( .A(n2953), .B(n2952), .ZN(n2979) );
  INV_X1 U3707 ( .A(n2979), .ZN(n2975) );
  NAND2_X1 U3708 ( .A1(n3106), .A2(B_REG_SCAN_IN), .ZN(n2955) );
  MUX2_X1 U3709 ( .A(n2955), .B(B_REG_SCAN_IN), .S(n2954), .Z(n2956) );
  NOR2_X1 U3710 ( .A1(D_REG_13__SCAN_IN), .A2(D_REG_11__SCAN_IN), .ZN(n2960)
         );
  NOR4_X1 U3711 ( .A1(D_REG_28__SCAN_IN), .A2(D_REG_30__SCAN_IN), .A3(
        D_REG_4__SCAN_IN), .A4(D_REG_12__SCAN_IN), .ZN(n2959) );
  NOR4_X1 U3712 ( .A1(D_REG_19__SCAN_IN), .A2(D_REG_18__SCAN_IN), .A3(
        D_REG_17__SCAN_IN), .A4(D_REG_7__SCAN_IN), .ZN(n2958) );
  NOR4_X1 U3713 ( .A1(D_REG_10__SCAN_IN), .A2(D_REG_29__SCAN_IN), .A3(
        D_REG_24__SCAN_IN), .A4(D_REG_5__SCAN_IN), .ZN(n2957) );
  NAND4_X1 U3714 ( .A1(n2960), .A2(n2959), .A3(n2958), .A4(n2957), .ZN(n2966)
         );
  NOR4_X1 U3715 ( .A1(D_REG_21__SCAN_IN), .A2(D_REG_2__SCAN_IN), .A3(
        D_REG_3__SCAN_IN), .A4(D_REG_6__SCAN_IN), .ZN(n2964) );
  NOR4_X1 U3716 ( .A1(D_REG_9__SCAN_IN), .A2(D_REG_8__SCAN_IN), .A3(
        D_REG_26__SCAN_IN), .A4(D_REG_25__SCAN_IN), .ZN(n2963) );
  NOR4_X1 U3717 ( .A1(D_REG_22__SCAN_IN), .A2(D_REG_23__SCAN_IN), .A3(
        D_REG_27__SCAN_IN), .A4(D_REG_31__SCAN_IN), .ZN(n2962) );
  NOR4_X1 U3718 ( .A1(D_REG_14__SCAN_IN), .A2(D_REG_15__SCAN_IN), .A3(
        D_REG_16__SCAN_IN), .A4(D_REG_20__SCAN_IN), .ZN(n2961) );
  NAND4_X1 U3719 ( .A1(n2964), .A2(n2963), .A3(n2962), .A4(n2961), .ZN(n2965)
         );
  NOR2_X1 U3720 ( .A1(n2966), .A2(n2965), .ZN(n2967) );
  NAND2_X1 U3721 ( .A1(n2507), .A2(n3106), .ZN(n3116) );
  INV_X1 U3722 ( .A(n2954), .ZN(n2968) );
  NAND2_X1 U3723 ( .A1(n2968), .A2(n2507), .ZN(n3114) );
  NAND3_X1 U3724 ( .A1(n3205), .A2(n3098), .A3(n3203), .ZN(n2989) );
  INV_X1 U3725 ( .A(n3202), .ZN(n2973) );
  INV_X1 U3726 ( .A(n2972), .ZN(n4568) );
  NAND2_X1 U3727 ( .A1(n3785), .A2(n4379), .ZN(n3082) );
  OAI211_X1 U3728 ( .C1(n4568), .C2(n3959), .A(n4255), .B(n3082), .ZN(n2981)
         );
  NOR2_X1 U3729 ( .A1(n2973), .A2(n2981), .ZN(n2974) );
  NAND2_X1 U3730 ( .A1(n2975), .A2(n4405), .ZN(n3016) );
  NAND2_X1 U3731 ( .A1(n2977), .A2(n2976), .ZN(n2978) );
  NAND2_X1 U3732 ( .A1(n3017), .A2(n2469), .ZN(n3015) );
  INV_X1 U3733 ( .A(n2978), .ZN(n2980) );
  NAND3_X1 U3734 ( .A1(n2980), .A2(n4405), .A3(n2975), .ZN(n3013) );
  NAND2_X1 U3735 ( .A1(n2981), .A2(n4255), .ZN(n2982) );
  NAND2_X1 U3736 ( .A1(n2989), .A2(n2982), .ZN(n2984) );
  NAND2_X1 U3737 ( .A1(n3848), .A2(n3959), .ZN(n2983) );
  NAND2_X1 U3738 ( .A1(n3121), .A2(n2983), .ZN(n3201) );
  NAND2_X1 U3739 ( .A1(n2984), .A2(n3201), .ZN(n3154) );
  NAND2_X1 U3740 ( .A1(n2544), .A2(n3120), .ZN(n2985) );
  OAI21_X1 U3741 ( .B1(n3154), .B2(n2985), .A(STATE_REG_SCAN_IN), .ZN(n2990)
         );
  INV_X1 U3742 ( .A(n3900), .ZN(n2988) );
  NAND2_X1 U3743 ( .A1(n2989), .A2(n2988), .ZN(n3152) );
  INV_X1 U3744 ( .A(n4410), .ZN(n3011) );
  INV_X1 U3745 ( .A(n3610), .ZN(n2997) );
  INV_X1 U3746 ( .A(REG2_REG_29__SCAN_IN), .ZN(n2994) );
  NAND2_X1 U3747 ( .A1(n2991), .A2(REG0_REG_29__SCAN_IN), .ZN(n2993) );
  NAND2_X1 U3748 ( .A1(n2563), .A2(REG1_REG_29__SCAN_IN), .ZN(n2992) );
  OAI211_X1 U3749 ( .C1(n2994), .C2(n3230), .A(n2993), .B(n2992), .ZN(n2995)
         );
  AOI21_X1 U3750 ( .B1(n2997), .B2(n2996), .A(n2995), .ZN(n3969) );
  NAND2_X1 U3751 ( .A1(n2248), .A2(IR_REG_31__SCAN_IN), .ZN(n2998) );
  MUX2_X1 U3752 ( .A(IR_REG_31__SCAN_IN), .B(n2998), .S(IR_REG_28__SCAN_IN), 
        .Z(n3001) );
  INV_X1 U3753 ( .A(n2999), .ZN(n3000) );
  NAND2_X1 U3754 ( .A1(n3001), .A2(n3000), .ZN(n3083) );
  INV_X1 U3755 ( .A(n3083), .ZN(n4377) );
  NOR2_X1 U3756 ( .A1(n3900), .A2(n4377), .ZN(n3002) );
  INV_X2 U3757 ( .A(n3618), .ZN(n3720) );
  OAI22_X1 U3758 ( .A1(n3969), .A2(n3720), .B1(STATE_REG_SCAN_IN), .B2(n3003), 
        .ZN(n3010) );
  AND2_X1 U3759 ( .A1(n3202), .A2(n4055), .ZN(n3004) );
  NAND2_X1 U3760 ( .A1(n3008), .A2(n3004), .ZN(n3006) );
  OR2_X1 U3761 ( .A1(n2542), .A2(n3959), .ZN(n4576) );
  INV_X1 U3762 ( .A(n4576), .ZN(n3005) );
  NAND2_X1 U3763 ( .A1(n3005), .A2(n3897), .ZN(n4614) );
  NOR2_X1 U3764 ( .A1(n4614), .A2(n3785), .ZN(n3087) );
  AND2_X2 U3765 ( .A1(n3006), .A2(n4213), .ZN(n3733) );
  NOR2_X1 U3766 ( .A1(n3900), .A2(n3083), .ZN(n3007) );
  NAND2_X2 U3767 ( .A1(n3008), .A2(n3007), .ZN(n3722) );
  OAI22_X1 U3768 ( .A1(n3733), .A2(n3968), .B1(n3779), .B2(n3722), .ZN(n3009)
         );
  AOI211_X1 U3769 ( .C1(n3976), .C2(n3011), .A(n3010), .B(n3009), .ZN(n3012)
         );
  OAI211_X1 U3770 ( .C1(n3017), .C2(n3016), .A(n3015), .B(n3014), .ZN(U3217)
         );
  INV_X1 U3771 ( .A(REG1_REG_26__SCAN_IN), .ZN(n3092) );
  INV_X1 U3772 ( .A(n3905), .ZN(n3462) );
  INV_X1 U3773 ( .A(n3906), .ZN(n3414) );
  INV_X1 U3774 ( .A(n3384), .ZN(n3395) );
  NAND2_X1 U3775 ( .A1(n3018), .A2(n3253), .ZN(n3783) );
  NAND2_X1 U3776 ( .A1(n3787), .A2(n3783), .ZN(n3053) );
  NAND2_X1 U3777 ( .A1(n3053), .A2(n3241), .ZN(n3240) );
  NAND2_X1 U3778 ( .A1(n3018), .A2(n3243), .ZN(n3019) );
  NAND2_X1 U3779 ( .A1(n2576), .A2(n4232), .ZN(n3791) );
  NAND2_X1 U3780 ( .A1(n3788), .A2(n3791), .ZN(n4224) );
  OR2_X1 U3781 ( .A1(n2576), .A2(n4239), .ZN(n3020) );
  NOR2_X1 U3782 ( .A1(n4229), .A2(n3220), .ZN(n3021) );
  INV_X1 U3783 ( .A(n4229), .ZN(n3266) );
  INV_X1 U3784 ( .A(n3220), .ZN(n3173) );
  OR2_X1 U3785 ( .A1(n3909), .A2(n3267), .ZN(n3794) );
  NAND2_X1 U3786 ( .A1(n3909), .A2(n3267), .ZN(n3798) );
  NAND2_X1 U3787 ( .A1(n3794), .A2(n3798), .ZN(n3193) );
  INV_X1 U3788 ( .A(n3196), .ZN(n3336) );
  OR2_X1 U3789 ( .A1(n3908), .A2(n3345), .ZN(n3022) );
  INV_X1 U3790 ( .A(n3908), .ZN(n3312) );
  OR2_X1 U3791 ( .A1(n3366), .A2(n3310), .ZN(n3058) );
  NAND2_X1 U3792 ( .A1(n3366), .A2(n3310), .ZN(n3805) );
  NAND2_X1 U3793 ( .A1(n3058), .A2(n3805), .ZN(n3296) );
  NAND2_X1 U3794 ( .A1(n3301), .A2(n3296), .ZN(n3024) );
  NAND2_X1 U3795 ( .A1(n3366), .A2(n3302), .ZN(n3023) );
  NAND2_X1 U3796 ( .A1(n3024), .A2(n3023), .ZN(n3372) );
  INV_X1 U3797 ( .A(n3907), .ZN(n3394) );
  NAND2_X1 U3798 ( .A1(n3028), .A2(n3027), .ZN(n3447) );
  OR2_X1 U3799 ( .A1(n3473), .A2(n3459), .ZN(n3468) );
  NAND2_X1 U3800 ( .A1(n3473), .A2(n3459), .ZN(n3470) );
  NAND2_X1 U3801 ( .A1(n3468), .A2(n3470), .ZN(n3446) );
  INV_X1 U3802 ( .A(n3473), .ZN(n3489) );
  INV_X1 U3803 ( .A(n3543), .ZN(n3561) );
  NAND2_X1 U3804 ( .A1(n3561), .A2(n3488), .ZN(n3030) );
  NOR2_X1 U3805 ( .A1(n4203), .A2(n3093), .ZN(n3533) );
  AND2_X1 U3806 ( .A1(n4203), .A2(n3093), .ZN(n3567) );
  INV_X1 U3807 ( .A(n3567), .ZN(n3032) );
  NAND2_X1 U3808 ( .A1(n3904), .A2(n4201), .ZN(n3811) );
  INV_X1 U3809 ( .A(n4187), .ZN(n4394) );
  NOR2_X1 U3810 ( .A1(n4394), .A2(n3732), .ZN(n3035) );
  OR2_X1 U3811 ( .A1(n3904), .A2(n4210), .ZN(n3569) );
  OAI22_X1 U3812 ( .A1(n3035), .A2(n3569), .B1(n3034), .B2(n4187), .ZN(n3036)
         );
  OR2_X1 U3813 ( .A1(n4169), .A2(n4395), .ZN(n3863) );
  NAND2_X1 U3814 ( .A1(n4169), .A2(n4395), .ZN(n3832) );
  NAND2_X1 U3815 ( .A1(n3863), .A2(n3832), .ZN(n4190) );
  NAND2_X1 U3816 ( .A1(n4398), .A2(n4173), .ZN(n3037) );
  AOI22_X1 U3817 ( .A1(n4165), .A2(n3037), .B1(n3094), .B2(n4151), .ZN(n4154)
         );
  NAND2_X1 U3818 ( .A1(n4133), .A2(n4145), .ZN(n4127) );
  NAND2_X1 U3819 ( .A1(n4126), .A2(n4127), .ZN(n4153) );
  NAND2_X1 U3820 ( .A1(n4154), .A2(n4153), .ZN(n4152) );
  NAND2_X1 U3821 ( .A1(n4146), .A2(n4138), .ZN(n3041) );
  INV_X1 U3822 ( .A(n4114), .ZN(n3042) );
  NAND2_X1 U3823 ( .A1(n4091), .A2(n3042), .ZN(n3757) );
  OR2_X1 U3824 ( .A1(n4091), .A2(n3042), .ZN(n3758) );
  NAND2_X1 U3825 ( .A1(n3043), .A2(n3758), .ZN(n4086) );
  INV_X1 U3826 ( .A(n4081), .ZN(n3046) );
  OR2_X1 U3827 ( .A1(n4089), .A2(n3046), .ZN(n3077) );
  NAND2_X1 U3828 ( .A1(n4089), .A2(n3046), .ZN(n4050) );
  NAND2_X1 U3829 ( .A1(n4070), .A2(n3045), .ZN(n4069) );
  INV_X1 U3830 ( .A(n4089), .ZN(n4056) );
  NAND2_X1 U3831 ( .A1(n4056), .A2(n3046), .ZN(n3047) );
  NAND2_X1 U3832 ( .A1(n4069), .A2(n3047), .ZN(n4045) );
  NAND2_X1 U3833 ( .A1(n4072), .A2(n4054), .ZN(n3048) );
  NOR2_X1 U3834 ( .A1(n4059), .A2(n3679), .ZN(n3049) );
  INV_X1 U3835 ( .A(n4021), .ZN(n3078) );
  NOR2_X1 U3836 ( .A1(n3232), .A2(n3078), .ZN(n3592) );
  NAND2_X1 U3837 ( .A1(n3232), .A2(n3078), .ZN(n3593) );
  INV_X1 U3838 ( .A(n3721), .ZN(n3604) );
  XNOR2_X1 U3839 ( .A(n3996), .B(n3604), .ZN(n3755) );
  XNOR2_X1 U3840 ( .A(n3050), .B(n3755), .ZN(n4002) );
  XNOR2_X1 U3841 ( .A(n3051), .B(n3897), .ZN(n3052) );
  NAND2_X1 U3842 ( .A1(n3052), .A2(n3959), .ZN(n4226) );
  OR2_X1 U3843 ( .A1(n3750), .A2(n4569), .ZN(n3782) );
  OAI21_X1 U3844 ( .B1(n3053), .B2(n3782), .A(n3787), .ZN(n4223) );
  INV_X1 U3845 ( .A(n4224), .ZN(n3766) );
  NAND2_X1 U3846 ( .A1(n4223), .A2(n3766), .ZN(n3054) );
  NAND2_X1 U3847 ( .A1(n3054), .A2(n3788), .ZN(n3214) );
  OR2_X1 U3848 ( .A1(n4229), .A2(n3173), .ZN(n3793) );
  NAND2_X1 U3849 ( .A1(n4229), .A2(n3173), .ZN(n3790) );
  NAND2_X1 U3850 ( .A1(n3214), .A2(n3769), .ZN(n3055) );
  INV_X1 U3851 ( .A(n3794), .ZN(n3056) );
  AND2_X1 U3852 ( .A1(n3196), .A2(n3277), .ZN(n3318) );
  OR2_X1 U3853 ( .A1(n3196), .A2(n3277), .ZN(n3814) );
  NAND2_X1 U3854 ( .A1(n3057), .A2(n3814), .ZN(n3334) );
  NAND2_X1 U3855 ( .A1(n3908), .A2(n3289), .ZN(n3796) );
  NOR2_X1 U3856 ( .A1(n3908), .A2(n3289), .ZN(n3800) );
  AOI21_X1 U3857 ( .B1(n3334), .B2(n3796), .A(n3800), .ZN(n3297) );
  NAND2_X1 U3858 ( .A1(n3297), .A2(n3058), .ZN(n3059) );
  NAND2_X1 U3859 ( .A1(n3059), .A2(n3805), .ZN(n3362) );
  OR2_X1 U3860 ( .A1(n3907), .A2(n3367), .ZN(n3806) );
  NAND2_X1 U3861 ( .A1(n3907), .A2(n3367), .ZN(n3804) );
  AND2_X1 U3862 ( .A1(n3906), .A2(n3395), .ZN(n3823) );
  OR2_X1 U3863 ( .A1(n3906), .A2(n3395), .ZN(n3807) );
  NAND2_X1 U3864 ( .A1(n3905), .A2(n3420), .ZN(n3825) );
  NAND2_X1 U3865 ( .A1(n3419), .A2(n3825), .ZN(n3060) );
  NAND2_X1 U3866 ( .A1(n3543), .A2(n3488), .ZN(n3535) );
  NAND2_X1 U3867 ( .A1(n4203), .A2(n3558), .ZN(n3061) );
  NAND2_X1 U3868 ( .A1(n3535), .A2(n3061), .ZN(n3063) );
  INV_X1 U3869 ( .A(n3470), .ZN(n3062) );
  NOR2_X1 U3870 ( .A1(n3063), .A2(n3062), .ZN(n3826) );
  INV_X1 U3871 ( .A(n3063), .ZN(n3066) );
  OR2_X1 U3872 ( .A1(n3543), .A2(n3488), .ZN(n3537) );
  NAND2_X1 U3873 ( .A1(n3468), .A2(n3537), .ZN(n3065) );
  NOR2_X1 U3874 ( .A1(n4203), .A2(n3558), .ZN(n3064) );
  AOI21_X1 U3875 ( .B1(n3066), .B2(n3065), .A(n3064), .ZN(n3828) );
  OR2_X1 U3876 ( .A1(n4187), .A2(n3732), .ZN(n3829) );
  NAND2_X1 U3877 ( .A1(n4187), .A2(n3732), .ZN(n3812) );
  NAND2_X1 U3878 ( .A1(n3829), .A2(n3812), .ZN(n3743) );
  INV_X1 U3879 ( .A(n3830), .ZN(n3067) );
  NOR2_X1 U3880 ( .A1(n3743), .A2(n3067), .ZN(n3068) );
  NAND2_X1 U3881 ( .A1(n4204), .A2(n3068), .ZN(n3069) );
  INV_X1 U3882 ( .A(n4190), .ZN(n4182) );
  NAND2_X1 U3883 ( .A1(n4112), .A2(n4138), .ZN(n3070) );
  NAND2_X1 U3884 ( .A1(n4127), .A2(n3070), .ZN(n3071) );
  AND2_X1 U3885 ( .A1(n4151), .A2(n4173), .ZN(n4125) );
  INV_X1 U3886 ( .A(n3071), .ZN(n3074) );
  OR2_X1 U3887 ( .A1(n4151), .A2(n4173), .ZN(n4124) );
  NAND2_X1 U3888 ( .A1(n4126), .A2(n4124), .ZN(n3073) );
  NOR2_X1 U3889 ( .A1(n4112), .A2(n4138), .ZN(n3072) );
  AOI21_X1 U3890 ( .B1(n3074), .B2(n3073), .A(n3072), .ZN(n4105) );
  OR2_X1 U3891 ( .A1(n4091), .A2(n4114), .ZN(n3075) );
  AND2_X1 U3892 ( .A1(n4091), .A2(n4114), .ZN(n3866) );
  NAND2_X1 U3893 ( .A1(n4104), .A2(n2382), .ZN(n4046) );
  NAND2_X1 U3894 ( .A1(n4050), .A2(n4046), .ZN(n3870) );
  AND2_X1 U3895 ( .A1(n4073), .A2(n4094), .ZN(n3838) );
  NAND2_X1 U3896 ( .A1(n4072), .A2(n4061), .ZN(n3076) );
  NAND2_X1 U3897 ( .A1(n3077), .A2(n3076), .ZN(n3841) );
  AOI21_X1 U3898 ( .B1(n3838), .B2(n4050), .A(n3841), .ZN(n3869) );
  OAI21_X1 U3899 ( .B1(n4087), .B2(n3870), .A(n3869), .ZN(n4030) );
  NOR2_X1 U3900 ( .A1(n4016), .A2(n3679), .ZN(n3753) );
  NOR2_X1 U3901 ( .A1(n4072), .A2(n4061), .ZN(n4028) );
  NOR2_X1 U3902 ( .A1(n3753), .A2(n4028), .ZN(n3874) );
  AND2_X1 U3903 ( .A1(n4016), .A2(n3679), .ZN(n3780) );
  NAND2_X1 U3904 ( .A1(n3232), .A2(n4021), .ZN(n3781) );
  INV_X1 U3905 ( .A(n3232), .ZN(n4036) );
  NAND2_X1 U3906 ( .A1(n4036), .A2(n3078), .ZN(n3754) );
  NAND2_X1 U3907 ( .A1(n3606), .A2(n3754), .ZN(n3079) );
  XNOR2_X1 U3908 ( .A(n3079), .B(n3755), .ZN(n3081) );
  NAND2_X1 U3909 ( .A1(n3785), .A2(n2542), .ZN(n3888) );
  OR2_X1 U3910 ( .A1(n3897), .A2(n3959), .ZN(n3080) );
  NAND2_X1 U3911 ( .A1(n3081), .A2(n4571), .ZN(n3085) );
  AOI22_X1 U3912 ( .A1(n3232), .A2(n4227), .B1(n4055), .B2(n3604), .ZN(n3084)
         );
  OAI211_X1 U3913 ( .C1(n3779), .C2(n4574), .A(n3085), .B(n3084), .ZN(n4008)
         );
  AOI21_X1 U3914 ( .B1(n4002), .B2(n4642), .A(n4008), .ZN(n3100) );
  NAND2_X1 U3915 ( .A1(n3203), .A2(n3116), .ZN(n3091) );
  INV_X1 U3916 ( .A(n3201), .ZN(n3086) );
  NOR2_X1 U3917 ( .A1(n3087), .A2(n3086), .ZN(n3088) );
  AND2_X1 U3918 ( .A1(n3088), .A2(n3202), .ZN(n3090) );
  MUX2_X1 U3919 ( .A(n3092), .B(n3100), .S(n4658), .Z(n3097) );
  AND2_X1 U3920 ( .A1(n3253), .A2(n4569), .ZN(n3235) );
  NAND2_X1 U3921 ( .A1(n3235), .A2(n4232), .ZN(n4609) );
  NAND2_X1 U3922 ( .A1(n3368), .A2(n3367), .ZN(n3385) );
  OAI21_X1 U3923 ( .B1(n4019), .B2(n3721), .A(n2245), .ZN(n4003) );
  NAND2_X1 U3924 ( .A1(n3097), .A2(n3096), .ZN(U3544) );
  INV_X1 U3925 ( .A(REG0_REG_26__SCAN_IN), .ZN(n3101) );
  MUX2_X1 U3926 ( .A(n3101), .B(n3100), .S(n4645), .Z(n3103) );
  NAND2_X1 U3927 ( .A1(n3103), .A2(n3102), .ZN(U3512) );
  INV_X2 U3928 ( .A(n3910), .ZN(U4043) );
  INV_X2 U3929 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  INV_X1 U3930 ( .A(DATAI_14_), .ZN(n4914) );
  NAND2_X1 U3931 ( .A1(n4512), .A2(STATE_REG_SCAN_IN), .ZN(n3104) );
  OAI21_X1 U3932 ( .B1(STATE_REG_SCAN_IN), .B2(n4914), .A(n3104), .ZN(U3338)
         );
  NAND2_X1 U3933 ( .A1(U3149), .A2(DATAI_25_), .ZN(n3105) );
  OAI21_X1 U3934 ( .B1(n3106), .B2(U3149), .A(n3105), .ZN(U3327) );
  NAND3_X1 U3935 ( .A1(n3108), .A2(STATE_REG_SCAN_IN), .A3(IR_REG_31__SCAN_IN), 
        .ZN(n3109) );
  INV_X1 U3936 ( .A(DATAI_31_), .ZN(n4769) );
  OAI22_X1 U3937 ( .A1(n3107), .A2(n3109), .B1(STATE_REG_SCAN_IN), .B2(n4769), 
        .ZN(U3321) );
  INV_X1 U3938 ( .A(DATAI_21_), .ZN(n4973) );
  NAND2_X1 U3939 ( .A1(n3785), .A2(STATE_REG_SCAN_IN), .ZN(n3110) );
  OAI21_X1 U3940 ( .B1(STATE_REG_SCAN_IN), .B2(n4973), .A(n3110), .ZN(U3331)
         );
  INV_X1 U3941 ( .A(DATAI_30_), .ZN(n4980) );
  NAND2_X1 U3942 ( .A1(n3111), .A2(STATE_REG_SCAN_IN), .ZN(n3112) );
  OAI21_X1 U3943 ( .B1(STATE_REG_SCAN_IN), .B2(n4980), .A(n3112), .ZN(U3322)
         );
  INV_X1 U3944 ( .A(D_REG_0__SCAN_IN), .ZN(n4961) );
  INV_X1 U3945 ( .A(n3114), .ZN(n3115) );
  AOI22_X1 U3946 ( .A1(n4583), .A2(n4961), .B1(n3115), .B2(n3117), .ZN(U3458)
         );
  INV_X1 U3947 ( .A(D_REG_1__SCAN_IN), .ZN(n3119) );
  INV_X1 U3948 ( .A(n3116), .ZN(n3118) );
  AOI22_X1 U3949 ( .A1(n4583), .A2(n3119), .B1(n3118), .B2(n3117), .ZN(U3459)
         );
  OR2_X1 U3950 ( .A1(n3120), .A2(U3149), .ZN(n3902) );
  INV_X1 U3951 ( .A(n3902), .ZN(n3898) );
  OR2_X1 U3952 ( .A1(n3202), .A2(n3898), .ZN(n3128) );
  AOI21_X1 U3953 ( .B1(n3121), .B2(n3120), .A(n2572), .ZN(n3127) );
  INV_X1 U3954 ( .A(n3127), .ZN(n3122) );
  NOR2_X1 U3955 ( .A1(n5045), .A2(U4043), .ZN(U3148) );
  INV_X1 U3956 ( .A(DATAO_REG_7__SCAN_IN), .ZN(n4841) );
  NAND2_X1 U3957 ( .A1(n3366), .A2(U4043), .ZN(n3123) );
  OAI21_X1 U3958 ( .B1(U4043), .B2(n4841), .A(n3123), .ZN(U3557) );
  INV_X1 U3959 ( .A(DATAO_REG_5__SCAN_IN), .ZN(n4979) );
  NAND2_X1 U3960 ( .A1(n3196), .A2(U4043), .ZN(n3124) );
  OAI21_X1 U3961 ( .B1(U4043), .B2(n4979), .A(n3124), .ZN(U3555) );
  INV_X1 U3962 ( .A(DATAO_REG_11__SCAN_IN), .ZN(n4982) );
  NAND2_X1 U3963 ( .A1(n3473), .A2(U4043), .ZN(n3125) );
  OAI21_X1 U3964 ( .B1(U4043), .B2(n4982), .A(n3125), .ZN(U3561) );
  INV_X1 U3965 ( .A(DATAO_REG_2__SCAN_IN), .ZN(n4839) );
  NAND2_X1 U3966 ( .A1(n2576), .A2(U4043), .ZN(n3126) );
  OAI21_X1 U3967 ( .B1(U4043), .B2(n4839), .A(n3126), .ZN(U3552) );
  NAND2_X1 U3968 ( .A1(n3128), .A2(n3127), .ZN(n4422) );
  AND2_X1 U3969 ( .A1(U3149), .A2(REG3_REG_5__SCAN_IN), .ZN(n3278) );
  INV_X1 U3970 ( .A(n5045), .ZN(n4560) );
  INV_X1 U3971 ( .A(ADDR_REG_5__SCAN_IN), .ZN(n4837) );
  MUX2_X1 U3972 ( .A(REG2_REG_5__SCAN_IN), .B(n3129), .S(n4382), .Z(n3139) );
  MUX2_X1 U3973 ( .A(REG2_REG_2__SCAN_IN), .B(n3130), .S(n3144), .Z(n3913) );
  AND2_X1 U3974 ( .A1(REG2_REG_0__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n5044)
         );
  NAND2_X1 U3975 ( .A1(n3143), .A2(REG2_REG_1__SCAN_IN), .ZN(n3131) );
  NAND2_X1 U3976 ( .A1(REG2_REG_3__SCAN_IN), .A2(n4390), .ZN(n4389) );
  OAI21_X1 U3977 ( .B1(n3132), .B2(n2419), .A(n4389), .ZN(n3133) );
  XNOR2_X1 U3978 ( .A(n3133), .B(n4432), .ZN(n4427) );
  INV_X1 U3979 ( .A(n4432), .ZN(n3134) );
  NOR2_X1 U3980 ( .A1(n3137), .A2(n3136), .ZN(n4419) );
  NAND2_X1 U3981 ( .A1(n4377), .A2(n4419), .ZN(n3922) );
  NAND2_X1 U3982 ( .A1(n3508), .A2(n3139), .ZN(n3138) );
  OAI211_X1 U3983 ( .C1(n3139), .C2(n3508), .A(n5042), .B(n3138), .ZN(n3140)
         );
  OAI21_X1 U3984 ( .B1(n4560), .B2(n4837), .A(n3140), .ZN(n3141) );
  NOR2_X1 U3985 ( .A1(n3278), .A2(n3141), .ZN(n3151) );
  MUX2_X1 U3986 ( .A(REG1_REG_5__SCAN_IN), .B(n3142), .S(n4382), .Z(n3149) );
  INV_X1 U3987 ( .A(REG1_REG_1__SCAN_IN), .ZN(n4647) );
  AOI21_X1 U3988 ( .B1(n3143), .B2(REG1_REG_1__SCAN_IN), .A(n5036), .ZN(n3917)
         );
  MUX2_X1 U3989 ( .A(n4879), .B(REG1_REG_2__SCAN_IN), .S(n3144), .Z(n3916) );
  XNOR2_X1 U3990 ( .A(n3146), .B(n4383), .ZN(n4388) );
  NAND2_X1 U3991 ( .A1(REG1_REG_3__SCAN_IN), .A2(n4388), .ZN(n4387) );
  NAND2_X1 U3992 ( .A1(n4387), .A2(n2467), .ZN(n3147) );
  MUX2_X1 U3993 ( .A(n3142), .B(REG1_REG_5__SCAN_IN), .S(n4382), .Z(n3148) );
  OAI211_X1 U3994 ( .C1(n3149), .C2(n2280), .A(n5038), .B(n3495), .ZN(n3150)
         );
  OAI211_X1 U3995 ( .C1(n4547), .C2(n3509), .A(n3151), .B(n3150), .ZN(U3245)
         );
  NAND2_X1 U3996 ( .A1(n3152), .A2(n3202), .ZN(n3153) );
  NOR2_X1 U3997 ( .A1(n3154), .A2(n3153), .ZN(n3261) );
  INV_X1 U3998 ( .A(n4405), .ZN(n3704) );
  XNOR2_X1 U3999 ( .A(n3156), .B(n3155), .ZN(n3921) );
  INV_X1 U4000 ( .A(n3018), .ZN(n4575) );
  OAI22_X1 U4001 ( .A1(n3704), .A2(n3921), .B1(n4575), .B2(n3720), .ZN(n3157)
         );
  AOI21_X1 U4002 ( .B1(n3236), .B2(n3165), .A(n3157), .ZN(n3158) );
  OAI21_X1 U4003 ( .B1(n3261), .B2(n3159), .A(n3158), .ZN(U3229) );
  OAI21_X1 U4004 ( .B1(n3160), .B2(n3162), .A(n3161), .ZN(n3163) );
  NAND2_X1 U4005 ( .A1(n3163), .A2(n4405), .ZN(n3167) );
  OAI22_X1 U4006 ( .A1(n3266), .A2(n3720), .B1(n3722), .B2(n4575), .ZN(n3164)
         );
  AOI21_X1 U4007 ( .B1(n4239), .B2(n3165), .A(n3164), .ZN(n3166) );
  OAI211_X1 U4008 ( .C1(n3261), .C2(n3168), .A(n3167), .B(n3166), .ZN(U3234)
         );
  OAI21_X1 U4009 ( .B1(n3171), .B2(n3170), .A(n3169), .ZN(n3172) );
  NAND2_X1 U4010 ( .A1(n3172), .A2(n4405), .ZN(n3179) );
  INV_X1 U4011 ( .A(n2576), .ZN(n3254) );
  OAI22_X1 U4012 ( .A1(n3733), .A2(n3173), .B1(n3254), .B2(n3722), .ZN(n3177)
         );
  INV_X1 U4013 ( .A(n3909), .ZN(n3321) );
  INV_X1 U4014 ( .A(REG3_REG_3__SCAN_IN), .ZN(n3174) );
  NOR2_X1 U4015 ( .A1(STATE_REG_SCAN_IN), .A2(n3174), .ZN(n4384) );
  INV_X1 U4016 ( .A(n4384), .ZN(n3175) );
  OAI21_X1 U4017 ( .B1(n3720), .B2(n3321), .A(n3175), .ZN(n3176) );
  NOR2_X1 U4018 ( .A1(n3177), .A2(n3176), .ZN(n3178) );
  OAI211_X1 U4019 ( .C1(REG3_REG_3__SCAN_IN), .C2(n4410), .A(n3179), .B(n3178), 
        .ZN(U3215) );
  INV_X1 U4020 ( .A(DATAO_REG_19__SCAN_IN), .ZN(n4983) );
  NAND2_X1 U4021 ( .A1(n4112), .A2(U4043), .ZN(n3180) );
  OAI21_X1 U4022 ( .B1(U4043), .B2(n4983), .A(n3180), .ZN(U3569) );
  INV_X1 U4023 ( .A(DATAO_REG_12__SCAN_IN), .ZN(n4843) );
  NAND2_X1 U4024 ( .A1(n3543), .A2(U4043), .ZN(n3181) );
  OAI21_X1 U4025 ( .B1(U4043), .B2(n4843), .A(n3181), .ZN(U3562) );
  INV_X1 U4026 ( .A(DATAO_REG_29__SCAN_IN), .ZN(n3184) );
  INV_X1 U4027 ( .A(n3969), .ZN(n3182) );
  NAND2_X1 U4028 ( .A1(n3182), .A2(U4043), .ZN(n3183) );
  OAI21_X1 U4029 ( .B1(U4043), .B2(n3184), .A(n3183), .ZN(U3579) );
  INV_X1 U4030 ( .A(DATAO_REG_31__SCAN_IN), .ZN(n4960) );
  INV_X1 U4031 ( .A(REG2_REG_31__SCAN_IN), .ZN(n3188) );
  NAND2_X1 U4032 ( .A1(n2563), .A2(REG1_REG_31__SCAN_IN), .ZN(n3187) );
  INV_X1 U4033 ( .A(REG0_REG_31__SCAN_IN), .ZN(n3185) );
  OR2_X1 U4034 ( .A1(n2566), .A2(n3185), .ZN(n3186) );
  OAI211_X1 U4035 ( .C1(n3230), .C2(n3188), .A(n3187), .B(n3186), .ZN(n4245)
         );
  NAND2_X1 U4036 ( .A1(n4245), .A2(U4043), .ZN(n3189) );
  OAI21_X1 U4037 ( .B1(U4043), .B2(n4960), .A(n3189), .ZN(U3581) );
  INV_X1 U4038 ( .A(DATAO_REG_13__SCAN_IN), .ZN(n4966) );
  NAND2_X1 U4039 ( .A1(n4203), .A2(U4043), .ZN(n3191) );
  OAI21_X1 U4040 ( .B1(U4043), .B2(n4966), .A(n3191), .ZN(U3563) );
  XNOR2_X1 U4041 ( .A(n3192), .B(n3193), .ZN(n3209) );
  INV_X1 U4042 ( .A(n3193), .ZN(n3771) );
  XNOR2_X1 U40430 ( .A(n3194), .B(n3771), .ZN(n3199) );
  INV_X1 U4044 ( .A(n4188), .ZN(n3445) );
  INV_X1 U4045 ( .A(n4574), .ZN(n4228) );
  AOI22_X1 U4046 ( .A1(n3196), .A2(n4228), .B1(n4055), .B2(n3195), .ZN(n3197)
         );
  OAI21_X1 U4047 ( .B1(n3266), .B2(n3445), .A(n3197), .ZN(n3198) );
  AOI21_X1 U4048 ( .B1(n3199), .B2(n4571), .A(n3198), .ZN(n3200) );
  OAI21_X1 U4049 ( .B1(n3209), .B2(n4226), .A(n3200), .ZN(n4621) );
  OAI211_X1 U4050 ( .C1(n3219), .C2(n3267), .A(n3326), .B(n4619), .ZN(n4620)
         );
  OAI22_X1 U4051 ( .A1(n4620), .A2(n4380), .B1(n4213), .B2(n3273), .ZN(n3208)
         );
  AND3_X1 U4052 ( .A1(n3203), .A2(n3202), .A3(n3201), .ZN(n3204) );
  NAND3_X1 U4053 ( .A1(n3206), .A2(n3205), .A3(n3204), .ZN(n3207) );
  OAI21_X1 U4054 ( .B1(n4621), .B2(n3208), .A(n3576), .ZN(n3212) );
  INV_X1 U4055 ( .A(n3209), .ZN(n4624) );
  NAND2_X1 U4056 ( .A1(n3051), .A2(n4380), .ZN(n3238) );
  INV_X1 U4057 ( .A(n3238), .ZN(n3210) );
  NAND2_X1 U4058 ( .A1(n3576), .A2(n3210), .ZN(n4221) );
  INV_X1 U4059 ( .A(n4221), .ZN(n4578) );
  AOI22_X1 U4060 ( .A1(n4624), .A2(n4578), .B1(REG2_REG_4__SCAN_IN), .B2(n4581), .ZN(n3211) );
  NAND2_X1 U4061 ( .A1(n3212), .A2(n3211), .ZN(U3286) );
  XNOR2_X1 U4062 ( .A(n3213), .B(n3769), .ZN(n4615) );
  XNOR2_X1 U4063 ( .A(n3214), .B(n3769), .ZN(n3217) );
  AOI22_X1 U4064 ( .A1(n3909), .A2(n4228), .B1(n4055), .B2(n3220), .ZN(n3215)
         );
  OAI21_X1 U4065 ( .B1(n3254), .B2(n3445), .A(n3215), .ZN(n3216) );
  AOI21_X1 U4066 ( .B1(n3217), .B2(n4571), .A(n3216), .ZN(n3218) );
  OAI21_X1 U4067 ( .B1(n4615), .B2(n4226), .A(n3218), .ZN(n4616) );
  NAND2_X1 U4068 ( .A1(n4616), .A2(n3576), .ZN(n3224) );
  AOI21_X1 U4069 ( .B1(n3220), .B2(n4609), .A(n3219), .ZN(n4618) );
  OAI22_X1 U4071 ( .A1(n3576), .A2(n3221), .B1(n4213), .B2(REG3_REG_3__SCAN_IN), .ZN(n3222) );
  AOI21_X1 U4072 ( .B1(n4563), .B2(n4618), .A(n3222), .ZN(n3223) );
  OAI211_X1 U4073 ( .C1(n4615), .C2(n4221), .A(n3224), .B(n3223), .ZN(U3287)
         );
  INV_X1 U4074 ( .A(DATAO_REG_23__SCAN_IN), .ZN(n4958) );
  NAND2_X1 U4075 ( .A1(n4072), .A2(U4043), .ZN(n3225) );
  OAI21_X1 U4076 ( .B1(U4043), .B2(n4958), .A(n3225), .ZN(U3573) );
  INV_X1 U4077 ( .A(DATAO_REG_30__SCAN_IN), .ZN(n4850) );
  INV_X1 U4078 ( .A(REG2_REG_30__SCAN_IN), .ZN(n3229) );
  NAND2_X1 U4079 ( .A1(n2563), .A2(REG1_REG_30__SCAN_IN), .ZN(n3228) );
  INV_X1 U4080 ( .A(REG0_REG_30__SCAN_IN), .ZN(n3226) );
  OR2_X1 U4081 ( .A1(n2566), .A2(n3226), .ZN(n3227) );
  OAI211_X1 U4082 ( .C1(n3230), .C2(n3229), .A(n3228), .B(n3227), .ZN(n3751)
         );
  NAND2_X1 U4083 ( .A1(n3751), .A2(U4043), .ZN(n3231) );
  OAI21_X1 U4084 ( .B1(U4043), .B2(n4850), .A(n3231), .ZN(U3580) );
  INV_X1 U4085 ( .A(DATAO_REG_25__SCAN_IN), .ZN(n4974) );
  NAND2_X1 U4086 ( .A1(n3232), .A2(U4043), .ZN(n3233) );
  OAI21_X1 U4087 ( .B1(U4043), .B2(n4974), .A(n3233), .ZN(U3575) );
  INV_X1 U4088 ( .A(DATAO_REG_0__SCAN_IN), .ZN(n4951) );
  NAND2_X1 U4089 ( .A1(n3750), .A2(U4043), .ZN(n3234) );
  OAI21_X1 U4090 ( .B1(U4043), .B2(n4951), .A(n3234), .ZN(U3550) );
  INV_X1 U4091 ( .A(n3235), .ZN(n4240) );
  NAND2_X1 U4092 ( .A1(n3236), .A2(n3243), .ZN(n3237) );
  NAND2_X1 U4093 ( .A1(n4240), .A2(n3237), .ZN(n4604) );
  NAND2_X1 U4094 ( .A1(n4226), .A2(n3238), .ZN(n3239) );
  OAI21_X1 U4095 ( .B1(n3053), .B2(n3241), .A(n3240), .ZN(n4606) );
  INV_X1 U4096 ( .A(n4606), .ZN(n3242) );
  AOI22_X1 U4097 ( .A1(n4196), .A2(n3242), .B1(REG3_REG_1__SCAN_IN), .B2(n4577), .ZN(n3249) );
  XNOR2_X1 U4098 ( .A(n3053), .B(n3782), .ZN(n3246) );
  INV_X1 U4099 ( .A(n3750), .ZN(n3255) );
  AOI22_X1 U4100 ( .A1(n2576), .A2(n4228), .B1(n4055), .B2(n3243), .ZN(n3244)
         );
  OAI21_X1 U4101 ( .B1(n3255), .B2(n3445), .A(n3244), .ZN(n3245) );
  AOI21_X1 U4102 ( .B1(n3246), .B2(n4571), .A(n3245), .ZN(n4603) );
  MUX2_X1 U4103 ( .A(n4603), .B(n3247), .S(n4581), .Z(n3248) );
  OAI211_X1 U4104 ( .C1(n4175), .C2(n4604), .A(n3249), .B(n3248), .ZN(U3289)
         );
  XOR2_X1 U4105 ( .A(n3250), .B(n3251), .Z(n3252) );
  NAND2_X1 U4106 ( .A1(n3252), .A2(n4405), .ZN(n3259) );
  NOR2_X1 U4107 ( .A1(n3733), .A2(n3253), .ZN(n3257) );
  OAI22_X1 U4108 ( .A1(n3255), .A2(n3722), .B1(n3720), .B2(n3254), .ZN(n3256)
         );
  NOR2_X1 U4109 ( .A1(n3257), .A2(n3256), .ZN(n3258) );
  OAI211_X1 U4110 ( .C1(n3261), .C2(n3260), .A(n3259), .B(n3258), .ZN(U3219)
         );
  AND2_X1 U4111 ( .A1(n3169), .A2(n3262), .ZN(n3265) );
  OAI211_X1 U4112 ( .C1(n3265), .C2(n3264), .A(n3263), .B(n4405), .ZN(n3272)
         );
  OAI22_X1 U4113 ( .A1(n3733), .A2(n3267), .B1(n3266), .B2(n3722), .ZN(n3270)
         );
  AND2_X1 U4114 ( .A1(U3149), .A2(REG3_REG_4__SCAN_IN), .ZN(n4424) );
  INV_X1 U4115 ( .A(n4424), .ZN(n3268) );
  OAI21_X1 U4116 ( .B1(n3720), .B2(n3336), .A(n3268), .ZN(n3269) );
  NOR2_X1 U4117 ( .A1(n3270), .A2(n3269), .ZN(n3271) );
  OAI211_X1 U4118 ( .C1(n4410), .C2(n3273), .A(n3272), .B(n3271), .ZN(U3227)
         );
  XOR2_X1 U4119 ( .A(n3275), .B(n3274), .Z(n3276) );
  NAND2_X1 U4120 ( .A1(n3276), .A2(n4405), .ZN(n3283) );
  OAI22_X1 U4121 ( .A1(n3733), .A2(n3277), .B1(n3321), .B2(n3722), .ZN(n3281)
         );
  INV_X1 U4122 ( .A(n3278), .ZN(n3279) );
  OAI21_X1 U4123 ( .B1(n3720), .B2(n3312), .A(n3279), .ZN(n3280) );
  NOR2_X1 U4124 ( .A1(n3281), .A2(n3280), .ZN(n3282) );
  OAI211_X1 U4125 ( .C1(n4410), .C2(n3328), .A(n3283), .B(n3282), .ZN(U3224)
         );
  INV_X1 U4126 ( .A(n3284), .ZN(n3286) );
  NOR2_X1 U4127 ( .A1(n3286), .A2(n3285), .ZN(n3287) );
  XNOR2_X1 U4128 ( .A(n2276), .B(n3287), .ZN(n3288) );
  NAND2_X1 U4129 ( .A1(n3288), .A2(n4405), .ZN(n3294) );
  OAI22_X1 U4130 ( .A1(n3733), .A2(n3289), .B1(n3336), .B2(n3722), .ZN(n3292)
         );
  INV_X1 U4131 ( .A(n3366), .ZN(n3357) );
  NOR2_X1 U4132 ( .A1(STATE_REG_SCAN_IN), .A2(n4963), .ZN(n4435) );
  INV_X1 U4133 ( .A(n4435), .ZN(n3290) );
  OAI21_X1 U4134 ( .B1(n3720), .B2(n3357), .A(n3290), .ZN(n3291) );
  NOR2_X1 U4135 ( .A1(n3292), .A2(n3291), .ZN(n3293) );
  OAI211_X1 U4136 ( .C1(n4410), .C2(n3295), .A(n3294), .B(n3293), .ZN(U3236)
         );
  INV_X1 U4137 ( .A(n3296), .ZN(n3802) );
  XNOR2_X1 U4138 ( .A(n3297), .B(n3802), .ZN(n3300) );
  OAI22_X1 U4139 ( .A1(n3394), .A2(n4574), .B1(n4255), .B2(n3310), .ZN(n3298)
         );
  AOI21_X1 U4140 ( .B1(n4227), .B2(n3908), .A(n3298), .ZN(n3299) );
  OAI21_X1 U4141 ( .B1(n3300), .B2(n4236), .A(n3299), .ZN(n4631) );
  INV_X1 U4142 ( .A(n4631), .ZN(n3306) );
  XNOR2_X1 U4143 ( .A(n3301), .B(n3802), .ZN(n4633) );
  NAND2_X1 U4144 ( .A1(n4633), .A2(n4196), .ZN(n3305) );
  AOI211_X1 U4145 ( .C1(n3302), .C2(n3342), .A(n4638), .B(n3368), .ZN(n4632)
         );
  OAI22_X1 U4146 ( .A1(n3576), .A2(n2654), .B1(n3317), .B2(n4213), .ZN(n3303)
         );
  AOI21_X1 U4147 ( .B1(n4632), .B2(n4158), .A(n3303), .ZN(n3304) );
  OAI211_X1 U4148 ( .C1(n3306), .C2(n4581), .A(n3305), .B(n3304), .ZN(U3283)
         );
  OAI211_X1 U4149 ( .C1(n3309), .C2(n3308), .A(n3307), .B(n4405), .ZN(n3316)
         );
  OAI22_X1 U4150 ( .A1(n3733), .A2(n3310), .B1(n3394), .B2(n3720), .ZN(n3314)
         );
  NOR2_X1 U4151 ( .A1(n2651), .A2(STATE_REG_SCAN_IN), .ZN(n4449) );
  INV_X1 U4152 ( .A(n4449), .ZN(n3311) );
  OAI21_X1 U4153 ( .B1(n3722), .B2(n3312), .A(n3311), .ZN(n3313) );
  NOR2_X1 U4154 ( .A1(n3314), .A2(n3313), .ZN(n3315) );
  OAI211_X1 U4155 ( .C1(n4410), .C2(n3317), .A(n3316), .B(n3315), .ZN(U3210)
         );
  INV_X1 U4156 ( .A(n3318), .ZN(n3797) );
  AND2_X1 U4157 ( .A1(n3797), .A2(n3814), .ZN(n3768) );
  XOR2_X1 U4158 ( .A(n3768), .B(n3319), .Z(n3323) );
  AOI22_X1 U4159 ( .A1(n3908), .A2(n4228), .B1(n4055), .B2(n3325), .ZN(n3320)
         );
  OAI21_X1 U4160 ( .B1(n3321), .B2(n3445), .A(n3320), .ZN(n3322) );
  AOI21_X1 U4161 ( .B1(n3323), .B2(n4571), .A(n3322), .ZN(n4626) );
  XOR2_X1 U4162 ( .A(n3768), .B(n3324), .Z(n4629) );
  NAND2_X1 U4163 ( .A1(n3326), .A2(n3325), .ZN(n3327) );
  NAND2_X1 U4164 ( .A1(n3344), .A2(n3327), .ZN(n4627) );
  NOR2_X1 U4165 ( .A1(n4175), .A2(n4627), .ZN(n3330) );
  OAI22_X1 U4166 ( .A1(n3576), .A2(n3129), .B1(n3328), .B2(n4213), .ZN(n3329)
         );
  AOI211_X1 U4167 ( .C1(n4629), .C2(n4196), .A(n3330), .B(n3329), .ZN(n3331)
         );
  OAI21_X1 U4168 ( .B1(n4581), .B2(n4626), .A(n3331), .ZN(U3285) );
  INV_X1 U4169 ( .A(n4614), .ZN(n4623) );
  INV_X1 U4170 ( .A(n3796), .ZN(n3815) );
  OR2_X1 U4171 ( .A1(n3815), .A2(n3800), .ZN(n3333) );
  XNOR2_X1 U4172 ( .A(n3332), .B(n3333), .ZN(n3337) );
  INV_X1 U4173 ( .A(n3337), .ZN(n4564) );
  INV_X1 U4174 ( .A(n3333), .ZN(n3745) );
  XNOR2_X1 U4175 ( .A(n3334), .B(n3745), .ZN(n3340) );
  AOI22_X1 U4176 ( .A1(n3366), .A2(n4228), .B1(n4055), .B2(n3345), .ZN(n3335)
         );
  OAI21_X1 U4177 ( .B1(n3336), .B2(n3445), .A(n3335), .ZN(n3339) );
  NOR2_X1 U4178 ( .A1(n3337), .A2(n4226), .ZN(n3338) );
  AOI211_X1 U4179 ( .C1(n3340), .C2(n4571), .A(n3339), .B(n3338), .ZN(n4567)
         );
  INV_X1 U4180 ( .A(n4567), .ZN(n3341) );
  AOI21_X1 U4181 ( .B1(n4623), .B2(n4564), .A(n3341), .ZN(n3350) );
  INV_X1 U4182 ( .A(n3342), .ZN(n3343) );
  AOI21_X1 U4183 ( .B1(n3345), .B2(n3344), .A(n3343), .ZN(n4562) );
  AOI22_X1 U4184 ( .A1(n4562), .A2(n4264), .B1(n4656), .B2(REG1_REG_6__SCAN_IN), .ZN(n3346) );
  OAI21_X1 U4185 ( .B1(n3350), .B2(n4656), .A(n3346), .ZN(U3524) );
  INV_X1 U4186 ( .A(REG0_REG_6__SCAN_IN), .ZN(n3347) );
  NOR2_X1 U4187 ( .A1(n4645), .A2(n3347), .ZN(n3348) );
  AOI21_X1 U4188 ( .B1(n4562), .B2(n4329), .A(n3348), .ZN(n3349) );
  OAI21_X1 U4189 ( .B1(n3350), .B2(n4644), .A(n3349), .ZN(U3479) );
  XNOR2_X1 U4190 ( .A(n3352), .B(n3351), .ZN(n3353) );
  XNOR2_X1 U4191 ( .A(n3354), .B(n3353), .ZN(n3355) );
  NAND2_X1 U4192 ( .A1(n3355), .A2(n4405), .ZN(n3361) );
  OAI22_X1 U4193 ( .A1(n3733), .A2(n3367), .B1(n3414), .B2(n3720), .ZN(n3359)
         );
  INV_X1 U4194 ( .A(REG3_REG_8__SCAN_IN), .ZN(n4948) );
  NOR2_X1 U4195 ( .A1(STATE_REG_SCAN_IN), .A2(n4948), .ZN(n4458) );
  INV_X1 U4196 ( .A(n4458), .ZN(n3356) );
  OAI21_X1 U4197 ( .B1(n3722), .B2(n3357), .A(n3356), .ZN(n3358) );
  NOR2_X1 U4198 ( .A1(n3359), .A2(n3358), .ZN(n3360) );
  OAI211_X1 U4199 ( .C1(n4410), .C2(n3370), .A(n3361), .B(n3360), .ZN(U3218)
         );
  OAI22_X1 U4200 ( .A1(n3414), .A2(n4574), .B1(n4255), .B2(n3367), .ZN(n3365)
         );
  AND2_X1 U4201 ( .A1(n3806), .A2(n3804), .ZN(n3747) );
  XNOR2_X1 U4202 ( .A(n3362), .B(n3747), .ZN(n3363) );
  NOR2_X1 U4203 ( .A1(n3363), .A2(n4236), .ZN(n3364) );
  AOI211_X1 U4204 ( .C1(n4227), .C2(n3366), .A(n3365), .B(n3364), .ZN(n3400)
         );
  OR2_X1 U4205 ( .A1(n3368), .A2(n3367), .ZN(n3369) );
  NAND2_X1 U4206 ( .A1(n3385), .A2(n3369), .ZN(n3404) );
  INV_X1 U4207 ( .A(n3404), .ZN(n3376) );
  OAI22_X1 U4208 ( .A1(n3576), .A2(n3371), .B1(n3370), .B2(n4213), .ZN(n3375)
         );
  XNOR2_X1 U4209 ( .A(n3373), .B(n3747), .ZN(n3401) );
  NOR2_X1 U4210 ( .A1(n3401), .A2(n4180), .ZN(n3374) );
  AOI211_X1 U4211 ( .C1(n3376), .C2(n4563), .A(n3375), .B(n3374), .ZN(n3377)
         );
  OAI21_X1 U4212 ( .B1(n4581), .B2(n3400), .A(n3377), .ZN(U3282) );
  INV_X1 U4213 ( .A(n3823), .ZN(n3378) );
  AND2_X1 U4214 ( .A1(n3378), .A2(n3807), .ZN(n3749) );
  XOR2_X1 U4215 ( .A(n3749), .B(n3379), .Z(n3382) );
  AOI22_X1 U4216 ( .A1(n3905), .A2(n4228), .B1(n4055), .B2(n3384), .ZN(n3380)
         );
  OAI21_X1 U4217 ( .B1(n3394), .B2(n3445), .A(n3380), .ZN(n3381) );
  AOI21_X1 U4218 ( .B1(n3382), .B2(n4571), .A(n3381), .ZN(n4634) );
  XOR2_X1 U4219 ( .A(n3749), .B(n3383), .Z(n4637) );
  NAND2_X1 U4220 ( .A1(n3385), .A2(n3384), .ZN(n3386) );
  NAND2_X1 U4221 ( .A1(n3426), .A2(n3386), .ZN(n4635) );
  NOR2_X1 U4222 ( .A1(n4635), .A2(n4175), .ZN(n3388) );
  INV_X1 U4223 ( .A(REG2_REG_9__SCAN_IN), .ZN(n3506) );
  OAI22_X1 U4224 ( .A1(n3576), .A2(n3506), .B1(n3399), .B2(n4213), .ZN(n3387)
         );
  AOI211_X1 U4225 ( .C1(n4637), .C2(n4196), .A(n3388), .B(n3387), .ZN(n3389)
         );
  OAI21_X1 U4226 ( .B1(n4581), .B2(n4634), .A(n3389), .ZN(U3281) );
  OAI21_X1 U4227 ( .B1(n3392), .B2(n3390), .A(n3391), .ZN(n3393) );
  NAND2_X1 U4228 ( .A1(n3393), .A2(n4405), .ZN(n3398) );
  AND2_X1 U4229 ( .A1(U3149), .A2(REG3_REG_9__SCAN_IN), .ZN(n4467) );
  OAI22_X1 U4230 ( .A1(n3733), .A2(n3395), .B1(n3394), .B2(n3722), .ZN(n3396)
         );
  AOI211_X1 U4231 ( .C1(n3618), .C2(n3905), .A(n4467), .B(n3396), .ZN(n3397)
         );
  OAI211_X1 U4232 ( .C1(n4410), .C2(n3399), .A(n3398), .B(n3397), .ZN(U3228)
         );
  OAI21_X1 U4233 ( .B1(n4605), .B2(n3401), .A(n3400), .ZN(n3406) );
  INV_X1 U4234 ( .A(REG0_REG_8__SCAN_IN), .ZN(n4803) );
  OAI22_X1 U4235 ( .A1(n3404), .A2(n4374), .B1(n4645), .B2(n4803), .ZN(n3402)
         );
  AOI21_X1 U4236 ( .B1(n3406), .B2(n4645), .A(n3402), .ZN(n3403) );
  INV_X1 U4237 ( .A(n3403), .ZN(U3483) );
  OAI22_X1 U4238 ( .A1(n3404), .A2(n4323), .B1(n4658), .B2(n2669), .ZN(n3405)
         );
  AOI21_X1 U4239 ( .B1(n3406), .B2(n4658), .A(n3405), .ZN(n3407) );
  INV_X1 U4240 ( .A(n3407), .ZN(U3526) );
  AND2_X1 U4241 ( .A1(n3391), .A2(n3408), .ZN(n3411) );
  OAI211_X1 U4242 ( .C1(n3411), .C2(n3410), .A(n4405), .B(n3409), .ZN(n3418)
         );
  OAI22_X1 U4243 ( .A1(n3733), .A2(n3420), .B1(n3489), .B2(n3720), .ZN(n3416)
         );
  NOR2_X1 U4244 ( .A1(STATE_REG_SCAN_IN), .A2(n3412), .ZN(n4477) );
  INV_X1 U4245 ( .A(n4477), .ZN(n3413) );
  OAI21_X1 U4246 ( .B1(n3722), .B2(n3414), .A(n3413), .ZN(n3415) );
  NOR2_X1 U4247 ( .A1(n3416), .A2(n3415), .ZN(n3417) );
  OAI211_X1 U4248 ( .C1(n4410), .C2(n3429), .A(n3418), .B(n3417), .ZN(U3214)
         );
  AND2_X1 U4249 ( .A1(n3822), .A2(n3825), .ZN(n3770) );
  XOR2_X1 U4250 ( .A(n3770), .B(n3419), .Z(n3423) );
  OAI22_X1 U4251 ( .A1(n3489), .A2(n4574), .B1(n4255), .B2(n3420), .ZN(n3421)
         );
  AOI21_X1 U4252 ( .B1(n4188), .B2(n3906), .A(n3421), .ZN(n3422) );
  OAI21_X1 U4253 ( .B1(n3423), .B2(n4236), .A(n3422), .ZN(n3435) );
  INV_X1 U4254 ( .A(n3435), .ZN(n3434) );
  XOR2_X1 U4255 ( .A(n3770), .B(n3424), .Z(n3436) );
  INV_X1 U4256 ( .A(n3449), .ZN(n3428) );
  NAND2_X1 U4257 ( .A1(n3426), .A2(n3425), .ZN(n3427) );
  NAND2_X1 U4258 ( .A1(n3428), .A2(n3427), .ZN(n3440) );
  NOR2_X1 U4259 ( .A1(n3440), .A2(n4175), .ZN(n3432) );
  OAI22_X1 U4260 ( .A1(n3576), .A2(n3430), .B1(n3429), .B2(n4213), .ZN(n3431)
         );
  AOI211_X1 U4261 ( .C1(n3436), .C2(n4196), .A(n3432), .B(n3431), .ZN(n3433)
         );
  OAI21_X1 U4262 ( .B1(n4581), .B2(n3434), .A(n3433), .ZN(U3280) );
  AOI21_X1 U4263 ( .B1(n3436), .B2(n4642), .A(n3435), .ZN(n3438) );
  MUX2_X1 U4264 ( .A(n2700), .B(n3438), .S(n4645), .Z(n3437) );
  OAI21_X1 U4265 ( .B1(n3440), .B2(n4374), .A(n3437), .ZN(U3487) );
  INV_X1 U4266 ( .A(REG1_REG_10__SCAN_IN), .ZN(n4476) );
  MUX2_X1 U4267 ( .A(n4476), .B(n3438), .S(n4658), .Z(n3439) );
  OAI21_X1 U4268 ( .B1(n3440), .B2(n4323), .A(n3439), .ZN(U3528) );
  INV_X1 U4269 ( .A(n3446), .ZN(n3767) );
  XNOR2_X1 U4270 ( .A(n3471), .B(n3767), .ZN(n3441) );
  NAND2_X1 U4271 ( .A1(n3441), .A2(n4571), .ZN(n3444) );
  AOI22_X1 U4272 ( .A1(n3543), .A2(n4228), .B1(n4055), .B2(n3442), .ZN(n3443)
         );
  OAI211_X1 U4273 ( .C1(n3462), .C2(n3445), .A(n3444), .B(n3443), .ZN(n4640)
         );
  INV_X1 U4274 ( .A(n4640), .ZN(n3454) );
  XNOR2_X1 U4275 ( .A(n3447), .B(n3446), .ZN(n4643) );
  INV_X1 U4276 ( .A(n3477), .ZN(n3448) );
  OAI21_X1 U4277 ( .B1(n3449), .B2(n3459), .A(n3448), .ZN(n4639) );
  NOR2_X1 U4278 ( .A1(n4639), .A2(n4175), .ZN(n3452) );
  OAI22_X1 U4279 ( .A1(n3576), .A2(n3450), .B1(n3467), .B2(n4213), .ZN(n3451)
         );
  AOI211_X1 U4280 ( .C1(n4643), .C2(n4196), .A(n3452), .B(n3451), .ZN(n3453)
         );
  OAI21_X1 U4281 ( .B1(n4581), .B2(n3454), .A(n3453), .ZN(U3279) );
  NAND2_X1 U4282 ( .A1(n2278), .A2(n3455), .ZN(n3456) );
  XNOR2_X1 U4283 ( .A(n3457), .B(n3456), .ZN(n3458) );
  NAND2_X1 U4284 ( .A1(n3458), .A2(n4405), .ZN(n3466) );
  OAI22_X1 U4285 ( .A1(n3733), .A2(n3459), .B1(n3561), .B2(n3720), .ZN(n3464)
         );
  NOR2_X1 U4286 ( .A1(STATE_REG_SCAN_IN), .A2(n3460), .ZN(n4486) );
  INV_X1 U4287 ( .A(n4486), .ZN(n3461) );
  OAI21_X1 U4288 ( .B1(n3722), .B2(n3462), .A(n3461), .ZN(n3463) );
  NOR2_X1 U4289 ( .A1(n3464), .A2(n3463), .ZN(n3465) );
  OAI211_X1 U4290 ( .C1(n4410), .C2(n3467), .A(n3466), .B(n3465), .ZN(U3233)
         );
  INV_X1 U4291 ( .A(n3468), .ZN(n3469) );
  AOI21_X1 U4292 ( .B1(n3471), .B2(n3470), .A(n3469), .ZN(n3538) );
  AND2_X1 U4293 ( .A1(n3537), .A2(n3535), .ZN(n3748) );
  XNOR2_X1 U4294 ( .A(n3538), .B(n3748), .ZN(n3475) );
  INV_X1 U4295 ( .A(n4203), .ZN(n3586) );
  OAI22_X1 U4296 ( .A1(n3586), .A2(n4574), .B1(n4255), .B2(n3488), .ZN(n3472)
         );
  AOI21_X1 U4297 ( .B1(n4227), .B2(n3473), .A(n3472), .ZN(n3474) );
  OAI21_X1 U4298 ( .B1(n3475), .B2(n4236), .A(n3474), .ZN(n3526) );
  INV_X1 U4299 ( .A(n3526), .ZN(n3483) );
  XNOR2_X1 U4300 ( .A(n3476), .B(n3748), .ZN(n3527) );
  OR2_X1 U4301 ( .A1(n3477), .A2(n3488), .ZN(n3478) );
  NAND2_X1 U4302 ( .A1(n3545), .A2(n3478), .ZN(n3532) );
  NOR2_X1 U4303 ( .A1(n3532), .A2(n4175), .ZN(n3481) );
  OAI22_X1 U4304 ( .A1(n3576), .A2(n3479), .B1(n3494), .B2(n4213), .ZN(n3480)
         );
  AOI211_X1 U4305 ( .C1(n3527), .C2(n4196), .A(n3481), .B(n3480), .ZN(n3482)
         );
  OAI21_X1 U4306 ( .B1(n4581), .B2(n3483), .A(n3482), .ZN(U3278) );
  XNOR2_X1 U4307 ( .A(n2263), .B(n3484), .ZN(n3485) );
  XNOR2_X1 U4308 ( .A(n3486), .B(n3485), .ZN(n3487) );
  NAND2_X1 U4309 ( .A1(n3487), .A2(n4405), .ZN(n3493) );
  OAI22_X1 U4310 ( .A1(n3733), .A2(n3488), .B1(n3586), .B2(n3720), .ZN(n3491)
         );
  NAND2_X1 U4311 ( .A1(REG3_REG_12__SCAN_IN), .A2(U3149), .ZN(n3520) );
  OAI21_X1 U4312 ( .B1(n3722), .B2(n3489), .A(n3520), .ZN(n3490) );
  NOR2_X1 U4313 ( .A1(n3491), .A2(n3490), .ZN(n3492) );
  OAI211_X1 U4314 ( .C1(n4410), .C2(n3494), .A(n3493), .B(n3492), .ZN(U3221)
         );
  INV_X1 U4315 ( .A(n4440), .ZN(n4598) );
  XNOR2_X1 U4316 ( .A(n4598), .B(n3496), .ZN(n4437) );
  NAND2_X1 U4317 ( .A1(REG1_REG_6__SCAN_IN), .A2(n4437), .ZN(n4436) );
  NAND2_X1 U4318 ( .A1(n4440), .A2(n3496), .ZN(n3497) );
  NOR2_X1 U4319 ( .A1(n3499), .A2(n3500), .ZN(n3501) );
  XNOR2_X1 U4320 ( .A(n3500), .B(n3499), .ZN(n4457) );
  NOR2_X1 U4321 ( .A1(n2669), .A2(n4457), .ZN(n4456) );
  NOR2_X1 U4322 ( .A1(n3501), .A2(n4456), .ZN(n4466) );
  NAND2_X1 U4323 ( .A1(n3507), .A2(REG1_REG_9__SCAN_IN), .ZN(n3502) );
  OAI21_X1 U4324 ( .B1(n3507), .B2(REG1_REG_9__SCAN_IN), .A(n3502), .ZN(n4465)
         );
  NOR2_X1 U4325 ( .A1(n4466), .A2(n4465), .ZN(n4464) );
  INV_X1 U4326 ( .A(n4591), .ZN(n4493) );
  INV_X1 U4327 ( .A(REG1_REG_11__SCAN_IN), .ZN(n4880) );
  AOI22_X1 U4328 ( .A1(REG1_REG_11__SCAN_IN), .A2(n4493), .B1(n4591), .B2(
        n4880), .ZN(n4484) );
  NOR2_X1 U4329 ( .A1(n4485), .A2(n4484), .ZN(n4483) );
  AND2_X1 U4330 ( .A1(n4591), .A2(REG1_REG_11__SCAN_IN), .ZN(n3504) );
  AOI211_X1 U4331 ( .C1(n2487), .C2(n3505), .A(n3930), .B(n4548), .ZN(n3525)
         );
  NAND2_X1 U4332 ( .A1(n3507), .A2(REG2_REG_9__SCAN_IN), .ZN(n3516) );
  INV_X1 U4333 ( .A(n3507), .ZN(n4596) );
  AOI22_X1 U4334 ( .A1(n3507), .A2(REG2_REG_9__SCAN_IN), .B1(n3506), .B2(n4596), .ZN(n4471) );
  NAND2_X1 U4335 ( .A1(n4440), .A2(n3510), .ZN(n3511) );
  INV_X1 U4336 ( .A(n4445), .ZN(n4597) );
  AOI22_X1 U4337 ( .A1(REG2_REG_7__SCAN_IN), .A2(n4445), .B1(n4597), .B2(n2654), .ZN(n4453) );
  NAND2_X1 U4338 ( .A1(REG2_REG_7__SCAN_IN), .A2(n4445), .ZN(n3512) );
  NAND2_X1 U4339 ( .A1(n3513), .A2(n3514), .ZN(n3515) );
  NAND2_X1 U4340 ( .A1(REG2_REG_8__SCAN_IN), .A2(n4461), .ZN(n4460) );
  NAND2_X1 U4341 ( .A1(n4593), .A2(n3517), .ZN(n3518) );
  NAND2_X1 U4342 ( .A1(REG2_REG_10__SCAN_IN), .A2(n4480), .ZN(n4479) );
  NAND2_X1 U4343 ( .A1(n3518), .A2(n4479), .ZN(n4489) );
  AOI22_X1 U4344 ( .A1(REG2_REG_11__SCAN_IN), .A2(n4591), .B1(n4493), .B2(
        n3450), .ZN(n4490) );
  OAI211_X1 U4345 ( .C1(n3519), .C2(REG2_REG_12__SCAN_IN), .A(n5042), .B(n3945), .ZN(n3523) );
  INV_X1 U4346 ( .A(n3520), .ZN(n3521) );
  AOI21_X1 U4347 ( .B1(n5045), .B2(ADDR_REG_12__SCAN_IN), .A(n3521), .ZN(n3522) );
  OAI211_X1 U4348 ( .C1(n4547), .C2(n2417), .A(n3523), .B(n3522), .ZN(n3524)
         );
  OR2_X1 U4349 ( .A1(n3525), .A2(n3524), .ZN(U3252) );
  INV_X1 U4350 ( .A(REG0_REG_12__SCAN_IN), .ZN(n3528) );
  AOI21_X1 U4351 ( .B1(n3527), .B2(n4642), .A(n3526), .ZN(n3530) );
  MUX2_X1 U4352 ( .A(n3528), .B(n3530), .S(n4645), .Z(n3529) );
  OAI21_X1 U4353 ( .B1(n3532), .B2(n4374), .A(n3529), .ZN(U3491) );
  MUX2_X1 U4354 ( .A(n2487), .B(n3530), .S(n4658), .Z(n3531) );
  OAI21_X1 U4355 ( .B1(n3532), .B2(n4323), .A(n3531), .ZN(U3530) );
  OR2_X1 U4356 ( .A1(n3533), .A2(n3567), .ZN(n3746) );
  XNOR2_X1 U4357 ( .A(n3534), .B(n3746), .ZN(n4318) );
  OAI22_X1 U4358 ( .A1(n3731), .A2(n4574), .B1(n4255), .B2(n3558), .ZN(n3542)
         );
  INV_X1 U4359 ( .A(n3535), .ZN(n3536) );
  AOI21_X1 U4360 ( .B1(n3538), .B2(n3537), .A(n3536), .ZN(n3539) );
  XOR2_X1 U4361 ( .A(n3746), .B(n3539), .Z(n3540) );
  NOR2_X1 U4362 ( .A1(n3540), .A2(n4236), .ZN(n3541) );
  AOI211_X1 U4363 ( .C1(n4188), .C2(n3543), .A(n3542), .B(n3541), .ZN(n3544)
         );
  OAI21_X1 U4364 ( .B1(n4318), .B2(n4226), .A(n3544), .ZN(n4319) );
  NAND2_X1 U4365 ( .A1(n4319), .A2(n3576), .ZN(n3551) );
  INV_X1 U4366 ( .A(n3545), .ZN(n3546) );
  OAI21_X1 U4367 ( .B1(n3546), .B2(n3558), .A(n4211), .ZN(n4375) );
  INV_X1 U4368 ( .A(n4375), .ZN(n3549) );
  INV_X1 U4369 ( .A(REG2_REG_13__SCAN_IN), .ZN(n3547) );
  OAI22_X1 U4370 ( .A1(n3576), .A2(n3547), .B1(n3566), .B2(n4213), .ZN(n3548)
         );
  AOI21_X1 U4371 ( .B1(n3549), .B2(n4563), .A(n3548), .ZN(n3550) );
  OAI211_X1 U4372 ( .C1(n4318), .C2(n4221), .A(n3551), .B(n3550), .ZN(U3277)
         );
  INV_X1 U4373 ( .A(n3553), .ZN(n3555) );
  NOR2_X1 U4374 ( .A1(n3555), .A2(n3554), .ZN(n3556) );
  XNOR2_X1 U4375 ( .A(n3552), .B(n3556), .ZN(n3557) );
  NAND2_X1 U4376 ( .A1(n3557), .A2(n4405), .ZN(n3565) );
  OAI22_X1 U4377 ( .A1(n3733), .A2(n3558), .B1(n3731), .B2(n3720), .ZN(n3563)
         );
  INV_X1 U4378 ( .A(REG3_REG_13__SCAN_IN), .ZN(n3559) );
  NOR2_X1 U4379 ( .A1(STATE_REG_SCAN_IN), .A2(n3559), .ZN(n4498) );
  INV_X1 U4380 ( .A(n4498), .ZN(n3560) );
  OAI21_X1 U4381 ( .B1(n3722), .B2(n3561), .A(n3560), .ZN(n3562) );
  NOR2_X1 U4382 ( .A1(n3563), .A2(n3562), .ZN(n3564) );
  OAI211_X1 U4383 ( .C1(n4410), .C2(n3566), .A(n3565), .B(n3564), .ZN(U3231)
         );
  NOR2_X1 U4384 ( .A1(n3568), .A2(n3567), .ZN(n4200) );
  NAND2_X1 U4385 ( .A1(n4200), .A2(n3031), .ZN(n4199) );
  NAND2_X1 U4386 ( .A1(n4199), .A2(n3569), .ZN(n3570) );
  XNOR2_X1 U4387 ( .A(n3570), .B(n3743), .ZN(n4312) );
  INV_X1 U4388 ( .A(n4312), .ZN(n3580) );
  NAND2_X1 U4389 ( .A1(n4204), .A2(n3830), .ZN(n3571) );
  XNOR2_X1 U4390 ( .A(n3571), .B(n3743), .ZN(n3574) );
  OAI22_X1 U4391 ( .A1(n3735), .A2(n4574), .B1(n4255), .B2(n3732), .ZN(n3572)
         );
  AOI21_X1 U4392 ( .B1(n4227), .B2(n3904), .A(n3572), .ZN(n3573) );
  OAI21_X1 U4393 ( .B1(n3574), .B2(n4236), .A(n3573), .ZN(n4311) );
  INV_X1 U4394 ( .A(n3575), .ZN(n4192) );
  OAI21_X1 U4395 ( .B1(n2273), .B2(n3732), .A(n4192), .ZN(n4366) );
  NOR2_X1 U4396 ( .A1(n4366), .A2(n4175), .ZN(n3578) );
  OAI22_X1 U4397 ( .A1(n3576), .A2(n3950), .B1(n3740), .B2(n4213), .ZN(n3577)
         );
  AOI211_X1 U4398 ( .C1(n4311), .C2(n3576), .A(n3578), .B(n3577), .ZN(n3579)
         );
  OAI21_X1 U4399 ( .B1(n3580), .B2(n4180), .A(n3579), .ZN(U3275) );
  XNOR2_X1 U4400 ( .A(n3582), .B(n3581), .ZN(n3583) );
  XNOR2_X1 U4401 ( .A(n3584), .B(n3583), .ZN(n3585) );
  NAND2_X1 U4402 ( .A1(n3585), .A2(n4405), .ZN(n3590) );
  OAI22_X1 U4403 ( .A1(n3733), .A2(n4201), .B1(n3586), .B2(n3722), .ZN(n3588)
         );
  NAND2_X1 U4404 ( .A1(REG3_REG_14__SCAN_IN), .A2(U3149), .ZN(n4513) );
  OAI21_X1 U4405 ( .B1(n3720), .B2(n4394), .A(n4513), .ZN(n3587) );
  NOR2_X1 U4406 ( .A1(n3588), .A2(n3587), .ZN(n3589) );
  OAI211_X1 U4407 ( .C1(n4410), .C2(n4214), .A(n3590), .B(n3589), .ZN(U3212)
         );
  INV_X1 U4408 ( .A(DATAI_24_), .ZN(n4771) );
  NAND2_X1 U4409 ( .A1(n2954), .A2(STATE_REG_SCAN_IN), .ZN(n3591) );
  OAI21_X1 U4410 ( .B1(STATE_REG_SCAN_IN), .B2(n4771), .A(n3591), .ZN(U3328)
         );
  INV_X1 U4411 ( .A(n3996), .ZN(n4014) );
  AND2_X1 U4412 ( .A1(n4014), .A2(n3721), .ZN(n3596) );
  OR2_X1 U4413 ( .A1(n3592), .A2(n3596), .ZN(n3983) );
  NOR2_X1 U4414 ( .A1(n3971), .A2(n3995), .ZN(n3597) );
  OR2_X1 U4415 ( .A1(n3983), .A2(n3597), .ZN(n3600) );
  NAND2_X1 U4416 ( .A1(n3996), .A2(n3604), .ZN(n3594) );
  AND2_X1 U4417 ( .A1(n3594), .A2(n3593), .ZN(n3595) );
  OR2_X1 U4418 ( .A1(n3597), .A2(n3982), .ZN(n3599) );
  NAND2_X1 U4419 ( .A1(n3971), .A2(n3995), .ZN(n3598) );
  OR2_X1 U4420 ( .A1(n3990), .A2(n3968), .ZN(n3876) );
  NAND2_X1 U4421 ( .A1(n3990), .A2(n3968), .ZN(n3845) );
  INV_X1 U4422 ( .A(n3968), .ZN(n3975) );
  NAND2_X1 U4423 ( .A1(n3741), .A2(DATAI_29_), .ZN(n3602) );
  XNOR2_X1 U4424 ( .A(n3969), .B(n3602), .ZN(n3778) );
  XNOR2_X1 U4425 ( .A(n3601), .B(n3778), .ZN(n4261) );
  INV_X1 U4426 ( .A(n3602), .ZN(n3855) );
  NOR2_X2 U4427 ( .A1(n3986), .A2(n3975), .ZN(n3974) );
  INV_X1 U4428 ( .A(n3974), .ZN(n3603) );
  AND2_X2 U4429 ( .A1(n3974), .A2(n3602), .ZN(n4249) );
  AOI21_X1 U4430 ( .B1(n3855), .B2(n3603), .A(n4249), .ZN(n4260) );
  AOI22_X1 U4431 ( .A1(n4260), .A2(n4563), .B1(REG2_REG_29__SCAN_IN), .B2(
        n4581), .ZN(n3613) );
  NAND2_X1 U4432 ( .A1(n4014), .A2(n3604), .ZN(n3605) );
  AND2_X1 U4433 ( .A1(n3996), .A2(n3721), .ZN(n3881) );
  XNOR2_X1 U4434 ( .A(n3779), .B(n3616), .ZN(n3993) );
  NAND2_X1 U4435 ( .A1(n3779), .A2(n3995), .ZN(n3875) );
  NAND2_X1 U4436 ( .A1(n3991), .A2(n3875), .ZN(n3967) );
  INV_X1 U4437 ( .A(n3876), .ZN(n3852) );
  AOI21_X1 U4438 ( .B1(n3967), .B2(n3845), .A(n3852), .ZN(n3607) );
  AOI21_X1 U4439 ( .B1(B_REG_SCAN_IN), .B2(n4419), .A(n4574), .ZN(n4244) );
  AOI22_X1 U4440 ( .A1(n3751), .A2(n4244), .B1(n4055), .B2(n3855), .ZN(n3609)
         );
  NAND2_X1 U4441 ( .A1(n3990), .A2(n4188), .ZN(n3608) );
  NOR2_X1 U4442 ( .A1(n3610), .A2(n4213), .ZN(n3611) );
  OAI21_X1 U4443 ( .B1(n4259), .B2(n3611), .A(n3576), .ZN(n3612) );
  OAI211_X1 U4444 ( .C1(n4261), .C2(n4180), .A(n3613), .B(n3612), .ZN(U3354)
         );
  XNOR2_X1 U4445 ( .A(n3615), .B(n3614), .ZN(n3623) );
  OAI22_X1 U4446 ( .A1(n3733), .A2(n3616), .B1(n4014), .B2(n3722), .ZN(n3617)
         );
  INV_X1 U4447 ( .A(n3617), .ZN(n3620) );
  AOI22_X1 U4448 ( .A1(n3990), .A2(n3618), .B1(REG3_REG_27__SCAN_IN), .B2(
        U3149), .ZN(n3619) );
  OAI211_X1 U4449 ( .C1(n4410), .C2(n3987), .A(n3620), .B(n3619), .ZN(n3621)
         );
  INV_X1 U4450 ( .A(n3621), .ZN(n3622) );
  OAI21_X1 U4451 ( .B1(n3623), .B2(n3704), .A(n3622), .ZN(U3211) );
  INV_X1 U4452 ( .A(n3624), .ZN(n3695) );
  OAI21_X1 U4453 ( .B1(n3695), .B2(n3626), .A(n3625), .ZN(n3628) );
  NAND3_X1 U4454 ( .A1(n3628), .A2(n4405), .A3(n3627), .ZN(n3633) );
  OAI22_X1 U4455 ( .A1(n3733), .A2(n4061), .B1(n4089), .B2(n3722), .ZN(n3631)
         );
  OAI22_X1 U4456 ( .A1(n3720), .A2(n4059), .B1(STATE_REG_SCAN_IN), .B2(n3629), 
        .ZN(n3630) );
  NOR2_X1 U4457 ( .A1(n3631), .A2(n3630), .ZN(n3632) );
  OAI211_X1 U4458 ( .C1(n4410), .C2(n4063), .A(n3633), .B(n3632), .ZN(U3213)
         );
  OAI21_X1 U4459 ( .B1(n3636), .B2(n3635), .A(n3634), .ZN(n3637) );
  NAND2_X1 U4460 ( .A1(n3637), .A2(n4405), .ZN(n3641) );
  INV_X1 U4461 ( .A(n4091), .ZN(n4131) );
  OAI22_X1 U4462 ( .A1(n3733), .A2(n4138), .B1(n4131), .B2(n3720), .ZN(n3639)
         );
  NAND2_X1 U4463 ( .A1(U3149), .A2(REG3_REG_19__SCAN_IN), .ZN(n3958) );
  OAI21_X1 U4464 ( .B1(n3722), .B2(n3038), .A(n3958), .ZN(n3638) );
  NOR2_X1 U4465 ( .A1(n3639), .A2(n3638), .ZN(n3640) );
  OAI211_X1 U4466 ( .C1(n4410), .C2(n4139), .A(n3641), .B(n3640), .ZN(U3216)
         );
  INV_X1 U4467 ( .A(n3642), .ZN(n3644) );
  NAND2_X1 U4468 ( .A1(n3644), .A2(n3643), .ZN(n3647) );
  OAI211_X1 U4469 ( .C1(n3645), .C2(n2458), .A(n3688), .B(n3647), .ZN(n3646)
         );
  OAI211_X1 U4470 ( .C1(n3648), .C2(n3647), .A(n4405), .B(n3646), .ZN(n3653)
         );
  OAI22_X1 U4471 ( .A1(n3733), .A2(n4094), .B1(n4131), .B2(n3722), .ZN(n3651)
         );
  OAI22_X1 U4472 ( .A1(n3720), .A2(n4089), .B1(STATE_REG_SCAN_IN), .B2(n3649), 
        .ZN(n3650) );
  NOR2_X1 U4473 ( .A1(n3651), .A2(n3650), .ZN(n3652) );
  OAI211_X1 U4474 ( .C1(n4410), .C2(n4097), .A(n3653), .B(n3652), .ZN(U3220)
         );
  INV_X1 U4475 ( .A(n4022), .ZN(n3663) );
  NAND2_X1 U4476 ( .A1(n2264), .A2(n3654), .ZN(n3655) );
  XNOR2_X1 U4477 ( .A(n3656), .B(n3655), .ZN(n3657) );
  NAND2_X1 U4478 ( .A1(n3657), .A2(n4405), .ZN(n3662) );
  OAI22_X1 U4479 ( .A1(n3733), .A2(n4021), .B1(n4014), .B2(n3720), .ZN(n3660)
         );
  OAI22_X1 U4480 ( .A1(n3722), .A2(n4059), .B1(STATE_REG_SCAN_IN), .B2(n3658), 
        .ZN(n3659) );
  NOR2_X1 U4481 ( .A1(n3660), .A2(n3659), .ZN(n3661) );
  OAI211_X1 U4482 ( .C1(n4410), .C2(n3663), .A(n3662), .B(n3661), .ZN(U3222)
         );
  XOR2_X1 U4483 ( .A(n3666), .B(n3665), .Z(n3667) );
  XNOR2_X1 U4484 ( .A(n3664), .B(n3667), .ZN(n3668) );
  NAND2_X1 U4485 ( .A1(n3668), .A2(n4405), .ZN(n3673) );
  OAI22_X1 U4486 ( .A1(n3733), .A2(n4173), .B1(n3038), .B2(n3720), .ZN(n3671)
         );
  NOR2_X1 U4487 ( .A1(STATE_REG_SCAN_IN), .A2(n2803), .ZN(n4536) );
  INV_X1 U4488 ( .A(n4536), .ZN(n3669) );
  OAI21_X1 U4489 ( .B1(n3722), .B2(n3735), .A(n3669), .ZN(n3670) );
  NOR2_X1 U4490 ( .A1(n3671), .A2(n3670), .ZN(n3672) );
  OAI211_X1 U4491 ( .C1(n4410), .C2(n4176), .A(n3673), .B(n3672), .ZN(U3225)
         );
  INV_X1 U4492 ( .A(n4040), .ZN(n3685) );
  NAND2_X1 U4493 ( .A1(n3675), .A2(n3674), .ZN(n3677) );
  XNOR2_X1 U4494 ( .A(n3677), .B(n3676), .ZN(n3678) );
  NAND2_X1 U4495 ( .A1(n3678), .A2(n4405), .ZN(n3684) );
  OAI22_X1 U4496 ( .A1(n3733), .A2(n3679), .B1(n4036), .B2(n3720), .ZN(n3682)
         );
  INV_X1 U4497 ( .A(n4072), .ZN(n3699) );
  OAI22_X1 U4498 ( .A1(n3722), .A2(n3699), .B1(STATE_REG_SCAN_IN), .B2(n3680), 
        .ZN(n3681) );
  NOR2_X1 U4499 ( .A1(n3682), .A2(n3681), .ZN(n3683) );
  OAI211_X1 U4500 ( .C1(n4410), .C2(n3685), .A(n3684), .B(n3683), .ZN(U3226)
         );
  NOR2_X1 U4501 ( .A1(n3686), .A2(n2458), .ZN(n3690) );
  AOI21_X1 U4502 ( .B1(n3688), .B2(n3687), .A(n3645), .ZN(n3689) );
  OAI21_X1 U4503 ( .B1(n3690), .B2(n3689), .A(n4405), .ZN(n3694) );
  OAI22_X1 U4504 ( .A1(n3733), .A2(n4114), .B1(n4104), .B2(n3720), .ZN(n3692)
         );
  OAI22_X1 U4505 ( .A1(n3722), .A2(n4146), .B1(STATE_REG_SCAN_IN), .B2(n4867), 
        .ZN(n3691) );
  NOR2_X1 U4506 ( .A1(n3692), .A2(n3691), .ZN(n3693) );
  OAI211_X1 U4507 ( .C1(n4410), .C2(n4117), .A(n3694), .B(n3693), .ZN(U3230)
         );
  AOI21_X1 U4508 ( .B1(n3697), .B2(n3696), .A(n3695), .ZN(n3705) );
  OAI22_X1 U4509 ( .A1(n3733), .A2(n4081), .B1(n4104), .B2(n3722), .ZN(n3701)
         );
  OAI22_X1 U4510 ( .A1(n3720), .A2(n3699), .B1(STATE_REG_SCAN_IN), .B2(n3698), 
        .ZN(n3700) );
  NOR2_X1 U4511 ( .A1(n3701), .A2(n3700), .ZN(n3703) );
  OR2_X1 U4512 ( .A1(n4410), .A2(n4078), .ZN(n3702) );
  OAI211_X1 U4513 ( .C1(n3705), .C2(n3704), .A(n3703), .B(n3702), .ZN(U3232)
         );
  NAND2_X1 U4514 ( .A1(n2274), .A2(n3707), .ZN(n3708) );
  XNOR2_X1 U4515 ( .A(n3706), .B(n3708), .ZN(n3709) );
  NAND2_X1 U4516 ( .A1(n3709), .A2(n4405), .ZN(n3713) );
  OAI22_X1 U4517 ( .A1(n3733), .A2(n4145), .B1(n4146), .B2(n3720), .ZN(n3711)
         );
  NAND2_X1 U4518 ( .A1(U3149), .A2(REG3_REG_18__SCAN_IN), .ZN(n4559) );
  OAI21_X1 U4519 ( .B1(n3722), .B2(n4398), .A(n4559), .ZN(n3710) );
  NOR2_X1 U4520 ( .A1(n3711), .A2(n3710), .ZN(n3712) );
  OAI211_X1 U4521 ( .C1(n4410), .C2(n4160), .A(n3713), .B(n3712), .ZN(U3235)
         );
  INV_X1 U4522 ( .A(n3714), .ZN(n3716) );
  NOR2_X1 U4523 ( .A1(n3716), .A2(n3715), .ZN(n3717) );
  XNOR2_X1 U4524 ( .A(n3718), .B(n3717), .ZN(n3719) );
  NAND2_X1 U4525 ( .A1(n3719), .A2(n4405), .ZN(n3726) );
  OAI22_X1 U4526 ( .A1(n3733), .A2(n3721), .B1(n3779), .B2(n3720), .ZN(n3724)
         );
  OAI22_X1 U4527 ( .A1(n3722), .A2(n4036), .B1(STATE_REG_SCAN_IN), .B2(n4852), 
        .ZN(n3723) );
  NOR2_X1 U4528 ( .A1(n3724), .A2(n3723), .ZN(n3725) );
  OAI211_X1 U4529 ( .C1(n4410), .C2(n4004), .A(n3726), .B(n3725), .ZN(U3237)
         );
  NAND2_X1 U4530 ( .A1(n3727), .A2(n3728), .ZN(n3729) );
  XNOR2_X1 U4531 ( .A(n3729), .B(n4401), .ZN(n3730) );
  NAND2_X1 U4532 ( .A1(n3730), .A2(n4405), .ZN(n3739) );
  OAI22_X1 U4533 ( .A1(n3733), .A2(n3732), .B1(n3731), .B2(n3722), .ZN(n3737)
         );
  NOR2_X1 U4534 ( .A1(STATE_REG_SCAN_IN), .A2(n2763), .ZN(n4520) );
  INV_X1 U4535 ( .A(n4520), .ZN(n3734) );
  OAI21_X1 U4536 ( .B1(n3720), .B2(n3735), .A(n3734), .ZN(n3736) );
  NOR2_X1 U4537 ( .A1(n3737), .A2(n3736), .ZN(n3738) );
  OAI211_X1 U4538 ( .C1(n4410), .C2(n3740), .A(n3739), .B(n3738), .ZN(U3238)
         );
  NAND2_X1 U4539 ( .A1(n3741), .A2(DATAI_30_), .ZN(n4256) );
  NAND2_X1 U4540 ( .A1(n3751), .A2(n4256), .ZN(n3887) );
  NAND2_X1 U4541 ( .A1(n3741), .A2(DATAI_31_), .ZN(n4246) );
  OR2_X1 U4542 ( .A1(n4245), .A2(n4246), .ZN(n3742) );
  NAND2_X1 U4543 ( .A1(n3887), .A2(n3742), .ZN(n3858) );
  INV_X1 U4544 ( .A(n3858), .ZN(n3895) );
  INV_X1 U4545 ( .A(n3743), .ZN(n3744) );
  AND4_X1 U4546 ( .A1(n3745), .A2(n4182), .A3(n4206), .A4(n3744), .ZN(n3777)
         );
  NAND4_X1 U4547 ( .A1(n3749), .A2(n3748), .A3(n3747), .A4(n3746), .ZN(n3765)
         );
  NAND2_X1 U4548 ( .A1(n3750), .A2(n4569), .ZN(n3784) );
  AND2_X1 U4549 ( .A1(n3782), .A2(n3784), .ZN(n4570) );
  NAND2_X1 U4550 ( .A1(n4245), .A2(n4246), .ZN(n3859) );
  OR2_X1 U4551 ( .A1(n3751), .A2(n4256), .ZN(n3752) );
  AND2_X1 U4552 ( .A1(n3859), .A2(n3752), .ZN(n3853) );
  NOR2_X1 U4553 ( .A1(n3753), .A2(n3780), .ZN(n4031) );
  XNOR2_X1 U4554 ( .A(n4072), .B(n4054), .ZN(n4051) );
  INV_X1 U4555 ( .A(n3838), .ZN(n4048) );
  AND2_X1 U4556 ( .A1(n4048), .A2(n4046), .ZN(n4088) );
  NAND4_X1 U4557 ( .A1(n4049), .A2(n4031), .A3(n4051), .A4(n4088), .ZN(n3761)
         );
  AND2_X1 U4558 ( .A1(n3754), .A2(n3781), .ZN(n4013) );
  NAND4_X1 U4559 ( .A1(n3993), .A2(n3964), .A3(n4013), .A4(n3755), .ZN(n3760)
         );
  XNOR2_X1 U4560 ( .A(n4112), .B(n4138), .ZN(n4130) );
  INV_X1 U4561 ( .A(n4125), .ZN(n3756) );
  NAND2_X1 U4562 ( .A1(n3756), .A2(n4124), .ZN(n4167) );
  NAND2_X1 U4563 ( .A1(n3758), .A2(n3757), .ZN(n4103) );
  INV_X1 U4564 ( .A(n4103), .ZN(n4107) );
  OR4_X1 U4565 ( .A1(n4153), .A2(n4130), .A3(n4167), .A4(n4107), .ZN(n3759) );
  NOR3_X1 U4566 ( .A1(n3761), .A2(n3760), .A3(n3759), .ZN(n3763) );
  NAND4_X1 U4567 ( .A1(n4570), .A2(n3853), .A3(n3763), .A4(n3762), .ZN(n3764)
         );
  NOR2_X1 U4568 ( .A1(n3765), .A2(n3764), .ZN(n3776) );
  NAND4_X1 U4569 ( .A1(n3768), .A2(n3767), .A3(n3802), .A4(n3766), .ZN(n3774)
         );
  INV_X1 U4570 ( .A(n3053), .ZN(n3772) );
  NAND4_X1 U4571 ( .A1(n3772), .A2(n3771), .A3(n3770), .A4(n3769), .ZN(n3773)
         );
  NOR2_X1 U4572 ( .A1(n3774), .A2(n3773), .ZN(n3775) );
  AND4_X1 U4573 ( .A1(n3778), .A2(n3777), .A3(n3776), .A4(n3775), .ZN(n3850)
         );
  NOR2_X1 U4574 ( .A1(n3779), .A2(n3995), .ZN(n3847) );
  AND2_X1 U4575 ( .A1(n2306), .A2(n3781), .ZN(n3872) );
  INV_X1 U4576 ( .A(n3782), .ZN(n3786) );
  OAI211_X1 U4577 ( .C1(n3786), .C2(n3785), .A(n3784), .B(n3783), .ZN(n3789)
         );
  NAND3_X1 U4578 ( .A1(n3789), .A2(n3788), .A3(n3787), .ZN(n3792) );
  NAND3_X1 U4579 ( .A1(n3792), .A2(n3791), .A3(n3790), .ZN(n3795) );
  NAND3_X1 U4580 ( .A1(n3795), .A2(n3794), .A3(n3793), .ZN(n3799) );
  NAND4_X1 U4581 ( .A1(n3799), .A2(n3798), .A3(n3797), .A4(n3796), .ZN(n3803)
         );
  INV_X1 U4582 ( .A(n3800), .ZN(n3801) );
  NAND3_X1 U4583 ( .A1(n3803), .A2(n3802), .A3(n3801), .ZN(n3810) );
  AND2_X1 U4584 ( .A1(n3805), .A2(n3804), .ZN(n3813) );
  INV_X1 U4585 ( .A(n3806), .ZN(n3809) );
  INV_X1 U4586 ( .A(n3807), .ZN(n3808) );
  AOI211_X1 U4587 ( .C1(n3810), .C2(n3813), .A(n3809), .B(n3808), .ZN(n3821)
         );
  NAND2_X1 U4588 ( .A1(n3812), .A2(n3811), .ZN(n3820) );
  INV_X1 U4589 ( .A(n3813), .ZN(n3816) );
  NOR3_X1 U4590 ( .A1(n3816), .A2(n3815), .A3(n3814), .ZN(n3818) );
  INV_X1 U4591 ( .A(n3822), .ZN(n3817) );
  NAND2_X1 U4592 ( .A1(n3820), .A2(n3829), .ZN(n3860) );
  OAI21_X1 U4593 ( .B1(n3818), .B2(n3817), .A(n3860), .ZN(n3819) );
  OAI21_X1 U4594 ( .B1(n3821), .B2(n3820), .A(n3819), .ZN(n3827) );
  NAND2_X1 U4595 ( .A1(n3823), .A2(n3822), .ZN(n3824) );
  NAND4_X1 U4596 ( .A1(n3827), .A2(n3826), .A3(n3825), .A4(n3824), .ZN(n3834)
         );
  INV_X1 U4597 ( .A(n3828), .ZN(n3831) );
  NAND2_X1 U4598 ( .A1(n3830), .A2(n3829), .ZN(n3861) );
  OAI21_X1 U4599 ( .B1(n3831), .B2(n3861), .A(n3860), .ZN(n3833) );
  AOI21_X1 U4600 ( .B1(n3834), .B2(n3833), .A(n2314), .ZN(n3837) );
  INV_X1 U4601 ( .A(n3863), .ZN(n3836) );
  INV_X1 U4602 ( .A(n3862), .ZN(n3835) );
  OAI21_X1 U4603 ( .B1(n3837), .B2(n3836), .A(n3835), .ZN(n3839) );
  AOI211_X1 U4604 ( .C1(n3839), .C2(n3867), .A(n3866), .B(n3838), .ZN(n3840)
         );
  NOR2_X1 U4605 ( .A1(n3840), .A2(n3870), .ZN(n3842) );
  OAI21_X1 U4606 ( .B1(n3842), .B2(n3841), .A(n3874), .ZN(n3844) );
  INV_X1 U4607 ( .A(n3878), .ZN(n3843) );
  AOI21_X1 U4608 ( .B1(n3872), .B2(n3844), .A(n3843), .ZN(n3846) );
  OAI21_X1 U4609 ( .B1(n3969), .B2(n3855), .A(n3845), .ZN(n3879) );
  NOR4_X1 U4610 ( .A1(n3847), .A2(n3881), .A3(n3846), .A4(n3879), .ZN(n3849)
         );
  MUX2_X1 U4611 ( .A(n3850), .B(n3849), .S(n3848), .Z(n3894) );
  INV_X1 U4612 ( .A(n3875), .ZN(n3851) );
  NOR2_X1 U4613 ( .A1(n3852), .A2(n3851), .ZN(n3856) );
  INV_X1 U4614 ( .A(n3853), .ZN(n3854) );
  AOI21_X1 U4615 ( .B1(n3969), .B2(n3855), .A(n3854), .ZN(n3877) );
  OAI21_X1 U4616 ( .B1(n3856), .B2(n3879), .A(n3877), .ZN(n3882) );
  INV_X1 U4617 ( .A(n3882), .ZN(n3857) );
  AOI211_X1 U4618 ( .C1(n3859), .C2(n3858), .A(n2542), .B(n3857), .ZN(n3893)
         );
  OAI21_X1 U4619 ( .B1(n4205), .B2(n3861), .A(n3860), .ZN(n3864) );
  AOI211_X1 U4620 ( .C1(n3864), .C2(n3863), .A(n2314), .B(n3862), .ZN(n3865)
         );
  INV_X1 U4621 ( .A(n3865), .ZN(n3868) );
  AOI21_X1 U4622 ( .B1(n3868), .B2(n3867), .A(n3866), .ZN(n3871) );
  OAI21_X1 U4623 ( .B1(n3871), .B2(n3870), .A(n3869), .ZN(n3873) );
  AOI21_X1 U4624 ( .B1(n3874), .B2(n3873), .A(n2303), .ZN(n3885) );
  NAND4_X1 U4625 ( .A1(n3878), .A2(n3877), .A3(n3876), .A4(n3875), .ZN(n3884)
         );
  INV_X1 U4626 ( .A(n3993), .ZN(n3880) );
  NOR3_X1 U4627 ( .A1(n3881), .A2(n3880), .A3(n3879), .ZN(n3883) );
  OAI22_X1 U4628 ( .A1(n3885), .A2(n3884), .B1(n3883), .B2(n3882), .ZN(n3891)
         );
  INV_X1 U4629 ( .A(n4245), .ZN(n3886) );
  INV_X1 U4630 ( .A(n4256), .ZN(n4253) );
  NAND2_X1 U4631 ( .A1(n3886), .A2(n4253), .ZN(n3890) );
  AOI21_X1 U4632 ( .B1(n3887), .B2(n4245), .A(n4246), .ZN(n3889) );
  AOI211_X1 U4633 ( .C1(n3891), .C2(n3890), .A(n3889), .B(n3888), .ZN(n3892)
         );
  AOI211_X1 U4634 ( .C1(n3895), .C2(n3894), .A(n3893), .B(n3892), .ZN(n3896)
         );
  XNOR2_X1 U4635 ( .A(n3896), .B(n3959), .ZN(n3903) );
  NAND2_X1 U4636 ( .A1(n3898), .A2(n3897), .ZN(n3899) );
  OAI211_X1 U4637 ( .C1(n3900), .C2(n3922), .A(B_REG_SCAN_IN), .B(n3899), .ZN(
        n3901) );
  OAI21_X1 U4638 ( .B1(n3903), .B2(n3902), .A(n3901), .ZN(U3239) );
  MUX2_X1 U4639 ( .A(n3990), .B(DATAO_REG_28__SCAN_IN), .S(n3910), .Z(U3578)
         );
  MUX2_X1 U4640 ( .A(n3971), .B(DATAO_REG_27__SCAN_IN), .S(n3910), .Z(U3577)
         );
  MUX2_X1 U4641 ( .A(n3996), .B(DATAO_REG_26__SCAN_IN), .S(n3910), .Z(U3576)
         );
  MUX2_X1 U4642 ( .A(n4016), .B(DATAO_REG_24__SCAN_IN), .S(n3910), .Z(U3574)
         );
  MUX2_X1 U4643 ( .A(DATAO_REG_22__SCAN_IN), .B(n4056), .S(U4043), .Z(U3572)
         );
  MUX2_X1 U4644 ( .A(n4073), .B(DATAO_REG_21__SCAN_IN), .S(n3910), .Z(U3571)
         );
  MUX2_X1 U4645 ( .A(n4091), .B(DATAO_REG_20__SCAN_IN), .S(n3910), .Z(U3570)
         );
  MUX2_X1 U4646 ( .A(n4133), .B(DATAO_REG_18__SCAN_IN), .S(n3910), .Z(U3568)
         );
  MUX2_X1 U4647 ( .A(n4151), .B(DATAO_REG_17__SCAN_IN), .S(n3910), .Z(U3567)
         );
  MUX2_X1 U4648 ( .A(n4169), .B(DATAO_REG_16__SCAN_IN), .S(n3910), .Z(U3566)
         );
  MUX2_X1 U4649 ( .A(n4187), .B(DATAO_REG_15__SCAN_IN), .S(n3910), .Z(U3565)
         );
  MUX2_X1 U4650 ( .A(n3904), .B(DATAO_REG_14__SCAN_IN), .S(n3910), .Z(U3564)
         );
  MUX2_X1 U4651 ( .A(n3905), .B(DATAO_REG_10__SCAN_IN), .S(n3910), .Z(U3560)
         );
  MUX2_X1 U4652 ( .A(n3906), .B(DATAO_REG_9__SCAN_IN), .S(n3910), .Z(U3559) );
  MUX2_X1 U4653 ( .A(n3907), .B(DATAO_REG_8__SCAN_IN), .S(n3910), .Z(U3558) );
  MUX2_X1 U4654 ( .A(n3908), .B(DATAO_REG_6__SCAN_IN), .S(n3910), .Z(U3556) );
  MUX2_X1 U4655 ( .A(n3909), .B(DATAO_REG_4__SCAN_IN), .S(n3910), .Z(U3554) );
  MUX2_X1 U4656 ( .A(n4229), .B(DATAO_REG_3__SCAN_IN), .S(n3910), .Z(U3553) );
  MUX2_X1 U4657 ( .A(n3018), .B(DATAO_REG_1__SCAN_IN), .S(n3910), .Z(U3551) );
  OAI21_X1 U4658 ( .B1(n3913), .B2(n3912), .A(n3911), .ZN(n3914) );
  NOR2_X1 U4659 ( .A1(n4551), .A2(n3914), .ZN(n3919) );
  AOI211_X1 U4660 ( .C1(n3917), .C2(n3916), .A(n3915), .B(n4548), .ZN(n3918)
         );
  AOI211_X1 U4661 ( .C1(n5046), .C2(n3144), .A(n3919), .B(n3918), .ZN(n3928)
         );
  AOI22_X1 U4662 ( .A1(ADDR_REG_2__SCAN_IN), .A2(n5045), .B1(
        REG3_REG_2__SCAN_IN), .B2(U3149), .ZN(n3927) );
  INV_X1 U4663 ( .A(n4419), .ZN(n3920) );
  NAND3_X1 U4664 ( .A1(n3921), .A2(n4377), .A3(n3920), .ZN(n3926) );
  INV_X1 U4665 ( .A(n3922), .ZN(n3924) );
  INV_X1 U4666 ( .A(REG2_REG_0__SCAN_IN), .ZN(n4977) );
  NAND2_X1 U4667 ( .A1(n4419), .A2(n4977), .ZN(n3923) );
  NAND2_X1 U4668 ( .A1(n4377), .A2(n3923), .ZN(n4417) );
  AOI22_X1 U4669 ( .A1(n3924), .A2(n5044), .B1(n5035), .B2(n4417), .ZN(n3925)
         );
  NAND3_X1 U4670 ( .A1(n3926), .A2(U4043), .A3(n3925), .ZN(n4433) );
  NAND3_X1 U4671 ( .A1(n3928), .A2(n3927), .A3(n4433), .ZN(U3242) );
  AOI22_X1 U4672 ( .A1(n3954), .A2(REG1_REG_17__SCAN_IN), .B1(n4304), .B2(
        n4586), .ZN(n4539) );
  INV_X1 U4673 ( .A(n3929), .ZN(n3931) );
  NOR2_X1 U4674 ( .A1(n3931), .A2(n3930), .ZN(n4496) );
  INV_X1 U4675 ( .A(n4499), .ZN(n4590) );
  AOI22_X1 U4676 ( .A1(REG1_REG_13__SCAN_IN), .A2(n4590), .B1(n4499), .B2(
        n4321), .ZN(n4495) );
  NOR2_X1 U4677 ( .A1(n4496), .A2(n4495), .ZN(n4494) );
  AND2_X1 U4678 ( .A1(n4499), .A2(REG1_REG_13__SCAN_IN), .ZN(n3932) );
  NAND2_X1 U4679 ( .A1(n3934), .A2(n4512), .ZN(n3933) );
  INV_X1 U4680 ( .A(n3933), .ZN(n3935) );
  OAI21_X1 U4681 ( .B1(n3934), .B2(n4512), .A(n3933), .ZN(n4509) );
  INV_X1 U4682 ( .A(n3951), .ZN(n4589) );
  AOI22_X1 U4683 ( .A1(REG1_REG_15__SCAN_IN), .A2(n4589), .B1(n3951), .B2(
        n4313), .ZN(n4522) );
  INV_X1 U4684 ( .A(n3937), .ZN(n3936) );
  NAND2_X1 U4685 ( .A1(n3936), .A2(n4587), .ZN(n3938) );
  NAND2_X1 U4686 ( .A1(n4529), .A2(n4528), .ZN(n4527) );
  NAND2_X1 U4687 ( .A1(n3938), .A2(n4527), .ZN(n4538) );
  NAND2_X1 U4688 ( .A1(n4554), .A2(REG1_REG_18__SCAN_IN), .ZN(n3940) );
  OR2_X1 U4689 ( .A1(n4554), .A2(REG1_REG_18__SCAN_IN), .ZN(n3939) );
  NAND2_X1 U4690 ( .A1(n3940), .A2(n3939), .ZN(n4549) );
  XNOR2_X1 U4691 ( .A(n3959), .B(REG1_REG_19__SCAN_IN), .ZN(n3941) );
  XNOR2_X1 U4692 ( .A(n3942), .B(n3941), .ZN(n3963) );
  NOR2_X1 U4693 ( .A1(n3954), .A2(REG2_REG_17__SCAN_IN), .ZN(n3943) );
  AOI21_X1 U4694 ( .B1(REG2_REG_17__SCAN_IN), .B2(n3954), .A(n3943), .ZN(n4542) );
  NAND2_X1 U4695 ( .A1(n4381), .A2(n3944), .ZN(n3946) );
  NAND2_X1 U4696 ( .A1(n4499), .A2(REG2_REG_13__SCAN_IN), .ZN(n3947) );
  NOR2_X1 U4697 ( .A1(n3949), .A2(n4505), .ZN(n4518) );
  AOI22_X1 U4698 ( .A1(REG2_REG_15__SCAN_IN), .A2(n4589), .B1(n3951), .B2(
        n3950), .ZN(n4517) );
  NAND2_X1 U4699 ( .A1(n3952), .A2(n4587), .ZN(n3953) );
  NAND2_X1 U4700 ( .A1(n3953), .A2(n4530), .ZN(n4541) );
  XNOR2_X1 U4701 ( .A(n4554), .B(REG2_REG_18__SCAN_IN), .ZN(n4552) );
  XNOR2_X1 U4702 ( .A(n3959), .B(REG2_REG_19__SCAN_IN), .ZN(n3955) );
  XNOR2_X1 U4703 ( .A(n3956), .B(n3955), .ZN(n3961) );
  NAND2_X1 U4704 ( .A1(n5045), .A2(ADDR_REG_19__SCAN_IN), .ZN(n3957) );
  OAI211_X1 U4705 ( .C1(n4547), .C2(n3959), .A(n3958), .B(n3957), .ZN(n3960)
         );
  AOI21_X1 U4706 ( .B1(n3961), .B2(n5042), .A(n3960), .ZN(n3962) );
  OAI21_X1 U4707 ( .B1(n3963), .B2(n4548), .A(n3962), .ZN(U3259) );
  XNOR2_X1 U4708 ( .A(n3965), .B(n3964), .ZN(n4263) );
  INV_X1 U4709 ( .A(n4263), .ZN(n3981) );
  XNOR2_X1 U4710 ( .A(n3967), .B(n3966), .ZN(n3973) );
  OAI22_X1 U4711 ( .A1(n3969), .A2(n4574), .B1(n4255), .B2(n3968), .ZN(n3970)
         );
  AOI21_X1 U4712 ( .B1(n4227), .B2(n3971), .A(n3970), .ZN(n3972) );
  OAI21_X1 U4713 ( .B1(n3973), .B2(n4236), .A(n3972), .ZN(n4262) );
  AOI21_X1 U4714 ( .B1(n3975), .B2(n3986), .A(n3974), .ZN(n4330) );
  INV_X1 U4715 ( .A(n4330), .ZN(n3978) );
  AOI22_X1 U4716 ( .A1(n4581), .A2(REG2_REG_28__SCAN_IN), .B1(n3976), .B2(
        n4577), .ZN(n3977) );
  OAI21_X1 U4717 ( .B1(n3978), .B2(n4175), .A(n3977), .ZN(n3979) );
  AOI21_X1 U4718 ( .B1(n4262), .B2(n3576), .A(n3979), .ZN(n3980) );
  OAI21_X1 U4719 ( .B1(n3981), .B2(n4180), .A(n3980), .ZN(U3262) );
  XNOR2_X1 U4720 ( .A(n3985), .B(n3993), .ZN(n4270) );
  AOI21_X1 U4721 ( .B1(n3995), .B2(n2245), .A(n2377), .ZN(n4268) );
  INV_X1 U4723 ( .A(REG2_REG_27__SCAN_IN), .ZN(n3988) );
  OAI22_X1 U4724 ( .A1(n3576), .A2(n3988), .B1(n3987), .B2(n4213), .ZN(n3989)
         );
  AOI21_X1 U4725 ( .B1(n4268), .B2(n4563), .A(n3989), .ZN(n4001) );
  INV_X1 U4726 ( .A(n3990), .ZN(n3999) );
  OAI21_X1 U4727 ( .B1(n3993), .B2(n3992), .A(n3991), .ZN(n3994) );
  NAND2_X1 U4728 ( .A1(n3994), .A2(n4571), .ZN(n3998) );
  AOI22_X1 U4729 ( .A1(n3996), .A2(n4227), .B1(n4055), .B2(n3995), .ZN(n3997)
         );
  OAI211_X1 U4730 ( .C1(n3999), .C2(n4574), .A(n3998), .B(n3997), .ZN(n4267)
         );
  NAND2_X1 U4731 ( .A1(n4267), .A2(n3576), .ZN(n4000) );
  OAI211_X1 U4732 ( .C1(n4270), .C2(n4180), .A(n4001), .B(n4000), .ZN(U3263)
         );
  INV_X1 U4733 ( .A(n4002), .ZN(n4010) );
  NOR2_X1 U4734 ( .A1(n4003), .A2(n4175), .ZN(n4007) );
  OAI22_X1 U4735 ( .A1(n3576), .A2(n4005), .B1(n4004), .B2(n4213), .ZN(n4006)
         );
  AOI211_X1 U4736 ( .C1(n4008), .C2(n3576), .A(n4007), .B(n4006), .ZN(n4009)
         );
  OAI21_X1 U4737 ( .B1(n4010), .B2(n4180), .A(n4009), .ZN(U3264) );
  XOR2_X1 U4738 ( .A(n4013), .B(n4011), .Z(n4272) );
  INV_X1 U4739 ( .A(n4272), .ZN(n4026) );
  XOR2_X1 U4740 ( .A(n4013), .B(n4012), .Z(n4018) );
  OAI22_X1 U4741 ( .A1(n4014), .A2(n4574), .B1(n4255), .B2(n4021), .ZN(n4015)
         );
  AOI21_X1 U4742 ( .B1(n4227), .B2(n4016), .A(n4015), .ZN(n4017) );
  OAI21_X1 U4743 ( .B1(n4018), .B2(n4236), .A(n4017), .ZN(n4271) );
  INV_X1 U4744 ( .A(n4019), .ZN(n4020) );
  OAI21_X1 U4745 ( .B1(n4038), .B2(n4021), .A(n4020), .ZN(n4337) );
  AOI22_X1 U4746 ( .A1(n4581), .A2(REG2_REG_25__SCAN_IN), .B1(n4022), .B2(
        n4577), .ZN(n4023) );
  OAI21_X1 U4747 ( .B1(n4337), .B2(n4175), .A(n4023), .ZN(n4024) );
  AOI21_X1 U4748 ( .B1(n4271), .B2(n3576), .A(n4024), .ZN(n4025) );
  OAI21_X1 U4749 ( .B1(n4026), .B2(n4180), .A(n4025), .ZN(U3265) );
  XNOR2_X1 U4750 ( .A(n4027), .B(n4031), .ZN(n4276) );
  INV_X1 U4751 ( .A(n4276), .ZN(n4044) );
  INV_X1 U4752 ( .A(n4028), .ZN(n4029) );
  NAND2_X1 U4753 ( .A1(n4030), .A2(n4029), .ZN(n4032) );
  XNOR2_X1 U4754 ( .A(n4032), .B(n4031), .ZN(n4033) );
  NAND2_X1 U4755 ( .A1(n4033), .A2(n4571), .ZN(n4035) );
  AOI22_X1 U4756 ( .A1(n4072), .A2(n4188), .B1(n4055), .B2(n4037), .ZN(n4034)
         );
  OAI211_X1 U4757 ( .C1(n4036), .C2(n4574), .A(n4035), .B(n4034), .ZN(n4275)
         );
  AND2_X1 U4758 ( .A1(n4060), .A2(n4037), .ZN(n4039) );
  OR2_X1 U4759 ( .A1(n4039), .A2(n4038), .ZN(n4341) );
  AOI22_X1 U4760 ( .A1(n4581), .A2(REG2_REG_24__SCAN_IN), .B1(n4040), .B2(
        n4577), .ZN(n4041) );
  OAI21_X1 U4761 ( .B1(n4341), .B2(n4175), .A(n4041), .ZN(n4042) );
  AOI21_X1 U4762 ( .B1(n4275), .B2(n3576), .A(n4042), .ZN(n4043) );
  OAI21_X1 U4763 ( .B1(n4044), .B2(n4180), .A(n4043), .ZN(U3266) );
  XNOR2_X1 U4764 ( .A(n4045), .B(n4051), .ZN(n4279) );
  INV_X1 U4765 ( .A(n4279), .ZN(n4068) );
  INV_X1 U4766 ( .A(n4046), .ZN(n4047) );
  AOI21_X1 U4767 ( .B1(n4087), .B2(n4048), .A(n4047), .ZN(n4071) );
  OAI21_X1 U4768 ( .B1(n4071), .B2(n3045), .A(n4050), .ZN(n4052) );
  XNOR2_X1 U4769 ( .A(n4052), .B(n4051), .ZN(n4053) );
  NAND2_X1 U4770 ( .A1(n4053), .A2(n4571), .ZN(n4058) );
  AOI22_X1 U4771 ( .A1(n4056), .A2(n4188), .B1(n4055), .B2(n4054), .ZN(n4057)
         );
  OAI211_X1 U4772 ( .C1(n4059), .C2(n4574), .A(n4058), .B(n4057), .ZN(n4278)
         );
  INV_X1 U4773 ( .A(n4281), .ZN(n4062) );
  OAI21_X1 U4774 ( .B1(n4062), .B2(n4061), .A(n4060), .ZN(n4345) );
  NOR2_X1 U4775 ( .A1(n4345), .A2(n4175), .ZN(n4066) );
  OAI22_X1 U4776 ( .A1(n3576), .A2(n4064), .B1(n4063), .B2(n4213), .ZN(n4065)
         );
  AOI211_X1 U4777 ( .C1(n4278), .C2(n3576), .A(n4066), .B(n4065), .ZN(n4067)
         );
  OAI21_X1 U4778 ( .B1(n4068), .B2(n4180), .A(n4067), .ZN(U3267) );
  OAI21_X1 U4779 ( .B1(n4070), .B2(n3045), .A(n4069), .ZN(n4285) );
  XNOR2_X1 U4780 ( .A(n4071), .B(n3045), .ZN(n4077) );
  NAND2_X1 U4781 ( .A1(n4072), .A2(n4228), .ZN(n4075) );
  NAND2_X1 U4782 ( .A1(n4073), .A2(n4227), .ZN(n4074) );
  OAI211_X1 U4783 ( .C1(n4081), .C2(n4255), .A(n4075), .B(n4074), .ZN(n4076)
         );
  AOI21_X1 U4784 ( .B1(n4077), .B2(n4571), .A(n4076), .ZN(n4284) );
  OAI22_X1 U4785 ( .A1(n3576), .A2(n4079), .B1(n4078), .B2(n4213), .ZN(n4080)
         );
  INV_X1 U4786 ( .A(n4080), .ZN(n4083) );
  OR2_X1 U4787 ( .A1(n4096), .A2(n4081), .ZN(n4282) );
  NAND3_X1 U4788 ( .A1(n4282), .A2(n4563), .A3(n4281), .ZN(n4082) );
  OAI211_X1 U4789 ( .C1(n4284), .C2(n4581), .A(n4083), .B(n4082), .ZN(n4084)
         );
  INV_X1 U4790 ( .A(n4084), .ZN(n4085) );
  OAI21_X1 U4791 ( .B1(n4285), .B2(n4180), .A(n4085), .ZN(U3268) );
  XOR2_X1 U4792 ( .A(n4088), .B(n4086), .Z(n4287) );
  INV_X1 U4793 ( .A(n4287), .ZN(n4101) );
  XOR2_X1 U4794 ( .A(n4088), .B(n4087), .Z(n4093) );
  OAI22_X1 U4795 ( .A1(n4089), .A2(n4574), .B1(n4255), .B2(n4094), .ZN(n4090)
         );
  AOI21_X1 U4796 ( .B1(n4188), .B2(n4091), .A(n4090), .ZN(n4092) );
  OAI21_X1 U4797 ( .B1(n4093), .B2(n4236), .A(n4092), .ZN(n4286) );
  NOR2_X1 U4798 ( .A1(n4116), .A2(n4094), .ZN(n4095) );
  OR2_X1 U4799 ( .A1(n4096), .A2(n4095), .ZN(n4350) );
  NOR2_X1 U4800 ( .A1(n4350), .A2(n4175), .ZN(n4099) );
  OAI22_X1 U4801 ( .A1(n3576), .A2(n4831), .B1(n4097), .B2(n4213), .ZN(n4098)
         );
  AOI211_X1 U4802 ( .C1(n4286), .C2(n3576), .A(n4099), .B(n4098), .ZN(n4100)
         );
  OAI21_X1 U4803 ( .B1(n4101), .B2(n4180), .A(n4100), .ZN(U3269) );
  XNOR2_X1 U4804 ( .A(n4102), .B(n4103), .ZN(n4290) );
  OAI22_X1 U4805 ( .A1(n4104), .A2(n4574), .B1(n4255), .B2(n4114), .ZN(n4111)
         );
  NAND2_X1 U4806 ( .A1(n4106), .A2(n4105), .ZN(n4108) );
  XNOR2_X1 U4807 ( .A(n4108), .B(n4107), .ZN(n4109) );
  NOR2_X1 U4808 ( .A1(n4109), .A2(n4236), .ZN(n4110) );
  AOI211_X1 U4809 ( .C1(n4188), .C2(n4112), .A(n4111), .B(n4110), .ZN(n4113)
         );
  OAI21_X1 U4810 ( .B1(n4290), .B2(n4226), .A(n4113), .ZN(n4291) );
  NAND2_X1 U4811 ( .A1(n4291), .A2(n3576), .ZN(n4122) );
  NOR2_X1 U4812 ( .A1(n4136), .A2(n4114), .ZN(n4115) );
  OR2_X1 U4813 ( .A1(n4116), .A2(n4115), .ZN(n4354) );
  INV_X1 U4814 ( .A(n4354), .ZN(n4120) );
  OAI22_X1 U4815 ( .A1(n3576), .A2(n4118), .B1(n4117), .B2(n4213), .ZN(n4119)
         );
  AOI21_X1 U4816 ( .B1(n4120), .B2(n4563), .A(n4119), .ZN(n4121) );
  OAI211_X1 U4817 ( .C1(n4290), .C2(n4221), .A(n4122), .B(n4121), .ZN(U3270)
         );
  XNOR2_X1 U4818 ( .A(n4123), .B(n4130), .ZN(n4295) );
  INV_X1 U4819 ( .A(n4295), .ZN(n4144) );
  OAI21_X1 U4820 ( .B1(n4166), .B2(n4125), .A(n4124), .ZN(n4147) );
  INV_X1 U4821 ( .A(n4126), .ZN(n4128) );
  OAI21_X1 U4822 ( .B1(n4147), .B2(n4128), .A(n4127), .ZN(n4129) );
  XOR2_X1 U4823 ( .A(n4130), .B(n4129), .Z(n4135) );
  OAI22_X1 U4824 ( .A1(n4131), .A2(n4574), .B1(n4255), .B2(n4138), .ZN(n4132)
         );
  AOI21_X1 U4825 ( .B1(n4188), .B2(n4133), .A(n4132), .ZN(n4134) );
  OAI21_X1 U4826 ( .B1(n4135), .B2(n4236), .A(n4134), .ZN(n4294) );
  INV_X1 U4827 ( .A(n4136), .ZN(n4137) );
  OAI21_X1 U4828 ( .B1(n2381), .B2(n4138), .A(n4137), .ZN(n4358) );
  NOR2_X1 U4829 ( .A1(n4358), .A2(n4175), .ZN(n4142) );
  OAI22_X1 U4830 ( .A1(n3576), .A2(n4140), .B1(n4139), .B2(n4213), .ZN(n4141)
         );
  AOI211_X1 U4831 ( .C1(n4294), .C2(n3576), .A(n4142), .B(n4141), .ZN(n4143)
         );
  OAI21_X1 U4832 ( .B1(n4144), .B2(n4180), .A(n4143), .ZN(U3271) );
  OAI22_X1 U4833 ( .A1(n4146), .A2(n4574), .B1(n4255), .B2(n4145), .ZN(n4150)
         );
  XNOR2_X1 U4834 ( .A(n4147), .B(n4153), .ZN(n4148) );
  NOR2_X1 U4835 ( .A1(n4148), .A2(n4236), .ZN(n4149) );
  AOI211_X1 U4836 ( .C1(n4227), .C2(n4151), .A(n4150), .B(n4149), .ZN(n4300)
         );
  OAI21_X1 U4837 ( .B1(n4154), .B2(n4153), .A(n4152), .ZN(n4298) );
  AOI21_X1 U4838 ( .B1(n4172), .B2(n4155), .A(n4638), .ZN(n4157) );
  NAND2_X1 U4839 ( .A1(n4157), .A2(n4156), .ZN(n4299) );
  INV_X1 U4840 ( .A(n4158), .ZN(n4159) );
  NOR2_X1 U4841 ( .A1(n4299), .A2(n4159), .ZN(n4163) );
  OAI22_X1 U4842 ( .A1(n3576), .A2(n4161), .B1(n4160), .B2(n4213), .ZN(n4162)
         );
  AOI211_X1 U4843 ( .C1(n4298), .C2(n4196), .A(n4163), .B(n4162), .ZN(n4164)
         );
  OAI21_X1 U4844 ( .B1(n4581), .B2(n4300), .A(n4164), .ZN(U3272) );
  XOR2_X1 U4845 ( .A(n4167), .B(n4165), .Z(n4303) );
  INV_X1 U4846 ( .A(n4303), .ZN(n4181) );
  XOR2_X1 U4847 ( .A(n4167), .B(n4166), .Z(n4171) );
  OAI22_X1 U4848 ( .A1(n3038), .A2(n4574), .B1(n4255), .B2(n4173), .ZN(n4168)
         );
  AOI21_X1 U4849 ( .B1(n4188), .B2(n4169), .A(n4168), .ZN(n4170) );
  OAI21_X1 U4850 ( .B1(n4171), .B2(n4236), .A(n4170), .ZN(n4302) );
  INV_X1 U4851 ( .A(n4306), .ZN(n4174) );
  OAI21_X1 U4852 ( .B1(n4174), .B2(n4173), .A(n4172), .ZN(n4362) );
  NOR2_X1 U4853 ( .A1(n4362), .A2(n4175), .ZN(n4178) );
  OAI22_X1 U4854 ( .A1(n3576), .A2(n4829), .B1(n4176), .B2(n4213), .ZN(n4177)
         );
  AOI211_X1 U4855 ( .C1(n4302), .C2(n3576), .A(n4178), .B(n4177), .ZN(n4179)
         );
  OAI21_X1 U4856 ( .B1(n4181), .B2(n4180), .A(n4179), .ZN(U3273) );
  OAI22_X1 U4857 ( .A1(n4398), .A2(n4574), .B1(n4255), .B2(n4395), .ZN(n4186)
         );
  XNOR2_X1 U4858 ( .A(n4183), .B(n4182), .ZN(n4184) );
  NOR2_X1 U4859 ( .A1(n4184), .A2(n4236), .ZN(n4185) );
  AOI211_X1 U4860 ( .C1(n4188), .C2(n4187), .A(n4186), .B(n4185), .ZN(n4309)
         );
  OAI21_X1 U4861 ( .B1(n2272), .B2(n4190), .A(n4189), .ZN(n4310) );
  INV_X1 U4862 ( .A(n4310), .ZN(n4197) );
  NAND2_X1 U4863 ( .A1(n4192), .A2(n4191), .ZN(n4307) );
  AND3_X1 U4864 ( .A1(n4307), .A2(n4563), .A3(n4306), .ZN(n4195) );
  OAI22_X1 U4865 ( .A1(n3576), .A2(n4193), .B1(n4409), .B2(n4213), .ZN(n4194)
         );
  AOI211_X1 U4866 ( .C1(n4197), .C2(n4196), .A(n4195), .B(n4194), .ZN(n4198)
         );
  OAI21_X1 U4867 ( .B1(n4581), .B2(n4309), .A(n4198), .ZN(U3274) );
  OAI21_X1 U4868 ( .B1(n4200), .B2(n3031), .A(n4199), .ZN(n4316) );
  INV_X1 U4869 ( .A(n4316), .ZN(n4222) );
  OAI22_X1 U4870 ( .A1(n4394), .A2(n4574), .B1(n4255), .B2(n4201), .ZN(n4202)
         );
  AOI21_X1 U4871 ( .B1(n4227), .B2(n4203), .A(n4202), .ZN(n4209) );
  OAI21_X1 U4872 ( .B1(n4206), .B2(n4205), .A(n4204), .ZN(n4207) );
  NAND2_X1 U4873 ( .A1(n4207), .A2(n4571), .ZN(n4208) );
  OAI211_X1 U4874 ( .C1(n4222), .C2(n4226), .A(n4209), .B(n4208), .ZN(n4315)
         );
  NAND2_X1 U4875 ( .A1(n4315), .A2(n3576), .ZN(n4220) );
  AND2_X1 U4876 ( .A1(n4211), .A2(n4210), .ZN(n4212) );
  OR2_X1 U4877 ( .A1(n4212), .A2(n2273), .ZN(n4370) );
  INV_X1 U4878 ( .A(n4370), .ZN(n4218) );
  OAI22_X1 U4879 ( .A1(n3576), .A2(n4215), .B1(n4214), .B2(n4213), .ZN(n4217)
         );
  AOI21_X1 U4880 ( .B1(n4218), .B2(n4563), .A(n4217), .ZN(n4219) );
  OAI211_X1 U4881 ( .C1(n4222), .C2(n4221), .A(n4220), .B(n4219), .ZN(U3276)
         );
  XNOR2_X1 U4882 ( .A(n4223), .B(n4224), .ZN(n4237) );
  INV_X1 U4883 ( .A(n4226), .ZN(n4572) );
  NAND2_X1 U4884 ( .A1(n4613), .A2(n4572), .ZN(n4235) );
  NAND2_X1 U4885 ( .A1(n3018), .A2(n4227), .ZN(n4231) );
  NAND2_X1 U4886 ( .A1(n4229), .A2(n4228), .ZN(n4230) );
  OAI211_X1 U4887 ( .C1(n4232), .C2(n4255), .A(n4231), .B(n4230), .ZN(n4233)
         );
  INV_X1 U4888 ( .A(n4233), .ZN(n4234) );
  OAI211_X1 U4889 ( .C1(n4237), .C2(n4236), .A(n4235), .B(n4234), .ZN(n4611)
         );
  MUX2_X1 U4890 ( .A(n4611), .B(REG2_REG_2__SCAN_IN), .S(n4581), .Z(n4238) );
  INV_X1 U4891 ( .A(n4238), .ZN(n4243) );
  AOI22_X1 U4892 ( .A1(n4613), .A2(n4578), .B1(REG3_REG_2__SCAN_IN), .B2(n4577), .ZN(n4242) );
  NAND2_X1 U4893 ( .A1(n4240), .A2(n4239), .ZN(n4610) );
  NAND3_X1 U4894 ( .A1(n4563), .A2(n4609), .A3(n4610), .ZN(n4241) );
  NAND3_X1 U4895 ( .A1(n4243), .A2(n4242), .A3(n4241), .ZN(U3288) );
  INV_X1 U4896 ( .A(REG1_REG_31__SCAN_IN), .ZN(n4944) );
  NAND2_X1 U4897 ( .A1(n4249), .A2(n4256), .ZN(n4250) );
  XNOR2_X1 U4898 ( .A(n4250), .B(n4246), .ZN(n4412) );
  NAND2_X1 U4899 ( .A1(n4412), .A2(n4264), .ZN(n4248) );
  NAND2_X1 U4900 ( .A1(n4245), .A2(n4244), .ZN(n4254) );
  OAI21_X1 U4901 ( .B1(n4246), .B2(n4255), .A(n4254), .ZN(n4411) );
  NAND2_X1 U4902 ( .A1(n4658), .A2(n4411), .ZN(n4247) );
  OAI211_X1 U4903 ( .C1(n4658), .C2(n4944), .A(n4248), .B(n4247), .ZN(U3549)
         );
  INV_X1 U4904 ( .A(REG1_REG_30__SCAN_IN), .ZN(n4821) );
  INV_X1 U4905 ( .A(n4249), .ZN(n4252) );
  INV_X1 U4906 ( .A(n4250), .ZN(n4251) );
  NAND2_X1 U4907 ( .A1(n4415), .A2(n4264), .ZN(n4258) );
  OAI21_X1 U4908 ( .B1(n4256), .B2(n4255), .A(n4254), .ZN(n4414) );
  NAND2_X1 U4909 ( .A1(n4658), .A2(n4414), .ZN(n4257) );
  OAI211_X1 U4910 ( .C1(n4658), .C2(n4821), .A(n4258), .B(n4257), .ZN(U3548)
         );
  MUX2_X1 U4911 ( .A(REG1_REG_29__SCAN_IN), .B(n2260), .S(n4658), .Z(U3547) );
  AOI21_X1 U4912 ( .B1(n4263), .B2(n4642), .A(n4262), .ZN(n4328) );
  MUX2_X1 U4913 ( .A(n4819), .B(n4328), .S(n4658), .Z(n4266) );
  NAND2_X1 U4914 ( .A1(n4330), .A2(n4264), .ZN(n4265) );
  NAND2_X1 U4915 ( .A1(n4266), .A2(n4265), .ZN(U3546) );
  AOI21_X1 U4916 ( .B1(n4619), .B2(n4268), .A(n4267), .ZN(n4269) );
  OAI21_X1 U4917 ( .B1(n4270), .B2(n4605), .A(n4269), .ZN(n4333) );
  MUX2_X1 U4918 ( .A(REG1_REG_27__SCAN_IN), .B(n4333), .S(n4658), .Z(U3545) );
  INV_X1 U4919 ( .A(REG1_REG_25__SCAN_IN), .ZN(n4273) );
  AOI21_X1 U4920 ( .B1(n4272), .B2(n4642), .A(n4271), .ZN(n4334) );
  MUX2_X1 U4921 ( .A(n4273), .B(n4334), .S(n4658), .Z(n4274) );
  OAI21_X1 U4922 ( .B1(n4323), .B2(n4337), .A(n4274), .ZN(U3543) );
  AOI21_X1 U4923 ( .B1(n4276), .B2(n4642), .A(n4275), .ZN(n4338) );
  MUX2_X1 U4924 ( .A(n4941), .B(n4338), .S(n4658), .Z(n4277) );
  OAI21_X1 U4925 ( .B1(n4323), .B2(n4341), .A(n4277), .ZN(U3542) );
  AOI21_X1 U4926 ( .B1(n4279), .B2(n4642), .A(n4278), .ZN(n4342) );
  MUX2_X1 U4927 ( .A(n4942), .B(n4342), .S(n4658), .Z(n4280) );
  OAI21_X1 U4928 ( .B1(n4323), .B2(n4345), .A(n4280), .ZN(U3541) );
  NAND3_X1 U4929 ( .A1(n4282), .A2(n4619), .A3(n4281), .ZN(n4283) );
  OAI211_X1 U4930 ( .C1(n4285), .C2(n4605), .A(n4284), .B(n4283), .ZN(n4346)
         );
  MUX2_X1 U4931 ( .A(REG1_REG_22__SCAN_IN), .B(n4346), .S(n4658), .Z(U3540) );
  AOI21_X1 U4932 ( .B1(n4287), .B2(n4642), .A(n4286), .ZN(n4347) );
  MUX2_X1 U4933 ( .A(n4288), .B(n4347), .S(n4658), .Z(n4289) );
  OAI21_X1 U4934 ( .B1(n4323), .B2(n4350), .A(n4289), .ZN(U3539) );
  INV_X1 U4935 ( .A(n4290), .ZN(n4292) );
  AOI21_X1 U4936 ( .B1(n4623), .B2(n4292), .A(n4291), .ZN(n4351) );
  MUX2_X1 U4937 ( .A(n4935), .B(n4351), .S(n4658), .Z(n4293) );
  OAI21_X1 U4938 ( .B1(n4323), .B2(n4354), .A(n4293), .ZN(U3538) );
  AOI21_X1 U4939 ( .B1(n4295), .B2(n4642), .A(n4294), .ZN(n4355) );
  MUX2_X1 U4940 ( .A(n4296), .B(n4355), .S(n4658), .Z(n4297) );
  OAI21_X1 U4941 ( .B1(n4323), .B2(n4358), .A(n4297), .ZN(U3537) );
  INV_X1 U4942 ( .A(n4298), .ZN(n4301) );
  OAI211_X1 U4943 ( .C1(n4301), .C2(n4605), .A(n4300), .B(n4299), .ZN(n4359)
         );
  MUX2_X1 U4944 ( .A(REG1_REG_18__SCAN_IN), .B(n4359), .S(n4658), .Z(U3536) );
  AOI21_X1 U4945 ( .B1(n4303), .B2(n4642), .A(n4302), .ZN(n4360) );
  MUX2_X1 U4946 ( .A(n4304), .B(n4360), .S(n4658), .Z(n4305) );
  OAI21_X1 U4947 ( .B1(n4323), .B2(n4362), .A(n4305), .ZN(U3535) );
  NAND3_X1 U4948 ( .A1(n4307), .A2(n4619), .A3(n4306), .ZN(n4308) );
  OAI211_X1 U4949 ( .C1(n4310), .C2(n4605), .A(n4309), .B(n4308), .ZN(n4363)
         );
  MUX2_X1 U4950 ( .A(REG1_REG_16__SCAN_IN), .B(n4363), .S(n4658), .Z(U3534) );
  AOI21_X1 U4951 ( .B1(n4312), .B2(n4642), .A(n4311), .ZN(n4364) );
  MUX2_X1 U4952 ( .A(n4313), .B(n4364), .S(n4658), .Z(n4314) );
  OAI21_X1 U4953 ( .B1(n4323), .B2(n4366), .A(n4314), .ZN(U3533) );
  AOI21_X1 U4954 ( .B1(n4623), .B2(n4316), .A(n4315), .ZN(n4367) );
  MUX2_X1 U4955 ( .A(n4508), .B(n4367), .S(n4658), .Z(n4317) );
  OAI21_X1 U4956 ( .B1(n4323), .B2(n4370), .A(n4317), .ZN(U3532) );
  INV_X1 U4957 ( .A(n4318), .ZN(n4320) );
  AOI21_X1 U4958 ( .B1(n4623), .B2(n4320), .A(n4319), .ZN(n4371) );
  MUX2_X1 U4959 ( .A(n4321), .B(n4371), .S(n4658), .Z(n4322) );
  OAI21_X1 U4960 ( .B1(n4323), .B2(n4375), .A(n4322), .ZN(U3531) );
  NAND2_X1 U4961 ( .A1(n4412), .A2(n4329), .ZN(n4325) );
  NAND2_X1 U4962 ( .A1(n4645), .A2(n4411), .ZN(n4324) );
  OAI211_X1 U4963 ( .C1(n4645), .C2(n3185), .A(n4325), .B(n4324), .ZN(U3517)
         );
  NAND2_X1 U4964 ( .A1(n4415), .A2(n4329), .ZN(n4327) );
  NAND2_X1 U4965 ( .A1(n4645), .A2(n4414), .ZN(n4326) );
  OAI211_X1 U4966 ( .C1(n4645), .C2(n3226), .A(n4327), .B(n4326), .ZN(U3516)
         );
  MUX2_X1 U4967 ( .A(REG0_REG_29__SCAN_IN), .B(n2260), .S(n4645), .Z(U3515) );
  MUX2_X1 U4968 ( .A(n4945), .B(n4328), .S(n4645), .Z(n4332) );
  NAND2_X1 U4969 ( .A1(n4330), .A2(n4329), .ZN(n4331) );
  NAND2_X1 U4970 ( .A1(n4332), .A2(n4331), .ZN(U3514) );
  MUX2_X1 U4971 ( .A(REG0_REG_27__SCAN_IN), .B(n4333), .S(n4645), .Z(U3513) );
  INV_X1 U4972 ( .A(REG0_REG_25__SCAN_IN), .ZN(n4335) );
  MUX2_X1 U4973 ( .A(n4335), .B(n4334), .S(n4645), .Z(n4336) );
  OAI21_X1 U4974 ( .B1(n4337), .B2(n4374), .A(n4336), .ZN(U3511) );
  INV_X1 U4975 ( .A(REG0_REG_24__SCAN_IN), .ZN(n4339) );
  MUX2_X1 U4976 ( .A(n4339), .B(n4338), .S(n4645), .Z(n4340) );
  OAI21_X1 U4977 ( .B1(n4341), .B2(n4374), .A(n4340), .ZN(U3510) );
  MUX2_X1 U4978 ( .A(n4343), .B(n4342), .S(n4645), .Z(n4344) );
  OAI21_X1 U4979 ( .B1(n4345), .B2(n4374), .A(n4344), .ZN(U3509) );
  MUX2_X1 U4980 ( .A(REG0_REG_22__SCAN_IN), .B(n4346), .S(n4645), .Z(U3508) );
  MUX2_X1 U4981 ( .A(n4348), .B(n4347), .S(n4645), .Z(n4349) );
  OAI21_X1 U4982 ( .B1(n4350), .B2(n4374), .A(n4349), .ZN(U3507) );
  INV_X1 U4983 ( .A(REG0_REG_20__SCAN_IN), .ZN(n4352) );
  MUX2_X1 U4984 ( .A(n4352), .B(n4351), .S(n4645), .Z(n4353) );
  OAI21_X1 U4985 ( .B1(n4354), .B2(n4374), .A(n4353), .ZN(U3506) );
  INV_X1 U4986 ( .A(REG0_REG_19__SCAN_IN), .ZN(n4356) );
  MUX2_X1 U4987 ( .A(n4356), .B(n4355), .S(n4645), .Z(n4357) );
  OAI21_X1 U4988 ( .B1(n4358), .B2(n4374), .A(n4357), .ZN(U3505) );
  MUX2_X1 U4989 ( .A(REG0_REG_18__SCAN_IN), .B(n4359), .S(n4645), .Z(U3503) );
  MUX2_X1 U4990 ( .A(n4932), .B(n4360), .S(n4645), .Z(n4361) );
  OAI21_X1 U4991 ( .B1(n4362), .B2(n4374), .A(n4361), .ZN(U3501) );
  MUX2_X1 U4992 ( .A(REG0_REG_16__SCAN_IN), .B(n4363), .S(n4645), .Z(U3499) );
  MUX2_X1 U4993 ( .A(n4892), .B(n4364), .S(n4645), .Z(n4365) );
  OAI21_X1 U4994 ( .B1(n4366), .B2(n4374), .A(n4365), .ZN(U3497) );
  INV_X1 U4995 ( .A(REG0_REG_14__SCAN_IN), .ZN(n4368) );
  MUX2_X1 U4996 ( .A(n4368), .B(n4367), .S(n4645), .Z(n4369) );
  OAI21_X1 U4997 ( .B1(n4370), .B2(n4374), .A(n4369), .ZN(U3495) );
  MUX2_X1 U4998 ( .A(n4372), .B(n4371), .S(n4645), .Z(n4373) );
  OAI21_X1 U4999 ( .B1(n4375), .B2(n4374), .A(n4373), .ZN(U3493) );
  MUX2_X1 U5000 ( .A(DATAI_29_), .B(n4376), .S(STATE_REG_SCAN_IN), .Z(U3323)
         );
  MUX2_X1 U5001 ( .A(DATAI_28_), .B(n4377), .S(STATE_REG_SCAN_IN), .Z(U3324)
         );
  MUX2_X1 U5002 ( .A(DATAI_27_), .B(n4419), .S(STATE_REG_SCAN_IN), .Z(U3325)
         );
  MUX2_X1 U5003 ( .A(n4378), .B(DATAI_26_), .S(U3149), .Z(U3326) );
  MUX2_X1 U5004 ( .A(DATAI_22_), .B(n4379), .S(STATE_REG_SCAN_IN), .Z(U3330)
         );
  MUX2_X1 U5005 ( .A(n2542), .B(DATAI_20_), .S(U3149), .Z(U3332) );
  MUX2_X1 U5006 ( .A(n4380), .B(DATAI_19_), .S(U3149), .Z(U3333) );
  MUX2_X1 U5007 ( .A(DATAI_18_), .B(n4554), .S(STATE_REG_SCAN_IN), .Z(U3334)
         );
  MUX2_X1 U5008 ( .A(n4381), .B(DATAI_12_), .S(U3149), .Z(U3340) );
  MUX2_X1 U5009 ( .A(n4382), .B(DATAI_5_), .S(U3149), .Z(U3347) );
  MUX2_X1 U5010 ( .A(DATAI_4_), .B(n4432), .S(STATE_REG_SCAN_IN), .Z(U3348) );
  MUX2_X1 U5011 ( .A(n4383), .B(DATAI_3_), .S(U3149), .Z(U3349) );
  MUX2_X1 U5012 ( .A(n3144), .B(DATAI_2_), .S(U3149), .Z(U3350) );
  MUX2_X1 U5013 ( .A(n3143), .B(DATAI_1_), .S(U3149), .Z(U3351) );
  AOI21_X1 U5014 ( .B1(n5045), .B2(ADDR_REG_3__SCAN_IN), .A(n4384), .ZN(n4385)
         );
  OAI21_X1 U5015 ( .B1(n4547), .B2(n2419), .A(n4385), .ZN(n4386) );
  INV_X1 U5016 ( .A(n4386), .ZN(n4393) );
  OAI211_X1 U5017 ( .C1(REG1_REG_3__SCAN_IN), .C2(n4388), .A(n5038), .B(n4387), 
        .ZN(n4392) );
  OAI211_X1 U5018 ( .C1(REG2_REG_3__SCAN_IN), .C2(n4390), .A(n5042), .B(n4389), 
        .ZN(n4391) );
  NAND3_X1 U5019 ( .A1(n4393), .A2(n4392), .A3(n4391), .ZN(U3243) );
  OAI22_X1 U5020 ( .A1(n3733), .A2(n4395), .B1(n4394), .B2(n3722), .ZN(n4400)
         );
  NOR2_X1 U5021 ( .A1(STATE_REG_SCAN_IN), .A2(n4396), .ZN(n4526) );
  INV_X1 U5022 ( .A(n4526), .ZN(n4397) );
  OAI21_X1 U5023 ( .B1(n3720), .B2(n4398), .A(n4397), .ZN(n4399) );
  NOR2_X1 U5024 ( .A1(n4400), .A2(n4399), .ZN(n4408) );
  INV_X1 U5025 ( .A(n3728), .ZN(n4402) );
  OAI21_X1 U5026 ( .B1(n4402), .B2(n4401), .A(n3727), .ZN(n4404) );
  XNOR2_X1 U5027 ( .A(n4404), .B(n4403), .ZN(n4406) );
  NAND2_X1 U5028 ( .A1(n4406), .A2(n4405), .ZN(n4407) );
  OAI211_X1 U5029 ( .C1(n4410), .C2(n4409), .A(n4408), .B(n4407), .ZN(U3223)
         );
  AOI22_X1 U5030 ( .A1(n4412), .A2(n4563), .B1(n3576), .B2(n4411), .ZN(n4413)
         );
  OAI21_X1 U5031 ( .B1(n3576), .B2(n3188), .A(n4413), .ZN(U3260) );
  AOI22_X1 U5032 ( .A1(n4415), .A2(n4563), .B1(n3576), .B2(n4414), .ZN(n4416)
         );
  OAI21_X1 U5033 ( .B1(n3229), .B2(n3576), .A(n4416), .ZN(U3261) );
  INV_X1 U5034 ( .A(n4417), .ZN(n4418) );
  OAI21_X1 U5035 ( .B1(REG1_REG_0__SCAN_IN), .B2(n4419), .A(n4418), .ZN(n4420)
         );
  XNOR2_X1 U5036 ( .A(n4420), .B(n5035), .ZN(n4423) );
  AOI22_X1 U5037 ( .A1(ADDR_REG_0__SCAN_IN), .A2(n5045), .B1(
        REG3_REG_0__SCAN_IN), .B2(U3149), .ZN(n4421) );
  OAI21_X1 U5038 ( .B1(n4423), .B2(n4422), .A(n4421), .ZN(U3240) );
  AOI21_X1 U5039 ( .B1(n5045), .B2(ADDR_REG_4__SCAN_IN), .A(n4424), .ZN(n4425)
         );
  INV_X1 U5040 ( .A(n4425), .ZN(n4431) );
  XNOR2_X1 U5041 ( .A(n4426), .B(REG1_REG_4__SCAN_IN), .ZN(n4429) );
  XOR2_X1 U5042 ( .A(REG2_REG_4__SCAN_IN), .B(n4427), .Z(n4428) );
  OAI22_X1 U5043 ( .A1(n4429), .A2(n4548), .B1(n4551), .B2(n4428), .ZN(n4430)
         );
  AOI211_X1 U5044 ( .C1(n4432), .C2(n5046), .A(n4431), .B(n4430), .ZN(n4434)
         );
  NAND2_X1 U5045 ( .A1(n4434), .A2(n4433), .ZN(U3244) );
  AOI21_X1 U5046 ( .B1(n5045), .B2(ADDR_REG_6__SCAN_IN), .A(n4435), .ZN(n4444)
         );
  OAI211_X1 U5047 ( .C1(REG1_REG_6__SCAN_IN), .C2(n4437), .A(n5038), .B(n4436), 
        .ZN(n4443) );
  OAI211_X1 U5048 ( .C1(REG2_REG_6__SCAN_IN), .C2(n4439), .A(n5042), .B(n4438), 
        .ZN(n4442) );
  NAND2_X1 U5049 ( .A1(n4440), .A2(n5046), .ZN(n4441) );
  NAND4_X1 U5050 ( .A1(n4444), .A2(n4443), .A3(n4442), .A4(n4441), .ZN(U3246)
         );
  AOI22_X1 U5051 ( .A1(REG1_REG_7__SCAN_IN), .A2(n4445), .B1(n4597), .B2(n2650), .ZN(n4448) );
  OAI21_X1 U5052 ( .B1(n4448), .B2(n4447), .A(n5038), .ZN(n4446) );
  AOI21_X1 U5053 ( .B1(n4448), .B2(n4447), .A(n4446), .ZN(n4450) );
  AOI211_X1 U5054 ( .C1(n5045), .C2(ADDR_REG_7__SCAN_IN), .A(n4450), .B(n4449), 
        .ZN(n4455) );
  OAI211_X1 U5055 ( .C1(n4453), .C2(n4452), .A(n5042), .B(n4451), .ZN(n4454)
         );
  OAI211_X1 U5056 ( .C1(n4547), .C2(n4597), .A(n4455), .B(n4454), .ZN(U3247)
         );
  AOI211_X1 U5057 ( .C1(n2669), .C2(n4457), .A(n4456), .B(n4548), .ZN(n4459)
         );
  AOI211_X1 U5058 ( .C1(n5045), .C2(ADDR_REG_8__SCAN_IN), .A(n4459), .B(n4458), 
        .ZN(n4463) );
  OAI211_X1 U5059 ( .C1(REG2_REG_8__SCAN_IN), .C2(n4461), .A(n5042), .B(n4460), 
        .ZN(n4462) );
  OAI211_X1 U5060 ( .C1(n4547), .C2(n3499), .A(n4463), .B(n4462), .ZN(U3248)
         );
  AOI211_X1 U5061 ( .C1(n4466), .C2(n4465), .A(n4464), .B(n4548), .ZN(n4468)
         );
  AOI211_X1 U5062 ( .C1(n5045), .C2(ADDR_REG_9__SCAN_IN), .A(n4468), .B(n4467), 
        .ZN(n4473) );
  OAI211_X1 U5063 ( .C1(n4471), .C2(n4470), .A(n5042), .B(n4469), .ZN(n4472)
         );
  OAI211_X1 U5064 ( .C1(n4547), .C2(n4596), .A(n4473), .B(n4472), .ZN(U3249)
         );
  AOI211_X1 U5065 ( .C1(n4476), .C2(n4475), .A(n4474), .B(n4548), .ZN(n4478)
         );
  AOI211_X1 U5066 ( .C1(n5045), .C2(ADDR_REG_10__SCAN_IN), .A(n4478), .B(n4477), .ZN(n4482) );
  OAI211_X1 U5067 ( .C1(REG2_REG_10__SCAN_IN), .C2(n4480), .A(n5042), .B(n4479), .ZN(n4481) );
  OAI211_X1 U5068 ( .C1(n4547), .C2(n2411), .A(n4482), .B(n4481), .ZN(U3250)
         );
  AOI211_X1 U5069 ( .C1(n4485), .C2(n4484), .A(n4483), .B(n4548), .ZN(n4487)
         );
  AOI211_X1 U5070 ( .C1(n5045), .C2(ADDR_REG_11__SCAN_IN), .A(n4487), .B(n4486), .ZN(n4492) );
  OAI211_X1 U5071 ( .C1(n4490), .C2(n4489), .A(n5042), .B(n4488), .ZN(n4491)
         );
  OAI211_X1 U5072 ( .C1(n4547), .C2(n4493), .A(n4492), .B(n4491), .ZN(U3251)
         );
  AOI211_X1 U5073 ( .C1(n4496), .C2(n4495), .A(n4494), .B(n4548), .ZN(n4497)
         );
  AOI211_X1 U5074 ( .C1(n5045), .C2(ADDR_REG_13__SCAN_IN), .A(n4498), .B(n4497), .ZN(n4504) );
  AOI22_X1 U5075 ( .A1(REG2_REG_13__SCAN_IN), .A2(n4499), .B1(n4590), .B2(
        n3547), .ZN(n4502) );
  AOI21_X1 U5076 ( .B1(n4502), .B2(n4501), .A(n4551), .ZN(n4500) );
  OAI21_X1 U5077 ( .B1(n4502), .B2(n4501), .A(n4500), .ZN(n4503) );
  OAI211_X1 U5078 ( .C1(n4547), .C2(n4590), .A(n4504), .B(n4503), .ZN(U3253)
         );
  NAND2_X1 U5079 ( .A1(ADDR_REG_14__SCAN_IN), .A2(n5045), .ZN(n4515) );
  AOI211_X1 U5080 ( .C1(n4215), .C2(n4506), .A(n4505), .B(n4551), .ZN(n4511)
         );
  AOI211_X1 U5081 ( .C1(n4509), .C2(n4508), .A(n4507), .B(n4548), .ZN(n4510)
         );
  AOI211_X1 U5082 ( .C1(n5046), .C2(n4512), .A(n4511), .B(n4510), .ZN(n4514)
         );
  NAND3_X1 U5083 ( .A1(n4515), .A2(n4514), .A3(n4513), .ZN(U3254) );
  AOI211_X1 U5084 ( .C1(n4518), .C2(n4517), .A(n4516), .B(n4551), .ZN(n4519)
         );
  AOI211_X1 U5085 ( .C1(n5045), .C2(ADDR_REG_15__SCAN_IN), .A(n4520), .B(n4519), .ZN(n4525) );
  AOI21_X1 U5086 ( .B1(n4522), .B2(n2238), .A(n4521), .ZN(n4523) );
  NAND2_X1 U5087 ( .A1(n5038), .A2(n4523), .ZN(n4524) );
  OAI211_X1 U5088 ( .C1(n4547), .C2(n4589), .A(n4525), .B(n4524), .ZN(U3255)
         );
  AOI21_X1 U5089 ( .B1(n5045), .B2(ADDR_REG_16__SCAN_IN), .A(n4526), .ZN(n4535) );
  OAI21_X1 U5090 ( .B1(n4529), .B2(n4528), .A(n4527), .ZN(n4533) );
  OAI21_X1 U5091 ( .B1(n4531), .B2(n4193), .A(n4530), .ZN(n4532) );
  AOI22_X1 U5092 ( .A1(n5038), .A2(n4533), .B1(n5042), .B2(n4532), .ZN(n4534)
         );
  OAI211_X1 U5093 ( .C1(n4587), .C2(n4547), .A(n4535), .B(n4534), .ZN(U3256)
         );
  AOI21_X1 U5094 ( .B1(n5045), .B2(ADDR_REG_17__SCAN_IN), .A(n4536), .ZN(n4546) );
  OAI21_X1 U5095 ( .B1(n4539), .B2(n4538), .A(n4537), .ZN(n4544) );
  OAI21_X1 U5096 ( .B1(n4542), .B2(n4541), .A(n4540), .ZN(n4543) );
  AOI22_X1 U5097 ( .A1(n5038), .A2(n4544), .B1(n5042), .B2(n4543), .ZN(n4545)
         );
  OAI211_X1 U5098 ( .C1(n4586), .C2(n4547), .A(n4546), .B(n4545), .ZN(U3257)
         );
  INV_X1 U5099 ( .A(ADDR_REG_18__SCAN_IN), .ZN(n4950) );
  AOI21_X1 U5100 ( .B1(n4550), .B2(n4549), .A(n4548), .ZN(n4557) );
  INV_X1 U5101 ( .A(n4554), .ZN(n4555) );
  AOI22_X1 U5102 ( .A1(n4561), .A2(n4577), .B1(REG2_REG_6__SCAN_IN), .B2(n4581), .ZN(n4566) );
  AOI22_X1 U5103 ( .A1(n4564), .A2(n4578), .B1(n4563), .B2(n4562), .ZN(n4565)
         );
  OAI211_X1 U5104 ( .C1(n4581), .C2(n4567), .A(n4566), .B(n4565), .ZN(U3284)
         );
  NOR2_X1 U5105 ( .A1(n4569), .A2(n4568), .ZN(n4601) );
  INV_X1 U5106 ( .A(n4570), .ZN(n4602) );
  OAI21_X1 U5107 ( .B1(n4572), .B2(n4571), .A(n4602), .ZN(n4573) );
  OAI21_X1 U5108 ( .B1(n4575), .B2(n4574), .A(n4573), .ZN(n4600) );
  AOI21_X1 U5109 ( .B1(n4601), .B2(n4576), .A(n4600), .ZN(n4580) );
  AOI22_X1 U5110 ( .A1(n4578), .A2(n4602), .B1(REG3_REG_0__SCAN_IN), .B2(n4577), .ZN(n4579) );
  OAI221_X1 U5111 ( .B1(n4581), .B2(n4580), .C1(n3576), .C2(n4977), .A(n4579), 
        .ZN(U3290) );
  AND2_X1 U5112 ( .A1(D_REG_31__SCAN_IN), .A2(n4583), .ZN(U3291) );
  AND2_X1 U5113 ( .A1(D_REG_30__SCAN_IN), .A2(n4583), .ZN(U3292) );
  INV_X1 U5114 ( .A(D_REG_29__SCAN_IN), .ZN(n4800) );
  NOR2_X1 U5115 ( .A1(n4582), .A2(n4800), .ZN(U3293) );
  AND2_X1 U5116 ( .A1(D_REG_28__SCAN_IN), .A2(n4583), .ZN(U3294) );
  AND2_X1 U5117 ( .A1(D_REG_27__SCAN_IN), .A2(n4583), .ZN(U3295) );
  INV_X1 U5118 ( .A(D_REG_26__SCAN_IN), .ZN(n4926) );
  NOR2_X1 U5119 ( .A1(n4582), .A2(n4926), .ZN(U3296) );
  INV_X1 U5120 ( .A(D_REG_25__SCAN_IN), .ZN(n4930) );
  NOR2_X1 U5121 ( .A1(n4582), .A2(n4930), .ZN(U3297) );
  INV_X1 U5122 ( .A(D_REG_24__SCAN_IN), .ZN(n4801) );
  NOR2_X1 U5123 ( .A1(n4582), .A2(n4801), .ZN(U3298) );
  AND2_X1 U5124 ( .A1(D_REG_23__SCAN_IN), .A2(n4583), .ZN(U3299) );
  AND2_X1 U5125 ( .A1(D_REG_22__SCAN_IN), .A2(n4583), .ZN(U3300) );
  INV_X1 U5126 ( .A(D_REG_21__SCAN_IN), .ZN(n4929) );
  NOR2_X1 U5127 ( .A1(n4582), .A2(n4929), .ZN(U3301) );
  AND2_X1 U5128 ( .A1(D_REG_20__SCAN_IN), .A2(n4583), .ZN(U3302) );
  INV_X1 U5129 ( .A(D_REG_19__SCAN_IN), .ZN(n4909) );
  NOR2_X1 U5130 ( .A1(n4582), .A2(n4909), .ZN(U3303) );
  INV_X1 U5131 ( .A(D_REG_18__SCAN_IN), .ZN(n4913) );
  NOR2_X1 U5132 ( .A1(n4582), .A2(n4913), .ZN(U3304) );
  INV_X1 U5133 ( .A(D_REG_17__SCAN_IN), .ZN(n4912) );
  NOR2_X1 U5134 ( .A1(n4582), .A2(n4912), .ZN(U3305) );
  AND2_X1 U5135 ( .A1(D_REG_16__SCAN_IN), .A2(n4583), .ZN(U3306) );
  AND2_X1 U5136 ( .A1(D_REG_15__SCAN_IN), .A2(n4583), .ZN(U3307) );
  AND2_X1 U5137 ( .A1(D_REG_14__SCAN_IN), .A2(n4583), .ZN(U3308) );
  AND2_X1 U5138 ( .A1(n4583), .A2(D_REG_13__SCAN_IN), .ZN(U3309) );
  INV_X1 U5139 ( .A(D_REG_12__SCAN_IN), .ZN(n4791) );
  NOR2_X1 U5140 ( .A1(n4582), .A2(n4791), .ZN(U3310) );
  AND2_X1 U5141 ( .A1(n4583), .A2(D_REG_11__SCAN_IN), .ZN(U3311) );
  INV_X1 U5142 ( .A(D_REG_10__SCAN_IN), .ZN(n4792) );
  NOR2_X1 U5143 ( .A1(n4582), .A2(n4792), .ZN(U3312) );
  INV_X1 U5144 ( .A(D_REG_9__SCAN_IN), .ZN(n4906) );
  NOR2_X1 U5145 ( .A1(n4582), .A2(n4906), .ZN(U3313) );
  INV_X1 U5146 ( .A(D_REG_8__SCAN_IN), .ZN(n4927) );
  NOR2_X1 U5147 ( .A1(n4582), .A2(n4927), .ZN(U3314) );
  INV_X1 U5148 ( .A(D_REG_7__SCAN_IN), .ZN(n4907) );
  NOR2_X1 U5149 ( .A1(n4582), .A2(n4907), .ZN(U3315) );
  AND2_X1 U5150 ( .A1(D_REG_6__SCAN_IN), .A2(n4583), .ZN(U3316) );
  INV_X1 U5151 ( .A(D_REG_5__SCAN_IN), .ZN(n4910) );
  NOR2_X1 U5152 ( .A1(n4582), .A2(n4910), .ZN(U3317) );
  AND2_X1 U5153 ( .A1(n4583), .A2(D_REG_4__SCAN_IN), .ZN(U3318) );
  AND2_X1 U5154 ( .A1(D_REG_3__SCAN_IN), .A2(n4583), .ZN(U3319) );
  AND2_X1 U5155 ( .A1(D_REG_2__SCAN_IN), .A2(n4583), .ZN(U3320) );
  OAI21_X1 U5156 ( .B1(STATE_REG_SCAN_IN), .B2(DATAI_23_), .A(n4584), .ZN(
        n4585) );
  INV_X1 U5157 ( .A(n4585), .ZN(U3329) );
  INV_X1 U5158 ( .A(DATAI_17_), .ZN(n4883) );
  AOI22_X1 U5159 ( .A1(STATE_REG_SCAN_IN), .A2(n4586), .B1(n4883), .B2(U3149), 
        .ZN(U3335) );
  INV_X1 U5160 ( .A(DATAI_16_), .ZN(n4774) );
  AOI22_X1 U5161 ( .A1(STATE_REG_SCAN_IN), .A2(n4587), .B1(n4774), .B2(U3149), 
        .ZN(U3336) );
  INV_X1 U5162 ( .A(DATAI_15_), .ZN(n4588) );
  AOI22_X1 U5163 ( .A1(STATE_REG_SCAN_IN), .A2(n4589), .B1(n4588), .B2(U3149), 
        .ZN(U3337) );
  INV_X1 U5164 ( .A(DATAI_13_), .ZN(n4957) );
  AOI22_X1 U5165 ( .A1(STATE_REG_SCAN_IN), .A2(n4590), .B1(n4957), .B2(U3149), 
        .ZN(U3339) );
  OAI22_X1 U5166 ( .A1(U3149), .A2(n4591), .B1(DATAI_11_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4592) );
  INV_X1 U5167 ( .A(n4592), .ZN(U3341) );
  OAI22_X1 U5168 ( .A1(U3149), .A2(n4593), .B1(DATAI_10_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4594) );
  INV_X1 U5169 ( .A(n4594), .ZN(U3342) );
  INV_X1 U5170 ( .A(DATAI_9_), .ZN(n4595) );
  AOI22_X1 U5171 ( .A1(STATE_REG_SCAN_IN), .A2(n4596), .B1(n4595), .B2(U3149), 
        .ZN(U3343) );
  INV_X1 U5172 ( .A(DATAI_8_), .ZN(n4899) );
  AOI22_X1 U5173 ( .A1(STATE_REG_SCAN_IN), .A2(n3499), .B1(n4899), .B2(U3149), 
        .ZN(U3344) );
  INV_X1 U5174 ( .A(DATAI_7_), .ZN(n4773) );
  AOI22_X1 U5175 ( .A1(STATE_REG_SCAN_IN), .A2(n4597), .B1(n4773), .B2(U3149), 
        .ZN(U3345) );
  INV_X1 U5176 ( .A(DATAI_6_), .ZN(n4900) );
  AOI22_X1 U5177 ( .A1(STATE_REG_SCAN_IN), .A2(n4598), .B1(n4900), .B2(U3149), 
        .ZN(U3346) );
  OAI22_X1 U5178 ( .A1(U3149), .A2(IR_REG_0__SCAN_IN), .B1(DATAI_0_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4599) );
  INV_X1 U5179 ( .A(n4599), .ZN(U3352) );
  AOI211_X1 U5180 ( .C1(n4623), .C2(n4602), .A(n4601), .B(n4600), .ZN(n4646)
         );
  AOI22_X1 U5181 ( .A1(n4645), .A2(n4646), .B1(n2537), .B2(n4644), .ZN(U3467)
         );
  INV_X1 U5182 ( .A(n4603), .ZN(n4608) );
  OAI22_X1 U5183 ( .A1(n4606), .A2(n4605), .B1(n4638), .B2(n4604), .ZN(n4607)
         );
  NOR2_X1 U5184 ( .A1(n4608), .A2(n4607), .ZN(n4648) );
  AOI22_X1 U5185 ( .A1(n4645), .A2(n4648), .B1(n2549), .B2(n4644), .ZN(U3469)
         );
  AND3_X1 U5186 ( .A1(n4610), .A2(n4619), .A3(n4609), .ZN(n4612) );
  AOI211_X1 U5187 ( .C1(n4623), .C2(n4613), .A(n4612), .B(n4611), .ZN(n4649)
         );
  AOI22_X1 U5188 ( .A1(n4645), .A2(n4649), .B1(n2565), .B2(n4644), .ZN(U3471)
         );
  NOR2_X1 U5189 ( .A1(n4615), .A2(n4614), .ZN(n4617) );
  AOI211_X1 U5190 ( .C1(n4619), .C2(n4618), .A(n4617), .B(n4616), .ZN(n4651)
         );
  AOI22_X1 U5191 ( .A1(n4645), .A2(n4651), .B1(n2583), .B2(n4644), .ZN(U3473)
         );
  INV_X1 U5192 ( .A(n4620), .ZN(n4622) );
  AOI211_X1 U5193 ( .C1(n4624), .C2(n4623), .A(n4622), .B(n4621), .ZN(n4652)
         );
  INV_X1 U5194 ( .A(REG0_REG_4__SCAN_IN), .ZN(n4625) );
  AOI22_X1 U5195 ( .A1(n4645), .A2(n4652), .B1(n4625), .B2(n4644), .ZN(U3475)
         );
  OAI21_X1 U5196 ( .B1(n4638), .B2(n4627), .A(n4626), .ZN(n4628) );
  AOI21_X1 U5197 ( .B1(n4629), .B2(n4642), .A(n4628), .ZN(n4653) );
  INV_X1 U5198 ( .A(REG0_REG_5__SCAN_IN), .ZN(n4630) );
  AOI22_X1 U5199 ( .A1(n4645), .A2(n4653), .B1(n4630), .B2(n4644), .ZN(U3477)
         );
  AOI211_X1 U5200 ( .C1(n4633), .C2(n4642), .A(n4632), .B(n4631), .ZN(n4654)
         );
  INV_X1 U5201 ( .A(REG0_REG_7__SCAN_IN), .ZN(n4804) );
  AOI22_X1 U5202 ( .A1(n4645), .A2(n4654), .B1(n4804), .B2(n4644), .ZN(U3481)
         );
  OAI21_X1 U5203 ( .B1(n4638), .B2(n4635), .A(n4634), .ZN(n4636) );
  AOI21_X1 U5204 ( .B1(n4637), .B2(n4642), .A(n4636), .ZN(n4655) );
  AOI22_X1 U5205 ( .A1(n4645), .A2(n4655), .B1(n2686), .B2(n4644), .ZN(U3485)
         );
  NOR2_X1 U5206 ( .A1(n4639), .A2(n4638), .ZN(n4641) );
  AOI211_X1 U5207 ( .C1(n4643), .C2(n4642), .A(n4641), .B(n4640), .ZN(n4657)
         );
  AOI22_X1 U5208 ( .A1(n4645), .A2(n4657), .B1(n2720), .B2(n4644), .ZN(U3489)
         );
  AOI22_X1 U5209 ( .A1(n4658), .A2(n4646), .B1(n5034), .B2(n4656), .ZN(U3518)
         );
  AOI22_X1 U5210 ( .A1(n4658), .A2(n4648), .B1(n4647), .B2(n4656), .ZN(U3519)
         );
  AOI22_X1 U5211 ( .A1(n4658), .A2(n4649), .B1(n4879), .B2(n4656), .ZN(U3520)
         );
  INV_X1 U5212 ( .A(REG1_REG_3__SCAN_IN), .ZN(n4650) );
  AOI22_X1 U5213 ( .A1(n4658), .A2(n4651), .B1(n4650), .B2(n4656), .ZN(U3521)
         );
  AOI22_X1 U5214 ( .A1(n4658), .A2(n4652), .B1(n2403), .B2(n4656), .ZN(U3522)
         );
  AOI22_X1 U5215 ( .A1(n4658), .A2(n4653), .B1(n3142), .B2(n4656), .ZN(U3523)
         );
  AOI22_X1 U5216 ( .A1(n4658), .A2(n4654), .B1(n2650), .B2(n4656), .ZN(U3525)
         );
  AOI22_X1 U5217 ( .A1(n4658), .A2(n4655), .B1(n2685), .B2(n4656), .ZN(U3527)
         );
  AOI22_X1 U5218 ( .A1(n4658), .A2(n4657), .B1(n4880), .B2(n4656), .ZN(U3529)
         );
  OAI22_X1 U5219 ( .A1(REG2_REG_21__SCAN_IN), .A2(keyinput26), .B1(
        REG2_REG_20__SCAN_IN), .B2(keyinput89), .ZN(n4659) );
  AOI221_X1 U5220 ( .B1(REG2_REG_21__SCAN_IN), .B2(keyinput26), .C1(keyinput89), .C2(REG2_REG_20__SCAN_IN), .A(n4659), .ZN(n4666) );
  OAI22_X1 U5221 ( .A1(REG3_REG_26__SCAN_IN), .A2(keyinput112), .B1(
        keyinput104), .B2(DATAO_REG_14__SCAN_IN), .ZN(n4660) );
  AOI221_X1 U5222 ( .B1(REG3_REG_26__SCAN_IN), .B2(keyinput112), .C1(
        DATAO_REG_14__SCAN_IN), .C2(keyinput104), .A(n4660), .ZN(n4665) );
  OAI22_X1 U5223 ( .A1(REG0_REG_27__SCAN_IN), .A2(keyinput33), .B1(DATAI_24_), 
        .B2(keyinput58), .ZN(n4661) );
  AOI221_X1 U5224 ( .B1(REG0_REG_27__SCAN_IN), .B2(keyinput33), .C1(keyinput58), .C2(DATAI_24_), .A(n4661), .ZN(n4664) );
  OAI22_X1 U5225 ( .A1(REG2_REG_16__SCAN_IN), .A2(keyinput21), .B1(
        REG0_REG_31__SCAN_IN), .B2(keyinput102), .ZN(n4662) );
  AOI221_X1 U5226 ( .B1(REG2_REG_16__SCAN_IN), .B2(keyinput21), .C1(
        keyinput102), .C2(REG0_REG_31__SCAN_IN), .A(n4662), .ZN(n4663) );
  NAND4_X1 U5227 ( .A1(n4666), .A2(n4665), .A3(n4664), .A4(n4663), .ZN(n4694)
         );
  OAI22_X1 U5228 ( .A1(REG2_REG_25__SCAN_IN), .A2(keyinput115), .B1(
        REG2_REG_17__SCAN_IN), .B2(keyinput117), .ZN(n4667) );
  AOI221_X1 U5229 ( .B1(REG2_REG_25__SCAN_IN), .B2(keyinput115), .C1(
        keyinput117), .C2(REG2_REG_17__SCAN_IN), .A(n4667), .ZN(n4674) );
  OAI22_X1 U5230 ( .A1(REG3_REG_25__SCAN_IN), .A2(keyinput103), .B1(DATAI_1_), 
        .B2(keyinput70), .ZN(n4668) );
  AOI221_X1 U5231 ( .B1(REG3_REG_25__SCAN_IN), .B2(keyinput103), .C1(
        keyinput70), .C2(DATAI_1_), .A(n4668), .ZN(n4673) );
  OAI22_X1 U5232 ( .A1(DATAO_REG_9__SCAN_IN), .A2(keyinput20), .B1(
        DATAO_REG_15__SCAN_IN), .B2(keyinput10), .ZN(n4669) );
  AOI221_X1 U5233 ( .B1(DATAO_REG_9__SCAN_IN), .B2(keyinput20), .C1(keyinput10), .C2(DATAO_REG_15__SCAN_IN), .A(n4669), .ZN(n4672) );
  OAI22_X1 U5234 ( .A1(REG2_REG_3__SCAN_IN), .A2(keyinput93), .B1(keyinput78), 
        .B2(DATAI_2_), .ZN(n4670) );
  AOI221_X1 U5235 ( .B1(REG2_REG_3__SCAN_IN), .B2(keyinput93), .C1(DATAI_2_), 
        .C2(keyinput78), .A(n4670), .ZN(n4671) );
  NAND4_X1 U5236 ( .A1(n4674), .A2(n4673), .A3(n4672), .A4(n4671), .ZN(n4693)
         );
  OAI22_X1 U5237 ( .A1(IR_REG_31__SCAN_IN), .A2(keyinput121), .B1(keyinput46), 
        .B2(D_REG_4__SCAN_IN), .ZN(n4675) );
  AOI221_X1 U5238 ( .B1(IR_REG_31__SCAN_IN), .B2(keyinput121), .C1(
        D_REG_4__SCAN_IN), .C2(keyinput46), .A(n4675), .ZN(n4682) );
  OAI22_X1 U5239 ( .A1(D_REG_13__SCAN_IN), .A2(keyinput42), .B1(
        D_REG_11__SCAN_IN), .B2(keyinput85), .ZN(n4676) );
  AOI221_X1 U5240 ( .B1(D_REG_13__SCAN_IN), .B2(keyinput42), .C1(keyinput85), 
        .C2(D_REG_11__SCAN_IN), .A(n4676), .ZN(n4681) );
  OAI22_X1 U5241 ( .A1(REG0_REG_3__SCAN_IN), .A2(keyinput116), .B1(keyinput23), 
        .B2(DATAI_0_), .ZN(n4677) );
  AOI221_X1 U5242 ( .B1(REG0_REG_3__SCAN_IN), .B2(keyinput116), .C1(DATAI_0_), 
        .C2(keyinput23), .A(n4677), .ZN(n4680) );
  OAI22_X1 U5243 ( .A1(IR_REG_14__SCAN_IN), .A2(keyinput28), .B1(DATAI_10_), 
        .B2(keyinput90), .ZN(n4678) );
  AOI221_X1 U5244 ( .B1(IR_REG_14__SCAN_IN), .B2(keyinput28), .C1(keyinput90), 
        .C2(DATAI_10_), .A(n4678), .ZN(n4679) );
  NAND4_X1 U5245 ( .A1(n4682), .A2(n4681), .A3(n4680), .A4(n4679), .ZN(n4692)
         );
  OAI22_X1 U5246 ( .A1(REG1_REG_6__SCAN_IN), .A2(keyinput82), .B1(keyinput86), 
        .B2(ADDR_REG_0__SCAN_IN), .ZN(n4683) );
  AOI221_X1 U5247 ( .B1(REG1_REG_6__SCAN_IN), .B2(keyinput82), .C1(
        ADDR_REG_0__SCAN_IN), .C2(keyinput86), .A(n4683), .ZN(n4690) );
  OAI22_X1 U5248 ( .A1(REG0_REG_23__SCAN_IN), .A2(keyinput11), .B1(DATAI_23_), 
        .B2(keyinput113), .ZN(n4684) );
  AOI221_X1 U5249 ( .B1(REG0_REG_23__SCAN_IN), .B2(keyinput11), .C1(
        keyinput113), .C2(DATAI_23_), .A(n4684), .ZN(n4689) );
  OAI22_X1 U5250 ( .A1(REG1_REG_16__SCAN_IN), .A2(keyinput88), .B1(
        REG1_REG_5__SCAN_IN), .B2(keyinput1), .ZN(n4685) );
  AOI221_X1 U5251 ( .B1(REG1_REG_16__SCAN_IN), .B2(keyinput88), .C1(keyinput1), 
        .C2(REG1_REG_5__SCAN_IN), .A(n4685), .ZN(n4688) );
  OAI22_X1 U5252 ( .A1(REG2_REG_10__SCAN_IN), .A2(keyinput66), .B1(
        REG2_REG_2__SCAN_IN), .B2(keyinput107), .ZN(n4686) );
  AOI221_X1 U5253 ( .B1(REG2_REG_10__SCAN_IN), .B2(keyinput66), .C1(
        keyinput107), .C2(REG2_REG_2__SCAN_IN), .A(n4686), .ZN(n4687) );
  NAND4_X1 U5254 ( .A1(n4690), .A2(n4689), .A3(n4688), .A4(n4687), .ZN(n4691)
         );
  NOR4_X1 U5255 ( .A1(n4694), .A2(n4693), .A3(n4692), .A4(n4691), .ZN(n5033)
         );
  AOI22_X1 U5256 ( .A1(DATAI_23_), .A2(keyinput241), .B1(DATAI_28_), .B2(
        keyinput219), .ZN(n4695) );
  OAI221_X1 U5257 ( .B1(DATAI_23_), .B2(keyinput241), .C1(DATAI_28_), .C2(
        keyinput219), .A(n4695), .ZN(n4702) );
  AOI22_X1 U5258 ( .A1(DATAI_20_), .A2(keyinput132), .B1(DATAI_21_), .B2(
        keyinput199), .ZN(n4696) );
  OAI221_X1 U5259 ( .B1(DATAI_20_), .B2(keyinput132), .C1(DATAI_21_), .C2(
        keyinput199), .A(n4696), .ZN(n4701) );
  AOI22_X1 U5260 ( .A1(DATAI_17_), .A2(keyinput143), .B1(DATAI_19_), .B2(
        keyinput238), .ZN(n4697) );
  OAI221_X1 U5261 ( .B1(DATAI_17_), .B2(keyinput143), .C1(DATAI_19_), .C2(
        keyinput238), .A(n4697), .ZN(n4700) );
  AOI22_X1 U5262 ( .A1(DATAI_14_), .A2(keyinput181), .B1(DATAI_10_), .B2(
        keyinput218), .ZN(n4698) );
  OAI221_X1 U5263 ( .B1(DATAI_14_), .B2(keyinput181), .C1(DATAI_10_), .C2(
        keyinput218), .A(n4698), .ZN(n4699) );
  NOR4_X1 U5264 ( .A1(n4702), .A2(n4701), .A3(n4700), .A4(n4699), .ZN(n4730)
         );
  AOI22_X1 U5265 ( .A1(DATAI_13_), .A2(keyinput160), .B1(DATAI_4_), .B2(
        keyinput171), .ZN(n4703) );
  OAI221_X1 U5266 ( .B1(DATAI_13_), .B2(keyinput160), .C1(DATAI_4_), .C2(
        keyinput171), .A(n4703), .ZN(n4710) );
  AOI22_X1 U5267 ( .A1(DATAI_2_), .A2(keyinput206), .B1(DATAI_3_), .B2(
        keyinput140), .ZN(n4704) );
  OAI221_X1 U5268 ( .B1(DATAI_2_), .B2(keyinput206), .C1(DATAI_3_), .C2(
        keyinput140), .A(n4704), .ZN(n4709) );
  AOI22_X1 U5269 ( .A1(DATAI_0_), .A2(keyinput151), .B1(DATAI_1_), .B2(
        keyinput198), .ZN(n4705) );
  OAI221_X1 U5270 ( .B1(DATAI_0_), .B2(keyinput151), .C1(DATAI_1_), .C2(
        keyinput198), .A(n4705), .ZN(n4708) );
  AOI22_X1 U5271 ( .A1(REG3_REG_7__SCAN_IN), .A2(keyinput179), .B1(
        REG3_REG_8__SCAN_IN), .B2(keyinput227), .ZN(n4706) );
  OAI221_X1 U5272 ( .B1(REG3_REG_7__SCAN_IN), .B2(keyinput179), .C1(
        REG3_REG_8__SCAN_IN), .C2(keyinput227), .A(n4706), .ZN(n4707) );
  NOR4_X1 U5273 ( .A1(n4710), .A2(n4709), .A3(n4708), .A4(n4707), .ZN(n4729)
         );
  AOI22_X1 U5274 ( .A1(REG3_REG_20__SCAN_IN), .A2(keyinput146), .B1(
        IR_REG_3__SCAN_IN), .B2(keyinput202), .ZN(n4711) );
  OAI221_X1 U5275 ( .B1(REG3_REG_20__SCAN_IN), .B2(keyinput146), .C1(
        IR_REG_3__SCAN_IN), .C2(keyinput202), .A(n4711), .ZN(n4718) );
  AOI22_X1 U5276 ( .A1(IR_REG_4__SCAN_IN), .A2(keyinput201), .B1(
        IR_REG_18__SCAN_IN), .B2(keyinput236), .ZN(n4712) );
  OAI221_X1 U5277 ( .B1(IR_REG_4__SCAN_IN), .B2(keyinput201), .C1(
        IR_REG_18__SCAN_IN), .C2(keyinput236), .A(n4712), .ZN(n4717) );
  AOI22_X1 U5278 ( .A1(IR_REG_20__SCAN_IN), .A2(keyinput196), .B1(
        IR_REG_31__SCAN_IN), .B2(keyinput249), .ZN(n4713) );
  OAI221_X1 U5279 ( .B1(IR_REG_20__SCAN_IN), .B2(keyinput196), .C1(
        IR_REG_31__SCAN_IN), .C2(keyinput249), .A(n4713), .ZN(n4716) );
  AOI22_X1 U5280 ( .A1(IR_REG_28__SCAN_IN), .A2(keyinput128), .B1(
        D_REG_4__SCAN_IN), .B2(keyinput174), .ZN(n4714) );
  OAI221_X1 U5281 ( .B1(IR_REG_28__SCAN_IN), .B2(keyinput128), .C1(
        D_REG_4__SCAN_IN), .C2(keyinput174), .A(n4714), .ZN(n4715) );
  NOR4_X1 U5282 ( .A1(n4718), .A2(n4717), .A3(n4716), .A4(n4715), .ZN(n4728)
         );
  AOI22_X1 U5283 ( .A1(D_REG_7__SCAN_IN), .A2(keyinput135), .B1(
        D_REG_5__SCAN_IN), .B2(keyinput233), .ZN(n4719) );
  OAI221_X1 U5284 ( .B1(D_REG_7__SCAN_IN), .B2(keyinput135), .C1(
        D_REG_5__SCAN_IN), .C2(keyinput233), .A(n4719), .ZN(n4726) );
  AOI22_X1 U5285 ( .A1(D_REG_11__SCAN_IN), .A2(keyinput213), .B1(
        D_REG_13__SCAN_IN), .B2(keyinput170), .ZN(n4720) );
  OAI221_X1 U5286 ( .B1(D_REG_11__SCAN_IN), .B2(keyinput213), .C1(
        D_REG_13__SCAN_IN), .C2(keyinput170), .A(n4720), .ZN(n4725) );
  AOI22_X1 U5287 ( .A1(D_REG_21__SCAN_IN), .A2(keyinput188), .B1(
        D_REG_26__SCAN_IN), .B2(keyinput137), .ZN(n4721) );
  OAI221_X1 U5288 ( .B1(D_REG_21__SCAN_IN), .B2(keyinput188), .C1(
        D_REG_26__SCAN_IN), .C2(keyinput137), .A(n4721), .ZN(n4724) );
  AOI22_X1 U5289 ( .A1(REG0_REG_3__SCAN_IN), .A2(keyinput244), .B1(
        REG0_REG_9__SCAN_IN), .B2(keyinput167), .ZN(n4722) );
  OAI221_X1 U5290 ( .B1(REG0_REG_3__SCAN_IN), .B2(keyinput244), .C1(
        REG0_REG_9__SCAN_IN), .C2(keyinput167), .A(n4722), .ZN(n4723) );
  NOR4_X1 U5291 ( .A1(n4726), .A2(n4725), .A3(n4724), .A4(n4723), .ZN(n4727)
         );
  NAND4_X1 U5292 ( .A1(n4730), .A2(n4729), .A3(n4728), .A4(n4727), .ZN(n4865)
         );
  AOI22_X1 U5293 ( .A1(REG0_REG_13__SCAN_IN), .A2(keyinput145), .B1(
        REG0_REG_10__SCAN_IN), .B2(keyinput189), .ZN(n4731) );
  OAI221_X1 U5294 ( .B1(REG0_REG_13__SCAN_IN), .B2(keyinput145), .C1(
        REG0_REG_10__SCAN_IN), .C2(keyinput189), .A(n4731), .ZN(n4738) );
  AOI22_X1 U5295 ( .A1(REG0_REG_17__SCAN_IN), .A2(keyinput226), .B1(
        REG0_REG_23__SCAN_IN), .B2(keyinput139), .ZN(n4732) );
  OAI221_X1 U5296 ( .B1(REG0_REG_17__SCAN_IN), .B2(keyinput226), .C1(
        REG0_REG_23__SCAN_IN), .C2(keyinput139), .A(n4732), .ZN(n4737) );
  AOI22_X1 U5297 ( .A1(REG0_REG_31__SCAN_IN), .A2(keyinput230), .B1(
        REG0_REG_27__SCAN_IN), .B2(keyinput161), .ZN(n4733) );
  OAI221_X1 U5298 ( .B1(REG0_REG_31__SCAN_IN), .B2(keyinput230), .C1(
        REG0_REG_27__SCAN_IN), .C2(keyinput161), .A(n4733), .ZN(n4736) );
  AOI22_X1 U5299 ( .A1(REG1_REG_4__SCAN_IN), .A2(keyinput133), .B1(
        REG1_REG_5__SCAN_IN), .B2(keyinput129), .ZN(n4734) );
  OAI221_X1 U5300 ( .B1(REG1_REG_4__SCAN_IN), .B2(keyinput133), .C1(
        REG1_REG_5__SCAN_IN), .C2(keyinput129), .A(n4734), .ZN(n4735) );
  NOR4_X1 U5301 ( .A1(n4738), .A2(n4737), .A3(n4736), .A4(n4735), .ZN(n4766)
         );
  AOI22_X1 U5302 ( .A1(REG1_REG_11__SCAN_IN), .A2(keyinput255), .B1(
        REG1_REG_8__SCAN_IN), .B2(keyinput183), .ZN(n4739) );
  OAI221_X1 U5303 ( .B1(REG1_REG_11__SCAN_IN), .B2(keyinput255), .C1(
        REG1_REG_8__SCAN_IN), .C2(keyinput183), .A(n4739), .ZN(n4746) );
  AOI22_X1 U5304 ( .A1(REG1_REG_14__SCAN_IN), .A2(keyinput251), .B1(
        REG1_REG_16__SCAN_IN), .B2(keyinput216), .ZN(n4740) );
  OAI221_X1 U5305 ( .B1(REG1_REG_14__SCAN_IN), .B2(keyinput251), .C1(
        REG1_REG_16__SCAN_IN), .C2(keyinput216), .A(n4740), .ZN(n4745) );
  AOI22_X1 U5306 ( .A1(REG2_REG_2__SCAN_IN), .A2(keyinput235), .B1(
        REG1_REG_23__SCAN_IN), .B2(keyinput176), .ZN(n4741) );
  OAI221_X1 U5307 ( .B1(REG2_REG_2__SCAN_IN), .B2(keyinput235), .C1(
        REG1_REG_23__SCAN_IN), .C2(keyinput176), .A(n4741), .ZN(n4744) );
  AOI22_X1 U5308 ( .A1(REG2_REG_18__SCAN_IN), .A2(keyinput190), .B1(
        REG2_REG_16__SCAN_IN), .B2(keyinput149), .ZN(n4742) );
  OAI221_X1 U5309 ( .B1(REG2_REG_18__SCAN_IN), .B2(keyinput190), .C1(
        REG2_REG_16__SCAN_IN), .C2(keyinput149), .A(n4742), .ZN(n4743) );
  NOR4_X1 U5310 ( .A1(n4746), .A2(n4745), .A3(n4744), .A4(n4743), .ZN(n4765)
         );
  AOI22_X1 U5311 ( .A1(REG2_REG_20__SCAN_IN), .A2(keyinput217), .B1(
        REG2_REG_25__SCAN_IN), .B2(keyinput243), .ZN(n4747) );
  OAI221_X1 U5312 ( .B1(REG2_REG_20__SCAN_IN), .B2(keyinput217), .C1(
        REG2_REG_25__SCAN_IN), .C2(keyinput243), .A(n4747), .ZN(n4754) );
  AOI22_X1 U5313 ( .A1(ADDR_REG_13__SCAN_IN), .A2(keyinput163), .B1(
        ADDR_REG_18__SCAN_IN), .B2(keyinput215), .ZN(n4748) );
  OAI221_X1 U5314 ( .B1(ADDR_REG_13__SCAN_IN), .B2(keyinput163), .C1(
        ADDR_REG_18__SCAN_IN), .C2(keyinput215), .A(n4748), .ZN(n4753) );
  AOI22_X1 U5315 ( .A1(ADDR_REG_0__SCAN_IN), .A2(keyinput214), .B1(
        ADDR_REG_3__SCAN_IN), .B2(keyinput144), .ZN(n4749) );
  OAI221_X1 U5316 ( .B1(ADDR_REG_0__SCAN_IN), .B2(keyinput214), .C1(
        ADDR_REG_3__SCAN_IN), .C2(keyinput144), .A(n4749), .ZN(n4752) );
  AOI22_X1 U5317 ( .A1(DATAO_REG_0__SCAN_IN), .A2(keyinput239), .B1(
        ADDR_REG_1__SCAN_IN), .B2(keyinput197), .ZN(n4750) );
  OAI221_X1 U5318 ( .B1(DATAO_REG_0__SCAN_IN), .B2(keyinput239), .C1(
        ADDR_REG_1__SCAN_IN), .C2(keyinput197), .A(n4750), .ZN(n4751) );
  NOR4_X1 U5319 ( .A1(n4754), .A2(n4753), .A3(n4752), .A4(n4751), .ZN(n4764)
         );
  AOI22_X1 U5320 ( .A1(DATAO_REG_15__SCAN_IN), .A2(keyinput138), .B1(
        DATAO_REG_9__SCAN_IN), .B2(keyinput148), .ZN(n4755) );
  OAI221_X1 U5321 ( .B1(DATAO_REG_15__SCAN_IN), .B2(keyinput138), .C1(
        DATAO_REG_9__SCAN_IN), .C2(keyinput148), .A(n4755), .ZN(n4762) );
  AOI22_X1 U5322 ( .A1(DATAO_REG_29__SCAN_IN), .A2(keyinput172), .B1(
        DATAO_REG_14__SCAN_IN), .B2(keyinput232), .ZN(n4756) );
  OAI221_X1 U5323 ( .B1(DATAO_REG_29__SCAN_IN), .B2(keyinput172), .C1(
        DATAO_REG_14__SCAN_IN), .C2(keyinput232), .A(n4756), .ZN(n4761) );
  AOI22_X1 U5324 ( .A1(DATAO_REG_25__SCAN_IN), .A2(keyinput191), .B1(
        REG3_REG_6__SCAN_IN), .B2(keyinput130), .ZN(n4757) );
  OAI221_X1 U5325 ( .B1(DATAO_REG_25__SCAN_IN), .B2(keyinput191), .C1(
        REG3_REG_6__SCAN_IN), .C2(keyinput130), .A(n4757), .ZN(n4760) );
  AOI22_X1 U5326 ( .A1(REG3_REG_18__SCAN_IN), .A2(keyinput147), .B1(
        REG3_REG_25__SCAN_IN), .B2(keyinput231), .ZN(n4758) );
  OAI221_X1 U5327 ( .B1(REG3_REG_18__SCAN_IN), .B2(keyinput147), .C1(
        REG3_REG_25__SCAN_IN), .C2(keyinput231), .A(n4758), .ZN(n4759) );
  NOR4_X1 U5328 ( .A1(n4762), .A2(n4761), .A3(n4760), .A4(n4759), .ZN(n4763)
         );
  NAND4_X1 U5329 ( .A1(n4766), .A2(n4765), .A3(n4764), .A4(n4763), .ZN(n4864)
         );
  AOI22_X1 U5330 ( .A1(REG2_REG_26__SCAN_IN), .A2(keyinput195), .B1(
        D_REG_8__SCAN_IN), .B2(keyinput228), .ZN(n4767) );
  OAI221_X1 U5331 ( .B1(REG2_REG_26__SCAN_IN), .B2(keyinput195), .C1(
        D_REG_8__SCAN_IN), .C2(keyinput228), .A(n4767), .ZN(n4778) );
  AOI22_X1 U5332 ( .A1(n4769), .A2(keyinput165), .B1(n4980), .B2(keyinput205), 
        .ZN(n4768) );
  OAI221_X1 U5333 ( .B1(n4769), .B2(keyinput165), .C1(n4980), .C2(keyinput205), 
        .A(n4768), .ZN(n4777) );
  INV_X1 U5334 ( .A(DATAI_18_), .ZN(n4872) );
  AOI22_X1 U5335 ( .A1(n4771), .A2(keyinput186), .B1(n4872), .B2(keyinput185), 
        .ZN(n4770) );
  OAI221_X1 U5336 ( .B1(n4771), .B2(keyinput186), .C1(n4872), .C2(keyinput185), 
        .A(n4770), .ZN(n4776) );
  AOI22_X1 U5337 ( .A1(n4774), .A2(keyinput254), .B1(keyinput220), .B2(n4773), 
        .ZN(n4772) );
  OAI221_X1 U5338 ( .B1(n4774), .B2(keyinput254), .C1(n4773), .C2(keyinput220), 
        .A(n4772), .ZN(n4775) );
  NOR4_X1 U5339 ( .A1(n4778), .A2(n4777), .A3(n4776), .A4(n4775), .ZN(n4815)
         );
  AOI22_X1 U5340 ( .A1(n4899), .A2(keyinput131), .B1(keyinput211), .B2(n4900), 
        .ZN(n4779) );
  OAI221_X1 U5341 ( .B1(n4899), .B2(keyinput131), .C1(n4900), .C2(keyinput211), 
        .A(n4779), .ZN(n4787) );
  XNOR2_X1 U5342 ( .A(keyinput150), .B(n2803), .ZN(n4786) );
  XNOR2_X1 U5343 ( .A(keyinput204), .B(n2789), .ZN(n4785) );
  XNOR2_X1 U5344 ( .A(IR_REG_12__SCAN_IN), .B(keyinput209), .ZN(n4783) );
  XNOR2_X1 U5345 ( .A(IR_REG_5__SCAN_IN), .B(keyinput175), .ZN(n4782) );
  XNOR2_X1 U5346 ( .A(IR_REG_19__SCAN_IN), .B(keyinput158), .ZN(n4781) );
  XNOR2_X1 U5347 ( .A(IR_REG_14__SCAN_IN), .B(keyinput156), .ZN(n4780) );
  NAND4_X1 U5348 ( .A1(n4783), .A2(n4782), .A3(n4781), .A4(n4780), .ZN(n4784)
         );
  NOR4_X1 U5349 ( .A1(n4787), .A2(n4786), .A3(n4785), .A4(n4784), .ZN(n4814)
         );
  AOI22_X1 U5350 ( .A1(n4909), .A2(keyinput169), .B1(keyinput212), .B2(n4930), 
        .ZN(n4788) );
  OAI221_X1 U5351 ( .B1(n4909), .B2(keyinput169), .C1(n4930), .C2(keyinput212), 
        .A(n4788), .ZN(n4798) );
  AOI22_X1 U5352 ( .A1(n4913), .A2(keyinput225), .B1(keyinput166), .B2(n4912), 
        .ZN(n4789) );
  OAI221_X1 U5353 ( .B1(n4913), .B2(keyinput225), .C1(n4912), .C2(keyinput166), 
        .A(n4789), .ZN(n4797) );
  AOI22_X1 U5354 ( .A1(n4792), .A2(keyinput162), .B1(n4791), .B2(keyinput178), 
        .ZN(n4790) );
  OAI221_X1 U5355 ( .B1(n4792), .B2(keyinput162), .C1(n4791), .C2(keyinput178), 
        .A(n4790), .ZN(n4796) );
  XNOR2_X1 U5356 ( .A(D_REG_0__SCAN_IN), .B(keyinput184), .ZN(n4794) );
  XNOR2_X1 U5357 ( .A(IR_REG_26__SCAN_IN), .B(keyinput153), .ZN(n4793) );
  NAND2_X1 U5358 ( .A1(n4794), .A2(n4793), .ZN(n4795) );
  NOR4_X1 U5359 ( .A1(n4798), .A2(n4797), .A3(n4796), .A4(n4795), .ZN(n4813)
         );
  AOI22_X1 U5360 ( .A1(n4801), .A2(keyinput203), .B1(n4800), .B2(keyinput223), 
        .ZN(n4799) );
  OAI221_X1 U5361 ( .B1(n4801), .B2(keyinput203), .C1(n4800), .C2(keyinput223), 
        .A(n4799), .ZN(n4811) );
  AOI22_X1 U5362 ( .A1(n4804), .A2(keyinput200), .B1(n4803), .B2(keyinput152), 
        .ZN(n4802) );
  OAI221_X1 U5363 ( .B1(n4804), .B2(keyinput200), .C1(n4803), .C2(keyinput152), 
        .A(n4802), .ZN(n4810) );
  AOI22_X1 U5364 ( .A1(n2720), .A2(keyinput253), .B1(keyinput248), .B2(n4892), 
        .ZN(n4805) );
  OAI221_X1 U5365 ( .B1(n2720), .B2(keyinput253), .C1(n4892), .C2(keyinput248), 
        .A(n4805), .ZN(n4809) );
  AOI22_X1 U5366 ( .A1(n4807), .A2(keyinput180), .B1(n4934), .B2(keyinput136), 
        .ZN(n4806) );
  OAI221_X1 U5367 ( .B1(n4807), .B2(keyinput180), .C1(n4934), .C2(keyinput136), 
        .A(n4806), .ZN(n4808) );
  NOR4_X1 U5368 ( .A1(n4811), .A2(n4810), .A3(n4809), .A4(n4808), .ZN(n4812)
         );
  NAND4_X1 U5369 ( .A1(n4815), .A2(n4814), .A3(n4813), .A4(n4812), .ZN(n4863)
         );
  AOI22_X1 U5370 ( .A1(n4945), .A2(keyinput242), .B1(keyinput159), .B2(n4879), 
        .ZN(n4816) );
  OAI221_X1 U5371 ( .B1(n4945), .B2(keyinput242), .C1(n4879), .C2(keyinput159), 
        .A(n4816), .ZN(n4825) );
  AOI22_X1 U5372 ( .A1(n2635), .A2(keyinput210), .B1(n4935), .B2(keyinput234), 
        .ZN(n4817) );
  OAI221_X1 U5373 ( .B1(n2635), .B2(keyinput210), .C1(n4935), .C2(keyinput234), 
        .A(n4817), .ZN(n4824) );
  AOI22_X1 U5374 ( .A1(n4941), .A2(keyinput187), .B1(n4819), .B2(keyinput229), 
        .ZN(n4818) );
  OAI221_X1 U5375 ( .B1(n4941), .B2(keyinput187), .C1(n4819), .C2(keyinput229), 
        .A(n4818), .ZN(n4823) );
  AOI22_X1 U5376 ( .A1(n4821), .A2(keyinput168), .B1(keyinput157), .B2(n4944), 
        .ZN(n4820) );
  OAI221_X1 U5377 ( .B1(n4821), .B2(keyinput168), .C1(n4944), .C2(keyinput157), 
        .A(n4820), .ZN(n4822) );
  NOR4_X1 U5378 ( .A1(n4825), .A2(n4824), .A3(n4823), .A4(n4822), .ZN(n4861)
         );
  AOI22_X1 U5379 ( .A1(n4977), .A2(keyinput182), .B1(n3221), .B2(keyinput221), 
        .ZN(n4826) );
  OAI221_X1 U5380 ( .B1(n4977), .B2(keyinput182), .C1(n3221), .C2(keyinput221), 
        .A(n4826), .ZN(n4835) );
  AOI22_X1 U5381 ( .A1(n2636), .A2(keyinput134), .B1(n3430), .B2(keyinput194), 
        .ZN(n4827) );
  OAI221_X1 U5382 ( .B1(n2636), .B2(keyinput134), .C1(n3430), .C2(keyinput194), 
        .A(n4827), .ZN(n4834) );
  AOI22_X1 U5383 ( .A1(n4829), .A2(keyinput245), .B1(n4079), .B2(keyinput246), 
        .ZN(n4828) );
  OAI221_X1 U5384 ( .B1(n4829), .B2(keyinput245), .C1(n4079), .C2(keyinput246), 
        .A(n4828), .ZN(n4833) );
  AOI22_X1 U5385 ( .A1(n4831), .A2(keyinput154), .B1(keyinput141), .B2(n3229), 
        .ZN(n4830) );
  OAI221_X1 U5386 ( .B1(n4831), .B2(keyinput154), .C1(n3229), .C2(keyinput141), 
        .A(n4830), .ZN(n4832) );
  NOR4_X1 U5387 ( .A1(n4835), .A2(n4834), .A3(n4833), .A4(n4832), .ZN(n4860)
         );
  AOI22_X1 U5388 ( .A1(n3188), .A2(keyinput224), .B1(keyinput247), .B2(n4837), 
        .ZN(n4836) );
  OAI221_X1 U5389 ( .B1(n3188), .B2(keyinput224), .C1(n4837), .C2(keyinput247), 
        .A(n4836), .ZN(n4847) );
  INV_X1 U5390 ( .A(ADDR_REG_2__SCAN_IN), .ZN(n4882) );
  AOI22_X1 U5391 ( .A1(n4882), .A2(keyinput164), .B1(keyinput207), .B2(n4839), 
        .ZN(n4838) );
  OAI221_X1 U5392 ( .B1(n4882), .B2(keyinput164), .C1(n4839), .C2(keyinput207), 
        .A(n4838), .ZN(n4846) );
  AOI22_X1 U5393 ( .A1(n4841), .A2(keyinput237), .B1(keyinput193), .B2(n4979), 
        .ZN(n4840) );
  OAI221_X1 U5394 ( .B1(n4841), .B2(keyinput237), .C1(n4979), .C2(keyinput193), 
        .A(n4840), .ZN(n4845) );
  AOI22_X1 U5395 ( .A1(n4982), .A2(keyinput177), .B1(keyinput192), .B2(n4843), 
        .ZN(n4842) );
  OAI221_X1 U5396 ( .B1(n4982), .B2(keyinput177), .C1(n4843), .C2(keyinput192), 
        .A(n4842), .ZN(n4844) );
  NOR4_X1 U5397 ( .A1(n4847), .A2(n4846), .A3(n4845), .A4(n4844), .ZN(n4859)
         );
  AOI22_X1 U5398 ( .A1(n4966), .A2(keyinput142), .B1(keyinput173), .B2(n4983), 
        .ZN(n4848) );
  OAI221_X1 U5399 ( .B1(n4966), .B2(keyinput142), .C1(n4983), .C2(keyinput173), 
        .A(n4848), .ZN(n4857) );
  AOI22_X1 U5400 ( .A1(n4958), .A2(keyinput222), .B1(keyinput250), .B2(n4850), 
        .ZN(n4849) );
  OAI221_X1 U5401 ( .B1(n4958), .B2(keyinput222), .C1(n4850), .C2(keyinput250), 
        .A(n4849), .ZN(n4856) );
  AOI22_X1 U5402 ( .A1(n4960), .A2(keyinput155), .B1(n4852), .B2(keyinput240), 
        .ZN(n4851) );
  OAI221_X1 U5403 ( .B1(n4960), .B2(keyinput155), .C1(n4852), .C2(keyinput240), 
        .A(n4851), .ZN(n4855) );
  AOI22_X1 U5404 ( .A1(n2763), .A2(keyinput252), .B1(n4906), .B2(keyinput208), 
        .ZN(n4853) );
  OAI221_X1 U5405 ( .B1(n2763), .B2(keyinput252), .C1(n4906), .C2(keyinput208), 
        .A(n4853), .ZN(n4854) );
  NOR4_X1 U5406 ( .A1(n4857), .A2(n4856), .A3(n4855), .A4(n4854), .ZN(n4858)
         );
  NAND4_X1 U5407 ( .A1(n4861), .A2(n4860), .A3(n4859), .A4(n4858), .ZN(n4862)
         );
  NOR4_X1 U5408 ( .A1(n4865), .A2(n4864), .A3(n4863), .A4(n4862), .ZN(n4994)
         );
  AOI22_X1 U5409 ( .A1(n4867), .A2(keyinput18), .B1(keyinput96), .B2(n3188), 
        .ZN(n4866) );
  OAI221_X1 U5410 ( .B1(n4867), .B2(keyinput18), .C1(n3188), .C2(keyinput96), 
        .A(n4866), .ZN(n4877) );
  AOI22_X1 U5411 ( .A1(n3229), .A2(keyinput13), .B1(n4005), .B2(keyinput67), 
        .ZN(n4868) );
  OAI221_X1 U5412 ( .B1(n3229), .B2(keyinput13), .C1(n4005), .C2(keyinput67), 
        .A(n4868), .ZN(n4876) );
  INV_X1 U5413 ( .A(DATAI_28_), .ZN(n4870) );
  AOI22_X1 U5414 ( .A1(n4079), .A2(keyinput118), .B1(n4870), .B2(keyinput91), 
        .ZN(n4869) );
  OAI221_X1 U5415 ( .B1(n4079), .B2(keyinput118), .C1(n4870), .C2(keyinput91), 
        .A(n4869), .ZN(n4875) );
  INV_X1 U5416 ( .A(DATAI_20_), .ZN(n4873) );
  AOI22_X1 U5417 ( .A1(n4873), .A2(keyinput4), .B1(keyinput57), .B2(n4872), 
        .ZN(n4871) );
  OAI221_X1 U5418 ( .B1(n4873), .B2(keyinput4), .C1(n4872), .C2(keyinput57), 
        .A(n4871), .ZN(n4874) );
  NOR4_X1 U5419 ( .A1(n4877), .A2(n4876), .A3(n4875), .A4(n4874), .ZN(n4924)
         );
  AOI22_X1 U5420 ( .A1(n4880), .A2(keyinput127), .B1(n4879), .B2(keyinput31), 
        .ZN(n4878) );
  OAI221_X1 U5421 ( .B1(n4880), .B2(keyinput127), .C1(n4879), .C2(keyinput31), 
        .A(n4878), .ZN(n4890) );
  AOI22_X1 U5422 ( .A1(n4883), .A2(keyinput15), .B1(keyinput36), .B2(n4882), 
        .ZN(n4881) );
  OAI221_X1 U5423 ( .B1(n4883), .B2(keyinput15), .C1(n4882), .C2(keyinput36), 
        .A(n4881), .ZN(n4889) );
  AOI22_X1 U5424 ( .A1(n2403), .A2(keyinput5), .B1(n2636), .B2(keyinput6), 
        .ZN(n4884) );
  OAI221_X1 U5425 ( .B1(n2403), .B2(keyinput5), .C1(n2636), .C2(keyinput6), 
        .A(n4884), .ZN(n4888) );
  XOR2_X1 U5426 ( .A(n2789), .B(keyinput76), .Z(n4886) );
  XNOR2_X1 U5427 ( .A(IR_REG_18__SCAN_IN), .B(keyinput108), .ZN(n4885) );
  NAND2_X1 U5428 ( .A1(n4886), .A2(n4885), .ZN(n4887) );
  NOR4_X1 U5429 ( .A1(n4890), .A2(n4889), .A3(n4888), .A4(n4887), .ZN(n4923)
         );
  AOI22_X1 U5430 ( .A1(n4892), .A2(keyinput120), .B1(n2700), .B2(keyinput61), 
        .ZN(n4891) );
  OAI221_X1 U5431 ( .B1(n4892), .B2(keyinput120), .C1(n2700), .C2(keyinput61), 
        .A(n4891), .ZN(n4904) );
  INV_X1 U5432 ( .A(DATAI_3_), .ZN(n4894) );
  AOI22_X1 U5433 ( .A1(n2651), .A2(keyinput51), .B1(keyinput12), .B2(n4894), 
        .ZN(n4893) );
  OAI221_X1 U5434 ( .B1(n2651), .B2(keyinput51), .C1(n4894), .C2(keyinput12), 
        .A(n4893), .ZN(n4903) );
  INV_X1 U5435 ( .A(DATAI_4_), .ZN(n4897) );
  AOI22_X1 U5436 ( .A1(n4897), .A2(keyinput43), .B1(n4896), .B2(keyinput73), 
        .ZN(n4895) );
  OAI221_X1 U5437 ( .B1(n4897), .B2(keyinput43), .C1(n4896), .C2(keyinput73), 
        .A(n4895), .ZN(n4902) );
  AOI22_X1 U5438 ( .A1(n4900), .A2(keyinput83), .B1(n4899), .B2(keyinput3), 
        .ZN(n4898) );
  OAI221_X1 U5439 ( .B1(n4900), .B2(keyinput83), .C1(n4899), .C2(keyinput3), 
        .A(n4898), .ZN(n4901) );
  NOR4_X1 U5440 ( .A1(n4904), .A2(n4903), .A3(n4902), .A4(n4901), .ZN(n4922)
         );
  AOI22_X1 U5441 ( .A1(n4907), .A2(keyinput7), .B1(keyinput80), .B2(n4906), 
        .ZN(n4905) );
  OAI221_X1 U5442 ( .B1(n4907), .B2(keyinput7), .C1(n4906), .C2(keyinput80), 
        .A(n4905), .ZN(n4920) );
  AOI22_X1 U5443 ( .A1(n4910), .A2(keyinput105), .B1(keyinput41), .B2(n4909), 
        .ZN(n4908) );
  OAI221_X1 U5444 ( .B1(n4910), .B2(keyinput105), .C1(n4909), .C2(keyinput41), 
        .A(n4908), .ZN(n4919) );
  AOI22_X1 U5445 ( .A1(n4913), .A2(keyinput97), .B1(keyinput38), .B2(n4912), 
        .ZN(n4911) );
  OAI221_X1 U5446 ( .B1(n4913), .B2(keyinput97), .C1(n4912), .C2(keyinput38), 
        .A(n4911), .ZN(n4918) );
  XOR2_X1 U5447 ( .A(n4914), .B(keyinput53), .Z(n4916) );
  XNOR2_X1 U5448 ( .A(IR_REG_20__SCAN_IN), .B(keyinput68), .ZN(n4915) );
  NAND2_X1 U5449 ( .A1(n4916), .A2(n4915), .ZN(n4917) );
  NOR4_X1 U5450 ( .A1(n4920), .A2(n4919), .A3(n4918), .A4(n4917), .ZN(n4921)
         );
  NAND4_X1 U5451 ( .A1(n4924), .A2(n4923), .A3(n4922), .A4(n4921), .ZN(n4993)
         );
  AOI22_X1 U5452 ( .A1(n4927), .A2(keyinput100), .B1(keyinput9), .B2(n4926), 
        .ZN(n4925) );
  OAI221_X1 U5453 ( .B1(n4927), .B2(keyinput100), .C1(n4926), .C2(keyinput9), 
        .A(n4925), .ZN(n4939) );
  AOI22_X1 U5454 ( .A1(n4930), .A2(keyinput84), .B1(keyinput60), .B2(n4929), 
        .ZN(n4928) );
  OAI221_X1 U5455 ( .B1(n4930), .B2(keyinput84), .C1(n4929), .C2(keyinput60), 
        .A(n4928), .ZN(n4938) );
  AOI22_X1 U5456 ( .A1(n4932), .A2(keyinput98), .B1(n2803), .B2(keyinput22), 
        .ZN(n4931) );
  OAI221_X1 U5457 ( .B1(n4932), .B2(keyinput98), .C1(n2803), .C2(keyinput22), 
        .A(n4931), .ZN(n4937) );
  AOI22_X1 U5458 ( .A1(n4935), .A2(keyinput106), .B1(n4934), .B2(keyinput8), 
        .ZN(n4933) );
  OAI221_X1 U5459 ( .B1(n4935), .B2(keyinput106), .C1(n4934), .C2(keyinput8), 
        .A(n4933), .ZN(n4936) );
  NOR4_X1 U5460 ( .A1(n4939), .A2(n4938), .A3(n4937), .A4(n4936), .ZN(n4991)
         );
  AOI22_X1 U5461 ( .A1(n4942), .A2(keyinput48), .B1(keyinput59), .B2(n4941), 
        .ZN(n4940) );
  OAI221_X1 U5462 ( .B1(n4942), .B2(keyinput48), .C1(n4941), .C2(keyinput59), 
        .A(n4940), .ZN(n4955) );
  AOI22_X1 U5463 ( .A1(n4945), .A2(keyinput114), .B1(keyinput29), .B2(n4944), 
        .ZN(n4943) );
  OAI221_X1 U5464 ( .B1(n4945), .B2(keyinput114), .C1(n4944), .C2(keyinput29), 
        .A(n4943), .ZN(n4954) );
  INV_X1 U5465 ( .A(DATAI_19_), .ZN(n4947) );
  AOI22_X1 U5466 ( .A1(n4948), .A2(keyinput99), .B1(keyinput110), .B2(n4947), 
        .ZN(n4946) );
  OAI221_X1 U5467 ( .B1(n4948), .B2(keyinput99), .C1(n4947), .C2(keyinput110), 
        .A(n4946), .ZN(n4953) );
  AOI22_X1 U5468 ( .A1(n4951), .A2(keyinput111), .B1(n4950), .B2(keyinput87), 
        .ZN(n4949) );
  OAI221_X1 U5469 ( .B1(n4951), .B2(keyinput111), .C1(n4950), .C2(keyinput87), 
        .A(n4949), .ZN(n4952) );
  NOR4_X1 U5470 ( .A1(n4955), .A2(n4954), .A3(n4953), .A4(n4952), .ZN(n4990)
         );
  AOI22_X1 U5471 ( .A1(n4958), .A2(keyinput94), .B1(n4957), .B2(keyinput32), 
        .ZN(n4956) );
  OAI221_X1 U5472 ( .B1(n4958), .B2(keyinput94), .C1(n4957), .C2(keyinput32), 
        .A(n4956), .ZN(n4971) );
  AOI22_X1 U5473 ( .A1(n4961), .A2(keyinput56), .B1(keyinput27), .B2(n4960), 
        .ZN(n4959) );
  OAI221_X1 U5474 ( .B1(n4961), .B2(keyinput56), .C1(n4960), .C2(keyinput27), 
        .A(n4959), .ZN(n4970) );
  INV_X1 U5475 ( .A(ADDR_REG_13__SCAN_IN), .ZN(n4964) );
  AOI22_X1 U5476 ( .A1(n4964), .A2(keyinput35), .B1(n4963), .B2(keyinput2), 
        .ZN(n4962) );
  OAI221_X1 U5477 ( .B1(n4964), .B2(keyinput35), .C1(n4963), .C2(keyinput2), 
        .A(n4962), .ZN(n4969) );
  AOI22_X1 U5478 ( .A1(n4967), .A2(keyinput19), .B1(keyinput14), .B2(n4966), 
        .ZN(n4965) );
  OAI221_X1 U5479 ( .B1(n4967), .B2(keyinput19), .C1(n4966), .C2(keyinput14), 
        .A(n4965), .ZN(n4968) );
  NOR4_X1 U5480 ( .A1(n4971), .A2(n4970), .A3(n4969), .A4(n4968), .ZN(n4989)
         );
  AOI22_X1 U5481 ( .A1(n4974), .A2(keyinput63), .B1(n4973), .B2(keyinput71), 
        .ZN(n4972) );
  OAI221_X1 U5482 ( .B1(n4974), .B2(keyinput63), .C1(n4973), .C2(keyinput71), 
        .A(n4972), .ZN(n4987) );
  INV_X1 U5483 ( .A(ADDR_REG_3__SCAN_IN), .ZN(n4976) );
  AOI22_X1 U5484 ( .A1(n4977), .A2(keyinput54), .B1(keyinput16), .B2(n4976), 
        .ZN(n4975) );
  OAI221_X1 U5485 ( .B1(n4977), .B2(keyinput54), .C1(n4976), .C2(keyinput16), 
        .A(n4975), .ZN(n4986) );
  AOI22_X1 U5486 ( .A1(n4980), .A2(keyinput77), .B1(keyinput65), .B2(n4979), 
        .ZN(n4978) );
  OAI221_X1 U5487 ( .B1(n4980), .B2(keyinput77), .C1(n4979), .C2(keyinput65), 
        .A(n4978), .ZN(n4985) );
  AOI22_X1 U5488 ( .A1(n4983), .A2(keyinput45), .B1(n4982), .B2(keyinput49), 
        .ZN(n4981) );
  OAI221_X1 U5489 ( .B1(n4983), .B2(keyinput45), .C1(n4982), .C2(keyinput49), 
        .A(n4981), .ZN(n4984) );
  NOR4_X1 U5490 ( .A1(n4987), .A2(n4986), .A3(n4985), .A4(n4984), .ZN(n4988)
         );
  NAND4_X1 U5491 ( .A1(n4991), .A2(n4990), .A3(n4989), .A4(n4988), .ZN(n4992)
         );
  NOR3_X1 U5492 ( .A1(n4994), .A2(n4993), .A3(n4992), .ZN(n5032) );
  OAI22_X1 U5493 ( .A1(IR_REG_12__SCAN_IN), .A2(keyinput81), .B1(keyinput92), 
        .B2(DATAI_7_), .ZN(n4995) );
  AOI221_X1 U5494 ( .B1(IR_REG_12__SCAN_IN), .B2(keyinput81), .C1(DATAI_7_), 
        .C2(keyinput92), .A(n4995), .ZN(n5002) );
  OAI22_X1 U5495 ( .A1(IR_REG_5__SCAN_IN), .A2(keyinput47), .B1(keyinput74), 
        .B2(IR_REG_3__SCAN_IN), .ZN(n4996) );
  AOI221_X1 U5496 ( .B1(IR_REG_5__SCAN_IN), .B2(keyinput47), .C1(
        IR_REG_3__SCAN_IN), .C2(keyinput74), .A(n4996), .ZN(n5001) );
  OAI22_X1 U5497 ( .A1(D_REG_10__SCAN_IN), .A2(keyinput34), .B1(
        D_REG_29__SCAN_IN), .B2(keyinput95), .ZN(n4997) );
  AOI221_X1 U5498 ( .B1(D_REG_10__SCAN_IN), .B2(keyinput34), .C1(keyinput95), 
        .C2(D_REG_29__SCAN_IN), .A(n4997), .ZN(n5000) );
  OAI22_X1 U5499 ( .A1(IR_REG_19__SCAN_IN), .A2(keyinput30), .B1(
        D_REG_12__SCAN_IN), .B2(keyinput50), .ZN(n4998) );
  AOI221_X1 U5500 ( .B1(IR_REG_19__SCAN_IN), .B2(keyinput30), .C1(keyinput50), 
        .C2(D_REG_12__SCAN_IN), .A(n4998), .ZN(n4999) );
  NAND4_X1 U5501 ( .A1(n5002), .A2(n5001), .A3(n5000), .A4(n4999), .ZN(n5030)
         );
  OAI22_X1 U5502 ( .A1(REG1_REG_8__SCAN_IN), .A2(keyinput55), .B1(
        REG1_REG_14__SCAN_IN), .B2(keyinput123), .ZN(n5003) );
  AOI221_X1 U5503 ( .B1(REG1_REG_8__SCAN_IN), .B2(keyinput55), .C1(keyinput123), .C2(REG1_REG_14__SCAN_IN), .A(n5003), .ZN(n5010) );
  OAI22_X1 U5504 ( .A1(REG0_REG_9__SCAN_IN), .A2(keyinput39), .B1(
        REG0_REG_13__SCAN_IN), .B2(keyinput17), .ZN(n5004) );
  AOI221_X1 U5505 ( .B1(REG0_REG_9__SCAN_IN), .B2(keyinput39), .C1(keyinput17), 
        .C2(REG0_REG_13__SCAN_IN), .A(n5004), .ZN(n5009) );
  OAI22_X1 U5506 ( .A1(REG0_REG_8__SCAN_IN), .A2(keyinput24), .B1(
        REG0_REG_11__SCAN_IN), .B2(keyinput125), .ZN(n5005) );
  AOI221_X1 U5507 ( .B1(REG0_REG_8__SCAN_IN), .B2(keyinput24), .C1(keyinput125), .C2(REG0_REG_11__SCAN_IN), .A(n5005), .ZN(n5008) );
  OAI22_X1 U5508 ( .A1(REG3_REG_15__SCAN_IN), .A2(keyinput124), .B1(
        REG0_REG_7__SCAN_IN), .B2(keyinput72), .ZN(n5006) );
  AOI221_X1 U5509 ( .B1(REG3_REG_15__SCAN_IN), .B2(keyinput124), .C1(
        keyinput72), .C2(REG0_REG_7__SCAN_IN), .A(n5006), .ZN(n5007) );
  NAND4_X1 U5510 ( .A1(n5010), .A2(n5009), .A3(n5008), .A4(n5007), .ZN(n5029)
         );
  OAI22_X1 U5511 ( .A1(DATAI_16_), .A2(keyinput126), .B1(keyinput64), .B2(
        DATAO_REG_12__SCAN_IN), .ZN(n5011) );
  AOI221_X1 U5512 ( .B1(DATAI_16_), .B2(keyinput126), .C1(
        DATAO_REG_12__SCAN_IN), .C2(keyinput64), .A(n5011), .ZN(n5018) );
  OAI22_X1 U5513 ( .A1(IR_REG_26__SCAN_IN), .A2(keyinput25), .B1(keyinput37), 
        .B2(DATAI_31_), .ZN(n5012) );
  AOI221_X1 U5514 ( .B1(IR_REG_26__SCAN_IN), .B2(keyinput25), .C1(DATAI_31_), 
        .C2(keyinput37), .A(n5012), .ZN(n5017) );
  OAI22_X1 U5515 ( .A1(n4161), .A2(keyinput62), .B1(keyinput119), .B2(
        ADDR_REG_5__SCAN_IN), .ZN(n5013) );
  AOI221_X1 U5516 ( .B1(n4161), .B2(keyinput62), .C1(ADDR_REG_5__SCAN_IN), 
        .C2(keyinput119), .A(n5013), .ZN(n5016) );
  OAI22_X1 U5517 ( .A1(DATAO_REG_2__SCAN_IN), .A2(keyinput79), .B1(keyinput122), .B2(DATAO_REG_30__SCAN_IN), .ZN(n5014) );
  AOI221_X1 U5518 ( .B1(DATAO_REG_2__SCAN_IN), .B2(keyinput79), .C1(
        DATAO_REG_30__SCAN_IN), .C2(keyinput122), .A(n5014), .ZN(n5015) );
  NAND4_X1 U5519 ( .A1(n5018), .A2(n5017), .A3(n5016), .A4(n5015), .ZN(n5028)
         );
  OAI22_X1 U5520 ( .A1(REG1_REG_28__SCAN_IN), .A2(keyinput101), .B1(
        DATAO_REG_29__SCAN_IN), .B2(keyinput44), .ZN(n5019) );
  AOI221_X1 U5521 ( .B1(REG1_REG_28__SCAN_IN), .B2(keyinput101), .C1(
        keyinput44), .C2(DATAO_REG_29__SCAN_IN), .A(n5019), .ZN(n5026) );
  OAI22_X1 U5522 ( .A1(D_REG_24__SCAN_IN), .A2(keyinput75), .B1(
        REG0_REG_16__SCAN_IN), .B2(keyinput52), .ZN(n5020) );
  AOI221_X1 U5523 ( .B1(D_REG_24__SCAN_IN), .B2(keyinput75), .C1(keyinput52), 
        .C2(REG0_REG_16__SCAN_IN), .A(n5020), .ZN(n5025) );
  OAI22_X1 U5524 ( .A1(ADDR_REG_1__SCAN_IN), .A2(keyinput69), .B1(
        DATAO_REG_7__SCAN_IN), .B2(keyinput109), .ZN(n5021) );
  AOI221_X1 U5525 ( .B1(ADDR_REG_1__SCAN_IN), .B2(keyinput69), .C1(keyinput109), .C2(DATAO_REG_7__SCAN_IN), .A(n5021), .ZN(n5024) );
  OAI22_X1 U5526 ( .A1(IR_REG_28__SCAN_IN), .A2(keyinput0), .B1(keyinput40), 
        .B2(REG1_REG_30__SCAN_IN), .ZN(n5022) );
  AOI221_X1 U5527 ( .B1(IR_REG_28__SCAN_IN), .B2(keyinput0), .C1(
        REG1_REG_30__SCAN_IN), .C2(keyinput40), .A(n5022), .ZN(n5023) );
  NAND4_X1 U5528 ( .A1(n5026), .A2(n5025), .A3(n5024), .A4(n5023), .ZN(n5027)
         );
  NOR4_X1 U5529 ( .A1(n5030), .A2(n5029), .A3(n5028), .A4(n5027), .ZN(n5031)
         );
  NAND3_X1 U5530 ( .A1(n5033), .A2(n5032), .A3(n5031), .ZN(n5052) );
  NOR2_X1 U5531 ( .A1(n5035), .A2(n5034), .ZN(n5040) );
  INV_X1 U5532 ( .A(n5036), .ZN(n5037) );
  OAI211_X1 U5533 ( .C1(n5040), .C2(n5039), .A(n5038), .B(n5037), .ZN(n5050)
         );
  OAI211_X1 U5534 ( .C1(n5044), .C2(n5043), .A(n5042), .B(n5041), .ZN(n5049)
         );
  AOI22_X1 U5535 ( .A1(n5045), .A2(ADDR_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(U3149), .ZN(n5048) );
  NAND2_X1 U5536 ( .A1(n5046), .A2(n3143), .ZN(n5047) );
  NAND4_X1 U5537 ( .A1(n5050), .A2(n5049), .A3(n5048), .A4(n5047), .ZN(n5051)
         );
  XNOR2_X1 U5538 ( .A(n5052), .B(n5051), .ZN(U3241) );
  CLKBUF_X1 U2480 ( .A(n2944), .Z(n2987) );
  INV_X2 U4070 ( .A(n4581), .ZN(n3576) );
endmodule

