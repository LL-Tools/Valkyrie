

module b15_C_SARLock_k_64_9 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, 
        READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, 
        CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, 
        REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, 
        FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, U3445, U3446, U3447, U3448, U3213, U3212, 
        U3211, U3210, U3209, U3208, U3207, U3206, U3205, U3204, U3203, U3202, 
        U3201, U3200, U3199, U3198, U3197, U3196, U3195, U3194, U3193, U3192, 
        U3191, U3190, U3189, U3188, U3187, U3186, U3185, U3184, U3183, U3182, 
        U3181, U3451, U3452, U3180, U3179, U3178, U3177, U3176, U3175, U3174, 
        U3173, U3172, U3171, U3170, U3169, U3168, U3167, U3166, U3165, U3164, 
        U3163, U3162, U3161, U3160, U3159, U3158, U3157, U3156, U3155, U3154, 
        U3153, U3152, U3151, U3453, U3150, U3149, U3148, U3147, U3146, U3145, 
        U3144, U3143, U3142, U3141, U3140, U3139, U3138, U3137, U3136, U3135, 
        U3134, U3133, U3132, U3131, U3130, U3129, U3128, U3127, U3126, U3125, 
        U3124, U3123, U3122, U3121, U3120, U3119, U3118, U3117, U3116, U3115, 
        U3114, U3113, U3112, U3111, U3110, U3109, U3108, U3107, U3106, U3105, 
        U3104, U3103, U3102, U3101, U3100, U3099, U3098, U3097, U3096, U3095, 
        U3094, U3093, U3092, U3091, U3090, U3089, U3088, U3087, U3086, U3085, 
        U3084, U3083, U3082, U3081, U3080, U3079, U3078, U3077, U3076, U3075, 
        U3074, U3073, U3072, U3071, U3070, U3069, U3068, U3067, U3066, U3065, 
        U3064, U3063, U3062, U3061, U3060, U3059, U3058, U3057, U3056, U3055, 
        U3054, U3053, U3052, U3051, U3050, U3049, U3048, U3047, U3046, U3045, 
        U3044, U3043, U3042, U3041, U3040, U3039, U3038, U3037, U3036, U3035, 
        U3034, U3033, U3032, U3031, U3030, U3029, U3028, U3027, U3026, U3025, 
        U3024, U3023, U3022, U3021, U3020, U3455, U3456, U3459, U3460, U3461, 
        U3019, U3462, U3463, U3464, U3465, U3018, U3017, U3016, U3015, U3014, 
        U3013, U3012, U3011, U3010, U3009, U3008, U3007, U3006, U3005, U3004, 
        U3003, U3002, U3001, U3000, U2999, U2998, U2997, U2996, U2995, U2994, 
        U2993, U2992, U2991, U2990, U2989, U2988, U2987, U2986, U2985, U2984, 
        U2983, U2982, U2981, U2980, U2979, U2978, U2977, U2976, U2975, U2974, 
        U2973, U2972, U2971, U2970, U2969, U2968, U2967, U2966, U2965, U2964, 
        U2963, U2962, U2961, U2960, U2959, U2958, U2957, U2956, U2955, U2954, 
        U2953, U2952, U2951, U2950, U2949, U2948, U2947, U2946, U2945, U2944, 
        U2943, U2942, U2941, U2940, U2939, U2938, U2937, U2936, U2935, U2934, 
        U2933, U2932, U2931, U2930, U2929, U2928, U2927, U2926, U2925, U2924, 
        U2923, U2922, U2921, U2920, U2919, U2918, U2917, U2916, U2915, U2914, 
        U2913, U2912, U2911, U2910, U2909, U2908, U2907, U2906, U2905, U2904, 
        U2903, U2902, U2901, U2900, U2899, U2898, U2897, U2896, U2895, U2894, 
        U2893, U2892, U2891, U2890, U2889, U2888, U2887, U2886, U2885, U2884, 
        U2883, U2882, U2881, U2880, U2879, U2878, U2877, U2876, U2875, U2874, 
        U2873, U2872, U2871, U2870, U2869, U2868, U2867, U2866, U2865, U2864, 
        U2863, U2862, U2861, U2860, U2859, U2858, U2857, U2856, U2855, U2854, 
        U2853, U2852, U2851, U2850, U2849, U2848, U2847, U2846, U2845, U2844, 
        U2843, U2842, U2841, U2840, U2839, U2838, U2837, U2836, U2835, U2834, 
        U2833, U2832, U2831, U2830, U2829, U2828, U2827, U2826, U2825, U2824, 
        U2823, U2822, U2821, U2820, U2819, U2818, U2817, U2816, U2815, U2814, 
        U2813, U2812, U2811, U2810, U2809, U2808, U2807, U2806, U2805, U2804, 
        U2803, U2802, U2801, U2800, U2799, U2798, U2797, U2796, U2795, U3468, 
        U2794, U3469, U3470, U2793, U3471, U2792, U3472, U2791, U3473, U2790, 
        U2789, U3474, U2788 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
         READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
         M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
         STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
         W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput0, keyinput1,
         keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7,
         keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13,
         keyinput14, keyinput15, keyinput16, keyinput17, keyinput18,
         keyinput19, keyinput20, keyinput21, keyinput22, keyinput23,
         keyinput24, keyinput25, keyinput26, keyinput27, keyinput28,
         keyinput29, keyinput30, keyinput31, keyinput32, keyinput33,
         keyinput34, keyinput35, keyinput36, keyinput37, keyinput38,
         keyinput39, keyinput40, keyinput41, keyinput42, keyinput43,
         keyinput44, keyinput45, keyinput46, keyinput47, keyinput48,
         keyinput49, keyinput50, keyinput51, keyinput52, keyinput53,
         keyinput54, keyinput55, keyinput56, keyinput57, keyinput58,
         keyinput59, keyinput60, keyinput61, keyinput62, keyinput63;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n2963, n2964, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973,
         n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983,
         n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993,
         n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003,
         n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013,
         n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023,
         n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033,
         n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043,
         n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053,
         n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063,
         n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073,
         n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083,
         n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093,
         n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103,
         n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113,
         n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123,
         n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133,
         n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143,
         n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153,
         n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163,
         n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173,
         n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183,
         n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193,
         n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203,
         n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213,
         n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223,
         n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233,
         n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243,
         n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253,
         n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263,
         n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273,
         n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283,
         n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293,
         n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303,
         n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313,
         n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323,
         n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333,
         n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343,
         n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353,
         n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363,
         n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373,
         n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383,
         n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393,
         n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403,
         n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413,
         n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423,
         n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433,
         n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443,
         n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453,
         n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463,
         n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473,
         n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483,
         n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493,
         n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503,
         n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513,
         n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523,
         n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533,
         n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543,
         n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553,
         n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563,
         n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573,
         n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583,
         n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593,
         n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603,
         n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613,
         n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623,
         n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633,
         n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643,
         n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653,
         n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663,
         n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673,
         n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683,
         n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693,
         n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703,
         n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713,
         n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723,
         n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733,
         n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743,
         n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753,
         n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763,
         n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773,
         n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783,
         n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793,
         n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803,
         n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813,
         n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823,
         n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833,
         n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843,
         n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853,
         n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863,
         n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873,
         n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883,
         n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893,
         n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903,
         n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913,
         n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923,
         n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933,
         n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943,
         n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953,
         n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963,
         n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973,
         n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983,
         n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993,
         n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003,
         n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013,
         n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023,
         n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033,
         n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043,
         n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053,
         n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063,
         n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073,
         n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083,
         n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093,
         n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103,
         n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113,
         n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123,
         n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133,
         n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143,
         n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153,
         n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163,
         n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173,
         n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183,
         n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193,
         n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203,
         n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213,
         n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223,
         n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233,
         n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243,
         n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253,
         n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263,
         n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273,
         n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283,
         n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293,
         n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303,
         n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313,
         n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323,
         n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333,
         n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343,
         n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353,
         n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363,
         n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373,
         n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383,
         n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393,
         n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403,
         n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413,
         n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423,
         n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433,
         n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443,
         n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453,
         n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463,
         n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473,
         n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483,
         n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493,
         n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503,
         n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513,
         n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523,
         n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533,
         n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543,
         n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553,
         n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563,
         n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573,
         n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583,
         n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593,
         n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603,
         n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613,
         n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623,
         n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633,
         n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643,
         n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653,
         n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663,
         n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673,
         n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683,
         n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693,
         n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703,
         n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713,
         n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723,
         n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733,
         n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743,
         n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753,
         n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763,
         n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773,
         n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783,
         n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793,
         n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803,
         n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813,
         n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823,
         n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833,
         n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843,
         n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853,
         n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863,
         n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873,
         n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883,
         n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893,
         n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903,
         n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913,
         n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923,
         n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933,
         n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943,
         n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953,
         n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963,
         n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973,
         n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983,
         n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993,
         n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003,
         n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013,
         n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023,
         n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033,
         n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043,
         n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053,
         n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063,
         n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073,
         n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083,
         n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093,
         n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103,
         n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113,
         n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123,
         n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133,
         n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143,
         n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153,
         n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163,
         n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173,
         n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183,
         n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193,
         n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203,
         n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213,
         n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223,
         n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233,
         n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243,
         n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253,
         n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263,
         n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273,
         n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283,
         n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293,
         n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303,
         n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313,
         n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323,
         n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333,
         n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343,
         n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353,
         n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363,
         n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373,
         n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383,
         n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393,
         n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403,
         n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413,
         n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423,
         n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433,
         n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443,
         n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453,
         n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463,
         n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473,
         n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483,
         n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493,
         n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503,
         n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513,
         n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523,
         n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533,
         n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543,
         n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553,
         n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563,
         n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573,
         n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583,
         n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593,
         n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603,
         n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613,
         n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623,
         n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633,
         n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643,
         n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653,
         n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663,
         n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673,
         n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683,
         n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693,
         n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703,
         n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713,
         n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723,
         n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733,
         n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743,
         n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753,
         n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763,
         n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773,
         n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783,
         n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793,
         n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803,
         n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813,
         n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823,
         n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833,
         n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843,
         n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853,
         n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863,
         n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873,
         n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883,
         n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893,
         n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903,
         n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913,
         n5914, n5915, n5916, n5917, n5919, n5920, n5921, n5922, n5923, n5924,
         n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934,
         n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944,
         n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954,
         n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964,
         n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974,
         n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984,
         n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994,
         n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004,
         n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014,
         n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024,
         n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034,
         n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044,
         n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054,
         n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064,
         n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074,
         n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084,
         n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094,
         n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104,
         n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114,
         n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124,
         n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134,
         n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144,
         n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154,
         n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164,
         n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174,
         n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184,
         n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194,
         n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204,
         n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214,
         n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224,
         n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234,
         n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244,
         n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254,
         n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264,
         n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274,
         n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284,
         n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294,
         n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304,
         n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314,
         n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324,
         n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334,
         n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344,
         n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354,
         n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364,
         n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374,
         n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384,
         n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394,
         n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404,
         n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414,
         n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424,
         n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434,
         n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444,
         n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454,
         n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464,
         n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474,
         n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484,
         n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494,
         n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504,
         n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514,
         n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524,
         n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534,
         n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544,
         n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554,
         n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564,
         n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574,
         n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584,
         n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594,
         n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604,
         n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614,
         n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624,
         n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634,
         n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644,
         n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654,
         n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664,
         n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672;

  INV_X1 U3412 ( .A(n5813), .ZN(n5868) );
  OR2_X1 U3413 ( .A1(n4695), .A2(n3682), .ZN(n3525) );
  CLKBUF_X2 U3414 ( .A(n4012), .Z(n4110) );
  AOI21_X1 U3415 ( .B1(n4344), .B2(n6382), .A(n3189), .ZN(n3243) );
  INV_X1 U3416 ( .A(n3432), .ZN(n3471) );
  CLKBUF_X2 U3417 ( .A(n3043), .Z(n3878) );
  CLKBUF_X2 U3418 ( .A(n3851), .Z(n3963) );
  CLKBUF_X2 U3419 ( .A(n3164), .Z(n3925) );
  AND2_X2 U3421 ( .A1(n3109), .A2(n4391), .ZN(n4192) );
  INV_X4 U3422 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n6382) );
  BUF_X1 U3423 ( .A(n4013), .Z(n4382) );
  AND4_X1 U3424 ( .A1(n3009), .A2(n3008), .A3(n3007), .A4(n3006), .ZN(n3015)
         );
  INV_X1 U3425 ( .A(n3109), .ZN(n5272) );
  AND2_X1 U3426 ( .A1(n5285), .A2(n4534), .ZN(n3210) );
  AND2_X1 U3427 ( .A1(n2990), .A2(n4509), .ZN(n3164) );
  BUF_X2 U3428 ( .A(n3037), .Z(n2963) );
  BUF_X2 U3429 ( .A(n3074), .Z(n3853) );
  AND4_X1 U3430 ( .A1(n3078), .A2(n3077), .A3(n3076), .A4(n3075), .ZN(n3094)
         );
  AOI22_X1 U3431 ( .A1(n3243), .A2(n3232), .B1(n3231), .B2(n3230), .ZN(n3233)
         );
  OR2_X1 U3432 ( .A1(n4333), .A2(n5301), .ZN(n4277) );
  AOI22_X1 U3433 ( .A1(n6605), .A2(keyinput2), .B1(n5187), .B2(keyinput58), 
        .ZN(n6604) );
  AOI22_X1 U3434 ( .A1(keyinput7), .A2(n6534), .B1(keyinput10), .B2(n6532), 
        .ZN(n6533) );
  NAND2_X1 U3435 ( .A1(n3234), .A2(n3233), .ZN(n3298) );
  NAND2_X1 U3436 ( .A1(n4217), .A2(n4220), .ZN(n5301) );
  NAND2_X1 U3437 ( .A1(n3097), .A2(n4013), .ZN(n4012) );
  OAI221_X1 U3438 ( .B1(n6605), .B2(keyinput2), .C1(n5187), .C2(keyinput58), 
        .A(n6604), .ZN(n6609) );
  OAI21_X1 U3439 ( .B1(n6534), .B2(keyinput7), .A(n6533), .ZN(n6547) );
  XNOR2_X1 U3440 ( .A(n3328), .B(n3326), .ZN(n3534) );
  OR2_X1 U3441 ( .A1(n3027), .A2(n3026), .ZN(n3496) );
  CLKBUF_X2 U3442 ( .A(n3097), .Z(n4391) );
  AND2_X1 U3443 ( .A1(n2968), .A2(n4081), .ZN(n5403) );
  XNOR2_X1 U3444 ( .A(n4113), .B(n4112), .ZN(n5356) );
  INV_X1 U34450 ( .A(n6047), .ZN(n6032) );
  AND2_X2 U34460 ( .A1(n2982), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n5285) );
  INV_X1 U34470 ( .A(n5838), .ZN(n5826) );
  AOI22_X1 U34480 ( .A1(n4175), .A2(n4174), .B1(n4173), .B2(n4172), .ZN(n5216)
         );
  AOI21_X1 U3449 ( .B1(n5431), .B2(n5515), .A(n4009), .ZN(n4010) );
  NAND2_X1 U34510 ( .A1(n3110), .A2(n3109), .ZN(n3438) );
  AOI21_X2 U34520 ( .B1(n5617), .B2(n5241), .A(n2969), .ZN(n5504) );
  MUX2_X2 U34530 ( .A(n3258), .B(n3257), .S(n3256), .Z(n4764) );
  NAND2_X1 U3454 ( .A1(n5244), .A2(n5243), .ZN(n5246) );
  OR2_X1 U34550 ( .A1(n5401), .A2(n5400), .ZN(n5705) );
  NOR2_X1 U34560 ( .A1(n5259), .A2(n5383), .ZN(n4097) );
  NAND2_X1 U3457 ( .A1(n4735), .A2(n4737), .ZN(n4809) );
  NOR2_X1 U3458 ( .A1(n6543), .A2(n5331), .ZN(n5328) );
  NAND2_X1 U34590 ( .A1(n3546), .A2(n3545), .ZN(n4611) );
  CLKBUF_X1 U34600 ( .A(n4972), .Z(n4993) );
  AND2_X1 U34610 ( .A1(n3495), .A2(n3997), .ZN(n3513) );
  AOI21_X1 U34620 ( .B1(n4317), .B2(n4316), .A(n3267), .ZN(n5966) );
  AND2_X2 U34640 ( .A1(n5770), .A2(n4001), .ZN(n5963) );
  NAND2_X2 U34650 ( .A1(n5427), .A2(n5271), .ZN(n5417) );
  NAND2_X1 U3466 ( .A1(n3147), .A2(n3176), .ZN(n3272) );
  AOI21_X1 U3467 ( .B1(n3154), .B2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(n3153), 
        .ZN(n3273) );
  NAND2_X1 U34680 ( .A1(n4030), .A2(n4029), .ZN(n4555) );
  NAND2_X1 U34690 ( .A1(n3120), .A2(n3389), .ZN(n4230) );
  OAI211_X1 U34700 ( .C1(n3471), .C2(n3221), .A(n3220), .B(n3219), .ZN(n3255)
         );
  INV_X1 U34710 ( .A(n4277), .ZN(n4214) );
  CLKBUF_X1 U34720 ( .A(n4116), .Z(n4218) );
  CLKBUF_X1 U34730 ( .A(n4277), .Z(n4504) );
  NAND2_X1 U34740 ( .A1(n3282), .A2(n3281), .ZN(n3485) );
  INV_X1 U3475 ( .A(n4110), .ZN(n4208) );
  NOR2_X1 U3477 ( .A1(n4382), .A2(n3123), .ZN(n3134) );
  AND2_X2 U3478 ( .A1(n3496), .A2(n4276), .ZN(n4221) );
  CLKBUF_X1 U3479 ( .A(n3496), .Z(n5271) );
  AND4_X1 U3480 ( .A1(n3082), .A2(n3081), .A3(n3080), .A4(n3079), .ZN(n3093)
         );
  AND4_X1 U3481 ( .A1(n3090), .A2(n3089), .A3(n3088), .A4(n3087), .ZN(n3091)
         );
  NOR2_X1 U3482 ( .A1(n2996), .A2(n2995), .ZN(n2997) );
  AND4_X1 U3483 ( .A1(n3013), .A2(n3012), .A3(n3011), .A4(n3010), .ZN(n3014)
         );
  BUF_X2 U3484 ( .A(n2963), .Z(n3852) );
  AND4_X1 U3485 ( .A1(n3086), .A2(n3085), .A3(n3084), .A4(n3083), .ZN(n3092)
         );
  BUF_X2 U3486 ( .A(n3205), .Z(n3965) );
  BUF_X2 U3487 ( .A(n3036), .Z(n3156) );
  INV_X2 U3488 ( .A(n5542), .ZN(n5515) );
  BUF_X2 U3489 ( .A(n3210), .Z(n3973) );
  BUF_X2 U3490 ( .A(n3283), .Z(n3197) );
  NAND2_X2 U3491 ( .A1(n4923), .A2(n6382), .ZN(n6047) );
  CLKBUF_X2 U3492 ( .A(n3037), .Z(n2964) );
  XNOR2_X2 U3493 ( .A(n4151), .B(n3999), .ZN(n5431) );
  AND2_X4 U3494 ( .A1(n4519), .A2(n5285), .ZN(n3283) );
  OAI21_X2 U3495 ( .B1(n4091), .B2(EBX_REG_1__SCAN_IN), .A(n4015), .ZN(n4018)
         );
  OAI21_X2 U3496 ( .B1(n5021), .B2(n5024), .A(n5022), .ZN(n5076) );
  OAI21_X2 U3497 ( .B1(n4964), .B2(n3401), .A(n2971), .ZN(n5021) );
  AND2_X4 U3499 ( .A1(n2988), .A2(n4509), .ZN(n2966) );
  AND2_X1 U3500 ( .A1(n4377), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3435) );
  AND2_X2 U3501 ( .A1(n3435), .A2(n4370), .ZN(n3432) );
  INV_X1 U3502 ( .A(n4023), .ZN(n4043) );
  AND2_X1 U3503 ( .A1(n4103), .A2(n4110), .ZN(n4219) );
  INV_X1 U3504 ( .A(n4043), .ZN(n4334) );
  NOR2_X1 U3505 ( .A1(n3097), .A2(n4131), .ZN(n3137) );
  NAND2_X1 U3506 ( .A1(n3351), .A2(n3350), .ZN(n3368) );
  OR2_X1 U3507 ( .A1(n3170), .A2(n3169), .ZN(n3238) );
  AOI22_X1 U3508 ( .A1(n2963), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3036), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3020) );
  NAND2_X1 U3509 ( .A1(n4413), .A2(n6382), .ZN(n3295) );
  CLKBUF_X1 U3510 ( .A(n3124), .Z(n4282) );
  INV_X1 U3511 ( .A(n5505), .ZN(n5243) );
  INV_X1 U3512 ( .A(n5504), .ZN(n5244) );
  OAI211_X1 U3513 ( .C1(n3471), .C2(n3229), .A(n3228), .B(n3227), .ZN(n3245)
         );
  AND2_X1 U3514 ( .A1(n4493), .A2(n4236), .ZN(n5289) );
  AOI22_X1 U3515 ( .A1(n3037), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3036), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3031) );
  AOI22_X1 U3516 ( .A1(n3205), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3964), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3030) );
  INV_X1 U3517 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n6571) );
  AND4_X1 U3518 ( .A1(n3005), .A2(n3004), .A3(n3003), .A4(n3002), .ZN(n3016)
         );
  AND2_X1 U3519 ( .A1(n3422), .A2(n5083), .ZN(n3408) );
  NOR2_X2 U3520 ( .A1(n5073), .A2(n5058), .ZN(n5118) );
  NOR2_X2 U3521 ( .A1(n4555), .A2(n4554), .ZN(n4610) );
  AOI21_X1 U3522 ( .B1(n4107), .B2(n4022), .A(n4021), .ZN(n4480) );
  NAND2_X1 U3523 ( .A1(n4028), .A2(n4027), .ZN(n4479) );
  AND2_X1 U3524 ( .A1(n4026), .A2(n4025), .ZN(n4027) );
  NAND2_X1 U3525 ( .A1(n3483), .A2(n3482), .ZN(n3487) );
  INV_X1 U3526 ( .A(n6165), .ZN(n4701) );
  INV_X1 U3527 ( .A(n4165), .ZN(n4166) );
  AND2_X1 U3528 ( .A1(n4334), .A2(n4127), .ZN(n5866) );
  AND2_X1 U3529 ( .A1(n5016), .A2(STATE2_REG_3__SCAN_IN), .ZN(n5870) );
  INV_X1 U3530 ( .A(n5646), .ZN(n5438) );
  XNOR2_X1 U3531 ( .A(n4181), .B(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5172)
         );
  OR2_X1 U3532 ( .A1(n5644), .A2(n6024), .ZN(n4263) );
  AND2_X1 U3533 ( .A1(n4245), .A2(n4206), .ZN(n6050) );
  AND2_X1 U3534 ( .A1(n3124), .A2(n4370), .ZN(n3114) );
  NAND2_X1 U3535 ( .A1(n3109), .A2(n3494), .ZN(n3124) );
  CLKBUF_X2 U3536 ( .A(n3163), .Z(n3966) );
  NOR2_X1 U3537 ( .A1(n4217), .A2(n4220), .ZN(n4023) );
  XNOR2_X1 U3538 ( .A(n3174), .B(n3173), .ZN(n3234) );
  NAND2_X1 U3539 ( .A1(n3073), .A2(n3072), .ZN(n3126) );
  NAND2_X1 U3540 ( .A1(n3155), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3282) );
  NAND2_X1 U3541 ( .A1(n3432), .A2(n4192), .ZN(n3463) );
  INV_X1 U3542 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n2983) );
  NAND4_X1 U3543 ( .A1(n3134), .A2(n4221), .A3(n3073), .A4(n4363), .ZN(n4116)
         );
  INV_X1 U3544 ( .A(n4808), .ZN(n3585) );
  INV_X1 U3545 ( .A(n4809), .ZN(n3586) );
  AND2_X1 U3546 ( .A1(n4747), .A2(n4746), .ZN(n4735) );
  INV_X1 U3547 ( .A(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3526) );
  NAND2_X1 U3548 ( .A1(n3517), .A2(n3516), .ZN(n4326) );
  OR2_X1 U3549 ( .A1(n5237), .A2(n5520), .ZN(n5483) );
  INV_X1 U3550 ( .A(n3367), .ZN(n3365) );
  INV_X1 U3551 ( .A(n3368), .ZN(n3366) );
  INV_X1 U3552 ( .A(n3282), .ZN(n3226) );
  CLKBUF_X1 U3553 ( .A(n4183), .Z(n4184) );
  NAND2_X1 U3554 ( .A1(n3280), .A2(n3279), .ZN(n4346) );
  AND2_X2 U3555 ( .A1(n4503), .A2(n4519), .ZN(n3163) );
  INV_X1 U3556 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4864) );
  CLKBUF_X1 U3557 ( .A(n4114), .Z(n4115) );
  INV_X1 U3558 ( .A(n4116), .ZN(n5292) );
  INV_X1 U3559 ( .A(n5330), .ZN(n5853) );
  OR2_X1 U3560 ( .A1(n3148), .A2(n5288), .ZN(n3141) );
  NOR2_X1 U3561 ( .A1(n4157), .A2(n4955), .ZN(n4128) );
  INV_X1 U3562 ( .A(n5336), .ZN(n4073) );
  NAND2_X1 U3563 ( .A1(n3538), .A2(n3537), .ZN(n4560) );
  INV_X1 U3564 ( .A(n5920), .ZN(n4288) );
  OR3_X2 U3565 ( .A1(n5302), .A2(n4115), .A3(n6369), .ZN(n4392) );
  CLKBUF_X1 U3566 ( .A(n3239), .Z(n4394) );
  NOR2_X1 U3567 ( .A1(n3936), .A2(n5309), .ZN(n3937) );
  CLKBUF_X1 U3568 ( .A(n5227), .Z(n5228) );
  AND2_X1 U3569 ( .A1(n5425), .A2(n5229), .ZN(n5373) );
  INV_X1 U3570 ( .A(n3808), .ZN(n3797) );
  NAND2_X1 U3571 ( .A1(n3898), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n3808)
         );
  AND2_X1 U3572 ( .A1(n3892), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n3898)
         );
  AND2_X1 U3573 ( .A1(n5425), .A2(n5253), .ZN(n5381) );
  AND2_X1 U3574 ( .A1(n5425), .A2(n5313), .ZN(n5393) );
  AND2_X1 U3575 ( .A1(PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n3796), .ZN(n3848)
         );
  INV_X1 U3576 ( .A(n3870), .ZN(n3796) );
  NOR2_X1 U3577 ( .A1(n3730), .A2(n5534), .ZN(n3731) );
  NAND2_X1 U3578 ( .A1(n3731), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n3870)
         );
  CLKBUF_X1 U3579 ( .A(n5129), .Z(n5423) );
  NOR2_X1 U3580 ( .A1(n6605), .A2(n3666), .ZN(n3713) );
  INV_X1 U3581 ( .A(n5034), .ZN(n3648) );
  AND2_X1 U3582 ( .A1(n3422), .A2(n5988), .ZN(n3401) );
  NOR2_X1 U3583 ( .A1(n3422), .A2(n3402), .ZN(n5024) );
  NOR2_X1 U3584 ( .A1(n4984), .A2(n4985), .ZN(n4983) );
  NAND2_X1 U3585 ( .A1(n4937), .A2(n4936), .ZN(n4984) );
  NOR2_X1 U3586 ( .A1(n6534), .A2(n3588), .ZN(n3618) );
  NOR2_X2 U3587 ( .A1(n4807), .A2(n4918), .ZN(n4937) );
  NOR2_X1 U3588 ( .A1(n6636), .A2(n3554), .ZN(n3587) );
  CLKBUF_X1 U3589 ( .A(n4807), .Z(n4919) );
  NOR2_X1 U3590 ( .A1(n6571), .A2(n3540), .ZN(n3549) );
  NAND2_X1 U3591 ( .A1(n3549), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3554)
         );
  NOR2_X2 U3592 ( .A1(n4612), .A2(n3547), .ZN(n4747) );
  NAND2_X1 U3593 ( .A1(n4560), .A2(n4611), .ZN(n3547) );
  NOR2_X1 U3594 ( .A1(n3527), .A2(n3526), .ZN(n3541) );
  INV_X1 U3595 ( .A(n3519), .ZN(n3520) );
  NAND2_X1 U3596 ( .A1(n3520), .A2(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3527)
         );
  NAND2_X1 U3597 ( .A1(PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n3519) );
  NAND2_X1 U3598 ( .A1(n3513), .A2(n4298), .ZN(n4328) );
  INV_X1 U3599 ( .A(n4178), .ZN(n5457) );
  OR2_X1 U3600 ( .A1(n3419), .A2(n3426), .ZN(n3420) );
  CLKBUF_X1 U3601 ( .A(n5259), .Z(n5382) );
  NOR2_X2 U3602 ( .A1(n5395), .A2(n5318), .ZN(n5317) );
  NOR2_X1 U3603 ( .A1(n3422), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5494)
         );
  INV_X1 U3604 ( .A(n5246), .ZN(n5503) );
  XNOR2_X1 U3606 ( .A(n3422), .B(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5075)
         );
  NAND2_X1 U3607 ( .A1(n4060), .A2(n4059), .ZN(n5071) );
  INV_X1 U3608 ( .A(n4987), .ZN(n4060) );
  NOR2_X2 U3609 ( .A1(n4939), .A2(n4940), .ZN(n4989) );
  OR2_X1 U3610 ( .A1(n3422), .A2(n3399), .ZN(n4963) );
  OR2_X1 U3611 ( .A1(n3422), .A2(n5997), .ZN(n4912) );
  INV_X1 U3612 ( .A(n4481), .ZN(n4030) );
  NAND2_X1 U3613 ( .A1(n5013), .A2(n4334), .ZN(n4318) );
  CLKBUF_X1 U3614 ( .A(n3502), .Z(n3503) );
  XNOR2_X1 U3615 ( .A(n3248), .B(n3247), .ZN(n4343) );
  XNOR2_X1 U3616 ( .A(n3246), .B(n3245), .ZN(n3247) );
  BUF_X1 U3617 ( .A(n3244), .Z(n3246) );
  CLKBUF_X1 U3618 ( .A(n3493), .Z(n4694) );
  OR3_X1 U3619 ( .A1(n4497), .A2(n4496), .A3(n4495), .ZN(n6349) );
  AND2_X1 U3620 ( .A1(n4758), .A2(n6197), .ZN(n4760) );
  OR2_X1 U3621 ( .A1(n6057), .A2(n5627), .ZN(n4765) );
  AND2_X1 U3622 ( .A1(n5627), .A2(n6232), .ZN(n6118) );
  INV_X1 U3623 ( .A(n4352), .ZN(n6119) );
  OR2_X1 U3624 ( .A1(n4695), .A2(n5631), .ZN(n6191) );
  CLKBUF_X1 U3625 ( .A(n4413), .Z(n6237) );
  INV_X1 U3626 ( .A(n4764), .ZN(n6232) );
  INV_X1 U3627 ( .A(n5428), .ZN(n5415) );
  AND2_X1 U3628 ( .A1(n5435), .A2(n5273), .ZN(n5885) );
  AND2_X1 U3629 ( .A1(n5435), .A2(n4284), .ZN(n5060) );
  CLKBUF_X1 U3630 ( .A(n4463), .Z(n6668) );
  INV_X1 U3631 ( .A(n5928), .ZN(n5936) );
  AND2_X1 U3632 ( .A1(n5175), .A2(n5174), .ZN(n5646) );
  OAI21_X1 U3633 ( .B1(n5381), .B2(n5380), .A(n5379), .ZN(n5673) );
  INV_X1 U3634 ( .A(n5732), .ZN(n5878) );
  OR2_X1 U3635 ( .A1(n5963), .A2(n4304), .ZN(n5973) );
  XNOR2_X1 U3636 ( .A(n3430), .B(n6623), .ZN(n5201) );
  AOI21_X1 U3637 ( .B1(n5185), .B2(INSTADDRPOINTER_REG_30__SCAN_IN), .A(n3429), 
        .ZN(n3430) );
  OR2_X1 U3638 ( .A1(n5572), .A2(n4259), .ZN(n5564) );
  XNOR2_X1 U3639 ( .A(n5251), .B(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5269)
         );
  NAND2_X1 U3640 ( .A1(n5250), .A2(n5249), .ZN(n5251) );
  NAND2_X1 U3641 ( .A1(n5248), .A2(n5247), .ZN(n5249) );
  OR2_X1 U3642 ( .A1(n5741), .A2(n4256), .ZN(n5602) );
  CLKBUF_X1 U3643 ( .A(n5138), .Z(n5140) );
  AND2_X1 U3644 ( .A1(n5984), .A2(n5159), .ZN(n5742) );
  INV_X1 U3645 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6635) );
  CLKBUF_X1 U3647 ( .A(n4345), .Z(n5632) );
  INV_X1 U3648 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n5288) );
  INV_X1 U3649 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n2982) );
  OR2_X1 U3650 ( .A1(n5302), .A2(n6470), .ZN(n5637) );
  INV_X1 U3651 ( .A(n6117), .ZN(n6081) );
  OR4_X1 U3652 ( .A1(n6095), .A2(n6156), .A3(n6094), .A4(n6093), .ZN(n6114) );
  INV_X1 U3653 ( .A(n4663), .ZN(n4688) );
  INV_X1 U3654 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n6391) );
  AND2_X1 U3655 ( .A1(n6375), .A2(n6374), .ZN(n6467) );
  NOR3_X1 U3656 ( .A1(n4168), .A2(n4167), .A3(n4166), .ZN(n4176) );
  OR2_X1 U3657 ( .A1(n5276), .A2(n5826), .ZN(n4177) );
  AND2_X1 U3658 ( .A1(n4263), .A2(n4262), .ZN(n4264) );
  NAND2_X4 U3659 ( .A1(n3391), .A2(n3390), .ZN(n3422) );
  AND2_X2 U3660 ( .A1(n4534), .A2(n4509), .ZN(n3198) );
  NOR2_X1 U3661 ( .A1(n4480), .A2(n4479), .ZN(n4029) );
  AND4_X1 U3662 ( .A1(n2987), .A2(n2986), .A3(n2985), .A4(n2984), .ZN(n2967)
         );
  AND2_X1 U3663 ( .A1(n5131), .A2(n4073), .ZN(n2968) );
  INV_X1 U3664 ( .A(n4220), .ZN(n3123) );
  INV_X1 U3665 ( .A(n4983), .ZN(n5035) );
  NAND2_X1 U3666 ( .A1(n5482), .A2(n2973), .ZN(n2969) );
  AND2_X1 U3667 ( .A1(n5379), .A2(n5372), .ZN(n2970) );
  AND2_X1 U3668 ( .A1(n4963), .A2(n3400), .ZN(n2971) );
  AND4_X1 U3669 ( .A1(n3055), .A2(n3054), .A3(n3053), .A4(n3052), .ZN(n2972)
         );
  NAND2_X1 U3670 ( .A1(n3422), .A2(n5510), .ZN(n2973) );
  NOR2_X1 U3671 ( .A1(n3425), .A2(n3419), .ZN(n2974) );
  OR2_X1 U3672 ( .A1(n3403), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n2975)
         );
  AND3_X1 U3673 ( .A1(n3058), .A2(n3057), .A3(n3056), .ZN(n2976) );
  AND2_X1 U3674 ( .A1(n4740), .A2(n4741), .ZN(n4739) );
  OR2_X1 U3675 ( .A1(n4309), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n2977)
         );
  INV_X1 U3676 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3117) );
  OR2_X1 U3677 ( .A1(n5366), .A2(n4207), .ZN(n2978) );
  OR2_X1 U3678 ( .A1(n5216), .A2(n5863), .ZN(n2979) );
  AND4_X1 U3679 ( .A1(n3128), .A2(n4527), .A3(n3127), .A4(n4506), .ZN(n2980)
         );
  INV_X1 U3680 ( .A(n3297), .ZN(n4417) );
  INV_X1 U3681 ( .A(n3143), .ZN(n3140) );
  INV_X1 U3682 ( .A(n3422), .ZN(n3403) );
  NOR2_X1 U3683 ( .A1(n3102), .A2(n3135), .ZN(n3099) );
  CLKBUF_X1 U3684 ( .A(n3038), .Z(n3944) );
  NAND2_X1 U3685 ( .A1(n3104), .A2(n3050), .ZN(n3112) );
  INV_X1 U3686 ( .A(n3326), .ZN(n3327) );
  AND2_X1 U3687 ( .A1(n6635), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3449)
         );
  BUF_X1 U3688 ( .A(n3051), .Z(n3162) );
  NOR2_X2 U3689 ( .A1(n3328), .A2(n3327), .ZN(n3351) );
  NAND2_X1 U3690 ( .A1(n3223), .A2(n3222), .ZN(n3244) );
  NAND2_X1 U3691 ( .A1(n3403), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n3400) );
  XNOR2_X1 U3692 ( .A(n3391), .B(n3379), .ZN(n3548) );
  OR2_X1 U3693 ( .A1(n3316), .A2(n3315), .ZN(n3342) );
  INV_X1 U3694 ( .A(n4565), .ZN(n4038) );
  AND2_X1 U3695 ( .A1(n3364), .A2(n3363), .ZN(n3367) );
  OR2_X1 U3696 ( .A1(n3188), .A2(n3187), .ZN(n3249) );
  NAND2_X1 U3697 ( .A1(n3295), .A2(n3294), .ZN(n3297) );
  NAND3_X1 U3698 ( .A1(n4230), .A2(n2980), .A3(n3130), .ZN(n3190) );
  AOI22_X1 U3699 ( .A1(n3858), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3043), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3018) );
  AND4_X1 U3700 ( .A1(n3001), .A2(n3000), .A3(n2999), .A4(n2998), .ZN(n3017)
         );
  INV_X1 U3701 ( .A(n3463), .ZN(n3481) );
  OR2_X1 U3702 ( .A1(n3992), .A2(n3991), .ZN(n4004) );
  NOR2_X1 U3703 ( .A1(n3847), .A2(n5702), .ZN(n3890) );
  NAND2_X1 U3704 ( .A1(n3548), .A2(n3662), .ZN(n3553) );
  AND2_X1 U3705 ( .A1(n3416), .A2(n5527), .ZN(n5481) );
  OR2_X1 U3706 ( .A1(n3422), .A2(n5083), .ZN(n3407) );
  NAND2_X1 U3707 ( .A1(n3366), .A2(n3365), .ZN(n3391) );
  INV_X1 U3708 ( .A(n4020), .ZN(n4021) );
  OR2_X1 U3709 ( .A1(n3204), .A2(n3203), .ZN(n3237) );
  OR2_X1 U3710 ( .A1(n3216), .A2(n3215), .ZN(n3392) );
  INV_X1 U3711 ( .A(n3135), .ZN(n3121) );
  NOR2_X1 U3712 ( .A1(n5649), .A2(n6458), .ZN(n4164) );
  INV_X1 U3713 ( .A(n5695), .ZN(n4135) );
  INV_X1 U3714 ( .A(n5040), .ZN(n4059) );
  AND2_X1 U3715 ( .A1(n4023), .A2(n4110), .ZN(n4100) );
  AND2_X1 U3716 ( .A1(PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n3797), .ZN(n3913)
         );
  AND2_X1 U3717 ( .A1(n3890), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n3892)
         );
  OR2_X1 U3718 ( .A1(n3633), .A2(n5808), .ZN(n3650) );
  NAND2_X1 U3719 ( .A1(n3553), .A2(n3552), .ZN(n4746) );
  AND2_X1 U3720 ( .A1(n5517), .A2(n3412), .ZN(n5472) );
  INV_X1 U3721 ( .A(n4091), .ZN(n4107) );
  NAND2_X1 U3722 ( .A1(n3272), .A2(n3274), .ZN(n4486) );
  XNOR2_X1 U3723 ( .A(n4486), .B(n4346), .ZN(n4413) );
  AND2_X1 U3725 ( .A1(n4354), .A2(n4353), .ZN(n4383) );
  AND2_X1 U3726 ( .A1(n4217), .A2(n3123), .ZN(n3239) );
  AND2_X1 U3727 ( .A1(n6384), .A2(n6382), .ZN(n4000) );
  AND2_X1 U3728 ( .A1(n4144), .A2(n4143), .ZN(n4145) );
  NAND2_X1 U3729 ( .A1(n5704), .A2(n4135), .ZN(n5315) );
  INV_X1 U3730 ( .A(n5870), .ZN(n5834) );
  NAND2_X1 U3731 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n5016), .ZN(n4955) );
  OR2_X1 U3732 ( .A1(n5407), .A2(n5408), .ZN(n5405) );
  AND2_X1 U3733 ( .A1(n5326), .A2(n3917), .ZN(n5227) );
  INV_X1 U3734 ( .A(n4334), .ZN(n4202) );
  NAND2_X1 U3735 ( .A1(n3913), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n3936)
         );
  NAND2_X1 U3736 ( .A1(n3848), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n3847)
         );
  AND2_X1 U3737 ( .A1(n5129), .A2(n5422), .ZN(n5326) );
  NOR2_X1 U3738 ( .A1(n3650), .A2(n3649), .ZN(n3665) );
  NAND2_X1 U3739 ( .A1(n3586), .A2(n3585), .ZN(n4807) );
  AOI21_X1 U3740 ( .B1(n3534), .B2(n3662), .A(n3533), .ZN(n4553) );
  NAND2_X1 U3741 ( .A1(n4111), .A2(n4174), .ZN(n4113) );
  AND3_X1 U3742 ( .A1(n5211), .A2(n3403), .A3(n5210), .ZN(n5456) );
  OR2_X1 U3743 ( .A1(n5496), .A2(n5245), .ZN(n5250) );
  INV_X1 U3744 ( .A(n5131), .ZN(n5419) );
  CLKBUF_X1 U3745 ( .A(n4740), .Z(n4753) );
  AND2_X1 U3746 ( .A1(n4198), .A2(n6383), .ZN(n4245) );
  NAND2_X1 U3748 ( .A1(n5292), .A2(n4217), .ZN(n4505) );
  BUF_X1 U3749 ( .A(n3518), .Z(n4695) );
  INV_X1 U3750 ( .A(n4696), .ZN(n4729) );
  INV_X1 U3751 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n4699) );
  NAND2_X1 U3752 ( .A1(n4392), .A2(n4266), .ZN(n6490) );
  NAND2_X1 U3753 ( .A1(n4146), .A2(n4145), .ZN(n4147) );
  NOR2_X1 U3754 ( .A1(n6436), .A2(n5062), .ZN(n5342) );
  NOR2_X1 U3755 ( .A1(n5818), .A2(n4134), .ZN(n5807) );
  AND2_X1 U3756 ( .A1(n5016), .A2(n4148), .ZN(n5838) );
  AND2_X1 U3757 ( .A1(n5016), .A2(n4155), .ZN(n5813) );
  AND2_X1 U3758 ( .A1(n5425), .A2(n5390), .ZN(n5400) );
  INV_X1 U3759 ( .A(n4219), .ZN(n4309) );
  BUF_X1 U3760 ( .A(n3123), .Z(n4377) );
  NAND2_X1 U3761 ( .A1(n3487), .A2(n3486), .ZN(n5302) );
  INV_X1 U3762 ( .A(n5497), .ZN(n5719) );
  AND2_X1 U3763 ( .A1(n4983), .A2(n3648), .ZN(n5050) );
  NAND2_X1 U3764 ( .A1(n3541), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3540)
         );
  NAND2_X1 U3765 ( .A1(n5246), .A2(n2975), .ZN(n5496) );
  AND2_X1 U3766 ( .A1(n5484), .A2(n5483), .ZN(n5512) );
  AND2_X1 U3767 ( .A1(n4245), .A2(n4216), .ZN(n6044) );
  AND2_X1 U3768 ( .A1(n5627), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6192) );
  INV_X1 U3769 ( .A(n4909), .ZN(n4866) );
  INV_X1 U3770 ( .A(n6087), .ZN(n6072) );
  INV_X1 U3771 ( .A(n6096), .ZN(n6113) );
  AND2_X1 U3772 ( .A1(n4356), .A2(n6232), .ZN(n4619) );
  INV_X1 U3773 ( .A(n6154), .ZN(n6144) );
  OR2_X1 U3774 ( .A1(n6167), .A2(n6166), .ZN(n6185) );
  AND2_X1 U3775 ( .A1(n4588), .A2(n4764), .ZN(n6184) );
  OR2_X1 U3776 ( .A1(n6241), .A2(n6240), .ZN(n6272) );
  NOR2_X1 U3777 ( .A1(n6233), .A2(n4764), .ZN(n6335) );
  NOR2_X1 U3778 ( .A1(n4421), .A2(n4865), .ZN(n4663) );
  NAND2_X1 U3779 ( .A1(n5431), .A2(n5838), .ZN(n4149) );
  INV_X1 U3780 ( .A(n5866), .ZN(n5863) );
  OR2_X1 U3781 ( .A1(n5393), .A2(n5392), .ZN(n5497) );
  NAND2_X1 U3782 ( .A1(n4338), .A2(n4337), .ZN(n5427) );
  OR2_X1 U3783 ( .A1(n2970), .A2(n5373), .ZN(n5467) );
  NAND2_X1 U3784 ( .A1(n4281), .A2(n4280), .ZN(n5435) );
  NOR2_X1 U3785 ( .A1(n6493), .A2(n4288), .ZN(n5888) );
  OR3_X1 U3786 ( .A1(n5302), .A2(n4287), .A3(n4286), .ZN(n5920) );
  OR3_X1 U3787 ( .A1(n5302), .A2(n4490), .A3(n4278), .ZN(n5928) );
  INV_X1 U3788 ( .A(n6667), .ZN(n4470) );
  OR2_X1 U3789 ( .A1(n5228), .A2(n5231), .ZN(n5443) );
  OR2_X1 U3790 ( .A1(n6363), .A2(n6369), .ZN(n5770) );
  INV_X1 U3791 ( .A(n6044), .ZN(n6024) );
  INV_X1 U3792 ( .A(n6050), .ZN(n6023) );
  INV_X1 U3793 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6358) );
  OR2_X1 U3794 ( .A1(n4765), .A2(n6232), .ZN(n4785) );
  OR2_X1 U3795 ( .A1(n4765), .A2(n4764), .ZN(n4909) );
  OR2_X1 U3796 ( .A1(n6057), .A2(n6190), .ZN(n6117) );
  INV_X1 U3797 ( .A(n4619), .ZN(n4653) );
  NAND2_X1 U3798 ( .A1(n6119), .A2(n6118), .ZN(n6188) );
  OR2_X1 U3799 ( .A1(n6191), .A2(n4865), .ZN(n6226) );
  OR2_X1 U3800 ( .A1(n6191), .A2(n6190), .ZN(n6275) );
  INV_X1 U3801 ( .A(n6335), .ZN(n4693) );
  NAND2_X1 U3802 ( .A1(n4150), .A2(n4149), .ZN(U2796) );
  INV_X1 U3803 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n2981) );
  AND2_X2 U3804 ( .A1(n2981), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n2989)
         );
  AND2_X2 U3805 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4534) );
  AND2_X2 U3806 ( .A1(n2989), .A2(n4534), .ZN(n3051) );
  BUF_X8 U3807 ( .A(n3051), .Z(n3971) );
  NOR2_X4 U3808 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4503) );
  AND2_X2 U3809 ( .A1(n4503), .A2(n4534), .ZN(n3074) );
  BUF_X4 U3810 ( .A(n3074), .Z(n3972) );
  AOI22_X1 U3811 ( .A1(n3971), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3972), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n2987) );
  INV_X1 U3812 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3510) );
  AND2_X2 U3813 ( .A1(n3510), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4519)
         );
  AND2_X4 U3814 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4509) );
  AND2_X2 U3815 ( .A1(n4519), .A2(n4509), .ZN(n3851) );
  NOR2_X4 U3816 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n2988) );
  AND2_X2 U3817 ( .A1(n5285), .A2(n2988), .ZN(n3037) );
  AOI22_X1 U3818 ( .A1(n3851), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n2963), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n2986) );
  NOR2_X2 U3819 ( .A1(n2983), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n2990)
         );
  AND2_X2 U3820 ( .A1(n2989), .A2(n2990), .ZN(n3061) );
  AOI22_X1 U3821 ( .A1(n3061), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3043), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n2985) );
  AND2_X2 U3822 ( .A1(n5285), .A2(n2990), .ZN(n3964) );
  AND2_X4 U3823 ( .A1(n2988), .A2(n4509), .ZN(n3157) );
  AOI22_X1 U3824 ( .A1(n3964), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3157), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n2984) );
  AND2_X2 U3825 ( .A1(n2989), .A2(n2988), .ZN(n3036) );
  AND2_X2 U3826 ( .A1(n2990), .A2(n4503), .ZN(n3038) );
  AOI22_X1 U3827 ( .A1(n3036), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n3038), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n2993) );
  AND2_X2 U3828 ( .A1(n4519), .A2(n2989), .ZN(n3205) );
  AOI22_X1 U3829 ( .A1(n3205), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3198), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n2992) );
  AOI22_X1 U3830 ( .A1(n3210), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3164), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n2991) );
  NAND3_X1 U3831 ( .A1(n2993), .A2(n2992), .A3(n2991), .ZN(n2996) );
  AOI22_X1 U3832 ( .A1(n3283), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3163), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n2994) );
  INV_X1 U3833 ( .A(n2994), .ZN(n2995) );
  NAND2_X2 U3834 ( .A1(n2967), .A2(n2997), .ZN(n3097) );
  NAND2_X1 U3835 ( .A1(n2963), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3001) );
  NAND2_X1 U3836 ( .A1(n3205), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3000) );
  NAND2_X1 U3837 ( .A1(n3964), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n2999) );
  NAND2_X1 U3838 ( .A1(n2966), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n2998) );
  NAND2_X1 U3839 ( .A1(n3061), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3005) );
  NAND2_X1 U3840 ( .A1(n3162), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3004)
         );
  NAND2_X1 U3841 ( .A1(n3074), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3003)
         );
  NAND2_X1 U3842 ( .A1(n3043), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3002) );
  NAND2_X1 U3843 ( .A1(n3851), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3009)
         );
  NAND2_X1 U3844 ( .A1(n3036), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3008) );
  BUF_X4 U3845 ( .A(n3038), .Z(n3858) );
  NAND2_X1 U3846 ( .A1(n3858), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3007) );
  NAND2_X1 U3847 ( .A1(n3198), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3006)
         );
  NAND2_X1 U3848 ( .A1(n3210), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3013)
         );
  NAND2_X1 U3849 ( .A1(n3283), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3012)
         );
  NAND2_X1 U3850 ( .A1(n3163), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3011) );
  NAND2_X1 U3851 ( .A1(n3164), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3010) );
  AND4_X4 U3852 ( .A1(n3017), .A2(n3016), .A3(n3015), .A4(n3014), .ZN(n4220)
         );
  AOI22_X1 U3853 ( .A1(n3163), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3061), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3021) );
  AOI22_X1 U3854 ( .A1(n3164), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3074), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3019) );
  NAND4_X1 U3855 ( .A1(n3021), .A2(n3020), .A3(n3019), .A4(n3018), .ZN(n3027)
         );
  AOI22_X1 U3856 ( .A1(n3210), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3051), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3025) );
  AOI22_X1 U3857 ( .A1(n3283), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3851), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3024) );
  AOI22_X1 U3858 ( .A1(n3205), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3964), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3023) );
  AOI22_X1 U3859 ( .A1(n2966), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n3198), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3022) );
  NAND4_X1 U3860 ( .A1(n3025), .A2(n3024), .A3(n3023), .A4(n3022), .ZN(n3026)
         );
  AOI22_X1 U3861 ( .A1(n3851), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3038), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3029) );
  AOI22_X1 U3862 ( .A1(n3157), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n3198), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3028) );
  NAND4_X1 U3863 ( .A1(n3031), .A2(n3030), .A3(n3029), .A4(n3028), .ZN(n3101)
         );
  AOI22_X1 U3864 ( .A1(n3210), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3051), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3035) );
  AOI22_X1 U3865 ( .A1(n3163), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3061), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3034) );
  AOI22_X1 U3866 ( .A1(n3164), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3074), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3033) );
  AOI22_X1 U3867 ( .A1(n3283), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3043), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3032) );
  NAND4_X1 U3868 ( .A1(n3035), .A2(n3034), .A3(n3033), .A4(n3032), .ZN(n3100)
         );
  NOR2_X2 U3869 ( .A1(n3101), .A2(n3100), .ZN(n3494) );
  NAND2_X1 U3870 ( .A1(n3496), .A2(n3494), .ZN(n3104) );
  AOI22_X1 U3871 ( .A1(n3037), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3036), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3042) );
  AOI22_X1 U3872 ( .A1(n3205), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3964), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3041) );
  AOI22_X1 U3873 ( .A1(n3851), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3038), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3040) );
  AOI22_X1 U3874 ( .A1(n2966), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n3198), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3039) );
  NAND4_X1 U3875 ( .A1(n3042), .A2(n3041), .A3(n3040), .A4(n3039), .ZN(n3049)
         );
  AOI22_X1 U3876 ( .A1(n3163), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3061), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3047) );
  AOI22_X1 U3877 ( .A1(n3210), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3051), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3046) );
  AOI22_X1 U3878 ( .A1(n3164), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3074), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3045) );
  AOI22_X1 U3879 ( .A1(n3283), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3043), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3044) );
  NAND4_X1 U3880 ( .A1(n3047), .A2(n3046), .A3(n3045), .A4(n3044), .ZN(n3048)
         );
  OR2_X4 U3881 ( .A1(n3049), .A2(n3048), .ZN(n3109) );
  NAND2_X1 U3882 ( .A1(n3496), .A2(n3109), .ZN(n3050) );
  AOI22_X1 U3883 ( .A1(n3858), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n3043), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3055) );
  AOI22_X1 U3884 ( .A1(n3210), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3164), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3054) );
  AOI22_X1 U3885 ( .A1(n3283), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3051), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3053) );
  AOI22_X1 U3886 ( .A1(n3036), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n3157), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3052) );
  AOI22_X1 U3887 ( .A1(n3205), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3964), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3058) );
  AOI22_X1 U3888 ( .A1(n2964), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n3198), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3057) );
  AOI22_X1 U3889 ( .A1(n3163), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3972), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3056) );
  AOI22_X1 U3890 ( .A1(n3851), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3061), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3059) );
  NAND3_X2 U3891 ( .A1(n2972), .A2(n2976), .A3(n3059), .ZN(n3102) );
  BUF_X2 U3892 ( .A(n3102), .Z(n4370) );
  NAND2_X1 U3894 ( .A1(n3112), .A2(n3155), .ZN(n4191) );
  INV_X1 U3895 ( .A(STATE_REG_1__SCAN_IN), .ZN(n6572) );
  INV_X1 U3896 ( .A(STATE_REG_2__SCAN_IN), .ZN(n6584) );
  NOR2_X1 U3897 ( .A1(n6572), .A2(n6584), .ZN(n6398) );
  NOR2_X1 U3898 ( .A1(STATE_REG_1__SCAN_IN), .A2(STATE_REG_2__SCAN_IN), .ZN(
        n3060) );
  NOR2_X1 U3899 ( .A1(n6398), .A2(n3060), .ZN(n4131) );
  INV_X1 U3900 ( .A(n3102), .ZN(n3110) );
  INV_X1 U3901 ( .A(n3438), .ZN(n3073) );
  AOI22_X1 U3902 ( .A1(n3851), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n2963), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3065) );
  AOI22_X1 U3903 ( .A1(n3283), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3061), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3064) );
  AOI22_X1 U3904 ( .A1(n3163), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3210), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3063) );
  AOI22_X1 U3905 ( .A1(n3164), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3972), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3062) );
  NAND4_X1 U3906 ( .A1(n3065), .A2(n3064), .A3(n3063), .A4(n3062), .ZN(n3071)
         );
  AOI22_X1 U3907 ( .A1(n3162), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3043), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3069) );
  AOI22_X1 U3908 ( .A1(n3036), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3038), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3068) );
  AOI22_X1 U3909 ( .A1(n3205), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3964), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3067) );
  AOI22_X1 U3910 ( .A1(n3157), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n3198), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3066) );
  NAND4_X1 U3911 ( .A1(n3069), .A2(n3068), .A3(n3067), .A4(n3066), .ZN(n3070)
         );
  OR2_X2 U3912 ( .A1(n3071), .A2(n3070), .ZN(n4013) );
  INV_X1 U3913 ( .A(n4012), .ZN(n3072) );
  NAND2_X1 U3914 ( .A1(n3971), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3078)
         );
  NAND2_X1 U3915 ( .A1(n3210), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3077)
         );
  NAND2_X1 U3916 ( .A1(n3164), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3076) );
  NAND2_X1 U3917 ( .A1(n3853), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3075)
         );
  NAND2_X1 U3918 ( .A1(n3851), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3082)
         );
  NAND2_X1 U3919 ( .A1(n2963), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3081) );
  NAND2_X1 U3920 ( .A1(n3036), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3080) );
  NAND2_X1 U3921 ( .A1(n3858), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3079) );
  NAND2_X1 U3922 ( .A1(n3205), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3086) );
  NAND2_X1 U3923 ( .A1(n3964), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3085) );
  NAND2_X1 U3924 ( .A1(n2966), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3084) );
  NAND2_X1 U3925 ( .A1(n3198), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3083)
         );
  NAND2_X1 U3926 ( .A1(n3061), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3090) );
  NAND2_X1 U3927 ( .A1(n3283), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3089)
         );
  NAND2_X1 U3928 ( .A1(n3163), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3088) );
  NAND2_X1 U3929 ( .A1(n3043), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3087) );
  AND4_X4 U3930 ( .A1(n3094), .A2(n3093), .A3(n3092), .A4(n3091), .ZN(n3135)
         );
  NAND2_X1 U3931 ( .A1(n3135), .A2(n4013), .ZN(n4223) );
  INV_X1 U3932 ( .A(n4223), .ZN(n3095) );
  OAI211_X1 U3933 ( .C1(n3137), .C2(n3109), .A(n3126), .B(n3095), .ZN(n3096)
         );
  AOI21_X1 U3934 ( .B1(n3239), .B2(n4191), .A(n3096), .ZN(n3115) );
  INV_X1 U3935 ( .A(n3104), .ZN(n3501) );
  NAND2_X1 U3936 ( .A1(n3501), .A2(n3109), .ZN(n3489) );
  AOI21_X1 U3937 ( .B1(n3489), .B2(n4382), .A(n4391), .ZN(n3107) );
  NAND2_X1 U3938 ( .A1(n5272), .A2(n3121), .ZN(n3098) );
  OAI21_X1 U3939 ( .B1(n3099), .B2(n5272), .A(n3098), .ZN(n3105) );
  OR2_X2 U3940 ( .A1(n3101), .A2(n3100), .ZN(n4276) );
  NAND2_X1 U3941 ( .A1(n3135), .A2(n3102), .ZN(n3103) );
  OR2_X2 U3942 ( .A1(n3104), .A2(n3103), .ZN(n3684) );
  OAI21_X1 U3943 ( .B1(n3105), .B2(n5270), .A(n3684), .ZN(n3106) );
  NAND2_X1 U3944 ( .A1(n3107), .A2(n3106), .ZN(n3108) );
  NAND2_X1 U3945 ( .A1(n3108), .A2(n4220), .ZN(n3119) );
  INV_X1 U3946 ( .A(n3124), .ZN(n3111) );
  NAND2_X1 U3947 ( .A1(n3111), .A2(n3110), .ZN(n3113) );
  NAND2_X1 U3948 ( .A1(n3113), .A2(n3112), .ZN(n3488) );
  NOR2_X2 U3949 ( .A1(n3488), .A2(n3114), .ZN(n3132) );
  NAND3_X1 U3950 ( .A1(n3115), .A2(n3119), .A3(n3132), .ZN(n3116) );
  NAND2_X2 U3951 ( .A1(n3116), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3148) );
  AND2_X1 U3952 ( .A1(n6391), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3491) );
  NOR2_X1 U3953 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_3__SCAN_IN), .ZN(
        n6384) );
  INV_X1 U3954 ( .A(n4000), .ZN(n3152) );
  MUX2_X1 U3955 ( .A(n3491), .B(n3152), .S(n6635), .Z(n3118) );
  OAI21_X2 U3956 ( .B1(n3148), .B2(n3117), .A(n3118), .ZN(n3192) );
  INV_X1 U3957 ( .A(n3119), .ZN(n3120) );
  NAND2_X1 U3958 ( .A1(n4192), .A2(n3155), .ZN(n3389) );
  NAND2_X1 U3959 ( .A1(n6384), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3122) );
  AOI21_X1 U3960 ( .B1(n4363), .B2(n4377), .A(n3122), .ZN(n3128) );
  INV_X1 U3961 ( .A(n3684), .ZN(n5277) );
  NAND2_X1 U3962 ( .A1(n5277), .A2(n3134), .ZN(n4527) );
  NAND2_X1 U3963 ( .A1(n4282), .A2(n4382), .ZN(n3125) );
  OAI21_X1 U3964 ( .B1(n4191), .B2(n3125), .A(n3239), .ZN(n3127) );
  INV_X1 U3966 ( .A(n3132), .ZN(n3129) );
  INV_X1 U3967 ( .A(n4382), .ZN(n3136) );
  OAI21_X1 U3968 ( .B1(n3129), .B2(n3136), .A(n4391), .ZN(n3130) );
  AND2_X2 U3969 ( .A1(n3192), .A2(n3190), .ZN(n3177) );
  NOR2_X1 U3970 ( .A1(n4223), .A2(n3109), .ZN(n3131) );
  NAND2_X1 U3971 ( .A1(n3132), .A2(n3131), .ZN(n4183) );
  INV_X1 U3972 ( .A(n4183), .ZN(n3133) );
  NAND2_X1 U3973 ( .A1(n3133), .A2(n3123), .ZN(n4114) );
  NAND3_X1 U3974 ( .A1(n3135), .A2(n5272), .A3(n3136), .ZN(n4333) );
  NAND2_X1 U3975 ( .A1(n4214), .A2(n4221), .ZN(n4203) );
  OAI211_X2 U3976 ( .C1(n4114), .C2(n3137), .A(n4505), .B(n4203), .ZN(n3145)
         );
  NAND2_X1 U3977 ( .A1(n6635), .A2(n4699), .ZN(n3138) );
  NAND2_X1 U3978 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3150) );
  AND2_X1 U3979 ( .A1(n3138), .A2(n3150), .ZN(n4700) );
  INV_X1 U3980 ( .A(n3491), .ZN(n3278) );
  AND2_X1 U3981 ( .A1(n3278), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3139)
         );
  AOI21_X1 U3982 ( .B1(n4000), .B2(n4700), .A(n3139), .ZN(n3143) );
  AOI21_X1 U3983 ( .B1(n3145), .B2(STATE2_REG_0__SCAN_IN), .A(n3140), .ZN(
        n3142) );
  NAND2_X1 U3984 ( .A1(n3142), .A2(n3141), .ZN(n3175) );
  NAND2_X1 U3985 ( .A1(n3177), .A2(n3175), .ZN(n3147) );
  NOR2_X1 U3986 ( .A1(n3140), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3144)
         );
  NOR2_X1 U3987 ( .A1(n3144), .A2(n6382), .ZN(n3146) );
  NAND2_X1 U3988 ( .A1(n3146), .A2(n3145), .ZN(n3176) );
  INV_X1 U3989 ( .A(n3148), .ZN(n3154) );
  INV_X1 U3990 ( .A(n3150), .ZN(n3149) );
  NAND2_X1 U3991 ( .A1(n3149), .A2(n4864), .ZN(n6189) );
  NAND2_X1 U3992 ( .A1(n3150), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3151) );
  AND2_X1 U3993 ( .A1(n6189), .A2(n3151), .ZN(n4623) );
  OAI22_X1 U3994 ( .A1(n4623), .A2(n3152), .B1(n3491), .B2(n4864), .ZN(n3153)
         );
  XNOR2_X1 U3995 ( .A(n3272), .B(n3273), .ZN(n4345) );
  NAND2_X1 U3996 ( .A1(n4345), .A2(n6382), .ZN(n3172) );
  AOI22_X1 U3997 ( .A1(n3852), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n3156), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3161) );
  AOI22_X1 U3998 ( .A1(n3965), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3859), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3160) );
  AOI22_X1 U3999 ( .A1(n3963), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3944), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3159) );
  AOI22_X1 U4000 ( .A1(n2966), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3974), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3158) );
  NAND4_X1 U4001 ( .A1(n3161), .A2(n3160), .A3(n3159), .A4(n3158), .ZN(n3170)
         );
  AOI22_X1 U4002 ( .A1(n3973), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n3162), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3168) );
  AOI22_X1 U4003 ( .A1(n3966), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3949), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3167) );
  AOI22_X1 U4004 ( .A1(n3925), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3972), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3166) );
  AOI22_X1 U4005 ( .A1(n3197), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3043), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3165) );
  NAND4_X1 U4006 ( .A1(n3168), .A2(n3167), .A3(n3166), .A4(n3165), .ZN(n3169)
         );
  NAND2_X1 U4007 ( .A1(n3226), .A2(n3238), .ZN(n3171) );
  NAND2_X1 U4008 ( .A1(n3172), .A2(n3171), .ZN(n3174) );
  NAND2_X1 U4009 ( .A1(n4220), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3281) );
  INV_X1 U4010 ( .A(n3281), .ZN(n3224) );
  AOI22_X1 U4011 ( .A1(n3432), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3224), 
        .B2(n3238), .ZN(n3173) );
  NAND2_X1 U4012 ( .A1(n3175), .A2(n3176), .ZN(n3178) );
  XNOR2_X2 U4013 ( .A(n3178), .B(n3177), .ZN(n4344) );
  BUF_X2 U4014 ( .A(n3061), .Z(n3949) );
  AOI22_X1 U4015 ( .A1(n3949), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3971), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3182) );
  AOI22_X1 U4016 ( .A1(n3965), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3852), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3181) );
  AOI22_X1 U4017 ( .A1(n3156), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n3944), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3180) );
  AOI22_X1 U4018 ( .A1(n3963), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3878), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3179) );
  NAND4_X1 U4019 ( .A1(n3182), .A2(n3181), .A3(n3180), .A4(n3179), .ZN(n3188)
         );
  AOI22_X1 U4020 ( .A1(n3966), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3973), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3186) );
  AOI22_X1 U4021 ( .A1(n3925), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3972), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3185) );
  AOI22_X1 U4022 ( .A1(n3859), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3157), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3184) );
  BUF_X1 U4023 ( .A(n3198), .Z(n3974) );
  AOI22_X1 U4024 ( .A1(n3197), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3974), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3183) );
  NAND4_X1 U4025 ( .A1(n3186), .A2(n3185), .A3(n3184), .A4(n3183), .ZN(n3187)
         );
  AND2_X1 U4026 ( .A1(n3226), .A2(n3249), .ZN(n3189) );
  INV_X1 U4027 ( .A(n3190), .ZN(n3191) );
  XNOR2_X1 U4028 ( .A(n3192), .B(n3191), .ZN(n3502) );
  NAND2_X1 U4029 ( .A1(n3502), .A2(n6382), .ZN(n3218) );
  AOI22_X1 U4030 ( .A1(n3966), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3971), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3196) );
  AOI22_X1 U4031 ( .A1(n3205), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3036), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3195) );
  AOI22_X1 U4032 ( .A1(n3963), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3944), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3194) );
  AOI22_X1 U4034 ( .A1(n3925), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3879), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3193) );
  NAND4_X1 U4035 ( .A1(n3196), .A2(n3195), .A3(n3194), .A4(n3193), .ZN(n3204)
         );
  AOI22_X1 U4036 ( .A1(n3949), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n3973), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3202) );
  AOI22_X1 U4037 ( .A1(n3197), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3878), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3201) );
  AOI22_X1 U4038 ( .A1(n3859), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3157), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3200) );
  AOI22_X1 U4039 ( .A1(n3852), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n3198), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3199) );
  NAND4_X1 U4040 ( .A1(n3202), .A2(n3201), .A3(n3200), .A4(n3199), .ZN(n3203)
         );
  INV_X1 U4041 ( .A(n3237), .ZN(n3260) );
  AOI22_X1 U4042 ( .A1(n3852), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n3036), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3209) );
  AOI22_X1 U4043 ( .A1(n3205), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3964), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3208) );
  INV_X1 U4044 ( .A(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n6614) );
  AOI22_X1 U4045 ( .A1(n3963), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3944), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3207) );
  AOI22_X1 U4046 ( .A1(n2966), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3198), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3206) );
  NAND4_X1 U4047 ( .A1(n3209), .A2(n3208), .A3(n3207), .A4(n3206), .ZN(n3216)
         );
  AOI22_X1 U4048 ( .A1(n3973), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n3971), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3214) );
  AOI22_X1 U4049 ( .A1(n3966), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3949), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3213) );
  AOI22_X1 U4050 ( .A1(n3925), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3879), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3212) );
  AOI22_X1 U4051 ( .A1(n3197), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3878), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3211) );
  NAND4_X1 U4052 ( .A1(n3214), .A2(n3213), .A3(n3212), .A4(n3211), .ZN(n3215)
         );
  XNOR2_X1 U4053 ( .A(n3260), .B(n3392), .ZN(n3217) );
  NAND2_X1 U4054 ( .A1(n3217), .A2(n3226), .ZN(n3257) );
  NAND2_X1 U4055 ( .A1(n3218), .A2(n3257), .ZN(n3258) );
  INV_X1 U4056 ( .A(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3221) );
  AOI21_X1 U4057 ( .B1(n3155), .B2(n3392), .A(n6382), .ZN(n3220) );
  NAND2_X1 U4058 ( .A1(n4220), .A2(n3237), .ZN(n3219) );
  NAND2_X1 U4059 ( .A1(n3258), .A2(n3255), .ZN(n3223) );
  NAND2_X1 U4060 ( .A1(n3226), .A2(n3392), .ZN(n3222) );
  INV_X1 U4061 ( .A(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3229) );
  NAND2_X1 U4062 ( .A1(n3224), .A2(n3249), .ZN(n3228) );
  INV_X1 U4063 ( .A(n3392), .ZN(n3225) );
  NAND2_X1 U4064 ( .A1(n3226), .A2(n3225), .ZN(n3227) );
  NAND2_X1 U4065 ( .A1(n3244), .A2(n3245), .ZN(n3232) );
  INV_X1 U4066 ( .A(n3244), .ZN(n3231) );
  INV_X1 U4067 ( .A(n3245), .ZN(n3230) );
  NAND2_X1 U4069 ( .A1(n3298), .A2(n3235), .ZN(n3493) );
  INV_X1 U4070 ( .A(n3493), .ZN(n3236) );
  NAND2_X1 U4071 ( .A1(n3236), .A2(n4192), .ZN(n3242) );
  NAND2_X1 U4072 ( .A1(n3237), .A2(n3249), .ZN(n3301) );
  INV_X1 U4073 ( .A(n3238), .ZN(n3300) );
  XNOR2_X1 U4074 ( .A(n3301), .B(n3300), .ZN(n3240) );
  AND2_X1 U4075 ( .A1(n4220), .A2(n4382), .ZN(n3259) );
  AOI21_X1 U4076 ( .B1(n3240), .B2(n4394), .A(n3259), .ZN(n3241) );
  NAND2_X1 U4077 ( .A1(n3242), .A2(n3241), .ZN(n5965) );
  NAND2_X1 U4078 ( .A1(n5965), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3268)
         );
  INV_X1 U4079 ( .A(n3243), .ZN(n3248) );
  NAND2_X1 U4080 ( .A1(n4343), .A2(n4192), .ZN(n3254) );
  XNOR2_X1 U4081 ( .A(n3260), .B(n3249), .ZN(n3250) );
  NAND2_X1 U4082 ( .A1(n3250), .A2(n4394), .ZN(n3252) );
  NOR2_X1 U4083 ( .A1(n4223), .A2(n5272), .ZN(n3251) );
  AND2_X1 U4084 ( .A1(n3252), .A2(n3251), .ZN(n3253) );
  NAND2_X1 U4085 ( .A1(n3254), .A2(n3253), .ZN(n4317) );
  INV_X1 U4086 ( .A(n3255), .ZN(n3256) );
  INV_X1 U4087 ( .A(n4192), .ZN(n3262) );
  AOI21_X1 U4088 ( .B1(n3260), .B2(n4394), .A(n3259), .ZN(n3261) );
  OAI21_X2 U4089 ( .B1(n4764), .B2(n3262), .A(n3261), .ZN(n4302) );
  NAND2_X1 U4090 ( .A1(n4302), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n3263)
         );
  INV_X1 U4091 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n5149) );
  NAND2_X1 U4092 ( .A1(n3263), .A2(n5149), .ZN(n3265) );
  AND2_X1 U4093 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n3264) );
  NAND2_X1 U4094 ( .A1(n4302), .A2(n3264), .ZN(n3266) );
  AND2_X1 U4095 ( .A1(n3265), .A2(n3266), .ZN(n4316) );
  INV_X1 U4096 ( .A(n3266), .ZN(n3267) );
  NAND2_X1 U4097 ( .A1(n3268), .A2(n5966), .ZN(n3271) );
  INV_X1 U4098 ( .A(n5965), .ZN(n3269) );
  INV_X1 U4099 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n5964) );
  NAND2_X1 U4100 ( .A1(n3269), .A2(n5964), .ZN(n3270) );
  AND2_X1 U4101 ( .A1(n3271), .A2(n3270), .ZN(n5956) );
  INV_X1 U4102 ( .A(n3298), .ZN(n3296) );
  INV_X1 U4103 ( .A(n3273), .ZN(n3274) );
  INV_X1 U4104 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3275) );
  OR2_X1 U4105 ( .A1(n3148), .A2(n3275), .ZN(n3280) );
  NAND3_X1 U4106 ( .A1(n6358), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6126) );
  INV_X1 U4107 ( .A(n6126), .ZN(n3276) );
  NAND2_X1 U4108 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n3276), .ZN(n6122) );
  NAND2_X1 U4109 ( .A1(n6358), .A2(n6122), .ZN(n3277) );
  NOR3_X1 U4110 ( .A1(n6358), .A2(n4864), .A3(n4699), .ZN(n4656) );
  NAND2_X1 U4111 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4656), .ZN(n4446) );
  AND2_X1 U4112 ( .A1(n3277), .A2(n4446), .ZN(n6157) );
  AOI22_X1 U4113 ( .A1(n4000), .A2(n6157), .B1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n3278), .ZN(n3279) );
  AOI22_X1 U4114 ( .A1(n3973), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n3925), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3287) );
  AOI22_X1 U4115 ( .A1(n3197), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3966), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3286) );
  AOI22_X1 U4116 ( .A1(n3156), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3944), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3285) );
  AOI22_X1 U4117 ( .A1(n3963), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3878), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3284) );
  NAND4_X1 U4118 ( .A1(n3287), .A2(n3286), .A3(n3285), .A4(n3284), .ZN(n3293)
         );
  AOI22_X1 U4119 ( .A1(n3949), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3852), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3291) );
  AOI22_X1 U4120 ( .A1(n3965), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3964), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3290) );
  AOI22_X1 U4121 ( .A1(n3971), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3879), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3289) );
  AOI22_X1 U4122 ( .A1(n3157), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3974), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3288) );
  NAND4_X1 U4123 ( .A1(n3291), .A2(n3290), .A3(n3289), .A4(n3288), .ZN(n3292)
         );
  OR2_X1 U4124 ( .A1(n3293), .A2(n3292), .ZN(n3319) );
  AOI22_X1 U4125 ( .A1(n3485), .A2(n3319), .B1(n3432), .B2(
        INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3294) );
  NAND2_X2 U4126 ( .A1(n3296), .A2(n3297), .ZN(n3328) );
  NAND2_X1 U4127 ( .A1(n3298), .A2(n4417), .ZN(n3299) );
  NAND2_X1 U4128 ( .A1(n3328), .A2(n3299), .ZN(n3518) );
  NAND2_X1 U4129 ( .A1(n3301), .A2(n3300), .ZN(n3320) );
  INV_X1 U4130 ( .A(n3319), .ZN(n3302) );
  XNOR2_X1 U4131 ( .A(n3320), .B(n3302), .ZN(n3303) );
  NAND2_X1 U4132 ( .A1(n3303), .A2(n4394), .ZN(n3304) );
  OAI21_X1 U4133 ( .B1(n3518), .B2(n3262), .A(n3304), .ZN(n3305) );
  INV_X1 U4134 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n6038) );
  XNOR2_X1 U4135 ( .A(n3305), .B(n6038), .ZN(n5955) );
  NAND2_X1 U4136 ( .A1(n5956), .A2(n5955), .ZN(n5958) );
  NAND2_X1 U4137 ( .A1(n3305), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n3306)
         );
  NAND2_X1 U4138 ( .A1(n5958), .A2(n3306), .ZN(n4794) );
  AOI22_X1 U4139 ( .A1(n3852), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n3156), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3310) );
  AOI22_X1 U4140 ( .A1(n3965), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3964), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3309) );
  AOI22_X1 U4141 ( .A1(INSTQUEUE_REG_12__4__SCAN_IN), .A2(n3963), .B1(n3944), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3308) );
  AOI22_X1 U4142 ( .A1(n2966), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n3974), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3307) );
  NAND4_X1 U4143 ( .A1(n3310), .A2(n3309), .A3(n3308), .A4(n3307), .ZN(n3316)
         );
  AOI22_X1 U4144 ( .A1(INSTQUEUE_REG_15__4__SCAN_IN), .A2(n3973), .B1(n3971), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3314) );
  AOI22_X1 U4145 ( .A1(n3966), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3949), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3313) );
  AOI22_X1 U4146 ( .A1(INSTQUEUE_REG_8__4__SCAN_IN), .A2(n3925), .B1(n3879), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3312) );
  AOI22_X1 U4147 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n3197), .B1(n3878), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3311) );
  NAND4_X1 U4148 ( .A1(n3314), .A2(n3313), .A3(n3312), .A4(n3311), .ZN(n3315)
         );
  NAND2_X1 U4149 ( .A1(n3485), .A2(n3342), .ZN(n3318) );
  NAND2_X1 U4150 ( .A1(n3432), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3317) );
  NAND2_X1 U4151 ( .A1(n3318), .A2(n3317), .ZN(n3326) );
  NAND2_X1 U4152 ( .A1(n3534), .A2(n4192), .ZN(n3323) );
  NAND2_X1 U4153 ( .A1(n3320), .A2(n3319), .ZN(n3344) );
  XNOR2_X1 U4154 ( .A(n3344), .B(n3342), .ZN(n3321) );
  NAND2_X1 U4155 ( .A1(n3321), .A2(n4394), .ZN(n3322) );
  NAND2_X1 U4156 ( .A1(n3323), .A2(n3322), .ZN(n3324) );
  INV_X1 U4157 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n6031) );
  XNOR2_X1 U4158 ( .A(n3324), .B(n6031), .ZN(n4793) );
  NAND2_X1 U4159 ( .A1(n4794), .A2(n4793), .ZN(n4792) );
  NAND2_X1 U4160 ( .A1(n3324), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n3325)
         );
  NAND2_X1 U4161 ( .A1(n4792), .A2(n3325), .ZN(n5949) );
  INV_X1 U4162 ( .A(n3351), .ZN(n3341) );
  AOI22_X1 U4163 ( .A1(n3966), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3971), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3332) );
  AOI22_X1 U4164 ( .A1(n3197), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3949), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3331) );
  AOI22_X1 U4165 ( .A1(n3965), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3964), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3330) );
  AOI22_X1 U4166 ( .A1(n3156), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3974), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3329) );
  NAND4_X1 U4167 ( .A1(n3332), .A2(n3331), .A3(n3330), .A4(n3329), .ZN(n3338)
         );
  AOI22_X1 U4168 ( .A1(n3963), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3944), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3336) );
  AOI22_X1 U4169 ( .A1(n3925), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3879), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3335) );
  AOI22_X1 U4170 ( .A1(n3973), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n3878), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3334) );
  AOI22_X1 U4171 ( .A1(n3852), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n3157), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3333) );
  NAND4_X1 U4172 ( .A1(n3336), .A2(n3335), .A3(n3334), .A4(n3333), .ZN(n3337)
         );
  OR2_X1 U4173 ( .A1(n3338), .A2(n3337), .ZN(n3370) );
  NAND2_X1 U4174 ( .A1(n3485), .A2(n3370), .ZN(n3340) );
  NAND2_X1 U4175 ( .A1(n3432), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3339) );
  NAND2_X1 U4176 ( .A1(n3340), .A2(n3339), .ZN(n3350) );
  XNOR2_X1 U4177 ( .A(n3341), .B(n3350), .ZN(n3539) );
  NAND2_X1 U4178 ( .A1(n3539), .A2(n4192), .ZN(n3347) );
  INV_X1 U4179 ( .A(n3342), .ZN(n3343) );
  OR2_X1 U4180 ( .A1(n3344), .A2(n3343), .ZN(n3369) );
  XNOR2_X1 U4181 ( .A(n3369), .B(n3370), .ZN(n3345) );
  NAND2_X1 U4182 ( .A1(n3345), .A2(n4394), .ZN(n3346) );
  NAND2_X1 U4183 ( .A1(n3347), .A2(n3346), .ZN(n3348) );
  INV_X1 U4184 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4241) );
  XNOR2_X1 U4185 ( .A(n3348), .B(n4241), .ZN(n5948) );
  NAND2_X1 U4186 ( .A1(n5949), .A2(n5948), .ZN(n5947) );
  NAND2_X1 U4187 ( .A1(n3348), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n3349)
         );
  NAND2_X1 U4188 ( .A1(n5947), .A2(n3349), .ZN(n4570) );
  INV_X1 U4189 ( .A(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n6645) );
  AOI22_X1 U4190 ( .A1(n3852), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n3156), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3355) );
  AOI22_X1 U4191 ( .A1(n3965), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3859), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3354) );
  AOI22_X1 U4192 ( .A1(n3963), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3944), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3353) );
  AOI22_X1 U4193 ( .A1(n3157), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3974), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3352) );
  NAND4_X1 U4194 ( .A1(n3355), .A2(n3354), .A3(n3353), .A4(n3352), .ZN(n3362)
         );
  INV_X1 U4195 ( .A(n3971), .ZN(n3356) );
  INV_X1 U4196 ( .A(n3356), .ZN(n3924) );
  AOI22_X1 U4197 ( .A1(n3973), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n3924), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3360) );
  AOI22_X1 U4198 ( .A1(n3966), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3949), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3359) );
  AOI22_X1 U4199 ( .A1(n3925), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3879), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3358) );
  AOI22_X1 U4200 ( .A1(n3197), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3878), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3357) );
  NAND4_X1 U4201 ( .A1(n3360), .A2(n3359), .A3(n3358), .A4(n3357), .ZN(n3361)
         );
  OR2_X1 U4202 ( .A1(n3362), .A2(n3361), .ZN(n3381) );
  NAND2_X1 U4203 ( .A1(n3485), .A2(n3381), .ZN(n3364) );
  NAND2_X1 U4204 ( .A1(n3432), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3363) );
  NAND2_X1 U4205 ( .A1(n3368), .A2(n3367), .ZN(n3535) );
  NAND3_X1 U4206 ( .A1(n3391), .A2(n3535), .A3(n4192), .ZN(n3374) );
  INV_X1 U4207 ( .A(n3369), .ZN(n3371) );
  NAND2_X1 U4208 ( .A1(n3371), .A2(n3370), .ZN(n3380) );
  XNOR2_X1 U4209 ( .A(n3380), .B(n3381), .ZN(n3372) );
  NAND2_X1 U4210 ( .A1(n3372), .A2(n4394), .ZN(n3373) );
  NAND2_X1 U4211 ( .A1(n3374), .A2(n3373), .ZN(n3375) );
  INV_X1 U4212 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n4240) );
  XNOR2_X1 U4213 ( .A(n3375), .B(n4240), .ZN(n4569) );
  NAND2_X1 U4214 ( .A1(n4570), .A2(n4569), .ZN(n4568) );
  NAND2_X1 U4215 ( .A1(n3375), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n3376)
         );
  NAND2_X1 U4216 ( .A1(n4568), .A2(n3376), .ZN(n5941) );
  INV_X1 U4217 ( .A(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3378) );
  NAND2_X1 U4218 ( .A1(n3485), .A2(n3392), .ZN(n3377) );
  OAI21_X1 U4219 ( .B1(n3378), .B2(n3471), .A(n3377), .ZN(n3379) );
  NAND2_X1 U4220 ( .A1(n3548), .A2(n4192), .ZN(n3385) );
  INV_X1 U4221 ( .A(n3380), .ZN(n3382) );
  NAND2_X1 U4222 ( .A1(n3382), .A2(n3381), .ZN(n3394) );
  XNOR2_X1 U4223 ( .A(n3394), .B(n3392), .ZN(n3383) );
  NAND2_X1 U4224 ( .A1(n3383), .A2(n4394), .ZN(n3384) );
  NAND2_X1 U4225 ( .A1(n3385), .A2(n3384), .ZN(n3386) );
  INV_X1 U4226 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n6570) );
  XNOR2_X1 U4227 ( .A(n3386), .B(n6570), .ZN(n5940) );
  NAND2_X1 U4228 ( .A1(n5941), .A2(n5940), .ZN(n5939) );
  NAND2_X1 U4229 ( .A1(n3386), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n3387)
         );
  NAND2_X1 U4230 ( .A1(n5939), .A2(n3387), .ZN(n4858) );
  NAND2_X1 U4231 ( .A1(n3392), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3388) );
  NOR2_X1 U4232 ( .A1(n3389), .A2(n3388), .ZN(n3390) );
  NAND2_X1 U4233 ( .A1(n4394), .A2(n3392), .ZN(n3393) );
  OR2_X1 U4234 ( .A1(n3394), .A2(n3393), .ZN(n3395) );
  NAND2_X1 U4235 ( .A1(n3422), .A2(n3395), .ZN(n3396) );
  INV_X1 U4236 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n6006) );
  XNOR2_X1 U4237 ( .A(n3396), .B(n6006), .ZN(n4857) );
  NAND2_X1 U4238 ( .A1(n4858), .A2(n4857), .ZN(n4856) );
  NAND2_X1 U4239 ( .A1(n3396), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n3397)
         );
  NAND2_X1 U4240 ( .A1(n4856), .A2(n3397), .ZN(n4910) );
  INV_X1 U4241 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n5997) );
  NAND2_X1 U4242 ( .A1(n3422), .A2(n5997), .ZN(n4911) );
  NAND2_X1 U4243 ( .A1(n4910), .A2(n4911), .ZN(n3398) );
  NAND2_X1 U4244 ( .A1(n3398), .A2(n4912), .ZN(n4943) );
  INV_X1 U4245 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n3399) );
  NAND2_X1 U4246 ( .A1(n3422), .A2(n3399), .ZN(n4942) );
  NAND2_X1 U4247 ( .A1(n4943), .A2(n4942), .ZN(n4964) );
  INV_X1 U4248 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n5988) );
  INV_X1 U4249 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n3402) );
  NAND2_X1 U4250 ( .A1(n3422), .A2(n3402), .ZN(n5022) );
  NAND2_X1 U4251 ( .A1(n5076), .A2(n5075), .ZN(n3406) );
  INV_X1 U4252 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n3404) );
  NAND2_X1 U4253 ( .A1(n3422), .A2(n3404), .ZN(n3405) );
  NAND2_X1 U4254 ( .A1(n3406), .A2(n3405), .ZN(n5082) );
  INV_X1 U4255 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5083) );
  OAI21_X2 U4256 ( .B1(n5082), .B2(n3408), .A(n3407), .ZN(n5138) );
  INV_X1 U4257 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5162) );
  NOR2_X1 U4258 ( .A1(n3422), .A2(n5162), .ZN(n3410) );
  NAND2_X1 U4259 ( .A1(n3422), .A2(n5162), .ZN(n3409) );
  OAI21_X1 U4260 ( .B1(n5138), .B2(n3410), .A(n3409), .ZN(n5205) );
  BUF_X2 U4261 ( .A(n5205), .Z(n5529) );
  INV_X1 U4262 ( .A(n5529), .ZN(n3414) );
  INV_X1 U4263 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5161) );
  AND2_X1 U4264 ( .A1(n3422), .A2(n5161), .ZN(n5204) );
  NAND2_X1 U4265 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n4256) );
  NAND2_X1 U4266 ( .A1(n3422), .A2(n4256), .ZN(n5517) );
  AND2_X1 U4267 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5579) );
  AND2_X1 U4268 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n4239) );
  AND2_X1 U4269 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n4258) );
  NAND3_X1 U4270 ( .A1(n5579), .A2(n4239), .A3(n4258), .ZN(n3411) );
  NAND2_X1 U4271 ( .A1(n3422), .A2(n3411), .ZN(n3412) );
  INV_X1 U4272 ( .A(n5472), .ZN(n3413) );
  OR2_X1 U4273 ( .A1(n5204), .A2(n3413), .ZN(n3425) );
  INV_X1 U4274 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5209) );
  AND2_X1 U4275 ( .A1(n3422), .A2(n5209), .ZN(n3419) );
  NAND2_X1 U4276 ( .A1(n3414), .A2(n2974), .ZN(n3421) );
  NOR2_X1 U4277 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n3415) );
  OR2_X1 U4278 ( .A1(n3422), .A2(n3415), .ZN(n3416) );
  OR2_X1 U4279 ( .A1(n3422), .A2(n5161), .ZN(n5527) );
  NOR2_X1 U4280 ( .A1(INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5263) );
  NOR2_X1 U4281 ( .A1(INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5580) );
  INV_X1 U4282 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5510) );
  INV_X1 U4283 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5613) );
  NAND4_X1 U4284 ( .A1(n5263), .A2(n5580), .A3(n5510), .A4(n5613), .ZN(n3417)
         );
  NAND2_X1 U4285 ( .A1(n3403), .A2(n3417), .ZN(n3418) );
  AND2_X1 U4286 ( .A1(n5481), .A2(n3418), .ZN(n5207) );
  XNOR2_X1 U4287 ( .A(n3422), .B(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5475)
         );
  AND2_X1 U4288 ( .A1(n5207), .A2(n5475), .ZN(n3426) );
  AND2_X2 U4289 ( .A1(n3421), .A2(n3420), .ZN(n5466) );
  INV_X1 U4290 ( .A(n5466), .ZN(n3423) );
  NAND3_X1 U4291 ( .A1(n3423), .A2(n3422), .A3(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n4178) );
  AND2_X1 U4292 ( .A1(INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5543) );
  NAND2_X1 U4293 ( .A1(n5543), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n3424) );
  NOR2_X1 U4294 ( .A1(n4178), .A2(n3424), .ZN(n5185) );
  OR2_X1 U4295 ( .A1(n5529), .A2(n3425), .ZN(n3427) );
  NAND2_X1 U4296 ( .A1(n3427), .A2(n3426), .ZN(n5474) );
  INV_X1 U4297 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5455) );
  INV_X1 U4298 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n6586) );
  NAND2_X1 U4299 ( .A1(n5455), .A2(n6586), .ZN(n5545) );
  OR2_X1 U4300 ( .A1(n3422), .A2(n5545), .ZN(n4179) );
  INV_X1 U4301 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5195) );
  INV_X1 U4302 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5208) );
  NAND2_X1 U4303 ( .A1(n5195), .A2(n5208), .ZN(n3428) );
  OR2_X1 U4304 ( .A1(n4179), .A2(n3428), .ZN(n5182) );
  NOR3_X1 U4305 ( .A1(n5474), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .A3(n5182), 
        .ZN(n3429) );
  INV_X1 U4306 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n6623) );
  INV_X1 U4307 ( .A(n5201), .ZN(n3492) );
  NAND2_X1 U4308 ( .A1(n3485), .A2(n4391), .ZN(n3431) );
  NAND2_X1 U4309 ( .A1(n3431), .A2(n3109), .ZN(n3444) );
  XNOR2_X1 U4310 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3448) );
  XNOR2_X1 U4311 ( .A(n3448), .B(n3449), .ZN(n4119) );
  INV_X1 U4312 ( .A(n4119), .ZN(n3443) );
  AND2_X1 U4313 ( .A1(n3117), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n3433)
         );
  NOR2_X1 U4314 ( .A1(n3449), .A2(n3433), .ZN(n3437) );
  NAND2_X1 U4315 ( .A1(n3485), .A2(n3437), .ZN(n3434) );
  NAND2_X1 U4316 ( .A1(n3463), .A2(n3434), .ZN(n3442) );
  INV_X1 U4317 ( .A(n3435), .ZN(n3436) );
  AOI21_X1 U4318 ( .B1(n3438), .B2(n3437), .A(n3436), .ZN(n3440) );
  NAND2_X1 U4319 ( .A1(n4217), .A2(n3109), .ZN(n3439) );
  NAND2_X1 U4320 ( .A1(n5301), .A2(n3439), .ZN(n3452) );
  OR2_X1 U4321 ( .A1(n3440), .A2(n3452), .ZN(n3441) );
  OAI211_X1 U4322 ( .C1(n3444), .C2(n3443), .A(n3442), .B(n3441), .ZN(n3447)
         );
  NAND3_X1 U4323 ( .A1(n3444), .A2(STATE2_REG_0__SCAN_IN), .A3(n3443), .ZN(
        n3446) );
  NAND2_X1 U4324 ( .A1(n3481), .A2(n4119), .ZN(n3445) );
  NAND3_X1 U4325 ( .A1(n3447), .A2(n3446), .A3(n3445), .ZN(n3458) );
  NAND2_X1 U4326 ( .A1(n3449), .A2(n3448), .ZN(n3451) );
  NAND2_X1 U4327 ( .A1(n4699), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3450) );
  NAND2_X1 U4328 ( .A1(n3451), .A2(n3450), .ZN(n3460) );
  XNOR2_X1 U4329 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3459) );
  XNOR2_X1 U4330 ( .A(n3460), .B(n3459), .ZN(n4118) );
  INV_X1 U4331 ( .A(n4118), .ZN(n3453) );
  NAND2_X1 U4332 ( .A1(n3485), .A2(n3453), .ZN(n3455) );
  INV_X1 U4333 ( .A(n3452), .ZN(n3454) );
  OAI211_X1 U4334 ( .C1(n3453), .C2(n3471), .A(n3455), .B(n3454), .ZN(n3457)
         );
  NOR2_X1 U4335 ( .A1(n3455), .A2(n3454), .ZN(n3456) );
  AOI21_X1 U4336 ( .B1(n3458), .B2(n3457), .A(n3456), .ZN(n3466) );
  NAND2_X1 U4337 ( .A1(n3460), .A2(n3459), .ZN(n3462) );
  NAND2_X1 U4338 ( .A1(n4864), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3461) );
  NAND2_X1 U4339 ( .A1(n3462), .A2(n3461), .ZN(n3469) );
  XNOR2_X1 U4340 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3468) );
  XNOR2_X1 U4341 ( .A(n3469), .B(n3468), .ZN(n4120) );
  AND2_X1 U4342 ( .A1(n3471), .A2(n4120), .ZN(n3465) );
  INV_X1 U4343 ( .A(n4120), .ZN(n3464) );
  OAI22_X1 U4344 ( .A1(n3466), .A2(n3465), .B1(n3464), .B2(n3463), .ZN(n3473)
         );
  NOR2_X1 U4345 ( .A1(n3275), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3467)
         );
  AOI21_X1 U4346 ( .B1(n3469), .B2(n3468), .A(n3467), .ZN(n3476) );
  INV_X1 U4347 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n6056) );
  NOR2_X1 U4348 ( .A1(n6056), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n3470)
         );
  AND2_X1 U4349 ( .A1(n3476), .A2(n3470), .ZN(n4117) );
  NAND2_X1 U4350 ( .A1(n3471), .A2(n4117), .ZN(n3472) );
  NAND2_X1 U4351 ( .A1(n3473), .A2(n3472), .ZN(n3475) );
  AOI22_X1 U4352 ( .A1(n3481), .A2(n4117), .B1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n6382), .ZN(n3474) );
  NAND2_X1 U4353 ( .A1(n3475), .A2(n3474), .ZN(n3483) );
  INV_X1 U4354 ( .A(n3476), .ZN(n3478) );
  AND2_X1 U4355 ( .A1(n6056), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n3477)
         );
  OR2_X1 U4356 ( .A1(n3478), .A2(n3477), .ZN(n3480) );
  NAND2_X1 U4357 ( .A1(n4498), .A2(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n3479) );
  NAND2_X1 U4358 ( .A1(n3480), .A2(n3479), .ZN(n4122) );
  INV_X1 U4359 ( .A(n4122), .ZN(n3484) );
  NAND2_X1 U4360 ( .A1(n3481), .A2(n3484), .ZN(n3482) );
  NAND2_X1 U4361 ( .A1(n3485), .A2(n3484), .ZN(n3486) );
  INV_X1 U4362 ( .A(n3488), .ZN(n4227) );
  AOI21_X1 U4363 ( .B1(n3489), .B2(n4220), .A(n4223), .ZN(n3490) );
  AND2_X1 U4364 ( .A1(n4227), .A2(n3490), .ZN(n4200) );
  NAND2_X1 U4365 ( .A1(n4200), .A2(n3073), .ZN(n4201) );
  OR2_X1 U4366 ( .A1(n5302), .A2(n4201), .ZN(n6363) );
  AND2_X1 U4367 ( .A1(n3491), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6383) );
  INV_X1 U4368 ( .A(n6383), .ZN(n6369) );
  NAND2_X1 U4369 ( .A1(n3492), .A2(n5968), .ZN(n4011) );
  NAND2_X1 U4370 ( .A1(n3494), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3682) );
  NAND2_X1 U4371 ( .A1(n3236), .A2(n3662), .ZN(n3495) );
  INV_X2 U4372 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n6379) );
  NAND2_X1 U4373 ( .A1(n6379), .A2(STATEBS16_REG_SCAN_IN), .ZN(n3997) );
  INV_X1 U4374 ( .A(n3682), .ZN(n3662) );
  NAND2_X1 U4375 ( .A1(n4343), .A2(n3662), .ZN(n3500) );
  AND2_X1 U4376 ( .A1(n4221), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3509) );
  NAND2_X1 U4377 ( .A1(n3509), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3498) );
  OR2_X1 U4378 ( .A1(n5271), .A2(n6379), .ZN(n3998) );
  AOI22_X1 U4379 ( .A1(n3987), .A2(EAX_REG_1__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n6379), .ZN(n3497) );
  AND2_X1 U4380 ( .A1(n3498), .A2(n3497), .ZN(n3499) );
  NAND2_X1 U4381 ( .A1(n3500), .A2(n3499), .ZN(n4300) );
  AOI21_X1 U4382 ( .B1(n4764), .B2(n3501), .A(n6379), .ZN(n4273) );
  INV_X1 U4383 ( .A(n3503), .ZN(n6346) );
  NAND2_X1 U4384 ( .A1(n3503), .A2(n3662), .ZN(n3507) );
  NAND2_X1 U4385 ( .A1(n3509), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3505) );
  AOI22_X1 U4386 ( .A1(n3987), .A2(EAX_REG_0__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n6379), .ZN(n3504) );
  AND2_X1 U4387 ( .A1(n3505), .A2(n3504), .ZN(n3506) );
  NAND2_X1 U4388 ( .A1(n3507), .A2(n3506), .ZN(n4272) );
  NAND2_X1 U4389 ( .A1(n4273), .A2(n4272), .ZN(n4271) );
  INV_X1 U4390 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n6234) );
  NAND2_X1 U4391 ( .A1(n6379), .A2(n6234), .ZN(n4123) );
  OR2_X1 U4392 ( .A1(n4272), .A2(n4123), .ZN(n3508) );
  NAND2_X1 U4393 ( .A1(n4271), .A2(n3508), .ZN(n4299) );
  NAND2_X1 U4394 ( .A1(n4300), .A2(n4299), .ZN(n4298) );
  INV_X1 U4395 ( .A(n3509), .ZN(n3530) );
  CLKBUF_X1 U4396 ( .A(n3510), .Z(n5156) );
  INV_X1 U4397 ( .A(n4123), .ZN(n3993) );
  OAI21_X1 U4398 ( .B1(PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .A(n3519), .ZN(n5972) );
  INV_X1 U4399 ( .A(n3997), .ZN(n3899) );
  AOI22_X1 U4400 ( .A1(n3993), .A2(n5972), .B1(n3899), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3512) );
  NAND2_X1 U4401 ( .A1(n3987), .A2(EAX_REG_2__SCAN_IN), .ZN(n3511) );
  OAI211_X1 U4402 ( .C1(n3530), .C2(n5156), .A(n3512), .B(n3511), .ZN(n4327)
         );
  NAND2_X1 U4403 ( .A1(n4328), .A2(n4327), .ZN(n3517) );
  INV_X1 U4404 ( .A(n4298), .ZN(n3515) );
  INV_X1 U4405 ( .A(n3513), .ZN(n3514) );
  NAND2_X1 U4406 ( .A1(n3515), .A2(n3514), .ZN(n3516) );
  OAI21_X1 U4407 ( .B1(PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n3520), .A(n3527), 
        .ZN(n5962) );
  AOI22_X1 U4408 ( .A1(n3993), .A2(n5962), .B1(n3899), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3522) );
  INV_X2 U4409 ( .A(n3998), .ZN(n3987) );
  NAND2_X1 U4410 ( .A1(n3987), .A2(EAX_REG_3__SCAN_IN), .ZN(n3521) );
  OAI211_X1 U4411 ( .C1(n3530), .C2(n3275), .A(n3522), .B(n3521), .ZN(n3523)
         );
  INV_X1 U4412 ( .A(n3523), .ZN(n3524) );
  NAND2_X1 U4414 ( .A1(n4326), .A2(n4476), .ZN(n4552) );
  AOI21_X1 U4415 ( .B1(n3527), .B2(n3526), .A(n3541), .ZN(n4795) );
  INV_X1 U4416 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4498) );
  NAND2_X1 U4417 ( .A1(n6379), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3529)
         );
  NAND2_X1 U4418 ( .A1(n3987), .A2(EAX_REG_4__SCAN_IN), .ZN(n3528) );
  OAI211_X1 U4419 ( .C1(n3530), .C2(n4498), .A(n3529), .B(n3528), .ZN(n3531)
         );
  NAND2_X1 U4420 ( .A1(n3531), .A2(n4123), .ZN(n3532) );
  OAI21_X1 U4421 ( .B1(n4795), .B2(n4123), .A(n3532), .ZN(n3533) );
  OR2_X2 U4422 ( .A1(n4552), .A2(n4553), .ZN(n4612) );
  NAND2_X1 U4423 ( .A1(n3535), .A2(n3662), .ZN(n3538) );
  AOI21_X1 U4424 ( .B1(n6571), .B2(n3540), .A(n3549), .ZN(n4801) );
  AOI22_X1 U4425 ( .A1(n3987), .A2(EAX_REG_6__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n6379), .ZN(n3536) );
  MUX2_X1 U4426 ( .A(n4801), .B(n3536), .S(n4123), .Z(n3537) );
  NAND2_X1 U4427 ( .A1(n3539), .A2(n3662), .ZN(n3546) );
  INV_X1 U4428 ( .A(EAX_REG_5__SCAN_IN), .ZN(n4614) );
  OAI21_X1 U4429 ( .B1(n3541), .B2(PHYADDRPOINTER_REG_5__SCAN_IN), .A(n3540), 
        .ZN(n5954) );
  NAND2_X1 U4430 ( .A1(n5954), .A2(n3993), .ZN(n3543) );
  NAND2_X1 U4431 ( .A1(n3899), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3542)
         );
  OAI211_X1 U4432 ( .C1(n3998), .C2(n4614), .A(n3543), .B(n3542), .ZN(n3544)
         );
  INV_X1 U4433 ( .A(n3544), .ZN(n3545) );
  OAI21_X1 U4434 ( .B1(n3549), .B2(PHYADDRPOINTER_REG_7__SCAN_IN), .A(n3554), 
        .ZN(n5946) );
  NAND2_X1 U4435 ( .A1(n5946), .A2(n3993), .ZN(n3551) );
  AOI22_X1 U4436 ( .A1(n3987), .A2(EAX_REG_7__SCAN_IN), .B1(n3899), .B2(
        PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3550) );
  AND2_X1 U4437 ( .A1(n3551), .A2(n3550), .ZN(n3552) );
  INV_X1 U4438 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n6636) );
  AOI21_X1 U4439 ( .B1(n6636), .B2(n3554), .A(n3587), .ZN(n4859) );
  OR2_X1 U4440 ( .A1(n4859), .A2(n4123), .ZN(n3570) );
  AOI22_X1 U4441 ( .A1(n3965), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3859), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3558) );
  AOI22_X1 U4442 ( .A1(n3963), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n3944), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3557) );
  AOI22_X1 U4443 ( .A1(n3973), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n3879), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3556) );
  AOI22_X1 U4444 ( .A1(n3156), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n3974), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3555) );
  NAND4_X1 U4445 ( .A1(n3558), .A2(n3557), .A3(n3556), .A4(n3555), .ZN(n3564)
         );
  AOI22_X1 U4446 ( .A1(n3966), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3949), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3562) );
  AOI22_X1 U4447 ( .A1(n3971), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n3925), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3561) );
  AOI22_X1 U4448 ( .A1(n3197), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3878), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3560) );
  AOI22_X1 U4449 ( .A1(n3852), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n3157), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3559) );
  NAND4_X1 U4450 ( .A1(n3562), .A2(n3561), .A3(n3560), .A4(n3559), .ZN(n3563)
         );
  NOR2_X1 U4451 ( .A1(n3564), .A2(n3563), .ZN(n3567) );
  NAND2_X1 U4452 ( .A1(n3987), .A2(EAX_REG_8__SCAN_IN), .ZN(n3566) );
  NAND2_X1 U4453 ( .A1(n3899), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3565)
         );
  OAI211_X1 U4454 ( .C1(n3682), .C2(n3567), .A(n3566), .B(n3565), .ZN(n3568)
         );
  INV_X1 U4455 ( .A(n3568), .ZN(n3569) );
  NAND2_X1 U4456 ( .A1(n3570), .A2(n3569), .ZN(n4737) );
  XNOR2_X1 U4457 ( .A(n3587), .B(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n4932) );
  AOI22_X1 U4458 ( .A1(n3949), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3973), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3574) );
  AOI22_X1 U4459 ( .A1(n3197), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3851), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3573) );
  AOI22_X1 U4460 ( .A1(n3852), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n3944), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3572) );
  AOI22_X1 U4461 ( .A1(n3859), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3157), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3571) );
  NAND4_X1 U4462 ( .A1(n3574), .A2(n3573), .A3(n3572), .A4(n3571), .ZN(n3580)
         );
  AOI22_X1 U4463 ( .A1(n3966), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3924), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3578) );
  AOI22_X1 U4464 ( .A1(n3925), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3879), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3577) );
  AOI22_X1 U4465 ( .A1(n3156), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n3878), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3576) );
  AOI22_X1 U4466 ( .A1(n3965), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3974), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3575) );
  NAND4_X1 U4467 ( .A1(n3578), .A2(n3577), .A3(n3576), .A4(n3575), .ZN(n3579)
         );
  NOR2_X1 U4468 ( .A1(n3580), .A2(n3579), .ZN(n3583) );
  NAND2_X1 U4469 ( .A1(n3987), .A2(EAX_REG_9__SCAN_IN), .ZN(n3582) );
  NAND2_X1 U4470 ( .A1(n3899), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3581)
         );
  OAI211_X1 U4471 ( .C1(n3682), .C2(n3583), .A(n3582), .B(n3581), .ZN(n3584)
         );
  AOI21_X1 U4472 ( .B1(n4932), .B2(n3993), .A(n3584), .ZN(n4808) );
  INV_X1 U4473 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n6534) );
  NAND2_X1 U4474 ( .A1(n3587), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3588)
         );
  AOI21_X1 U4475 ( .B1(n6534), .B2(n3588), .A(n3618), .ZN(n5824) );
  OR2_X1 U4476 ( .A1(n5824), .A2(n4123), .ZN(n3604) );
  AOI22_X1 U4477 ( .A1(n3973), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3925), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3592) );
  AOI22_X1 U4478 ( .A1(n3966), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3971), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3591) );
  AOI22_X1 U4479 ( .A1(n3197), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3944), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3590) );
  AOI22_X1 U4480 ( .A1(n3156), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n3974), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3589) );
  NAND4_X1 U4481 ( .A1(n3592), .A2(n3591), .A3(n3590), .A4(n3589), .ZN(n3598)
         );
  AOI22_X1 U4482 ( .A1(n3965), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3859), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3596) );
  AOI22_X1 U4483 ( .A1(n3949), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3879), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3595) );
  AOI22_X1 U4484 ( .A1(n3963), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3878), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3594) );
  AOI22_X1 U4485 ( .A1(n3852), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n2966), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3593) );
  NAND4_X1 U4486 ( .A1(n3596), .A2(n3595), .A3(n3594), .A4(n3593), .ZN(n3597)
         );
  NOR2_X1 U4487 ( .A1(n3598), .A2(n3597), .ZN(n3601) );
  NAND2_X1 U4488 ( .A1(n3987), .A2(EAX_REG_10__SCAN_IN), .ZN(n3600) );
  NAND2_X1 U4489 ( .A1(n3899), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3599)
         );
  OAI211_X1 U4490 ( .C1(n3682), .C2(n3601), .A(n3600), .B(n3599), .ZN(n3602)
         );
  INV_X1 U4491 ( .A(n3602), .ZN(n3603) );
  AND2_X1 U4492 ( .A1(n3604), .A2(n3603), .ZN(n4918) );
  AOI22_X1 U4493 ( .A1(n3973), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3924), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3608) );
  AOI22_X1 U4494 ( .A1(n3197), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3949), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3607) );
  AOI22_X1 U4495 ( .A1(n3878), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3974), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3606) );
  AOI22_X1 U4496 ( .A1(n3965), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3157), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3605) );
  NAND4_X1 U4497 ( .A1(n3608), .A2(n3607), .A3(n3606), .A4(n3605), .ZN(n3614)
         );
  AOI22_X1 U4498 ( .A1(n3966), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3851), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3612) );
  AOI22_X1 U4499 ( .A1(n3852), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3859), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3611) );
  AOI22_X1 U4500 ( .A1(n3036), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n3944), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3610) );
  AOI22_X1 U4501 ( .A1(n3925), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3879), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3609) );
  NAND4_X1 U4502 ( .A1(n3612), .A2(n3611), .A3(n3610), .A4(n3609), .ZN(n3613)
         );
  NOR2_X1 U4503 ( .A1(n3614), .A2(n3613), .ZN(n3617) );
  XNOR2_X1 U4504 ( .A(n3618), .B(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n5347)
         );
  NAND2_X1 U4505 ( .A1(n5347), .A2(n3993), .ZN(n3616) );
  AOI22_X1 U4506 ( .A1(n3987), .A2(EAX_REG_11__SCAN_IN), .B1(n3899), .B2(
        PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3615) );
  OAI211_X1 U4507 ( .C1(n3617), .C2(n3682), .A(n3616), .B(n3615), .ZN(n4936)
         );
  INV_X1 U4508 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n5808) );
  NAND2_X1 U4509 ( .A1(n3618), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3633)
         );
  XOR2_X1 U4510 ( .A(n5808), .B(n3633), .Z(n5812) );
  INV_X1 U4511 ( .A(n5812), .ZN(n5027) );
  AOI22_X1 U4512 ( .A1(n3966), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3949), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3622) );
  AOI22_X1 U4513 ( .A1(INSTQUEUE_REG_12__4__SCAN_IN), .A2(n3197), .B1(n3156), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3621) );
  AOI22_X1 U4514 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n3925), .B1(n3879), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3620) );
  AOI22_X1 U4515 ( .A1(n3965), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n2966), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3619) );
  NAND4_X1 U4516 ( .A1(n3622), .A2(n3621), .A3(n3620), .A4(n3619), .ZN(n3628)
         );
  AOI22_X1 U4517 ( .A1(INSTQUEUE_REG_15__4__SCAN_IN), .A2(n3971), .B1(n3973), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3626) );
  AOI22_X1 U4518 ( .A1(n3852), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n3944), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3625) );
  AOI22_X1 U4519 ( .A1(n3963), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3878), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3624) );
  AOI22_X1 U4520 ( .A1(n3859), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3974), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3623) );
  NAND4_X1 U4521 ( .A1(n3626), .A2(n3625), .A3(n3624), .A4(n3623), .ZN(n3627)
         );
  NOR2_X1 U4522 ( .A1(n3628), .A2(n3627), .ZN(n3631) );
  NAND2_X1 U4523 ( .A1(n3987), .A2(EAX_REG_12__SCAN_IN), .ZN(n3630) );
  NAND2_X1 U4524 ( .A1(n3899), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3629)
         );
  OAI211_X1 U4525 ( .C1(n3682), .C2(n3631), .A(n3630), .B(n3629), .ZN(n3632)
         );
  AOI21_X1 U4526 ( .B1(n5027), .B2(n3993), .A(n3632), .ZN(n4985) );
  INV_X1 U4527 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3649) );
  XNOR2_X1 U4528 ( .A(n3650), .B(n3649), .ZN(n5077) );
  AOI22_X1 U4529 ( .A1(n3197), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3973), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3637) );
  AOI22_X1 U4530 ( .A1(n3965), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3859), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3636) );
  AOI22_X1 U4531 ( .A1(n3852), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3944), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3635) );
  AOI22_X1 U4532 ( .A1(n2966), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3974), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3634) );
  NAND4_X1 U4533 ( .A1(n3637), .A2(n3636), .A3(n3635), .A4(n3634), .ZN(n3643)
         );
  AOI22_X1 U4534 ( .A1(n3966), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3971), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3641) );
  AOI22_X1 U4535 ( .A1(n3963), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3156), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3640) );
  AOI22_X1 U4536 ( .A1(n3925), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3853), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3639) );
  AOI22_X1 U4537 ( .A1(n3949), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3878), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3638) );
  NAND4_X1 U4538 ( .A1(n3641), .A2(n3640), .A3(n3639), .A4(n3638), .ZN(n3642)
         );
  NOR2_X1 U4539 ( .A1(n3643), .A2(n3642), .ZN(n3646) );
  NAND2_X1 U4540 ( .A1(n3987), .A2(EAX_REG_13__SCAN_IN), .ZN(n3645) );
  NAND2_X1 U4541 ( .A1(n3899), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3644)
         );
  OAI211_X1 U4542 ( .C1(n3682), .C2(n3646), .A(n3645), .B(n3644), .ZN(n3647)
         );
  AOI21_X1 U4543 ( .B1(n5077), .B2(n3993), .A(n3647), .ZN(n5034) );
  XOR2_X1 U4544 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .B(n3665), .Z(n5801) );
  AOI22_X1 U4545 ( .A1(n3973), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n3925), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3654) );
  AOI22_X1 U4546 ( .A1(n3966), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3851), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3653) );
  AOI22_X1 U4547 ( .A1(n3156), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n3944), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3652) );
  AOI22_X1 U4548 ( .A1(n3965), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3974), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3651) );
  NAND4_X1 U4549 ( .A1(n3654), .A2(n3653), .A3(n3652), .A4(n3651), .ZN(n3660)
         );
  AOI22_X1 U4550 ( .A1(n3197), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3949), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3658) );
  AOI22_X1 U4551 ( .A1(n3971), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n3853), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3657) );
  AOI22_X1 U4552 ( .A1(n3852), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3878), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3656) );
  AOI22_X1 U4553 ( .A1(n3859), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3157), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3655) );
  NAND4_X1 U4554 ( .A1(n3658), .A2(n3657), .A3(n3656), .A4(n3655), .ZN(n3659)
         );
  OR2_X1 U4555 ( .A1(n3660), .A2(n3659), .ZN(n3661) );
  AOI22_X1 U4556 ( .A1(n3662), .A2(n3661), .B1(n3899), .B2(
        PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n3664) );
  NAND2_X1 U4557 ( .A1(n3987), .A2(EAX_REG_14__SCAN_IN), .ZN(n3663) );
  OAI211_X1 U4558 ( .C1(n5801), .C2(n4123), .A(n3664), .B(n3663), .ZN(n5049)
         );
  NAND2_X1 U4559 ( .A1(n5050), .A2(n5049), .ZN(n5051) );
  NAND2_X1 U4560 ( .A1(n3665), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n3666)
         );
  INV_X1 U4561 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n6605) );
  NAND2_X1 U4562 ( .A1(n3666), .A2(n6605), .ZN(n3668) );
  INV_X1 U4563 ( .A(n3713), .ZN(n3667) );
  NAND2_X1 U4564 ( .A1(n3668), .A2(n3667), .ZN(n5141) );
  AOI22_X1 U4565 ( .A1(n3197), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3949), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3672) );
  AOI22_X1 U4566 ( .A1(n3965), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3859), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3671) );
  AOI22_X1 U4567 ( .A1(n3971), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n3925), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3670) );
  AOI22_X1 U4568 ( .A1(n3156), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n3157), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3669) );
  NAND4_X1 U4569 ( .A1(n3672), .A2(n3671), .A3(n3670), .A4(n3669), .ZN(n3678)
         );
  AOI22_X1 U4570 ( .A1(n3963), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3944), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3676) );
  AOI22_X1 U4571 ( .A1(n3966), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3878), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3675) );
  AOI22_X1 U4572 ( .A1(n3973), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n3853), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3674) );
  AOI22_X1 U4573 ( .A1(n3852), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3974), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3673) );
  NAND4_X1 U4574 ( .A1(n3676), .A2(n3675), .A3(n3674), .A4(n3673), .ZN(n3677)
         );
  NOR2_X1 U4575 ( .A1(n3678), .A2(n3677), .ZN(n3681) );
  NAND2_X1 U4576 ( .A1(n3987), .A2(EAX_REG_15__SCAN_IN), .ZN(n3680) );
  NAND2_X1 U4577 ( .A1(n3899), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3679)
         );
  OAI211_X1 U4578 ( .C1(n3682), .C2(n3681), .A(n3680), .B(n3679), .ZN(n3683)
         );
  AOI21_X1 U4579 ( .B1(n5141), .B2(n3993), .A(n3683), .ZN(n5055) );
  OR2_X2 U4580 ( .A1(n5051), .A2(n5055), .ZN(n5111) );
  NOR2_X1 U4581 ( .A1(n3684), .A2(n6382), .ZN(n3956) );
  AOI22_X1 U4582 ( .A1(n3973), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n3924), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3688) );
  AOI22_X1 U4583 ( .A1(n3283), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n3156), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3687) );
  AOI22_X1 U4584 ( .A1(n3965), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n2964), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3686) );
  AOI22_X1 U4585 ( .A1(n3925), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3853), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3685) );
  NAND4_X1 U4586 ( .A1(n3688), .A2(n3687), .A3(n3686), .A4(n3685), .ZN(n3694)
         );
  AOI22_X1 U4587 ( .A1(n3966), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3949), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3692) );
  AOI22_X1 U4588 ( .A1(n3963), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n3878), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3691) );
  AOI22_X1 U4589 ( .A1(n3859), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3157), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3690) );
  AOI22_X1 U4590 ( .A1(n3858), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3198), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3689) );
  NAND4_X1 U4591 ( .A1(n3692), .A2(n3691), .A3(n3690), .A4(n3689), .ZN(n3693)
         );
  OR2_X1 U4592 ( .A1(n3694), .A2(n3693), .ZN(n3698) );
  INV_X1 U4593 ( .A(EAX_REG_16__SCAN_IN), .ZN(n3696) );
  XOR2_X1 U4594 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .B(n3713), .Z(n5120) );
  INV_X1 U4595 ( .A(n5120), .ZN(n5168) );
  AOI22_X1 U4596 ( .A1(n3993), .A2(n5168), .B1(n3899), .B2(
        PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3695) );
  OAI21_X1 U4597 ( .B1(n3998), .B2(n3696), .A(n3695), .ZN(n3697) );
  AOI21_X1 U4598 ( .B1(n3956), .B2(n3698), .A(n3697), .ZN(n5112) );
  NOR2_X2 U4599 ( .A1(n5111), .A2(n5112), .ZN(n3699) );
  INV_X1 U4600 ( .A(n3699), .ZN(n5128) );
  INV_X1 U4601 ( .A(n3956), .ZN(n3989) );
  AOI22_X1 U4602 ( .A1(n3973), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n3971), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3703) );
  AOI22_X1 U4603 ( .A1(n3966), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3949), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3702) );
  AOI22_X1 U4604 ( .A1(n3925), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3853), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3701) );
  AOI22_X1 U4605 ( .A1(n3283), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3043), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3700) );
  NAND4_X1 U4606 ( .A1(n3703), .A2(n3702), .A3(n3701), .A4(n3700), .ZN(n3709)
         );
  AOI22_X1 U4607 ( .A1(n3852), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3156), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3707) );
  AOI22_X1 U4608 ( .A1(n3965), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3859), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3706) );
  AOI22_X1 U4609 ( .A1(n3963), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3858), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3705) );
  INV_X1 U4610 ( .A(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n6532) );
  AOI22_X1 U4611 ( .A1(n3157), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3198), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3704) );
  NAND4_X1 U4612 ( .A1(n3707), .A2(n3706), .A3(n3705), .A4(n3704), .ZN(n3708)
         );
  NOR2_X1 U4613 ( .A1(n3709), .A2(n3708), .ZN(n3712) );
  INV_X1 U4614 ( .A(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5534) );
  AOI21_X1 U4615 ( .B1(n5534), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3710) );
  AOI21_X1 U4616 ( .B1(n3987), .B2(EAX_REG_17__SCAN_IN), .A(n3710), .ZN(n3711)
         );
  OAI21_X1 U4617 ( .B1(n3989), .B2(n3712), .A(n3711), .ZN(n3715) );
  NAND2_X1 U4618 ( .A1(n3713), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3730)
         );
  XNOR2_X1 U4619 ( .A(PHYADDRPOINTER_REG_17__SCAN_IN), .B(n3730), .ZN(n5537)
         );
  NAND2_X1 U4620 ( .A1(n3993), .A2(n5537), .ZN(n3714) );
  NAND2_X1 U4621 ( .A1(n3715), .A2(n3714), .ZN(n5127) );
  NOR2_X2 U4622 ( .A1(n5128), .A2(n5127), .ZN(n5129) );
  AOI22_X1 U4623 ( .A1(n3966), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3949), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3719) );
  AOI22_X1 U4624 ( .A1(n3283), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3156), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3718) );
  AOI22_X1 U4625 ( .A1(n3973), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n3925), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3717) );
  AOI22_X1 U4626 ( .A1(n2966), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3198), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3716) );
  NAND4_X1 U4627 ( .A1(n3719), .A2(n3718), .A3(n3717), .A4(n3716), .ZN(n3725)
         );
  AOI22_X1 U4628 ( .A1(n3965), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3964), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3723) );
  AOI22_X1 U4629 ( .A1(n3852), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3858), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3722) );
  AOI22_X1 U4630 ( .A1(n3963), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3043), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3721) );
  AOI22_X1 U4631 ( .A1(n3971), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3853), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3720) );
  NAND4_X1 U4632 ( .A1(n3723), .A2(n3722), .A3(n3721), .A4(n3720), .ZN(n3724)
         );
  NOR2_X1 U4633 ( .A1(n3725), .A2(n3724), .ZN(n3729) );
  NAND2_X1 U4634 ( .A1(n6379), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n3726)
         );
  NAND2_X1 U4635 ( .A1(n4123), .A2(n3726), .ZN(n3727) );
  AOI21_X1 U4636 ( .B1(n3987), .B2(EAX_REG_18__SCAN_IN), .A(n3727), .ZN(n3728)
         );
  OAI21_X1 U4637 ( .B1(n3989), .B2(n3729), .A(n3728), .ZN(n3733) );
  OAI21_X1 U4638 ( .B1(PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n3731), .A(n3870), 
        .ZN(n5791) );
  OR2_X1 U4639 ( .A1(n4123), .A2(n5791), .ZN(n3732) );
  AND2_X1 U4640 ( .A1(n3733), .A2(n3732), .ZN(n5422) );
  AOI22_X1 U4641 ( .A1(n3973), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3971), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3737) );
  AOI22_X1 U4642 ( .A1(n3966), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3949), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3736) );
  AOI22_X1 U4643 ( .A1(n3925), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3853), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3735) );
  AOI22_X1 U4644 ( .A1(n3283), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3878), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3734) );
  NAND4_X1 U4645 ( .A1(n3737), .A2(n3736), .A3(n3735), .A4(n3734), .ZN(n3743)
         );
  AOI22_X1 U4646 ( .A1(n3852), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3156), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3741) );
  AOI22_X1 U4647 ( .A1(n3965), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3859), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3740) );
  AOI22_X1 U4648 ( .A1(n3963), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n3858), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3739) );
  AOI22_X1 U4649 ( .A1(n2966), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3974), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3738) );
  NAND4_X1 U4650 ( .A1(n3741), .A2(n3740), .A3(n3739), .A4(n3738), .ZN(n3742)
         );
  NOR2_X1 U4651 ( .A1(n3743), .A2(n3742), .ZN(n3802) );
  AOI22_X1 U4652 ( .A1(n3197), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n3851), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3747) );
  AOI22_X1 U4653 ( .A1(n3949), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3879), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3746) );
  AOI22_X1 U4654 ( .A1(n3859), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n2966), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3745) );
  AOI22_X1 U4655 ( .A1(n3852), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n3974), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3744) );
  NAND4_X1 U4656 ( .A1(n3747), .A2(n3746), .A3(n3745), .A4(n3744), .ZN(n3753)
         );
  AOI22_X1 U4657 ( .A1(n3966), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3924), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3751) );
  AOI22_X1 U4658 ( .A1(n3965), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n3156), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3750) );
  AOI22_X1 U4659 ( .A1(n3973), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n3925), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3749) );
  AOI22_X1 U4660 ( .A1(n3858), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3878), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3748) );
  NAND4_X1 U4661 ( .A1(n3751), .A2(n3750), .A3(n3749), .A4(n3748), .ZN(n3752)
         );
  NOR2_X1 U4662 ( .A1(n3753), .A2(n3752), .ZN(n3812) );
  AOI22_X1 U4663 ( .A1(n3851), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3944), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3757) );
  AOI22_X1 U4664 ( .A1(n3971), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n3879), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3756) );
  AOI22_X1 U4665 ( .A1(n3197), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3878), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3755) );
  AOI22_X1 U4666 ( .A1(n3036), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n2966), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3754) );
  NAND4_X1 U4667 ( .A1(n3757), .A2(n3756), .A3(n3755), .A4(n3754), .ZN(n3763)
         );
  AOI22_X1 U4668 ( .A1(n3966), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3061), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3761) );
  AOI22_X1 U4669 ( .A1(n3965), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3859), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3760) );
  AOI22_X1 U4670 ( .A1(n3973), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3925), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3759) );
  AOI22_X1 U4671 ( .A1(n2964), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3974), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3758) );
  NAND4_X1 U4672 ( .A1(n3761), .A2(n3760), .A3(n3759), .A4(n3758), .ZN(n3762)
         );
  NOR2_X1 U4673 ( .A1(n3763), .A2(n3762), .ZN(n3811) );
  OR2_X1 U4674 ( .A1(n3812), .A2(n3811), .ZN(n3897) );
  AOI22_X1 U4675 ( .A1(n2964), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3036), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3767) );
  AOI22_X1 U4676 ( .A1(n3965), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3973), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3766) );
  AOI22_X1 U4677 ( .A1(n3859), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3971), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3765) );
  AOI22_X1 U4678 ( .A1(n3157), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3974), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3764) );
  NAND4_X1 U4679 ( .A1(n3767), .A2(n3766), .A3(n3765), .A4(n3764), .ZN(n3773)
         );
  AOI22_X1 U4680 ( .A1(n3966), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3061), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3771) );
  AOI22_X1 U4681 ( .A1(n3197), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3944), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3770) );
  AOI22_X1 U4682 ( .A1(n3925), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3878), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3769) );
  AOI22_X1 U4683 ( .A1(n3851), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n3879), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3768) );
  NAND4_X1 U4684 ( .A1(n3771), .A2(n3770), .A3(n3769), .A4(n3768), .ZN(n3772)
         );
  NOR2_X1 U4685 ( .A1(n3773), .A2(n3772), .ZN(n3895) );
  OR2_X1 U4686 ( .A1(n3897), .A2(n3895), .ZN(n3801) );
  NOR2_X1 U4687 ( .A1(n3802), .A2(n3801), .ZN(n3908) );
  AOI22_X1 U4688 ( .A1(n2963), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3036), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3777) );
  AOI22_X1 U4689 ( .A1(n3965), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3859), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3776) );
  AOI22_X1 U4690 ( .A1(n3963), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n3944), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3775) );
  AOI22_X1 U4691 ( .A1(n2966), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3198), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3774) );
  NAND4_X1 U4692 ( .A1(n3777), .A2(n3776), .A3(n3775), .A4(n3774), .ZN(n3783)
         );
  AOI22_X1 U4693 ( .A1(n3973), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3924), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3781) );
  AOI22_X1 U4694 ( .A1(n3966), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3061), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3780) );
  AOI22_X1 U4695 ( .A1(n3925), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3879), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3779) );
  AOI22_X1 U4696 ( .A1(n3283), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3878), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3778) );
  NAND4_X1 U4697 ( .A1(n3781), .A2(n3780), .A3(n3779), .A4(n3778), .ZN(n3782)
         );
  OR2_X1 U4698 ( .A1(n3783), .A2(n3782), .ZN(n3906) );
  NAND2_X1 U4699 ( .A1(n3908), .A2(n3906), .ZN(n3918) );
  AOI22_X1 U4700 ( .A1(INSTQUEUE_REG_14__4__SCAN_IN), .A2(n3197), .B1(n3966), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3787) );
  AOI22_X1 U4701 ( .A1(n3924), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n3972), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3786) );
  AOI22_X1 U4702 ( .A1(INSTQUEUE_REG_5__4__SCAN_IN), .A2(n3156), .B1(n3878), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3785) );
  AOI22_X1 U4703 ( .A1(n3965), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3198), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3784) );
  NAND4_X1 U4704 ( .A1(n3787), .A2(n3786), .A3(n3785), .A4(n3784), .ZN(n3793)
         );
  AOI22_X1 U4705 ( .A1(INSTQUEUE_REG_2__4__SCAN_IN), .A2(n3973), .B1(n3925), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3791) );
  AOI22_X1 U4706 ( .A1(n3963), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n3061), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3790) );
  AOI22_X1 U4707 ( .A1(n2963), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3944), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3789) );
  AOI22_X1 U4708 ( .A1(n3859), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n2966), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3788) );
  NAND4_X1 U4709 ( .A1(n3791), .A2(n3790), .A3(n3789), .A4(n3788), .ZN(n3792)
         );
  NOR2_X1 U4710 ( .A1(n3793), .A2(n3792), .ZN(n3919) );
  XOR2_X1 U4711 ( .A(n3918), .B(n3919), .Z(n3794) );
  NAND2_X1 U4712 ( .A1(n3794), .A2(n3956), .ZN(n3800) );
  INV_X1 U4713 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5309) );
  OAI21_X1 U4714 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n5309), .A(n4123), .ZN(
        n3795) );
  AOI21_X1 U4715 ( .B1(n3987), .B2(EAX_REG_27__SCAN_IN), .A(n3795), .ZN(n3799)
         );
  INV_X1 U4716 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n5702) );
  XNOR2_X1 U4717 ( .A(n3936), .B(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5307)
         );
  AND2_X1 U4718 ( .A1(n5307), .A2(n3993), .ZN(n3798) );
  AOI21_X1 U4719 ( .B1(n3800), .B2(n3799), .A(n3798), .ZN(n5230) );
  XOR2_X1 U4720 ( .A(n3802), .B(n3801), .Z(n3806) );
  INV_X1 U4721 ( .A(EAX_REG_25__SCAN_IN), .ZN(n3804) );
  NAND2_X1 U4722 ( .A1(n6379), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n3803)
         );
  OAI211_X1 U4723 ( .C1(n3998), .C2(n3804), .A(n4123), .B(n3803), .ZN(n3805)
         );
  AOI21_X1 U4724 ( .B1(n3806), .B2(n3956), .A(n3805), .ZN(n3807) );
  INV_X1 U4725 ( .A(n3807), .ZN(n3810) );
  XNOR2_X1 U4726 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .B(n3808), .ZN(n5672)
         );
  NAND2_X1 U4727 ( .A1(n3993), .A2(n5672), .ZN(n3809) );
  AND2_X1 U4728 ( .A1(n3810), .A2(n3809), .ZN(n5380) );
  XOR2_X1 U4729 ( .A(n3812), .B(n3811), .Z(n3813) );
  NAND2_X1 U4730 ( .A1(n3813), .A2(n3956), .ZN(n3817) );
  INV_X1 U4731 ( .A(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5490) );
  AOI21_X1 U4732 ( .B1(n5490), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3814) );
  AOI21_X1 U4733 ( .B1(n3987), .B2(EAX_REG_23__SCAN_IN), .A(n3814), .ZN(n3816)
         );
  XNOR2_X1 U4734 ( .A(n3892), .B(n5490), .ZN(n5488) );
  AND2_X1 U4735 ( .A1(n5488), .A2(n3993), .ZN(n3815) );
  AOI21_X1 U4736 ( .B1(n3817), .B2(n3816), .A(n3815), .ZN(n5314) );
  AOI22_X1 U4737 ( .A1(n3973), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3924), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3821) );
  AOI22_X1 U4738 ( .A1(n3197), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3966), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3820) );
  AOI22_X1 U4739 ( .A1(n3965), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n2963), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3819) );
  AOI22_X1 U4740 ( .A1(n3963), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3944), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3818) );
  NAND4_X1 U4741 ( .A1(n3821), .A2(n3820), .A3(n3819), .A4(n3818), .ZN(n3827)
         );
  AOI22_X1 U4742 ( .A1(n3925), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3853), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3825) );
  AOI22_X1 U4743 ( .A1(n3949), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3878), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3824) );
  AOI22_X1 U4744 ( .A1(n3859), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3157), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3823) );
  AOI22_X1 U4745 ( .A1(n3156), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3974), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3822) );
  NAND4_X1 U4746 ( .A1(n3825), .A2(n3824), .A3(n3823), .A4(n3822), .ZN(n3826)
         );
  NOR2_X1 U4747 ( .A1(n3827), .A2(n3826), .ZN(n3830) );
  OAI21_X1 U4748 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n5702), .A(n4123), .ZN(
        n3828) );
  AOI21_X1 U4749 ( .B1(n3987), .B2(EAX_REG_21__SCAN_IN), .A(n3828), .ZN(n3829)
         );
  OAI21_X1 U4750 ( .B1(n3989), .B2(n3830), .A(n3829), .ZN(n3832) );
  XNOR2_X1 U4751 ( .A(n3847), .B(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n5700)
         );
  NAND2_X1 U4752 ( .A1(n5700), .A2(n3993), .ZN(n3831) );
  NAND2_X1 U4753 ( .A1(n3832), .A2(n3831), .ZN(n5399) );
  AOI22_X1 U4754 ( .A1(n3197), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3971), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3836) );
  AOI22_X1 U4755 ( .A1(INSTQUEUE_REG_12__4__SCAN_IN), .A2(n3965), .B1(n3859), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3835) );
  AOI22_X1 U4756 ( .A1(n3973), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n3853), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3834) );
  AOI22_X1 U4757 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n3858), .B1(n2966), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3833) );
  NAND4_X1 U4758 ( .A1(n3836), .A2(n3835), .A3(n3834), .A4(n3833), .ZN(n3842)
         );
  AOI22_X1 U4759 ( .A1(n3963), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3156), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3840) );
  AOI22_X1 U4760 ( .A1(n3966), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3925), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3839) );
  AOI22_X1 U4761 ( .A1(INSTQUEUE_REG_8__4__SCAN_IN), .A2(n3949), .B1(n3878), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3838) );
  AOI22_X1 U4762 ( .A1(n3852), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3974), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3837) );
  NAND4_X1 U4763 ( .A1(n3840), .A2(n3839), .A3(n3838), .A4(n3837), .ZN(n3841)
         );
  NOR2_X1 U4764 ( .A1(n3842), .A2(n3841), .ZN(n3846) );
  NAND2_X1 U4765 ( .A1(n6379), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n3843)
         );
  NAND2_X1 U4766 ( .A1(n4123), .A2(n3843), .ZN(n3844) );
  AOI21_X1 U4767 ( .B1(n3987), .B2(EAX_REG_20__SCAN_IN), .A(n3844), .ZN(n3845)
         );
  OAI21_X1 U4768 ( .B1(n3989), .B2(n3846), .A(n3845), .ZN(n3850) );
  OAI21_X1 U4769 ( .B1(n3848), .B2(PHYADDRPOINTER_REG_20__SCAN_IN), .A(n3847), 
        .ZN(n5710) );
  OR2_X1 U4770 ( .A1(n5710), .A2(n4123), .ZN(n3849) );
  NAND2_X1 U4771 ( .A1(n3850), .A2(n3849), .ZN(n5408) );
  NOR2_X1 U4772 ( .A1(n5399), .A2(n5408), .ZN(n3873) );
  AOI22_X1 U4773 ( .A1(n3197), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3851), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3857) );
  AOI22_X1 U4774 ( .A1(n3852), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3156), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3856) );
  AOI22_X1 U4775 ( .A1(n3924), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3853), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3855) );
  AOI22_X1 U4776 ( .A1(n3965), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3974), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3854) );
  NAND4_X1 U4777 ( .A1(n3857), .A2(n3856), .A3(n3855), .A4(n3854), .ZN(n3865)
         );
  AOI22_X1 U4778 ( .A1(n3966), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3949), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3863) );
  AOI22_X1 U4779 ( .A1(n3973), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3925), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3862) );
  AOI22_X1 U4780 ( .A1(n3858), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3878), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3861) );
  AOI22_X1 U4781 ( .A1(n3859), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n2966), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3860) );
  NAND4_X1 U4782 ( .A1(n3863), .A2(n3862), .A3(n3861), .A4(n3860), .ZN(n3864)
         );
  NOR2_X1 U4783 ( .A1(n3865), .A2(n3864), .ZN(n3869) );
  NAND2_X1 U4784 ( .A1(n6379), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n3866)
         );
  NAND2_X1 U4785 ( .A1(n4123), .A2(n3866), .ZN(n3867) );
  AOI21_X1 U4786 ( .B1(n3987), .B2(EAX_REG_19__SCAN_IN), .A(n3867), .ZN(n3868)
         );
  OAI21_X1 U4787 ( .B1(n3989), .B2(n3869), .A(n3868), .ZN(n3872) );
  XNOR2_X1 U4788 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .B(n3870), .ZN(n5524)
         );
  NAND2_X1 U4789 ( .A1(n3993), .A2(n5524), .ZN(n3871) );
  AND2_X1 U4790 ( .A1(n3872), .A2(n3871), .ZN(n5327) );
  AND2_X1 U4791 ( .A1(n3873), .A2(n5327), .ZN(n5390) );
  AOI22_X1 U4792 ( .A1(n3973), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3971), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3877) );
  AOI22_X1 U4793 ( .A1(n3283), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3966), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3876) );
  AOI22_X1 U4794 ( .A1(n3852), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3156), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3875) );
  AOI22_X1 U4795 ( .A1(n3965), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3859), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3874) );
  NAND4_X1 U4796 ( .A1(n3877), .A2(n3876), .A3(n3875), .A4(n3874), .ZN(n3885)
         );
  AOI22_X1 U4797 ( .A1(n3963), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3944), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3883) );
  AOI22_X1 U4798 ( .A1(n3949), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3878), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3882) );
  AOI22_X1 U4799 ( .A1(n3925), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3879), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3881) );
  AOI22_X1 U4800 ( .A1(n2966), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3974), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3880) );
  NAND4_X1 U4801 ( .A1(n3883), .A2(n3882), .A3(n3881), .A4(n3880), .ZN(n3884)
         );
  NOR2_X1 U4802 ( .A1(n3885), .A2(n3884), .ZN(n3889) );
  NAND2_X1 U4803 ( .A1(n6379), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n3886)
         );
  NAND2_X1 U4804 ( .A1(n4123), .A2(n3886), .ZN(n3887) );
  AOI21_X1 U4805 ( .B1(n3987), .B2(EAX_REG_22__SCAN_IN), .A(n3887), .ZN(n3888)
         );
  OAI21_X1 U4806 ( .B1(n3989), .B2(n3889), .A(n3888), .ZN(n3894) );
  NOR2_X1 U4807 ( .A1(n3890), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n3891)
         );
  OR2_X1 U4808 ( .A1(n3892), .A2(n3891), .ZN(n5500) );
  INV_X1 U4809 ( .A(n5500), .ZN(n5693) );
  NAND2_X1 U4810 ( .A1(n5693), .A2(n3993), .ZN(n3893) );
  AND2_X1 U4811 ( .A1(n3894), .A2(n3893), .ZN(n5391) );
  AND2_X1 U4812 ( .A1(n5390), .A2(n5391), .ZN(n5313) );
  AND2_X1 U4813 ( .A1(n5314), .A2(n5313), .ZN(n5252) );
  INV_X1 U4814 ( .A(n3895), .ZN(n3896) );
  XNOR2_X1 U4815 ( .A(n3897), .B(n3896), .ZN(n3904) );
  INV_X1 U4816 ( .A(EAX_REG_24__SCAN_IN), .ZN(n3902) );
  XNOR2_X1 U4817 ( .A(n3898), .B(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5683)
         );
  NAND2_X1 U4818 ( .A1(n5683), .A2(n3993), .ZN(n3901) );
  NAND2_X1 U4819 ( .A1(n3899), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n3900)
         );
  OAI211_X1 U4820 ( .C1(n3998), .C2(n3902), .A(n3901), .B(n3900), .ZN(n3903)
         );
  AOI21_X1 U4821 ( .B1(n3904), .B2(n3956), .A(n3903), .ZN(n5255) );
  INV_X1 U4822 ( .A(n5255), .ZN(n3905) );
  AND2_X1 U4823 ( .A1(n5252), .A2(n3905), .ZN(n5253) );
  AND2_X1 U4824 ( .A1(n5380), .A2(n5253), .ZN(n5371) );
  INV_X1 U4825 ( .A(n3906), .ZN(n3907) );
  XNOR2_X1 U4826 ( .A(n3908), .B(n3907), .ZN(n3912) );
  INV_X1 U4827 ( .A(EAX_REG_26__SCAN_IN), .ZN(n3910) );
  NAND2_X1 U4828 ( .A1(n6379), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n3909)
         );
  OAI211_X1 U4829 ( .C1(n3998), .C2(n3910), .A(n4123), .B(n3909), .ZN(n3911)
         );
  AOI21_X1 U4830 ( .B1(n3912), .B2(n3956), .A(n3911), .ZN(n3915) );
  OAI21_X1 U4831 ( .B1(n3913), .B2(PHYADDRPOINTER_REG_26__SCAN_IN), .A(n3936), 
        .ZN(n5661) );
  NOR2_X1 U4832 ( .A1(n5661), .A2(n4123), .ZN(n3914) );
  OR2_X1 U4833 ( .A1(n3915), .A2(n3914), .ZN(n5372) );
  INV_X1 U4834 ( .A(n5372), .ZN(n3916) );
  AND2_X1 U4835 ( .A1(n5371), .A2(n3916), .ZN(n5229) );
  AND2_X1 U4836 ( .A1(n5230), .A2(n5229), .ZN(n3917) );
  NOR2_X1 U4837 ( .A1(n3919), .A2(n3918), .ZN(n3943) );
  AOI22_X1 U4838 ( .A1(n2964), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3036), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3923) );
  AOI22_X1 U4839 ( .A1(n3965), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3964), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3922) );
  AOI22_X1 U4840 ( .A1(n3963), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n3944), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3921) );
  AOI22_X1 U4841 ( .A1(n2966), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3198), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3920) );
  NAND4_X1 U4842 ( .A1(n3923), .A2(n3922), .A3(n3921), .A4(n3920), .ZN(n3931)
         );
  AOI22_X1 U4843 ( .A1(n3973), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3924), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3929) );
  AOI22_X1 U4844 ( .A1(n3966), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3061), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3928) );
  AOI22_X1 U4845 ( .A1(n3925), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3972), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3927) );
  AOI22_X1 U4846 ( .A1(n3197), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3878), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3926) );
  NAND4_X1 U4847 ( .A1(n3929), .A2(n3928), .A3(n3927), .A4(n3926), .ZN(n3930)
         );
  OR2_X1 U4848 ( .A1(n3931), .A2(n3930), .ZN(n3942) );
  INV_X1 U4849 ( .A(n3942), .ZN(n3932) );
  XNOR2_X1 U4850 ( .A(n3943), .B(n3932), .ZN(n3933) );
  NAND2_X1 U4851 ( .A1(n3933), .A2(n3956), .ZN(n3941) );
  NAND2_X1 U4852 ( .A1(n6379), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n3934)
         );
  NAND2_X1 U4853 ( .A1(n4123), .A2(n3934), .ZN(n3935) );
  AOI21_X1 U4854 ( .B1(n3987), .B2(EAX_REG_28__SCAN_IN), .A(n3935), .ZN(n3940)
         );
  NAND2_X1 U4855 ( .A1(n3937), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n3992)
         );
  OR2_X1 U4856 ( .A1(n3937), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n3938)
         );
  NAND2_X1 U4857 ( .A1(n3992), .A2(n3938), .ZN(n5650) );
  NOR2_X1 U4858 ( .A1(n5650), .A2(n4123), .ZN(n3939) );
  AOI21_X1 U4859 ( .B1(n3941), .B2(n3940), .A(n3939), .ZN(n5360) );
  AND2_X2 U4860 ( .A1(n5227), .A2(n5360), .ZN(n5362) );
  NAND2_X1 U4861 ( .A1(n3943), .A2(n3942), .ZN(n3981) );
  AOI22_X1 U4862 ( .A1(n3966), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3971), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3948) );
  AOI22_X1 U4863 ( .A1(n3156), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3944), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3947) );
  AOI22_X1 U4864 ( .A1(n3973), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3972), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3946) );
  AOI22_X1 U4865 ( .A1(n3852), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3157), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3945) );
  NAND4_X1 U4866 ( .A1(n3948), .A2(n3947), .A3(n3946), .A4(n3945), .ZN(n3955)
         );
  AOI22_X1 U4867 ( .A1(n3965), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3964), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3953) );
  AOI22_X1 U4868 ( .A1(n3949), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3925), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3952) );
  AOI22_X1 U4869 ( .A1(n3283), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3878), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3951) );
  AOI22_X1 U4870 ( .A1(n3963), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n3974), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3950) );
  NAND4_X1 U4871 ( .A1(n3953), .A2(n3952), .A3(n3951), .A4(n3950), .ZN(n3954)
         );
  NOR2_X1 U4872 ( .A1(n3955), .A2(n3954), .ZN(n3982) );
  XOR2_X1 U4873 ( .A(n3981), .B(n3982), .Z(n3957) );
  NAND2_X1 U4874 ( .A1(n3957), .A2(n3956), .ZN(n3962) );
  NAND2_X1 U4875 ( .A1(n6379), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n3958)
         );
  NAND2_X1 U4876 ( .A1(n4123), .A2(n3958), .ZN(n3959) );
  AOI21_X1 U4877 ( .B1(n3987), .B2(EAX_REG_29__SCAN_IN), .A(n3959), .ZN(n3961)
         );
  XNOR2_X1 U4878 ( .A(n3992), .B(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5643)
         );
  AND2_X1 U4879 ( .A1(n5643), .A2(n3993), .ZN(n3960) );
  AOI21_X1 U4880 ( .B1(n3962), .B2(n3961), .A(n3960), .ZN(n5173) );
  NAND2_X1 U4881 ( .A1(n5362), .A2(n5173), .ZN(n5174) );
  AOI22_X1 U4882 ( .A1(n3283), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3949), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3970) );
  AOI22_X1 U4883 ( .A1(n3963), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n2963), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3969) );
  AOI22_X1 U4884 ( .A1(n3965), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3964), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3968) );
  AOI22_X1 U4885 ( .A1(n3966), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3925), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3967) );
  NAND4_X1 U4886 ( .A1(n3970), .A2(n3969), .A3(n3968), .A4(n3967), .ZN(n3980)
         );
  AOI22_X1 U4887 ( .A1(n3156), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3858), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3978) );
  AOI22_X1 U4888 ( .A1(n3971), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3043), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3977) );
  AOI22_X1 U4889 ( .A1(n3973), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3972), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3976) );
  AOI22_X1 U4890 ( .A1(n2966), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3974), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3975) );
  NAND4_X1 U4891 ( .A1(n3978), .A2(n3977), .A3(n3976), .A4(n3975), .ZN(n3979)
         );
  NOR2_X1 U4892 ( .A1(n3980), .A2(n3979), .ZN(n3984) );
  NOR2_X1 U4893 ( .A1(n3982), .A2(n3981), .ZN(n3983) );
  XOR2_X1 U4894 ( .A(n3984), .B(n3983), .Z(n3990) );
  NAND2_X1 U4895 ( .A1(n6379), .A2(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n3985)
         );
  NAND2_X1 U4896 ( .A1(n4123), .A2(n3985), .ZN(n3986) );
  AOI21_X1 U4897 ( .B1(n3987), .B2(EAX_REG_30__SCAN_IN), .A(n3986), .ZN(n3988)
         );
  OAI21_X1 U4898 ( .B1(n3990), .B2(n3989), .A(n3988), .ZN(n3995) );
  INV_X1 U4899 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n3991) );
  XNOR2_X1 U4900 ( .A(n4004), .B(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n4156)
         );
  NAND2_X1 U4901 ( .A1(n4156), .A2(n3993), .ZN(n3994) );
  NAND2_X1 U4902 ( .A1(n3995), .A2(n3994), .ZN(n4153) );
  OR2_X2 U4903 ( .A1(n5174), .A2(n4153), .ZN(n4151) );
  INV_X1 U4904 ( .A(EAX_REG_31__SCAN_IN), .ZN(n5434) );
  INV_X1 U4905 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n3996) );
  OAI22_X1 U4906 ( .A1(n3998), .A2(n5434), .B1(n3997), .B2(n3996), .ZN(n3999)
         );
  NAND3_X1 U4907 ( .A1(n6382), .A2(STATEBS16_REG_SCAN_IN), .A3(
        STATE2_REG_1__SCAN_IN), .ZN(n6395) );
  INV_X1 U4908 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n6470) );
  NAND2_X1 U4909 ( .A1(n6470), .A2(n6379), .ZN(n6286) );
  OR2_X1 U4910 ( .A1(n6395), .A2(n6286), .ZN(n5542) );
  INV_X1 U4911 ( .A(n6286), .ZN(n6197) );
  OR2_X1 U4912 ( .A1(n4000), .A2(n6197), .ZN(n6491) );
  NAND2_X1 U4913 ( .A1(n6491), .A2(n6382), .ZN(n4001) );
  NAND2_X1 U4914 ( .A1(n6382), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4003) );
  NAND2_X1 U4915 ( .A1(n6234), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4002) );
  AND2_X1 U4916 ( .A1(n4003), .A2(n4002), .ZN(n4304) );
  INV_X1 U4917 ( .A(n4004), .ZN(n4005) );
  NAND2_X1 U4918 ( .A1(n4005), .A2(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n4006)
         );
  XNOR2_X1 U4919 ( .A(n4006), .B(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4154)
         );
  INV_X1 U4920 ( .A(n4154), .ZN(n4008) );
  NOR2_X1 U4921 ( .A1(n6286), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4923) );
  INV_X1 U4922 ( .A(REIP_REG_31__SCAN_IN), .ZN(n6462) );
  NOR2_X1 U4923 ( .A1(n6047), .A2(n6462), .ZN(n5197) );
  AOI21_X1 U4924 ( .B1(n5963), .B2(PHYADDRPOINTER_REG_31__SCAN_IN), .A(n5197), 
        .ZN(n4007) );
  OAI21_X1 U4925 ( .B1(n5973), .B2(n4008), .A(n4007), .ZN(n4009) );
  NAND2_X1 U4926 ( .A1(n4011), .A2(n4010), .ZN(U2955) );
  OR2_X2 U4927 ( .A1(n4043), .A2(n4110), .ZN(n4091) );
  OR2_X2 U4928 ( .A1(n4013), .A2(n4220), .ZN(n4103) );
  NAND2_X1 U4929 ( .A1(n4103), .A2(n5149), .ZN(n4014) );
  OAI211_X1 U4930 ( .C1(n4043), .C2(EBX_REG_1__SCAN_IN), .A(n4110), .B(n4014), 
        .ZN(n4015) );
  NAND2_X1 U4931 ( .A1(n4103), .A2(EBX_REG_0__SCAN_IN), .ZN(n4017) );
  INV_X1 U4932 ( .A(EBX_REG_0__SCAN_IN), .ZN(n6652) );
  NAND2_X1 U4933 ( .A1(n4110), .A2(n6652), .ZN(n4016) );
  NAND2_X1 U4934 ( .A1(n4017), .A2(n4016), .ZN(n4308) );
  XNOR2_X1 U4935 ( .A(n4018), .B(n4308), .ZN(n5013) );
  NAND2_X1 U4936 ( .A1(n4318), .A2(n4018), .ZN(n4481) );
  INV_X1 U4937 ( .A(EBX_REG_2__SCAN_IN), .ZN(n4022) );
  NAND2_X1 U4938 ( .A1(n4103), .A2(n5964), .ZN(n4019) );
  OAI211_X1 U4939 ( .C1(n4043), .C2(EBX_REG_2__SCAN_IN), .A(n4110), .B(n4019), 
        .ZN(n4020) );
  NAND2_X1 U4940 ( .A1(n4219), .A2(n6038), .ZN(n4028) );
  INV_X1 U4941 ( .A(EBX_REG_3__SCAN_IN), .ZN(n4024) );
  NAND2_X1 U4942 ( .A1(n4100), .A2(n4024), .ZN(n4026) );
  NAND2_X1 U4943 ( .A1(n4208), .A2(EBX_REG_3__SCAN_IN), .ZN(n4025) );
  INV_X1 U4944 ( .A(EBX_REG_4__SCAN_IN), .ZN(n4033) );
  NAND2_X1 U4945 ( .A1(n4334), .A2(n4033), .ZN(n4032) );
  AOI21_X1 U4946 ( .B1(n4103), .B2(n6031), .A(n4208), .ZN(n4031) );
  AOI22_X1 U4947 ( .A1(n4107), .A2(n4033), .B1(n4032), .B2(n4031), .ZN(n4554)
         );
  INV_X1 U4948 ( .A(EBX_REG_5__SCAN_IN), .ZN(n4613) );
  MUX2_X1 U4949 ( .A(n4208), .B(n4100), .S(n4613), .Z(n4035) );
  NOR2_X1 U4950 ( .A1(n4309), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4034)
         );
  NOR2_X1 U4951 ( .A1(n4035), .A2(n4034), .ZN(n4609) );
  NAND2_X1 U4952 ( .A1(n4610), .A2(n4609), .ZN(n4608) );
  INV_X1 U4953 ( .A(n4608), .ZN(n4039) );
  INV_X1 U4954 ( .A(EBX_REG_6__SCAN_IN), .ZN(n6633) );
  NAND2_X1 U4955 ( .A1(n4334), .A2(n6633), .ZN(n4037) );
  AOI21_X1 U4956 ( .B1(n4103), .B2(n4240), .A(n4208), .ZN(n4036) );
  AOI22_X1 U4957 ( .A1(n4107), .A2(n6633), .B1(n4037), .B2(n4036), .ZN(n4565)
         );
  NAND2_X1 U4958 ( .A1(n4039), .A2(n4038), .ZN(n4564) );
  MUX2_X1 U4959 ( .A(n4100), .B(n4208), .S(EBX_REG_7__SCAN_IN), .Z(n4040) );
  INV_X1 U4960 ( .A(n4040), .ZN(n4041) );
  NAND2_X1 U4961 ( .A1(n4041), .A2(n2977), .ZN(n4750) );
  NOR2_X2 U4962 ( .A1(n4564), .A2(n4750), .ZN(n4740) );
  NAND2_X1 U4963 ( .A1(n4103), .A2(n6006), .ZN(n4042) );
  OAI211_X1 U4964 ( .C1(n4043), .C2(EBX_REG_8__SCAN_IN), .A(n4110), .B(n4042), 
        .ZN(n4044) );
  OAI21_X1 U4965 ( .B1(n4091), .B2(EBX_REG_8__SCAN_IN), .A(n4044), .ZN(n4741)
         );
  INV_X1 U4966 ( .A(EBX_REG_9__SCAN_IN), .ZN(n4855) );
  MUX2_X1 U4967 ( .A(n4208), .B(n4100), .S(n4855), .Z(n4046) );
  NOR2_X1 U4968 ( .A1(n4309), .A2(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n4045)
         );
  NOR2_X1 U4969 ( .A1(n4046), .A2(n4045), .ZN(n4850) );
  NAND2_X1 U4970 ( .A1(n4739), .A2(n4850), .ZN(n4851) );
  MUX2_X1 U4971 ( .A(n4091), .B(n4103), .S(EBX_REG_10__SCAN_IN), .Z(n4050) );
  INV_X1 U4972 ( .A(n4103), .ZN(n4047) );
  NAND2_X1 U4973 ( .A1(n4047), .A2(n4202), .ZN(n4085) );
  NAND2_X1 U4974 ( .A1(INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n4202), .ZN(n4048) );
  AND2_X1 U4975 ( .A1(n4085), .A2(n4048), .ZN(n4049) );
  NAND2_X1 U4976 ( .A1(n4050), .A2(n4049), .ZN(n4933) );
  INV_X1 U4977 ( .A(n4933), .ZN(n4051) );
  OR2_X2 U4978 ( .A1(n4851), .A2(n4051), .ZN(n4939) );
  INV_X1 U4979 ( .A(n4100), .ZN(n4090) );
  NAND2_X1 U4980 ( .A1(n4110), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n4052) );
  OAI211_X1 U4981 ( .C1(n4202), .C2(EBX_REG_11__SCAN_IN), .A(n4103), .B(n4052), 
        .ZN(n4053) );
  OAI21_X1 U4982 ( .B1(n4090), .B2(EBX_REG_11__SCAN_IN), .A(n4053), .ZN(n4940)
         );
  MUX2_X1 U4983 ( .A(n4091), .B(n4103), .S(EBX_REG_12__SCAN_IN), .Z(n4056) );
  NAND2_X1 U4984 ( .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n4202), .ZN(n4054) );
  AND2_X1 U4985 ( .A1(n4085), .A2(n4054), .ZN(n4055) );
  NAND2_X1 U4986 ( .A1(n4056), .A2(n4055), .ZN(n4988) );
  NAND2_X1 U4987 ( .A1(n4989), .A2(n4988), .ZN(n4987) );
  NAND2_X1 U4988 ( .A1(n4110), .A2(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n4057) );
  OAI211_X1 U4989 ( .C1(n4202), .C2(EBX_REG_13__SCAN_IN), .A(n4103), .B(n4057), 
        .ZN(n4058) );
  OAI21_X1 U4990 ( .B1(n4090), .B2(EBX_REG_13__SCAN_IN), .A(n4058), .ZN(n5040)
         );
  MUX2_X1 U4991 ( .A(n4091), .B(n4103), .S(EBX_REG_14__SCAN_IN), .Z(n4063) );
  NAND2_X1 U4992 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n4202), .ZN(n4061) );
  AND2_X1 U4993 ( .A1(n4085), .A2(n4061), .ZN(n4062) );
  AND2_X1 U4994 ( .A1(n4063), .A2(n4062), .ZN(n5070) );
  OR2_X2 U4995 ( .A1(n5071), .A2(n5070), .ZN(n5073) );
  NAND2_X1 U4996 ( .A1(n4110), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n4064) );
  OAI211_X1 U4997 ( .C1(n4202), .C2(EBX_REG_15__SCAN_IN), .A(n4103), .B(n4064), 
        .ZN(n4065) );
  OAI21_X1 U4998 ( .B1(n4090), .B2(EBX_REG_15__SCAN_IN), .A(n4065), .ZN(n5058)
         );
  MUX2_X1 U4999 ( .A(n4091), .B(n4103), .S(EBX_REG_16__SCAN_IN), .Z(n4068) );
  NAND2_X1 U5000 ( .A1(INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n4202), .ZN(n4066) );
  AND2_X1 U5001 ( .A1(n4085), .A2(n4066), .ZN(n4067) );
  NAND2_X1 U5002 ( .A1(n4068), .A2(n4067), .ZN(n5117) );
  NAND2_X1 U5003 ( .A1(n5118), .A2(n5117), .ZN(n5116) );
  NAND2_X1 U5004 ( .A1(n4110), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n4069) );
  OAI211_X1 U5005 ( .C1(n4202), .C2(EBX_REG_17__SCAN_IN), .A(n4103), .B(n4069), 
        .ZN(n4070) );
  OAI21_X1 U5006 ( .B1(n4090), .B2(EBX_REG_17__SCAN_IN), .A(n4070), .ZN(n5132)
         );
  NOR2_X2 U5007 ( .A1(n5116), .A2(n5132), .ZN(n5131) );
  INV_X1 U5008 ( .A(EBX_REG_19__SCAN_IN), .ZN(n5338) );
  NAND2_X1 U5009 ( .A1(n4334), .A2(n5338), .ZN(n4072) );
  AOI21_X1 U5010 ( .B1(n4103), .B2(n5613), .A(n4208), .ZN(n4071) );
  AOI22_X1 U5011 ( .A1(n4107), .A2(n5338), .B1(n4072), .B2(n4071), .ZN(n5336)
         );
  NAND2_X1 U5012 ( .A1(n4309), .A2(EBX_REG_18__SCAN_IN), .ZN(n4075) );
  NAND2_X1 U5013 ( .A1(n4202), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n4074) );
  AND2_X1 U5014 ( .A1(n4075), .A2(n4074), .ZN(n5409) );
  NAND2_X1 U5015 ( .A1(n5409), .A2(n4208), .ZN(n5335) );
  OR2_X1 U5016 ( .A1(n4202), .A2(EBX_REG_20__SCAN_IN), .ZN(n4076) );
  OAI21_X1 U5017 ( .B1(n4309), .B2(INSTADDRPOINTER_REG_20__SCAN_IN), .A(n4076), 
        .ZN(n5410) );
  NAND2_X1 U5018 ( .A1(n5335), .A2(n5410), .ZN(n4080) );
  INV_X1 U5019 ( .A(n5410), .ZN(n4078) );
  INV_X1 U5020 ( .A(n5409), .ZN(n4077) );
  NAND2_X1 U5021 ( .A1(n4077), .A2(n4110), .ZN(n5334) );
  NAND2_X1 U5022 ( .A1(n4078), .A2(n5334), .ZN(n4079) );
  AND2_X1 U5023 ( .A1(n4080), .A2(n4079), .ZN(n4081) );
  INV_X1 U5024 ( .A(EBX_REG_21__SCAN_IN), .ZN(n5404) );
  MUX2_X1 U5025 ( .A(n4208), .B(n4100), .S(n5404), .Z(n4083) );
  NOR2_X1 U5026 ( .A1(n4309), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n4082)
         );
  NOR2_X1 U5027 ( .A1(n4083), .A2(n4082), .ZN(n5402) );
  NAND2_X1 U5028 ( .A1(n5403), .A2(n5402), .ZN(n5394) );
  MUX2_X1 U5029 ( .A(n4091), .B(n4103), .S(EBX_REG_22__SCAN_IN), .Z(n4087) );
  NAND2_X1 U5030 ( .A1(n4202), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n4084) );
  AND2_X1 U5031 ( .A1(n4085), .A2(n4084), .ZN(n4086) );
  AND2_X1 U5032 ( .A1(n4087), .A2(n4086), .ZN(n5397) );
  OR2_X2 U5033 ( .A1(n5394), .A2(n5397), .ZN(n5395) );
  NAND2_X1 U5034 ( .A1(n4110), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4088) );
  OAI211_X1 U5035 ( .C1(n4202), .C2(EBX_REG_23__SCAN_IN), .A(n4103), .B(n4088), 
        .ZN(n4089) );
  OAI21_X1 U5036 ( .B1(n4090), .B2(EBX_REG_23__SCAN_IN), .A(n4089), .ZN(n5318)
         );
  MUX2_X1 U5037 ( .A(n4091), .B(n4103), .S(EBX_REG_24__SCAN_IN), .Z(n4093) );
  NAND2_X1 U5038 ( .A1(INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n4202), .ZN(n4092) );
  NAND2_X1 U5039 ( .A1(n4093), .A2(n4092), .ZN(n5260) );
  NAND2_X1 U5040 ( .A1(n5317), .A2(n5260), .ZN(n5259) );
  MUX2_X1 U5041 ( .A(n4100), .B(n4208), .S(EBX_REG_25__SCAN_IN), .Z(n4094) );
  INV_X1 U5042 ( .A(n4094), .ZN(n4096) );
  NAND2_X1 U5043 ( .A1(n4219), .A2(n5209), .ZN(n4095) );
  NAND2_X1 U5044 ( .A1(n4096), .A2(n4095), .ZN(n5383) );
  INV_X1 U5045 ( .A(n4097), .ZN(n5384) );
  INV_X1 U5046 ( .A(EBX_REG_26__SCAN_IN), .ZN(n5663) );
  NAND2_X1 U5047 ( .A1(n4334), .A2(n5663), .ZN(n4099) );
  AOI21_X1 U5048 ( .B1(n4103), .B2(n5208), .A(n4208), .ZN(n4098) );
  AOI22_X1 U5049 ( .A1(n4107), .A2(n5663), .B1(n4099), .B2(n4098), .ZN(n5374)
         );
  NOR2_X2 U5050 ( .A1(n5384), .A2(n5374), .ZN(n5376) );
  INV_X1 U5051 ( .A(EBX_REG_27__SCAN_IN), .ZN(n5370) );
  MUX2_X1 U5052 ( .A(n4208), .B(n4100), .S(n5370), .Z(n4102) );
  NOR2_X1 U5053 ( .A1(n4309), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n4101)
         );
  NOR2_X1 U5054 ( .A1(n4102), .A2(n4101), .ZN(n5202) );
  NAND2_X1 U5055 ( .A1(n5376), .A2(n5202), .ZN(n5364) );
  INV_X1 U5056 ( .A(EBX_REG_28__SCAN_IN), .ZN(n6607) );
  NAND2_X1 U5057 ( .A1(n4334), .A2(n6607), .ZN(n4105) );
  AOI21_X1 U5058 ( .B1(n4103), .B2(n6586), .A(n4208), .ZN(n4104) );
  AOI22_X1 U5059 ( .A1(n4107), .A2(n6607), .B1(n4105), .B2(n4104), .ZN(n5363)
         );
  OR2_X2 U5060 ( .A1(n5364), .A2(n5363), .ZN(n5366) );
  OR2_X1 U5061 ( .A1(n4202), .A2(EBX_REG_29__SCAN_IN), .ZN(n4106) );
  OAI21_X1 U5062 ( .B1(n4309), .B2(INSTADDRPOINTER_REG_29__SCAN_IN), .A(n4106), 
        .ZN(n4209) );
  OR2_X2 U5063 ( .A1(n5366), .A2(n4209), .ZN(n4172) );
  INV_X1 U5064 ( .A(EBX_REG_29__SCAN_IN), .ZN(n5359) );
  NAND2_X1 U5065 ( .A1(n4107), .A2(n5359), .ZN(n4207) );
  OAI21_X2 U5066 ( .B1(n4172), .B2(n4208), .A(n2978), .ZN(n4213) );
  NAND2_X1 U5067 ( .A1(n4309), .A2(EBX_REG_30__SCAN_IN), .ZN(n4109) );
  NAND2_X1 U5068 ( .A1(n4202), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4108) );
  AND2_X1 U5069 ( .A1(n4109), .A2(n4108), .ZN(n4171) );
  NAND2_X1 U5070 ( .A1(n4213), .A2(n4171), .ZN(n4111) );
  NAND2_X1 U5071 ( .A1(n4172), .A2(n4110), .ZN(n4174) );
  INV_X1 U5072 ( .A(EBX_REG_31__SCAN_IN), .ZN(n5357) );
  AOI22_X1 U5073 ( .A1(n4219), .A2(n6623), .B1(n4334), .B2(n5357), .ZN(n4112)
         );
  INV_X1 U5074 ( .A(READY_N), .ZN(n6492) );
  NAND2_X1 U5075 ( .A1(n6492), .A2(n6234), .ZN(n4157) );
  OR4_X1 U5076 ( .A1(n4120), .A2(n4119), .A3(n4118), .A4(n4117), .ZN(n4121) );
  NAND2_X1 U5077 ( .A1(n4122), .A2(n4121), .ZN(n5291) );
  NOR2_X1 U5078 ( .A1(n4218), .A2(n5291), .ZN(n5298) );
  NAND2_X1 U5079 ( .A1(n5298), .A2(n6383), .ZN(n4266) );
  NOR2_X1 U5080 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n6497) );
  INV_X1 U5081 ( .A(n6497), .ZN(n6392) );
  NOR3_X1 U5082 ( .A1(n6382), .A2(n6470), .A3(n6392), .ZN(n6377) );
  NOR3_X1 U5083 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n6391), .A3(n4123), .ZN(
        n6387) );
  INV_X1 U5084 ( .A(n6387), .ZN(n4124) );
  NAND2_X1 U5085 ( .A1(n6047), .A2(n4124), .ZN(n4125) );
  OR2_X1 U5086 ( .A1(n6377), .A2(n4125), .ZN(n4126) );
  OR2_X2 U5087 ( .A1(n6490), .A2(n4126), .ZN(n5016) );
  INV_X1 U5088 ( .A(n4955), .ZN(n4161) );
  AND2_X1 U5089 ( .A1(EBX_REG_31__SCAN_IN), .A2(n4161), .ZN(n4142) );
  AND2_X1 U5090 ( .A1(n4157), .A2(n4142), .ZN(n4127) );
  INV_X1 U5091 ( .A(REIP_REG_26__SCAN_IN), .ZN(n6451) );
  INV_X1 U5092 ( .A(REIP_REG_20__SCAN_IN), .ZN(n6632) );
  INV_X1 U5093 ( .A(REIP_REG_18__SCAN_IN), .ZN(n6543) );
  INV_X1 U5094 ( .A(REIP_REG_15__SCAN_IN), .ZN(n6436) );
  INV_X1 U5095 ( .A(n4128), .ZN(n4129) );
  NOR2_X1 U5096 ( .A1(n4220), .A2(n4129), .ZN(n4132) );
  INV_X1 U5097 ( .A(STATE_REG_0__SCAN_IN), .ZN(n4130) );
  NAND2_X1 U5098 ( .A1(n4131), .A2(n4130), .ZN(n6402) );
  NAND2_X1 U5099 ( .A1(n4217), .A2(n6402), .ZN(n4185) );
  NAND2_X1 U5100 ( .A1(n4132), .A2(n4185), .ZN(n5003) );
  NAND3_X1 U5101 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_3__SCAN_IN), .A3(
        REIP_REG_2__SCAN_IN), .ZN(n4133) );
  NOR2_X2 U5102 ( .A1(n5003), .A2(n4133), .ZN(n4972) );
  INV_X1 U5103 ( .A(REIP_REG_8__SCAN_IN), .ZN(n6424) );
  NAND4_X1 U5104 ( .A1(REIP_REG_7__SCAN_IN), .A2(REIP_REG_6__SCAN_IN), .A3(
        REIP_REG_5__SCAN_IN), .A4(REIP_REG_4__SCAN_IN), .ZN(n4994) );
  NOR2_X1 U5105 ( .A1(n6424), .A2(n4994), .ZN(n4136) );
  NAND2_X1 U5106 ( .A1(n4972), .A2(n4136), .ZN(n5818) );
  NAND3_X1 U5107 ( .A1(REIP_REG_11__SCAN_IN), .A2(REIP_REG_10__SCAN_IN), .A3(
        REIP_REG_9__SCAN_IN), .ZN(n4134) );
  NAND4_X1 U5108 ( .A1(n5807), .A2(REIP_REG_14__SCAN_IN), .A3(
        REIP_REG_13__SCAN_IN), .A4(REIP_REG_12__SCAN_IN), .ZN(n5062) );
  NAND3_X1 U5109 ( .A1(n5342), .A2(REIP_REG_17__SCAN_IN), .A3(
        REIP_REG_16__SCAN_IN), .ZN(n5331) );
  NAND2_X1 U5110 ( .A1(REIP_REG_19__SCAN_IN), .A2(n5328), .ZN(n5712) );
  NOR2_X2 U5111 ( .A1(n6632), .A2(n5712), .ZN(n5704) );
  NAND2_X1 U5112 ( .A1(REIP_REG_22__SCAN_IN), .A2(REIP_REG_21__SCAN_IN), .ZN(
        n5695) );
  INV_X1 U5113 ( .A(REIP_REG_23__SCAN_IN), .ZN(n6446) );
  NOR2_X2 U5114 ( .A1(n5315), .A2(n6446), .ZN(n5689) );
  NAND3_X1 U5115 ( .A1(REIP_REG_24__SCAN_IN), .A2(REIP_REG_25__SCAN_IN), .A3(
        n5689), .ZN(n5665) );
  NOR2_X2 U5116 ( .A1(n6451), .A2(n5665), .ZN(n5657) );
  NAND3_X1 U5117 ( .A1(n5657), .A2(REIP_REG_28__SCAN_IN), .A3(
        REIP_REG_27__SCAN_IN), .ZN(n5649) );
  INV_X1 U5118 ( .A(REIP_REG_29__SCAN_IN), .ZN(n6458) );
  NAND3_X1 U5119 ( .A1(REIP_REG_30__SCAN_IN), .A2(n4164), .A3(n6462), .ZN(
        n4146) );
  NAND2_X1 U5120 ( .A1(n5016), .A2(n5003), .ZN(n5330) );
  NAND2_X1 U5121 ( .A1(REIP_REG_28__SCAN_IN), .A2(REIP_REG_27__SCAN_IN), .ZN(
        n4139) );
  NAND2_X1 U5122 ( .A1(REIP_REG_24__SCAN_IN), .A2(REIP_REG_25__SCAN_IN), .ZN(
        n5677) );
  INV_X1 U5123 ( .A(REIP_REG_19__SCAN_IN), .ZN(n6441) );
  NAND3_X1 U5124 ( .A1(REIP_REG_14__SCAN_IN), .A2(REIP_REG_13__SCAN_IN), .A3(
        REIP_REG_12__SCAN_IN), .ZN(n4137) );
  INV_X1 U5125 ( .A(REIP_REG_1__SCAN_IN), .ZN(n6580) );
  INV_X1 U5126 ( .A(REIP_REG_3__SCAN_IN), .ZN(n6590) );
  INV_X1 U5127 ( .A(REIP_REG_2__SCAN_IN), .ZN(n6416) );
  INV_X1 U5128 ( .A(n5016), .ZN(n5002) );
  NOR4_X1 U5129 ( .A1(n6580), .A2(n6590), .A3(n6416), .A4(n5002), .ZN(n5852)
         );
  AND2_X1 U5130 ( .A1(n4136), .A2(n5852), .ZN(n4922) );
  NAND4_X1 U5131 ( .A1(REIP_REG_11__SCAN_IN), .A2(REIP_REG_10__SCAN_IN), .A3(
        REIP_REG_9__SCAN_IN), .A4(n4922), .ZN(n5043) );
  NOR2_X1 U5132 ( .A1(n4137), .A2(n5043), .ZN(n5066) );
  NAND4_X1 U5133 ( .A1(REIP_REG_15__SCAN_IN), .A2(REIP_REG_17__SCAN_IN), .A3(
        REIP_REG_16__SCAN_IN), .A4(n5066), .ZN(n5329) );
  NOR4_X1 U5134 ( .A1(n6632), .A2(n6441), .A3(n6543), .A4(n5329), .ZN(n5692)
         );
  NAND4_X1 U5135 ( .A1(REIP_REG_23__SCAN_IN), .A2(REIP_REG_22__SCAN_IN), .A3(
        REIP_REG_21__SCAN_IN), .A4(n5692), .ZN(n5316) );
  NOR2_X1 U5136 ( .A1(n5677), .A2(n5316), .ZN(n4138) );
  AOI21_X1 U5137 ( .B1(n4138), .B2(REIP_REG_26__SCAN_IN), .A(n5853), .ZN(n5667) );
  AOI21_X1 U5138 ( .B1(n4139), .B2(n5330), .A(n5667), .ZN(n5654) );
  OAI211_X1 U5139 ( .C1(REIP_REG_29__SCAN_IN), .C2(n5853), .A(n5654), .B(
        REIP_REG_30__SCAN_IN), .ZN(n4163) );
  NAND3_X1 U5140 ( .A1(REIP_REG_31__SCAN_IN), .A2(n5330), .A3(n4163), .ZN(
        n4144) );
  INV_X1 U5141 ( .A(n6402), .ZN(n4488) );
  INV_X1 U5142 ( .A(n4157), .ZN(n4140) );
  NAND2_X1 U5143 ( .A1(n4488), .A2(n4140), .ZN(n6371) );
  NAND2_X1 U5144 ( .A1(n4394), .A2(n6371), .ZN(n4160) );
  INV_X1 U5145 ( .A(n4160), .ZN(n4141) );
  AOI22_X1 U5146 ( .A1(n5870), .A2(PHYADDRPOINTER_REG_31__SCAN_IN), .B1(n4142), 
        .B2(n4141), .ZN(n4143) );
  AOI21_X1 U5147 ( .B1(n5356), .B2(n5866), .A(n4147), .ZN(n4150) );
  AND2_X1 U5148 ( .A1(n4154), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4148) );
  INV_X1 U5149 ( .A(n4151), .ZN(n4152) );
  AOI21_X1 U5150 ( .B1(n4153), .B2(n5174), .A(n4152), .ZN(n5191) );
  INV_X1 U5151 ( .A(n5191), .ZN(n5276) );
  NOR2_X1 U5152 ( .A1(n4154), .A2(n6391), .ZN(n4155) );
  INV_X1 U5153 ( .A(n4156), .ZN(n5189) );
  INV_X1 U5154 ( .A(EBX_REG_30__SCAN_IN), .ZN(n5146) );
  NAND2_X1 U5155 ( .A1(n4157), .A2(n5357), .ZN(n4158) );
  OR2_X1 U5156 ( .A1(n4220), .A2(n4158), .ZN(n4159) );
  NAND2_X1 U5157 ( .A1(n4160), .A2(n4159), .ZN(n4162) );
  AND2_X2 U5158 ( .A1(n4162), .A2(n4161), .ZN(n5865) );
  INV_X1 U5159 ( .A(n5865), .ZN(n5662) );
  OAI22_X1 U5160 ( .A1(n5868), .A2(n5189), .B1(n5146), .B2(n5662), .ZN(n4168)
         );
  AND2_X1 U5161 ( .A1(n5870), .A2(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n4167)
         );
  OAI21_X1 U5162 ( .B1(n4164), .B2(REIP_REG_30__SCAN_IN), .A(n4163), .ZN(n4165) );
  INV_X1 U5163 ( .A(n5366), .ZN(n4170) );
  INV_X1 U5164 ( .A(n4171), .ZN(n4169) );
  AOI21_X1 U5165 ( .B1(n4172), .B2(n4170), .A(n4169), .ZN(n4175) );
  AOI21_X1 U5166 ( .B1(n5366), .B2(n4208), .A(n4171), .ZN(n4173) );
  NAND3_X1 U5167 ( .A1(n4177), .A2(n4176), .A3(n2979), .ZN(U2797) );
  NOR2_X1 U5168 ( .A1(n4179), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n4180)
         );
  AOI22_X1 U5169 ( .A1(n5457), .A2(n5543), .B1(n4180), .B2(n5466), .ZN(n4181)
         );
  NAND2_X1 U5170 ( .A1(n4391), .A2(n6402), .ZN(n4182) );
  NOR2_X1 U5171 ( .A1(READY_N), .A2(n5291), .ZN(n4274) );
  NAND2_X1 U5172 ( .A1(n4182), .A2(n4274), .ZN(n4190) );
  NAND2_X1 U5173 ( .A1(n4185), .A2(n6492), .ZN(n4186) );
  OAI211_X1 U5174 ( .C1(n4184), .C2(n4186), .A(n4377), .B(n5270), .ZN(n4187)
         );
  INV_X1 U5175 ( .A(n4187), .ZN(n4188) );
  OR2_X1 U5176 ( .A1(n5302), .A2(n4188), .ZN(n4189) );
  MUX2_X1 U5177 ( .A(n4190), .B(n4189), .S(n3135), .Z(n4197) );
  OR2_X1 U5178 ( .A1(n4191), .A2(n3111), .ZN(n4194) );
  NAND2_X1 U5179 ( .A1(n4192), .A2(n3494), .ZN(n4235) );
  AND2_X1 U5180 ( .A1(n4235), .A2(n4377), .ZN(n4193) );
  NAND2_X1 U5181 ( .A1(n4194), .A2(n4193), .ZN(n4225) );
  NAND2_X1 U5182 ( .A1(n4200), .A2(n4225), .ZN(n4195) );
  NAND2_X1 U5183 ( .A1(n4195), .A2(n4218), .ZN(n4234) );
  NAND3_X1 U5184 ( .A1(n5302), .A2(n5277), .A3(n4391), .ZN(n4196) );
  NAND3_X1 U5185 ( .A1(n4197), .A2(n4234), .A3(n4196), .ZN(n4198) );
  INV_X1 U5186 ( .A(n5301), .ZN(n4199) );
  NAND2_X1 U5187 ( .A1(n4200), .A2(n4199), .ZN(n4512) );
  AND2_X1 U5188 ( .A1(n4512), .A2(n4201), .ZN(n5293) );
  OR2_X1 U5189 ( .A1(n4184), .A2(n4202), .ZN(n4490) );
  INV_X1 U5190 ( .A(n4203), .ZN(n4204) );
  NAND2_X1 U5191 ( .A1(n4204), .A2(n4370), .ZN(n4205) );
  NAND4_X1 U5192 ( .A1(n5293), .A2(n4505), .A3(n4490), .A4(n4205), .ZN(n4206)
         );
  NAND2_X1 U5193 ( .A1(n5172), .A2(n6050), .ZN(n4265) );
  OAI21_X1 U5194 ( .B1(n4209), .B2(n4208), .A(n4207), .ZN(n4210) );
  INV_X1 U5195 ( .A(n4210), .ZN(n4211) );
  AND2_X1 U5196 ( .A1(n5366), .A2(n4211), .ZN(n4212) );
  OR2_X1 U5197 ( .A1(n4213), .A2(n4212), .ZN(n5644) );
  INV_X1 U5198 ( .A(n4394), .ZN(n6496) );
  OR2_X1 U5199 ( .A1(n4184), .A2(n6496), .ZN(n6370) );
  NAND3_X1 U5200 ( .A1(n4214), .A2(n3155), .A3(n4221), .ZN(n4215) );
  NAND2_X1 U5201 ( .A1(n6370), .A2(n4215), .ZN(n4216) );
  NOR2_X1 U5202 ( .A1(n4218), .A2(n4217), .ZN(n6347) );
  NAND2_X1 U5203 ( .A1(n4245), .A2(n6347), .ZN(n5085) );
  NAND2_X1 U5204 ( .A1(n4220), .A2(n4391), .ZN(n4956) );
  OR2_X1 U5205 ( .A1(n4956), .A2(n4363), .ZN(n4233) );
  NAND2_X1 U5206 ( .A1(n4219), .A2(n4233), .ZN(n4224) );
  AOI21_X1 U5207 ( .B1(n4221), .B2(n4220), .A(n3135), .ZN(n4222) );
  AOI21_X1 U5208 ( .B1(n4224), .B2(n4223), .A(n4222), .ZN(n4226) );
  OAI211_X1 U5209 ( .C1(n4227), .C2(n4110), .A(n4226), .B(n4225), .ZN(n4228)
         );
  INV_X1 U5210 ( .A(n4228), .ZN(n4229) );
  NAND2_X1 U5211 ( .A1(n4230), .A2(n4229), .ZN(n4508) );
  OAI21_X1 U5212 ( .B1(n4506), .B2(n4377), .A(n4527), .ZN(n4231) );
  OR2_X1 U5213 ( .A1(n4508), .A2(n4231), .ZN(n4232) );
  NAND2_X1 U5214 ( .A1(n4245), .A2(n4232), .ZN(n4313) );
  NAND2_X1 U5215 ( .A1(n5085), .A2(n4313), .ZN(n5600) );
  AND2_X1 U5216 ( .A1(n4234), .A2(n4233), .ZN(n4493) );
  INV_X1 U5217 ( .A(n4235), .ZN(n4236) );
  NAND2_X1 U5218 ( .A1(n4245), .A2(n5289), .ZN(n5598) );
  INV_X1 U5219 ( .A(n5598), .ZN(n6040) );
  OR2_X1 U5220 ( .A1(n5600), .A2(n6040), .ZN(n5194) );
  INV_X1 U5221 ( .A(n5194), .ZN(n5601) );
  NAND2_X1 U5222 ( .A1(INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5556) );
  NOR2_X1 U5223 ( .A1(n6570), .A2(n6006), .ZN(n6001) );
  INV_X1 U5224 ( .A(n6001), .ZN(n4945) );
  NAND2_X1 U5225 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n4946) );
  NOR2_X1 U5226 ( .A1(n4945), .A2(n4946), .ZN(n4242) );
  AOI21_X1 U5227 ( .B1(INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .A(INSTADDRPOINTER_REG_2__SCAN_IN), 
        .ZN(n6041) );
  NAND2_X1 U5228 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n6028) );
  NOR2_X1 U5229 ( .A1(n6041), .A2(n6028), .ZN(n6015) );
  NAND2_X1 U5230 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n6015), .ZN(n4575)
         );
  NOR2_X1 U5231 ( .A1(n4240), .A2(n4575), .ZN(n4947) );
  NAND2_X1 U5232 ( .A1(n4242), .A2(n4947), .ZN(n5087) );
  INV_X1 U5233 ( .A(n5087), .ZN(n4238) );
  NAND2_X1 U5234 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n4252) );
  NAND2_X1 U5235 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n5974) );
  INV_X1 U5236 ( .A(n5974), .ZN(n5092) );
  NAND2_X1 U5237 ( .A1(INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n5092), .ZN(n5099) );
  NOR2_X1 U5238 ( .A1(n5083), .A2(n5099), .ZN(n5159) );
  INV_X1 U5239 ( .A(n5159), .ZN(n4237) );
  NOR2_X1 U5240 ( .A1(n4252), .A2(n4237), .ZN(n4244) );
  NAND2_X1 U5241 ( .A1(n4238), .A2(n4244), .ZN(n5596) );
  INV_X1 U5242 ( .A(n4239), .ZN(n4257) );
  OR3_X1 U5243 ( .A1(n5596), .A2(n4256), .A3(n4257), .ZN(n4249) );
  NAND2_X1 U5244 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4573) );
  NOR4_X1 U5245 ( .A1(n4241), .A2(n4240), .A3(n4573), .A4(n6028), .ZN(n4948)
         );
  NAND2_X1 U5246 ( .A1(n4948), .A2(n4242), .ZN(n5090) );
  INV_X1 U5247 ( .A(n5090), .ZN(n4243) );
  INV_X1 U5248 ( .A(n5600), .ZN(n4949) );
  AOI21_X1 U5249 ( .B1(n4244), .B2(n4243), .A(n4949), .ZN(n4247) );
  OR2_X1 U5250 ( .A1(n4313), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4246)
         );
  OR2_X1 U5251 ( .A1(n4245), .A2(n6032), .ZN(n4321) );
  NAND2_X1 U5252 ( .A1(n4246), .A2(n4321), .ZN(n5086) );
  NOR2_X1 U5253 ( .A1(n4247), .A2(n5086), .ZN(n5597) );
  INV_X1 U5254 ( .A(n5597), .ZN(n4248) );
  AOI21_X1 U5255 ( .B1(n5194), .B2(n4249), .A(n4248), .ZN(n5577) );
  OAI21_X1 U5256 ( .B1(n5579), .B2(n5601), .A(n5577), .ZN(n5569) );
  INV_X1 U5257 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4250) );
  NAND2_X1 U5258 ( .A1(n4250), .A2(n5085), .ZN(n4319) );
  NAND2_X1 U5259 ( .A1(n5600), .A2(n4319), .ZN(n4571) );
  AOI21_X1 U5260 ( .B1(n4571), .B2(n5598), .A(n4258), .ZN(n4251) );
  NOR2_X1 U5261 ( .A1(n5569), .A2(n4251), .ZN(n5262) );
  INV_X1 U5262 ( .A(n5262), .ZN(n5566) );
  AOI21_X1 U5263 ( .B1(n5194), .B2(n5556), .A(n5566), .ZN(n5549) );
  OAI21_X1 U5264 ( .B1(n5543), .B2(n5601), .A(n5549), .ZN(n5193) );
  NOR2_X1 U5265 ( .A1(n6047), .A2(n6458), .ZN(n5176) );
  INV_X1 U5266 ( .A(n4252), .ZN(n4255) );
  NOR2_X1 U5267 ( .A1(n4571), .A2(n5090), .ZN(n5975) );
  INV_X1 U5268 ( .A(n5975), .ZN(n4254) );
  NOR2_X1 U5269 ( .A1(n5598), .A2(n5087), .ZN(n5095) );
  INV_X1 U5270 ( .A(n5095), .ZN(n4253) );
  NAND2_X1 U5271 ( .A1(n4254), .A2(n4253), .ZN(n5984) );
  NAND2_X1 U5272 ( .A1(n4255), .A2(n5742), .ZN(n5741) );
  NOR2_X1 U5273 ( .A1(n5602), .A2(n4257), .ZN(n5578) );
  NAND2_X1 U5274 ( .A1(n5578), .A2(n5579), .ZN(n5572) );
  INV_X1 U5275 ( .A(n4258), .ZN(n4259) );
  NOR2_X1 U5276 ( .A1(n5564), .A2(n5556), .ZN(n5546) );
  AND2_X1 U5277 ( .A1(n5546), .A2(n5543), .ZN(n5218) );
  INV_X1 U5278 ( .A(n5218), .ZN(n4260) );
  NOR2_X1 U5279 ( .A1(n4260), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4261)
         );
  AOI211_X1 U5280 ( .C1(n5193), .C2(INSTADDRPOINTER_REG_29__SCAN_IN), .A(n5176), .B(n4261), .ZN(n4262) );
  NAND2_X1 U5281 ( .A1(n4265), .A2(n4264), .ZN(U2989) );
  INV_X1 U5282 ( .A(n4392), .ZN(n4393) );
  AOI211_X1 U5283 ( .C1(MEMORYFETCH_REG_SCAN_IN), .C2(n4266), .A(n4923), .B(
        n4393), .ZN(n4267) );
  INV_X1 U5284 ( .A(n4267), .ZN(U2788) );
  INV_X1 U5285 ( .A(n6490), .ZN(n4270) );
  INV_X1 U5286 ( .A(n4956), .ZN(n4268) );
  OR2_X1 U5287 ( .A1(n4394), .A2(n4268), .ZN(n5303) );
  OAI21_X1 U5288 ( .B1(n4923), .B2(READREQUEST_REG_SCAN_IN), .A(n4270), .ZN(
        n4269) );
  OAI21_X1 U5289 ( .B1(n4270), .B2(n5303), .A(n4269), .ZN(U3474) );
  OAI21_X1 U5290 ( .B1(n4273), .B2(n4272), .A(n4271), .ZN(n4962) );
  INV_X1 U5291 ( .A(n4274), .ZN(n4275) );
  OAI22_X1 U5292 ( .A1(n5302), .A2(n4512), .B1(n4505), .B2(n4275), .ZN(n4497)
         );
  NAND2_X1 U5293 ( .A1(n4497), .A2(n6383), .ZN(n4281) );
  INV_X1 U5294 ( .A(n5271), .ZN(n5429) );
  NAND4_X1 U5295 ( .A1(n5429), .A2(n3155), .A3(n6383), .A4(n4276), .ZN(n4332)
         );
  NAND2_X1 U5296 ( .A1(n6383), .A2(n6492), .ZN(n4278) );
  OAI21_X1 U5297 ( .B1(n4332), .B2(n4504), .A(n5928), .ZN(n4279) );
  INV_X1 U5298 ( .A(n4279), .ZN(n4280) );
  NAND2_X1 U5299 ( .A1(n4282), .A2(n5271), .ZN(n4283) );
  NAND2_X2 U5300 ( .A1(n5435), .A2(n4283), .ZN(n5718) );
  INV_X1 U5301 ( .A(n4283), .ZN(n4284) );
  INV_X2 U5302 ( .A(n5435), .ZN(n5884) );
  AOI22_X1 U5303 ( .A1(n5060), .A2(DATAI_0_), .B1(n5884), .B2(
        EAX_REG_0__SCAN_IN), .ZN(n4285) );
  OAI21_X1 U5304 ( .B1(n4962), .B2(n5718), .A(n4285), .ZN(U2891) );
  INV_X1 U5305 ( .A(EAX_REG_27__SCAN_IN), .ZN(n4456) );
  INV_X1 U5306 ( .A(n6347), .ZN(n5280) );
  AND2_X1 U5307 ( .A1(n6370), .A2(n5280), .ZN(n4287) );
  NAND2_X1 U5308 ( .A1(n4488), .A2(n6383), .ZN(n4286) );
  NAND2_X1 U5309 ( .A1(n4288), .A2(n4377), .ZN(n4474) );
  NOR2_X1 U5310 ( .A1(n6391), .A2(n6379), .ZN(n6388) );
  NAND2_X1 U5311 ( .A1(n6382), .A2(n6388), .ZN(n6368) );
  AOI22_X1 U5313 ( .A1(n6493), .A2(UWORD_REG_11__SCAN_IN), .B1(n5888), .B2(
        DATAO_REG_27__SCAN_IN), .ZN(n4289) );
  OAI21_X1 U5314 ( .B1(n4456), .B2(n4474), .A(n4289), .ZN(U2896) );
  AOI22_X1 U5315 ( .A1(n6493), .A2(UWORD_REG_8__SCAN_IN), .B1(n5888), .B2(
        DATAO_REG_24__SCAN_IN), .ZN(n4290) );
  OAI21_X1 U5316 ( .B1(n3902), .B2(n4474), .A(n4290), .ZN(U2899) );
  AOI22_X1 U5317 ( .A1(n6493), .A2(UWORD_REG_10__SCAN_IN), .B1(n5888), .B2(
        DATAO_REG_26__SCAN_IN), .ZN(n4291) );
  OAI21_X1 U5318 ( .B1(n3910), .B2(n4474), .A(n4291), .ZN(U2897) );
  INV_X1 U5319 ( .A(EAX_REG_22__SCAN_IN), .ZN(n4467) );
  AOI22_X1 U5321 ( .A1(n6493), .A2(UWORD_REG_6__SCAN_IN), .B1(n5888), .B2(
        DATAO_REG_22__SCAN_IN), .ZN(n4292) );
  OAI21_X1 U5322 ( .B1(n4467), .B2(n4474), .A(n4292), .ZN(U2901) );
  INV_X1 U5323 ( .A(EAX_REG_19__SCAN_IN), .ZN(n4410) );
  AOI22_X1 U5324 ( .A1(n6493), .A2(UWORD_REG_3__SCAN_IN), .B1(n5888), .B2(
        DATAO_REG_19__SCAN_IN), .ZN(n4293) );
  OAI21_X1 U5325 ( .B1(n4410), .B2(n4474), .A(n4293), .ZN(U2904) );
  INV_X1 U5326 ( .A(EAX_REG_20__SCAN_IN), .ZN(n4404) );
  AOI22_X1 U5327 ( .A1(n6493), .A2(UWORD_REG_4__SCAN_IN), .B1(n5888), .B2(
        DATAO_REG_20__SCAN_IN), .ZN(n4294) );
  OAI21_X1 U5328 ( .B1(n4404), .B2(n4474), .A(n4294), .ZN(U2903) );
  INV_X1 U5329 ( .A(EAX_REG_21__SCAN_IN), .ZN(n4471) );
  AOI22_X1 U5330 ( .A1(n6493), .A2(UWORD_REG_5__SCAN_IN), .B1(n5888), .B2(
        DATAO_REG_21__SCAN_IN), .ZN(n4295) );
  OAI21_X1 U5331 ( .B1(n4471), .B2(n4474), .A(n4295), .ZN(U2902) );
  INV_X1 U5332 ( .A(EAX_REG_17__SCAN_IN), .ZN(n4407) );
  AOI22_X1 U5333 ( .A1(n6493), .A2(UWORD_REG_1__SCAN_IN), .B1(n5888), .B2(
        DATAO_REG_17__SCAN_IN), .ZN(n4296) );
  OAI21_X1 U5334 ( .B1(n4407), .B2(n4474), .A(n4296), .ZN(U2906) );
  INV_X1 U5335 ( .A(EAX_REG_23__SCAN_IN), .ZN(n4461) );
  AOI22_X1 U5336 ( .A1(n6493), .A2(UWORD_REG_7__SCAN_IN), .B1(n5888), .B2(
        DATAO_REG_23__SCAN_IN), .ZN(n4297) );
  OAI21_X1 U5337 ( .B1(n4461), .B2(n4474), .A(n4297), .ZN(U2900) );
  OAI21_X1 U5338 ( .B1(n4300), .B2(n4299), .A(n4298), .ZN(n5020) );
  INV_X1 U5339 ( .A(n5060), .ZN(n4616) );
  INV_X1 U5340 ( .A(DATAI_1_), .ZN(n4301) );
  INV_X1 U5341 ( .A(EAX_REG_1__SCAN_IN), .ZN(n6540) );
  OAI222_X1 U5342 ( .A1(n5020), .A2(n5718), .B1(n4616), .B2(n4301), .C1(n5435), 
        .C2(n6540), .ZN(U2890) );
  XNOR2_X1 U5343 ( .A(n4302), .B(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4315)
         );
  INV_X1 U5344 ( .A(n4962), .ZN(n4306) );
  AND2_X1 U5345 ( .A1(n6032), .A2(REIP_REG_0__SCAN_IN), .ZN(n4311) );
  INV_X1 U5346 ( .A(n5963), .ZN(n5535) );
  INV_X1 U5347 ( .A(PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n4303) );
  AOI21_X1 U5348 ( .B1(n5535), .B2(n4304), .A(n4303), .ZN(n4305) );
  AOI211_X1 U5349 ( .C1(n4306), .C2(n5515), .A(n4311), .B(n4305), .ZN(n4307)
         );
  OAI21_X1 U5350 ( .B1(n4315), .B2(n5770), .A(n4307), .ZN(U2986) );
  OAI21_X1 U5351 ( .B1(n4309), .B2(INSTADDRPOINTER_REG_0__SCAN_IN), .A(n4308), 
        .ZN(n4957) );
  INV_X1 U5352 ( .A(n4957), .ZN(n4312) );
  AOI21_X1 U5353 ( .B1(n4321), .B2(n5085), .A(n4250), .ZN(n4310) );
  AOI211_X1 U5354 ( .C1(n6044), .C2(n4312), .A(n4311), .B(n4310), .ZN(n4314)
         );
  INV_X1 U5355 ( .A(n4313), .ZN(n5096) );
  NOR2_X1 U5356 ( .A1(n6040), .A2(n5096), .ZN(n5091) );
  OR2_X1 U5357 ( .A1(n5091), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4322)
         );
  OAI211_X1 U5358 ( .C1(n4315), .C2(n6023), .A(n4314), .B(n4322), .ZN(U3018)
         );
  XNOR2_X1 U5359 ( .A(n4317), .B(n4316), .ZN(n4791) );
  OAI21_X1 U5360 ( .B1(n5013), .B2(n4334), .A(n4318), .ZN(n4339) );
  NAND3_X1 U5361 ( .A1(n5149), .A2(n4319), .A3(n5194), .ZN(n4320) );
  OAI21_X1 U5362 ( .B1(n6047), .B2(n6580), .A(n4320), .ZN(n4324) );
  AOI21_X1 U5363 ( .B1(n4322), .B2(n4321), .A(n5149), .ZN(n4323) );
  AOI211_X1 U5364 ( .C1(n6044), .C2(n4339), .A(n4324), .B(n4323), .ZN(n4325)
         );
  OAI21_X1 U5365 ( .B1(n4791), .B2(n6023), .A(n4325), .ZN(U3017) );
  CLKBUF_X1 U5366 ( .A(n4326), .Z(n4477) );
  NOR2_X1 U5367 ( .A1(n4328), .A2(n4327), .ZN(n4329) );
  NOR2_X1 U5368 ( .A1(n4477), .A2(n4329), .ZN(n5969) );
  INV_X1 U5369 ( .A(n5969), .ZN(n5011) );
  AOI22_X1 U5370 ( .A1(n5060), .A2(DATAI_2_), .B1(n5884), .B2(
        EAX_REG_2__SCAN_IN), .ZN(n4330) );
  OAI21_X1 U5371 ( .B1(n5011), .B2(n5718), .A(n4330), .ZN(U2889) );
  AND2_X1 U5372 ( .A1(n5289), .A2(n6383), .ZN(n4331) );
  NAND2_X1 U5373 ( .A1(n5302), .A2(n4331), .ZN(n4338) );
  INV_X1 U5374 ( .A(n4332), .ZN(n4336) );
  INV_X1 U5375 ( .A(n4333), .ZN(n4335) );
  NAND3_X1 U5376 ( .A1(n4336), .A2(n4335), .A3(n4334), .ZN(n4337) );
  NAND2_X1 U5377 ( .A1(n5427), .A2(n5429), .ZN(n5428) );
  INV_X1 U5378 ( .A(n5427), .ZN(n5414) );
  AOI22_X1 U5379 ( .A1(n5415), .A2(n4339), .B1(n5414), .B2(EBX_REG_1__SCAN_IN), 
        .ZN(n4340) );
  OAI21_X1 U5380 ( .B1(n5020), .B2(n5417), .A(n4340), .ZN(U2858) );
  INV_X1 U5381 ( .A(n4480), .ZN(n4341) );
  XNOR2_X1 U5382 ( .A(n4481), .B(n4341), .ZN(n6043) );
  AOI22_X1 U5383 ( .A1(n5415), .A2(n6043), .B1(n5414), .B2(EBX_REG_2__SCAN_IN), 
        .ZN(n4342) );
  OAI21_X1 U5384 ( .B1(n5011), .B2(n5417), .A(n4342), .ZN(U2857) );
  OAI222_X1 U5385 ( .A1(n4962), .A2(n5417), .B1(n5427), .B2(n6652), .C1(n5428), 
        .C2(n4957), .ZN(U2859) );
  OR2_X1 U5386 ( .A1(n4694), .A2(n3297), .ZN(n4352) );
  OR2_X1 U5387 ( .A1(n5627), .A2(n6234), .ZN(n4582) );
  INV_X1 U5388 ( .A(n4582), .ZN(n4541) );
  AOI21_X1 U5389 ( .B1(n6119), .B2(n4541), .A(n6286), .ZN(n4350) );
  INV_X1 U5390 ( .A(n4350), .ZN(n4347) );
  INV_X1 U5391 ( .A(n4344), .ZN(n5628) );
  AND2_X1 U5392 ( .A1(n5628), .A2(n5632), .ZN(n6278) );
  INV_X1 U5393 ( .A(n4346), .ZN(n4485) );
  AND2_X1 U5394 ( .A1(n6278), .A2(n4485), .ZN(n6091) );
  NOR2_X1 U5395 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n4864), .ZN(n6282)
         );
  NAND2_X1 U5396 ( .A1(n6282), .A2(n6358), .ZN(n6090) );
  NOR2_X1 U5397 ( .A1(n6635), .A2(n6090), .ZN(n4355) );
  AOI21_X1 U5398 ( .B1(n6091), .B2(n3503), .A(n4355), .ZN(n4349) );
  OAI22_X1 U5399 ( .A1(n4347), .A2(n4349), .B1(n6090), .B2(n6379), .ZN(n4348)
         );
  INV_X1 U5400 ( .A(n4348), .ZN(n4388) );
  OAI21_X1 U5401 ( .B1(n6497), .B2(n6388), .A(n5637), .ZN(n4353) );
  NAND2_X1 U5402 ( .A1(n6382), .A2(n4353), .ZN(n6165) );
  NAND2_X1 U5403 ( .A1(DATAI_5_), .A2(n4701), .ZN(n6324) );
  AOI21_X1 U5404 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n6635), .A(n6165), .ZN(
        n6290) );
  AOI22_X1 U5405 ( .A1(n4350), .A2(n4349), .B1(n6090), .B2(n6286), .ZN(n4351)
         );
  NAND2_X1 U5406 ( .A1(n6290), .A2(n4351), .ZN(n4381) );
  NAND2_X1 U5407 ( .A1(n4381), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4359) );
  NAND2_X1 U5408 ( .A1(n5515), .A2(DATAI_21_), .ZN(n6143) );
  INV_X1 U5409 ( .A(n6143), .ZN(n6321) );
  NOR2_X1 U5410 ( .A1(n4352), .A2(n5627), .ZN(n4356) );
  NAND2_X1 U5411 ( .A1(n6382), .A2(STATE2_REG_3__SCAN_IN), .ZN(n5148) );
  INV_X1 U5412 ( .A(n5148), .ZN(n4354) );
  NAND2_X1 U5413 ( .A1(n4383), .A2(n3109), .ZN(n4886) );
  INV_X1 U5414 ( .A(n4355), .ZN(n4384) );
  NAND2_X1 U5415 ( .A1(n4356), .A2(n4764), .ZN(n6096) );
  NAND2_X1 U5416 ( .A1(n5515), .A2(DATAI_29_), .ZN(n6264) );
  OAI22_X1 U5417 ( .A1(n4886), .A2(n4384), .B1(n6096), .B2(n6264), .ZN(n4357)
         );
  AOI21_X1 U5418 ( .B1(n6321), .B2(n4619), .A(n4357), .ZN(n4358) );
  OAI211_X1 U5419 ( .C1(n4388), .C2(n6324), .A(n4359), .B(n4358), .ZN(U3065)
         );
  NAND2_X1 U5420 ( .A1(DATAI_6_), .A2(n4701), .ZN(n6330) );
  NAND2_X1 U5421 ( .A1(n4381), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4362) );
  NAND2_X1 U5422 ( .A1(n5515), .A2(DATAI_22_), .ZN(n6147) );
  INV_X1 U5423 ( .A(n6147), .ZN(n6325) );
  NAND2_X1 U5424 ( .A1(n4383), .A2(n4276), .ZN(n4874) );
  NAND2_X1 U5425 ( .A1(n5515), .A2(DATAI_30_), .ZN(n6268) );
  OAI22_X1 U5426 ( .A1(n4874), .A2(n4384), .B1(n6096), .B2(n6268), .ZN(n4360)
         );
  AOI21_X1 U5427 ( .B1(n6325), .B2(n4619), .A(n4360), .ZN(n4361) );
  OAI211_X1 U5428 ( .C1(n4388), .C2(n6330), .A(n4362), .B(n4361), .ZN(U3066)
         );
  NAND2_X1 U5429 ( .A1(DATAI_2_), .A2(n4701), .ZN(n6306) );
  NAND2_X1 U5430 ( .A1(n4381), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4366) );
  NAND2_X1 U5431 ( .A1(n5515), .A2(DATAI_18_), .ZN(n6209) );
  INV_X1 U5432 ( .A(n6209), .ZN(n6301) );
  NAND2_X1 U5433 ( .A1(n4383), .A2(n4363), .ZN(n4894) );
  NAND2_X1 U5434 ( .A1(n5515), .A2(DATAI_26_), .ZN(n6252) );
  OAI22_X1 U5435 ( .A1(n4894), .A2(n4384), .B1(n6096), .B2(n6252), .ZN(n4364)
         );
  AOI21_X1 U5436 ( .B1(n6301), .B2(n4619), .A(n4364), .ZN(n4365) );
  OAI211_X1 U5437 ( .C1(n4388), .C2(n6306), .A(n4366), .B(n4365), .ZN(U3062)
         );
  NAND2_X1 U5438 ( .A1(DATAI_7_), .A2(n4701), .ZN(n6340) );
  NAND2_X1 U5439 ( .A1(n4381), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4369) );
  NAND2_X1 U5440 ( .A1(n5515), .A2(DATAI_23_), .ZN(n4824) );
  INV_X1 U5441 ( .A(n4824), .ZN(n6336) );
  NAND2_X1 U5442 ( .A1(n4383), .A2(n5271), .ZN(n4904) );
  NAND2_X1 U5443 ( .A1(n5515), .A2(DATAI_31_), .ZN(n6276) );
  OAI22_X1 U5444 ( .A1(n4904), .A2(n4384), .B1(n6096), .B2(n6276), .ZN(n4367)
         );
  AOI21_X1 U5445 ( .B1(n6336), .B2(n4619), .A(n4367), .ZN(n4368) );
  OAI211_X1 U5446 ( .C1(n4388), .C2(n6340), .A(n4369), .B(n4368), .ZN(U3067)
         );
  NAND2_X1 U5447 ( .A1(DATAI_4_), .A2(n4701), .ZN(n6318) );
  NAND2_X1 U5448 ( .A1(n4381), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4373) );
  NAND2_X1 U5449 ( .A1(n5515), .A2(DATAI_20_), .ZN(n6140) );
  INV_X1 U5450 ( .A(n6140), .ZN(n6315) );
  NAND2_X1 U5451 ( .A1(n4383), .A2(n4370), .ZN(n4898) );
  NAND2_X1 U5452 ( .A1(n5515), .A2(DATAI_28_), .ZN(n6260) );
  OAI22_X1 U5453 ( .A1(n4898), .A2(n4384), .B1(n6096), .B2(n6260), .ZN(n4371)
         );
  AOI21_X1 U5454 ( .B1(n6315), .B2(n4619), .A(n4371), .ZN(n4372) );
  OAI211_X1 U5455 ( .C1(n4388), .C2(n6318), .A(n4373), .B(n4372), .ZN(U3064)
         );
  NAND2_X1 U5456 ( .A1(DATAI_1_), .A2(n4701), .ZN(n6300) );
  NAND2_X1 U5457 ( .A1(n4381), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n4376) );
  NAND2_X1 U5458 ( .A1(n5515), .A2(DATAI_17_), .ZN(n6206) );
  INV_X1 U5459 ( .A(n6206), .ZN(n6295) );
  NAND2_X1 U5460 ( .A1(n4383), .A2(n4391), .ZN(n4878) );
  NAND2_X1 U5461 ( .A1(n5515), .A2(DATAI_25_), .ZN(n6248) );
  OAI22_X1 U5462 ( .A1(n4878), .A2(n4384), .B1(n6096), .B2(n6248), .ZN(n4374)
         );
  AOI21_X1 U5463 ( .B1(n6295), .B2(n4619), .A(n4374), .ZN(n4375) );
  OAI211_X1 U5464 ( .C1(n4388), .C2(n6300), .A(n4376), .B(n4375), .ZN(U3061)
         );
  NAND2_X1 U5465 ( .A1(DATAI_0_), .A2(n4701), .ZN(n6294) );
  NAND2_X1 U5466 ( .A1(n4381), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n4380) );
  NAND2_X1 U5467 ( .A1(n5515), .A2(DATAI_16_), .ZN(n6131) );
  INV_X1 U5468 ( .A(n6131), .ZN(n6291) );
  NAND2_X1 U5469 ( .A1(n4383), .A2(n4377), .ZN(n4882) );
  NAND2_X1 U5470 ( .A1(n5515), .A2(DATAI_24_), .ZN(n6244) );
  OAI22_X1 U5471 ( .A1(n4882), .A2(n4384), .B1(n6096), .B2(n6244), .ZN(n4378)
         );
  AOI21_X1 U5472 ( .B1(n6291), .B2(n4619), .A(n4378), .ZN(n4379) );
  OAI211_X1 U5473 ( .C1(n4388), .C2(n6294), .A(n4380), .B(n4379), .ZN(U3060)
         );
  NAND2_X1 U5474 ( .A1(DATAI_3_), .A2(n4701), .ZN(n6312) );
  NAND2_X1 U5475 ( .A1(n4381), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4387) );
  NAND2_X1 U5476 ( .A1(n5515), .A2(DATAI_19_), .ZN(n6213) );
  INV_X1 U5477 ( .A(n6213), .ZN(n6309) );
  NAND2_X1 U5478 ( .A1(n4383), .A2(n4382), .ZN(n4890) );
  NAND2_X1 U5479 ( .A1(n5515), .A2(DATAI_27_), .ZN(n6256) );
  OAI22_X1 U5480 ( .A1(n4890), .A2(n4384), .B1(n6096), .B2(n6256), .ZN(n4385)
         );
  AOI21_X1 U5481 ( .B1(n6309), .B2(n4619), .A(n4385), .ZN(n4386) );
  OAI211_X1 U5482 ( .C1(n4388), .C2(n6312), .A(n4387), .B(n4386), .ZN(U3063)
         );
  INV_X1 U5483 ( .A(EAX_REG_29__SCAN_IN), .ZN(n4452) );
  AOI22_X1 U5484 ( .A1(n6493), .A2(UWORD_REG_13__SCAN_IN), .B1(
        DATAO_REG_29__SCAN_IN), .B2(n5917), .ZN(n4389) );
  OAI21_X1 U5485 ( .B1(n4452), .B2(n4474), .A(n4389), .ZN(U2894) );
  INV_X1 U5486 ( .A(EAX_REG_28__SCAN_IN), .ZN(n4454) );
  AOI22_X1 U5487 ( .A1(n6493), .A2(UWORD_REG_12__SCAN_IN), .B1(
        DATAO_REG_28__SCAN_IN), .B2(n5917), .ZN(n4390) );
  OAI21_X1 U5488 ( .B1(n4454), .B2(n4474), .A(n4390), .ZN(U2895) );
  NOR2_X1 U5489 ( .A1(n4392), .A2(n4391), .ZN(n6667) );
  INV_X1 U5490 ( .A(EAX_REG_18__SCAN_IN), .ZN(n4475) );
  OAI21_X1 U5491 ( .B1(n4394), .B2(n6492), .A(n4393), .ZN(n4463) );
  NAND2_X1 U5492 ( .A1(n4463), .A2(UWORD_REG_2__SCAN_IN), .ZN(n4395) );
  NAND2_X1 U5493 ( .A1(n5936), .A2(DATAI_2_), .ZN(n4399) );
  OAI211_X1 U5494 ( .C1(n4470), .C2(n4475), .A(n4395), .B(n4399), .ZN(U2926)
         );
  INV_X1 U5495 ( .A(EAX_REG_3__SCAN_IN), .ZN(n5913) );
  NAND2_X1 U5496 ( .A1(n5936), .A2(DATAI_3_), .ZN(n4408) );
  NAND2_X1 U5497 ( .A1(n6668), .A2(LWORD_REG_3__SCAN_IN), .ZN(n4396) );
  OAI211_X1 U5498 ( .C1(n4470), .C2(n5913), .A(n4408), .B(n4396), .ZN(U2942)
         );
  NAND2_X1 U5499 ( .A1(n6668), .A2(LWORD_REG_1__SCAN_IN), .ZN(n4397) );
  NAND2_X1 U5500 ( .A1(n5936), .A2(DATAI_1_), .ZN(n4405) );
  OAI211_X1 U5501 ( .C1(n4470), .C2(n6540), .A(n4397), .B(n4405), .ZN(U2940)
         );
  INV_X1 U5502 ( .A(EAX_REG_2__SCAN_IN), .ZN(n5915) );
  NAND2_X1 U5503 ( .A1(n6668), .A2(LWORD_REG_2__SCAN_IN), .ZN(n4398) );
  OAI211_X1 U5504 ( .C1(n4470), .C2(n5915), .A(n4399), .B(n4398), .ZN(U2941)
         );
  NAND2_X1 U5505 ( .A1(n6668), .A2(UWORD_REG_0__SCAN_IN), .ZN(n4400) );
  NAND2_X1 U5506 ( .A1(n5936), .A2(DATAI_0_), .ZN(n4402) );
  OAI211_X1 U5507 ( .C1(n4470), .C2(n3696), .A(n4400), .B(n4402), .ZN(U2924)
         );
  INV_X1 U5508 ( .A(EAX_REG_0__SCAN_IN), .ZN(n5921) );
  NAND2_X1 U5509 ( .A1(n6668), .A2(LWORD_REG_0__SCAN_IN), .ZN(n4401) );
  OAI211_X1 U5510 ( .C1(n4470), .C2(n5921), .A(n4402), .B(n4401), .ZN(U2939)
         );
  NAND2_X1 U5511 ( .A1(n6668), .A2(UWORD_REG_4__SCAN_IN), .ZN(n4403) );
  NAND2_X1 U5512 ( .A1(n5936), .A2(DATAI_4_), .ZN(n4411) );
  OAI211_X1 U5513 ( .C1(n4470), .C2(n4404), .A(n4403), .B(n4411), .ZN(U2928)
         );
  NAND2_X1 U5514 ( .A1(n6668), .A2(UWORD_REG_1__SCAN_IN), .ZN(n4406) );
  OAI211_X1 U5515 ( .C1(n4470), .C2(n4407), .A(n4406), .B(n4405), .ZN(U2925)
         );
  NAND2_X1 U5516 ( .A1(n4463), .A2(UWORD_REG_3__SCAN_IN), .ZN(n4409) );
  OAI211_X1 U5517 ( .C1(n4470), .C2(n4410), .A(n4409), .B(n4408), .ZN(U2927)
         );
  INV_X1 U5518 ( .A(EAX_REG_4__SCAN_IN), .ZN(n5911) );
  NAND2_X1 U5519 ( .A1(n6668), .A2(LWORD_REG_4__SCAN_IN), .ZN(n4412) );
  OAI211_X1 U5520 ( .C1(n4470), .C2(n5911), .A(n4412), .B(n4411), .ZN(U2943)
         );
  AND2_X1 U5521 ( .A1(n6237), .A2(n3503), .ZN(n6279) );
  NAND2_X1 U5522 ( .A1(n5632), .A2(n4344), .ZN(n6121) );
  INV_X1 U5523 ( .A(n6121), .ZN(n4415) );
  INV_X1 U5524 ( .A(n4446), .ZN(n4414) );
  AOI21_X1 U5525 ( .B1(n6279), .B2(n4415), .A(n4414), .ZN(n4418) );
  INV_X1 U5526 ( .A(n4418), .ZN(n4416) );
  AOI22_X1 U5527 ( .A1(n4416), .A2(n6197), .B1(n4656), .B2(
        STATE2_REG_2__SCAN_IN), .ZN(n4450) );
  NOR2_X1 U5528 ( .A1(n4694), .A2(n4417), .ZN(n4655) );
  AOI21_X1 U5529 ( .B1(n4655), .B2(n5627), .A(n5542), .ZN(n4419) );
  NOR2_X1 U5530 ( .A1(n6286), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4697) );
  OAI21_X1 U5531 ( .B1(n4419), .B2(n4697), .A(n4418), .ZN(n4420) );
  OAI211_X1 U5532 ( .C1(n4656), .C2(n6197), .A(n6290), .B(n4420), .ZN(n4445)
         );
  NAND2_X1 U5533 ( .A1(n4445), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4424)
         );
  INV_X1 U5534 ( .A(n6252), .ZN(n6303) );
  INV_X1 U5535 ( .A(n4655), .ZN(n4421) );
  NAND2_X1 U5536 ( .A1(n5627), .A2(n4764), .ZN(n4865) );
  AND2_X1 U5537 ( .A1(n4655), .A2(n6118), .ZN(n4696) );
  OAI22_X1 U5538 ( .A1(n4894), .A2(n4446), .B1(n4729), .B2(n6209), .ZN(n4422)
         );
  AOI21_X1 U5539 ( .B1(n6303), .B2(n4663), .A(n4422), .ZN(n4423) );
  OAI211_X1 U5540 ( .C1(n4450), .C2(n6306), .A(n4424), .B(n4423), .ZN(U3142)
         );
  NAND2_X1 U5541 ( .A1(n4445), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4427)
         );
  INV_X1 U5542 ( .A(n6244), .ZN(n6283) );
  OAI22_X1 U5543 ( .A1(n4882), .A2(n4446), .B1(n4729), .B2(n6131), .ZN(n4425)
         );
  AOI21_X1 U5544 ( .B1(n6283), .B2(n4663), .A(n4425), .ZN(n4426) );
  OAI211_X1 U5545 ( .C1(n4450), .C2(n6294), .A(n4427), .B(n4426), .ZN(U3140)
         );
  NAND2_X1 U5546 ( .A1(n4445), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4430)
         );
  INV_X1 U5547 ( .A(n6260), .ZN(n6313) );
  OAI22_X1 U5548 ( .A1(n4898), .A2(n4446), .B1(n4729), .B2(n6140), .ZN(n4428)
         );
  AOI21_X1 U5549 ( .B1(n6313), .B2(n4663), .A(n4428), .ZN(n4429) );
  OAI211_X1 U5550 ( .C1(n4450), .C2(n6318), .A(n4430), .B(n4429), .ZN(U3144)
         );
  NAND2_X1 U5551 ( .A1(n4445), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4433)
         );
  INV_X1 U5552 ( .A(n6248), .ZN(n6297) );
  OAI22_X1 U5553 ( .A1(n4878), .A2(n4446), .B1(n4729), .B2(n6206), .ZN(n4431)
         );
  AOI21_X1 U5554 ( .B1(n6297), .B2(n4663), .A(n4431), .ZN(n4432) );
  OAI211_X1 U5555 ( .C1(n4450), .C2(n6300), .A(n4433), .B(n4432), .ZN(U3141)
         );
  NAND2_X1 U5556 ( .A1(n4445), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4436)
         );
  INV_X1 U5557 ( .A(n6268), .ZN(n6327) );
  OAI22_X1 U5558 ( .A1(n4874), .A2(n4446), .B1(n4729), .B2(n6147), .ZN(n4434)
         );
  AOI21_X1 U5559 ( .B1(n6327), .B2(n4663), .A(n4434), .ZN(n4435) );
  OAI211_X1 U5560 ( .C1(n4450), .C2(n6330), .A(n4436), .B(n4435), .ZN(U3146)
         );
  NAND2_X1 U5561 ( .A1(n4445), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4439)
         );
  INV_X1 U5562 ( .A(n6276), .ZN(n6331) );
  OAI22_X1 U5563 ( .A1(n4904), .A2(n4446), .B1(n4729), .B2(n4824), .ZN(n4437)
         );
  AOI21_X1 U5564 ( .B1(n6331), .B2(n4663), .A(n4437), .ZN(n4438) );
  OAI211_X1 U5565 ( .C1(n4450), .C2(n6340), .A(n4439), .B(n4438), .ZN(U3147)
         );
  NAND2_X1 U5566 ( .A1(n4445), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4442)
         );
  INV_X1 U5567 ( .A(n6264), .ZN(n6319) );
  OAI22_X1 U5568 ( .A1(n4886), .A2(n4446), .B1(n4729), .B2(n6143), .ZN(n4440)
         );
  AOI21_X1 U5569 ( .B1(n6319), .B2(n4663), .A(n4440), .ZN(n4441) );
  OAI211_X1 U5570 ( .C1(n4450), .C2(n6324), .A(n4442), .B(n4441), .ZN(U3145)
         );
  INV_X1 U5571 ( .A(EAX_REG_30__SCAN_IN), .ZN(n4459) );
  AOI22_X1 U5572 ( .A1(n6493), .A2(UWORD_REG_14__SCAN_IN), .B1(n5917), .B2(
        DATAO_REG_30__SCAN_IN), .ZN(n4443) );
  OAI21_X1 U5573 ( .B1(n4459), .B2(n4474), .A(n4443), .ZN(U2893) );
  AOI22_X1 U5574 ( .A1(n6493), .A2(UWORD_REG_9__SCAN_IN), .B1(n5917), .B2(
        DATAO_REG_25__SCAN_IN), .ZN(n4444) );
  OAI21_X1 U5575 ( .B1(n3804), .B2(n4474), .A(n4444), .ZN(U2898) );
  NAND2_X1 U5576 ( .A1(n4445), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4449)
         );
  INV_X1 U5577 ( .A(n6256), .ZN(n6307) );
  OAI22_X1 U5578 ( .A1(n4890), .A2(n4446), .B1(n4729), .B2(n6213), .ZN(n4447)
         );
  AOI21_X1 U5579 ( .B1(n6307), .B2(n4663), .A(n4447), .ZN(n4448) );
  OAI211_X1 U5580 ( .C1(n4450), .C2(n6312), .A(n4449), .B(n4448), .ZN(U3143)
         );
  AOI22_X1 U5581 ( .A1(n4463), .A2(UWORD_REG_13__SCAN_IN), .B1(n5936), .B2(
        DATAI_13_), .ZN(n4451) );
  OAI21_X1 U5582 ( .B1(n4452), .B2(n4470), .A(n4451), .ZN(U2937) );
  AOI22_X1 U5583 ( .A1(n4463), .A2(UWORD_REG_12__SCAN_IN), .B1(n5936), .B2(
        DATAI_12_), .ZN(n4453) );
  OAI21_X1 U5584 ( .B1(n4454), .B2(n4470), .A(n4453), .ZN(U2936) );
  AOI22_X1 U5585 ( .A1(n4463), .A2(UWORD_REG_11__SCAN_IN), .B1(n5936), .B2(
        DATAI_11_), .ZN(n4455) );
  OAI21_X1 U5586 ( .B1(n4456), .B2(n4470), .A(n4455), .ZN(U2935) );
  AOI22_X1 U5587 ( .A1(n4463), .A2(UWORD_REG_9__SCAN_IN), .B1(n5936), .B2(
        DATAI_9_), .ZN(n4457) );
  OAI21_X1 U5588 ( .B1(n3804), .B2(n4470), .A(n4457), .ZN(U2933) );
  AOI22_X1 U5589 ( .A1(n4463), .A2(UWORD_REG_14__SCAN_IN), .B1(n5936), .B2(
        DATAI_14_), .ZN(n4458) );
  OAI21_X1 U5590 ( .B1(n4459), .B2(n4470), .A(n4458), .ZN(U2938) );
  AOI22_X1 U5591 ( .A1(n4463), .A2(UWORD_REG_7__SCAN_IN), .B1(n5936), .B2(
        DATAI_7_), .ZN(n4460) );
  OAI21_X1 U5592 ( .B1(n4461), .B2(n4470), .A(n4460), .ZN(U2931) );
  INV_X1 U5593 ( .A(EAX_REG_15__SCAN_IN), .ZN(n5890) );
  AOI22_X1 U5594 ( .A1(n4463), .A2(LWORD_REG_15__SCAN_IN), .B1(n5936), .B2(
        DATAI_15_), .ZN(n4462) );
  OAI21_X1 U5595 ( .B1(n5890), .B2(n4470), .A(n4462), .ZN(U2954) );
  AOI22_X1 U5596 ( .A1(n4463), .A2(UWORD_REG_8__SCAN_IN), .B1(n5936), .B2(
        DATAI_8_), .ZN(n4464) );
  OAI21_X1 U5597 ( .B1(n3902), .B2(n4470), .A(n4464), .ZN(U2932) );
  INV_X1 U5598 ( .A(DATAI_5_), .ZN(n4617) );
  NOR2_X1 U5599 ( .A1(n5928), .A2(n4617), .ZN(n4468) );
  AOI21_X1 U5600 ( .B1(LWORD_REG_5__SCAN_IN), .B2(n6668), .A(n4468), .ZN(n4465) );
  OAI21_X1 U5601 ( .B1(n4614), .B2(n4470), .A(n4465), .ZN(U2944) );
  AOI22_X1 U5602 ( .A1(n6668), .A2(UWORD_REG_6__SCAN_IN), .B1(n5936), .B2(
        DATAI_6_), .ZN(n4466) );
  OAI21_X1 U5603 ( .B1(n4467), .B2(n4470), .A(n4466), .ZN(U2930) );
  AOI21_X1 U5604 ( .B1(UWORD_REG_5__SCAN_IN), .B2(n6668), .A(n4468), .ZN(n4469) );
  OAI21_X1 U5605 ( .B1(n4471), .B2(n4470), .A(n4469), .ZN(U2929) );
  AOI22_X1 U5606 ( .A1(n6493), .A2(UWORD_REG_0__SCAN_IN), .B1(
        DATAO_REG_16__SCAN_IN), .B2(n5917), .ZN(n4472) );
  OAI21_X1 U5607 ( .B1(n3696), .B2(n4474), .A(n4472), .ZN(U2907) );
  AOI22_X1 U5608 ( .A1(n6493), .A2(UWORD_REG_2__SCAN_IN), .B1(
        DATAO_REG_18__SCAN_IN), .B2(n5917), .ZN(n4473) );
  OAI21_X1 U5609 ( .B1(n4475), .B2(n4474), .A(n4473), .ZN(U2905) );
  XOR2_X1 U5610 ( .A(n4477), .B(n4476), .Z(n5959) );
  INV_X1 U5611 ( .A(n5959), .ZN(n4484) );
  AOI22_X1 U5612 ( .A1(n5060), .A2(DATAI_3_), .B1(n5884), .B2(
        EAX_REG_3__SCAN_IN), .ZN(n4478) );
  OAI21_X1 U5613 ( .B1(n4484), .B2(n5718), .A(n4478), .ZN(U2888) );
  OAI21_X1 U5614 ( .B1(n4481), .B2(n4480), .A(n4479), .ZN(n4482) );
  AND2_X1 U5615 ( .A1(n4482), .A2(n4555), .ZN(n6033) );
  AOI22_X1 U5616 ( .A1(n5415), .A2(n6033), .B1(n5414), .B2(EBX_REG_3__SCAN_IN), 
        .ZN(n4483) );
  OAI21_X1 U5617 ( .B1(n4484), .B2(n5417), .A(n4483), .ZN(U2856) );
  OR2_X1 U5618 ( .A1(n4486), .A2(n4485), .ZN(n4487) );
  XNOR2_X1 U5619 ( .A(n4487), .B(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n5851)
         );
  INV_X1 U5620 ( .A(n4505), .ZN(n5758) );
  NAND2_X1 U5621 ( .A1(n5851), .A2(n5758), .ZN(n4500) );
  AND2_X1 U5622 ( .A1(n5302), .A2(n5289), .ZN(n4496) );
  NAND2_X1 U5623 ( .A1(n5280), .A2(n4184), .ZN(n4489) );
  NAND2_X1 U5624 ( .A1(n4489), .A2(n4488), .ZN(n4491) );
  NAND2_X1 U5625 ( .A1(n4491), .A2(n4490), .ZN(n4492) );
  NAND2_X1 U5626 ( .A1(n4492), .A2(n6492), .ZN(n4494) );
  OAI21_X1 U5627 ( .B1(n5302), .B2(n4494), .A(n4493), .ZN(n4495) );
  OR2_X1 U5628 ( .A1(n6349), .A2(n4498), .ZN(n4499) );
  NAND2_X1 U5629 ( .A1(n4500), .A2(n4499), .ZN(n4502) );
  INV_X1 U5630 ( .A(FLUSH_REG_SCAN_IN), .ZN(n5771) );
  NAND2_X1 U5631 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n5771), .ZN(n4533) );
  NOR2_X1 U5632 ( .A1(n4533), .A2(n4498), .ZN(n4501) );
  AOI21_X1 U5633 ( .B1(n4502), .B2(n6391), .A(n4501), .ZN(n4539) );
  NAND4_X1 U5634 ( .A1(n4184), .A2(n4506), .A3(n4505), .A4(n4504), .ZN(n4507)
         );
  OR2_X1 U5635 ( .A1(n4508), .A2(n4507), .ZN(n6344) );
  NAND2_X1 U5636 ( .A1(n6237), .A2(n6344), .ZN(n4524) );
  INV_X1 U5637 ( .A(n4519), .ZN(n4510) );
  OAI21_X1 U5638 ( .B1(n4509), .B2(n3275), .A(n4510), .ZN(n4511) );
  NOR2_X1 U5639 ( .A1(n4511), .A2(n3925), .ZN(n5638) );
  INV_X1 U5640 ( .A(n4512), .ZN(n4513) );
  OR2_X1 U5641 ( .A1(n5289), .A2(n4513), .ZN(n4530) );
  INV_X1 U5642 ( .A(n4509), .ZN(n5150) );
  NAND2_X1 U5643 ( .A1(n5150), .A2(n5156), .ZN(n4515) );
  NAND2_X1 U5644 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4516) );
  INV_X1 U5645 ( .A(n4516), .ZN(n4514) );
  AOI22_X1 U5646 ( .A1(n4530), .A2(n4515), .B1(n6347), .B2(n4514), .ZN(n4518)
         );
  NAND2_X1 U5647 ( .A1(n6347), .A2(n4516), .ZN(n4517) );
  MUX2_X1 U5648 ( .A(n4518), .B(n4517), .S(INSTQUEUERD_ADDR_REG_3__SCAN_IN), 
        .Z(n4521) );
  NAND2_X1 U5649 ( .A1(n5150), .A2(n4519), .ZN(n4520) );
  OAI211_X1 U5650 ( .C1(n5638), .C2(n4527), .A(n4521), .B(n4520), .ZN(n4522)
         );
  INV_X1 U5651 ( .A(n4522), .ZN(n4523) );
  NAND2_X1 U5652 ( .A1(n4524), .A2(n4523), .ZN(n6342) );
  NAND2_X1 U5653 ( .A1(n5632), .A2(n6344), .ZN(n4532) );
  XNOR2_X1 U5654 ( .A(n4509), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4529)
         );
  XNOR2_X1 U5655 ( .A(n5288), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4525)
         );
  NAND2_X1 U5656 ( .A1(n6347), .A2(n4525), .ZN(n4526) );
  OAI21_X1 U5657 ( .B1(n4529), .B2(n4527), .A(n4526), .ZN(n4528) );
  AOI21_X1 U5658 ( .B1(n4530), .B2(n4529), .A(n4528), .ZN(n4531) );
  NAND2_X1 U5659 ( .A1(n4532), .A2(n4531), .ZN(n5151) );
  NAND4_X1 U5660 ( .A1(n6342), .A2(n6391), .A3(n6349), .A4(n5151), .ZN(n4537)
         );
  OAI21_X1 U5661 ( .B1(n6349), .B2(STATE2_REG_1__SCAN_IN), .A(n4533), .ZN(
        n4535) );
  NAND2_X1 U5662 ( .A1(n4535), .A2(n4534), .ZN(n4536) );
  AND2_X1 U5663 ( .A1(n4537), .A2(n4536), .ZN(n4538) );
  AND2_X1 U5664 ( .A1(n4539), .A2(n4538), .ZN(n6365) );
  AOI21_X1 U5665 ( .B1(n4539), .B2(n4503), .A(n6365), .ZN(n4547) );
  NOR2_X1 U5666 ( .A1(n4547), .A2(FLUSH_REG_SCAN_IN), .ZN(n4540) );
  NAND2_X1 U5667 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n6388), .ZN(n6468) );
  OAI21_X1 U5668 ( .B1(n4540), .B2(n6468), .A(n6165), .ZN(n6055) );
  AND2_X1 U5669 ( .A1(n4655), .A2(n4541), .ZN(n6277) );
  INV_X1 U5670 ( .A(n4694), .ZN(n5631) );
  INV_X1 U5671 ( .A(n6191), .ZN(n6193) );
  NOR2_X1 U5672 ( .A1(n6277), .A2(n6193), .ZN(n4543) );
  AND2_X1 U5673 ( .A1(n6119), .A2(n6192), .ZN(n6120) );
  INV_X1 U5674 ( .A(n6120), .ZN(n4542) );
  AOI21_X1 U5675 ( .B1(n4543), .B2(n4542), .A(n6286), .ZN(n4545) );
  INV_X1 U5676 ( .A(n4697), .ZN(n6163) );
  INV_X1 U5677 ( .A(n6237), .ZN(n6229) );
  AND2_X1 U5678 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6470), .ZN(n5633) );
  OAI22_X1 U5679 ( .A1(n4695), .A2(n6163), .B1(n6229), .B2(n5633), .ZN(n4544)
         );
  OAI21_X1 U5680 ( .B1(n4545), .B2(n4544), .A(n6055), .ZN(n4546) );
  OAI21_X1 U5681 ( .B1(n6055), .B2(n6358), .A(n4546), .ZN(U3462) );
  INV_X1 U5682 ( .A(n4547), .ZN(n4548) );
  NAND2_X1 U5683 ( .A1(n4548), .A2(n6388), .ZN(n6381) );
  INV_X1 U5684 ( .A(n6381), .ZN(n4550) );
  OAI22_X1 U5685 ( .A1(n4764), .A2(n6286), .B1(n6346), .B2(n5633), .ZN(n4549)
         );
  OAI21_X1 U5686 ( .B1(n4550), .B2(n4549), .A(n6055), .ZN(n4551) );
  OAI21_X1 U5687 ( .B1(n6055), .B2(n6635), .A(n4551), .ZN(U3465) );
  INV_X1 U5688 ( .A(n4612), .ZN(n4561) );
  AOI21_X1 U5689 ( .B1(n4553), .B2(n4552), .A(n4561), .ZN(n4798) );
  INV_X1 U5690 ( .A(n4798), .ZN(n5858) );
  AND2_X1 U5691 ( .A1(n4555), .A2(n4554), .ZN(n4556) );
  OR2_X1 U5692 ( .A1(n4556), .A2(n4610), .ZN(n6025) );
  INV_X1 U5693 ( .A(n6025), .ZN(n4557) );
  AOI22_X1 U5694 ( .A1(n5415), .A2(n4557), .B1(n5414), .B2(EBX_REG_4__SCAN_IN), 
        .ZN(n4558) );
  OAI21_X1 U5695 ( .B1(n5858), .B2(n5417), .A(n4558), .ZN(U2855) );
  INV_X1 U5696 ( .A(DATAI_4_), .ZN(n4559) );
  OAI222_X1 U5697 ( .A1(n5858), .A2(n5718), .B1(n4616), .B2(n4559), .C1(n5435), 
        .C2(n5911), .ZN(U2887) );
  AOI21_X1 U5698 ( .B1(n4561), .B2(n4611), .A(n4560), .ZN(n4562) );
  OR2_X1 U5699 ( .A1(n4562), .A2(n4747), .ZN(n4800) );
  AOI22_X1 U5700 ( .A1(n5060), .A2(DATAI_6_), .B1(n5884), .B2(
        EAX_REG_6__SCAN_IN), .ZN(n4563) );
  OAI21_X1 U5701 ( .B1(n4800), .B2(n5718), .A(n4563), .ZN(U2885) );
  CLKBUF_X1 U5702 ( .A(n4564), .Z(n4751) );
  NAND2_X1 U5703 ( .A1(n4608), .A2(n4565), .ZN(n4566) );
  NAND2_X1 U5704 ( .A1(n4751), .A2(n4566), .ZN(n4973) );
  INV_X1 U5705 ( .A(n4973), .ZN(n4579) );
  AOI22_X1 U5706 ( .A1(n4579), .A2(n5415), .B1(n5414), .B2(EBX_REG_6__SCAN_IN), 
        .ZN(n4567) );
  OAI21_X1 U5707 ( .B1(n4800), .B2(n5417), .A(n4567), .ZN(U2853) );
  OAI21_X1 U5708 ( .B1(n4570), .B2(n4569), .A(n4568), .ZN(n4806) );
  INV_X1 U5709 ( .A(REIP_REG_6__SCAN_IN), .ZN(n4981) );
  NOR2_X1 U5710 ( .A1(n6047), .A2(n4981), .ZN(n4802) );
  INV_X1 U5711 ( .A(n4571), .ZN(n4572) );
  NAND2_X1 U5712 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n4572), .ZN(n6054)
         );
  OAI21_X1 U5713 ( .B1(n5964), .B2(n6054), .A(n5598), .ZN(n6014) );
  INV_X1 U5714 ( .A(n6014), .ZN(n6027) );
  NOR2_X1 U5715 ( .A1(n6027), .A2(n4575), .ZN(n4577) );
  INV_X1 U5716 ( .A(n4573), .ZN(n6042) );
  INV_X1 U5717 ( .A(n5086), .ZN(n4574) );
  OAI21_X1 U5718 ( .B1(n4949), .B2(n6042), .A(n4574), .ZN(n6049) );
  AOI21_X1 U5719 ( .B1(n4575), .B2(n5194), .A(n6049), .ZN(n6021) );
  INV_X1 U5720 ( .A(n6021), .ZN(n4576) );
  MUX2_X1 U5721 ( .A(n4577), .B(n4576), .S(INSTADDRPOINTER_REG_6__SCAN_IN), 
        .Z(n4578) );
  AOI211_X1 U5722 ( .C1(n6044), .C2(n4579), .A(n4802), .B(n4578), .ZN(n4580)
         );
  OAI21_X1 U5723 ( .B1(n6023), .B2(n4806), .A(n4580), .ZN(U3012) );
  NOR2_X1 U5724 ( .A1(n6191), .A2(n5627), .ZN(n4588) );
  NAND2_X1 U5725 ( .A1(n4588), .A2(n6232), .ZN(n4820) );
  OR2_X1 U5726 ( .A1(n5632), .A2(n4344), .ZN(n6155) );
  INV_X1 U5727 ( .A(n6155), .ZN(n4581) );
  NAND3_X1 U5728 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n4864), .A3(n4699), .ZN(n6160) );
  NOR2_X1 U5729 ( .A1(n6635), .A2(n6160), .ZN(n4605) );
  AOI21_X1 U5730 ( .B1(n6279), .B2(n4581), .A(n4605), .ZN(n4587) );
  OR2_X1 U5731 ( .A1(n6191), .A2(n4582), .ZN(n4583) );
  NAND2_X1 U5732 ( .A1(n4583), .A2(n6197), .ZN(n4586) );
  INV_X1 U5733 ( .A(n4586), .ZN(n4584) );
  AOI22_X1 U5734 ( .A1(n4587), .A2(n4584), .B1(n6286), .B2(n6160), .ZN(n4585)
         );
  NAND2_X1 U5735 ( .A1(n6290), .A2(n4585), .ZN(n4604) );
  INV_X1 U5736 ( .A(n6312), .ZN(n6253) );
  OAI22_X1 U5737 ( .A1(n4587), .A2(n4586), .B1(n6379), .B2(n6160), .ZN(n4603)
         );
  AOI22_X1 U5738 ( .A1(INSTQUEUE_REG_9__3__SCAN_IN), .A2(n4604), .B1(n6253), 
        .B2(n4603), .ZN(n4590) );
  INV_X1 U5739 ( .A(n4890), .ZN(n6308) );
  AOI22_X1 U5740 ( .A1(n6308), .A2(n4605), .B1(n6184), .B2(n6307), .ZN(n4589)
         );
  OAI211_X1 U5741 ( .C1(n4820), .C2(n6213), .A(n4590), .B(n4589), .ZN(U3095)
         );
  INV_X1 U5742 ( .A(n6294), .ZN(n6231) );
  AOI22_X1 U5743 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n4604), .B1(n6231), 
        .B2(n4603), .ZN(n4592) );
  INV_X1 U5744 ( .A(n4882), .ZN(n6284) );
  AOI22_X1 U5745 ( .A1(n6284), .A2(n4605), .B1(n6184), .B2(n6283), .ZN(n4591)
         );
  OAI211_X1 U5746 ( .C1(n4820), .C2(n6131), .A(n4592), .B(n4591), .ZN(U3092)
         );
  INV_X1 U5747 ( .A(n6330), .ZN(n6265) );
  AOI22_X1 U5748 ( .A1(INSTQUEUE_REG_9__6__SCAN_IN), .A2(n4604), .B1(n6265), 
        .B2(n4603), .ZN(n4594) );
  INV_X1 U5749 ( .A(n4874), .ZN(n6326) );
  AOI22_X1 U5750 ( .A1(n6326), .A2(n4605), .B1(n6184), .B2(n6327), .ZN(n4593)
         );
  OAI211_X1 U5751 ( .C1(n4820), .C2(n6147), .A(n4594), .B(n4593), .ZN(U3098)
         );
  INV_X1 U5752 ( .A(n6306), .ZN(n6249) );
  AOI22_X1 U5753 ( .A1(INSTQUEUE_REG_9__2__SCAN_IN), .A2(n4604), .B1(n6249), 
        .B2(n4603), .ZN(n4596) );
  INV_X1 U5754 ( .A(n4894), .ZN(n6302) );
  AOI22_X1 U5755 ( .A1(n6302), .A2(n4605), .B1(n6184), .B2(n6303), .ZN(n4595)
         );
  OAI211_X1 U5756 ( .C1(n4820), .C2(n6209), .A(n4596), .B(n4595), .ZN(U3094)
         );
  INV_X1 U5757 ( .A(n6340), .ZN(n6271) );
  AOI22_X1 U5758 ( .A1(INSTQUEUE_REG_9__7__SCAN_IN), .A2(n4604), .B1(n6271), 
        .B2(n4603), .ZN(n4598) );
  INV_X1 U5759 ( .A(n4904), .ZN(n6334) );
  AOI22_X1 U5760 ( .A1(n6334), .A2(n4605), .B1(n6184), .B2(n6331), .ZN(n4597)
         );
  OAI211_X1 U5761 ( .C1(n4820), .C2(n4824), .A(n4598), .B(n4597), .ZN(U3099)
         );
  INV_X1 U5762 ( .A(n6318), .ZN(n6257) );
  AOI22_X1 U5763 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n4604), .B1(n6257), 
        .B2(n4603), .ZN(n4600) );
  INV_X1 U5764 ( .A(n4898), .ZN(n6314) );
  AOI22_X1 U5765 ( .A1(n6314), .A2(n4605), .B1(n6184), .B2(n6313), .ZN(n4599)
         );
  OAI211_X1 U5766 ( .C1(n4820), .C2(n6140), .A(n4600), .B(n4599), .ZN(U3096)
         );
  INV_X1 U5767 ( .A(n6300), .ZN(n6245) );
  AOI22_X1 U5768 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(n4604), .B1(n6245), 
        .B2(n4603), .ZN(n4602) );
  INV_X1 U5769 ( .A(n4878), .ZN(n6296) );
  AOI22_X1 U5770 ( .A1(n6296), .A2(n4605), .B1(n6184), .B2(n6297), .ZN(n4601)
         );
  OAI211_X1 U5771 ( .C1(n4820), .C2(n6206), .A(n4602), .B(n4601), .ZN(U3093)
         );
  INV_X1 U5772 ( .A(n6324), .ZN(n6261) );
  AOI22_X1 U5773 ( .A1(INSTQUEUE_REG_9__5__SCAN_IN), .A2(n4604), .B1(n6261), 
        .B2(n4603), .ZN(n4607) );
  INV_X1 U5774 ( .A(n4886), .ZN(n6320) );
  AOI22_X1 U5775 ( .A1(n6320), .A2(n4605), .B1(n6184), .B2(n6319), .ZN(n4606)
         );
  OAI211_X1 U5776 ( .C1(n4820), .C2(n6143), .A(n4607), .B(n4606), .ZN(U3097)
         );
  OAI21_X1 U5777 ( .B1(n4610), .B2(n4609), .A(n4608), .ZN(n5842) );
  XNOR2_X1 U5778 ( .A(n4612), .B(n4611), .ZN(n5951) );
  INV_X1 U5779 ( .A(n5951), .ZN(n4615) );
  OAI222_X1 U5780 ( .A1(n5842), .A2(n5428), .B1(n5417), .B2(n4615), .C1(n4613), 
        .C2(n5427), .ZN(U2854) );
  OAI222_X1 U5781 ( .A1(n4617), .A2(n4616), .B1(n5718), .B2(n4615), .C1(n4614), 
        .C2(n5435), .ZN(U2886) );
  INV_X1 U5782 ( .A(n4865), .ZN(n4618) );
  NAND2_X1 U5783 ( .A1(n6119), .A2(n4618), .ZN(n6154) );
  OAI21_X1 U5784 ( .B1(n4619), .B2(n6144), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n4620) );
  NAND3_X1 U5785 ( .A1(n6121), .A2(n6197), .A3(n4620), .ZN(n4622) );
  OR2_X1 U5786 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6126), .ZN(n4648)
         );
  AND2_X1 U5787 ( .A1(n4623), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6156) );
  OAI21_X1 U5788 ( .B1(n4700), .B2(n6379), .A(n4701), .ZN(n4815) );
  AOI211_X1 U5789 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n4648), .A(n6156), .B(
        n4815), .ZN(n4621) );
  NAND3_X1 U5790 ( .A1(n6358), .A2(n4622), .A3(n4621), .ZN(n4647) );
  NAND2_X1 U5791 ( .A1(n4647), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4628) );
  OR2_X1 U5792 ( .A1(n6121), .A2(n6286), .ZN(n4662) );
  OR2_X1 U5793 ( .A1(n4662), .A2(n6237), .ZN(n4625) );
  NOR2_X1 U5794 ( .A1(n4623), .A2(n6379), .ZN(n4816) );
  AND2_X1 U5795 ( .A1(n4700), .A2(n6358), .ZN(n4872) );
  NAND2_X1 U5796 ( .A1(n4816), .A2(n4872), .ZN(n4624) );
  NAND2_X1 U5797 ( .A1(n4625), .A2(n4624), .ZN(n4650) );
  OAI22_X1 U5798 ( .A1(n4904), .A2(n4648), .B1(n4824), .B2(n6154), .ZN(n4626)
         );
  AOI21_X1 U5799 ( .B1(n6271), .B2(n4650), .A(n4626), .ZN(n4627) );
  OAI211_X1 U5800 ( .C1(n4653), .C2(n6276), .A(n4628), .B(n4627), .ZN(U3075)
         );
  NAND2_X1 U5801 ( .A1(n4647), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n4631) );
  OAI22_X1 U5802 ( .A1(n4878), .A2(n4648), .B1(n6206), .B2(n6154), .ZN(n4629)
         );
  AOI21_X1 U5803 ( .B1(n6245), .B2(n4650), .A(n4629), .ZN(n4630) );
  OAI211_X1 U5804 ( .C1(n4653), .C2(n6248), .A(n4631), .B(n4630), .ZN(U3069)
         );
  NAND2_X1 U5805 ( .A1(n4647), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n4634) );
  OAI22_X1 U5806 ( .A1(n4890), .A2(n4648), .B1(n6213), .B2(n6154), .ZN(n4632)
         );
  AOI21_X1 U5807 ( .B1(n6253), .B2(n4650), .A(n4632), .ZN(n4633) );
  OAI211_X1 U5808 ( .C1(n4653), .C2(n6256), .A(n4634), .B(n4633), .ZN(U3071)
         );
  NAND2_X1 U5809 ( .A1(n4647), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n4637) );
  OAI22_X1 U5810 ( .A1(n4882), .A2(n4648), .B1(n6131), .B2(n6154), .ZN(n4635)
         );
  AOI21_X1 U5811 ( .B1(n6231), .B2(n4650), .A(n4635), .ZN(n4636) );
  OAI211_X1 U5812 ( .C1(n4653), .C2(n6244), .A(n4637), .B(n4636), .ZN(U3068)
         );
  NAND2_X1 U5813 ( .A1(n4647), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n4640) );
  OAI22_X1 U5814 ( .A1(n4898), .A2(n4648), .B1(n6140), .B2(n6154), .ZN(n4638)
         );
  AOI21_X1 U5815 ( .B1(n6257), .B2(n4650), .A(n4638), .ZN(n4639) );
  OAI211_X1 U5816 ( .C1(n4653), .C2(n6260), .A(n4640), .B(n4639), .ZN(U3072)
         );
  NAND2_X1 U5817 ( .A1(n4647), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n4643) );
  OAI22_X1 U5818 ( .A1(n4894), .A2(n4648), .B1(n6209), .B2(n6154), .ZN(n4641)
         );
  AOI21_X1 U5819 ( .B1(n6249), .B2(n4650), .A(n4641), .ZN(n4642) );
  OAI211_X1 U5820 ( .C1(n4653), .C2(n6252), .A(n4643), .B(n4642), .ZN(U3070)
         );
  NAND2_X1 U5821 ( .A1(n4647), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n4646) );
  OAI22_X1 U5822 ( .A1(n4874), .A2(n4648), .B1(n6147), .B2(n6154), .ZN(n4644)
         );
  AOI21_X1 U5823 ( .B1(n6265), .B2(n4650), .A(n4644), .ZN(n4645) );
  OAI211_X1 U5824 ( .C1(n4653), .C2(n6268), .A(n4646), .B(n4645), .ZN(U3074)
         );
  NAND2_X1 U5825 ( .A1(n4647), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4652) );
  OAI22_X1 U5826 ( .A1(n4886), .A2(n4648), .B1(n6143), .B2(n6154), .ZN(n4649)
         );
  AOI21_X1 U5827 ( .B1(n6261), .B2(n4650), .A(n4649), .ZN(n4651) );
  OAI211_X1 U5828 ( .C1(n4653), .C2(n6264), .A(n4652), .B(n4651), .ZN(U3073)
         );
  INV_X1 U5829 ( .A(n5627), .ZN(n4654) );
  NAND2_X1 U5830 ( .A1(n4655), .A2(n4654), .ZN(n6233) );
  INV_X1 U5831 ( .A(n4656), .ZN(n4657) );
  NOR2_X1 U5832 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4657), .ZN(n4664)
         );
  NOR3_X1 U5833 ( .A1(n4815), .A2(n6358), .A3(n6156), .ZN(n4660) );
  OAI21_X1 U5834 ( .B1(n6335), .B2(n4663), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n4658) );
  NAND3_X1 U5835 ( .A1(n6121), .A2(n6197), .A3(n4658), .ZN(n4659) );
  OAI211_X1 U5836 ( .C1(n4664), .C2(n6470), .A(n4660), .B(n4659), .ZN(n4686)
         );
  NAND2_X1 U5837 ( .A1(n4686), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4667)
         );
  INV_X1 U5838 ( .A(n4816), .ZN(n6227) );
  INV_X1 U5839 ( .A(n4700), .ZN(n6158) );
  NOR2_X1 U5840 ( .A1(n6158), .A2(n6358), .ZN(n4814) );
  INV_X1 U5841 ( .A(n4814), .ZN(n4661) );
  OAI22_X1 U5842 ( .A1(n4662), .A2(n6229), .B1(n6227), .B2(n4661), .ZN(n4690)
         );
  INV_X1 U5843 ( .A(n4664), .ZN(n4687) );
  OAI22_X1 U5844 ( .A1(n4688), .A2(n6209), .B1(n4894), .B2(n4687), .ZN(n4665)
         );
  AOI21_X1 U5845 ( .B1(n6249), .B2(n4690), .A(n4665), .ZN(n4666) );
  OAI211_X1 U5846 ( .C1(n4693), .C2(n6252), .A(n4667), .B(n4666), .ZN(U3134)
         );
  NAND2_X1 U5847 ( .A1(n4686), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4670)
         );
  OAI22_X1 U5848 ( .A1(n4688), .A2(n6143), .B1(n4886), .B2(n4687), .ZN(n4668)
         );
  AOI21_X1 U5849 ( .B1(n6261), .B2(n4690), .A(n4668), .ZN(n4669) );
  OAI211_X1 U5850 ( .C1(n4693), .C2(n6264), .A(n4670), .B(n4669), .ZN(U3137)
         );
  NAND2_X1 U5851 ( .A1(n4686), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4673)
         );
  OAI22_X1 U5852 ( .A1(n4688), .A2(n4824), .B1(n4904), .B2(n4687), .ZN(n4671)
         );
  AOI21_X1 U5853 ( .B1(n6271), .B2(n4690), .A(n4671), .ZN(n4672) );
  OAI211_X1 U5854 ( .C1(n4693), .C2(n6276), .A(n4673), .B(n4672), .ZN(U3139)
         );
  NAND2_X1 U5855 ( .A1(n4686), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4676)
         );
  OAI22_X1 U5856 ( .A1(n4688), .A2(n6147), .B1(n4874), .B2(n4687), .ZN(n4674)
         );
  AOI21_X1 U5857 ( .B1(n6265), .B2(n4690), .A(n4674), .ZN(n4675) );
  OAI211_X1 U5858 ( .C1(n4693), .C2(n6268), .A(n4676), .B(n4675), .ZN(U3138)
         );
  NAND2_X1 U5859 ( .A1(n4686), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4679)
         );
  OAI22_X1 U5860 ( .A1(n4688), .A2(n6140), .B1(n4898), .B2(n4687), .ZN(n4677)
         );
  AOI21_X1 U5861 ( .B1(n6257), .B2(n4690), .A(n4677), .ZN(n4678) );
  OAI211_X1 U5862 ( .C1(n4693), .C2(n6260), .A(n4679), .B(n4678), .ZN(U3136)
         );
  NAND2_X1 U5863 ( .A1(n4686), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4682)
         );
  OAI22_X1 U5864 ( .A1(n4882), .A2(n4687), .B1(n6131), .B2(n4688), .ZN(n4680)
         );
  AOI21_X1 U5865 ( .B1(n6231), .B2(n4690), .A(n4680), .ZN(n4681) );
  OAI211_X1 U5866 ( .C1(n4693), .C2(n6244), .A(n4682), .B(n4681), .ZN(U3132)
         );
  NAND2_X1 U5867 ( .A1(n4686), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n4685)
         );
  OAI22_X1 U5868 ( .A1(n4688), .A2(n6206), .B1(n4878), .B2(n4687), .ZN(n4683)
         );
  AOI21_X1 U5869 ( .B1(n6245), .B2(n4690), .A(n4683), .ZN(n4684) );
  OAI211_X1 U5870 ( .C1(n4693), .C2(n6248), .A(n4685), .B(n4684), .ZN(U3133)
         );
  NAND2_X1 U5871 ( .A1(n4686), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4692)
         );
  OAI22_X1 U5872 ( .A1(n4688), .A2(n6213), .B1(n4890), .B2(n4687), .ZN(n4689)
         );
  AOI21_X1 U5873 ( .B1(n6253), .B2(n4690), .A(n4689), .ZN(n4691) );
  OAI211_X1 U5874 ( .C1(n4693), .C2(n6256), .A(n4692), .B(n4691), .ZN(U3135)
         );
  NAND2_X1 U5875 ( .A1(n4695), .A2(n4694), .ZN(n6057) );
  NOR2_X1 U5876 ( .A1(n6155), .A2(n6237), .ZN(n4757) );
  NOR2_X1 U5877 ( .A1(n4696), .A2(n6286), .ZN(n4698) );
  AOI21_X1 U5878 ( .B1(n4698), .B2(n4785), .A(n4697), .ZN(n4703) );
  NAND3_X1 U5879 ( .A1(n6358), .A2(n4864), .A3(n4699), .ZN(n4761) );
  OR2_X1 U5880 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4761), .ZN(n4730)
         );
  NOR2_X1 U5881 ( .A1(n4700), .A2(n6157), .ZN(n6088) );
  OAI21_X1 U5882 ( .B1(n6088), .B2(n6379), .A(n4701), .ZN(n6094) );
  AOI211_X1 U5883 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n4730), .A(n4816), .B(
        n6094), .ZN(n4702) );
  OAI21_X1 U5884 ( .B1(n4757), .B2(n4703), .A(n4702), .ZN(n4728) );
  NAND2_X1 U5885 ( .A1(n4728), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4709) );
  INV_X1 U5886 ( .A(n4757), .ZN(n4704) );
  OR2_X1 U5887 ( .A1(n4704), .A2(n6286), .ZN(n4706) );
  NAND2_X1 U5888 ( .A1(n6088), .A2(n6156), .ZN(n4705) );
  NAND2_X1 U5889 ( .A1(n4706), .A2(n4705), .ZN(n4732) );
  OAI22_X1 U5890 ( .A1(n4878), .A2(n4730), .B1(n4729), .B2(n6248), .ZN(n4707)
         );
  AOI21_X1 U5891 ( .B1(n6245), .B2(n4732), .A(n4707), .ZN(n4708) );
  OAI211_X1 U5892 ( .C1(n4785), .C2(n6206), .A(n4709), .B(n4708), .ZN(U3021)
         );
  NAND2_X1 U5893 ( .A1(n4728), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4712) );
  OAI22_X1 U5894 ( .A1(n4894), .A2(n4730), .B1(n4729), .B2(n6252), .ZN(n4710)
         );
  AOI21_X1 U5895 ( .B1(n6249), .B2(n4732), .A(n4710), .ZN(n4711) );
  OAI211_X1 U5896 ( .C1(n4785), .C2(n6209), .A(n4712), .B(n4711), .ZN(U3022)
         );
  NAND2_X1 U5897 ( .A1(n4728), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4715) );
  OAI22_X1 U5898 ( .A1(n4882), .A2(n4730), .B1(n6244), .B2(n4729), .ZN(n4713)
         );
  AOI21_X1 U5899 ( .B1(n6231), .B2(n4732), .A(n4713), .ZN(n4714) );
  OAI211_X1 U5900 ( .C1(n4785), .C2(n6131), .A(n4715), .B(n4714), .ZN(U3020)
         );
  NAND2_X1 U5901 ( .A1(n4728), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4718) );
  OAI22_X1 U5902 ( .A1(n4890), .A2(n4730), .B1(n4729), .B2(n6256), .ZN(n4716)
         );
  AOI21_X1 U5903 ( .B1(n6253), .B2(n4732), .A(n4716), .ZN(n4717) );
  OAI211_X1 U5904 ( .C1(n4785), .C2(n6213), .A(n4718), .B(n4717), .ZN(U3023)
         );
  NAND2_X1 U5905 ( .A1(n4728), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4721) );
  OAI22_X1 U5906 ( .A1(n4898), .A2(n4730), .B1(n4729), .B2(n6260), .ZN(n4719)
         );
  AOI21_X1 U5907 ( .B1(n6257), .B2(n4732), .A(n4719), .ZN(n4720) );
  OAI211_X1 U5908 ( .C1(n4785), .C2(n6140), .A(n4721), .B(n4720), .ZN(U3024)
         );
  NAND2_X1 U5909 ( .A1(n4728), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4724) );
  OAI22_X1 U5910 ( .A1(n4886), .A2(n4730), .B1(n4729), .B2(n6264), .ZN(n4722)
         );
  AOI21_X1 U5911 ( .B1(n6261), .B2(n4732), .A(n4722), .ZN(n4723) );
  OAI211_X1 U5912 ( .C1(n4785), .C2(n6143), .A(n4724), .B(n4723), .ZN(U3025)
         );
  NAND2_X1 U5913 ( .A1(n4728), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4727) );
  OAI22_X1 U5914 ( .A1(n4904), .A2(n4730), .B1(n4729), .B2(n6276), .ZN(n4725)
         );
  AOI21_X1 U5915 ( .B1(n6271), .B2(n4732), .A(n4725), .ZN(n4726) );
  OAI211_X1 U5916 ( .C1(n4785), .C2(n4824), .A(n4727), .B(n4726), .ZN(U3027)
         );
  NAND2_X1 U5917 ( .A1(n4728), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4734) );
  OAI22_X1 U5918 ( .A1(n4874), .A2(n4730), .B1(n4729), .B2(n6268), .ZN(n4731)
         );
  AOI21_X1 U5919 ( .B1(n6265), .B2(n4732), .A(n4731), .ZN(n4733) );
  OAI211_X1 U5920 ( .C1(n4785), .C2(n6147), .A(n4734), .B(n4733), .ZN(U3026)
         );
  CLKBUF_X1 U5921 ( .A(n4735), .Z(n4736) );
  OAI21_X1 U5922 ( .B1(n4736), .B2(n4737), .A(n4809), .ZN(n5001) );
  AOI22_X1 U5923 ( .A1(n5060), .A2(DATAI_8_), .B1(n5884), .B2(
        EAX_REG_8__SCAN_IN), .ZN(n4738) );
  OAI21_X1 U5924 ( .B1(n5001), .B2(n5718), .A(n4738), .ZN(U2883) );
  NOR2_X1 U5925 ( .A1(n4753), .A2(n4741), .ZN(n4742) );
  OR2_X1 U5926 ( .A1(n4739), .A2(n4742), .ZN(n6000) );
  INV_X1 U5927 ( .A(EBX_REG_8__SCAN_IN), .ZN(n4743) );
  OAI22_X1 U5928 ( .A1(n6000), .A2(n5428), .B1(n4743), .B2(n5427), .ZN(n4744)
         );
  INV_X1 U5929 ( .A(n4744), .ZN(n4745) );
  OAI21_X1 U5930 ( .B1(n5001), .B2(n5417), .A(n4745), .ZN(U2851) );
  INV_X1 U5931 ( .A(n4746), .ZN(n4749) );
  INV_X1 U5932 ( .A(n4747), .ZN(n4748) );
  AOI21_X1 U5933 ( .B1(n4749), .B2(n4748), .A(n4736), .ZN(n5943) );
  INV_X1 U5934 ( .A(n5943), .ZN(n4756) );
  AND2_X1 U5935 ( .A1(n4751), .A2(n4750), .ZN(n4752) );
  NOR2_X1 U5936 ( .A1(n4753), .A2(n4752), .ZN(n6007) );
  AOI22_X1 U5937 ( .A1(n6007), .A2(n5415), .B1(EBX_REG_7__SCAN_IN), .B2(n5414), 
        .ZN(n4754) );
  OAI21_X1 U5938 ( .B1(n4756), .B2(n5417), .A(n4754), .ZN(U2852) );
  AOI22_X1 U5939 ( .A1(n5060), .A2(DATAI_7_), .B1(n5884), .B2(
        EAX_REG_7__SCAN_IN), .ZN(n4755) );
  OAI21_X1 U5940 ( .B1(n4756), .B2(n5718), .A(n4755), .ZN(U2884) );
  NOR2_X1 U5941 ( .A1(n6635), .A2(n4761), .ZN(n4782) );
  AOI21_X1 U5942 ( .B1(n4757), .B2(n3503), .A(n4782), .ZN(n4762) );
  OR2_X1 U5943 ( .A1(n4765), .A2(n6234), .ZN(n4758) );
  AOI22_X1 U5944 ( .A1(n4762), .A2(n4760), .B1(n6286), .B2(n4761), .ZN(n4759)
         );
  NAND2_X1 U5945 ( .A1(n6290), .A2(n4759), .ZN(n4781) );
  INV_X1 U5946 ( .A(n4760), .ZN(n4763) );
  OAI22_X1 U5947 ( .A1(n4763), .A2(n4762), .B1(n6379), .B2(n4761), .ZN(n4780)
         );
  AOI22_X1 U5948 ( .A1(INSTQUEUE_REG_1__4__SCAN_IN), .A2(n4781), .B1(n6257), 
        .B2(n4780), .ZN(n4767) );
  AOI22_X1 U5949 ( .A1(n6314), .A2(n4782), .B1(n4866), .B2(n6315), .ZN(n4766)
         );
  OAI211_X1 U5950 ( .C1(n6260), .C2(n4785), .A(n4767), .B(n4766), .ZN(U3032)
         );
  AOI22_X1 U5951 ( .A1(INSTQUEUE_REG_1__3__SCAN_IN), .A2(n4781), .B1(n6253), 
        .B2(n4780), .ZN(n4769) );
  AOI22_X1 U5952 ( .A1(n6308), .A2(n4782), .B1(n4866), .B2(n6309), .ZN(n4768)
         );
  OAI211_X1 U5953 ( .C1(n6256), .C2(n4785), .A(n4769), .B(n4768), .ZN(U3031)
         );
  AOI22_X1 U5954 ( .A1(INSTQUEUE_REG_1__1__SCAN_IN), .A2(n4781), .B1(n6245), 
        .B2(n4780), .ZN(n4771) );
  AOI22_X1 U5955 ( .A1(n6296), .A2(n4782), .B1(n4866), .B2(n6295), .ZN(n4770)
         );
  OAI211_X1 U5956 ( .C1(n6248), .C2(n4785), .A(n4771), .B(n4770), .ZN(U3029)
         );
  AOI22_X1 U5957 ( .A1(INSTQUEUE_REG_1__7__SCAN_IN), .A2(n4781), .B1(n6271), 
        .B2(n4780), .ZN(n4773) );
  AOI22_X1 U5958 ( .A1(n6334), .A2(n4782), .B1(n4866), .B2(n6336), .ZN(n4772)
         );
  OAI211_X1 U5959 ( .C1(n6276), .C2(n4785), .A(n4773), .B(n4772), .ZN(U3035)
         );
  AOI22_X1 U5960 ( .A1(INSTQUEUE_REG_1__2__SCAN_IN), .A2(n4781), .B1(n6249), 
        .B2(n4780), .ZN(n4775) );
  AOI22_X1 U5961 ( .A1(n6302), .A2(n4782), .B1(n4866), .B2(n6301), .ZN(n4774)
         );
  OAI211_X1 U5962 ( .C1(n6252), .C2(n4785), .A(n4775), .B(n4774), .ZN(U3030)
         );
  AOI22_X1 U5963 ( .A1(INSTQUEUE_REG_1__0__SCAN_IN), .A2(n4781), .B1(n6231), 
        .B2(n4780), .ZN(n4777) );
  AOI22_X1 U5964 ( .A1(n6284), .A2(n4782), .B1(n4866), .B2(n6291), .ZN(n4776)
         );
  OAI211_X1 U5965 ( .C1(n6244), .C2(n4785), .A(n4777), .B(n4776), .ZN(U3028)
         );
  AOI22_X1 U5966 ( .A1(INSTQUEUE_REG_1__5__SCAN_IN), .A2(n4781), .B1(n6261), 
        .B2(n4780), .ZN(n4779) );
  AOI22_X1 U5967 ( .A1(n6320), .A2(n4782), .B1(n4866), .B2(n6321), .ZN(n4778)
         );
  OAI211_X1 U5968 ( .C1(n6264), .C2(n4785), .A(n4779), .B(n4778), .ZN(U3033)
         );
  AOI22_X1 U5969 ( .A1(INSTQUEUE_REG_1__6__SCAN_IN), .A2(n4781), .B1(n6265), 
        .B2(n4780), .ZN(n4784) );
  AOI22_X1 U5970 ( .A1(n6326), .A2(n4782), .B1(n4866), .B2(n6325), .ZN(n4783)
         );
  OAI211_X1 U5971 ( .C1(n6268), .C2(n4785), .A(n4784), .B(n4783), .ZN(U3034)
         );
  INV_X1 U5972 ( .A(n5020), .ZN(n4789) );
  NOR2_X1 U5973 ( .A1(n6047), .A2(n6580), .ZN(n4786) );
  AOI21_X1 U5974 ( .B1(n5963), .B2(PHYADDRPOINTER_REG_1__SCAN_IN), .A(n4786), 
        .ZN(n4787) );
  OAI21_X1 U5975 ( .B1(n5973), .B2(PHYADDRPOINTER_REG_1__SCAN_IN), .A(n4787), 
        .ZN(n4788) );
  AOI21_X1 U5976 ( .B1(n4789), .B2(n5515), .A(n4788), .ZN(n4790) );
  OAI21_X1 U5977 ( .B1(n4791), .B2(n5770), .A(n4790), .ZN(U2985) );
  OAI21_X1 U5978 ( .B1(n4794), .B2(n4793), .A(n4792), .ZN(n6022) );
  INV_X1 U5979 ( .A(n4795), .ZN(n5856) );
  AOI22_X1 U5980 ( .A1(n5963), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .B1(n6032), 
        .B2(REIP_REG_4__SCAN_IN), .ZN(n4796) );
  OAI21_X1 U5981 ( .B1(n5973), .B2(n5856), .A(n4796), .ZN(n4797) );
  AOI21_X1 U5982 ( .B1(n4798), .B2(n5515), .A(n4797), .ZN(n4799) );
  OAI21_X1 U5983 ( .B1(n5770), .B2(n6022), .A(n4799), .ZN(U2982) );
  INV_X1 U5984 ( .A(n4800), .ZN(n4979) );
  INV_X1 U5985 ( .A(n4801), .ZN(n4977) );
  AOI21_X1 U5986 ( .B1(n5963), .B2(PHYADDRPOINTER_REG_6__SCAN_IN), .A(n4802), 
        .ZN(n4803) );
  OAI21_X1 U5987 ( .B1(n5973), .B2(n4977), .A(n4803), .ZN(n4804) );
  AOI21_X1 U5988 ( .B1(n4979), .B2(n5515), .A(n4804), .ZN(n4805) );
  OAI21_X1 U5989 ( .B1(n4806), .B2(n5770), .A(n4805), .ZN(U2980) );
  NAND2_X1 U5990 ( .A1(n4809), .A2(n4808), .ZN(n4810) );
  NAND2_X1 U5991 ( .A1(n4919), .A2(n4810), .ZN(n4928) );
  AOI22_X1 U5992 ( .A1(n5060), .A2(DATAI_9_), .B1(n5884), .B2(
        EAX_REG_9__SCAN_IN), .ZN(n4811) );
  OAI21_X1 U5993 ( .B1(n4928), .B2(n5718), .A(n4811), .ZN(U2882) );
  NAND2_X1 U5994 ( .A1(n4820), .A2(n6226), .ZN(n4812) );
  AOI21_X1 U5995 ( .B1(n4812), .B2(STATEBS16_REG_SCAN_IN), .A(n6286), .ZN(
        n4818) );
  OR2_X1 U5996 ( .A1(n5628), .A2(n5632), .ZN(n4867) );
  INV_X1 U5997 ( .A(n4867), .ZN(n4813) );
  AND2_X1 U5998 ( .A1(n4813), .A2(n6237), .ZN(n6194) );
  AOI22_X1 U5999 ( .A1(n4818), .A2(n6194), .B1(n6156), .B2(n4814), .ZN(n4849)
         );
  NOR2_X1 U6000 ( .A1(n4816), .A2(n4815), .ZN(n4870) );
  INV_X1 U6001 ( .A(n6194), .ZN(n4817) );
  NAND3_X1 U6002 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n4864), .ZN(n6199) );
  OR2_X1 U6003 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6199), .ZN(n4844)
         );
  AOI22_X1 U6004 ( .A1(n4818), .A2(n4817), .B1(STATE2_REG_3__SCAN_IN), .B2(
        n4844), .ZN(n4819) );
  OAI211_X1 U6005 ( .C1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C2(n6379), .A(n4870), .B(n4819), .ZN(n4843) );
  NAND2_X1 U6006 ( .A1(n4843), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n4823)
         );
  INV_X1 U6007 ( .A(n4820), .ZN(n4846) );
  OAI22_X1 U6008 ( .A1(n4882), .A2(n4844), .B1(n6226), .B2(n6131), .ZN(n4821)
         );
  AOI21_X1 U6009 ( .B1(n4846), .B2(n6283), .A(n4821), .ZN(n4822) );
  OAI211_X1 U6010 ( .C1(n4849), .C2(n6294), .A(n4823), .B(n4822), .ZN(U3100)
         );
  NAND2_X1 U6011 ( .A1(n4843), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n4827)
         );
  OAI22_X1 U6012 ( .A1(n4904), .A2(n4844), .B1(n6226), .B2(n4824), .ZN(n4825)
         );
  AOI21_X1 U6013 ( .B1(n4846), .B2(n6331), .A(n4825), .ZN(n4826) );
  OAI211_X1 U6014 ( .C1(n4849), .C2(n6340), .A(n4827), .B(n4826), .ZN(U3107)
         );
  NAND2_X1 U6015 ( .A1(n4843), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n4830)
         );
  OAI22_X1 U6016 ( .A1(n4874), .A2(n4844), .B1(n6226), .B2(n6147), .ZN(n4828)
         );
  AOI21_X1 U6017 ( .B1(n4846), .B2(n6327), .A(n4828), .ZN(n4829) );
  OAI211_X1 U6018 ( .C1(n4849), .C2(n6330), .A(n4830), .B(n4829), .ZN(U3106)
         );
  NAND2_X1 U6019 ( .A1(n4843), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n4833)
         );
  OAI22_X1 U6020 ( .A1(n4886), .A2(n4844), .B1(n6226), .B2(n6143), .ZN(n4831)
         );
  AOI21_X1 U6021 ( .B1(n4846), .B2(n6319), .A(n4831), .ZN(n4832) );
  OAI211_X1 U6022 ( .C1(n4849), .C2(n6324), .A(n4833), .B(n4832), .ZN(U3105)
         );
  NAND2_X1 U6023 ( .A1(n4843), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n4836)
         );
  OAI22_X1 U6024 ( .A1(n4898), .A2(n4844), .B1(n6226), .B2(n6140), .ZN(n4834)
         );
  AOI21_X1 U6025 ( .B1(n4846), .B2(n6313), .A(n4834), .ZN(n4835) );
  OAI211_X1 U6026 ( .C1(n4849), .C2(n6318), .A(n4836), .B(n4835), .ZN(U3104)
         );
  NAND2_X1 U6027 ( .A1(n4843), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n4839)
         );
  OAI22_X1 U6028 ( .A1(n4890), .A2(n4844), .B1(n6226), .B2(n6213), .ZN(n4837)
         );
  AOI21_X1 U6029 ( .B1(n4846), .B2(n6307), .A(n4837), .ZN(n4838) );
  OAI211_X1 U6030 ( .C1(n4849), .C2(n6312), .A(n4839), .B(n4838), .ZN(U3103)
         );
  NAND2_X1 U6031 ( .A1(n4843), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n4842)
         );
  OAI22_X1 U6032 ( .A1(n4894), .A2(n4844), .B1(n6226), .B2(n6209), .ZN(n4840)
         );
  AOI21_X1 U6033 ( .B1(n4846), .B2(n6303), .A(n4840), .ZN(n4841) );
  OAI211_X1 U6034 ( .C1(n4849), .C2(n6306), .A(n4842), .B(n4841), .ZN(U3102)
         );
  NAND2_X1 U6035 ( .A1(n4843), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n4848)
         );
  OAI22_X1 U6036 ( .A1(n4878), .A2(n4844), .B1(n6226), .B2(n6206), .ZN(n4845)
         );
  AOI21_X1 U6037 ( .B1(n4846), .B2(n6297), .A(n4845), .ZN(n4847) );
  OAI211_X1 U6038 ( .C1(n4849), .C2(n6300), .A(n4848), .B(n4847), .ZN(U3101)
         );
  INV_X1 U6039 ( .A(n4850), .ZN(n4853) );
  INV_X1 U6040 ( .A(n4739), .ZN(n4852) );
  INV_X1 U6041 ( .A(n4851), .ZN(n4934) );
  AOI21_X1 U6042 ( .B1(n4853), .B2(n4852), .A(n4934), .ZN(n5992) );
  INV_X1 U6043 ( .A(n5992), .ZN(n4854) );
  OAI222_X1 U6044 ( .A1(n4928), .A2(n5417), .B1(n5427), .B2(n4855), .C1(n5428), 
        .C2(n4854), .ZN(U2850) );
  OAI21_X1 U6045 ( .B1(n4858), .B2(n4857), .A(n4856), .ZN(n5999) );
  INV_X1 U6046 ( .A(n5001), .ZN(n4862) );
  INV_X1 U6047 ( .A(n4859), .ZN(n4996) );
  AOI22_X1 U6048 ( .A1(n5963), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .B1(n6032), 
        .B2(REIP_REG_8__SCAN_IN), .ZN(n4860) );
  OAI21_X1 U6049 ( .B1(n5973), .B2(n4996), .A(n4860), .ZN(n4861) );
  AOI21_X1 U6050 ( .B1(n4862), .B2(n5515), .A(n4861), .ZN(n4863) );
  OAI21_X1 U6051 ( .B1(n5999), .B2(n5770), .A(n4863), .ZN(U2978) );
  NAND3_X1 U6052 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n6358), .A3(n4864), .ZN(n6063) );
  NOR2_X1 U6053 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6063), .ZN(n4873)
         );
  OR2_X1 U6054 ( .A1(n6057), .A2(n4865), .ZN(n6087) );
  OAI21_X1 U6055 ( .B1(n4866), .B2(n6072), .A(n6163), .ZN(n4869) );
  NOR2_X1 U6056 ( .A1(n4867), .A2(n6237), .ZN(n6059) );
  INV_X1 U6057 ( .A(n6059), .ZN(n4868) );
  NAND2_X1 U6058 ( .A1(n4869), .A2(n4868), .ZN(n4871) );
  OAI221_X1 U6059 ( .B1(n4873), .B2(n6470), .C1(n4873), .C2(n4871), .A(n4870), 
        .ZN(n4902) );
  NAND2_X1 U6060 ( .A1(n4902), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4877) );
  AOI22_X1 U6061 ( .A1(n6059), .A2(n6197), .B1(n6156), .B2(n4872), .ZN(n4905)
         );
  INV_X1 U6062 ( .A(n4873), .ZN(n4903) );
  OAI22_X1 U6063 ( .A1(n6330), .A2(n4905), .B1(n4874), .B2(n4903), .ZN(n4875)
         );
  AOI21_X1 U6064 ( .B1(n6325), .B2(n6072), .A(n4875), .ZN(n4876) );
  OAI211_X1 U6065 ( .C1(n4909), .C2(n6268), .A(n4877), .B(n4876), .ZN(U3042)
         );
  NAND2_X1 U6066 ( .A1(n4902), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4881) );
  OAI22_X1 U6067 ( .A1(n6300), .A2(n4905), .B1(n4878), .B2(n4903), .ZN(n4879)
         );
  AOI21_X1 U6068 ( .B1(n6295), .B2(n6072), .A(n4879), .ZN(n4880) );
  OAI211_X1 U6069 ( .C1(n4909), .C2(n6248), .A(n4881), .B(n4880), .ZN(U3037)
         );
  NAND2_X1 U6070 ( .A1(n4902), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4885) );
  OAI22_X1 U6071 ( .A1(n6294), .A2(n4905), .B1(n4882), .B2(n4903), .ZN(n4883)
         );
  AOI21_X1 U6072 ( .B1(n6291), .B2(n6072), .A(n4883), .ZN(n4884) );
  OAI211_X1 U6073 ( .C1(n6244), .C2(n4909), .A(n4885), .B(n4884), .ZN(U3036)
         );
  NAND2_X1 U6074 ( .A1(n4902), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4889) );
  OAI22_X1 U6075 ( .A1(n6324), .A2(n4905), .B1(n4886), .B2(n4903), .ZN(n4887)
         );
  AOI21_X1 U6076 ( .B1(n6321), .B2(n6072), .A(n4887), .ZN(n4888) );
  OAI211_X1 U6077 ( .C1(n4909), .C2(n6264), .A(n4889), .B(n4888), .ZN(U3041)
         );
  NAND2_X1 U6078 ( .A1(n4902), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4893) );
  OAI22_X1 U6079 ( .A1(n6312), .A2(n4905), .B1(n4890), .B2(n4903), .ZN(n4891)
         );
  AOI21_X1 U6080 ( .B1(n6309), .B2(n6072), .A(n4891), .ZN(n4892) );
  OAI211_X1 U6081 ( .C1(n4909), .C2(n6256), .A(n4893), .B(n4892), .ZN(U3039)
         );
  NAND2_X1 U6082 ( .A1(n4902), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4897) );
  OAI22_X1 U6083 ( .A1(n6306), .A2(n4905), .B1(n4894), .B2(n4903), .ZN(n4895)
         );
  AOI21_X1 U6084 ( .B1(n6301), .B2(n6072), .A(n4895), .ZN(n4896) );
  OAI211_X1 U6085 ( .C1(n4909), .C2(n6252), .A(n4897), .B(n4896), .ZN(U3038)
         );
  NAND2_X1 U6086 ( .A1(n4902), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4901) );
  OAI22_X1 U6087 ( .A1(n6318), .A2(n4905), .B1(n4898), .B2(n4903), .ZN(n4899)
         );
  AOI21_X1 U6088 ( .B1(n6315), .B2(n6072), .A(n4899), .ZN(n4900) );
  OAI211_X1 U6089 ( .C1(n4909), .C2(n6260), .A(n4901), .B(n4900), .ZN(U3040)
         );
  NAND2_X1 U6090 ( .A1(n4902), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4908) );
  OAI22_X1 U6091 ( .A1(n6340), .A2(n4905), .B1(n4904), .B2(n4903), .ZN(n4906)
         );
  AOI21_X1 U6092 ( .B1(n6336), .B2(n6072), .A(n4906), .ZN(n4907) );
  OAI211_X1 U6093 ( .C1(n4909), .C2(n6276), .A(n4908), .B(n4907), .ZN(U3043)
         );
  NAND2_X1 U6094 ( .A1(n4912), .A2(n4911), .ZN(n4913) );
  XNOR2_X1 U6095 ( .A(n4910), .B(n4913), .ZN(n5994) );
  INV_X1 U6096 ( .A(n5770), .ZN(n5968) );
  NAND2_X1 U6097 ( .A1(n5994), .A2(n5968), .ZN(n4917) );
  INV_X1 U6098 ( .A(REIP_REG_9__SCAN_IN), .ZN(n4914) );
  NOR2_X1 U6099 ( .A1(n6047), .A2(n4914), .ZN(n5991) );
  NOR2_X1 U6100 ( .A1(n5973), .A2(n4932), .ZN(n4915) );
  AOI211_X1 U6101 ( .C1(n5963), .C2(PHYADDRPOINTER_REG_9__SCAN_IN), .A(n5991), 
        .B(n4915), .ZN(n4916) );
  OAI211_X1 U6102 ( .C1(n5542), .C2(n4928), .A(n4917), .B(n4916), .ZN(U2977)
         );
  AND2_X1 U6103 ( .A1(n4919), .A2(n4918), .ZN(n4920) );
  OR2_X1 U6104 ( .A1(n4920), .A2(n4937), .ZN(n5827) );
  AOI22_X1 U6105 ( .A1(n5060), .A2(DATAI_10_), .B1(n5884), .B2(
        EAX_REG_10__SCAN_IN), .ZN(n4921) );
  OAI21_X1 U6106 ( .B1(n5827), .B2(n5718), .A(n4921), .ZN(U2881) );
  INV_X1 U6107 ( .A(n5818), .ZN(n4927) );
  NOR2_X1 U6108 ( .A1(n5853), .A2(n4922), .ZN(n5821) );
  INV_X1 U6109 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n4925) );
  AOI22_X1 U6110 ( .A1(EBX_REG_9__SCAN_IN), .A2(n5865), .B1(n5866), .B2(n5992), 
        .ZN(n4924) );
  NAND2_X1 U6111 ( .A1(n5016), .A2(n4923), .ZN(n5854) );
  OAI211_X1 U6112 ( .C1(n5834), .C2(n4925), .A(n4924), .B(n5854), .ZN(n4926)
         );
  AOI221_X1 U6113 ( .B1(n4927), .B2(n4914), .C1(n5821), .C2(
        REIP_REG_9__SCAN_IN), .A(n4926), .ZN(n4931) );
  INV_X1 U6114 ( .A(n4928), .ZN(n4929) );
  NAND2_X1 U6115 ( .A1(n4929), .A2(n5838), .ZN(n4930) );
  OAI211_X1 U6116 ( .C1(n5868), .C2(n4932), .A(n4931), .B(n4930), .ZN(U2818)
         );
  INV_X1 U6117 ( .A(EBX_REG_10__SCAN_IN), .ZN(n4935) );
  OAI21_X1 U6118 ( .B1(n4934), .B2(n4933), .A(n4939), .ZN(n5822) );
  OAI222_X1 U6119 ( .A1(n5827), .A2(n5417), .B1(n5427), .B2(n4935), .C1(n5428), 
        .C2(n5822), .ZN(U2849) );
  OAI21_X1 U6120 ( .B1(n4937), .B2(n4936), .A(n4984), .ZN(n5355) );
  AOI22_X1 U6121 ( .A1(n5060), .A2(DATAI_11_), .B1(n5884), .B2(
        EAX_REG_11__SCAN_IN), .ZN(n4938) );
  OAI21_X1 U6122 ( .B1(n5355), .B2(n5718), .A(n4938), .ZN(U2880) );
  AOI21_X1 U6123 ( .B1(n4940), .B2(n4939), .A(n4989), .ZN(n5983) );
  AOI22_X1 U6124 ( .A1(n5983), .A2(n5415), .B1(n5414), .B2(EBX_REG_11__SCAN_IN), .ZN(n4941) );
  OAI21_X1 U6125 ( .B1(n5355), .B2(n5417), .A(n4941), .ZN(U2848) );
  NAND2_X1 U6126 ( .A1(n4963), .A2(n4942), .ZN(n4944) );
  XOR2_X1 U6127 ( .A(n4944), .B(n4943), .Z(n5033) );
  NAND2_X1 U6128 ( .A1(n4947), .A2(n6014), .ZN(n6008) );
  NOR2_X1 U6129 ( .A1(n4945), .A2(n6008), .ZN(n5993) );
  OAI211_X1 U6130 ( .C1(INSTADDRPOINTER_REG_9__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .A(n5993), .B(n4946), .ZN(n4953) );
  OAI22_X1 U6131 ( .A1(n4949), .A2(n4948), .B1(n4947), .B2(n5598), .ZN(n4950)
         );
  NOR2_X1 U6132 ( .A1(n5086), .A2(n4950), .ZN(n6013) );
  OAI21_X1 U6133 ( .B1(n6001), .B2(n5601), .A(n6013), .ZN(n5990) );
  INV_X1 U6134 ( .A(REIP_REG_10__SCAN_IN), .ZN(n6427) );
  OAI22_X1 U6135 ( .A1(n5822), .A2(n6024), .B1(n6427), .B2(n6047), .ZN(n4951)
         );
  AOI21_X1 U6136 ( .B1(n5990), .B2(INSTADDRPOINTER_REG_10__SCAN_IN), .A(n4951), 
        .ZN(n4952) );
  OAI211_X1 U6137 ( .C1(n5033), .C2(n6023), .A(n4953), .B(n4952), .ZN(U3008)
         );
  NOR2_X1 U6138 ( .A1(n5301), .A2(n4955), .ZN(n4954) );
  OR2_X1 U6139 ( .A1(n5838), .A2(n4954), .ZN(n5874) );
  INV_X1 U6140 ( .A(n5874), .ZN(n5857) );
  NOR2_X1 U6141 ( .A1(n4956), .A2(n4955), .ZN(n5850) );
  INV_X1 U6142 ( .A(n5850), .ZN(n5872) );
  NOR2_X1 U6143 ( .A1(n6346), .A2(n5872), .ZN(n4959) );
  OAI22_X1 U6144 ( .A1(n4957), .A2(n5863), .B1(n5662), .B2(n6652), .ZN(n4958)
         );
  AOI211_X1 U6145 ( .C1(n5330), .C2(REIP_REG_0__SCAN_IN), .A(n4959), .B(n4958), 
        .ZN(n4961) );
  OAI21_X1 U6146 ( .B1(n5870), .B2(n5813), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n4960) );
  OAI211_X1 U6147 ( .C1(n4962), .C2(n5857), .A(n4961), .B(n4960), .ZN(U2827)
         );
  NAND2_X1 U6148 ( .A1(n4964), .A2(n4963), .ZN(n4966) );
  XNOR2_X1 U6149 ( .A(n3422), .B(n5988), .ZN(n4965) );
  XNOR2_X1 U6150 ( .A(n4966), .B(n4965), .ZN(n5985) );
  NAND2_X1 U6151 ( .A1(n5985), .A2(n5968), .ZN(n4970) );
  INV_X1 U6152 ( .A(REIP_REG_11__SCAN_IN), .ZN(n4967) );
  NOR2_X1 U6153 ( .A1(n6047), .A2(n4967), .ZN(n5982) );
  NOR2_X1 U6154 ( .A1(n5973), .A2(n5347), .ZN(n4968) );
  AOI211_X1 U6155 ( .C1(n5963), .C2(PHYADDRPOINTER_REG_11__SCAN_IN), .A(n5982), 
        .B(n4968), .ZN(n4969) );
  OAI211_X1 U6156 ( .C1(n5542), .C2(n5355), .A(n4970), .B(n4969), .ZN(U2975)
         );
  INV_X1 U6157 ( .A(REIP_REG_5__SCAN_IN), .ZN(n6421) );
  INV_X1 U6158 ( .A(REIP_REG_4__SCAN_IN), .ZN(n6419) );
  NOR2_X1 U6159 ( .A1(n6421), .A2(n6419), .ZN(n4971) );
  AOI21_X1 U6160 ( .B1(n5852), .B2(n4971), .A(n5853), .ZN(n5847) );
  INV_X1 U6161 ( .A(n5847), .ZN(n4982) );
  NAND3_X1 U6162 ( .A1(n4993), .A2(REIP_REG_5__SCAN_IN), .A3(
        REIP_REG_4__SCAN_IN), .ZN(n5835) );
  NOR2_X1 U6163 ( .A1(REIP_REG_6__SCAN_IN), .A2(n5835), .ZN(n5839) );
  OAI21_X1 U6164 ( .B1(n5834), .B2(n6571), .A(n5854), .ZN(n4975) );
  OAI22_X1 U6165 ( .A1(n6633), .A2(n5662), .B1(n5863), .B2(n4973), .ZN(n4974)
         );
  NOR3_X1 U6166 ( .A1(n5839), .A2(n4975), .A3(n4974), .ZN(n4976) );
  OAI21_X1 U6167 ( .B1(n4977), .B2(n5868), .A(n4976), .ZN(n4978) );
  AOI21_X1 U6168 ( .B1(n5838), .B2(n4979), .A(n4978), .ZN(n4980) );
  OAI21_X1 U6169 ( .B1(n4982), .B2(n4981), .A(n4980), .ZN(U2821) );
  AOI21_X1 U6170 ( .B1(n4985), .B2(n4984), .A(n4983), .ZN(n5814) );
  INV_X1 U6171 ( .A(n5814), .ZN(n4992) );
  AOI22_X1 U6172 ( .A1(n5060), .A2(DATAI_12_), .B1(n5884), .B2(
        EAX_REG_12__SCAN_IN), .ZN(n4986) );
  OAI21_X1 U6173 ( .B1(n4992), .B2(n5718), .A(n4986), .ZN(U2879) );
  INV_X1 U6174 ( .A(EBX_REG_12__SCAN_IN), .ZN(n4991) );
  CLKBUF_X1 U6175 ( .A(n4987), .Z(n5039) );
  OR2_X1 U6176 ( .A1(n4989), .A2(n4988), .ZN(n4990) );
  NAND2_X1 U6177 ( .A1(n5039), .A2(n4990), .ZN(n5976) );
  OAI222_X1 U6178 ( .A1(n4992), .A2(n5417), .B1(n5427), .B2(n4991), .C1(n5976), 
        .C2(n5428), .ZN(U2847) );
  INV_X1 U6179 ( .A(n4993), .ZN(n5855) );
  OAI21_X1 U6180 ( .B1(n5855), .B2(n4994), .A(n6424), .ZN(n4999) );
  INV_X1 U6181 ( .A(n5854), .ZN(n5845) );
  AOI21_X1 U6182 ( .B1(n5865), .B2(EBX_REG_8__SCAN_IN), .A(n5845), .ZN(n4995)
         );
  OAI21_X1 U6183 ( .B1(n5868), .B2(n4996), .A(n4995), .ZN(n4998) );
  OAI22_X1 U6184 ( .A1(n6636), .A2(n5834), .B1(n5863), .B2(n6000), .ZN(n4997)
         );
  AOI211_X1 U6185 ( .C1(n5821), .C2(n4999), .A(n4998), .B(n4997), .ZN(n5000)
         );
  OAI21_X1 U6186 ( .B1(n5826), .B2(n5001), .A(n5000), .ZN(U2819) );
  NOR2_X1 U6187 ( .A1(n5003), .A2(REIP_REG_1__SCAN_IN), .ZN(n5012) );
  NOR2_X1 U6188 ( .A1(n5002), .A2(n5012), .ZN(n5864) );
  NOR3_X1 U6189 ( .A1(n5003), .A2(REIP_REG_2__SCAN_IN), .A3(n6580), .ZN(n5004)
         );
  AOI21_X1 U6190 ( .B1(n5865), .B2(EBX_REG_2__SCAN_IN), .A(n5004), .ZN(n5006)
         );
  NAND2_X1 U6191 ( .A1(n6043), .A2(n5866), .ZN(n5005) );
  OAI211_X1 U6192 ( .C1(n5864), .C2(n6416), .A(n5006), .B(n5005), .ZN(n5009)
         );
  INV_X1 U6193 ( .A(PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n5007) );
  OAI22_X1 U6194 ( .A1(n5972), .A2(n5868), .B1(n5834), .B2(n5007), .ZN(n5008)
         );
  AOI211_X1 U6195 ( .C1(n5632), .C2(n5850), .A(n5009), .B(n5008), .ZN(n5010)
         );
  OAI21_X1 U6196 ( .B1(n5011), .B2(n5857), .A(n5010), .ZN(U2825) );
  AOI21_X1 U6197 ( .B1(n5865), .B2(EBX_REG_1__SCAN_IN), .A(n5012), .ZN(n5015)
         );
  NAND2_X1 U6198 ( .A1(n5013), .A2(n5866), .ZN(n5014) );
  OAI211_X1 U6199 ( .C1(n5016), .C2(n6580), .A(n5015), .B(n5014), .ZN(n5018)
         );
  MUX2_X1 U6200 ( .A(n5813), .B(n5870), .S(PHYADDRPOINTER_REG_1__SCAN_IN), .Z(
        n5017) );
  AOI211_X1 U6201 ( .C1(n4344), .C2(n5850), .A(n5018), .B(n5017), .ZN(n5019)
         );
  OAI21_X1 U6202 ( .B1(n5020), .B2(n5857), .A(n5019), .ZN(U2826) );
  INV_X1 U6203 ( .A(n5022), .ZN(n5023) );
  NOR2_X1 U6204 ( .A1(n5024), .A2(n5023), .ZN(n5025) );
  XNOR2_X1 U6205 ( .A(n5021), .B(n5025), .ZN(n5977) );
  AOI22_X1 U6206 ( .A1(n5963), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .B1(n6032), 
        .B2(REIP_REG_12__SCAN_IN), .ZN(n5026) );
  OAI21_X1 U6207 ( .B1(n5973), .B2(n5027), .A(n5026), .ZN(n5028) );
  AOI21_X1 U6208 ( .B1(n5814), .B2(n5515), .A(n5028), .ZN(n5029) );
  OAI21_X1 U6209 ( .B1(n5977), .B2(n5770), .A(n5029), .ZN(U2974) );
  INV_X1 U6210 ( .A(n5973), .ZN(n5538) );
  OAI22_X1 U6211 ( .A1(n5535), .A2(n6534), .B1(n6047), .B2(n6427), .ZN(n5031)
         );
  NOR2_X1 U6212 ( .A1(n5827), .A2(n5542), .ZN(n5030) );
  AOI211_X1 U6213 ( .C1(n5538), .C2(n5824), .A(n5031), .B(n5030), .ZN(n5032)
         );
  OAI21_X1 U6214 ( .B1(n5033), .B2(n5770), .A(n5032), .ZN(U2976) );
  AND2_X1 U6215 ( .A1(n5035), .A2(n5034), .ZN(n5036) );
  OR2_X1 U6216 ( .A1(n5050), .A2(n5036), .ZN(n5081) );
  AOI22_X1 U6217 ( .A1(n5060), .A2(DATAI_13_), .B1(n5884), .B2(
        EAX_REG_13__SCAN_IN), .ZN(n5037) );
  OAI21_X1 U6218 ( .B1(n5081), .B2(n5718), .A(n5037), .ZN(U2878) );
  INV_X1 U6219 ( .A(n5071), .ZN(n5038) );
  AOI21_X1 U6220 ( .B1(n5040), .B2(n5039), .A(n5038), .ZN(n5751) );
  AOI22_X1 U6221 ( .A1(n5751), .A2(n5415), .B1(n5414), .B2(EBX_REG_13__SCAN_IN), .ZN(n5041) );
  OAI21_X1 U6222 ( .B1(n5081), .B2(n5417), .A(n5041), .ZN(U2846) );
  INV_X1 U6223 ( .A(REIP_REG_13__SCAN_IN), .ZN(n6433) );
  INV_X1 U6224 ( .A(REIP_REG_12__SCAN_IN), .ZN(n6431) );
  NOR2_X1 U6225 ( .A1(n6433), .A2(n6431), .ZN(n5796) );
  AOI21_X1 U6226 ( .B1(n6433), .B2(n6431), .A(n5796), .ZN(n5047) );
  AOI21_X1 U6227 ( .B1(n5870), .B2(PHYADDRPOINTER_REG_13__SCAN_IN), .A(n5845), 
        .ZN(n5042) );
  OAI21_X1 U6228 ( .B1(n5868), .B2(n5077), .A(n5042), .ZN(n5046) );
  NAND2_X1 U6229 ( .A1(n5330), .A2(n5043), .ZN(n5809) );
  AOI22_X1 U6230 ( .A1(EBX_REG_13__SCAN_IN), .A2(n5865), .B1(n5866), .B2(n5751), .ZN(n5044) );
  OAI21_X1 U6231 ( .B1(n6433), .B2(n5809), .A(n5044), .ZN(n5045) );
  AOI211_X1 U6232 ( .C1(n5807), .C2(n5047), .A(n5046), .B(n5045), .ZN(n5048)
         );
  OAI21_X1 U6233 ( .B1(n5081), .B2(n5826), .A(n5048), .ZN(U2814) );
  INV_X1 U6234 ( .A(n5049), .ZN(n5053) );
  INV_X1 U6235 ( .A(n5050), .ZN(n5052) );
  INV_X1 U6236 ( .A(n5051), .ZN(n5057) );
  AOI21_X1 U6237 ( .B1(n5053), .B2(n5052), .A(n5057), .ZN(n5802) );
  INV_X1 U6238 ( .A(n5802), .ZN(n5074) );
  AOI22_X1 U6239 ( .A1(n5060), .A2(DATAI_14_), .B1(n5884), .B2(
        EAX_REG_14__SCAN_IN), .ZN(n5054) );
  OAI21_X1 U6240 ( .B1(n5074), .B2(n5718), .A(n5054), .ZN(U2877) );
  INV_X1 U6241 ( .A(n5055), .ZN(n5056) );
  OAI21_X1 U6242 ( .B1(n5057), .B2(n5056), .A(n5111), .ZN(n5145) );
  AOI21_X1 U6243 ( .B1(n5058), .B2(n5073), .A(n5118), .ZN(n5744) );
  AOI22_X1 U6244 ( .A1(n5744), .A2(n5415), .B1(n5414), .B2(EBX_REG_15__SCAN_IN), .ZN(n5059) );
  OAI21_X1 U6245 ( .B1(n5145), .B2(n5417), .A(n5059), .ZN(U2844) );
  AOI22_X1 U6246 ( .A1(n5060), .A2(DATAI_15_), .B1(n5884), .B2(
        EAX_REG_15__SCAN_IN), .ZN(n5061) );
  OAI21_X1 U6247 ( .B1(n5145), .B2(n5718), .A(n5061), .ZN(U2876) );
  NOR2_X1 U6248 ( .A1(REIP_REG_15__SCAN_IN), .A2(n5062), .ZN(n5113) );
  INV_X1 U6249 ( .A(EBX_REG_15__SCAN_IN), .ZN(n5064) );
  AOI22_X1 U6250 ( .A1(PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n5870), .B1(n5866), 
        .B2(n5744), .ZN(n5063) );
  OAI21_X1 U6251 ( .B1(n5064), .B2(n5662), .A(n5063), .ZN(n5065) );
  NOR3_X1 U6252 ( .A1(n5845), .A2(n5113), .A3(n5065), .ZN(n5069) );
  NOR2_X1 U6253 ( .A1(n5853), .A2(n5066), .ZN(n5797) );
  INV_X1 U6254 ( .A(n5141), .ZN(n5067) );
  AOI22_X1 U6255 ( .A1(n5797), .A2(REIP_REG_15__SCAN_IN), .B1(n5067), .B2(
        n5813), .ZN(n5068) );
  OAI211_X1 U6256 ( .C1(n5145), .C2(n5826), .A(n5069), .B(n5068), .ZN(U2812)
         );
  NAND2_X1 U6257 ( .A1(n5071), .A2(n5070), .ZN(n5072) );
  NAND2_X1 U6258 ( .A1(n5073), .A2(n5072), .ZN(n5798) );
  INV_X1 U6259 ( .A(EBX_REG_14__SCAN_IN), .ZN(n6550) );
  OAI222_X1 U6260 ( .A1(n5798), .A2(n5428), .B1(n5427), .B2(n6550), .C1(n5417), 
        .C2(n5074), .ZN(U2845) );
  XNOR2_X1 U6261 ( .A(n5076), .B(n5075), .ZN(n5753) );
  NAND2_X1 U6262 ( .A1(n5753), .A2(n5968), .ZN(n5080) );
  NOR2_X1 U6263 ( .A1(n6047), .A2(n6433), .ZN(n5750) );
  NOR2_X1 U6264 ( .A1(n5973), .A2(n5077), .ZN(n5078) );
  AOI211_X1 U6265 ( .C1(n5963), .C2(PHYADDRPOINTER_REG_13__SCAN_IN), .A(n5750), 
        .B(n5078), .ZN(n5079) );
  OAI211_X1 U6266 ( .C1(n5542), .C2(n5081), .A(n5080), .B(n5079), .ZN(U2973)
         );
  XNOR2_X1 U6267 ( .A(n3422), .B(n5083), .ZN(n5084) );
  XNOR2_X1 U6268 ( .A(n5082), .B(n5084), .ZN(n5109) );
  INV_X1 U6269 ( .A(n5085), .ZN(n5094) );
  AOI21_X1 U6270 ( .B1(n5087), .B2(n6040), .A(n5086), .ZN(n5088) );
  INV_X1 U6271 ( .A(n5088), .ZN(n5089) );
  AOI21_X1 U6272 ( .B1(n5600), .B2(n5090), .A(n5089), .ZN(n5989) );
  OAI21_X1 U6273 ( .B1(n5092), .B2(n5091), .A(n5989), .ZN(n5093) );
  AOI21_X1 U6274 ( .B1(n5094), .B2(n5099), .A(n5093), .ZN(n5756) );
  OAI21_X1 U6275 ( .B1(n5096), .B2(n5095), .A(n3404), .ZN(n5097) );
  AOI21_X1 U6276 ( .B1(n5756), .B2(n5097), .A(n5083), .ZN(n5103) );
  NOR2_X1 U6277 ( .A1(n5798), .A2(n6024), .ZN(n5102) );
  INV_X1 U6278 ( .A(REIP_REG_14__SCAN_IN), .ZN(n5098) );
  NOR2_X1 U6279 ( .A1(n6047), .A2(n5098), .ZN(n5106) );
  INV_X1 U6280 ( .A(n5984), .ZN(n5100) );
  NOR3_X1 U6281 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n5100), .A3(n5099), 
        .ZN(n5101) );
  NOR4_X1 U6282 ( .A1(n5103), .A2(n5102), .A3(n5106), .A4(n5101), .ZN(n5104)
         );
  OAI21_X1 U6283 ( .B1(n5109), .B2(n6023), .A(n5104), .ZN(U3004) );
  AND2_X1 U6284 ( .A1(n5963), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n5105)
         );
  AOI211_X1 U6285 ( .C1(n5538), .C2(n5801), .A(n5106), .B(n5105), .ZN(n5108)
         );
  NAND2_X1 U6286 ( .A1(n5802), .A2(n5515), .ZN(n5107) );
  OAI211_X1 U6287 ( .C1(n5109), .C2(n5770), .A(n5108), .B(n5107), .ZN(U2972)
         );
  INV_X1 U6288 ( .A(n5128), .ZN(n5110) );
  AOI21_X1 U6289 ( .B1(n5112), .B2(n5111), .A(n5110), .ZN(n5883) );
  INV_X1 U6290 ( .A(n5883), .ZN(n5125) );
  INV_X1 U6291 ( .A(n5342), .ZN(n5115) );
  NOR2_X1 U6292 ( .A1(n5797), .A2(n5113), .ZN(n5114) );
  MUX2_X1 U6293 ( .A(n5115), .B(n5114), .S(REIP_REG_16__SCAN_IN), .Z(n5124) );
  OR2_X1 U6294 ( .A1(n5118), .A2(n5117), .ZN(n5119) );
  NAND2_X1 U6295 ( .A1(n5133), .A2(n5119), .ZN(n5160) );
  AOI22_X1 U6296 ( .A1(EBX_REG_16__SCAN_IN), .A2(n5865), .B1(n5120), .B2(n5813), .ZN(n5121) );
  OAI21_X1 U6297 ( .B1(n5863), .B2(n5160), .A(n5121), .ZN(n5122) );
  AOI211_X1 U6298 ( .C1(n5870), .C2(PHYADDRPOINTER_REG_16__SCAN_IN), .A(n5845), 
        .B(n5122), .ZN(n5123) );
  OAI211_X1 U6299 ( .C1(n5125), .C2(n5826), .A(n5124), .B(n5123), .ZN(U2811)
         );
  INV_X1 U6300 ( .A(EBX_REG_16__SCAN_IN), .ZN(n5126) );
  OAI222_X1 U6301 ( .A1(n5428), .A2(n5160), .B1(n5427), .B2(n5126), .C1(n5125), 
        .C2(n5417), .ZN(U2843) );
  AND2_X1 U6302 ( .A1(n5128), .A2(n5127), .ZN(n5130) );
  OR2_X1 U6303 ( .A1(n5130), .A2(n5423), .ZN(n5541) );
  NAND2_X1 U6304 ( .A1(n5133), .A2(n5132), .ZN(n5134) );
  AND2_X1 U6305 ( .A1(n5419), .A2(n5134), .ZN(n5737) );
  INV_X1 U6306 ( .A(EBX_REG_17__SCAN_IN), .ZN(n5135) );
  NOR2_X1 U6307 ( .A1(n5427), .A2(n5135), .ZN(n5136) );
  AOI21_X1 U6308 ( .B1(n5737), .B2(n5415), .A(n5136), .ZN(n5137) );
  OAI21_X1 U6309 ( .B1(n5541), .B2(n5417), .A(n5137), .ZN(U2842) );
  XNOR2_X1 U6310 ( .A(n3422), .B(n5162), .ZN(n5139) );
  XNOR2_X1 U6311 ( .A(n5140), .B(n5139), .ZN(n5746) );
  NAND2_X1 U6312 ( .A1(n5746), .A2(n5968), .ZN(n5144) );
  AND2_X1 U6313 ( .A1(n6032), .A2(REIP_REG_15__SCAN_IN), .ZN(n5743) );
  NOR2_X1 U6314 ( .A1(n5973), .A2(n5141), .ZN(n5142) );
  AOI211_X1 U6315 ( .C1(n5963), .C2(PHYADDRPOINTER_REG_15__SCAN_IN), .A(n5743), 
        .B(n5142), .ZN(n5143) );
  OAI211_X1 U6316 ( .C1(n5542), .C2(n5145), .A(n5144), .B(n5143), .ZN(U2971)
         );
  OAI222_X1 U6317 ( .A1(n5417), .A2(n5276), .B1(n5428), .B2(n5216), .C1(n5146), 
        .C2(n5427), .ZN(U2829) );
  INV_X1 U6318 ( .A(n5637), .ZN(n6472) );
  NOR2_X1 U6319 ( .A1(n5771), .A2(n6468), .ZN(n5147) );
  AOI21_X1 U6320 ( .B1(n6349), .B2(n6383), .A(n5147), .ZN(n5757) );
  NAND2_X1 U6321 ( .A1(n5757), .A2(n5148), .ZN(n6477) );
  INV_X1 U6322 ( .A(n6477), .ZN(n5154) );
  AOI21_X1 U6323 ( .B1(n6472), .B2(n5150), .A(n5154), .ZN(n5157) );
  AOI22_X1 U6324 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B1(n6623), .B2(n5149), .ZN(n5283)
         );
  NAND2_X1 U6325 ( .A1(STATE2_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n5282) );
  INV_X1 U6326 ( .A(n5282), .ZN(n6475) );
  NOR3_X1 U6327 ( .A1(n5637), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n5150), 
        .ZN(n5153) );
  INV_X1 U6328 ( .A(n5151), .ZN(n6343) );
  INV_X1 U6329 ( .A(n6384), .ZN(n6479) );
  NOR2_X1 U6330 ( .A1(n6343), .A2(n6479), .ZN(n5152) );
  AOI211_X1 U6331 ( .C1(n5283), .C2(n6475), .A(n5153), .B(n5152), .ZN(n5155)
         );
  OAI22_X1 U6332 ( .A1(n5157), .A2(n5156), .B1(n5155), .B2(n5154), .ZN(U3459)
         );
  XNOR2_X1 U6333 ( .A(n3422), .B(n5161), .ZN(n5158) );
  XNOR2_X1 U6334 ( .A(n5529), .B(n5158), .ZN(n5171) );
  OAI21_X1 U6335 ( .B1(n5159), .B2(n5601), .A(n5989), .ZN(n5745) );
  NOR2_X1 U6336 ( .A1(n5160), .A2(n6024), .ZN(n5165) );
  INV_X1 U6337 ( .A(REIP_REG_16__SCAN_IN), .ZN(n6438) );
  OAI221_X1 U6338 ( .B1(INSTADDRPOINTER_REG_15__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .C1(n5162), .C2(n5161), .A(n5742), 
        .ZN(n5163) );
  OAI21_X1 U6339 ( .B1(n6047), .B2(n6438), .A(n5163), .ZN(n5164) );
  AOI211_X1 U6340 ( .C1(n5745), .C2(INSTADDRPOINTER_REG_16__SCAN_IN), .A(n5165), .B(n5164), .ZN(n5166) );
  OAI21_X1 U6341 ( .B1(n5171), .B2(n6023), .A(n5166), .ZN(U3002) );
  AOI22_X1 U6342 ( .A1(n5963), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .B1(n6032), 
        .B2(REIP_REG_16__SCAN_IN), .ZN(n5167) );
  OAI21_X1 U6343 ( .B1(n5973), .B2(n5168), .A(n5167), .ZN(n5169) );
  AOI21_X1 U6344 ( .B1(n5883), .B2(n5515), .A(n5169), .ZN(n5170) );
  OAI21_X1 U6345 ( .B1(n5171), .B2(n5770), .A(n5170), .ZN(U2970) );
  INV_X1 U6346 ( .A(n5172), .ZN(n5181) );
  OR2_X1 U6347 ( .A1(n5362), .A2(n5173), .ZN(n5175) );
  INV_X1 U6348 ( .A(n5643), .ZN(n5178) );
  AOI21_X1 U6349 ( .B1(n5963), .B2(PHYADDRPOINTER_REG_29__SCAN_IN), .A(n5176), 
        .ZN(n5177) );
  OAI21_X1 U6350 ( .B1(n5973), .B2(n5178), .A(n5177), .ZN(n5179) );
  AOI21_X1 U6351 ( .B1(n5646), .B2(n5515), .A(n5179), .ZN(n5180) );
  OAI21_X1 U6352 ( .B1(n5181), .B2(n5770), .A(n5180), .ZN(U2957) );
  INV_X1 U6353 ( .A(n5182), .ZN(n5183) );
  AND2_X1 U6354 ( .A1(n5466), .A2(n5183), .ZN(n5184) );
  OR2_X1 U6355 ( .A1(n5185), .A2(n5184), .ZN(n5186) );
  XNOR2_X1 U6356 ( .A(n5186), .B(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5226)
         );
  INV_X1 U6357 ( .A(REIP_REG_30__SCAN_IN), .ZN(n5187) );
  NOR2_X1 U6358 ( .A1(n6047), .A2(n5187), .ZN(n5217) );
  AOI21_X1 U6359 ( .B1(n5963), .B2(PHYADDRPOINTER_REG_30__SCAN_IN), .A(n5217), 
        .ZN(n5188) );
  OAI21_X1 U6360 ( .B1(n5973), .B2(n5189), .A(n5188), .ZN(n5190) );
  AOI21_X1 U6361 ( .B1(n5191), .B2(n5515), .A(n5190), .ZN(n5192) );
  OAI21_X1 U6362 ( .B1(n5226), .B2(n5770), .A(n5192), .ZN(U2956) );
  AOI21_X1 U6363 ( .B1(n5195), .B2(n5194), .A(n5193), .ZN(n5222) );
  OAI21_X1 U6364 ( .B1(INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n5601), .A(n5222), 
        .ZN(n5198) );
  AND4_X1 U6365 ( .A1(n5218), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_30__SCAN_IN), .A4(n6623), .ZN(n5196) );
  AOI211_X1 U6366 ( .C1(n5198), .C2(INSTADDRPOINTER_REG_31__SCAN_IN), .A(n5197), .B(n5196), .ZN(n5200) );
  NAND2_X1 U6367 ( .A1(n5356), .A2(n6044), .ZN(n5199) );
  OAI211_X1 U6368 ( .C1(n5201), .C2(n6023), .A(n5200), .B(n5199), .ZN(U2987)
         );
  OR2_X1 U6369 ( .A1(n5376), .A2(n5202), .ZN(n5203) );
  NAND2_X1 U6370 ( .A1(n5364), .A2(n5203), .ZN(n5369) );
  NOR2_X1 U6371 ( .A1(n5205), .A2(n5204), .ZN(n5206) );
  INV_X1 U6372 ( .A(n5206), .ZN(n5617) );
  NAND2_X1 U6373 ( .A1(n5617), .A2(n5207), .ZN(n5473) );
  INV_X1 U6374 ( .A(n5473), .ZN(n5211) );
  NAND2_X1 U6375 ( .A1(n5209), .A2(n5208), .ZN(n5555) );
  INV_X1 U6376 ( .A(n5555), .ZN(n5210) );
  NOR2_X1 U6377 ( .A1(n5457), .A2(n5456), .ZN(n5212) );
  XNOR2_X1 U6378 ( .A(n5212), .B(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5232)
         );
  NAND2_X1 U6379 ( .A1(n5232), .A2(n6050), .ZN(n5215) );
  NOR2_X1 U6380 ( .A1(n6047), .A2(n6620), .ZN(n5234) );
  NOR2_X1 U6381 ( .A1(n5549), .A2(n5455), .ZN(n5213) );
  AOI211_X1 U6382 ( .C1(n5546), .C2(n5455), .A(n5234), .B(n5213), .ZN(n5214)
         );
  OAI211_X1 U6383 ( .C1(n6024), .C2(n5369), .A(n5215), .B(n5214), .ZN(U2991)
         );
  INV_X1 U6384 ( .A(n5216), .ZN(n5224) );
  INV_X1 U6385 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5221) );
  INV_X1 U6386 ( .A(n5217), .ZN(n5220) );
  NAND3_X1 U6387 ( .A1(n5218), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .A3(n5221), .ZN(n5219) );
  OAI211_X1 U6388 ( .C1(n5222), .C2(n5221), .A(n5220), .B(n5219), .ZN(n5223)
         );
  AOI21_X1 U6389 ( .B1(n5224), .B2(n6044), .A(n5223), .ZN(n5225) );
  OAI21_X1 U6390 ( .B1(n5226), .B2(n6023), .A(n5225), .ZN(U2988) );
  CLKBUF_X3 U6391 ( .A(n5326), .Z(n5425) );
  NOR2_X1 U6392 ( .A1(n5373), .A2(n5230), .ZN(n5231) );
  NAND2_X1 U6393 ( .A1(n5232), .A2(n5968), .ZN(n5236) );
  NOR2_X1 U6394 ( .A1(n5535), .A2(n5309), .ZN(n5233) );
  AOI211_X1 U6395 ( .C1(n5538), .C2(n5307), .A(n5234), .B(n5233), .ZN(n5235)
         );
  OAI211_X1 U6396 ( .C1(n5542), .C2(n5443), .A(n5236), .B(n5235), .ZN(U2959)
         );
  NAND2_X1 U6397 ( .A1(n3422), .A2(n5613), .ZN(n5240) );
  INV_X1 U6398 ( .A(n5240), .ZN(n5237) );
  XNOR2_X1 U6399 ( .A(n3422), .B(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5520)
         );
  AND2_X1 U6400 ( .A1(n5481), .A2(n5483), .ZN(n5239) );
  OR2_X1 U6401 ( .A1(n3422), .A2(n5510), .ZN(n5238) );
  AND2_X1 U6402 ( .A1(n5239), .A2(n5238), .ZN(n5241) );
  AND2_X1 U6403 ( .A1(n5517), .A2(n5240), .ZN(n5482) );
  INV_X1 U6404 ( .A(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5242) );
  XNOR2_X1 U6405 ( .A(n3422), .B(n5242), .ZN(n5505) );
  NAND3_X1 U6406 ( .A1(n3422), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5245) );
  NAND2_X1 U6407 ( .A1(n5503), .A2(n5494), .ZN(n5485) );
  INV_X1 U6408 ( .A(n5485), .ZN(n5248) );
  INV_X1 U6409 ( .A(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5247) );
  NAND2_X1 U6410 ( .A1(n5425), .A2(n5252), .ZN(n5254) );
  AOI21_X1 U6411 ( .B1(n5255), .B2(n5254), .A(n5381), .ZN(n5388) );
  AND2_X1 U6412 ( .A1(n6032), .A2(REIP_REG_24__SCAN_IN), .ZN(n5266) );
  AOI21_X1 U6413 ( .B1(n5963), .B2(PHYADDRPOINTER_REG_24__SCAN_IN), .A(n5266), 
        .ZN(n5256) );
  OAI21_X1 U6414 ( .B1(n5973), .B2(n5683), .A(n5256), .ZN(n5257) );
  AOI21_X1 U6415 ( .B1(n5388), .B2(n5515), .A(n5257), .ZN(n5258) );
  OAI21_X1 U6416 ( .B1(n5269), .B2(n5770), .A(n5258), .ZN(U2962) );
  OR2_X1 U6417 ( .A1(n5317), .A2(n5260), .ZN(n5261) );
  NAND2_X1 U6418 ( .A1(n5382), .A2(n5261), .ZN(n5691) );
  INV_X1 U6419 ( .A(n5691), .ZN(n5267) );
  INV_X1 U6420 ( .A(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5264) );
  AOI211_X1 U6421 ( .C1(n5264), .C2(n5572), .A(n5263), .B(n5262), .ZN(n5265)
         );
  AOI211_X1 U6422 ( .C1(n5267), .C2(n6044), .A(n5266), .B(n5265), .ZN(n5268)
         );
  OAI21_X1 U6423 ( .B1(n5269), .B2(n6023), .A(n5268), .ZN(U2994) );
  NOR2_X2 U6424 ( .A1(n5884), .A2(n5270), .ZN(n5881) );
  AOI22_X1 U6425 ( .A1(n5881), .A2(DATAI_30_), .B1(EAX_REG_30__SCAN_IN), .B2(
        n5884), .ZN(n5275) );
  AND2_X1 U6426 ( .A1(n5272), .A2(n5271), .ZN(n5273) );
  NAND2_X1 U6427 ( .A1(n5885), .A2(DATAI_14_), .ZN(n5274) );
  OAI211_X1 U6428 ( .C1(n5276), .C2(n5718), .A(n5275), .B(n5274), .ZN(U2861)
         );
  CLKBUF_X1 U6429 ( .A(n2989), .Z(n5278) );
  INV_X1 U6430 ( .A(n5278), .ZN(n5284) );
  OAI21_X1 U6431 ( .B1(n5278), .B2(n5285), .A(n5277), .ZN(n5279) );
  OAI21_X1 U6432 ( .B1(n5280), .B2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(n5279), 
        .ZN(n5281) );
  AOI21_X1 U6433 ( .B1(n4344), .B2(n6344), .A(n5281), .ZN(n6350) );
  OAI222_X1 U6434 ( .A1(n5637), .A2(n5284), .B1(n5283), .B2(n5282), .C1(n6479), 
        .C2(n6350), .ZN(n5286) );
  AOI22_X1 U6435 ( .A1(n6477), .A2(n5286), .B1(n5285), .B2(n6472), .ZN(n5287)
         );
  OAI21_X1 U6436 ( .B1(n6477), .B2(n5288), .A(n5287), .ZN(U3460) );
  INV_X1 U6437 ( .A(n5289), .ZN(n5290) );
  OR2_X1 U6438 ( .A1(n5302), .A2(n5290), .ZN(n5297) );
  NAND2_X1 U6439 ( .A1(n5292), .A2(n5291), .ZN(n5296) );
  NAND2_X1 U6440 ( .A1(n5293), .A2(n4115), .ZN(n5294) );
  NAND2_X1 U6441 ( .A1(n5302), .A2(n5294), .ZN(n5295) );
  AND3_X1 U6442 ( .A1(n5297), .A2(n5296), .A3(n5295), .ZN(n6364) );
  INV_X1 U6443 ( .A(n6364), .ZN(n5305) );
  INV_X1 U6444 ( .A(n5298), .ZN(n5299) );
  AND2_X1 U6445 ( .A1(n4115), .A2(n5299), .ZN(n5300) );
  AOI21_X1 U6446 ( .B1(n5302), .B2(n5301), .A(n5300), .ZN(n5762) );
  NAND2_X1 U6447 ( .A1(n5303), .A2(n6402), .ZN(n5304) );
  NAND2_X1 U6448 ( .A1(n5304), .A2(n6492), .ZN(n6494) );
  AND2_X1 U6449 ( .A1(n5762), .A2(n6494), .ZN(n6360) );
  NOR2_X1 U6450 ( .A1(n6360), .A2(n6369), .ZN(n5772) );
  MUX2_X1 U6451 ( .A(MORE_REG_SCAN_IN), .B(n5305), .S(n5772), .Z(U3471) );
  INV_X1 U6452 ( .A(n5443), .ZN(n5306) );
  NAND2_X1 U6453 ( .A1(n5306), .A2(n5838), .ZN(n5312) );
  INV_X1 U6454 ( .A(REIP_REG_27__SCAN_IN), .ZN(n6620) );
  AOI22_X1 U6455 ( .A1(EBX_REG_27__SCAN_IN), .A2(n5865), .B1(n5307), .B2(n5813), .ZN(n5308) );
  OAI21_X1 U6456 ( .B1(n5309), .B2(n5834), .A(n5308), .ZN(n5310) );
  AOI221_X1 U6457 ( .B1(n5667), .B2(REIP_REG_27__SCAN_IN), .C1(n5657), .C2(
        n6620), .A(n5310), .ZN(n5311) );
  OAI211_X1 U6458 ( .C1(n5863), .C2(n5369), .A(n5312), .B(n5311), .ZN(U2800)
         );
  XOR2_X1 U6459 ( .A(n5314), .B(n5393), .Z(n5492) );
  INV_X1 U6460 ( .A(n5492), .ZN(n5452) );
  NAND2_X1 U6461 ( .A1(n6446), .A2(n5315), .ZN(n5324) );
  AND2_X1 U6462 ( .A1(n5330), .A2(n5316), .ZN(n5685) );
  AOI21_X1 U6463 ( .B1(n5318), .B2(n5395), .A(n5317), .ZN(n5574) );
  INV_X1 U6464 ( .A(n5574), .ZN(n5322) );
  INV_X1 U6465 ( .A(EBX_REG_23__SCAN_IN), .ZN(n5319) );
  OAI22_X1 U6466 ( .A1(n5319), .A2(n5662), .B1(n5490), .B2(n5834), .ZN(n5320)
         );
  AOI21_X1 U6467 ( .B1(n5813), .B2(n5488), .A(n5320), .ZN(n5321) );
  OAI21_X1 U6468 ( .B1(n5322), .B2(n5863), .A(n5321), .ZN(n5323) );
  AOI21_X1 U6469 ( .B1(n5324), .B2(n5685), .A(n5323), .ZN(n5325) );
  OAI21_X1 U6470 ( .B1(n5452), .B2(n5826), .A(n5325), .ZN(U2804) );
  NAND2_X1 U6471 ( .A1(n5326), .A2(n5327), .ZN(n5407) );
  OAI21_X1 U6472 ( .B1(n5425), .B2(n5327), .A(n5407), .ZN(n5728) );
  INV_X1 U6473 ( .A(n5328), .ZN(n5333) );
  AND2_X1 U6474 ( .A1(n5330), .A2(n5329), .ZN(n5788) );
  NOR2_X1 U6475 ( .A1(REIP_REG_18__SCAN_IN), .A2(n5331), .ZN(n5793) );
  NOR2_X1 U6476 ( .A1(n5788), .A2(n5793), .ZN(n5332) );
  MUX2_X1 U6477 ( .A(n5333), .B(n5332), .S(REIP_REG_19__SCAN_IN), .Z(n5341) );
  AND2_X1 U6478 ( .A1(n5335), .A2(n5334), .ZN(n5418) );
  NOR2_X1 U6479 ( .A1(n5419), .A2(n5418), .ZN(n5420) );
  XNOR2_X1 U6480 ( .A(n5420), .B(n5336), .ZN(n5610) );
  AOI22_X1 U6481 ( .A1(n5524), .A2(n5813), .B1(n5866), .B2(n5610), .ZN(n5337)
         );
  OAI21_X1 U6482 ( .B1(n5338), .B2(n5662), .A(n5337), .ZN(n5339) );
  AOI211_X1 U6483 ( .C1(n5870), .C2(PHYADDRPOINTER_REG_19__SCAN_IN), .A(n5845), 
        .B(n5339), .ZN(n5340) );
  OAI211_X1 U6484 ( .C1(n5728), .C2(n5826), .A(n5341), .B(n5340), .ZN(U2808)
         );
  OAI221_X1 U6485 ( .B1(REIP_REG_17__SCAN_IN), .B2(n5342), .C1(
        REIP_REG_17__SCAN_IN), .C2(REIP_REG_16__SCAN_IN), .A(n5788), .ZN(n5346) );
  AOI22_X1 U6486 ( .A1(EBX_REG_17__SCAN_IN), .A2(n5865), .B1(n5537), .B2(n5813), .ZN(n5343) );
  OAI21_X1 U6487 ( .B1(n5534), .B2(n5834), .A(n5343), .ZN(n5344) );
  AOI211_X1 U6488 ( .C1(n5737), .C2(n5866), .A(n5845), .B(n5344), .ZN(n5345)
         );
  OAI211_X1 U6489 ( .C1(n5541), .C2(n5826), .A(n5346), .B(n5345), .ZN(U2810)
         );
  INV_X1 U6490 ( .A(n5809), .ZN(n5353) );
  NAND2_X1 U6491 ( .A1(REIP_REG_10__SCAN_IN), .A2(REIP_REG_9__SCAN_IN), .ZN(
        n5819) );
  OAI21_X1 U6492 ( .B1(n5818), .B2(n5819), .A(n4967), .ZN(n5352) );
  AOI22_X1 U6493 ( .A1(EBX_REG_11__SCAN_IN), .A2(n5865), .B1(
        PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n5870), .ZN(n5350) );
  OAI21_X1 U6494 ( .B1(n5868), .B2(n5347), .A(n5854), .ZN(n5348) );
  AOI21_X1 U6495 ( .B1(n5983), .B2(n5866), .A(n5348), .ZN(n5349) );
  NAND2_X1 U6496 ( .A1(n5350), .A2(n5349), .ZN(n5351) );
  AOI21_X1 U6497 ( .B1(n5353), .B2(n5352), .A(n5351), .ZN(n5354) );
  OAI21_X1 U6498 ( .B1(n5355), .B2(n5826), .A(n5354), .ZN(U2816) );
  INV_X1 U6499 ( .A(n5356), .ZN(n5358) );
  OAI22_X1 U6500 ( .A1(n5358), .A2(n5428), .B1(n5357), .B2(n5427), .ZN(U2828)
         );
  OAI222_X1 U6501 ( .A1(n5417), .A2(n5438), .B1(n5427), .B2(n5359), .C1(n5644), 
        .C2(n5428), .ZN(U2830) );
  NOR2_X1 U6502 ( .A1(n5228), .A2(n5360), .ZN(n5361) );
  OR2_X1 U6503 ( .A1(n5362), .A2(n5361), .ZN(n5459) );
  NAND2_X1 U6504 ( .A1(n5364), .A2(n5363), .ZN(n5365) );
  NAND2_X1 U6505 ( .A1(n5366), .A2(n5365), .ZN(n5660) );
  OAI22_X1 U6506 ( .A1(n5660), .A2(n5428), .B1(n6607), .B2(n5427), .ZN(n5367)
         );
  INV_X1 U6507 ( .A(n5367), .ZN(n5368) );
  OAI21_X1 U6508 ( .B1(n5459), .B2(n5417), .A(n5368), .ZN(U2831) );
  OAI222_X1 U6509 ( .A1(n5417), .A2(n5443), .B1(n5427), .B2(n5370), .C1(n5369), 
        .C2(n5428), .ZN(U2832) );
  NAND2_X1 U6510 ( .A1(n5425), .A2(n5371), .ZN(n5379) );
  AND2_X1 U6511 ( .A1(n5384), .A2(n5374), .ZN(n5375) );
  OR2_X1 U6512 ( .A1(n5376), .A2(n5375), .ZN(n5671) );
  OAI22_X1 U6513 ( .A1(n5671), .A2(n5428), .B1(n5663), .B2(n5427), .ZN(n5377)
         );
  INV_X1 U6514 ( .A(n5377), .ZN(n5378) );
  OAI21_X1 U6515 ( .B1(n5467), .B2(n5417), .A(n5378), .ZN(U2833) );
  INV_X1 U6516 ( .A(EBX_REG_25__SCAN_IN), .ZN(n5387) );
  INV_X1 U6517 ( .A(n5382), .ZN(n5386) );
  INV_X1 U6518 ( .A(n5383), .ZN(n5385) );
  OAI21_X1 U6519 ( .B1(n5386), .B2(n5385), .A(n5384), .ZN(n5674) );
  OAI222_X1 U6520 ( .A1(n5417), .A2(n5673), .B1(n5427), .B2(n5387), .C1(n5674), 
        .C2(n5428), .ZN(U2834) );
  INV_X1 U6521 ( .A(n5388), .ZN(n5687) );
  INV_X1 U6522 ( .A(EBX_REG_24__SCAN_IN), .ZN(n6622) );
  OAI222_X1 U6523 ( .A1(n5417), .A2(n5687), .B1(n5427), .B2(n6622), .C1(n5691), 
        .C2(n5428), .ZN(U2835) );
  AOI22_X1 U6524 ( .A1(n5574), .A2(n5415), .B1(n5414), .B2(EBX_REG_23__SCAN_IN), .ZN(n5389) );
  OAI21_X1 U6525 ( .B1(n5452), .B2(n5417), .A(n5389), .ZN(U2836) );
  NOR2_X1 U6526 ( .A1(n5400), .A2(n5391), .ZN(n5392) );
  INV_X1 U6527 ( .A(n5395), .ZN(n5396) );
  AOI21_X1 U6528 ( .B1(n5397), .B2(n5394), .A(n5396), .ZN(n5694) );
  AOI22_X1 U6529 ( .A1(n5694), .A2(n5415), .B1(EBX_REG_22__SCAN_IN), .B2(n5414), .ZN(n5398) );
  OAI21_X1 U6530 ( .B1(n5497), .B2(n5417), .A(n5398), .ZN(U2837) );
  AND2_X1 U6531 ( .A1(n5405), .A2(n5399), .ZN(n5401) );
  OAI21_X1 U6532 ( .B1(n5403), .B2(n5402), .A(n5394), .ZN(n5706) );
  OAI222_X1 U6533 ( .A1(n5417), .A2(n5705), .B1(n5427), .B2(n5404), .C1(n5706), 
        .C2(n5428), .ZN(U2838) );
  INV_X1 U6534 ( .A(n5405), .ZN(n5406) );
  AOI21_X1 U6535 ( .B1(n5408), .B2(n5407), .A(n5406), .ZN(n5725) );
  INV_X1 U6536 ( .A(n5725), .ZN(n5413) );
  MUX2_X1 U6537 ( .A(n4110), .B(n5409), .S(n2968), .Z(n5411) );
  XNOR2_X1 U6538 ( .A(n5411), .B(n5410), .ZN(n5717) );
  INV_X1 U6539 ( .A(EBX_REG_20__SCAN_IN), .ZN(n5412) );
  OAI222_X1 U6540 ( .A1(n5417), .A2(n5413), .B1(n5428), .B2(n5717), .C1(n5412), 
        .C2(n5427), .ZN(U2839) );
  AOI22_X1 U6541 ( .A1(n5610), .A2(n5415), .B1(n5414), .B2(EBX_REG_19__SCAN_IN), .ZN(n5416) );
  OAI21_X1 U6542 ( .B1(n5728), .B2(n5417), .A(n5416), .ZN(U2840) );
  AND2_X1 U6543 ( .A1(n5419), .A2(n5418), .ZN(n5421) );
  OR2_X1 U6544 ( .A1(n5421), .A2(n5420), .ZN(n5795) );
  INV_X1 U6545 ( .A(EBX_REG_18__SCAN_IN), .ZN(n5426) );
  NOR2_X1 U6546 ( .A1(n5423), .A2(n5422), .ZN(n5424) );
  OR2_X1 U6547 ( .A1(n5425), .A2(n5424), .ZN(n5732) );
  OAI222_X1 U6548 ( .A1(n5428), .A2(n5795), .B1(n5427), .B2(n5426), .C1(n5417), 
        .C2(n5732), .ZN(U2841) );
  AND2_X1 U6549 ( .A1(n5435), .A2(n5429), .ZN(n5430) );
  NAND2_X1 U6550 ( .A1(n5431), .A2(n5430), .ZN(n5433) );
  NAND2_X1 U6551 ( .A1(n5881), .A2(DATAI_31_), .ZN(n5432) );
  OAI211_X1 U6552 ( .C1(n5435), .C2(n5434), .A(n5433), .B(n5432), .ZN(U2860)
         );
  AOI22_X1 U6553 ( .A1(n5885), .A2(DATAI_13_), .B1(n5884), .B2(
        EAX_REG_29__SCAN_IN), .ZN(n5437) );
  NAND2_X1 U6554 ( .A1(n5881), .A2(DATAI_29_), .ZN(n5436) );
  OAI211_X1 U6555 ( .C1(n5438), .C2(n5718), .A(n5437), .B(n5436), .ZN(U2862)
         );
  AOI22_X1 U6556 ( .A1(n5885), .A2(DATAI_12_), .B1(n5884), .B2(
        EAX_REG_28__SCAN_IN), .ZN(n5440) );
  NAND2_X1 U6557 ( .A1(n5881), .A2(DATAI_28_), .ZN(n5439) );
  OAI211_X1 U6558 ( .C1(n5459), .C2(n5718), .A(n5440), .B(n5439), .ZN(U2863)
         );
  AOI22_X1 U6559 ( .A1(n5881), .A2(DATAI_27_), .B1(EAX_REG_27__SCAN_IN), .B2(
        n5884), .ZN(n5442) );
  NAND2_X1 U6560 ( .A1(n5885), .A2(DATAI_11_), .ZN(n5441) );
  OAI211_X1 U6561 ( .C1(n5443), .C2(n5718), .A(n5442), .B(n5441), .ZN(U2864)
         );
  AOI22_X1 U6562 ( .A1(n5885), .A2(DATAI_10_), .B1(n5884), .B2(
        EAX_REG_26__SCAN_IN), .ZN(n5445) );
  NAND2_X1 U6563 ( .A1(n5881), .A2(DATAI_26_), .ZN(n5444) );
  OAI211_X1 U6564 ( .C1(n5467), .C2(n5718), .A(n5445), .B(n5444), .ZN(U2865)
         );
  AOI22_X1 U6565 ( .A1(n5885), .A2(DATAI_9_), .B1(n5884), .B2(
        EAX_REG_25__SCAN_IN), .ZN(n5447) );
  NAND2_X1 U6566 ( .A1(n5881), .A2(DATAI_25_), .ZN(n5446) );
  OAI211_X1 U6567 ( .C1(n5673), .C2(n5718), .A(n5447), .B(n5446), .ZN(U2866)
         );
  AOI22_X1 U6568 ( .A1(n5885), .A2(DATAI_8_), .B1(n5884), .B2(
        EAX_REG_24__SCAN_IN), .ZN(n5449) );
  NAND2_X1 U6569 ( .A1(n5881), .A2(DATAI_24_), .ZN(n5448) );
  OAI211_X1 U6570 ( .C1(n5687), .C2(n5718), .A(n5449), .B(n5448), .ZN(U2867)
         );
  AOI22_X1 U6571 ( .A1(n5881), .A2(DATAI_23_), .B1(EAX_REG_23__SCAN_IN), .B2(
        n5884), .ZN(n5451) );
  NAND2_X1 U6572 ( .A1(n5885), .A2(DATAI_7_), .ZN(n5450) );
  OAI211_X1 U6573 ( .C1(n5452), .C2(n5718), .A(n5451), .B(n5450), .ZN(U2868)
         );
  AOI22_X1 U6574 ( .A1(n5881), .A2(DATAI_17_), .B1(EAX_REG_17__SCAN_IN), .B2(
        n5884), .ZN(n5454) );
  NAND2_X1 U6575 ( .A1(n5885), .A2(DATAI_1_), .ZN(n5453) );
  OAI211_X1 U6576 ( .C1(n5541), .C2(n5718), .A(n5454), .B(n5453), .ZN(U2874)
         );
  AOI22_X1 U6577 ( .A1(n5457), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .B1(n5456), .B2(n5455), .ZN(n5458) );
  XNOR2_X1 U6578 ( .A(n5458), .B(n6586), .ZN(n5553) );
  INV_X1 U6579 ( .A(n5459), .ZN(n5656) );
  INV_X1 U6580 ( .A(REIP_REG_28__SCAN_IN), .ZN(n5460) );
  OR2_X1 U6581 ( .A1(n6047), .A2(n5460), .ZN(n5548) );
  INV_X1 U6582 ( .A(n5548), .ZN(n5461) );
  AOI21_X1 U6583 ( .B1(n5963), .B2(PHYADDRPOINTER_REG_28__SCAN_IN), .A(n5461), 
        .ZN(n5462) );
  OAI21_X1 U6584 ( .B1(n5973), .B2(n5650), .A(n5462), .ZN(n5463) );
  AOI21_X1 U6585 ( .B1(n5656), .B2(n5515), .A(n5463), .ZN(n5464) );
  OAI21_X1 U6586 ( .B1(n5553), .B2(n5770), .A(n5464), .ZN(U2958) );
  XNOR2_X1 U6587 ( .A(n3422), .B(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5465)
         );
  XNOR2_X1 U6588 ( .A(n5466), .B(n5465), .ZN(n5554) );
  INV_X1 U6589 ( .A(n5554), .ZN(n5471) );
  INV_X1 U6590 ( .A(n5467), .ZN(n5668) );
  NOR2_X1 U6591 ( .A1(n6047), .A2(n6451), .ZN(n5559) );
  AOI21_X1 U6592 ( .B1(n5963), .B2(PHYADDRPOINTER_REG_26__SCAN_IN), .A(n5559), 
        .ZN(n5468) );
  OAI21_X1 U6593 ( .B1(n5973), .B2(n5661), .A(n5468), .ZN(n5469) );
  AOI21_X1 U6594 ( .B1(n5668), .B2(n5515), .A(n5469), .ZN(n5470) );
  OAI21_X1 U6595 ( .B1(n5471), .B2(n5770), .A(n5470), .ZN(U2960) );
  NAND2_X1 U6596 ( .A1(n5473), .A2(n5472), .ZN(n5476) );
  OAI21_X1 U6597 ( .B1(n5476), .B2(n5475), .A(n5474), .ZN(n5562) );
  NAND2_X1 U6598 ( .A1(n5562), .A2(n5968), .ZN(n5480) );
  INV_X1 U6599 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5477) );
  NAND2_X1 U6600 ( .A1(n6032), .A2(REIP_REG_25__SCAN_IN), .ZN(n5563) );
  OAI21_X1 U6601 ( .B1(n5535), .B2(n5477), .A(n5563), .ZN(n5478) );
  AOI21_X1 U6602 ( .B1(n5538), .B2(n5672), .A(n5478), .ZN(n5479) );
  OAI211_X1 U6603 ( .C1(n5673), .C2(n5542), .A(n5480), .B(n5479), .ZN(U2961)
         );
  NAND2_X1 U6604 ( .A1(n5617), .A2(n5481), .ZN(n5518) );
  NAND2_X1 U6605 ( .A1(n5518), .A2(n5482), .ZN(n5484) );
  NAND3_X1 U6606 ( .A1(n3422), .A2(n5579), .A3(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5486) );
  OAI21_X1 U6607 ( .B1(n5512), .B2(n5486), .A(n5485), .ZN(n5487) );
  XNOR2_X1 U6608 ( .A(n5487), .B(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5576)
         );
  NAND2_X1 U6609 ( .A1(n5538), .A2(n5488), .ZN(n5489) );
  NAND2_X1 U6610 ( .A1(n6032), .A2(REIP_REG_23__SCAN_IN), .ZN(n5570) );
  OAI211_X1 U6611 ( .C1(n5535), .C2(n5490), .A(n5489), .B(n5570), .ZN(n5491)
         );
  AOI21_X1 U6612 ( .B1(n5492), .B2(n5515), .A(n5491), .ZN(n5493) );
  OAI21_X1 U6613 ( .B1(n5576), .B2(n5770), .A(n5493), .ZN(U2963) );
  AOI21_X1 U6614 ( .B1(INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n3422), .A(n5494), 
        .ZN(n5495) );
  XNOR2_X1 U6615 ( .A(n5496), .B(n5495), .ZN(n5585) );
  INV_X1 U6616 ( .A(REIP_REG_22__SCAN_IN), .ZN(n5498) );
  NOR2_X1 U6617 ( .A1(n6047), .A2(n5498), .ZN(n5582) );
  AOI21_X1 U6618 ( .B1(n5963), .B2(PHYADDRPOINTER_REG_22__SCAN_IN), .A(n5582), 
        .ZN(n5499) );
  OAI21_X1 U6619 ( .B1(n5973), .B2(n5500), .A(n5499), .ZN(n5501) );
  AOI21_X1 U6620 ( .B1(n5719), .B2(n5515), .A(n5501), .ZN(n5502) );
  OAI21_X1 U6621 ( .B1(n5585), .B2(n5770), .A(n5502), .ZN(U2964) );
  AOI21_X1 U6622 ( .B1(n5505), .B2(n5504), .A(n5503), .ZN(n5592) );
  INV_X1 U6623 ( .A(REIP_REG_21__SCAN_IN), .ZN(n5506) );
  OR2_X1 U6624 ( .A1(n6047), .A2(n5506), .ZN(n5586) );
  OAI21_X1 U6625 ( .B1(n5535), .B2(n5702), .A(n5586), .ZN(n5508) );
  NOR2_X1 U6626 ( .A1(n5705), .A2(n5542), .ZN(n5507) );
  AOI211_X1 U6627 ( .C1(n5538), .C2(n5700), .A(n5508), .B(n5507), .ZN(n5509)
         );
  OAI21_X1 U6628 ( .B1(n5592), .B2(n5770), .A(n5509), .ZN(U2965) );
  XNOR2_X1 U6629 ( .A(n3422), .B(n5510), .ZN(n5511) );
  XNOR2_X1 U6630 ( .A(n5512), .B(n5511), .ZN(n5605) );
  NOR2_X1 U6631 ( .A1(n6047), .A2(n6632), .ZN(n5594) );
  AOI21_X1 U6632 ( .B1(n5963), .B2(PHYADDRPOINTER_REG_20__SCAN_IN), .A(n5594), 
        .ZN(n5513) );
  OAI21_X1 U6633 ( .B1(n5973), .B2(n5710), .A(n5513), .ZN(n5514) );
  AOI21_X1 U6634 ( .B1(n5725), .B2(n5515), .A(n5514), .ZN(n5516) );
  OAI21_X1 U6635 ( .B1(n5605), .B2(n5770), .A(n5516), .ZN(U2966) );
  NAND2_X1 U6636 ( .A1(n5518), .A2(n5517), .ZN(n5521) );
  NAND2_X1 U6637 ( .A1(n5521), .A2(n5520), .ZN(n5519) );
  OAI21_X1 U6638 ( .B1(n5521), .B2(n5520), .A(n5519), .ZN(n5607) );
  NAND2_X1 U6639 ( .A1(n5607), .A2(n5968), .ZN(n5526) );
  NOR2_X1 U6640 ( .A1(n6047), .A2(n6441), .ZN(n5609) );
  INV_X1 U6641 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n5522) );
  NOR2_X1 U6642 ( .A1(n5535), .A2(n5522), .ZN(n5523) );
  AOI211_X1 U6643 ( .C1(n5538), .C2(n5524), .A(n5609), .B(n5523), .ZN(n5525)
         );
  OAI211_X1 U6644 ( .C1(n5542), .C2(n5728), .A(n5526), .B(n5525), .ZN(U2967)
         );
  AND2_X1 U6645 ( .A1(n5617), .A2(n5527), .ZN(n5532) );
  MUX2_X1 U6646 ( .A(n5619), .B(INSTADDRPOINTER_REG_17__SCAN_IN), .S(n3422), 
        .Z(n5531) );
  OR3_X1 U6647 ( .A1(n3422), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5616) );
  INV_X1 U6648 ( .A(n5616), .ZN(n5528) );
  AOI22_X1 U6649 ( .A1(n5529), .A2(n5528), .B1(INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n3422), .ZN(n5615) );
  INV_X1 U6650 ( .A(n5617), .ZN(n5530) );
  OAI22_X1 U6651 ( .A1(n5532), .A2(n5531), .B1(n5615), .B2(n5530), .ZN(n5738)
         );
  NAND2_X1 U6652 ( .A1(n5738), .A2(n5968), .ZN(n5540) );
  INV_X1 U6653 ( .A(REIP_REG_17__SCAN_IN), .ZN(n5533) );
  OAI22_X1 U6654 ( .A1(n5535), .A2(n5534), .B1(n6047), .B2(n5533), .ZN(n5536)
         );
  AOI21_X1 U6655 ( .B1(n5538), .B2(n5537), .A(n5536), .ZN(n5539) );
  OAI211_X1 U6656 ( .C1(n5542), .C2(n5541), .A(n5540), .B(n5539), .ZN(U2969)
         );
  INV_X1 U6657 ( .A(n5660), .ZN(n5551) );
  INV_X1 U6658 ( .A(n5543), .ZN(n5544) );
  NAND3_X1 U6659 ( .A1(n5546), .A2(n5545), .A3(n5544), .ZN(n5547) );
  OAI211_X1 U6660 ( .C1(n5549), .C2(n6586), .A(n5548), .B(n5547), .ZN(n5550)
         );
  AOI21_X1 U6661 ( .B1(n5551), .B2(n6044), .A(n5550), .ZN(n5552) );
  OAI21_X1 U6662 ( .B1(n5553), .B2(n6023), .A(n5552), .ZN(U2990) );
  NAND2_X1 U6663 ( .A1(n5554), .A2(n6050), .ZN(n5561) );
  INV_X1 U6664 ( .A(n5564), .ZN(n5557) );
  AND3_X1 U6665 ( .A1(n5557), .A2(n5556), .A3(n5555), .ZN(n5558) );
  AOI211_X1 U6666 ( .C1(n5566), .C2(INSTADDRPOINTER_REG_26__SCAN_IN), .A(n5559), .B(n5558), .ZN(n5560) );
  OAI211_X1 U6667 ( .C1(n6024), .C2(n5671), .A(n5561), .B(n5560), .ZN(U2992)
         );
  NAND2_X1 U6668 ( .A1(n5562), .A2(n6050), .ZN(n5568) );
  OAI21_X1 U6669 ( .B1(n5564), .B2(INSTADDRPOINTER_REG_25__SCAN_IN), .A(n5563), 
        .ZN(n5565) );
  AOI21_X1 U6670 ( .B1(n5566), .B2(INSTADDRPOINTER_REG_25__SCAN_IN), .A(n5565), 
        .ZN(n5567) );
  OAI211_X1 U6671 ( .C1(n6024), .C2(n5674), .A(n5568), .B(n5567), .ZN(U2993)
         );
  NAND2_X1 U6672 ( .A1(n5569), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5571) );
  OAI211_X1 U6673 ( .C1(INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n5572), .A(n5571), .B(n5570), .ZN(n5573) );
  AOI21_X1 U6674 ( .B1(n5574), .B2(n6044), .A(n5573), .ZN(n5575) );
  OAI21_X1 U6675 ( .B1(n5576), .B2(n6023), .A(n5575), .ZN(U2995) );
  INV_X1 U6676 ( .A(n5577), .ZN(n5590) );
  INV_X1 U6677 ( .A(n5578), .ZN(n5587) );
  NOR3_X1 U6678 ( .A1(n5587), .A2(n5580), .A3(n5579), .ZN(n5581) );
  AOI211_X1 U6679 ( .C1(n5590), .C2(INSTADDRPOINTER_REG_22__SCAN_IN), .A(n5582), .B(n5581), .ZN(n5584) );
  NAND2_X1 U6680 ( .A1(n5694), .A2(n6044), .ZN(n5583) );
  OAI211_X1 U6681 ( .C1(n5585), .C2(n6023), .A(n5584), .B(n5583), .ZN(U2996)
         );
  OAI21_X1 U6682 ( .B1(n5587), .B2(INSTADDRPOINTER_REG_21__SCAN_IN), .A(n5586), 
        .ZN(n5589) );
  NOR2_X1 U6683 ( .A1(n5706), .A2(n6024), .ZN(n5588) );
  AOI211_X1 U6684 ( .C1(INSTADDRPOINTER_REG_21__SCAN_IN), .C2(n5590), .A(n5589), .B(n5588), .ZN(n5591) );
  OAI21_X1 U6685 ( .B1(n5592), .B2(n6023), .A(n5591), .ZN(U2997) );
  INV_X1 U6686 ( .A(n5717), .ZN(n5595) );
  NOR3_X1 U6687 ( .A1(n5602), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .A3(n5613), 
        .ZN(n5593) );
  AOI211_X1 U6688 ( .C1(n5595), .C2(n6044), .A(n5594), .B(n5593), .ZN(n5604)
         );
  INV_X1 U6689 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5619) );
  NOR2_X1 U6690 ( .A1(n5596), .A2(n5619), .ZN(n5599) );
  OAI21_X1 U6691 ( .B1(n5599), .B2(n5598), .A(n5597), .ZN(n5736) );
  AOI21_X1 U6692 ( .B1(n5619), .B2(n5600), .A(n5736), .ZN(n5621) );
  OAI21_X1 U6693 ( .B1(INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n5601), .A(n5621), 
        .ZN(n5606) );
  NOR2_X1 U6694 ( .A1(n5602), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5608)
         );
  OAI21_X1 U6695 ( .B1(n5606), .B2(n5608), .A(INSTADDRPOINTER_REG_20__SCAN_IN), 
        .ZN(n5603) );
  OAI211_X1 U6696 ( .C1(n5605), .C2(n6023), .A(n5604), .B(n5603), .ZN(U2998)
         );
  INV_X1 U6697 ( .A(n5606), .ZN(n5614) );
  NAND2_X1 U6698 ( .A1(n5607), .A2(n6050), .ZN(n5612) );
  AOI211_X1 U6699 ( .C1(n5610), .C2(n6044), .A(n5609), .B(n5608), .ZN(n5611)
         );
  OAI211_X1 U6700 ( .C1(n5614), .C2(n5613), .A(n5612), .B(n5611), .ZN(U2999)
         );
  AOI21_X1 U6701 ( .B1(n5617), .B2(n5616), .A(n5615), .ZN(n5618) );
  INV_X1 U6702 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5620) );
  XNOR2_X1 U6703 ( .A(n5618), .B(n5620), .ZN(n5733) );
  INV_X1 U6704 ( .A(n5733), .ZN(n5626) );
  INV_X1 U6705 ( .A(n5795), .ZN(n5624) );
  NOR3_X1 U6706 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n5619), .A3(n5741), 
        .ZN(n5623) );
  OAI22_X1 U6707 ( .A1(n5621), .A2(n5620), .B1(n6047), .B2(n6543), .ZN(n5622)
         );
  AOI211_X1 U6708 ( .C1(n6044), .C2(n5624), .A(n5623), .B(n5622), .ZN(n5625)
         );
  OAI21_X1 U6709 ( .B1(n5626), .B2(n6023), .A(n5625), .ZN(U3000) );
  OAI21_X1 U6710 ( .B1(n5627), .B2(STATEBS16_REG_SCAN_IN), .A(n6197), .ZN(
        n5629) );
  OAI22_X1 U6711 ( .A1(n5629), .A2(n6192), .B1(n5628), .B2(n5633), .ZN(n5630)
         );
  MUX2_X1 U6712 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n5630), .S(n6055), 
        .Z(U3464) );
  XNOR2_X1 U6713 ( .A(n5631), .B(n6192), .ZN(n5635) );
  INV_X1 U6714 ( .A(n5632), .ZN(n5634) );
  OAI22_X1 U6715 ( .A1(n5635), .A2(n6286), .B1(n5634), .B2(n5633), .ZN(n5636)
         );
  MUX2_X1 U6716 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n5636), .S(n6055), 
        .Z(U3463) );
  INV_X1 U6717 ( .A(n6342), .ZN(n5639) );
  OAI22_X1 U6718 ( .A1(n5639), .A2(n6479), .B1(n5638), .B2(n5637), .ZN(n5640)
         );
  MUX2_X1 U6719 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n5640), .S(n6477), 
        .Z(U3456) );
  AND2_X1 U6720 ( .A1(n5888), .A2(DATAO_REG_31__SCAN_IN), .ZN(U2892) );
  AOI22_X1 U6721 ( .A1(EBX_REG_29__SCAN_IN), .A2(n5865), .B1(
        PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n5870), .ZN(n5641) );
  OAI21_X1 U6722 ( .B1(n5654), .B2(n6458), .A(n5641), .ZN(n5642) );
  AOI21_X1 U6723 ( .B1(n5643), .B2(n5813), .A(n5642), .ZN(n5648) );
  NOR2_X1 U6724 ( .A1(n5644), .A2(n5863), .ZN(n5645) );
  AOI21_X1 U6725 ( .B1(n5646), .B2(n5838), .A(n5645), .ZN(n5647) );
  OAI211_X1 U6726 ( .C1(REIP_REG_29__SCAN_IN), .C2(n5649), .A(n5648), .B(n5647), .ZN(U2798) );
  INV_X1 U6727 ( .A(n5650), .ZN(n5651) );
  AOI22_X1 U6728 ( .A1(n5813), .A2(n5651), .B1(n5865), .B2(EBX_REG_28__SCAN_IN), .ZN(n5653) );
  NAND2_X1 U6729 ( .A1(n5870), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5652)
         );
  OAI211_X1 U6730 ( .C1(n5654), .C2(n5460), .A(n5653), .B(n5652), .ZN(n5655)
         );
  AOI21_X1 U6731 ( .B1(n5656), .B2(n5838), .A(n5655), .ZN(n5659) );
  NAND3_X1 U6732 ( .A1(REIP_REG_27__SCAN_IN), .A2(n5657), .A3(n5460), .ZN(
        n5658) );
  OAI211_X1 U6733 ( .C1(n5863), .C2(n5660), .A(n5659), .B(n5658), .ZN(U2799)
         );
  OAI22_X1 U6734 ( .A1(n5663), .A2(n5662), .B1(n5661), .B2(n5868), .ZN(n5664)
         );
  AOI21_X1 U6735 ( .B1(PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n5870), .A(n5664), 
        .ZN(n5670) );
  NAND2_X1 U6736 ( .A1(n6451), .A2(n5665), .ZN(n5666) );
  AOI22_X1 U6737 ( .A1(n5668), .A2(n5838), .B1(n5667), .B2(n5666), .ZN(n5669)
         );
  OAI211_X1 U6738 ( .C1(n5671), .C2(n5863), .A(n5670), .B(n5669), .ZN(U2801)
         );
  AOI22_X1 U6739 ( .A1(EBX_REG_25__SCAN_IN), .A2(n5865), .B1(
        PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n5870), .ZN(n5681) );
  AOI22_X1 U6740 ( .A1(n5672), .A2(n5813), .B1(REIP_REG_25__SCAN_IN), .B2(
        n5685), .ZN(n5680) );
  INV_X1 U6741 ( .A(n5673), .ZN(n5676) );
  INV_X1 U6742 ( .A(n5674), .ZN(n5675) );
  AOI22_X1 U6743 ( .A1(n5676), .A2(n5838), .B1(n5675), .B2(n5866), .ZN(n5679)
         );
  OAI211_X1 U6744 ( .C1(REIP_REG_24__SCAN_IN), .C2(REIP_REG_25__SCAN_IN), .A(
        n5689), .B(n5677), .ZN(n5678) );
  NAND4_X1 U6745 ( .A1(n5681), .A2(n5680), .A3(n5679), .A4(n5678), .ZN(U2802)
         );
  INV_X1 U6746 ( .A(REIP_REG_24__SCAN_IN), .ZN(n6449) );
  AOI22_X1 U6747 ( .A1(n5870), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .B1(
        EBX_REG_24__SCAN_IN), .B2(n5865), .ZN(n5682) );
  OAI21_X1 U6748 ( .B1(n5868), .B2(n5683), .A(n5682), .ZN(n5684) );
  AOI21_X1 U6749 ( .B1(n5685), .B2(REIP_REG_24__SCAN_IN), .A(n5684), .ZN(n5686) );
  OAI21_X1 U6750 ( .B1(n5687), .B2(n5826), .A(n5686), .ZN(n5688) );
  AOI21_X1 U6751 ( .B1(n5689), .B2(n6449), .A(n5688), .ZN(n5690) );
  OAI21_X1 U6752 ( .B1(n5691), .B2(n5863), .A(n5690), .ZN(U2803) );
  AOI22_X1 U6753 ( .A1(EBX_REG_22__SCAN_IN), .A2(n5865), .B1(
        PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n5870), .ZN(n5699) );
  NOR2_X1 U6754 ( .A1(n5692), .A2(n5853), .ZN(n5714) );
  AOI22_X1 U6755 ( .A1(n5693), .A2(n5813), .B1(REIP_REG_22__SCAN_IN), .B2(
        n5714), .ZN(n5698) );
  AOI22_X1 U6756 ( .A1(n5719), .A2(n5838), .B1(n5694), .B2(n5866), .ZN(n5697)
         );
  OAI211_X1 U6757 ( .C1(REIP_REG_22__SCAN_IN), .C2(REIP_REG_21__SCAN_IN), .A(
        n5704), .B(n5695), .ZN(n5696) );
  NAND4_X1 U6758 ( .A1(n5699), .A2(n5698), .A3(n5697), .A4(n5696), .ZN(U2805)
         );
  AOI22_X1 U6759 ( .A1(EBX_REG_21__SCAN_IN), .A2(n5865), .B1(n5700), .B2(n5813), .ZN(n5701) );
  OAI21_X1 U6760 ( .B1(n5702), .B2(n5834), .A(n5701), .ZN(n5703) );
  AOI221_X1 U6761 ( .B1(n5714), .B2(REIP_REG_21__SCAN_IN), .C1(n5704), .C2(
        n5506), .A(n5703), .ZN(n5709) );
  INV_X1 U6762 ( .A(n5705), .ZN(n5722) );
  INV_X1 U6763 ( .A(n5706), .ZN(n5707) );
  AOI22_X1 U6764 ( .A1(n5722), .A2(n5838), .B1(n5707), .B2(n5866), .ZN(n5708)
         );
  NAND2_X1 U6765 ( .A1(n5709), .A2(n5708), .ZN(U2806) );
  INV_X1 U6766 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n6565) );
  OAI22_X1 U6767 ( .A1(n6565), .A2(n5834), .B1(n5710), .B2(n5868), .ZN(n5711)
         );
  AOI21_X1 U6768 ( .B1(EBX_REG_20__SCAN_IN), .B2(n5865), .A(n5711), .ZN(n5716)
         );
  NAND2_X1 U6769 ( .A1(n6632), .A2(n5712), .ZN(n5713) );
  AOI22_X1 U6770 ( .A1(n5725), .A2(n5838), .B1(n5714), .B2(n5713), .ZN(n5715)
         );
  OAI211_X1 U6771 ( .C1(n5717), .C2(n5863), .A(n5716), .B(n5715), .ZN(U2807)
         );
  INV_X1 U6772 ( .A(n5718), .ZN(n5882) );
  AOI22_X1 U6773 ( .A1(n5719), .A2(n5882), .B1(n5881), .B2(DATAI_22_), .ZN(
        n5721) );
  AOI22_X1 U6774 ( .A1(n5885), .A2(DATAI_6_), .B1(n5884), .B2(
        EAX_REG_22__SCAN_IN), .ZN(n5720) );
  NAND2_X1 U6775 ( .A1(n5721), .A2(n5720), .ZN(U2869) );
  AOI22_X1 U6776 ( .A1(n5722), .A2(n5882), .B1(n5881), .B2(DATAI_21_), .ZN(
        n5724) );
  AOI22_X1 U6777 ( .A1(n5885), .A2(DATAI_5_), .B1(n5884), .B2(
        EAX_REG_21__SCAN_IN), .ZN(n5723) );
  NAND2_X1 U6778 ( .A1(n5724), .A2(n5723), .ZN(U2870) );
  AOI22_X1 U6779 ( .A1(n5725), .A2(n5882), .B1(n5881), .B2(DATAI_20_), .ZN(
        n5727) );
  AOI22_X1 U6780 ( .A1(n5885), .A2(DATAI_4_), .B1(n5884), .B2(
        EAX_REG_20__SCAN_IN), .ZN(n5726) );
  NAND2_X1 U6781 ( .A1(n5727), .A2(n5726), .ZN(U2871) );
  INV_X1 U6782 ( .A(n5728), .ZN(n5729) );
  AOI22_X1 U6783 ( .A1(n5729), .A2(n5882), .B1(n5881), .B2(DATAI_19_), .ZN(
        n5731) );
  AOI22_X1 U6784 ( .A1(n5885), .A2(DATAI_3_), .B1(n5884), .B2(
        EAX_REG_19__SCAN_IN), .ZN(n5730) );
  NAND2_X1 U6785 ( .A1(n5731), .A2(n5730), .ZN(U2872) );
  AOI22_X1 U6786 ( .A1(n6032), .A2(REIP_REG_18__SCAN_IN), .B1(n5963), .B2(
        PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n5735) );
  AOI22_X1 U6787 ( .A1(n5733), .A2(n5968), .B1(n5515), .B2(n5878), .ZN(n5734)
         );
  OAI211_X1 U6788 ( .C1(n5973), .C2(n5791), .A(n5735), .B(n5734), .ZN(U2968)
         );
  AOI22_X1 U6789 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n5736), .B1(n6032), .B2(REIP_REG_17__SCAN_IN), .ZN(n5740) );
  AOI22_X1 U6790 ( .A1(n5738), .A2(n6050), .B1(n6044), .B2(n5737), .ZN(n5739)
         );
  OAI211_X1 U6791 ( .C1(INSTADDRPOINTER_REG_17__SCAN_IN), .C2(n5741), .A(n5740), .B(n5739), .ZN(U3001) );
  INV_X1 U6792 ( .A(n5742), .ZN(n5749) );
  AOI21_X1 U6793 ( .B1(n5744), .B2(n6044), .A(n5743), .ZN(n5748) );
  AOI22_X1 U6794 ( .A1(n5746), .A2(n6050), .B1(INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n5745), .ZN(n5747) );
  OAI211_X1 U6795 ( .C1(INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n5749), .A(n5748), .B(n5747), .ZN(U3003) );
  AOI21_X1 U6796 ( .B1(n5751), .B2(n6044), .A(n5750), .ZN(n5755) );
  NOR2_X1 U6797 ( .A1(INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n5974), .ZN(n5752)
         );
  AOI22_X1 U6798 ( .A1(n5753), .A2(n6050), .B1(n5752), .B2(n5984), .ZN(n5754)
         );
  OAI211_X1 U6799 ( .C1(n5756), .C2(n3404), .A(n5755), .B(n5754), .ZN(U3005)
         );
  INV_X1 U6800 ( .A(n5757), .ZN(n5759) );
  NAND4_X1 U6801 ( .A1(n5759), .A2(n5758), .A3(n6384), .A4(n5851), .ZN(n5760)
         );
  OAI21_X1 U6802 ( .B1(n6477), .B2(n4498), .A(n5760), .ZN(U3455) );
  AOI21_X1 U6803 ( .B1(STATE_REG_1__SCAN_IN), .B2(n6584), .A(n4130), .ZN(n5768) );
  INV_X1 U6804 ( .A(ADS_N_REG_SCAN_IN), .ZN(n5761) );
  NAND2_X1 U6805 ( .A1(n4130), .A2(STATE_REG_1__SCAN_IN), .ZN(n6489) );
  AOI21_X1 U6806 ( .B1(n5768), .B2(n5761), .A(n5766), .ZN(U2789) );
  NAND2_X1 U6807 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n6497), .ZN(n5765) );
  INV_X1 U6808 ( .A(n5762), .ZN(n5763) );
  OAI21_X1 U6809 ( .B1(n5763), .B2(n6369), .A(CODEFETCH_REG_SCAN_IN), .ZN(
        n5764) );
  OAI21_X1 U6810 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n5765), .A(n5764), .ZN(
        U2790) );
  NOR2_X1 U6811 ( .A1(STATE_REG_0__SCAN_IN), .A2(STATE_REG_2__SCAN_IN), .ZN(
        n5769) );
  INV_X1 U6812 ( .A(n6489), .ZN(n5766) );
  INV_X1 U6813 ( .A(n5766), .ZN(n6502) );
  OAI21_X1 U6814 ( .B1(D_C_N_REG_SCAN_IN), .B2(n5769), .A(n6502), .ZN(n5767)
         );
  OAI21_X1 U6815 ( .B1(CODEFETCH_REG_SCAN_IN), .B2(n6489), .A(n5767), .ZN(
        U2791) );
  NOR2_X1 U6816 ( .A1(n5766), .A2(n5768), .ZN(n6466) );
  OAI21_X1 U6817 ( .B1(BS16_N), .B2(n5769), .A(n6466), .ZN(n6464) );
  OAI21_X1 U6818 ( .B1(n6466), .B2(n6234), .A(n6464), .ZN(U2792) );
  OAI21_X1 U6819 ( .B1(n5772), .B2(n5771), .A(n5770), .ZN(U2793) );
  NOR4_X1 U6820 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(
        DATAWIDTH_REG_19__SCAN_IN), .A3(DATAWIDTH_REG_20__SCAN_IN), .A4(
        DATAWIDTH_REG_21__SCAN_IN), .ZN(n5776) );
  NOR4_X1 U6821 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(
        DATAWIDTH_REG_15__SCAN_IN), .A3(DATAWIDTH_REG_16__SCAN_IN), .A4(
        DATAWIDTH_REG_17__SCAN_IN), .ZN(n5775) );
  NOR4_X1 U6822 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(
        DATAWIDTH_REG_29__SCAN_IN), .A3(DATAWIDTH_REG_30__SCAN_IN), .A4(
        DATAWIDTH_REG_31__SCAN_IN), .ZN(n5774) );
  NOR4_X1 U6823 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(
        DATAWIDTH_REG_23__SCAN_IN), .A3(DATAWIDTH_REG_25__SCAN_IN), .A4(
        DATAWIDTH_REG_26__SCAN_IN), .ZN(n5773) );
  NAND4_X1 U6824 ( .A1(n5776), .A2(n5775), .A3(n5774), .A4(n5773), .ZN(n5782)
         );
  NOR4_X1 U6825 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(DATAWIDTH_REG_8__SCAN_IN), .A3(DATAWIDTH_REG_3__SCAN_IN), .A4(DATAWIDTH_REG_2__SCAN_IN), .ZN(n5780) );
  AOI211_X1 U6826 ( .C1(DATAWIDTH_REG_0__SCAN_IN), .C2(
        DATAWIDTH_REG_1__SCAN_IN), .A(DATAWIDTH_REG_24__SCAN_IN), .B(
        DATAWIDTH_REG_12__SCAN_IN), .ZN(n5779) );
  NOR4_X1 U6827 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(DATAWIDTH_REG_10__SCAN_IN), .A3(DATAWIDTH_REG_11__SCAN_IN), .A4(DATAWIDTH_REG_13__SCAN_IN), .ZN(n5778)
         );
  NOR4_X1 U6828 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(DATAWIDTH_REG_5__SCAN_IN), 
        .A3(DATAWIDTH_REG_6__SCAN_IN), .A4(DATAWIDTH_REG_7__SCAN_IN), .ZN(
        n5777) );
  NAND4_X1 U6829 ( .A1(n5780), .A2(n5779), .A3(n5778), .A4(n5777), .ZN(n5781)
         );
  NOR2_X1 U6830 ( .A1(n5782), .A2(n5781), .ZN(n6487) );
  INV_X1 U6831 ( .A(BYTEENABLE_REG_1__SCAN_IN), .ZN(n5784) );
  NOR3_X1 U6832 ( .A1(REIP_REG_0__SCAN_IN), .A2(DATAWIDTH_REG_0__SCAN_IN), 
        .A3(DATAWIDTH_REG_1__SCAN_IN), .ZN(n5785) );
  OAI21_X1 U6833 ( .B1(REIP_REG_1__SCAN_IN), .B2(n5785), .A(n6487), .ZN(n5783)
         );
  OAI21_X1 U6834 ( .B1(n6487), .B2(n5784), .A(n5783), .ZN(U2794) );
  INV_X1 U6835 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6465) );
  AOI21_X1 U6836 ( .B1(n6580), .B2(n6465), .A(n5785), .ZN(n5787) );
  INV_X1 U6837 ( .A(BYTEENABLE_REG_3__SCAN_IN), .ZN(n5786) );
  INV_X1 U6838 ( .A(n6487), .ZN(n6484) );
  AOI22_X1 U6839 ( .A1(n6487), .A2(n5787), .B1(n5786), .B2(n6484), .ZN(U2795)
         );
  AOI22_X1 U6840 ( .A1(EBX_REG_18__SCAN_IN), .A2(n5865), .B1(
        REIP_REG_18__SCAN_IN), .B2(n5788), .ZN(n5790) );
  AOI21_X1 U6841 ( .B1(n5870), .B2(PHYADDRPOINTER_REG_18__SCAN_IN), .A(n5845), 
        .ZN(n5789) );
  OAI211_X1 U6842 ( .C1(n5791), .C2(n5868), .A(n5790), .B(n5789), .ZN(n5792)
         );
  AOI211_X1 U6843 ( .C1(n5878), .C2(n5838), .A(n5793), .B(n5792), .ZN(n5794)
         );
  OAI21_X1 U6844 ( .B1(n5863), .B2(n5795), .A(n5794), .ZN(U2809) );
  AOI21_X1 U6845 ( .B1(n5807), .B2(n5796), .A(REIP_REG_14__SCAN_IN), .ZN(n5806) );
  INV_X1 U6846 ( .A(n5797), .ZN(n5805) );
  INV_X1 U6847 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n5799) );
  OAI22_X1 U6848 ( .A1(n5799), .A2(n5834), .B1(n5863), .B2(n5798), .ZN(n5800)
         );
  AOI211_X1 U6849 ( .C1(n5865), .C2(EBX_REG_14__SCAN_IN), .A(n5845), .B(n5800), 
        .ZN(n5804) );
  AOI22_X1 U6850 ( .A1(n5802), .A2(n5838), .B1(n5813), .B2(n5801), .ZN(n5803)
         );
  OAI211_X1 U6851 ( .C1(n5806), .C2(n5805), .A(n5804), .B(n5803), .ZN(U2813)
         );
  INV_X1 U6852 ( .A(n5807), .ZN(n5817) );
  OAI21_X1 U6853 ( .B1(n5834), .B2(n5808), .A(n5854), .ZN(n5811) );
  OAI22_X1 U6854 ( .A1(n5863), .A2(n5976), .B1(n6431), .B2(n5809), .ZN(n5810)
         );
  AOI211_X1 U6855 ( .C1(EBX_REG_12__SCAN_IN), .C2(n5865), .A(n5811), .B(n5810), 
        .ZN(n5816) );
  AOI22_X1 U6856 ( .A1(n5814), .A2(n5838), .B1(n5813), .B2(n5812), .ZN(n5815)
         );
  OAI211_X1 U6857 ( .C1(REIP_REG_12__SCAN_IN), .C2(n5817), .A(n5816), .B(n5815), .ZN(U2815) );
  AOI21_X1 U6858 ( .B1(n6427), .B2(n4914), .A(n5818), .ZN(n5820) );
  AOI22_X1 U6859 ( .A1(REIP_REG_10__SCAN_IN), .A2(n5821), .B1(n5820), .B2(
        n5819), .ZN(n5831) );
  OAI22_X1 U6860 ( .A1(n6534), .A2(n5834), .B1(n5863), .B2(n5822), .ZN(n5823)
         );
  AOI211_X1 U6861 ( .C1(n5865), .C2(EBX_REG_10__SCAN_IN), .A(n5845), .B(n5823), 
        .ZN(n5830) );
  INV_X1 U6862 ( .A(n5824), .ZN(n5825) );
  OAI22_X1 U6863 ( .A1(n5827), .A2(n5826), .B1(n5868), .B2(n5825), .ZN(n5828)
         );
  INV_X1 U6864 ( .A(n5828), .ZN(n5829) );
  NAND3_X1 U6865 ( .A1(n5831), .A2(n5830), .A3(n5829), .ZN(U2817) );
  INV_X1 U6866 ( .A(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n5833) );
  AOI22_X1 U6867 ( .A1(EBX_REG_7__SCAN_IN), .A2(n5865), .B1(n5866), .B2(n6007), 
        .ZN(n5832) );
  OAI211_X1 U6868 ( .C1(n5834), .C2(n5833), .A(n5854), .B(n5832), .ZN(n5837)
         );
  NOR3_X1 U6869 ( .A1(REIP_REG_7__SCAN_IN), .A2(n4981), .A3(n5835), .ZN(n5836)
         );
  AOI211_X1 U6870 ( .C1(n5943), .C2(n5838), .A(n5837), .B(n5836), .ZN(n5841)
         );
  OAI21_X1 U6871 ( .B1(n5839), .B2(n5847), .A(REIP_REG_7__SCAN_IN), .ZN(n5840)
         );
  OAI211_X1 U6872 ( .C1(n5868), .C2(n5946), .A(n5841), .B(n5840), .ZN(U2820)
         );
  INV_X1 U6873 ( .A(n5842), .ZN(n6016) );
  AOI22_X1 U6874 ( .A1(PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n5870), .B1(n5866), 
        .B2(n6016), .ZN(n5843) );
  INV_X1 U6875 ( .A(n5843), .ZN(n5844) );
  AOI211_X1 U6876 ( .C1(n5865), .C2(EBX_REG_5__SCAN_IN), .A(n5845), .B(n5844), 
        .ZN(n5849) );
  OAI21_X1 U6877 ( .B1(n5855), .B2(n6419), .A(n6421), .ZN(n5846) );
  AOI22_X1 U6878 ( .A1(n5847), .A2(n5846), .B1(n5951), .B2(n5874), .ZN(n5848)
         );
  OAI211_X1 U6879 ( .C1(n5954), .C2(n5868), .A(n5849), .B(n5848), .ZN(U2822)
         );
  AOI22_X1 U6880 ( .A1(EBX_REG_4__SCAN_IN), .A2(n5865), .B1(n5851), .B2(n5850), 
        .ZN(n5862) );
  OR2_X1 U6881 ( .A1(n5853), .A2(n5852), .ZN(n5877) );
  OAI221_X1 U6882 ( .B1(REIP_REG_4__SCAN_IN), .B2(n5855), .C1(n6419), .C2(
        n5877), .A(n5854), .ZN(n5860) );
  OAI22_X1 U6883 ( .A1(n5858), .A2(n5857), .B1(n5856), .B2(n5868), .ZN(n5859)
         );
  AOI211_X1 U6884 ( .C1(PHYADDRPOINTER_REG_4__SCAN_IN), .C2(n5870), .A(n5860), 
        .B(n5859), .ZN(n5861) );
  OAI211_X1 U6885 ( .C1(n5863), .C2(n6025), .A(n5862), .B(n5861), .ZN(U2823)
         );
  NAND2_X1 U6886 ( .A1(n5864), .A2(REIP_REG_2__SCAN_IN), .ZN(n5876) );
  AOI22_X1 U6887 ( .A1(n6033), .A2(n5866), .B1(n5865), .B2(EBX_REG_3__SCAN_IN), 
        .ZN(n5867) );
  OAI21_X1 U6888 ( .B1(n5868), .B2(n5962), .A(n5867), .ZN(n5869) );
  AOI21_X1 U6889 ( .B1(PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n5870), .A(n5869), 
        .ZN(n5871) );
  OAI21_X1 U6890 ( .B1(n6229), .B2(n5872), .A(n5871), .ZN(n5873) );
  AOI21_X1 U6891 ( .B1(n5959), .B2(n5874), .A(n5873), .ZN(n5875) );
  OAI221_X1 U6892 ( .B1(n5877), .B2(n6590), .C1(n5877), .C2(n5876), .A(n5875), 
        .ZN(U2824) );
  AOI22_X1 U6893 ( .A1(n5878), .A2(n5882), .B1(n5881), .B2(DATAI_18_), .ZN(
        n5880) );
  AOI22_X1 U6894 ( .A1(n5885), .A2(DATAI_2_), .B1(n5884), .B2(
        EAX_REG_18__SCAN_IN), .ZN(n5879) );
  NAND2_X1 U6895 ( .A1(n5880), .A2(n5879), .ZN(U2873) );
  AOI22_X1 U6896 ( .A1(n5883), .A2(n5882), .B1(n5881), .B2(DATAI_16_), .ZN(
        n5887) );
  AOI22_X1 U6897 ( .A1(n5885), .A2(DATAI_0_), .B1(n5884), .B2(
        EAX_REG_16__SCAN_IN), .ZN(n5886) );
  NAND2_X1 U6898 ( .A1(n5887), .A2(n5886), .ZN(U2875) );
  AOI22_X1 U6899 ( .A1(n6493), .A2(LWORD_REG_15__SCAN_IN), .B1(n5888), .B2(
        DATAO_REG_15__SCAN_IN), .ZN(n5889) );
  OAI21_X1 U6900 ( .B1(n5890), .B2(n5920), .A(n5889), .ZN(U2908) );
  INV_X1 U6901 ( .A(EAX_REG_14__SCAN_IN), .ZN(n5892) );
  AOI22_X1 U6902 ( .A1(n6493), .A2(LWORD_REG_14__SCAN_IN), .B1(n5917), .B2(
        DATAO_REG_14__SCAN_IN), .ZN(n5891) );
  OAI21_X1 U6903 ( .B1(n5892), .B2(n5920), .A(n5891), .ZN(U2909) );
  INV_X1 U6904 ( .A(EAX_REG_13__SCAN_IN), .ZN(n5894) );
  AOI22_X1 U6905 ( .A1(n6493), .A2(LWORD_REG_13__SCAN_IN), .B1(n5917), .B2(
        DATAO_REG_13__SCAN_IN), .ZN(n5893) );
  OAI21_X1 U6906 ( .B1(n5894), .B2(n5920), .A(n5893), .ZN(U2910) );
  INV_X1 U6907 ( .A(EAX_REG_12__SCAN_IN), .ZN(n5896) );
  AOI22_X1 U6908 ( .A1(n6493), .A2(LWORD_REG_12__SCAN_IN), .B1(n5917), .B2(
        DATAO_REG_12__SCAN_IN), .ZN(n5895) );
  OAI21_X1 U6909 ( .B1(n5896), .B2(n5920), .A(n5895), .ZN(U2911) );
  INV_X1 U6910 ( .A(EAX_REG_11__SCAN_IN), .ZN(n5898) );
  AOI22_X1 U6911 ( .A1(n6493), .A2(LWORD_REG_11__SCAN_IN), .B1(n5917), .B2(
        DATAO_REG_11__SCAN_IN), .ZN(n5897) );
  OAI21_X1 U6912 ( .B1(n5898), .B2(n5920), .A(n5897), .ZN(U2912) );
  INV_X1 U6913 ( .A(EAX_REG_10__SCAN_IN), .ZN(n5900) );
  AOI22_X1 U6914 ( .A1(n6493), .A2(LWORD_REG_10__SCAN_IN), .B1(n5917), .B2(
        DATAO_REG_10__SCAN_IN), .ZN(n5899) );
  OAI21_X1 U6915 ( .B1(n5900), .B2(n5920), .A(n5899), .ZN(U2913) );
  INV_X1 U6916 ( .A(EAX_REG_9__SCAN_IN), .ZN(n5902) );
  AOI22_X1 U6917 ( .A1(n6493), .A2(LWORD_REG_9__SCAN_IN), .B1(n5917), .B2(
        DATAO_REG_9__SCAN_IN), .ZN(n5901) );
  OAI21_X1 U6918 ( .B1(n5902), .B2(n5920), .A(n5901), .ZN(U2914) );
  INV_X1 U6919 ( .A(EAX_REG_8__SCAN_IN), .ZN(n5904) );
  AOI22_X1 U6920 ( .A1(n6493), .A2(LWORD_REG_8__SCAN_IN), .B1(n5917), .B2(
        DATAO_REG_8__SCAN_IN), .ZN(n5903) );
  OAI21_X1 U6921 ( .B1(n5904), .B2(n5920), .A(n5903), .ZN(U2915) );
  INV_X1 U6922 ( .A(EAX_REG_7__SCAN_IN), .ZN(n5906) );
  AOI22_X1 U6923 ( .A1(n6493), .A2(LWORD_REG_7__SCAN_IN), .B1(n5917), .B2(
        DATAO_REG_7__SCAN_IN), .ZN(n5905) );
  OAI21_X1 U6924 ( .B1(n5906), .B2(n5920), .A(n5905), .ZN(U2916) );
  INV_X1 U6925 ( .A(EAX_REG_6__SCAN_IN), .ZN(n5908) );
  AOI22_X1 U6926 ( .A1(n6493), .A2(LWORD_REG_6__SCAN_IN), .B1(n5917), .B2(
        DATAO_REG_6__SCAN_IN), .ZN(n5907) );
  OAI21_X1 U6927 ( .B1(n5908), .B2(n5920), .A(n5907), .ZN(U2917) );
  AOI22_X1 U6928 ( .A1(n6493), .A2(LWORD_REG_5__SCAN_IN), .B1(n5917), .B2(
        DATAO_REG_5__SCAN_IN), .ZN(n5909) );
  OAI21_X1 U6929 ( .B1(n4614), .B2(n5920), .A(n5909), .ZN(U2918) );
  AOI22_X1 U6930 ( .A1(n6493), .A2(LWORD_REG_4__SCAN_IN), .B1(n5917), .B2(
        DATAO_REG_4__SCAN_IN), .ZN(n5910) );
  OAI21_X1 U6931 ( .B1(n5911), .B2(n5920), .A(n5910), .ZN(U2919) );
  AOI22_X1 U6932 ( .A1(n6493), .A2(LWORD_REG_3__SCAN_IN), .B1(n5917), .B2(
        DATAO_REG_3__SCAN_IN), .ZN(n5912) );
  OAI21_X1 U6933 ( .B1(n5913), .B2(n5920), .A(n5912), .ZN(U2920) );
  AOI22_X1 U6934 ( .A1(n6493), .A2(LWORD_REG_2__SCAN_IN), .B1(
        DATAO_REG_2__SCAN_IN), .B2(n5917), .ZN(n5914) );
  OAI21_X1 U6935 ( .B1(n5915), .B2(n5920), .A(n5914), .ZN(U2921) );
  AOI22_X1 U6936 ( .A1(n6493), .A2(LWORD_REG_1__SCAN_IN), .B1(n5917), .B2(
        DATAO_REG_1__SCAN_IN), .ZN(n5916) );
  OAI21_X1 U6937 ( .B1(n6540), .B2(n5920), .A(n5916), .ZN(U2922) );
  AOI22_X1 U6938 ( .A1(n6493), .A2(LWORD_REG_0__SCAN_IN), .B1(n5917), .B2(
        DATAO_REG_0__SCAN_IN), .ZN(n5919) );
  OAI21_X1 U6939 ( .B1(n5921), .B2(n5920), .A(n5919), .ZN(U2923) );
  INV_X1 U6940 ( .A(DATAI_6_), .ZN(n6646) );
  AOI22_X1 U6941 ( .A1(LWORD_REG_6__SCAN_IN), .A2(n6668), .B1(n6667), .B2(
        EAX_REG_6__SCAN_IN), .ZN(n5922) );
  OAI21_X1 U6942 ( .B1(n5928), .B2(n6646), .A(n5922), .ZN(U2945) );
  INV_X1 U6943 ( .A(DATAI_7_), .ZN(n5924) );
  AOI22_X1 U6944 ( .A1(LWORD_REG_7__SCAN_IN), .A2(n6668), .B1(n6667), .B2(
        EAX_REG_7__SCAN_IN), .ZN(n5923) );
  OAI21_X1 U6945 ( .B1(n5928), .B2(n5924), .A(n5923), .ZN(U2946) );
  AOI22_X1 U6946 ( .A1(LWORD_REG_8__SCAN_IN), .A2(n6668), .B1(n6667), .B2(
        EAX_REG_8__SCAN_IN), .ZN(n5926) );
  NAND2_X1 U6947 ( .A1(n5936), .A2(DATAI_8_), .ZN(n5925) );
  NAND2_X1 U6948 ( .A1(n5926), .A2(n5925), .ZN(U2947) );
  INV_X1 U6949 ( .A(DATAI_9_), .ZN(n6557) );
  AOI22_X1 U6950 ( .A1(LWORD_REG_9__SCAN_IN), .A2(n6668), .B1(n6667), .B2(
        EAX_REG_9__SCAN_IN), .ZN(n5927) );
  OAI21_X1 U6951 ( .B1(n5928), .B2(n6557), .A(n5927), .ZN(U2948) );
  AOI22_X1 U6952 ( .A1(LWORD_REG_10__SCAN_IN), .A2(n6668), .B1(n6667), .B2(
        EAX_REG_10__SCAN_IN), .ZN(n5929) );
  NAND2_X1 U6953 ( .A1(n5936), .A2(DATAI_10_), .ZN(n6670) );
  NAND2_X1 U6954 ( .A1(n5929), .A2(n6670), .ZN(U2949) );
  AOI22_X1 U6955 ( .A1(LWORD_REG_11__SCAN_IN), .A2(n6668), .B1(n6667), .B2(
        EAX_REG_11__SCAN_IN), .ZN(n5931) );
  NAND2_X1 U6956 ( .A1(n5936), .A2(DATAI_11_), .ZN(n5930) );
  NAND2_X1 U6957 ( .A1(n5931), .A2(n5930), .ZN(U2950) );
  AOI22_X1 U6958 ( .A1(LWORD_REG_12__SCAN_IN), .A2(n6668), .B1(n6667), .B2(
        EAX_REG_12__SCAN_IN), .ZN(n5933) );
  NAND2_X1 U6959 ( .A1(n5936), .A2(DATAI_12_), .ZN(n5932) );
  NAND2_X1 U6960 ( .A1(n5933), .A2(n5932), .ZN(U2951) );
  AOI22_X1 U6961 ( .A1(LWORD_REG_13__SCAN_IN), .A2(n6668), .B1(n6667), .B2(
        EAX_REG_13__SCAN_IN), .ZN(n5935) );
  NAND2_X1 U6962 ( .A1(n5936), .A2(DATAI_13_), .ZN(n5934) );
  NAND2_X1 U6963 ( .A1(n5935), .A2(n5934), .ZN(U2952) );
  AOI22_X1 U6964 ( .A1(LWORD_REG_14__SCAN_IN), .A2(n6668), .B1(n6667), .B2(
        EAX_REG_14__SCAN_IN), .ZN(n5938) );
  NAND2_X1 U6965 ( .A1(n5936), .A2(DATAI_14_), .ZN(n5937) );
  NAND2_X1 U6966 ( .A1(n5938), .A2(n5937), .ZN(U2953) );
  AOI22_X1 U6967 ( .A1(n6032), .A2(REIP_REG_7__SCAN_IN), .B1(n5963), .B2(
        PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n5945) );
  OAI21_X1 U6968 ( .B1(n5941), .B2(n5940), .A(n5939), .ZN(n5942) );
  INV_X1 U6969 ( .A(n5942), .ZN(n6010) );
  AOI22_X1 U6970 ( .A1(n6010), .A2(n5968), .B1(n5515), .B2(n5943), .ZN(n5944)
         );
  OAI211_X1 U6971 ( .C1(n5973), .C2(n5946), .A(n5945), .B(n5944), .ZN(U2979)
         );
  AOI22_X1 U6972 ( .A1(n6032), .A2(REIP_REG_5__SCAN_IN), .B1(n5963), .B2(
        PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n5953) );
  OAI21_X1 U6973 ( .B1(n5949), .B2(n5948), .A(n5947), .ZN(n5950) );
  INV_X1 U6974 ( .A(n5950), .ZN(n6017) );
  AOI22_X1 U6975 ( .A1(n6017), .A2(n5968), .B1(n5515), .B2(n5951), .ZN(n5952)
         );
  OAI211_X1 U6976 ( .C1(n5973), .C2(n5954), .A(n5953), .B(n5952), .ZN(U2981)
         );
  AOI22_X1 U6977 ( .A1(n6032), .A2(REIP_REG_3__SCAN_IN), .B1(n5963), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n5961) );
  OR2_X1 U6978 ( .A1(n5956), .A2(n5955), .ZN(n5957) );
  AND2_X1 U6979 ( .A1(n5958), .A2(n5957), .ZN(n6034) );
  AOI22_X1 U6980 ( .A1(n5959), .A2(n5515), .B1(n5968), .B2(n6034), .ZN(n5960)
         );
  OAI211_X1 U6981 ( .C1(n5973), .C2(n5962), .A(n5961), .B(n5960), .ZN(U2983)
         );
  AOI22_X1 U6982 ( .A1(n6032), .A2(REIP_REG_2__SCAN_IN), .B1(n5963), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n5971) );
  XNOR2_X1 U6983 ( .A(n5965), .B(n5964), .ZN(n5967) );
  XNOR2_X1 U6984 ( .A(n5967), .B(n5966), .ZN(n6051) );
  AOI22_X1 U6985 ( .A1(n5969), .A2(n5515), .B1(n5968), .B2(n6051), .ZN(n5970)
         );
  OAI211_X1 U6986 ( .C1(n5973), .C2(n5972), .A(n5971), .B(n5970), .ZN(U2984)
         );
  AOI21_X1 U6987 ( .B1(INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n5984), .A(
        INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n5981) );
  OAI21_X1 U6988 ( .B1(n5975), .B2(n6040), .A(n5974), .ZN(n5980) );
  OAI22_X1 U6989 ( .A1(n5977), .A2(n6023), .B1(n6024), .B2(n5976), .ZN(n5978)
         );
  AOI21_X1 U6990 ( .B1(n6032), .B2(REIP_REG_12__SCAN_IN), .A(n5978), .ZN(n5979) );
  OAI221_X1 U6991 ( .B1(n5981), .B2(n5989), .C1(n5981), .C2(n5980), .A(n5979), 
        .ZN(U3006) );
  AOI21_X1 U6992 ( .B1(n5983), .B2(n6044), .A(n5982), .ZN(n5987) );
  AOI22_X1 U6993 ( .A1(n6050), .A2(n5985), .B1(n5988), .B2(n5984), .ZN(n5986)
         );
  OAI211_X1 U6994 ( .C1(n5989), .C2(n5988), .A(n5987), .B(n5986), .ZN(U3007)
         );
  INV_X1 U6995 ( .A(n5990), .ZN(n5998) );
  AOI21_X1 U6996 ( .B1(n5992), .B2(n6044), .A(n5991), .ZN(n5996) );
  AOI22_X1 U6997 ( .A1(n5994), .A2(n6050), .B1(n5993), .B2(n5997), .ZN(n5995)
         );
  OAI211_X1 U6998 ( .C1(n5998), .C2(n5997), .A(n5996), .B(n5995), .ZN(U3009)
         );
  INV_X1 U6999 ( .A(n5999), .ZN(n6004) );
  OAI22_X1 U7000 ( .A1(n6024), .A2(n6000), .B1(n6424), .B2(n6047), .ZN(n6003)
         );
  AOI211_X1 U7001 ( .C1(n6570), .C2(n6006), .A(n6001), .B(n6008), .ZN(n6002)
         );
  AOI211_X1 U7002 ( .C1(n6004), .C2(n6050), .A(n6003), .B(n6002), .ZN(n6005)
         );
  OAI21_X1 U7003 ( .B1(n6013), .B2(n6006), .A(n6005), .ZN(U3010) );
  AOI22_X1 U7004 ( .A1(n6007), .A2(n6044), .B1(n6032), .B2(REIP_REG_7__SCAN_IN), .ZN(n6012) );
  INV_X1 U7005 ( .A(n6008), .ZN(n6009) );
  AOI22_X1 U7006 ( .A1(n6010), .A2(n6050), .B1(n6009), .B2(n6570), .ZN(n6011)
         );
  OAI211_X1 U7007 ( .C1(n6013), .C2(n6570), .A(n6012), .B(n6011), .ZN(U3011)
         );
  AOI21_X1 U7008 ( .B1(n6015), .B2(n6014), .A(INSTADDRPOINTER_REG_5__SCAN_IN), 
        .ZN(n6020) );
  AOI22_X1 U7009 ( .A1(n6017), .A2(n6050), .B1(n6044), .B2(n6016), .ZN(n6019)
         );
  NAND2_X1 U7010 ( .A1(n6032), .A2(REIP_REG_5__SCAN_IN), .ZN(n6018) );
  OAI211_X1 U7011 ( .C1(n6021), .C2(n6020), .A(n6019), .B(n6018), .ZN(U3013)
         );
  AOI21_X1 U7012 ( .B1(n6040), .B2(n6041), .A(n6049), .ZN(n6039) );
  OAI222_X1 U7013 ( .A1(n6025), .A2(n6024), .B1(n6047), .B2(n6419), .C1(n6023), 
        .C2(n6022), .ZN(n6026) );
  INV_X1 U7014 ( .A(n6026), .ZN(n6030) );
  NOR2_X1 U7015 ( .A1(n6041), .A2(n6027), .ZN(n6035) );
  OAI211_X1 U7016 ( .C1(INSTADDRPOINTER_REG_3__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .A(n6035), .B(n6028), .ZN(n6029) );
  OAI211_X1 U7017 ( .C1(n6039), .C2(n6031), .A(n6030), .B(n6029), .ZN(U3014)
         );
  AOI22_X1 U7018 ( .A1(n6044), .A2(n6033), .B1(n6032), .B2(REIP_REG_3__SCAN_IN), .ZN(n6037) );
  AOI22_X1 U7019 ( .A1(n6035), .A2(n6038), .B1(n6034), .B2(n6050), .ZN(n6036)
         );
  OAI211_X1 U7020 ( .C1(n6039), .C2(n6038), .A(n6037), .B(n6036), .ZN(U3015)
         );
  OAI221_X1 U7021 ( .B1(n6042), .B2(n6041), .C1(INSTADDRPOINTER_REG_0__SCAN_IN), .C2(n6041), .A(n6040), .ZN(n6046) );
  NAND2_X1 U7022 ( .A1(n6044), .A2(n6043), .ZN(n6045) );
  OAI211_X1 U7023 ( .C1(n6416), .C2(n6047), .A(n6046), .B(n6045), .ZN(n6048)
         );
  INV_X1 U7024 ( .A(n6048), .ZN(n6053) );
  AOI22_X1 U7025 ( .A1(n6051), .A2(n6050), .B1(INSTADDRPOINTER_REG_2__SCAN_IN), 
        .B2(n6049), .ZN(n6052) );
  OAI211_X1 U7026 ( .C1(INSTADDRPOINTER_REG_2__SCAN_IN), .C2(n6054), .A(n6053), 
        .B(n6052), .ZN(U3016) );
  NOR2_X1 U7027 ( .A1(n6056), .A2(n6055), .ZN(U3019) );
  NOR2_X1 U7028 ( .A1(n6189), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6082)
         );
  INV_X1 U7029 ( .A(n6118), .ZN(n6190) );
  AOI22_X1 U7030 ( .A1(n6284), .A2(n6082), .B1(n6291), .B2(n6081), .ZN(n6067)
         );
  INV_X1 U7031 ( .A(n6063), .ZN(n6061) );
  INV_X1 U7032 ( .A(n6057), .ZN(n6058) );
  AOI21_X1 U7033 ( .B1(n6058), .B2(n6192), .A(n6286), .ZN(n6062) );
  AOI21_X1 U7034 ( .B1(n6059), .B2(n3503), .A(n6082), .ZN(n6064) );
  NAND2_X1 U7035 ( .A1(n6062), .A2(n6064), .ZN(n6060) );
  OAI211_X1 U7036 ( .C1(n6197), .C2(n6061), .A(n6290), .B(n6060), .ZN(n6084)
         );
  INV_X1 U7037 ( .A(n6062), .ZN(n6065) );
  OAI22_X1 U7038 ( .A1(n6065), .A2(n6064), .B1(n6063), .B2(n6379), .ZN(n6083)
         );
  AOI22_X1 U7039 ( .A1(INSTQUEUE_REG_3__0__SCAN_IN), .A2(n6084), .B1(n6231), 
        .B2(n6083), .ZN(n6066) );
  OAI211_X1 U7040 ( .C1(n6244), .C2(n6087), .A(n6067), .B(n6066), .ZN(U3044)
         );
  AOI22_X1 U7041 ( .A1(n6296), .A2(n6082), .B1(n6295), .B2(n6081), .ZN(n6069)
         );
  AOI22_X1 U7042 ( .A1(INSTQUEUE_REG_3__1__SCAN_IN), .A2(n6084), .B1(n6245), 
        .B2(n6083), .ZN(n6068) );
  OAI211_X1 U7043 ( .C1(n6087), .C2(n6248), .A(n6069), .B(n6068), .ZN(U3045)
         );
  AOI22_X1 U7044 ( .A1(n6302), .A2(n6082), .B1(n6301), .B2(n6081), .ZN(n6071)
         );
  AOI22_X1 U7045 ( .A1(INSTQUEUE_REG_3__2__SCAN_IN), .A2(n6084), .B1(n6249), 
        .B2(n6083), .ZN(n6070) );
  OAI211_X1 U7046 ( .C1(n6087), .C2(n6252), .A(n6071), .B(n6070), .ZN(U3046)
         );
  AOI22_X1 U7047 ( .A1(n6308), .A2(n6082), .B1(n6307), .B2(n6072), .ZN(n6074)
         );
  AOI22_X1 U7048 ( .A1(INSTQUEUE_REG_3__3__SCAN_IN), .A2(n6084), .B1(n6253), 
        .B2(n6083), .ZN(n6073) );
  OAI211_X1 U7049 ( .C1(n6213), .C2(n6117), .A(n6074), .B(n6073), .ZN(U3047)
         );
  AOI22_X1 U7050 ( .A1(n6314), .A2(n6082), .B1(n6315), .B2(n6081), .ZN(n6076)
         );
  AOI22_X1 U7051 ( .A1(INSTQUEUE_REG_3__4__SCAN_IN), .A2(n6084), .B1(n6257), 
        .B2(n6083), .ZN(n6075) );
  OAI211_X1 U7052 ( .C1(n6087), .C2(n6260), .A(n6076), .B(n6075), .ZN(U3048)
         );
  AOI22_X1 U7053 ( .A1(n6320), .A2(n6082), .B1(n6321), .B2(n6081), .ZN(n6078)
         );
  AOI22_X1 U7054 ( .A1(INSTQUEUE_REG_3__5__SCAN_IN), .A2(n6084), .B1(n6261), 
        .B2(n6083), .ZN(n6077) );
  OAI211_X1 U7055 ( .C1(n6087), .C2(n6264), .A(n6078), .B(n6077), .ZN(U3049)
         );
  AOI22_X1 U7056 ( .A1(n6326), .A2(n6082), .B1(n6325), .B2(n6081), .ZN(n6080)
         );
  AOI22_X1 U7057 ( .A1(INSTQUEUE_REG_3__6__SCAN_IN), .A2(n6084), .B1(n6265), 
        .B2(n6083), .ZN(n6079) );
  OAI211_X1 U7058 ( .C1(n6087), .C2(n6268), .A(n6080), .B(n6079), .ZN(U3050)
         );
  AOI22_X1 U7059 ( .A1(n6334), .A2(n6082), .B1(n6336), .B2(n6081), .ZN(n6086)
         );
  AOI22_X1 U7060 ( .A1(INSTQUEUE_REG_3__7__SCAN_IN), .A2(n6084), .B1(n6271), 
        .B2(n6083), .ZN(n6085) );
  OAI211_X1 U7061 ( .C1(n6087), .C2(n6276), .A(n6086), .B(n6085), .ZN(U3051)
         );
  NAND2_X1 U7062 ( .A1(n6278), .A2(n6197), .ZN(n6230) );
  INV_X1 U7063 ( .A(n6088), .ZN(n6089) );
  OAI22_X1 U7064 ( .A1(n6230), .A2(n6237), .B1(n6089), .B2(n6227), .ZN(n6112)
         );
  NOR2_X1 U7065 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6090), .ZN(n6111)
         );
  AOI22_X1 U7066 ( .A1(n6231), .A2(n6112), .B1(n6284), .B2(n6111), .ZN(n6098)
         );
  NAND3_X1 U7067 ( .A1(n6096), .A2(n6197), .A3(n6117), .ZN(n6092) );
  AOI21_X1 U7068 ( .B1(n6092), .B2(n6163), .A(n6091), .ZN(n6095) );
  NOR2_X1 U7069 ( .A1(n6470), .A2(n6111), .ZN(n6093) );
  AOI22_X1 U7070 ( .A1(n6114), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n6291), 
        .B2(n6113), .ZN(n6097) );
  OAI211_X1 U7071 ( .C1(n6244), .C2(n6117), .A(n6098), .B(n6097), .ZN(U3052)
         );
  AOI22_X1 U7072 ( .A1(n6245), .A2(n6112), .B1(n6296), .B2(n6111), .ZN(n6100)
         );
  AOI22_X1 U7073 ( .A1(n6114), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n6295), 
        .B2(n6113), .ZN(n6099) );
  OAI211_X1 U7074 ( .C1(n6248), .C2(n6117), .A(n6100), .B(n6099), .ZN(U3053)
         );
  AOI22_X1 U7075 ( .A1(n6249), .A2(n6112), .B1(n6302), .B2(n6111), .ZN(n6102)
         );
  AOI22_X1 U7076 ( .A1(n6114), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n6301), 
        .B2(n6113), .ZN(n6101) );
  OAI211_X1 U7077 ( .C1(n6252), .C2(n6117), .A(n6102), .B(n6101), .ZN(U3054)
         );
  AOI22_X1 U7078 ( .A1(n6253), .A2(n6112), .B1(n6308), .B2(n6111), .ZN(n6104)
         );
  AOI22_X1 U7079 ( .A1(n6114), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n6309), 
        .B2(n6113), .ZN(n6103) );
  OAI211_X1 U7080 ( .C1(n6256), .C2(n6117), .A(n6104), .B(n6103), .ZN(U3055)
         );
  AOI22_X1 U7081 ( .A1(n6257), .A2(n6112), .B1(n6314), .B2(n6111), .ZN(n6106)
         );
  AOI22_X1 U7082 ( .A1(n6114), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n6315), 
        .B2(n6113), .ZN(n6105) );
  OAI211_X1 U7083 ( .C1(n6260), .C2(n6117), .A(n6106), .B(n6105), .ZN(U3056)
         );
  AOI22_X1 U7084 ( .A1(n6261), .A2(n6112), .B1(n6320), .B2(n6111), .ZN(n6108)
         );
  AOI22_X1 U7085 ( .A1(n6114), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n6321), 
        .B2(n6113), .ZN(n6107) );
  OAI211_X1 U7086 ( .C1(n6264), .C2(n6117), .A(n6108), .B(n6107), .ZN(U3057)
         );
  AOI22_X1 U7087 ( .A1(n6265), .A2(n6112), .B1(n6326), .B2(n6111), .ZN(n6110)
         );
  AOI22_X1 U7088 ( .A1(n6114), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n6325), 
        .B2(n6113), .ZN(n6109) );
  OAI211_X1 U7089 ( .C1(n6268), .C2(n6117), .A(n6110), .B(n6109), .ZN(U3058)
         );
  AOI22_X1 U7090 ( .A1(n6271), .A2(n6112), .B1(n6334), .B2(n6111), .ZN(n6116)
         );
  AOI22_X1 U7091 ( .A1(n6114), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n6336), 
        .B2(n6113), .ZN(n6115) );
  OAI211_X1 U7092 ( .C1(n6276), .C2(n6117), .A(n6116), .B(n6115), .ZN(U3059)
         );
  INV_X1 U7093 ( .A(n6122), .ZN(n6149) );
  AOI22_X1 U7094 ( .A1(n6284), .A2(n6149), .B1(n6283), .B2(n6144), .ZN(n6130)
         );
  NOR2_X1 U7095 ( .A1(n6120), .A2(n6286), .ZN(n6125) );
  OR3_X1 U7096 ( .A1(n6121), .A2(n6237), .A3(n6346), .ZN(n6123) );
  AND2_X1 U7097 ( .A1(n6123), .A2(n6122), .ZN(n6128) );
  AOI22_X1 U7098 ( .A1(n6125), .A2(n6128), .B1(n6126), .B2(n6286), .ZN(n6124)
         );
  NAND2_X1 U7099 ( .A1(n6290), .A2(n6124), .ZN(n6151) );
  INV_X1 U7100 ( .A(n6125), .ZN(n6127) );
  OAI22_X1 U7101 ( .A1(n6128), .A2(n6127), .B1(n6379), .B2(n6126), .ZN(n6150)
         );
  AOI22_X1 U7102 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n6151), .B1(n6231), 
        .B2(n6150), .ZN(n6129) );
  OAI211_X1 U7103 ( .C1(n6131), .C2(n6188), .A(n6130), .B(n6129), .ZN(U3076)
         );
  INV_X1 U7104 ( .A(n6188), .ZN(n6148) );
  AOI22_X1 U7105 ( .A1(n6296), .A2(n6149), .B1(n6295), .B2(n6148), .ZN(n6133)
         );
  AOI22_X1 U7106 ( .A1(INSTQUEUE_REG_7__1__SCAN_IN), .A2(n6151), .B1(n6245), 
        .B2(n6150), .ZN(n6132) );
  OAI211_X1 U7107 ( .C1(n6248), .C2(n6154), .A(n6133), .B(n6132), .ZN(U3077)
         );
  AOI22_X1 U7108 ( .A1(n6302), .A2(n6149), .B1(n6301), .B2(n6148), .ZN(n6135)
         );
  AOI22_X1 U7109 ( .A1(INSTQUEUE_REG_7__2__SCAN_IN), .A2(n6151), .B1(n6249), 
        .B2(n6150), .ZN(n6134) );
  OAI211_X1 U7110 ( .C1(n6252), .C2(n6154), .A(n6135), .B(n6134), .ZN(U3078)
         );
  AOI22_X1 U7111 ( .A1(n6308), .A2(n6149), .B1(n6307), .B2(n6144), .ZN(n6137)
         );
  AOI22_X1 U7112 ( .A1(INSTQUEUE_REG_7__3__SCAN_IN), .A2(n6151), .B1(n6253), 
        .B2(n6150), .ZN(n6136) );
  OAI211_X1 U7113 ( .C1(n6213), .C2(n6188), .A(n6137), .B(n6136), .ZN(U3079)
         );
  AOI22_X1 U7114 ( .A1(n6314), .A2(n6149), .B1(n6313), .B2(n6144), .ZN(n6139)
         );
  AOI22_X1 U7115 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n6151), .B1(n6257), 
        .B2(n6150), .ZN(n6138) );
  OAI211_X1 U7116 ( .C1(n6140), .C2(n6188), .A(n6139), .B(n6138), .ZN(U3080)
         );
  AOI22_X1 U7117 ( .A1(n6320), .A2(n6149), .B1(n6319), .B2(n6144), .ZN(n6142)
         );
  AOI22_X1 U7118 ( .A1(INSTQUEUE_REG_7__5__SCAN_IN), .A2(n6151), .B1(n6261), 
        .B2(n6150), .ZN(n6141) );
  OAI211_X1 U7119 ( .C1(n6143), .C2(n6188), .A(n6142), .B(n6141), .ZN(U3081)
         );
  AOI22_X1 U7120 ( .A1(n6326), .A2(n6149), .B1(n6327), .B2(n6144), .ZN(n6146)
         );
  AOI22_X1 U7121 ( .A1(INSTQUEUE_REG_7__6__SCAN_IN), .A2(n6151), .B1(n6265), 
        .B2(n6150), .ZN(n6145) );
  OAI211_X1 U7122 ( .C1(n6147), .C2(n6188), .A(n6146), .B(n6145), .ZN(U3082)
         );
  AOI22_X1 U7123 ( .A1(n6334), .A2(n6149), .B1(n6336), .B2(n6148), .ZN(n6153)
         );
  AOI22_X1 U7124 ( .A1(INSTQUEUE_REG_7__7__SCAN_IN), .A2(n6151), .B1(n6271), 
        .B2(n6150), .ZN(n6152) );
  OAI211_X1 U7125 ( .C1(n6276), .C2(n6154), .A(n6153), .B(n6152), .ZN(U3083)
         );
  NOR2_X1 U7126 ( .A1(n6229), .A2(n6155), .ZN(n6162) );
  INV_X1 U7127 ( .A(n6162), .ZN(n6159) );
  INV_X1 U7128 ( .A(n6156), .ZN(n6239) );
  NAND2_X1 U7129 ( .A1(n6158), .A2(n6157), .ZN(n6228) );
  OAI22_X1 U7130 ( .A1(n6159), .A2(n6286), .B1(n6239), .B2(n6228), .ZN(n6183)
         );
  NOR2_X1 U7131 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6160), .ZN(n6182)
         );
  AOI22_X1 U7132 ( .A1(n6231), .A2(n6183), .B1(n6284), .B2(n6182), .ZN(n6169)
         );
  INV_X1 U7133 ( .A(n6184), .ZN(n6161) );
  NAND3_X1 U7134 ( .A1(n6161), .A2(n6197), .A3(n6188), .ZN(n6164) );
  AOI21_X1 U7135 ( .B1(n6164), .B2(n6163), .A(n6162), .ZN(n6167) );
  AOI21_X1 U7136 ( .B1(n6228), .B2(STATE2_REG_2__SCAN_IN), .A(n6165), .ZN(
        n6238) );
  OAI211_X1 U7137 ( .C1(n6470), .C2(n6182), .A(n6227), .B(n6238), .ZN(n6166)
         );
  AOI22_X1 U7138 ( .A1(n6185), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n6291), 
        .B2(n6184), .ZN(n6168) );
  OAI211_X1 U7139 ( .C1(n6244), .C2(n6188), .A(n6169), .B(n6168), .ZN(U3084)
         );
  AOI22_X1 U7140 ( .A1(n6245), .A2(n6183), .B1(n6296), .B2(n6182), .ZN(n6171)
         );
  AOI22_X1 U7141 ( .A1(n6185), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n6295), 
        .B2(n6184), .ZN(n6170) );
  OAI211_X1 U7142 ( .C1(n6248), .C2(n6188), .A(n6171), .B(n6170), .ZN(U3085)
         );
  AOI22_X1 U7143 ( .A1(n6249), .A2(n6183), .B1(n6302), .B2(n6182), .ZN(n6173)
         );
  AOI22_X1 U7144 ( .A1(n6185), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n6301), 
        .B2(n6184), .ZN(n6172) );
  OAI211_X1 U7145 ( .C1(n6252), .C2(n6188), .A(n6173), .B(n6172), .ZN(U3086)
         );
  AOI22_X1 U7146 ( .A1(n6253), .A2(n6183), .B1(n6308), .B2(n6182), .ZN(n6175)
         );
  AOI22_X1 U7147 ( .A1(n6185), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n6309), 
        .B2(n6184), .ZN(n6174) );
  OAI211_X1 U7148 ( .C1(n6256), .C2(n6188), .A(n6175), .B(n6174), .ZN(U3087)
         );
  AOI22_X1 U7149 ( .A1(n6257), .A2(n6183), .B1(n6314), .B2(n6182), .ZN(n6177)
         );
  AOI22_X1 U7150 ( .A1(n6185), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n6315), 
        .B2(n6184), .ZN(n6176) );
  OAI211_X1 U7151 ( .C1(n6260), .C2(n6188), .A(n6177), .B(n6176), .ZN(U3088)
         );
  AOI22_X1 U7152 ( .A1(n6261), .A2(n6183), .B1(n6320), .B2(n6182), .ZN(n6179)
         );
  AOI22_X1 U7153 ( .A1(n6185), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n6321), 
        .B2(n6184), .ZN(n6178) );
  OAI211_X1 U7154 ( .C1(n6264), .C2(n6188), .A(n6179), .B(n6178), .ZN(U3089)
         );
  AOI22_X1 U7155 ( .A1(n6265), .A2(n6183), .B1(n6326), .B2(n6182), .ZN(n6181)
         );
  AOI22_X1 U7156 ( .A1(n6185), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n6325), 
        .B2(n6184), .ZN(n6180) );
  OAI211_X1 U7157 ( .C1(n6268), .C2(n6188), .A(n6181), .B(n6180), .ZN(U3090)
         );
  AOI22_X1 U7158 ( .A1(n6271), .A2(n6183), .B1(n6334), .B2(n6182), .ZN(n6187)
         );
  AOI22_X1 U7159 ( .A1(n6185), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n6336), 
        .B2(n6184), .ZN(n6186) );
  OAI211_X1 U7160 ( .C1(n6276), .C2(n6188), .A(n6187), .B(n6186), .ZN(U3091)
         );
  NOR2_X1 U7161 ( .A1(n6189), .A2(n6358), .ZN(n6221) );
  INV_X1 U7162 ( .A(n6275), .ZN(n6220) );
  AOI22_X1 U7163 ( .A1(n6284), .A2(n6221), .B1(n6291), .B2(n6220), .ZN(n6203)
         );
  INV_X1 U7164 ( .A(n6199), .ZN(n6196) );
  AOI21_X1 U7165 ( .B1(n6193), .B2(n6192), .A(n6286), .ZN(n6198) );
  AOI21_X1 U7166 ( .B1(n6194), .B2(n3503), .A(n6221), .ZN(n6200) );
  NAND2_X1 U7167 ( .A1(n6198), .A2(n6200), .ZN(n6195) );
  OAI211_X1 U7168 ( .C1(n6197), .C2(n6196), .A(n6290), .B(n6195), .ZN(n6223)
         );
  INV_X1 U7169 ( .A(n6198), .ZN(n6201) );
  OAI22_X1 U7170 ( .A1(n6201), .A2(n6200), .B1(n6199), .B2(n6379), .ZN(n6222)
         );
  AOI22_X1 U7171 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n6223), .B1(n6231), 
        .B2(n6222), .ZN(n6202) );
  OAI211_X1 U7172 ( .C1(n6244), .C2(n6226), .A(n6203), .B(n6202), .ZN(U3108)
         );
  INV_X1 U7173 ( .A(n6226), .ZN(n6210) );
  AOI22_X1 U7174 ( .A1(n6296), .A2(n6221), .B1(n6210), .B2(n6297), .ZN(n6205)
         );
  AOI22_X1 U7175 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(n6223), .B1(n6245), 
        .B2(n6222), .ZN(n6204) );
  OAI211_X1 U7176 ( .C1(n6206), .C2(n6275), .A(n6205), .B(n6204), .ZN(U3109)
         );
  AOI22_X1 U7177 ( .A1(n6302), .A2(n6221), .B1(n6210), .B2(n6303), .ZN(n6208)
         );
  AOI22_X1 U7178 ( .A1(INSTQUEUE_REG_11__2__SCAN_IN), .A2(n6223), .B1(n6249), 
        .B2(n6222), .ZN(n6207) );
  OAI211_X1 U7179 ( .C1(n6209), .C2(n6275), .A(n6208), .B(n6207), .ZN(U3110)
         );
  AOI22_X1 U7180 ( .A1(n6308), .A2(n6221), .B1(n6210), .B2(n6307), .ZN(n6212)
         );
  AOI22_X1 U7181 ( .A1(INSTQUEUE_REG_11__3__SCAN_IN), .A2(n6223), .B1(n6253), 
        .B2(n6222), .ZN(n6211) );
  OAI211_X1 U7182 ( .C1(n6213), .C2(n6275), .A(n6212), .B(n6211), .ZN(U3111)
         );
  AOI22_X1 U7183 ( .A1(n6314), .A2(n6221), .B1(n6315), .B2(n6220), .ZN(n6215)
         );
  AOI22_X1 U7184 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n6223), .B1(n6257), 
        .B2(n6222), .ZN(n6214) );
  OAI211_X1 U7185 ( .C1(n6260), .C2(n6226), .A(n6215), .B(n6214), .ZN(U3112)
         );
  AOI22_X1 U7186 ( .A1(n6320), .A2(n6221), .B1(n6321), .B2(n6220), .ZN(n6217)
         );
  AOI22_X1 U7187 ( .A1(INSTQUEUE_REG_11__5__SCAN_IN), .A2(n6223), .B1(n6261), 
        .B2(n6222), .ZN(n6216) );
  OAI211_X1 U7188 ( .C1(n6264), .C2(n6226), .A(n6217), .B(n6216), .ZN(U3113)
         );
  AOI22_X1 U7189 ( .A1(n6326), .A2(n6221), .B1(n6325), .B2(n6220), .ZN(n6219)
         );
  AOI22_X1 U7190 ( .A1(INSTQUEUE_REG_11__6__SCAN_IN), .A2(n6223), .B1(n6265), 
        .B2(n6222), .ZN(n6218) );
  OAI211_X1 U7191 ( .C1(n6268), .C2(n6226), .A(n6219), .B(n6218), .ZN(U3114)
         );
  AOI22_X1 U7192 ( .A1(n6334), .A2(n6221), .B1(n6336), .B2(n6220), .ZN(n6225)
         );
  AOI22_X1 U7193 ( .A1(INSTQUEUE_REG_11__7__SCAN_IN), .A2(n6223), .B1(n6271), 
        .B2(n6222), .ZN(n6224) );
  OAI211_X1 U7194 ( .C1(n6276), .C2(n6226), .A(n6225), .B(n6224), .ZN(U3115)
         );
  OAI22_X1 U7195 ( .A1(n6230), .A2(n6229), .B1(n6228), .B2(n6227), .ZN(n6270)
         );
  NAND2_X1 U7196 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6282), .ZN(n6285) );
  NOR2_X1 U7197 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6285), .ZN(n6269)
         );
  AOI22_X1 U7198 ( .A1(n6231), .A2(n6270), .B1(n6284), .B2(n6269), .ZN(n6243)
         );
  NOR2_X2 U7199 ( .A1(n6233), .A2(n6232), .ZN(n6332) );
  INV_X1 U7200 ( .A(n6332), .ZN(n6235) );
  AOI21_X1 U7201 ( .B1(n6235), .B2(n6275), .A(n6234), .ZN(n6236) );
  AOI211_X1 U7202 ( .C1(n6278), .C2(n6237), .A(n6286), .B(n6236), .ZN(n6241)
         );
  OAI211_X1 U7203 ( .C1(n6470), .C2(n6269), .A(n6239), .B(n6238), .ZN(n6240)
         );
  AOI22_X1 U7204 ( .A1(n6272), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n6291), 
        .B2(n6332), .ZN(n6242) );
  OAI211_X1 U7205 ( .C1(n6244), .C2(n6275), .A(n6243), .B(n6242), .ZN(U3116)
         );
  AOI22_X1 U7206 ( .A1(n6245), .A2(n6270), .B1(n6296), .B2(n6269), .ZN(n6247)
         );
  AOI22_X1 U7207 ( .A1(n6272), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n6295), 
        .B2(n6332), .ZN(n6246) );
  OAI211_X1 U7208 ( .C1(n6248), .C2(n6275), .A(n6247), .B(n6246), .ZN(U3117)
         );
  AOI22_X1 U7209 ( .A1(n6249), .A2(n6270), .B1(n6302), .B2(n6269), .ZN(n6251)
         );
  AOI22_X1 U7210 ( .A1(n6272), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n6301), 
        .B2(n6332), .ZN(n6250) );
  OAI211_X1 U7211 ( .C1(n6252), .C2(n6275), .A(n6251), .B(n6250), .ZN(U3118)
         );
  AOI22_X1 U7212 ( .A1(n6253), .A2(n6270), .B1(n6308), .B2(n6269), .ZN(n6255)
         );
  AOI22_X1 U7213 ( .A1(n6272), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n6309), 
        .B2(n6332), .ZN(n6254) );
  OAI211_X1 U7214 ( .C1(n6256), .C2(n6275), .A(n6255), .B(n6254), .ZN(U3119)
         );
  AOI22_X1 U7215 ( .A1(n6257), .A2(n6270), .B1(n6314), .B2(n6269), .ZN(n6259)
         );
  AOI22_X1 U7216 ( .A1(n6272), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n6315), 
        .B2(n6332), .ZN(n6258) );
  OAI211_X1 U7217 ( .C1(n6260), .C2(n6275), .A(n6259), .B(n6258), .ZN(U3120)
         );
  AOI22_X1 U7218 ( .A1(n6261), .A2(n6270), .B1(n6320), .B2(n6269), .ZN(n6263)
         );
  AOI22_X1 U7219 ( .A1(n6272), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n6321), 
        .B2(n6332), .ZN(n6262) );
  OAI211_X1 U7220 ( .C1(n6264), .C2(n6275), .A(n6263), .B(n6262), .ZN(U3121)
         );
  AOI22_X1 U7221 ( .A1(n6265), .A2(n6270), .B1(n6326), .B2(n6269), .ZN(n6267)
         );
  AOI22_X1 U7222 ( .A1(n6272), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n6325), 
        .B2(n6332), .ZN(n6266) );
  OAI211_X1 U7223 ( .C1(n6268), .C2(n6275), .A(n6267), .B(n6266), .ZN(U3122)
         );
  AOI22_X1 U7224 ( .A1(n6271), .A2(n6270), .B1(n6334), .B2(n6269), .ZN(n6274)
         );
  AOI22_X1 U7225 ( .A1(n6272), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n6336), 
        .B2(n6332), .ZN(n6273) );
  OAI211_X1 U7226 ( .C1(n6276), .C2(n6275), .A(n6274), .B(n6273), .ZN(U3123)
         );
  NOR2_X1 U7227 ( .A1(n6379), .A2(n6358), .ZN(n6281) );
  NOR2_X1 U7228 ( .A1(n6277), .A2(n6286), .ZN(n6288) );
  NOR2_X1 U7229 ( .A1(n6635), .A2(n6285), .ZN(n6333) );
  AOI21_X1 U7230 ( .B1(n6279), .B2(n6278), .A(n6333), .ZN(n6287) );
  INV_X1 U7231 ( .A(n6287), .ZN(n6280) );
  AOI22_X1 U7232 ( .A1(n6282), .A2(n6281), .B1(n6288), .B2(n6280), .ZN(n6341)
         );
  AOI22_X1 U7233 ( .A1(n6284), .A2(n6333), .B1(n6332), .B2(n6283), .ZN(n6293)
         );
  AOI22_X1 U7234 ( .A1(n6288), .A2(n6287), .B1(n6286), .B2(n6285), .ZN(n6289)
         );
  NAND2_X1 U7235 ( .A1(n6290), .A2(n6289), .ZN(n6337) );
  AOI22_X1 U7236 ( .A1(n6337), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n6291), 
        .B2(n6335), .ZN(n6292) );
  OAI211_X1 U7237 ( .C1(n6341), .C2(n6294), .A(n6293), .B(n6292), .ZN(U3124)
         );
  AOI22_X1 U7238 ( .A1(n6296), .A2(n6333), .B1(n6335), .B2(n6295), .ZN(n6299)
         );
  AOI22_X1 U7239 ( .A1(n6337), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n6297), 
        .B2(n6332), .ZN(n6298) );
  OAI211_X1 U7240 ( .C1(n6341), .C2(n6300), .A(n6299), .B(n6298), .ZN(U3125)
         );
  AOI22_X1 U7241 ( .A1(n6302), .A2(n6333), .B1(n6335), .B2(n6301), .ZN(n6305)
         );
  AOI22_X1 U7242 ( .A1(n6337), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n6303), 
        .B2(n6332), .ZN(n6304) );
  OAI211_X1 U7243 ( .C1(n6341), .C2(n6306), .A(n6305), .B(n6304), .ZN(U3126)
         );
  AOI22_X1 U7244 ( .A1(n6308), .A2(n6333), .B1(n6332), .B2(n6307), .ZN(n6311)
         );
  AOI22_X1 U7245 ( .A1(n6337), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n6309), 
        .B2(n6335), .ZN(n6310) );
  OAI211_X1 U7246 ( .C1(n6341), .C2(n6312), .A(n6311), .B(n6310), .ZN(U3127)
         );
  AOI22_X1 U7247 ( .A1(n6314), .A2(n6333), .B1(n6332), .B2(n6313), .ZN(n6317)
         );
  AOI22_X1 U7248 ( .A1(n6337), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n6315), 
        .B2(n6335), .ZN(n6316) );
  OAI211_X1 U7249 ( .C1(n6341), .C2(n6318), .A(n6317), .B(n6316), .ZN(U3128)
         );
  AOI22_X1 U7250 ( .A1(n6320), .A2(n6333), .B1(n6332), .B2(n6319), .ZN(n6323)
         );
  AOI22_X1 U7251 ( .A1(n6337), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n6321), 
        .B2(n6335), .ZN(n6322) );
  OAI211_X1 U7252 ( .C1(n6341), .C2(n6324), .A(n6323), .B(n6322), .ZN(U3129)
         );
  AOI22_X1 U7253 ( .A1(n6326), .A2(n6333), .B1(n6335), .B2(n6325), .ZN(n6329)
         );
  AOI22_X1 U7254 ( .A1(n6337), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n6327), 
        .B2(n6332), .ZN(n6328) );
  OAI211_X1 U7255 ( .C1(n6341), .C2(n6330), .A(n6329), .B(n6328), .ZN(U3130)
         );
  AOI22_X1 U7256 ( .A1(n6334), .A2(n6333), .B1(n6332), .B2(n6331), .ZN(n6339)
         );
  AOI22_X1 U7257 ( .A1(n6337), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n6336), 
        .B2(n6335), .ZN(n6338) );
  OAI211_X1 U7258 ( .C1(n6341), .C2(n6340), .A(n6339), .B(n6338), .ZN(U3131)
         );
  AND2_X1 U7259 ( .A1(n6349), .A2(n6342), .ZN(n6359) );
  NAND2_X1 U7260 ( .A1(n6349), .A2(n5151), .ZN(n6356) );
  INV_X1 U7261 ( .A(n6344), .ZN(n6345) );
  OAI22_X1 U7262 ( .A1(n6346), .A2(n6345), .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n3684), .ZN(n6471) );
  NAND2_X1 U7263 ( .A1(n6347), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n6480) );
  INV_X1 U7264 ( .A(n6480), .ZN(n6348) );
  NOR3_X1 U7265 ( .A1(n6471), .A2(n6348), .A3(n6635), .ZN(n6352) );
  NAND2_X1 U7266 ( .A1(n6352), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6354) );
  INV_X1 U7267 ( .A(n6349), .ZN(n6351) );
  OAI22_X1 U7268 ( .A1(n6352), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B1(n6351), .B2(n6350), .ZN(n6353) );
  NAND2_X1 U7269 ( .A1(n6354), .A2(n6353), .ZN(n6355) );
  AOI222_X1 U7270 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n6356), .B1(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n6355), .C1(n6356), .C2(n6355), 
        .ZN(n6357) );
  AOI222_X1 U7271 ( .A1(n6359), .A2(n6358), .B1(n6359), .B2(n6357), .C1(n6358), 
        .C2(n6357), .ZN(n6362) );
  OAI21_X1 U7272 ( .B1(FLUSH_REG_SCAN_IN), .B2(MORE_REG_SCAN_IN), .A(n6360), 
        .ZN(n6361) );
  OAI21_X1 U7273 ( .B1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(n6362), .A(n6361), 
        .ZN(n6367) );
  NAND3_X1 U7274 ( .A1(n6365), .A2(n6364), .A3(n6363), .ZN(n6366) );
  OR2_X1 U7275 ( .A1(n6367), .A2(n6366), .ZN(n6378) );
  OAI22_X1 U7276 ( .A1(n6378), .A2(n6369), .B1(n6492), .B2(n6368), .ZN(n6375)
         );
  INV_X1 U7277 ( .A(n6370), .ZN(n6373) );
  INV_X1 U7278 ( .A(n6371), .ZN(n6372) );
  NAND2_X1 U7279 ( .A1(n6373), .A2(n6372), .ZN(n6374) );
  AOI211_X1 U7280 ( .C1(n6497), .C2(n6472), .A(STATE2_REG_0__SCAN_IN), .B(
        n6467), .ZN(n6376) );
  AOI211_X1 U7281 ( .C1(n6383), .C2(n6378), .A(n6377), .B(n6376), .ZN(n6380)
         );
  OAI221_X1 U7282 ( .B1(n6467), .B2(READY_N), .C1(n6467), .C2(n6379), .A(
        STATE2_REG_0__SCAN_IN), .ZN(n6390) );
  OAI211_X1 U7283 ( .C1(n6382), .C2(n6381), .A(n6380), .B(n6390), .ZN(U3148)
         );
  NOR2_X1 U7284 ( .A1(READY_N), .A2(n6382), .ZN(n6393) );
  AOI21_X1 U7285 ( .B1(n6384), .B2(n6393), .A(n6383), .ZN(n6385) );
  NOR2_X1 U7286 ( .A1(n6385), .A2(n6467), .ZN(n6386) );
  AOI211_X1 U7287 ( .C1(n6467), .C2(n6388), .A(n6387), .B(n6386), .ZN(n6389)
         );
  OAI21_X1 U7288 ( .B1(n6391), .B2(n6390), .A(n6389), .ZN(U3149) );
  OAI211_X1 U7289 ( .C1(STATE2_REG_2__SCAN_IN), .C2(n6393), .A(n6468), .B(
        n6392), .ZN(n6394) );
  NAND2_X1 U7290 ( .A1(n6395), .A2(n6394), .ZN(U3150) );
  INV_X1 U7291 ( .A(n6466), .ZN(n6396) );
  AND2_X1 U7292 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(n6396), .ZN(U3151) );
  AND2_X1 U7293 ( .A1(DATAWIDTH_REG_30__SCAN_IN), .A2(n6396), .ZN(U3152) );
  AND2_X1 U7294 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(n6396), .ZN(U3153) );
  AND2_X1 U7295 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(n6396), .ZN(U3154) );
  AND2_X1 U7296 ( .A1(n6396), .A2(DATAWIDTH_REG_27__SCAN_IN), .ZN(U3155) );
  AND2_X1 U7297 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(n6396), .ZN(U3156) );
  AND2_X1 U7298 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(n6396), .ZN(U3157) );
  AND2_X1 U7299 ( .A1(n6396), .A2(DATAWIDTH_REG_24__SCAN_IN), .ZN(U3158) );
  AND2_X1 U7300 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(n6396), .ZN(U3159) );
  AND2_X1 U7301 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(n6396), .ZN(U3160) );
  AND2_X1 U7302 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(n6396), .ZN(U3161) );
  AND2_X1 U7303 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(n6396), .ZN(U3162) );
  AND2_X1 U7304 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(n6396), .ZN(U3163) );
  AND2_X1 U7305 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(n6396), .ZN(U3164) );
  AND2_X1 U7306 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(n6396), .ZN(U3165) );
  AND2_X1 U7307 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(n6396), .ZN(U3166) );
  AND2_X1 U7308 ( .A1(DATAWIDTH_REG_15__SCAN_IN), .A2(n6396), .ZN(U3167) );
  AND2_X1 U7309 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(n6396), .ZN(U3168) );
  AND2_X1 U7310 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(n6396), .ZN(U3169) );
  AND2_X1 U7311 ( .A1(n6396), .A2(DATAWIDTH_REG_12__SCAN_IN), .ZN(U3170) );
  AND2_X1 U7312 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(n6396), .ZN(U3171) );
  AND2_X1 U7313 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(n6396), .ZN(U3172) );
  AND2_X1 U7314 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(n6396), .ZN(U3173) );
  AND2_X1 U7315 ( .A1(n6396), .A2(DATAWIDTH_REG_8__SCAN_IN), .ZN(U3174) );
  AND2_X1 U7316 ( .A1(DATAWIDTH_REG_7__SCAN_IN), .A2(n6396), .ZN(U3175) );
  AND2_X1 U7317 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(n6396), .ZN(U3176) );
  AND2_X1 U7318 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(n6396), .ZN(U3177) );
  AND2_X1 U7319 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(n6396), .ZN(U3178) );
  AND2_X1 U7320 ( .A1(n6396), .A2(DATAWIDTH_REG_3__SCAN_IN), .ZN(U3179) );
  AND2_X1 U7321 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(n6396), .ZN(U3180) );
  AOI22_X1 U7322 ( .A1(READY_N), .A2(STATE_REG_1__SCAN_IN), .B1(
        STATE_REG_2__SCAN_IN), .B2(HOLD), .ZN(n6413) );
  AND2_X1 U7323 ( .A1(STATE_REG_1__SCAN_IN), .A2(HOLD), .ZN(n6400) );
  INV_X1 U7324 ( .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6399) );
  OAI21_X1 U7325 ( .B1(n6400), .B2(n6399), .A(n6502), .ZN(n6397) );
  INV_X1 U7326 ( .A(n6398), .ZN(n6412) );
  OAI211_X1 U7327 ( .C1(NA_N), .C2(n6584), .A(n4130), .B(n6412), .ZN(n6410) );
  OAI211_X1 U7328 ( .C1(n6398), .C2(n6413), .A(n6397), .B(n6410), .ZN(U3181)
         );
  NOR2_X1 U7329 ( .A1(n4130), .A2(n6399), .ZN(n6406) );
  NAND2_X1 U7330 ( .A1(STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n6404) );
  OAI21_X1 U7331 ( .B1(n6406), .B2(n6400), .A(n6404), .ZN(n6401) );
  OAI211_X1 U7332 ( .C1(n6572), .C2(n6492), .A(n6402), .B(n6401), .ZN(U3182)
         );
  NOR2_X1 U7333 ( .A1(NA_N), .A2(n6492), .ZN(n6403) );
  OAI21_X1 U7334 ( .B1(n6403), .B2(n6572), .A(HOLD), .ZN(n6405) );
  OAI211_X1 U7335 ( .C1(REQUESTPENDING_REG_SCAN_IN), .C2(n6405), .A(
        STATE_REG_0__SCAN_IN), .B(n6404), .ZN(n6409) );
  INV_X1 U7336 ( .A(n6406), .ZN(n6407) );
  NOR4_X1 U7337 ( .A1(NA_N), .A2(n6572), .A3(n6492), .A4(n6407), .ZN(n6408) );
  AOI21_X1 U7338 ( .B1(n6410), .B2(n6409), .A(n6408), .ZN(n6411) );
  OAI21_X1 U7339 ( .B1(n6413), .B2(n6412), .A(n6411), .ZN(U3183) );
  NOR2_X2 U7340 ( .A1(n6584), .A2(n6502), .ZN(n6459) );
  INV_X1 U7341 ( .A(n6459), .ZN(n6457) );
  NAND2_X1 U7342 ( .A1(n6584), .A2(n5766), .ZN(n6461) );
  INV_X1 U7343 ( .A(n6461), .ZN(n6455) );
  AOI22_X1 U7344 ( .A1(REIP_REG_2__SCAN_IN), .A2(n6455), .B1(
        ADDRESS_REG_0__SCAN_IN), .B2(n6489), .ZN(n6414) );
  OAI21_X1 U7345 ( .B1(n6580), .B2(n6457), .A(n6414), .ZN(U3184) );
  AOI22_X1 U7346 ( .A1(REIP_REG_3__SCAN_IN), .A2(n6455), .B1(
        ADDRESS_REG_1__SCAN_IN), .B2(n6502), .ZN(n6415) );
  OAI21_X1 U7347 ( .B1(n6416), .B2(n6457), .A(n6415), .ZN(U3185) );
  AOI22_X1 U7348 ( .A1(REIP_REG_4__SCAN_IN), .A2(n6455), .B1(
        ADDRESS_REG_2__SCAN_IN), .B2(n6489), .ZN(n6417) );
  OAI21_X1 U7349 ( .B1(n6590), .B2(n6457), .A(n6417), .ZN(U3186) );
  AOI22_X1 U7350 ( .A1(REIP_REG_5__SCAN_IN), .A2(n6455), .B1(
        ADDRESS_REG_3__SCAN_IN), .B2(n6502), .ZN(n6418) );
  OAI21_X1 U7351 ( .B1(n6419), .B2(n6457), .A(n6418), .ZN(U3187) );
  AOI22_X1 U7352 ( .A1(REIP_REG_6__SCAN_IN), .A2(n6455), .B1(
        ADDRESS_REG_4__SCAN_IN), .B2(n6489), .ZN(n6420) );
  OAI21_X1 U7353 ( .B1(n6421), .B2(n6457), .A(n6420), .ZN(U3188) );
  AOI22_X1 U7354 ( .A1(REIP_REG_7__SCAN_IN), .A2(n6455), .B1(
        ADDRESS_REG_5__SCAN_IN), .B2(n6489), .ZN(n6422) );
  OAI21_X1 U7355 ( .B1(n4981), .B2(n6457), .A(n6422), .ZN(U3189) );
  AOI22_X1 U7356 ( .A1(REIP_REG_7__SCAN_IN), .A2(n6459), .B1(
        ADDRESS_REG_6__SCAN_IN), .B2(n6489), .ZN(n6423) );
  OAI21_X1 U7357 ( .B1(n6424), .B2(n6461), .A(n6423), .ZN(U3190) );
  AOI22_X1 U7358 ( .A1(REIP_REG_8__SCAN_IN), .A2(n6459), .B1(
        ADDRESS_REG_7__SCAN_IN), .B2(n6489), .ZN(n6425) );
  OAI21_X1 U7359 ( .B1(n4914), .B2(n6461), .A(n6425), .ZN(U3191) );
  AOI22_X1 U7360 ( .A1(REIP_REG_9__SCAN_IN), .A2(n6459), .B1(
        ADDRESS_REG_8__SCAN_IN), .B2(n6489), .ZN(n6426) );
  OAI21_X1 U7361 ( .B1(n6427), .B2(n6461), .A(n6426), .ZN(U3192) );
  AOI22_X1 U7362 ( .A1(REIP_REG_10__SCAN_IN), .A2(n6459), .B1(
        ADDRESS_REG_9__SCAN_IN), .B2(n6489), .ZN(n6428) );
  OAI21_X1 U7363 ( .B1(n4967), .B2(n6461), .A(n6428), .ZN(U3193) );
  AOI22_X1 U7364 ( .A1(REIP_REG_12__SCAN_IN), .A2(n6455), .B1(
        ADDRESS_REG_10__SCAN_IN), .B2(n6489), .ZN(n6429) );
  OAI21_X1 U7365 ( .B1(n4967), .B2(n6457), .A(n6429), .ZN(U3194) );
  AOI22_X1 U7366 ( .A1(REIP_REG_13__SCAN_IN), .A2(n6455), .B1(
        ADDRESS_REG_11__SCAN_IN), .B2(n6502), .ZN(n6430) );
  OAI21_X1 U7367 ( .B1(n6431), .B2(n6457), .A(n6430), .ZN(U3195) );
  AOI22_X1 U7368 ( .A1(REIP_REG_14__SCAN_IN), .A2(n6455), .B1(
        ADDRESS_REG_12__SCAN_IN), .B2(n6489), .ZN(n6432) );
  OAI21_X1 U7369 ( .B1(n6433), .B2(n6457), .A(n6432), .ZN(U3196) );
  AOI22_X1 U7370 ( .A1(REIP_REG_14__SCAN_IN), .A2(n6459), .B1(
        ADDRESS_REG_13__SCAN_IN), .B2(n6489), .ZN(n6434) );
  OAI21_X1 U7371 ( .B1(n6436), .B2(n6461), .A(n6434), .ZN(U3197) );
  AOI22_X1 U7372 ( .A1(REIP_REG_16__SCAN_IN), .A2(n6455), .B1(
        ADDRESS_REG_14__SCAN_IN), .B2(n6489), .ZN(n6435) );
  OAI21_X1 U7373 ( .B1(n6436), .B2(n6457), .A(n6435), .ZN(U3198) );
  AOI22_X1 U7374 ( .A1(REIP_REG_17__SCAN_IN), .A2(n6455), .B1(
        ADDRESS_REG_15__SCAN_IN), .B2(n6502), .ZN(n6437) );
  OAI21_X1 U7375 ( .B1(n6438), .B2(n6457), .A(n6437), .ZN(U3199) );
  AOI22_X1 U7376 ( .A1(REIP_REG_17__SCAN_IN), .A2(n6459), .B1(
        ADDRESS_REG_16__SCAN_IN), .B2(n6489), .ZN(n6439) );
  OAI21_X1 U7377 ( .B1(n6543), .B2(n6461), .A(n6439), .ZN(U3200) );
  AOI22_X1 U7378 ( .A1(REIP_REG_18__SCAN_IN), .A2(n6459), .B1(
        ADDRESS_REG_17__SCAN_IN), .B2(n6502), .ZN(n6440) );
  OAI21_X1 U7379 ( .B1(n6441), .B2(n6461), .A(n6440), .ZN(U3201) );
  AOI22_X1 U7380 ( .A1(REIP_REG_19__SCAN_IN), .A2(n6459), .B1(
        ADDRESS_REG_18__SCAN_IN), .B2(n6489), .ZN(n6442) );
  OAI21_X1 U7381 ( .B1(n6632), .B2(n6461), .A(n6442), .ZN(U3202) );
  AOI22_X1 U7382 ( .A1(REIP_REG_21__SCAN_IN), .A2(n6455), .B1(
        ADDRESS_REG_19__SCAN_IN), .B2(n6489), .ZN(n6443) );
  OAI21_X1 U7383 ( .B1(n6632), .B2(n6457), .A(n6443), .ZN(U3203) );
  AOI22_X1 U7384 ( .A1(REIP_REG_22__SCAN_IN), .A2(n6455), .B1(
        ADDRESS_REG_20__SCAN_IN), .B2(n6489), .ZN(n6444) );
  OAI21_X1 U7385 ( .B1(n5506), .B2(n6457), .A(n6444), .ZN(U3204) );
  AOI22_X1 U7386 ( .A1(REIP_REG_22__SCAN_IN), .A2(n6459), .B1(
        ADDRESS_REG_21__SCAN_IN), .B2(n6489), .ZN(n6445) );
  OAI21_X1 U7387 ( .B1(n6446), .B2(n6461), .A(n6445), .ZN(U3205) );
  AOI22_X1 U7388 ( .A1(REIP_REG_23__SCAN_IN), .A2(n6459), .B1(
        ADDRESS_REG_22__SCAN_IN), .B2(n6502), .ZN(n6447) );
  OAI21_X1 U7389 ( .B1(n6449), .B2(n6461), .A(n6447), .ZN(U3206) );
  AOI22_X1 U7390 ( .A1(REIP_REG_25__SCAN_IN), .A2(n6455), .B1(
        ADDRESS_REG_23__SCAN_IN), .B2(n6502), .ZN(n6448) );
  OAI21_X1 U7391 ( .B1(n6449), .B2(n6457), .A(n6448), .ZN(U3207) );
  AOI22_X1 U7392 ( .A1(REIP_REG_25__SCAN_IN), .A2(n6459), .B1(
        ADDRESS_REG_24__SCAN_IN), .B2(n6502), .ZN(n6450) );
  OAI21_X1 U7393 ( .B1(n6451), .B2(n6461), .A(n6450), .ZN(U3208) );
  AOI22_X1 U7394 ( .A1(REIP_REG_26__SCAN_IN), .A2(n6459), .B1(
        ADDRESS_REG_25__SCAN_IN), .B2(n6502), .ZN(n6452) );
  OAI21_X1 U7395 ( .B1(n6620), .B2(n6461), .A(n6452), .ZN(U3209) );
  AOI22_X1 U7396 ( .A1(REIP_REG_28__SCAN_IN), .A2(n6455), .B1(
        ADDRESS_REG_26__SCAN_IN), .B2(n6502), .ZN(n6453) );
  OAI21_X1 U7397 ( .B1(n6620), .B2(n6457), .A(n6453), .ZN(U3210) );
  AOI222_X1 U7398 ( .A1(n6459), .A2(REIP_REG_28__SCAN_IN), .B1(
        ADDRESS_REG_27__SCAN_IN), .B2(n6502), .C1(REIP_REG_29__SCAN_IN), .C2(
        n6455), .ZN(n6454) );
  INV_X1 U7399 ( .A(n6454), .ZN(U3211) );
  AOI22_X1 U7400 ( .A1(REIP_REG_30__SCAN_IN), .A2(n6455), .B1(
        ADDRESS_REG_28__SCAN_IN), .B2(n6502), .ZN(n6456) );
  OAI21_X1 U7401 ( .B1(n6458), .B2(n6457), .A(n6456), .ZN(U3212) );
  AOI22_X1 U7402 ( .A1(REIP_REG_30__SCAN_IN), .A2(n6459), .B1(
        ADDRESS_REG_29__SCAN_IN), .B2(n6502), .ZN(n6460) );
  OAI21_X1 U7403 ( .B1(n6462), .B2(n6461), .A(n6460), .ZN(U3213) );
  MUX2_X1 U7404 ( .A(BYTEENABLE_REG_3__SCAN_IN), .B(BE_N_REG_3__SCAN_IN), .S(
        n6502), .Z(U3445) );
  MUX2_X1 U7405 ( .A(BYTEENABLE_REG_2__SCAN_IN), .B(BE_N_REG_2__SCAN_IN), .S(
        n6502), .Z(U3446) );
  MUX2_X1 U7406 ( .A(BYTEENABLE_REG_1__SCAN_IN), .B(BE_N_REG_1__SCAN_IN), .S(
        n6502), .Z(U3447) );
  MUX2_X1 U7407 ( .A(BYTEENABLE_REG_0__SCAN_IN), .B(BE_N_REG_0__SCAN_IN), .S(
        n6502), .Z(U3448) );
  OAI21_X1 U7408 ( .B1(DATAWIDTH_REG_0__SCAN_IN), .B2(n6466), .A(n6464), .ZN(
        n6463) );
  INV_X1 U7409 ( .A(n6463), .ZN(U3451) );
  OAI21_X1 U7410 ( .B1(n6466), .B2(n6465), .A(n6464), .ZN(U3452) );
  INV_X1 U7411 ( .A(n6467), .ZN(n6469) );
  OAI221_X1 U7412 ( .B1(n6470), .B2(STATE2_REG_0__SCAN_IN), .C1(n6470), .C2(
        n6469), .A(n6468), .ZN(U3453) );
  AOI21_X1 U7413 ( .B1(n6471), .B2(n6470), .A(STATE2_REG_1__SCAN_IN), .ZN(
        n6474) );
  NAND2_X1 U7414 ( .A1(n6472), .A2(n3117), .ZN(n6473) );
  OAI211_X1 U7415 ( .C1(n6475), .C2(n6474), .A(n6477), .B(n6473), .ZN(n6476)
         );
  OAI21_X1 U7416 ( .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n6477), .A(n6476), 
        .ZN(n6478) );
  OAI21_X1 U7417 ( .B1(n6480), .B2(n6479), .A(n6478), .ZN(U3461) );
  AOI21_X1 U7418 ( .B1(REIP_REG_0__SCAN_IN), .B2(DATAWIDTH_REG_0__SCAN_IN), 
        .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6481) );
  OAI22_X1 U7419 ( .A1(REIP_REG_0__SCAN_IN), .A2(n6580), .B1(
        REIP_REG_1__SCAN_IN), .B2(n6481), .ZN(n6483) );
  INV_X1 U7420 ( .A(BYTEENABLE_REG_2__SCAN_IN), .ZN(n6482) );
  AOI22_X1 U7421 ( .A1(n6487), .A2(n6483), .B1(n6482), .B2(n6484), .ZN(U3468)
         );
  NOR2_X1 U7422 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_0__SCAN_IN), .ZN(
        n6486) );
  INV_X1 U7423 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n6485) );
  AOI22_X1 U7424 ( .A1(n6487), .A2(n6486), .B1(n6485), .B2(n6484), .ZN(U3469)
         );
  NAND2_X1 U7425 ( .A1(n6489), .A2(W_R_N_REG_SCAN_IN), .ZN(n6488) );
  OAI21_X1 U7426 ( .B1(n6489), .B2(READREQUEST_REG_SCAN_IN), .A(n6488), .ZN(
        U3470) );
  AOI211_X1 U7427 ( .C1(n6493), .C2(n6492), .A(n6491), .B(n6490), .ZN(n6501)
         );
  INV_X1 U7428 ( .A(n6494), .ZN(n6495) );
  OAI211_X1 U7429 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n6496), .A(n6495), .B(
        STATE2_REG_2__SCAN_IN), .ZN(n6498) );
  AOI21_X1 U7430 ( .B1(n6498), .B2(STATE2_REG_0__SCAN_IN), .A(n6497), .ZN(
        n6500) );
  NAND2_X1 U7431 ( .A1(n6501), .A2(REQUESTPENDING_REG_SCAN_IN), .ZN(n6499) );
  OAI21_X1 U7432 ( .B1(n6501), .B2(n6500), .A(n6499), .ZN(U3472) );
  MUX2_X1 U7433 ( .A(MEMORYFETCH_REG_SCAN_IN), .B(M_IO_N_REG_SCAN_IN), .S(
        n6502), .Z(U3473) );
  NOR3_X1 U7434 ( .A1(keyinput26), .A2(keyinput32), .A3(keyinput18), .ZN(n6508) );
  NAND2_X1 U7435 ( .A1(keyinput44), .A2(keyinput35), .ZN(n6503) );
  NOR3_X1 U7436 ( .A1(keyinput16), .A2(keyinput57), .A3(n6503), .ZN(n6507) );
  INV_X1 U7437 ( .A(keyinput33), .ZN(n6505) );
  NAND4_X1 U7438 ( .A1(keyinput28), .A2(keyinput11), .A3(keyinput8), .A4(
        keyinput0), .ZN(n6504) );
  NOR4_X1 U7439 ( .A1(keyinput7), .A2(keyinput24), .A3(n6505), .A4(n6504), 
        .ZN(n6506) );
  NAND4_X1 U7440 ( .A1(keyinput62), .A2(n6508), .A3(n6507), .A4(n6506), .ZN(
        n6531) );
  NOR3_X1 U7441 ( .A1(keyinput19), .A2(keyinput20), .A3(keyinput25), .ZN(n6529) );
  NAND3_X1 U7442 ( .A1(keyinput54), .A2(keyinput48), .A3(keyinput38), .ZN(
        n6513) );
  NOR2_X1 U7443 ( .A1(keyinput51), .A2(keyinput6), .ZN(n6509) );
  NAND3_X1 U7444 ( .A1(keyinput22), .A2(keyinput56), .A3(n6509), .ZN(n6512) );
  NOR2_X1 U7445 ( .A1(keyinput49), .A2(keyinput2), .ZN(n6510) );
  NAND3_X1 U7446 ( .A1(keyinput40), .A2(keyinput23), .A3(n6510), .ZN(n6511) );
  NOR4_X1 U7447 ( .A1(keyinput29), .A2(n6513), .A3(n6512), .A4(n6511), .ZN(
        n6528) );
  NAND3_X1 U7448 ( .A1(keyinput50), .A2(keyinput60), .A3(keyinput63), .ZN(
        n6526) );
  NOR4_X1 U7449 ( .A1(keyinput13), .A2(keyinput42), .A3(keyinput61), .A4(
        keyinput15), .ZN(n6517) );
  NOR3_X1 U7450 ( .A1(keyinput3), .A2(keyinput53), .A3(keyinput17), .ZN(n6516)
         );
  NAND2_X1 U7451 ( .A1(keyinput45), .A2(keyinput59), .ZN(n6514) );
  NOR3_X1 U7452 ( .A1(keyinput37), .A2(keyinput27), .A3(n6514), .ZN(n6515) );
  NAND4_X1 U7453 ( .A1(n6517), .A2(keyinput39), .A3(n6516), .A4(n6515), .ZN(
        n6525) );
  NOR3_X1 U7454 ( .A1(keyinput58), .A2(keyinput55), .A3(keyinput46), .ZN(n6523) );
  INV_X1 U7455 ( .A(keyinput5), .ZN(n6518) );
  NOR4_X1 U7456 ( .A1(keyinput36), .A2(keyinput41), .A3(keyinput43), .A4(n6518), .ZN(n6522) );
  NAND3_X1 U7457 ( .A1(keyinput14), .A2(keyinput31), .A3(keyinput34), .ZN(
        n6520) );
  NAND3_X1 U7458 ( .A1(keyinput21), .A2(keyinput9), .A3(keyinput52), .ZN(n6519) );
  NOR4_X1 U7459 ( .A1(keyinput1), .A2(keyinput12), .A3(n6520), .A4(n6519), 
        .ZN(n6521) );
  NAND4_X1 U7460 ( .A1(keyinput4), .A2(n6523), .A3(n6522), .A4(n6521), .ZN(
        n6524) );
  NOR4_X1 U7461 ( .A1(keyinput47), .A2(n6526), .A3(n6525), .A4(n6524), .ZN(
        n6527) );
  NAND4_X1 U7462 ( .A1(keyinput30), .A2(n6529), .A3(n6528), .A4(n6527), .ZN(
        n6530) );
  OAI21_X1 U7463 ( .B1(n6531), .B2(n6530), .A(keyinput10), .ZN(n6666) );
  INV_X1 U7464 ( .A(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n6537) );
  INV_X1 U7465 ( .A(keyinput28), .ZN(n6536) );
  AOI22_X1 U7466 ( .A1(n6537), .A2(keyinput24), .B1(LWORD_REG_1__SCAN_IN), 
        .B2(n6536), .ZN(n6535) );
  OAI221_X1 U7467 ( .B1(n6537), .B2(keyinput24), .C1(n6536), .C2(
        LWORD_REG_1__SCAN_IN), .A(n6535), .ZN(n6546) );
  INV_X1 U7468 ( .A(keyinput8), .ZN(n6539) );
  AOI22_X1 U7469 ( .A1(n6540), .A2(keyinput11), .B1(DATAWIDTH_REG_12__SCAN_IN), 
        .B2(n6539), .ZN(n6538) );
  OAI221_X1 U7470 ( .B1(n6540), .B2(keyinput11), .C1(n6539), .C2(
        DATAWIDTH_REG_12__SCAN_IN), .A(n6538), .ZN(n6545) );
  INV_X1 U7471 ( .A(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n6542) );
  AOI22_X1 U7472 ( .A1(n6543), .A2(keyinput0), .B1(n6542), .B2(keyinput62), 
        .ZN(n6541) );
  OAI221_X1 U7473 ( .B1(n6543), .B2(keyinput0), .C1(n6542), .C2(keyinput62), 
        .A(n6541), .ZN(n6544) );
  NOR4_X1 U7474 ( .A1(n6547), .A2(n6546), .A3(n6545), .A4(n6544), .ZN(n6598)
         );
  INV_X1 U7475 ( .A(keyinput35), .ZN(n6549) );
  AOI22_X1 U7476 ( .A1(n6550), .A2(keyinput44), .B1(DATAO_REG_2__SCAN_IN), 
        .B2(n6549), .ZN(n6548) );
  OAI221_X1 U7477 ( .B1(n6550), .B2(keyinput44), .C1(n6549), .C2(
        DATAO_REG_2__SCAN_IN), .A(n6548), .ZN(n6563) );
  INV_X1 U7478 ( .A(keyinput18), .ZN(n6553) );
  INV_X1 U7479 ( .A(keyinput16), .ZN(n6552) );
  AOI22_X1 U7480 ( .A1(n6553), .A2(DATAO_REG_29__SCAN_IN), .B1(
        ADDRESS_REG_23__SCAN_IN), .B2(n6552), .ZN(n6551) );
  OAI221_X1 U7481 ( .B1(n6553), .B2(DATAO_REG_29__SCAN_IN), .C1(n6552), .C2(
        ADDRESS_REG_23__SCAN_IN), .A(n6551), .ZN(n6562) );
  INV_X1 U7482 ( .A(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n6556) );
  INV_X1 U7483 ( .A(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n6555) );
  AOI22_X1 U7484 ( .A1(n6556), .A2(keyinput26), .B1(n6555), .B2(keyinput32), 
        .ZN(n6554) );
  OAI221_X1 U7485 ( .B1(n6556), .B2(keyinput26), .C1(n6555), .C2(keyinput32), 
        .A(n6554), .ZN(n6561) );
  XOR2_X1 U7486 ( .A(n6557), .B(keyinput57), .Z(n6559) );
  XNOR2_X1 U7487 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B(keyinput50), .ZN(
        n6558) );
  NAND2_X1 U7488 ( .A1(n6559), .A2(n6558), .ZN(n6560) );
  NOR4_X1 U7489 ( .A1(n6563), .A2(n6562), .A3(n6561), .A4(n6560), .ZN(n6597)
         );
  INV_X1 U7490 ( .A(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n6566) );
  AOI22_X1 U7491 ( .A1(n6566), .A2(keyinput15), .B1(keyinput3), .B2(n6565), 
        .ZN(n6564) );
  OAI221_X1 U7492 ( .B1(n6566), .B2(keyinput15), .C1(n6565), .C2(keyinput3), 
        .A(n6564), .ZN(n6578) );
  INV_X1 U7493 ( .A(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n6568) );
  AOI22_X1 U7494 ( .A1(n5007), .A2(keyinput47), .B1(n6568), .B2(keyinput13), 
        .ZN(n6567) );
  OAI221_X1 U7495 ( .B1(n5007), .B2(keyinput47), .C1(n6568), .C2(keyinput13), 
        .A(n6567), .ZN(n6577) );
  AOI22_X1 U7496 ( .A1(n6571), .A2(keyinput60), .B1(n6570), .B2(keyinput63), 
        .ZN(n6569) );
  OAI221_X1 U7497 ( .B1(n6571), .B2(keyinput60), .C1(n6570), .C2(keyinput63), 
        .A(n6569), .ZN(n6576) );
  XOR2_X1 U7498 ( .A(n6572), .B(keyinput42), .Z(n6574) );
  XNOR2_X1 U7499 ( .A(INSTQUEUE_REG_3__5__SCAN_IN), .B(keyinput61), .ZN(n6573)
         );
  NAND2_X1 U7500 ( .A1(n6574), .A2(n6573), .ZN(n6575) );
  NOR4_X1 U7501 ( .A1(n6578), .A2(n6577), .A3(n6576), .A4(n6575), .ZN(n6596)
         );
  INV_X1 U7502 ( .A(DATAI_19_), .ZN(n6581) );
  AOI22_X1 U7503 ( .A1(n6581), .A2(keyinput39), .B1(n6580), .B2(keyinput53), 
        .ZN(n6579) );
  OAI221_X1 U7504 ( .B1(n6581), .B2(keyinput39), .C1(n6580), .C2(keyinput53), 
        .A(n6579), .ZN(n6594) );
  INV_X1 U7505 ( .A(keyinput59), .ZN(n6583) );
  AOI22_X1 U7506 ( .A1(n6584), .A2(keyinput17), .B1(ADDRESS_REG_27__SCAN_IN), 
        .B2(n6583), .ZN(n6582) );
  OAI221_X1 U7507 ( .B1(n6584), .B2(keyinput17), .C1(n6583), .C2(
        ADDRESS_REG_27__SCAN_IN), .A(n6582), .ZN(n6593) );
  INV_X1 U7508 ( .A(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n6587) );
  AOI22_X1 U7509 ( .A1(n6587), .A2(keyinput27), .B1(keyinput37), .B2(n6586), 
        .ZN(n6585) );
  OAI221_X1 U7510 ( .B1(n6587), .B2(keyinput27), .C1(n6586), .C2(keyinput37), 
        .A(n6585), .ZN(n6592) );
  INV_X1 U7511 ( .A(keyinput45), .ZN(n6589) );
  AOI22_X1 U7512 ( .A1(n6590), .A2(keyinput54), .B1(DATAWIDTH_REG_24__SCAN_IN), 
        .B2(n6589), .ZN(n6588) );
  OAI221_X1 U7513 ( .B1(n6590), .B2(keyinput54), .C1(n6589), .C2(
        DATAWIDTH_REG_24__SCAN_IN), .A(n6588), .ZN(n6591) );
  NOR4_X1 U7514 ( .A1(n6594), .A2(n6593), .A3(n6592), .A4(n6591), .ZN(n6595)
         );
  NAND4_X1 U7515 ( .A1(n6598), .A2(n6597), .A3(n6596), .A4(n6595), .ZN(n6665)
         );
  INV_X1 U7516 ( .A(keyinput23), .ZN(n6600) );
  AOI22_X1 U7517 ( .A1(n4024), .A2(keyinput6), .B1(DATAWIDTH_REG_0__SCAN_IN), 
        .B2(n6600), .ZN(n6599) );
  OAI221_X1 U7518 ( .B1(n4024), .B2(keyinput6), .C1(n6600), .C2(
        DATAWIDTH_REG_0__SCAN_IN), .A(n6599), .ZN(n6611) );
  INV_X1 U7519 ( .A(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n6603) );
  INV_X1 U7520 ( .A(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n6602) );
  AOI22_X1 U7521 ( .A1(n6603), .A2(keyinput22), .B1(n6602), .B2(keyinput51), 
        .ZN(n6601) );
  OAI221_X1 U7522 ( .B1(n6603), .B2(keyinput22), .C1(n6602), .C2(keyinput51), 
        .A(n6601), .ZN(n6610) );
  AOI22_X1 U7523 ( .A1(n5370), .A2(keyinput40), .B1(n6607), .B2(keyinput49), 
        .ZN(n6606) );
  OAI221_X1 U7524 ( .B1(n5370), .B2(keyinput40), .C1(n6607), .C2(keyinput49), 
        .A(n6606), .ZN(n6608) );
  NOR4_X1 U7525 ( .A1(n6611), .A2(n6610), .A3(n6609), .A4(n6608), .ZN(n6663)
         );
  INV_X1 U7526 ( .A(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n6613) );
  AOI22_X1 U7527 ( .A1(n6614), .A2(keyinput38), .B1(n6613), .B2(keyinput19), 
        .ZN(n6612) );
  OAI221_X1 U7528 ( .B1(n6614), .B2(keyinput38), .C1(n6613), .C2(keyinput19), 
        .A(n6612), .ZN(n6627) );
  INV_X1 U7529 ( .A(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n6617) );
  INV_X1 U7530 ( .A(keyinput29), .ZN(n6616) );
  AOI22_X1 U7531 ( .A1(n6617), .A2(keyinput48), .B1(DATAWIDTH_REG_27__SCAN_IN), 
        .B2(n6616), .ZN(n6615) );
  OAI221_X1 U7532 ( .B1(n6617), .B2(keyinput48), .C1(n6616), .C2(
        DATAWIDTH_REG_27__SCAN_IN), .A(n6615), .ZN(n6626) );
  INV_X1 U7533 ( .A(keyinput56), .ZN(n6619) );
  AOI22_X1 U7534 ( .A1(n6620), .A2(keyinput30), .B1(DATAO_REG_28__SCAN_IN), 
        .B2(n6619), .ZN(n6618) );
  OAI221_X1 U7535 ( .B1(n6620), .B2(keyinput30), .C1(n6619), .C2(
        DATAO_REG_28__SCAN_IN), .A(n6618), .ZN(n6625) );
  AOI22_X1 U7536 ( .A1(n6623), .A2(keyinput20), .B1(n6622), .B2(keyinput25), 
        .ZN(n6621) );
  OAI221_X1 U7537 ( .B1(n6623), .B2(keyinput20), .C1(n6622), .C2(keyinput25), 
        .A(n6621), .ZN(n6624) );
  NOR4_X1 U7538 ( .A1(n6627), .A2(n6626), .A3(n6625), .A4(n6624), .ZN(n6662)
         );
  INV_X1 U7539 ( .A(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n6630) );
  INV_X1 U7540 ( .A(keyinput52), .ZN(n6629) );
  AOI22_X1 U7541 ( .A1(n6630), .A2(keyinput5), .B1(DATAO_REG_16__SCAN_IN), 
        .B2(n6629), .ZN(n6628) );
  OAI221_X1 U7542 ( .B1(n6630), .B2(keyinput5), .C1(n6629), .C2(
        DATAO_REG_16__SCAN_IN), .A(n6628), .ZN(n6643) );
  AOI22_X1 U7543 ( .A1(n6633), .A2(keyinput21), .B1(keyinput9), .B2(n6632), 
        .ZN(n6631) );
  OAI221_X1 U7544 ( .B1(n6633), .B2(keyinput21), .C1(n6632), .C2(keyinput9), 
        .A(n6631), .ZN(n6642) );
  AOI22_X1 U7545 ( .A1(n6636), .A2(keyinput33), .B1(n6635), .B2(keyinput43), 
        .ZN(n6634) );
  OAI221_X1 U7546 ( .B1(n6636), .B2(keyinput33), .C1(n6635), .C2(keyinput43), 
        .A(n6634), .ZN(n6641) );
  INV_X1 U7547 ( .A(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n6639) );
  INV_X1 U7548 ( .A(keyinput36), .ZN(n6638) );
  AOI22_X1 U7549 ( .A1(n6639), .A2(keyinput41), .B1(ADDRESS_REG_16__SCAN_IN), 
        .B2(n6638), .ZN(n6637) );
  OAI221_X1 U7550 ( .B1(n6639), .B2(keyinput41), .C1(n6638), .C2(
        ADDRESS_REG_16__SCAN_IN), .A(n6637), .ZN(n6640) );
  NOR4_X1 U7551 ( .A1(n6643), .A2(n6642), .A3(n6641), .A4(n6640), .ZN(n6661)
         );
  AOI22_X1 U7552 ( .A1(n6646), .A2(keyinput4), .B1(n6645), .B2(keyinput14), 
        .ZN(n6644) );
  OAI221_X1 U7553 ( .B1(n6646), .B2(keyinput4), .C1(n6645), .C2(keyinput14), 
        .A(n6644), .ZN(n6659) );
  INV_X1 U7554 ( .A(keyinput55), .ZN(n6649) );
  INV_X1 U7555 ( .A(keyinput46), .ZN(n6648) );
  AOI22_X1 U7556 ( .A1(n6649), .A2(DATAWIDTH_REG_8__SCAN_IN), .B1(
        DATAO_REG_18__SCAN_IN), .B2(n6648), .ZN(n6647) );
  OAI221_X1 U7557 ( .B1(n6649), .B2(DATAWIDTH_REG_8__SCAN_IN), .C1(n6648), 
        .C2(DATAO_REG_18__SCAN_IN), .A(n6647), .ZN(n6658) );
  INV_X1 U7558 ( .A(keyinput1), .ZN(n6651) );
  AOI22_X1 U7559 ( .A1(n6652), .A2(keyinput12), .B1(DATAWIDTH_REG_3__SCAN_IN), 
        .B2(n6651), .ZN(n6650) );
  OAI221_X1 U7560 ( .B1(n6652), .B2(keyinput12), .C1(n6651), .C2(
        DATAWIDTH_REG_3__SCAN_IN), .A(n6650), .ZN(n6657) );
  INV_X1 U7561 ( .A(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n6655) );
  INV_X1 U7562 ( .A(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n6654) );
  AOI22_X1 U7563 ( .A1(n6655), .A2(keyinput31), .B1(keyinput34), .B2(n6654), 
        .ZN(n6653) );
  OAI221_X1 U7564 ( .B1(n6655), .B2(keyinput31), .C1(n6654), .C2(keyinput34), 
        .A(n6653), .ZN(n6656) );
  NOR4_X1 U7565 ( .A1(n6659), .A2(n6658), .A3(n6657), .A4(n6656), .ZN(n6660)
         );
  NAND4_X1 U7566 ( .A1(n6663), .A2(n6662), .A3(n6661), .A4(n6660), .ZN(n6664)
         );
  AOI211_X1 U7567 ( .C1(INSTQUEUE_REG_2__1__SCAN_IN), .C2(n6666), .A(n6665), 
        .B(n6664), .ZN(n6672) );
  AOI22_X1 U7568 ( .A1(UWORD_REG_10__SCAN_IN), .A2(n6668), .B1(n6667), .B2(
        EAX_REG_26__SCAN_IN), .ZN(n6669) );
  NAND2_X1 U7569 ( .A1(n6670), .A2(n6669), .ZN(n6671) );
  XOR2_X1 U7570 ( .A(n6672), .B(n6671), .Z(U2934) );
  INV_X1 U3893 ( .A(n4370), .ZN(n3155) );
  CLKBUF_X1 U3420 ( .A(n3964), .Z(n3859) );
  OR2_X1 U4068 ( .A1(n3234), .A2(n3233), .ZN(n3235) );
  NAND2_X1 U4413 ( .A1(n3525), .A2(n3524), .ZN(n4476) );
  AND2_X2 U3450 ( .A1(n4503), .A2(n2988), .ZN(n3043) );
  INV_X1 U3747 ( .A(n3097), .ZN(n4217) );
  CLKBUF_X1 U34630 ( .A(n3972), .Z(n3879) );
  CLKBUF_X1 U3476 ( .A(n3126), .Z(n4506) );
  CLKBUF_X1 U3498 ( .A(n3121), .Z(n4363) );
  INV_X1 U3605 ( .A(n4221), .ZN(n5270) );
  CLKBUF_X1 U3646 ( .A(n4343), .Z(n5627) );
  CLKBUF_X1 U3724 ( .A(n5116), .Z(n5133) );
  CLKBUF_X1 U3965 ( .A(n5888), .Z(n5917) );
  INV_X2 U4033 ( .A(n6368), .ZN(n6493) );
endmodule

