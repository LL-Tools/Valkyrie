

module b21_C_SARLock_k_128_2 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3, 
        keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, 
        keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, 
        keyinput16, keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, 
        keyinput22, keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, 
        keyinput28, keyinput29, keyinput30, keyinput31, keyinput32, keyinput33, 
        keyinput34, keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, 
        keyinput40, keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, 
        keyinput46, keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, 
        keyinput52, keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, 
        keyinput58, keyinput59, keyinput60, keyinput61, keyinput62, keyinput63, 
        keyinput64, keyinput65, keyinput66, keyinput67, keyinput68, keyinput69, 
        keyinput70, keyinput71, keyinput72, keyinput73, keyinput74, keyinput75, 
        keyinput76, keyinput77, keyinput78, keyinput79, keyinput80, keyinput81, 
        keyinput82, keyinput83, keyinput84, keyinput85, keyinput86, keyinput87, 
        keyinput88, keyinput89, keyinput90, keyinput91, keyinput92, keyinput93, 
        keyinput94, keyinput95, keyinput96, keyinput97, keyinput98, keyinput99, 
        keyinput100, keyinput101, keyinput102, keyinput103, keyinput104, 
        keyinput105, keyinput106, keyinput107, keyinput108, keyinput109, 
        keyinput110, keyinput111, keyinput112, keyinput113, keyinput114, 
        keyinput115, keyinput116, keyinput117, keyinput118, keyinput119, 
        keyinput120, keyinput121, keyinput122, keyinput123, keyinput124, 
        keyinput125, keyinput126, keyinput127, ADD_1071_U4, ADD_1071_U55, 
        ADD_1071_U56, ADD_1071_U57, ADD_1071_U58, ADD_1071_U59, ADD_1071_U60, 
        ADD_1071_U61, ADD_1071_U62, ADD_1071_U63, ADD_1071_U47, ADD_1071_U48, 
        ADD_1071_U49, ADD_1071_U50, ADD_1071_U51, ADD_1071_U52, ADD_1071_U53, 
        ADD_1071_U54, ADD_1071_U5, ADD_1071_U46, U126, U123, P1_U3353, 
        P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, 
        P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, 
        P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, 
        P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, 
        P1_U3324, P1_U3323, P1_U3322, P1_U3440, P1_U3441, P1_U3321, P1_U3320, 
        P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, 
        P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, 
        P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, 
        P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, P1_U3293, P1_U3292, 
        P1_U3454, P1_U3457, P1_U3460, P1_U3463, P1_U3466, P1_U3469, P1_U3472, 
        P1_U3475, P1_U3478, P1_U3481, P1_U3484, P1_U3487, P1_U3490, P1_U3493, 
        P1_U3496, P1_U3499, P1_U3502, P1_U3505, P1_U3508, P1_U3510, P1_U3511, 
        P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, 
        P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, 
        P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, 
        P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, 
        P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, 
        P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, 
        P1_U3554, P1_U3291, P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, 
        P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, 
        P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, 
        P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, 
        P1_U3264, P1_U3263, P1_U3355, P1_U3262, P1_U3261, P1_U3260, P1_U3259, 
        P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, 
        P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, 
        P1_U3244, P1_U3243, P1_U3242, P1_U3241, P1_U3555, P1_U3556, P1_U3557, 
        P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, 
        P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, 
        P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, 
        P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, 
        P1_U3586, P1_U3240, P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, 
        P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, 
        P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, 
        P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, 
        P1_U3213, P1_U3212, P1_U3211, P1_U3084, P1_U3083, P1_U4006, P2_U3358, 
        P2_U3357, P2_U3356, P2_U3355, P2_U3354, P2_U3353, P2_U3352, P2_U3351, 
        P2_U3350, P2_U3349, P2_U3348, P2_U3347, P2_U3346, P2_U3345, P2_U3344, 
        P2_U3343, P2_U3342, P2_U3341, P2_U3340, P2_U3339, P2_U3338, P2_U3337, 
        P2_U3336, P2_U3335, P2_U3334, P2_U3333, P2_U3332, P2_U3331, P2_U3330, 
        P2_U3329, P2_U3328, P2_U3327, P2_U3437, P2_U3438, P2_U3326, P2_U3325, 
        P2_U3324, P2_U3323, P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, 
        P2_U3317, P2_U3316, P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, 
        P2_U3310, P2_U3309, P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, 
        P2_U3303, P2_U3302, P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, 
        P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, 
        P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, P2_U3487, P2_U3490, 
        P2_U3493, P2_U3496, P2_U3499, P2_U3502, P2_U3505, P2_U3507, P2_U3508, 
        P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, 
        P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, 
        P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, 
        P2_U3530, P2_U3531, P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, 
        P2_U3537, P2_U3538, P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, 
        P2_U3544, P2_U3545, P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, 
        P2_U3551, P2_U3296, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, 
        P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, 
        P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, 
        P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, 
        P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3263, 
        P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, 
        P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, 
        P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3552, P2_U3553, P2_U3554, 
        P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, 
        P2_U3562, P2_U3563, P2_U3564, P2_U3565, P2_U3566, P2_U3567, P2_U3568, 
        P2_U3569, P2_U3570, P2_U3571, P2_U3572, P2_U3573, P2_U3574, P2_U3575, 
        P2_U3576, P2_U3577, P2_U3578, P2_U3579, P2_U3580, P2_U3581, P2_U3582, 
        P2_U3583, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, 
        P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, 
        P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, 
        P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, 
        P2_U3217, P2_U3216, P2_U3215, P2_U3152, P2_U3151, P2_U3966 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n4387, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398,
         n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408,
         n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418,
         n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428,
         n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438,
         n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448,
         n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458,
         n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468,
         n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478,
         n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488,
         n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498,
         n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508,
         n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518,
         n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528,
         n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538,
         n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548,
         n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558,
         n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568,
         n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578,
         n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588,
         n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598,
         n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608,
         n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618,
         n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628,
         n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638,
         n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648,
         n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658,
         n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668,
         n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678,
         n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688,
         n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698,
         n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708,
         n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718,
         n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728,
         n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738,
         n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748,
         n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758,
         n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768,
         n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778,
         n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788,
         n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798,
         n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808,
         n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818,
         n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828,
         n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838,
         n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848,
         n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858,
         n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868,
         n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878,
         n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888,
         n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898,
         n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908,
         n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918,
         n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928,
         n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938,
         n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948,
         n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958,
         n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968,
         n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978,
         n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988,
         n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998,
         n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008,
         n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018,
         n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028,
         n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038,
         n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048,
         n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058,
         n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068,
         n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078,
         n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088,
         n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098,
         n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108,
         n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118,
         n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128,
         n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138,
         n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148,
         n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158,
         n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168,
         n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178,
         n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188,
         n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198,
         n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208,
         n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218,
         n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228,
         n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238,
         n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248,
         n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258,
         n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268,
         n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278,
         n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288,
         n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298,
         n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308,
         n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318,
         n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328,
         n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338,
         n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348,
         n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358,
         n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368,
         n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378,
         n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388,
         n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398,
         n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408,
         n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418,
         n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428,
         n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438,
         n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448,
         n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458,
         n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468,
         n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478,
         n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488,
         n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498,
         n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508,
         n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518,
         n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528,
         n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538,
         n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548,
         n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558,
         n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568,
         n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578,
         n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588,
         n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598,
         n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608,
         n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618,
         n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628,
         n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638,
         n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648,
         n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658,
         n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668,
         n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678,
         n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688,
         n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698,
         n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708,
         n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718,
         n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728,
         n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738,
         n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748,
         n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758,
         n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768,
         n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778,
         n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788,
         n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798,
         n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808,
         n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818,
         n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828,
         n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838,
         n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848,
         n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858,
         n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868,
         n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878,
         n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888,
         n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898,
         n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908,
         n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918,
         n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928,
         n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938,
         n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948,
         n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958,
         n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968,
         n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978,
         n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988,
         n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998,
         n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008,
         n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018,
         n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028,
         n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038,
         n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048,
         n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058,
         n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068,
         n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078,
         n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088,
         n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098,
         n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108,
         n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118,
         n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128,
         n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138,
         n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148,
         n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158,
         n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168,
         n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178,
         n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188,
         n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198,
         n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208,
         n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218,
         n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228,
         n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238,
         n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248,
         n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258,
         n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268,
         n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278,
         n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288,
         n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298,
         n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308,
         n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318,
         n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328,
         n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338,
         n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348,
         n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358,
         n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368,
         n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378,
         n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388,
         n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398,
         n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408,
         n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418,
         n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428,
         n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438,
         n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448,
         n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458,
         n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468,
         n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478,
         n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488,
         n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498,
         n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508,
         n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518,
         n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528,
         n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538,
         n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548,
         n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558,
         n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568,
         n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578,
         n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588,
         n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598,
         n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608,
         n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618,
         n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628,
         n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638,
         n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648,
         n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658,
         n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668,
         n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678,
         n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688,
         n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698,
         n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708,
         n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718,
         n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728,
         n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738,
         n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748,
         n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758,
         n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768,
         n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778,
         n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788,
         n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798,
         n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808,
         n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818,
         n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828,
         n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838,
         n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848,
         n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858,
         n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868,
         n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878,
         n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888,
         n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898,
         n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908,
         n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918,
         n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928,
         n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938,
         n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948,
         n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958,
         n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968,
         n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978,
         n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988,
         n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998,
         n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008,
         n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018,
         n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028,
         n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038,
         n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048,
         n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058,
         n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068,
         n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078,
         n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088,
         n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098,
         n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108,
         n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118,
         n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128,
         n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138,
         n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148,
         n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158,
         n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168,
         n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178,
         n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188,
         n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198,
         n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208,
         n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218,
         n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228,
         n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238,
         n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248,
         n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258,
         n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268,
         n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278,
         n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288,
         n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298,
         n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308,
         n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318,
         n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328,
         n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338,
         n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348,
         n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358,
         n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368,
         n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378,
         n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388,
         n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398,
         n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408,
         n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418,
         n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428,
         n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438,
         n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448,
         n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458,
         n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468,
         n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478,
         n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488,
         n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498,
         n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508,
         n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518,
         n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528,
         n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538,
         n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548,
         n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558,
         n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568,
         n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578,
         n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588,
         n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598,
         n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608,
         n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618,
         n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628,
         n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638,
         n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648,
         n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658,
         n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668,
         n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678,
         n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688,
         n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698,
         n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708,
         n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718,
         n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728,
         n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738,
         n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748,
         n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758,
         n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768,
         n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778,
         n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788,
         n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798,
         n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808,
         n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818,
         n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828,
         n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838,
         n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848,
         n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858,
         n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868,
         n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878,
         n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888,
         n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898,
         n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908,
         n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918,
         n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928,
         n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938,
         n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948,
         n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958,
         n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968,
         n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978,
         n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988,
         n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998,
         n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008,
         n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018,
         n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028,
         n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038,
         n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048,
         n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058,
         n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068,
         n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078,
         n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088,
         n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098,
         n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108,
         n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118,
         n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128,
         n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138,
         n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148,
         n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158,
         n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168,
         n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178,
         n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188,
         n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198,
         n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208,
         n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218,
         n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228,
         n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238,
         n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248,
         n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258,
         n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268,
         n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278,
         n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288,
         n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298,
         n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308,
         n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318,
         n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328,
         n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338,
         n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348,
         n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358,
         n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368,
         n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378,
         n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388,
         n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398,
         n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408,
         n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418,
         n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428,
         n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438,
         n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448,
         n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458,
         n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468,
         n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478,
         n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488,
         n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498,
         n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508,
         n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518,
         n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528,
         n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538,
         n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548,
         n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558,
         n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568,
         n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578,
         n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588,
         n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598,
         n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608,
         n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618,
         n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628,
         n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638,
         n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648,
         n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658,
         n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668,
         n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678,
         n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688,
         n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698,
         n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708,
         n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718,
         n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728,
         n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738,
         n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748,
         n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758,
         n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768,
         n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778,
         n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788,
         n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798,
         n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808,
         n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818,
         n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828,
         n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838,
         n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848,
         n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858,
         n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868,
         n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878,
         n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888,
         n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898,
         n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908,
         n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918,
         n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928,
         n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938,
         n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948,
         n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958,
         n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968,
         n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978,
         n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988,
         n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998,
         n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008,
         n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018,
         n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028,
         n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038,
         n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048,
         n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058,
         n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068,
         n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078,
         n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088,
         n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098,
         n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108,
         n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118,
         n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128,
         n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138,
         n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148,
         n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158,
         n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168,
         n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178,
         n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188,
         n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198,
         n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208,
         n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218,
         n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228,
         n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238,
         n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248,
         n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258,
         n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268,
         n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278,
         n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288,
         n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298,
         n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308,
         n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318,
         n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328,
         n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338,
         n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348,
         n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358,
         n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368,
         n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378,
         n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388,
         n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398,
         n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408,
         n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418,
         n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428,
         n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438,
         n9439, n9440, n9441, n9442, n9444, n9445, n9446, n9447, n9448, n9449,
         n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459,
         n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469,
         n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479,
         n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489,
         n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499,
         n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509,
         n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519,
         n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529,
         n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539,
         n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549,
         n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559,
         n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569,
         n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579,
         n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589,
         n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599,
         n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609,
         n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619,
         n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629,
         n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639,
         n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649,
         n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659,
         n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669,
         n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679,
         n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689,
         n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699,
         n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709,
         n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719,
         n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729,
         n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739,
         n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749,
         n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759,
         n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769,
         n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779,
         n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789,
         n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799,
         n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809,
         n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819,
         n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829,
         n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839,
         n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849,
         n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859,
         n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869,
         n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879,
         n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889,
         n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899,
         n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909,
         n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919,
         n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929,
         n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939,
         n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949,
         n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959,
         n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969,
         n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979,
         n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989,
         n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999,
         n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
         n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
         n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
         n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
         n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
         n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
         n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247,
         n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255,
         n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263,
         n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271;

  OAI21_X1 U4893 ( .B1(n7488), .B2(n7487), .A(n6755), .ZN(n7655) );
  CLKBUF_X2 U4894 ( .A(n6435), .Z(n6646) );
  INV_X2 U4895 ( .A(n6928), .ZN(n6186) );
  INV_X1 U4896 ( .A(n6315), .ZN(n6288) );
  OR2_X1 U4897 ( .A1(n8668), .A2(n5873), .ZN(n6315) );
  INV_X1 U4898 ( .A(n6726), .ZN(n8165) );
  INV_X2 U4899 ( .A(n6497), .ZN(n6547) );
  OR2_X1 U4900 ( .A1(n9117), .A2(n8112), .ZN(n4889) );
  INV_X1 U4901 ( .A(n6547), .ZN(n7466) );
  OAI21_X1 U4902 ( .B1(n7877), .B2(n4580), .A(n4578), .ZN(n7959) );
  INV_X2 U4903 ( .A(n8165), .ZN(n8212) );
  BUF_X1 U4904 ( .A(n5991), .Z(n6304) );
  NAND2_X1 U4905 ( .A1(n6065), .A2(n6045), .ZN(n10077) );
  AND3_X1 U4906 ( .A1(n5954), .A2(n5953), .A3(n5952), .ZN(n10141) );
  INV_X1 U4907 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n6416) );
  NAND2_X1 U4908 ( .A1(n8900), .A2(n8901), .ZN(n8899) );
  NAND2_X1 U4909 ( .A1(n8899), .A2(n4782), .ZN(n6631) );
  XNOR2_X1 U4911 ( .A(n5129), .B(P1_IR_REG_28__SCAN_IN), .ZN(n5803) );
  NAND2_X1 U4912 ( .A1(n8497), .A2(n8496), .ZN(n8517) );
  INV_X2 U4913 ( .A(n4975), .ZN(n5831) );
  INV_X1 U4914 ( .A(n6434), .ZN(n6437) );
  NAND2_X1 U4915 ( .A1(n5537), .A2(n5536), .ZN(n9849) );
  NAND2_X1 U4916 ( .A1(n5165), .A2(n9442), .ZN(n4387) );
  NAND2_X4 U4917 ( .A1(n4393), .A2(n4394), .ZN(n5388) );
  OAI21_X1 U4918 ( .B1(n4407), .B2(n4602), .A(n4601), .ZN(n4600) );
  NAND4_X4 U4919 ( .A1(n5980), .A2(n5978), .A3(n5979), .A4(n5981), .ZN(n6718)
         );
  NAND2_X1 U4921 ( .A1(n6930), .A2(n8464), .ZN(n4390) );
  NAND2_X1 U4922 ( .A1(n6930), .A2(n8464), .ZN(n6928) );
  OAI21_X2 U4923 ( .B1(n5558), .B2(P1_IR_REG_19__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5748) );
  XNOR2_X2 U4924 ( .A(n5529), .B(n5528), .ZN(n6919) );
  AOI22_X2 U4925 ( .A1(n8566), .A2(n8569), .B1(n8592), .B2(n8580), .ZN(n8550)
         );
  NAND2_X2 U4926 ( .A1(n4937), .A2(n4938), .ZN(n8566) );
  AND2_X1 U4927 ( .A1(n5166), .A2(n5165), .ZN(n4391) );
  NAND2_X4 U4928 ( .A1(n7680), .A2(n4489), .ZN(n6724) );
  NOR2_X1 U4929 ( .A1(n5740), .A2(n5739), .ZN(n5746) );
  NAND2_X1 U4930 ( .A1(n5756), .A2(n5757), .ZN(n7511) );
  INV_X1 U4931 ( .A(n7785), .ZN(n6740) );
  NAND2_X1 U4932 ( .A1(n6332), .A2(n7242), .ZN(n10101) );
  NAND2_X1 U4933 ( .A1(n6334), .A2(n6358), .ZN(n7773) );
  NAND2_X1 U4934 ( .A1(n8351), .A2(n10147), .ZN(n7242) );
  INV_X1 U4935 ( .A(n7566), .ZN(n10003) );
  INV_X1 U4936 ( .A(n7520), .ZN(n9997) );
  INV_X1 U4937 ( .A(n6718), .ZN(n4943) );
  OAI21_X1 U4938 ( .B1(n7005), .B2(n6887), .A(n4628), .ZN(n7520) );
  INV_X1 U4939 ( .A(n6694), .ZN(n7373) );
  INV_X1 U4940 ( .A(n5464), .ZN(n4589) );
  CLKBUF_X2 U4941 ( .A(n6202), .Z(n6251) );
  NAND2_X1 U4942 ( .A1(n6433), .A2(n7494), .ZN(n6694) );
  NAND2_X4 U4943 ( .A1(n5388), .A2(n5831), .ZN(n5464) );
  AND2_X1 U4944 ( .A1(n5166), .A2(n9447), .ZN(n5453) );
  NAND2_X1 U4945 ( .A1(n5830), .A2(n5829), .ZN(n8464) );
  CLKBUF_X2 U4946 ( .A(n5804), .Z(n4394) );
  NOR2_X1 U4947 ( .A1(n6004), .A2(n6003), .ZN(n9752) );
  INV_X4 U4948 ( .A(n5831), .ZN(n6891) );
  INV_X2 U4949 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  AOI21_X1 U4950 ( .B1(n4708), .B2(n9963), .A(n4707), .ZN(n9344) );
  AND2_X1 U4951 ( .A1(n5750), .A2(n7398), .ZN(n5751) );
  AND2_X1 U4952 ( .A1(n9141), .A2(n4596), .ZN(n9123) );
  NAND2_X1 U4953 ( .A1(n4599), .A2(n4598), .ZN(n9141) );
  OAI21_X1 U4954 ( .B1(n4603), .B2(n8087), .A(n4408), .ZN(n5735) );
  NAND2_X1 U4955 ( .A1(n8969), .A2(n8966), .ZN(n8893) );
  NAND2_X1 U4956 ( .A1(n8071), .A2(n9258), .ZN(n9263) );
  NAND2_X1 U4957 ( .A1(n8176), .A2(n6786), .ZN(n8249) );
  OR2_X1 U4958 ( .A1(n9276), .A2(n8099), .ZN(n8101) );
  NAND2_X1 U4959 ( .A1(n6247), .A2(n6246), .ZN(n8774) );
  INV_X1 U4960 ( .A(n8607), .ZN(n8789) );
  NAND2_X1 U4961 ( .A1(n6526), .A2(n4431), .ZN(n7723) );
  NAND2_X1 U4962 ( .A1(n7574), .A2(n7576), .ZN(n6526) );
  NAND2_X1 U4963 ( .A1(n7870), .A2(n7869), .ZN(n9840) );
  AOI21_X1 U4964 ( .B1(n4946), .B2(n4945), .A(n4439), .ZN(n4944) );
  NAND2_X1 U4965 ( .A1(n5294), .A2(n5293), .ZN(n9388) );
  OR2_X1 U4966 ( .A1(n7637), .A2(n7643), .ZN(n7870) );
  AND2_X1 U4967 ( .A1(n7807), .A2(n7806), .ZN(n7808) );
  AND2_X1 U4968 ( .A1(n7943), .A2(n4825), .ZN(n4824) );
  NAND2_X1 U4969 ( .A1(n8299), .A2(n6750), .ZN(n7488) );
  NAND2_X1 U4970 ( .A1(n6073), .A2(n6072), .ZN(n7950) );
  NAND2_X1 U4971 ( .A1(n7164), .A2(n6465), .ZN(n7198) );
  NAND2_X1 U4972 ( .A1(n5520), .A2(n5519), .ZN(n7868) );
  NAND2_X1 U4973 ( .A1(n6052), .A2(n6051), .ZN(n10178) );
  NAND2_X1 U4974 ( .A1(n4488), .A2(n7274), .ZN(n7278) );
  NAND2_X1 U4975 ( .A1(n7240), .A2(n7239), .ZN(n7665) );
  NAND2_X1 U4976 ( .A1(n7276), .A2(n6731), .ZN(n4488) );
  AND2_X1 U4977 ( .A1(n5630), .A2(n5631), .ZN(n7618) );
  XNOR2_X1 U4978 ( .A(n5501), .B(n5502), .ZN(n6902) );
  INV_X2 U4979 ( .A(n10053), .ZN(n4392) );
  BUF_X4 U4980 ( .A(n6458), .Z(n4395) );
  NAND4_X1 U4981 ( .A1(n5407), .A2(n5406), .A3(n5405), .A4(n5404), .ZN(n9016)
         );
  NAND2_X1 U4982 ( .A1(n5458), .A2(n5457), .ZN(n6440) );
  NAND2_X1 U4983 ( .A1(n5417), .A2(n4416), .ZN(n9018) );
  CLKBUF_X1 U4984 ( .A(n6716), .Z(n8059) );
  NAND4_X1 U4985 ( .A1(n5935), .A2(n5934), .A3(n5933), .A4(n5932), .ZN(n8351)
         );
  XNOR2_X1 U4986 ( .A(n4787), .B(P2_IR_REG_20__SCAN_IN), .ZN(n6716) );
  INV_X1 U4987 ( .A(n6322), .ZN(n8668) );
  INV_X2 U4988 ( .A(n5890), .ZN(n6305) );
  AND2_X4 U4989 ( .A1(n7373), .A2(n6834), .ZN(n6458) );
  NAND4_X1 U4990 ( .A1(n5948), .A2(n5947), .A3(n5946), .A4(n5945), .ZN(n8352)
         );
  INV_X2 U4991 ( .A(n5463), .ZN(n4613) );
  AND2_X2 U4992 ( .A1(n6860), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U4006) );
  INV_X4 U4993 ( .A(n4387), .ZN(n4397) );
  INV_X2 U4994 ( .A(n6307), .ZN(n6294) );
  XNOR2_X1 U4995 ( .A(n6319), .B(P2_IR_REG_19__SCAN_IN), .ZN(n6322) );
  OR2_X1 U4996 ( .A1(n6202), .A2(n7770), .ZN(n5979) );
  AND2_X2 U4997 ( .A1(n6694), .A2(n6834), .ZN(n6435) );
  INV_X2 U4998 ( .A(n5964), .ZN(n6234) );
  AND2_X2 U4999 ( .A1(n5166), .A2(n5165), .ZN(n5542) );
  NAND2_X1 U5000 ( .A1(n5857), .A2(n8850), .ZN(n5992) );
  NAND2_X1 U5001 ( .A1(n5388), .A2(n6891), .ZN(n5463) );
  AND2_X1 U5002 ( .A1(n4390), .A2(n5831), .ZN(n6001) );
  CLKBUF_X2 U5003 ( .A(n5803), .Z(n4393) );
  OAI21_X1 U5004 ( .B1(n5462), .B2(n4731), .A(n4972), .ZN(n5422) );
  MUX2_X1 U5005 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5828), .S(
        P2_IR_REG_27__SCAN_IN), .Z(n5830) );
  OAI21_X1 U5006 ( .B1(n5137), .B2(P1_IR_REG_27__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5136) );
  NAND2_X1 U5007 ( .A1(n4499), .A2(n4501), .ZN(n5829) );
  NAND2_X2 U5008 ( .A1(n5831), .A2(P2_U3152), .ZN(n8859) );
  NOR2_X1 U5009 ( .A1(n4451), .A2(n4910), .ZN(n4909) );
  AND2_X1 U5010 ( .A1(n5285), .A2(n4952), .ZN(n5786) );
  BUF_X2 U5011 ( .A(n5285), .Z(n5475) );
  AND3_X1 U5012 ( .A1(n5921), .A2(n5825), .A3(n5811), .ZN(n4501) );
  AND3_X1 U5013 ( .A1(n4791), .A2(n4789), .A3(n4788), .ZN(n5921) );
  NOR2_X1 U5014 ( .A1(n5126), .A2(n5125), .ZN(n4952) );
  AND2_X1 U5015 ( .A1(n4786), .A2(n5289), .ZN(n4785) );
  AND2_X1 U5016 ( .A1(n5808), .A2(n4793), .ZN(n4791) );
  AND2_X1 U5017 ( .A1(n4794), .A2(n5809), .ZN(n4789) );
  AND2_X1 U5018 ( .A1(n5127), .A2(n5796), .ZN(n4911) );
  AND2_X1 U5019 ( .A1(n4792), .A2(n5810), .ZN(n4788) );
  INV_X1 U5020 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5810) );
  INV_X1 U5021 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n5809) );
  INV_X1 U5022 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n5808) );
  INV_X1 U5023 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n4794) );
  INV_X1 U5024 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n4793) );
  INV_X1 U5025 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n6115) );
  NOR2_X1 U5026 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n5812) );
  NOR2_X1 U5027 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), .ZN(
        n5813) );
  INV_X1 U5028 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n6411) );
  INV_X1 U5029 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n6425) );
  INV_X1 U5030 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n6422) );
  INV_X1 U5031 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n6418) );
  NOR2_X1 U5032 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .ZN(
        n4527) );
  NOR2_X1 U5033 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n4526) );
  NOR2_X1 U5034 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n4525) );
  INV_X1 U5035 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n4696) );
  INV_X1 U5036 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n5822) );
  INV_X4 U5037 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  INV_X1 U5038 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5796) );
  AND2_X1 U5039 ( .A1(n4390), .A2(n6891), .ZN(n5999) );
  OAI21_X2 U5040 ( .B1(n8956), .B2(n8952), .A(n6629), .ZN(n8882) );
  OAI21_X2 U5041 ( .B1(n7198), .B2(n7194), .A(n7195), .ZN(n7351) );
  XNOR2_X1 U5042 ( .A(n6481), .B(n6547), .ZN(n7352) );
  INV_X1 U5043 ( .A(n4387), .ZN(n4396) );
  OR2_X1 U5044 ( .A1(n9346), .A2(n6706), .ZN(n5731) );
  INV_X1 U5045 ( .A(n9183), .ZN(n8110) );
  NAND2_X1 U5046 ( .A1(n5331), .A2(n5330), .ZN(n5045) );
  AND2_X1 U5047 ( .A1(n5119), .A2(n4767), .ZN(n4766) );
  INV_X1 U5048 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n4767) );
  AOI21_X1 U5049 ( .B1(n4398), .B2(n8609), .A(n4440), .ZN(n4938) );
  OR2_X1 U5050 ( .A1(n8795), .A2(n8230), .ZN(n6385) );
  NAND2_X1 U5051 ( .A1(n5163), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n5202) );
  INV_X1 U5052 ( .A(n5227), .ZN(n5163) );
  INV_X1 U5053 ( .A(n5542), .ZN(n5302) );
  INV_X1 U5054 ( .A(n9156), .ZN(n9126) );
  NAND2_X1 U5055 ( .A1(n6085), .A2(n6084), .ZN(n6101) );
  AOI21_X1 U5056 ( .B1(n5663), .B2(n5662), .A(n4608), .ZN(n4607) );
  NAND2_X1 U5057 ( .A1(n8064), .A2(n7399), .ZN(n4608) );
  NAND2_X1 U5058 ( .A1(n4552), .A2(n4551), .ZN(n6184) );
  NAND2_X1 U5059 ( .A1(n6183), .A2(n6288), .ZN(n4551) );
  NAND2_X1 U5060 ( .A1(n4553), .A2(n6315), .ZN(n4552) );
  NOR2_X1 U5061 ( .A1(n5676), .A2(n5675), .ZN(n4605) );
  AND2_X1 U5062 ( .A1(n8078), .A2(n7399), .ZN(n4611) );
  NAND2_X1 U5063 ( .A1(n5695), .A2(n9164), .ZN(n4610) );
  OAI21_X1 U5064 ( .B1(n5693), .B2(n5692), .A(n5691), .ZN(n4612) );
  OR2_X1 U5065 ( .A1(n8753), .A2(n6921), .ZN(n6314) );
  INV_X1 U5066 ( .A(n6324), .ZN(n4724) );
  OR2_X1 U5067 ( .A1(n8768), .A2(n8339), .ZN(n6393) );
  NOR2_X1 U5068 ( .A1(n5729), .A2(n4604), .ZN(n4603) );
  AND2_X1 U5069 ( .A1(n5720), .A2(n4965), .ZN(n5777) );
  NAND2_X1 U5070 ( .A1(n5019), .A2(n5018), .ZN(n5022) );
  NOR2_X1 U5071 ( .A1(n5017), .A2(n4839), .ZN(n4838) );
  INV_X1 U5072 ( .A(n5014), .ZN(n4839) );
  NAND2_X1 U5073 ( .A1(n6314), .A2(n6311), .ZN(n6400) );
  NAND2_X1 U5074 ( .A1(n8753), .A2(n6921), .ZN(n6403) );
  NOR2_X1 U5075 ( .A1(n6263), .A2(n6392), .ZN(n8493) );
  OR2_X1 U5076 ( .A1(n8783), .A2(n8263), .ZN(n6389) );
  OR2_X1 U5077 ( .A1(n8745), .A2(n8719), .ZN(n6376) );
  NOR2_X1 U5078 ( .A1(n5824), .A2(n5823), .ZN(n5825) );
  NOR2_X1 U5079 ( .A1(n6086), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n6102) );
  INV_X1 U5080 ( .A(n9442), .ZN(n5166) );
  OR2_X1 U5081 ( .A1(n9336), .A2(n5172), .ZN(n5726) );
  NOR2_X1 U5082 ( .A1(n9125), .A2(n4597), .ZN(n4596) );
  INV_X1 U5083 ( .A(n8085), .ZN(n4597) );
  OR2_X1 U5084 ( .A1(n9371), .A2(n9215), .ZN(n8078) );
  OR2_X1 U5085 ( .A1(n9388), .A2(n9269), .ZN(n4627) );
  AND2_X1 U5086 ( .A1(n7494), .A2(n9086), .ZN(n6668) );
  AND2_X1 U5087 ( .A1(n5093), .A2(n5092), .ZN(n5187) );
  NAND2_X1 U5088 ( .A1(n5237), .A2(n5080), .ZN(n5208) );
  AOI21_X1 U5089 ( .B1(n4854), .B2(n4856), .A(n4851), .ZN(n4850) );
  INV_X1 U5090 ( .A(n4546), .ZN(n4545) );
  OAI21_X1 U5091 ( .B1(n4549), .B2(n4547), .A(n5038), .ZN(n4546) );
  NAND2_X1 U5092 ( .A1(n4548), .A2(n5033), .ZN(n4547) );
  NAND2_X1 U5093 ( .A1(n5038), .A2(n5037), .ZN(n5341) );
  AOI21_X1 U5094 ( .B1(n4846), .B2(n4848), .A(n4844), .ZN(n4843) );
  INV_X1 U5095 ( .A(n4964), .ZN(n4844) );
  NAND2_X1 U5096 ( .A1(n4992), .A2(n4991), .ZN(n5435) );
  XNOR2_X1 U5097 ( .A(n4986), .B(SI_4_), .ZN(n5410) );
  INV_X1 U5098 ( .A(n5399), .ZN(n4981) );
  INV_X1 U5099 ( .A(n4812), .ZN(n4486) );
  NAND2_X1 U5100 ( .A1(n8249), .A2(n6787), .ZN(n4814) );
  NOR2_X1 U5101 ( .A1(n6819), .A2(n7662), .ZN(n4490) );
  INV_X1 U5102 ( .A(n5992), .ZN(n5890) );
  INV_X1 U5103 ( .A(n5991), .ZN(n5931) );
  NOR2_X1 U5104 ( .A1(n8423), .A2(n8424), .ZN(n8430) );
  NAND2_X1 U5105 ( .A1(n6389), .A2(n6326), .ZN(n8591) );
  NAND2_X1 U5106 ( .A1(n4518), .A2(n4436), .ZN(n8626) );
  NOR2_X1 U5107 ( .A1(n8800), .A2(n8652), .ZN(n8487) );
  AOI21_X1 U5108 ( .B1(n4932), .B2(n4930), .A(n4444), .ZN(n4929) );
  INV_X1 U5109 ( .A(n8482), .ZN(n4930) );
  NAND2_X1 U5110 ( .A1(n5839), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6091) );
  INV_X1 U5111 ( .A(n6074), .ZN(n5839) );
  XNOR2_X1 U5112 ( .A(n5854), .B(P2_IR_REG_29__SCAN_IN), .ZN(n5855) );
  OR2_X1 U5113 ( .A1(n5853), .A2(n6416), .ZN(n5854) );
  NOR2_X1 U5114 ( .A1(n5829), .A2(P2_IR_REG_28__SCAN_IN), .ZN(n5853) );
  NAND2_X1 U5115 ( .A1(n4827), .A2(n5816), .ZN(n4826) );
  INV_X1 U5116 ( .A(n4828), .ZN(n4827) );
  NAND2_X1 U5117 ( .A1(n6437), .A2(n6433), .ZN(n7118) );
  INV_X1 U5118 ( .A(n4885), .ZN(n4884) );
  OAI21_X1 U5119 ( .B1(n9108), .B2(n4886), .A(n4446), .ZN(n4885) );
  NAND2_X1 U5120 ( .A1(n8112), .A2(n4891), .ZN(n4886) );
  AND2_X1 U5121 ( .A1(n5731), .A2(n5730), .ZN(n8112) );
  NOR2_X1 U5122 ( .A1(n9108), .A2(n4888), .ZN(n4887) );
  INV_X1 U5123 ( .A(n4891), .ZN(n4888) );
  NAND2_X1 U5124 ( .A1(n4904), .A2(n4903), .ZN(n9133) );
  AOI21_X1 U5125 ( .B1(n4905), .B2(n4400), .A(n4452), .ZN(n4903) );
  NOR2_X1 U5126 ( .A1(n8109), .A2(n4908), .ZN(n4907) );
  AND2_X1 U5127 ( .A1(n9363), .A2(n9183), .ZN(n8109) );
  INV_X1 U5128 ( .A(n8107), .ZN(n4908) );
  NAND2_X1 U5129 ( .A1(n9269), .A2(n9286), .ZN(n4923) );
  NAND2_X1 U5130 ( .A1(n7959), .A2(n4706), .ZN(n9825) );
  AND2_X1 U5131 ( .A1(n9827), .A2(n7958), .ZN(n4706) );
  NAND2_X1 U5132 ( .A1(n4438), .A2(n7878), .ZN(n4581) );
  INV_X1 U5133 ( .A(n9963), .ZN(n9844) );
  AND2_X1 U5134 ( .A1(n6673), .A2(n6672), .ZN(n7365) );
  OAI21_X1 U5135 ( .B1(n5136), .B2(P1_IR_REG_29__SCAN_IN), .A(n5135), .ZN(
        n5165) );
  OAI21_X1 U5136 ( .B1(n5069), .B2(n4874), .A(n4872), .ZN(n5237) );
  INV_X1 U5137 ( .A(n4873), .ZN(n4872) );
  OAI21_X1 U5138 ( .B1(n4875), .B2(n4874), .A(n5234), .ZN(n4873) );
  INV_X1 U5139 ( .A(n5074), .ZN(n4874) );
  NAND2_X1 U5140 ( .A1(n6651), .A2(n6653), .ZN(n6654) );
  INV_X1 U5141 ( .A(n6652), .ZN(n6653) );
  NAND2_X1 U5142 ( .A1(n5196), .A2(n5195), .ZN(n9156) );
  INV_X1 U5143 ( .A(n9086), .ZN(n9250) );
  NAND2_X1 U5144 ( .A1(n5636), .A2(n4602), .ZN(n4601) );
  NAND2_X1 U5145 ( .A1(n4683), .A2(n4682), .ZN(n4681) );
  NAND2_X1 U5146 ( .A1(n4680), .A2(n4679), .ZN(n4678) );
  NOR2_X1 U5147 ( .A1(n6099), .A2(n6315), .ZN(n4682) );
  OAI21_X1 U5148 ( .B1(n5664), .B2(n7399), .A(n4606), .ZN(n5672) );
  INV_X1 U5149 ( .A(n4605), .ZN(n5682) );
  NAND2_X1 U5150 ( .A1(n4677), .A2(n4676), .ZN(n6227) );
  OAI21_X1 U5151 ( .B1(n4671), .B2(n4670), .A(n4668), .ZN(n6220) );
  AND2_X1 U5152 ( .A1(n6224), .A2(n6288), .ZN(n4542) );
  AOI21_X1 U5153 ( .B1(n4689), .B2(n4429), .A(n6262), .ZN(n4686) );
  OAI21_X1 U5154 ( .B1(n4543), .B2(n4539), .A(n4690), .ZN(n4689) );
  NAND2_X1 U5155 ( .A1(n4685), .A2(n8539), .ZN(n4684) );
  INV_X1 U5156 ( .A(n6270), .ZN(n4685) );
  OAI21_X1 U5157 ( .B1(n5694), .B2(n7399), .A(n4609), .ZN(n5705) );
  NOR2_X1 U5158 ( .A1(n8774), .A2(n8543), .ZN(n6263) );
  AND2_X1 U5159 ( .A1(n8774), .A2(n8543), .ZN(n6392) );
  AND2_X1 U5160 ( .A1(n10165), .A2(n4645), .ZN(n4644) );
  AOI21_X1 U5161 ( .B1(n4868), .B2(n4865), .A(n4864), .ZN(n4863) );
  INV_X1 U5162 ( .A(n5187), .ZN(n4864) );
  INV_X1 U5163 ( .A(n4870), .ZN(n4865) );
  INV_X1 U5164 ( .A(n4868), .ZN(n4866) );
  INV_X1 U5165 ( .A(n5272), .ZN(n4851) );
  NAND2_X1 U5166 ( .A1(n5035), .A2(n5034), .ZN(n5038) );
  NAND2_X1 U5167 ( .A1(n5000), .A2(n9625), .ZN(n5003) );
  OAI22_X1 U5168 ( .A1(n5831), .A2(n4973), .B1(n4975), .B2(n4974), .ZN(n4977)
         );
  NAND2_X1 U5169 ( .A1(n8238), .A2(n8237), .ZN(n4808) );
  INV_X1 U5170 ( .A(n4511), .ZN(n4510) );
  OAI21_X1 U5171 ( .B1(n4401), .B2(n8516), .A(n6396), .ZN(n4511) );
  AND2_X1 U5172 ( .A1(n9792), .A2(n4401), .ZN(n4507) );
  NAND2_X1 U5173 ( .A1(n7844), .A2(n4473), .ZN(n8393) );
  NOR2_X1 U5174 ( .A1(n8757), .A2(n8338), .ZN(n6395) );
  INV_X1 U5175 ( .A(n6271), .ZN(n4877) );
  OR2_X1 U5176 ( .A1(n8779), .A2(n8592), .ZN(n6390) );
  NOR2_X1 U5177 ( .A1(n8811), .A2(n4641), .ZN(n4640) );
  INV_X1 U5178 ( .A(n4642), .ZN(n4641) );
  AND2_X1 U5179 ( .A1(n4719), .A2(n6375), .ZN(n4516) );
  OR2_X1 U5180 ( .A1(n10178), .A2(n7947), .ZN(n6339) );
  OR2_X1 U5181 ( .A1(n8351), .A2(n10147), .ZN(n6332) );
  OR2_X1 U5182 ( .A1(n8352), .A2(n10141), .ZN(n6360) );
  NAND2_X1 U5183 ( .A1(n4943), .A2(n4942), .ZN(n6334) );
  NAND2_X1 U5184 ( .A1(n8521), .A2(n8516), .ZN(n8524) );
  NOR2_X1 U5185 ( .A1(n8602), .A2(n8783), .ZN(n8573) );
  NAND2_X1 U5186 ( .A1(n8661), .A2(n6381), .ZN(n8662) );
  AOI21_X1 U5187 ( .B1(n4717), .B2(n4716), .A(n6368), .ZN(n7923) );
  AND2_X1 U5188 ( .A1(n4410), .A2(n6369), .ZN(n4716) );
  NOR2_X1 U5189 ( .A1(n10083), .A2(n8303), .ZN(n4645) );
  NAND2_X1 U5190 ( .A1(n4644), .A2(n7743), .ZN(n7712) );
  NOR2_X1 U5191 ( .A1(n10094), .A2(n7785), .ZN(n7743) );
  AND2_X1 U5192 ( .A1(n4763), .A2(n6590), .ZN(n4762) );
  NAND2_X1 U5193 ( .A1(n8928), .A2(n4764), .ZN(n4763) );
  INV_X1 U5194 ( .A(n8928), .ZN(n4765) );
  NAND2_X1 U5195 ( .A1(n5563), .A2(n7573), .ZN(n5741) );
  INV_X1 U5196 ( .A(n4596), .ZN(n4595) );
  INV_X1 U5197 ( .A(n8086), .ZN(n4592) );
  AOI21_X1 U5198 ( .B1(n4596), .B2(n9140), .A(n8087), .ZN(n4594) );
  OR2_X1 U5199 ( .A1(n9341), .A2(n9127), .ZN(n5732) );
  NAND2_X1 U5200 ( .A1(n9175), .A2(n4623), .ZN(n4622) );
  OR2_X1 U5201 ( .A1(n9356), .A2(n5233), .ZN(n8084) );
  OR2_X1 U5202 ( .A1(n9363), .A2(n8110), .ZN(n8083) );
  AND2_X1 U5203 ( .A1(n8081), .A2(n8079), .ZN(n4702) );
  OR2_X1 U5204 ( .A1(n9366), .A2(n5249), .ZN(n8082) );
  OR2_X1 U5205 ( .A1(n4627), .A2(n9381), .ZN(n4626) );
  NAND2_X1 U5206 ( .A1(n4894), .A2(n4895), .ZN(n4893) );
  NOR2_X1 U5207 ( .A1(n8096), .A2(n4897), .ZN(n4896) );
  INV_X1 U5208 ( .A(n4902), .ZN(n4897) );
  INV_X1 U5209 ( .A(n7956), .ZN(n4901) );
  OR2_X1 U5210 ( .A1(n7991), .A2(n9845), .ZN(n5653) );
  OR2_X1 U5211 ( .A1(n7868), .A2(n9961), .ZN(n5644) );
  INV_X1 U5212 ( .A(n7635), .ZN(n4913) );
  NOR2_X1 U5213 ( .A1(n7631), .A2(n4915), .ZN(n4914) );
  INV_X1 U5214 ( .A(n7497), .ZN(n4915) );
  NAND2_X1 U5215 ( .A1(n4589), .A2(P2_DATAO_REG_7__SCAN_IN), .ZN(n4588) );
  NOR2_X1 U5216 ( .A1(n7613), .A2(n7481), .ZN(n7504) );
  OR2_X1 U5217 ( .A1(n7615), .A2(n7477), .ZN(n5624) );
  NAND2_X1 U5218 ( .A1(n7557), .A2(n7520), .ZN(n5756) );
  INV_X1 U5219 ( .A(n4911), .ZN(n4910) );
  NAND2_X1 U5220 ( .A1(n5098), .A2(n5097), .ZN(n5174) );
  NOR2_X1 U5221 ( .A1(n5258), .A2(n4876), .ZN(n4875) );
  INV_X1 U5222 ( .A(n5068), .ZN(n4876) );
  NOR2_X1 U5223 ( .A1(n4858), .A2(n4550), .ZN(n4549) );
  INV_X1 U5224 ( .A(n5028), .ZN(n4550) );
  INV_X1 U5225 ( .A(n5355), .ZN(n4858) );
  OAI21_X1 U5226 ( .B1(n5009), .B2(n4833), .A(n4554), .ZN(n5367) );
  AOI21_X1 U5227 ( .B1(n4832), .B2(n4556), .A(n4555), .ZN(n4554) );
  INV_X1 U5228 ( .A(n5022), .ZN(n4555) );
  AOI21_X1 U5229 ( .B1(n4836), .B2(n4838), .A(n4449), .ZN(n4835) );
  INV_X1 U5230 ( .A(n4962), .ZN(n4836) );
  NOR2_X1 U5231 ( .A1(n4837), .A2(n4558), .ZN(n4557) );
  INV_X1 U5232 ( .A(n5008), .ZN(n4558) );
  INV_X1 U5233 ( .A(n4838), .ZN(n4837) );
  NAND2_X1 U5234 ( .A1(n5009), .A2(n5008), .ZN(n5518) );
  INV_X1 U5235 ( .A(n4847), .ZN(n4846) );
  OAI21_X1 U5236 ( .B1(n4848), .B2(n4997), .A(n5003), .ZN(n4847) );
  NAND2_X1 U5237 ( .A1(n4849), .A2(n4999), .ZN(n4848) );
  INV_X1 U5238 ( .A(n5480), .ZN(n4849) );
  INV_X1 U5239 ( .A(n5502), .ZN(n4997) );
  XNOR2_X1 U5240 ( .A(n4998), .B(SI_7_), .ZN(n5502) );
  NAND2_X1 U5241 ( .A1(n4996), .A2(n4995), .ZN(n5501) );
  INV_X1 U5242 ( .A(n5434), .ZN(n4993) );
  XNOR2_X1 U5243 ( .A(n4994), .B(SI_6_), .ZN(n5434) );
  INV_X1 U5244 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4714) );
  NOR2_X1 U5245 ( .A1(n8311), .A2(n4810), .ZN(n4809) );
  NAND2_X1 U5246 ( .A1(n8172), .A2(n6782), .ZN(n8176) );
  AOI21_X1 U5247 ( .B1(n4805), .B2(n4806), .A(n4804), .ZN(n4803) );
  INV_X1 U5248 ( .A(n8210), .ZN(n4804) );
  INV_X1 U5249 ( .A(n4809), .ZN(n4805) );
  NOR2_X1 U5250 ( .A1(n4823), .A2(n4484), .ZN(n4483) );
  INV_X1 U5251 ( .A(n6765), .ZN(n4484) );
  INV_X1 U5252 ( .A(n4824), .ZN(n4823) );
  NOR2_X1 U5253 ( .A1(n7283), .A2(n4820), .ZN(n4819) );
  INV_X1 U5254 ( .A(n6735), .ZN(n4820) );
  AOI21_X1 U5255 ( .B1(n7655), .B2(n7654), .A(n6759), .ZN(n7822) );
  AND2_X1 U5256 ( .A1(n8141), .A2(n8136), .ZN(n4812) );
  NAND2_X1 U5257 ( .A1(n8194), .A2(n8132), .ZN(n8201) );
  AND2_X1 U5258 ( .A1(n6814), .A2(n6792), .ZN(n4813) );
  NAND2_X1 U5259 ( .A1(n4667), .A2(n6312), .ZN(n4666) );
  MUX2_X1 U5260 ( .A(n6400), .B(n6352), .S(n6315), .Z(n6312) );
  AND4_X1 U5261 ( .A1(n5894), .A2(n5893), .A3(n5892), .A4(n5891), .ZN(n8230)
         );
  AND4_X1 U5262 ( .A1(n6207), .A2(n6206), .A3(n6205), .A4(n6204), .ZN(n8229)
         );
  NAND2_X1 U5263 ( .A1(n8850), .A2(n5855), .ZN(n6202) );
  NOR2_X1 U5264 ( .A1(n9749), .A2(n9750), .ZN(n9748) );
  NOR2_X1 U5265 ( .A1(n9748), .A2(n4573), .ZN(n6972) );
  AND2_X1 U5266 ( .A1(n9752), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n4573) );
  OR2_X1 U5267 ( .A1(n6972), .A2(n6971), .ZN(n4572) );
  INV_X1 U5268 ( .A(n8374), .ZN(n4565) );
  AOI21_X1 U5269 ( .B1(n8374), .B2(n4564), .A(n4469), .ZN(n4563) );
  INV_X1 U5270 ( .A(n6937), .ZN(n4564) );
  XNOR2_X1 U5271 ( .A(n8393), .B(n8394), .ZN(n7846) );
  NOR2_X1 U5272 ( .A1(n7846), .A2(n9801), .ZN(n8395) );
  NAND2_X1 U5273 ( .A1(n8421), .A2(n8422), .ZN(n8423) );
  NAND2_X1 U5274 ( .A1(n8434), .A2(n8433), .ZN(n8442) );
  NAND2_X1 U5275 ( .A1(n5870), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6319) );
  NAND2_X1 U5276 ( .A1(n8445), .A2(n8446), .ZN(n8449) );
  NOR2_X1 U5277 ( .A1(n6395), .A2(n6394), .ZN(n8499) );
  NAND2_X1 U5278 ( .A1(n8524), .A2(n6324), .ZN(n8502) );
  OR2_X1 U5279 ( .A1(n8768), .A2(n8495), .ZN(n8496) );
  NOR2_X1 U5280 ( .A1(n8774), .A2(n8574), .ZN(n8551) );
  NAND2_X1 U5281 ( .A1(n8661), .A2(n4434), .ZN(n4518) );
  INV_X1 U5282 ( .A(n4727), .ZN(n4519) );
  INV_X1 U5283 ( .A(n4726), .ZN(n4725) );
  OAI21_X1 U5284 ( .B1(n4419), .B2(n4727), .A(n6384), .ZN(n4726) );
  OR2_X1 U5285 ( .A1(n8805), .A2(n8229), .ZN(n6383) );
  AND2_X1 U5286 ( .A1(n8699), .A2(n4639), .ZN(n8644) );
  AND2_X1 U5287 ( .A1(n8648), .A2(n4640), .ZN(n4639) );
  OR2_X1 U5288 ( .A1(n8811), .A2(n8687), .ZN(n8483) );
  NAND2_X1 U5289 ( .A1(n8699), .A2(n4642), .ZN(n8677) );
  NAND2_X1 U5290 ( .A1(n6136), .A2(n6135), .ZN(n8745) );
  OR2_X1 U5291 ( .A1(n4722), .A2(n4720), .ZN(n4719) );
  INV_X1 U5292 ( .A(n4464), .ZN(n4720) );
  AND2_X1 U5293 ( .A1(n4464), .A2(n4945), .ZN(n4721) );
  NOR2_X1 U5294 ( .A1(n4948), .A2(n4723), .ZN(n4722) );
  INV_X1 U5295 ( .A(n6374), .ZN(n4723) );
  INV_X1 U5296 ( .A(n6106), .ZN(n5840) );
  NAND2_X1 U5297 ( .A1(n7997), .A2(n7996), .ZN(n8028) );
  OR2_X1 U5298 ( .A1(n7950), .A2(n8020), .ZN(n7857) );
  OR2_X1 U5299 ( .A1(n6055), .A2(n5838), .ZN(n6074) );
  NAND2_X1 U5300 ( .A1(n5926), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n6030) );
  AND2_X1 U5301 ( .A1(n7245), .A2(n6717), .ZN(n10089) );
  OR2_X1 U5302 ( .A1(n8857), .A2(n7233), .ZN(n10070) );
  INV_X1 U5303 ( .A(n8684), .ZN(n10072) );
  INV_X1 U5304 ( .A(n7895), .ZN(n7892) );
  NAND2_X1 U5305 ( .A1(n7893), .A2(n7892), .ZN(n7891) );
  OR2_X1 U5306 ( .A1(n9806), .A2(n6819), .ZN(n7229) );
  AND2_X1 U5307 ( .A1(n6927), .A2(n8857), .ZN(n8684) );
  NAND2_X1 U5308 ( .A1(n5886), .A2(n5885), .ZN(n8795) );
  NAND2_X1 U5309 ( .A1(n6209), .A2(n6208), .ZN(n8800) );
  NAND2_X1 U5310 ( .A1(n6174), .A2(n6173), .ZN(n8815) );
  NAND2_X1 U5311 ( .A1(n8059), .A2(n6818), .ZN(n9806) );
  AND2_X1 U5312 ( .A1(n6322), .A2(n7662), .ZN(n6818) );
  NAND2_X1 U5313 ( .A1(n7662), .A2(n7552), .ZN(n10123) );
  INV_X1 U5314 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5849) );
  NAND2_X1 U5315 ( .A1(n8846), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4950) );
  AND2_X1 U5316 ( .A1(n5819), .A2(n4498), .ZN(n4499) );
  AND2_X1 U5317 ( .A1(n5862), .A2(n4500), .ZN(n4498) );
  INV_X1 U5318 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n4500) );
  NAND2_X1 U5319 ( .A1(n5867), .A2(n4831), .ZN(n4830) );
  INV_X1 U5320 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n4831) );
  NOR2_X1 U5321 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n5864) );
  CLKBUF_X1 U5322 ( .A(n5921), .Z(n5922) );
  INV_X1 U5323 ( .A(n8917), .ZN(n4521) );
  NAND2_X1 U5324 ( .A1(n4779), .A2(n4777), .ZN(n7585) );
  NOR2_X1 U5325 ( .A1(n7587), .A2(n4778), .ZN(n4777) );
  INV_X1 U5326 ( .A(n4780), .ZN(n4778) );
  AOI21_X1 U5327 ( .B1(n6458), .B2(n7521), .A(n4743), .ZN(n4742) );
  NAND2_X1 U5328 ( .A1(n8893), .A2(n4775), .ZN(n4773) );
  OR2_X1 U5329 ( .A1(n8890), .A2(n8891), .ZN(n4775) );
  NOR2_X1 U5330 ( .A1(n4749), .A2(n4748), .ZN(n4747) );
  INV_X1 U5331 ( .A(n8883), .ZN(n4748) );
  NAND2_X1 U5332 ( .A1(n8909), .A2(n4757), .ZN(n4756) );
  INV_X1 U5333 ( .A(n6639), .ZN(n4757) );
  AND2_X1 U5334 ( .A1(n4413), .A2(n8978), .ZN(n4759) );
  AND2_X1 U5335 ( .A1(n9442), .A2(n9447), .ZN(n5452) );
  NAND2_X1 U5336 ( .A1(n6846), .A2(n6845), .ZN(n4664) );
  NAND2_X1 U5337 ( .A1(n4664), .A2(n4663), .ZN(n4662) );
  NAND2_X1 U5338 ( .A1(n7034), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n4663) );
  AND2_X1 U5339 ( .A1(n7094), .A2(n9908), .ZN(n9916) );
  NOR2_X1 U5340 ( .A1(n9914), .A2(n4659), .ZN(n7099) );
  AND2_X1 U5341 ( .A1(n7095), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n4659) );
  NOR2_X1 U5342 ( .A1(n7098), .A2(n7099), .ZN(n7218) );
  NAND2_X1 U5343 ( .A1(n9933), .A2(n9934), .ZN(n9932) );
  OR2_X1 U5344 ( .A1(n7222), .A2(n7221), .ZN(n4658) );
  AND2_X1 U5345 ( .A1(n4658), .A2(n4657), .ZN(n7309) );
  NAND2_X1 U5346 ( .A1(n7306), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n4657) );
  OR2_X1 U5347 ( .A1(n7309), .A2(n7308), .ZN(n4656) );
  OR2_X1 U5348 ( .A1(n7919), .A2(n7918), .ZN(n4653) );
  OR2_X1 U5349 ( .A1(n5202), .A2(n5164), .ZN(n8115) );
  AND2_X1 U5350 ( .A1(n8118), .A2(n9110), .ZN(n9098) );
  NOR2_X1 U5351 ( .A1(n9341), .A2(n9118), .ZN(n9110) );
  NAND2_X1 U5352 ( .A1(n4619), .A2(n4618), .ZN(n9134) );
  AND2_X1 U5353 ( .A1(n8083), .A2(n5569), .ZN(n9164) );
  OR2_X1 U5354 ( .A1(n9366), .A2(n9203), .ZN(n8106) );
  NOR2_X1 U5355 ( .A1(n4922), .A2(n4921), .ZN(n4920) );
  NOR2_X1 U5356 ( .A1(n8102), .A2(n9264), .ZN(n4921) );
  NOR2_X1 U5357 ( .A1(n8103), .A2(n4923), .ZN(n4922) );
  NAND2_X1 U5358 ( .A1(n9263), .A2(n8072), .ZN(n9242) );
  AND2_X1 U5359 ( .A1(n5679), .A2(n8073), .ZN(n9243) );
  NAND2_X1 U5360 ( .A1(n5311), .A2(n5310), .ZN(n9269) );
  OR2_X1 U5361 ( .A1(n9255), .A2(n9258), .ZN(n4924) );
  NOR2_X1 U5362 ( .A1(n9319), .A2(n9405), .ZN(n9300) );
  OR2_X1 U5363 ( .A1(n5362), .A2(n5348), .ZN(n5350) );
  NAND2_X1 U5364 ( .A1(n9310), .A2(n8066), .ZN(n4701) );
  AND2_X1 U5365 ( .A1(n7961), .A2(n7960), .ZN(n4705) );
  AND2_X1 U5366 ( .A1(n8064), .A2(n5657), .ZN(n7961) );
  NAND2_X1 U5367 ( .A1(n7877), .A2(n4417), .ZN(n4577) );
  INV_X1 U5368 ( .A(n4579), .ZN(n4578) );
  OAI21_X1 U5369 ( .B1(n4580), .B2(n4417), .A(n7880), .ZN(n4579) );
  INV_X1 U5370 ( .A(n4581), .ZN(n4580) );
  NOR2_X1 U5371 ( .A1(n7639), .A2(n4704), .ZN(n4703) );
  INV_X1 U5372 ( .A(n5464), .ZN(n5535) );
  INV_X1 U5373 ( .A(n5388), .ZN(n5534) );
  INV_X1 U5374 ( .A(n9016), .ZN(n7558) );
  NAND2_X1 U5375 ( .A1(n7379), .A2(n7378), .ZN(n9963) );
  INV_X1 U5376 ( .A(n9960), .ZN(n9285) );
  NAND2_X1 U5377 ( .A1(n6668), .A2(n6434), .ZN(n7416) );
  NAND2_X1 U5378 ( .A1(n5152), .A2(n5151), .ZN(n9336) );
  NAND2_X1 U5379 ( .A1(n5262), .A2(n5261), .ZN(n9371) );
  NOR2_X1 U5380 ( .A1(n7108), .A2(n7107), .ZN(n7204) );
  XNOR2_X1 U5381 ( .A(n5143), .B(SI_30_), .ZN(n8849) );
  XNOR2_X1 U5382 ( .A(n5174), .B(n5173), .ZN(n8855) );
  XNOR2_X1 U5383 ( .A(n5188), .B(n5187), .ZN(n8040) );
  NAND2_X1 U5384 ( .A1(n4862), .A2(n4868), .ZN(n5188) );
  XNOR2_X1 U5385 ( .A(n5221), .B(n5220), .ZN(n8010) );
  NAND2_X1 U5386 ( .A1(n4867), .A2(n5083), .ZN(n5221) );
  XNOR2_X1 U5387 ( .A(n5208), .B(n5209), .ZN(n7938) );
  AND2_X1 U5388 ( .A1(n5080), .A2(n5079), .ZN(n5234) );
  NAND2_X1 U5389 ( .A1(n5069), .A2(n4875), .ZN(n4960) );
  NAND3_X1 U5390 ( .A1(n4422), .A2(n5475), .A3(n4959), .ZN(n5558) );
  NAND2_X1 U5391 ( .A1(n4853), .A2(n5053), .ZN(n5284) );
  XNOR2_X1 U5392 ( .A(n5435), .B(n5434), .ZN(n5960) );
  INV_X1 U5393 ( .A(n5410), .ZN(n4985) );
  NAND3_X1 U5394 ( .A1(n8158), .A2(n4491), .A3(n4954), .ZN(n8241) );
  OR2_X1 U5395 ( .A1(n8261), .A2(n8265), .ZN(n4954) );
  OAI21_X1 U5396 ( .B1(n7822), .B2(n4482), .A(n4479), .ZN(n8017) );
  INV_X1 U5397 ( .A(n4483), .ZN(n4482) );
  AND2_X1 U5398 ( .A1(n4480), .A2(n4821), .ZN(n4479) );
  AOI21_X1 U5399 ( .B1(n4824), .B2(n4822), .A(n4426), .ZN(n4821) );
  AND4_X1 U5400 ( .A1(n6156), .A2(n6155), .A3(n6154), .A4(n6153), .ZN(n8737)
         );
  NOR2_X1 U5401 ( .A1(n4538), .A2(n6926), .ZN(n4536) );
  XNOR2_X1 U5402 ( .A(n6354), .B(n8668), .ZN(n6355) );
  NAND2_X1 U5403 ( .A1(n4497), .A2(n6407), .ZN(n4494) );
  OAI21_X1 U5404 ( .B1(n6959), .B2(n6948), .A(n8366), .ZN(n6998) );
  XOR2_X1 U5405 ( .A(n8447), .B(n8442), .Z(n8435) );
  NAND2_X1 U5406 ( .A1(n4941), .A2(n4398), .ZN(n8584) );
  AND2_X1 U5407 ( .A1(n5880), .A2(n5879), .ZN(n8607) );
  NAND2_X1 U5408 ( .A1(n6152), .A2(n6151), .ZN(n8825) );
  NAND2_X1 U5409 ( .A1(n5201), .A2(n5200), .ZN(n9346) );
  NAND2_X1 U5410 ( .A1(n8055), .A2(n4613), .ZN(n5201) );
  INV_X1 U5411 ( .A(n6456), .ZN(n4769) );
  OR2_X1 U5412 ( .A1(n8862), .A2(n6688), .ZN(n6660) );
  INV_X1 U5413 ( .A(n9008), .ZN(n9845) );
  INV_X1 U5414 ( .A(n9017), .ZN(n7514) );
  NAND2_X1 U5415 ( .A1(n6703), .A2(n7043), .ZN(n8992) );
  AND2_X1 U5416 ( .A1(n5791), .A2(n5790), .ZN(n5792) );
  NAND2_X1 U5417 ( .A1(n5207), .A2(n5206), .ZN(n9142) );
  NAND2_X1 U5418 ( .A1(n5219), .A2(n5218), .ZN(n9183) );
  OR2_X1 U5419 ( .A1(n9171), .A2(n5302), .ZN(n5219) );
  NAND2_X1 U5420 ( .A1(n8113), .A2(n4884), .ZN(n4883) );
  AOI21_X1 U5421 ( .B1(n9117), .B2(n4406), .A(n4880), .ZN(n4879) );
  AND2_X1 U5422 ( .A1(n4586), .A2(n4585), .ZN(n9338) );
  INV_X1 U5423 ( .A(n8092), .ZN(n4585) );
  NAND2_X1 U5424 ( .A1(n8093), .A2(n9963), .ZN(n4586) );
  OAI21_X1 U5425 ( .B1(n9127), .B2(n9959), .A(n8091), .ZN(n8092) );
  NAND2_X1 U5426 ( .A1(n9141), .A2(n8085), .ZN(n9124) );
  OR2_X1 U5427 ( .A1(n10034), .A2(n6692), .ZN(n9249) );
  MUX2_X1 U5428 ( .A(n5943), .B(n5942), .S(n6315), .Z(n6023) );
  OAI211_X1 U5429 ( .C1(n4600), .C2(n5642), .A(n7640), .B(n5641), .ZN(n5649)
         );
  OAI21_X1 U5430 ( .B1(n4600), .B2(n7639), .A(n7642), .ZN(n5640) );
  NAND2_X1 U5431 ( .A1(n6101), .A2(n6098), .ZN(n4680) );
  NOR2_X1 U5432 ( .A1(n6097), .A2(n6288), .ZN(n4679) );
  NAND2_X1 U5433 ( .A1(n6101), .A2(n6100), .ZN(n4683) );
  NAND2_X1 U5434 ( .A1(n8660), .A2(n6379), .ZN(n4553) );
  MUX2_X1 U5435 ( .A(n4464), .B(n6132), .S(n6315), .Z(n6146) );
  NOR2_X1 U5436 ( .A1(n6184), .A2(n4448), .ZN(n4673) );
  NOR2_X1 U5437 ( .A1(n6184), .A2(n6185), .ZN(n4672) );
  INV_X1 U5438 ( .A(n6158), .ZN(n4671) );
  AOI21_X1 U5439 ( .B1(n4672), .B2(n6329), .A(n4669), .ZN(n4668) );
  OR2_X1 U5440 ( .A1(n4675), .A2(n4674), .ZN(n4669) );
  NAND2_X1 U5441 ( .A1(n6382), .A2(n6328), .ZN(n4674) );
  AND2_X1 U5442 ( .A1(n6329), .A2(n6196), .ZN(n4675) );
  NAND2_X1 U5443 ( .A1(n6329), .A2(n4673), .ZN(n4670) );
  OAI21_X1 U5444 ( .B1(n5684), .B2(n4699), .A(n5681), .ZN(n5686) );
  NAND2_X1 U5445 ( .A1(n6232), .A2(n6389), .ZN(n4543) );
  AOI21_X1 U5446 ( .B1(n4442), .B2(n4541), .A(n4540), .ZN(n4539) );
  NOR2_X1 U5447 ( .A1(n6387), .A2(n6288), .ZN(n4540) );
  NAND2_X1 U5448 ( .A1(n6223), .A2(n6315), .ZN(n4541) );
  INV_X1 U5449 ( .A(n4691), .ZN(n4690) );
  OAI21_X1 U5450 ( .B1(n6233), .B2(n6315), .A(n6326), .ZN(n4691) );
  NAND2_X1 U5451 ( .A1(n4688), .A2(n6288), .ZN(n4687) );
  INV_X1 U5452 ( .A(n6326), .ZN(n4688) );
  NOR3_X1 U5453 ( .A1(n6284), .A2(n6283), .A3(n6282), .ZN(n6286) );
  NOR2_X1 U5454 ( .A1(n4686), .A2(n4684), .ZN(n6284) );
  INV_X1 U5455 ( .A(n5730), .ZN(n4604) );
  INV_X1 U5456 ( .A(n5341), .ZN(n4548) );
  INV_X1 U5457 ( .A(n5506), .ZN(n4841) );
  INV_X1 U5458 ( .A(n4557), .ZN(n4556) );
  OAI21_X1 U5459 ( .B1(n5831), .B2(n4694), .A(n4693), .ZN(n4982) );
  NAND2_X1 U5460 ( .A1(n5831), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n4693) );
  NAND2_X1 U5461 ( .A1(n6402), .A2(n6401), .ZN(n6404) );
  NOR2_X1 U5462 ( .A1(n4633), .A2(n4635), .ZN(n4632) );
  INV_X1 U5463 ( .A(n4634), .ZN(n4633) );
  NOR2_X1 U5464 ( .A1(n8763), .A2(n8768), .ZN(n4634) );
  AND2_X1 U5465 ( .A1(n8663), .A2(n8660), .ZN(n6381) );
  OR2_X1 U5466 ( .A1(n8635), .A2(n4728), .ZN(n4727) );
  INV_X1 U5467 ( .A(n6383), .ZN(n4728) );
  INV_X1 U5468 ( .A(n4929), .ZN(n4927) );
  AND2_X1 U5469 ( .A1(n8805), .A2(n8486), .ZN(n4934) );
  NOR2_X1 U5470 ( .A1(n8815), .A2(n8822), .ZN(n4642) );
  OR2_X1 U5471 ( .A1(n8822), .A2(n8718), .ZN(n6379) );
  NOR2_X1 U5472 ( .A1(n8023), .A2(n7950), .ZN(n4638) );
  OR2_X1 U5473 ( .A1(n7701), .A2(n6366), .ZN(n4718) );
  OR2_X1 U5474 ( .A1(n10069), .A2(n4503), .ZN(n4502) );
  OR2_X1 U5475 ( .A1(n10077), .A2(n10068), .ZN(n4503) );
  AND2_X1 U5476 ( .A1(n7242), .A2(n6333), .ZN(n6363) );
  NAND2_X1 U5477 ( .A1(n7237), .A2(n7895), .ZN(n4477) );
  AND2_X1 U5478 ( .A1(n6429), .A2(n6819), .ZN(n6927) );
  OR2_X1 U5479 ( .A1(n8815), .A2(n8698), .ZN(n8660) );
  NOR2_X1 U5480 ( .A1(n7814), .A2(n10178), .ZN(n7931) );
  NAND3_X1 U5481 ( .A1(n4644), .A2(n10171), .A3(n7743), .ZN(n7814) );
  AND2_X1 U5482 ( .A1(n7899), .A2(n10136), .ZN(n7900) );
  NOR2_X1 U5483 ( .A1(n5818), .A2(n5817), .ZN(n5819) );
  NOR2_X1 U5484 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n5862) );
  AND2_X1 U5485 ( .A1(n5819), .A2(n5862), .ZN(n5820) );
  OR2_X1 U5486 ( .A1(n5871), .A2(P2_IR_REG_21__SCAN_IN), .ZN(n6413) );
  NAND2_X1 U5487 ( .A1(n6413), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6408) );
  AND3_X1 U5488 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n5423) );
  AND2_X1 U5489 ( .A1(n4656), .A2(n4655), .ZN(n7915) );
  NAND2_X1 U5490 ( .A1(n7600), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n4655) );
  NOR2_X1 U5491 ( .A1(n9154), .A2(n4906), .ZN(n4905) );
  NOR2_X1 U5492 ( .A1(n4907), .A2(n4400), .ZN(n4906) );
  OR2_X1 U5493 ( .A1(n9378), .A2(n8960), .ZN(n5690) );
  NOR2_X1 U5494 ( .A1(n7979), .A2(n7991), .ZN(n4617) );
  OR2_X1 U5495 ( .A1(n9949), .A2(n7868), .ZN(n7883) );
  NAND2_X1 U5496 ( .A1(n5156), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n5513) );
  INV_X1 U5497 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n5468) );
  AND2_X1 U5498 ( .A1(n7959), .A2(n7958), .ZN(n9826) );
  AND2_X1 U5499 ( .A1(n7504), .A2(n7546), .ZN(n9950) );
  AND2_X1 U5500 ( .A1(n7401), .A2(n7400), .ZN(n7512) );
  NAND2_X1 U5501 ( .A1(n4861), .A2(n4859), .ZN(n5197) );
  AOI21_X1 U5502 ( .B1(n4863), .B2(n4866), .A(n4860), .ZN(n4859) );
  INV_X1 U5503 ( .A(n5093), .ZN(n4860) );
  NOR2_X1 U5504 ( .A1(n5220), .A2(n4871), .ZN(n4870) );
  INV_X1 U5505 ( .A(n5083), .ZN(n4871) );
  AOI21_X1 U5506 ( .B1(n4870), .B2(n5084), .A(n4869), .ZN(n4868) );
  INV_X1 U5507 ( .A(n5088), .ZN(n4869) );
  AND2_X1 U5508 ( .A1(n5063), .A2(n5062), .ZN(n5272) );
  NAND2_X1 U5509 ( .A1(n4857), .A2(n5053), .ZN(n4856) );
  INV_X1 U5510 ( .A(n5283), .ZN(n4857) );
  INV_X1 U5511 ( .A(n4855), .ZN(n4854) );
  OAI21_X1 U5512 ( .B1(n4856), .B2(n5051), .A(n5058), .ZN(n4855) );
  INV_X1 U5513 ( .A(n5319), .ZN(n5050) );
  INV_X1 U5514 ( .A(SI_8_), .ZN(n9625) );
  XNOR2_X1 U5515 ( .A(n4982), .B(SI_3_), .ZN(n5399) );
  INV_X1 U5516 ( .A(n5461), .ZN(n4731) );
  XNOR2_X1 U5517 ( .A(n4971), .B(SI_1_), .ZN(n5462) );
  AND2_X1 U5518 ( .A1(n6274), .A2(n8509), .ZN(n8216) );
  AND2_X1 U5519 ( .A1(n8154), .A2(n8188), .ZN(n8155) );
  OR2_X1 U5520 ( .A1(n8156), .A2(n8599), .ZN(n8154) );
  AOI21_X1 U5521 ( .B1(n4803), .B2(n4807), .A(n4468), .ZN(n4801) );
  NAND2_X1 U5522 ( .A1(n8855), .A2(n6245), .ZN(n4878) );
  NAND2_X1 U5523 ( .A1(n7830), .A2(n6768), .ZN(n4825) );
  INV_X1 U5524 ( .A(n6768), .ZN(n4822) );
  NAND2_X1 U5525 ( .A1(n4483), .A2(n4481), .ZN(n4480) );
  INV_X1 U5526 ( .A(n7821), .ZN(n4481) );
  INV_X1 U5527 ( .A(n6165), .ZN(n5842) );
  OR2_X1 U5528 ( .A1(n5889), .A2(n8189), .ZN(n5882) );
  NAND2_X1 U5529 ( .A1(n7822), .A2(n7821), .ZN(n7820) );
  OR2_X1 U5530 ( .A1(n6210), .A2(n8231), .ZN(n6212) );
  NAND2_X1 U5531 ( .A1(n4815), .A2(n4816), .ZN(n8300) );
  OAI21_X1 U5532 ( .B1(n4817), .B2(n7315), .A(n4418), .ZN(n4816) );
  INV_X1 U5533 ( .A(n7285), .ZN(n4817) );
  NOR2_X1 U5534 ( .A1(n6352), .A2(n6351), .ZN(n6353) );
  OAI21_X1 U5535 ( .B1(n4509), .B2(n4508), .A(n4506), .ZN(n6397) );
  AOI21_X1 U5536 ( .B1(n4510), .B2(n4507), .A(n4476), .ZN(n4506) );
  NAND2_X1 U5537 ( .A1(n4510), .A2(n9792), .ZN(n4508) );
  NOR2_X1 U5538 ( .A1(n6403), .A2(n8668), .ZN(n4497) );
  NAND2_X1 U5539 ( .A1(n6404), .A2(n4399), .ZN(n4495) );
  AND4_X1 U5540 ( .A1(n6060), .A2(n6059), .A3(n6058), .A4(n6057), .ZN(n7947)
         );
  OR2_X1 U5541 ( .A1(n8354), .A2(n8353), .ZN(n8356) );
  NAND2_X1 U5542 ( .A1(n4562), .A2(n4566), .ZN(n4561) );
  NAND2_X1 U5543 ( .A1(n4563), .A2(n4565), .ZN(n4562) );
  NOR2_X1 U5544 ( .A1(n6943), .A2(n6942), .ZN(n7017) );
  OR2_X1 U5545 ( .A1(n7020), .A2(n7019), .ZN(n4569) );
  AND2_X1 U5546 ( .A1(n4569), .A2(n4568), .ZN(n7138) );
  NAND2_X1 U5547 ( .A1(n7141), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n4568) );
  NOR2_X1 U5548 ( .A1(n7338), .A2(n4560), .ZN(n8386) );
  NOR2_X1 U5549 ( .A1(n7334), .A2(n7182), .ZN(n4560) );
  NAND2_X1 U5550 ( .A1(n8386), .A2(n8387), .ZN(n8385) );
  NAND2_X1 U5551 ( .A1(n8385), .A2(n4559), .ZN(n7341) );
  NAND2_X1 U5552 ( .A1(n7335), .A2(n7340), .ZN(n4559) );
  NAND2_X1 U5553 ( .A1(n7341), .A2(n7342), .ZN(n7451) );
  NOR2_X1 U5554 ( .A1(n8395), .A2(n8396), .ZN(n8399) );
  NOR2_X1 U5555 ( .A1(n8406), .A2(n8405), .ZN(n8409) );
  AND2_X1 U5556 ( .A1(n8551), .A2(n4630), .ZN(n8469) );
  NOR2_X1 U5557 ( .A1(n8470), .A2(n4631), .ZN(n4630) );
  INV_X1 U5558 ( .A(n4632), .ZN(n4631) );
  NAND2_X1 U5559 ( .A1(n8551), .A2(n4632), .ZN(n8508) );
  NAND2_X1 U5560 ( .A1(n6324), .A2(n6325), .ZN(n8522) );
  INV_X1 U5561 ( .A(n8522), .ZN(n8516) );
  AND2_X1 U5562 ( .A1(n6257), .A2(n6256), .ZN(n8543) );
  NAND2_X1 U5563 ( .A1(n8551), .A2(n8536), .ZN(n8531) );
  NAND2_X1 U5564 ( .A1(n6390), .A2(n6259), .ZN(n8569) );
  INV_X1 U5565 ( .A(n8569), .ZN(n8565) );
  AND2_X1 U5566 ( .A1(n6244), .A2(n6243), .ZN(n8592) );
  INV_X1 U5567 ( .A(n8491), .ZN(n4940) );
  OR2_X1 U5568 ( .A1(n8614), .A2(n8789), .ZN(n8602) );
  NOR2_X1 U5569 ( .A1(n6386), .A2(n4736), .ZN(n4735) );
  INV_X1 U5570 ( .A(n6385), .ZN(n4736) );
  INV_X1 U5571 ( .A(n4925), .ZN(n8631) );
  OAI21_X1 U5572 ( .B1(n8676), .B2(n4928), .A(n4926), .ZN(n4925) );
  NAND2_X1 U5573 ( .A1(n4932), .A2(n8642), .ZN(n4928) );
  AOI21_X1 U5574 ( .B1(n4927), .B2(n8642), .A(n4934), .ZN(n4926) );
  INV_X1 U5575 ( .A(n8662), .ZN(n4730) );
  INV_X1 U5576 ( .A(n6382), .ZN(n4729) );
  OR2_X1 U5577 ( .A1(n6190), .A2(n6189), .ZN(n6200) );
  AOI211_X1 U5578 ( .C1(n4517), .C2(n4425), .A(n4514), .B(n6377), .ZN(n8696)
         );
  NOR2_X1 U5579 ( .A1(n4515), .A2(n6376), .ZN(n4514) );
  AND2_X1 U5580 ( .A1(n8740), .A2(n8461), .ZN(n8699) );
  NAND2_X1 U5581 ( .A1(n8699), .A2(n8704), .ZN(n8700) );
  AND2_X1 U5582 ( .A1(n8825), .A2(n8479), .ZN(n8480) );
  OAI21_X1 U5583 ( .B1(n4513), .B2(n4512), .A(n6376), .ZN(n8712) );
  INV_X1 U5584 ( .A(n4516), .ZN(n4512) );
  INV_X1 U5585 ( .A(n4517), .ZN(n4513) );
  NOR2_X1 U5586 ( .A1(n8739), .A2(n8745), .ZN(n8740) );
  NAND2_X1 U5587 ( .A1(n7931), .A2(n4636), .ZN(n8739) );
  AND2_X1 U5588 ( .A1(n4402), .A2(n4637), .ZN(n4636) );
  NAND2_X1 U5589 ( .A1(n7931), .A2(n4402), .ZN(n8033) );
  AND4_X1 U5590 ( .A1(n6145), .A2(n6144), .A3(n6143), .A4(n6142), .ZN(n8719)
         );
  NAND2_X1 U5591 ( .A1(n7998), .A2(n6374), .ZN(n8030) );
  NAND2_X1 U5592 ( .A1(n7999), .A2(n4945), .ZN(n7998) );
  AND4_X1 U5593 ( .A1(n6096), .A2(n6095), .A3(n6094), .A4(n6093), .ZN(n8049)
         );
  AND2_X1 U5594 ( .A1(n7931), .A2(n4638), .ZN(n8004) );
  AND2_X1 U5595 ( .A1(n7931), .A2(n10188), .ZN(n7933) );
  NOR2_X1 U5596 ( .A1(n7923), .A2(n6371), .ZN(n7859) );
  AND4_X1 U5597 ( .A1(n5898), .A2(n5897), .A3(n5896), .A4(n5895), .ZN(n7834)
         );
  AND4_X1 U5598 ( .A1(n6079), .A2(n6078), .A3(n6077), .A4(n6076), .ZN(n8020)
         );
  NAND2_X1 U5599 ( .A1(n4717), .A2(n4718), .ZN(n7707) );
  NAND2_X1 U5600 ( .A1(n5837), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n6055) );
  AND2_X1 U5601 ( .A1(n4502), .A2(n6045), .ZN(n7683) );
  INV_X1 U5602 ( .A(n4502), .ZN(n10067) );
  AND2_X1 U5603 ( .A1(n7743), .A2(n10151), .ZN(n10079) );
  NAND2_X1 U5604 ( .A1(n7241), .A2(n6363), .ZN(n7738) );
  AND2_X1 U5605 ( .A1(n4505), .A2(n4504), .ZN(n10069) );
  NAND2_X1 U5606 ( .A1(n7738), .A2(n6364), .ZN(n4505) );
  AND2_X1 U5607 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n5926) );
  NOR2_X1 U5608 ( .A1(n7755), .A2(n6361), .ZN(n10088) );
  OR2_X1 U5609 ( .A1(n6725), .A2(n10136), .ZN(n7751) );
  AND2_X1 U5610 ( .A1(n7265), .A2(n10122), .ZN(n7899) );
  INV_X1 U5611 ( .A(n10070), .ZN(n8686) );
  OR2_X1 U5612 ( .A1(n5990), .A2(n10122), .ZN(n7772) );
  NAND2_X1 U5613 ( .A1(n7743), .A2(n4645), .ZN(n7691) );
  AND3_X1 U5614 ( .A1(n5941), .A2(n5940), .A3(n5939), .ZN(n10147) );
  NAND2_X1 U5615 ( .A1(n6410), .A2(n7247), .ZN(n10192) );
  INV_X1 U5616 ( .A(n10194), .ZN(n10126) );
  INV_X1 U5617 ( .A(n10192), .ZN(n10128) );
  XNOR2_X1 U5618 ( .A(n5826), .B(n5849), .ZN(n6930) );
  NAND2_X1 U5619 ( .A1(n5829), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5826) );
  NAND2_X1 U5620 ( .A1(n5820), .A2(n4501), .ZN(n5827) );
  AOI21_X1 U5621 ( .B1(n6319), .B2(n6318), .A(n6416), .ZN(n4787) );
  NAND2_X1 U5622 ( .A1(n4829), .A2(n5868), .ZN(n4828) );
  INV_X1 U5623 ( .A(n4830), .ZN(n4829) );
  AND2_X1 U5624 ( .A1(n4792), .A2(n5809), .ZN(n4790) );
  AND2_X1 U5625 ( .A1(n4794), .A2(n4793), .ZN(n5983) );
  OR2_X1 U5626 ( .A1(n6638), .A2(n6637), .ZN(n6639) );
  NAND2_X1 U5627 ( .A1(n5161), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n5242) );
  INV_X1 U5628 ( .A(n5265), .ZN(n5161) );
  NAND2_X1 U5629 ( .A1(n7388), .A2(n7389), .ZN(n4780) );
  OR2_X1 U5630 ( .A1(n7388), .A2(n7389), .ZN(n4781) );
  NAND2_X1 U5631 ( .A1(n6435), .A2(n7521), .ZN(n4739) );
  INV_X1 U5632 ( .A(n5297), .ZN(n5160) );
  NOR2_X1 U5633 ( .A1(n4776), .A2(n4772), .ZN(n4771) );
  INV_X1 U5634 ( .A(n4968), .ZN(n4776) );
  INV_X1 U5635 ( .A(n4774), .ZN(n4772) );
  NAND2_X1 U5636 ( .A1(n8890), .A2(n8891), .ZN(n4774) );
  AND2_X1 U5637 ( .A1(n6619), .A2(n4783), .ZN(n4782) );
  INV_X1 U5638 ( .A(n6625), .ZN(n4783) );
  OR2_X1 U5639 ( .A1(n5278), .A2(n8903), .ZN(n5263) );
  AOI21_X1 U5640 ( .B1(n4762), .B2(n4765), .A(n4420), .ZN(n4760) );
  NAND2_X1 U5641 ( .A1(n6597), .A2(n4420), .ZN(n8966) );
  NAND2_X1 U5642 ( .A1(n4758), .A2(n4413), .ZN(n4752) );
  NAND2_X1 U5643 ( .A1(n4754), .A2(n8936), .ZN(n4753) );
  AND2_X1 U5644 ( .A1(n4413), .A2(n6639), .ZN(n4754) );
  AND2_X1 U5645 ( .A1(n6572), .A2(n6571), .ZN(n4523) );
  AOI21_X1 U5646 ( .B1(n5780), .B2(n5779), .A(n5778), .ZN(n5783) );
  NAND2_X1 U5647 ( .A1(n4396), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5381) );
  NAND2_X1 U5648 ( .A1(n6877), .A2(n6878), .ZN(n6876) );
  AND2_X1 U5649 ( .A1(n9917), .A2(n9916), .ZN(n9914) );
  NOR2_X1 U5650 ( .A1(n7218), .A2(n4462), .ZN(n9933) );
  AND2_X1 U5651 ( .A1(n5475), .A2(n5286), .ZN(n5368) );
  NOR2_X1 U5652 ( .A1(n9068), .A2(n4649), .ZN(n9072) );
  AND2_X1 U5653 ( .A1(n9069), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n4649) );
  NOR2_X1 U5654 ( .A1(n9072), .A2(n9071), .ZN(n9078) );
  AOI22_X1 U5655 ( .A1(n8113), .A2(n4881), .B1(n4890), .B2(n4884), .ZN(n4880)
         );
  NAND2_X1 U5656 ( .A1(n4882), .A2(n4884), .ZN(n4881) );
  OAI21_X1 U5657 ( .B1(n9139), .B2(n4593), .A(n4591), .ZN(n8088) );
  INV_X1 U5658 ( .A(n4594), .ZN(n4593) );
  AOI21_X1 U5659 ( .B1(n4594), .B2(n4595), .A(n4592), .ZN(n4591) );
  AND2_X1 U5660 ( .A1(n5180), .A2(n8115), .ZN(n9111) );
  OR2_X1 U5661 ( .A1(n9134), .A2(n9346), .ZN(n9118) );
  NOR2_X1 U5662 ( .A1(n9195), .A2(n4622), .ZN(n9169) );
  NAND2_X1 U5663 ( .A1(n9152), .A2(n4621), .ZN(n4620) );
  INV_X1 U5664 ( .A(n4622), .ZN(n4621) );
  NAND2_X1 U5665 ( .A1(n9184), .A2(n8082), .ZN(n9165) );
  NOR2_X1 U5666 ( .A1(n9195), .A2(n9366), .ZN(n9179) );
  NOR2_X1 U5667 ( .A1(n4626), .A2(n9378), .ZN(n4625) );
  OR2_X1 U5668 ( .A1(n9216), .A2(n9371), .ZN(n9195) );
  AOI21_X1 U5669 ( .B1(n9243), .B2(n4575), .A(n4453), .ZN(n4574) );
  INV_X1 U5670 ( .A(n9243), .ZN(n4576) );
  INV_X1 U5671 ( .A(n8072), .ZN(n4575) );
  AOI21_X1 U5672 ( .B1(n4403), .B2(n4920), .A(n4443), .ZN(n4919) );
  NOR2_X1 U5673 ( .A1(n9277), .A2(n4626), .ZN(n9227) );
  NOR2_X1 U5674 ( .A1(n9277), .A2(n4627), .ZN(n9247) );
  NAND2_X1 U5675 ( .A1(n5158), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n5336) );
  INV_X1 U5676 ( .A(n4896), .ZN(n4895) );
  AOI21_X1 U5677 ( .B1(n4896), .B2(n4900), .A(n4405), .ZN(n4894) );
  NAND2_X1 U5678 ( .A1(n4404), .A2(n9850), .ZN(n9317) );
  OR2_X1 U5679 ( .A1(n5513), .A2(n5373), .ZN(n5375) );
  NAND2_X1 U5680 ( .A1(n5157), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n5362) );
  INV_X1 U5681 ( .A(n5375), .ZN(n5157) );
  NAND2_X1 U5682 ( .A1(n9850), .A2(n4617), .ZN(n9823) );
  AND2_X1 U5683 ( .A1(n9850), .A2(n9865), .ZN(n9821) );
  OR2_X1 U5684 ( .A1(n5521), .A2(n7102), .ZN(n5539) );
  NAND2_X1 U5685 ( .A1(n5155), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n5541) );
  INV_X1 U5686 ( .A(n5539), .ZN(n5155) );
  AND2_X1 U5687 ( .A1(n5644), .A2(n5645), .ZN(n7643) );
  OAI21_X1 U5688 ( .B1(n4914), .B2(n4913), .A(n4450), .ZN(n4912) );
  NAND2_X1 U5689 ( .A1(n4916), .A2(n4914), .ZN(n9947) );
  NAND2_X1 U5690 ( .A1(n7496), .A2(n7495), .ZN(n4916) );
  NAND2_X1 U5691 ( .A1(n4590), .A2(n4432), .ZN(n7481) );
  NAND2_X1 U5692 ( .A1(n6902), .A2(n4613), .ZN(n4590) );
  NAND2_X1 U5693 ( .A1(n7473), .A2(n4587), .ZN(n7499) );
  INV_X1 U5694 ( .A(n7495), .ZN(n4587) );
  NAND2_X1 U5695 ( .A1(n5634), .A2(n7498), .ZN(n7495) );
  NAND2_X1 U5696 ( .A1(n5632), .A2(n5624), .ZN(n7609) );
  INV_X1 U5697 ( .A(n7609), .ZN(n7620) );
  NAND2_X1 U5698 ( .A1(n4614), .A2(n10019), .ZN(n7613) );
  NAND2_X1 U5699 ( .A1(n5960), .A2(n4613), .ZN(n5437) );
  NOR2_X1 U5700 ( .A1(n7564), .A2(n10009), .ZN(n7428) );
  OR2_X1 U5701 ( .A1(n5463), .A2(n6892), .ZN(n5402) );
  INV_X1 U5702 ( .A(n9018), .ZN(n7557) );
  NAND2_X1 U5703 ( .A1(n7376), .A2(n5575), .ZN(n4695) );
  NAND2_X1 U5704 ( .A1(n7362), .A2(n7363), .ZN(n7401) );
  NOR2_X1 U5705 ( .A1(n7361), .A2(n7408), .ZN(n7377) );
  NAND2_X1 U5706 ( .A1(n8040), .A2(n4613), .ZN(n5190) );
  NAND2_X1 U5707 ( .A1(n5323), .A2(n5322), .ZN(n9398) );
  NAND2_X1 U5708 ( .A1(n5334), .A2(n5333), .ZN(n9405) );
  AND2_X1 U5709 ( .A1(n6671), .A2(n6670), .ZN(n7112) );
  INV_X1 U5710 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n4710) );
  XNOR2_X1 U5711 ( .A(n5150), .B(n5149), .ZN(n8852) );
  XNOR2_X1 U5712 ( .A(n5197), .B(n5198), .ZN(n8055) );
  NAND2_X1 U5713 ( .A1(n4520), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5799) );
  NAND2_X1 U5714 ( .A1(n5069), .A2(n5068), .ZN(n5259) );
  NAND2_X1 U5715 ( .A1(n4544), .A2(n5033), .ZN(n5342) );
  NAND2_X1 U5716 ( .A1(n5029), .A2(n4549), .ZN(n4544) );
  NAND2_X1 U5717 ( .A1(n4834), .A2(n4835), .ZN(n5507) );
  NAND2_X1 U5718 ( .A1(n5009), .A2(n4557), .ZN(n4834) );
  NAND2_X1 U5719 ( .A1(n4840), .A2(n5014), .ZN(n5529) );
  NAND2_X1 U5720 ( .A1(n5518), .A2(n4962), .ZN(n4840) );
  OAI21_X1 U5721 ( .B1(n5501), .B2(n4848), .A(n4846), .ZN(n5474) );
  NAND2_X1 U5722 ( .A1(n5431), .A2(n5119), .ZN(n5482) );
  NAND2_X1 U5723 ( .A1(n4845), .A2(n4999), .ZN(n5481) );
  NAND2_X1 U5724 ( .A1(n5501), .A2(n4997), .ZN(n4845) );
  AND2_X1 U5725 ( .A1(n4528), .A2(n5460), .ZN(n5396) );
  NOR2_X1 U5726 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), .ZN(
        n5117) );
  INV_X1 U5727 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n5118) );
  INV_X1 U5728 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5419) );
  NAND2_X1 U5729 ( .A1(n4661), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5420) );
  INV_X1 U5730 ( .A(n5396), .ZN(n4661) );
  INV_X1 U5731 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4712) );
  NAND2_X1 U5732 ( .A1(n4802), .A2(n4806), .ZN(n8211) );
  AND4_X1 U5733 ( .A1(n6111), .A2(n6110), .A3(n6109), .A4(n6108), .ZN(n8179)
         );
  NAND2_X1 U5734 ( .A1(n7820), .A2(n6765), .ZN(n7831) );
  AND2_X1 U5735 ( .A1(n4803), .A2(n4811), .ZN(n4796) );
  OAI22_X1 U5736 ( .A1(n4799), .A2(n4798), .B1(n4801), .B2(n4811), .ZN(n4797)
         );
  NOR2_X1 U5737 ( .A1(n4803), .A2(n4811), .ZN(n4798) );
  INV_X1 U5738 ( .A(n4801), .ZN(n4799) );
  NAND2_X1 U5739 ( .A1(n4801), .A2(n8215), .ZN(n4800) );
  NAND2_X1 U5740 ( .A1(n4878), .A2(n6271), .ZN(n8763) );
  NAND2_X1 U5741 ( .A1(n4487), .A2(n8223), .ZN(n8226) );
  OAI21_X1 U5742 ( .B1(n8194), .B2(n4486), .A(n4447), .ZN(n4487) );
  OR2_X1 U5743 ( .A1(n4486), .A2(n8132), .ZN(n4485) );
  NAND2_X1 U5744 ( .A1(n6236), .A2(n6235), .ZN(n8779) );
  NAND2_X1 U5745 ( .A1(n4818), .A2(n7285), .ZN(n7316) );
  NAND2_X1 U5746 ( .A1(n7278), .A2(n4819), .ZN(n4818) );
  NAND2_X1 U5747 ( .A1(n4814), .A2(n6792), .ZN(n6817) );
  NAND2_X1 U5748 ( .A1(n5875), .A2(n5874), .ZN(n8783) );
  NAND2_X1 U5749 ( .A1(n7278), .A2(n6735), .ZN(n7292) );
  NAND2_X1 U5750 ( .A1(n8201), .A2(n4812), .ZN(n8274) );
  NAND2_X1 U5751 ( .A1(n8201), .A2(n8136), .ZN(n8273) );
  NAND2_X1 U5752 ( .A1(n8017), .A2(n8015), .ZN(n6776) );
  NAND2_X1 U5753 ( .A1(n8046), .A2(n8047), .ZN(n8172) );
  INV_X1 U5754 ( .A(n8321), .ZN(n8325) );
  NAND2_X1 U5755 ( .A1(n6827), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8317) );
  OAI21_X1 U5756 ( .B1(n8241), .B2(n8238), .A(n8237), .ZN(n8312) );
  NAND2_X1 U5757 ( .A1(n8040), .A2(n6245), .ZN(n6247) );
  NAND2_X1 U5758 ( .A1(n6820), .A2(n10096), .ZN(n8319) );
  NAND4_X1 U5759 ( .A1(n5959), .A2(n5958), .A3(n5957), .A4(n5956), .ZN(n8349)
         );
  OR2_X1 U5760 ( .A1(n5994), .A2(n5977), .ZN(n5980) );
  NAND4_X1 U5761 ( .A1(n5972), .A2(n5971), .A3(n5970), .A4(n5969), .ZN(n5990)
         );
  OR2_X1 U5762 ( .A1(n5994), .A2(n5967), .ZN(n5971) );
  OR2_X1 U5763 ( .A1(n6202), .A2(n7790), .ZN(n5970) );
  OR2_X1 U5764 ( .A1(n5992), .A2(n5968), .ZN(n5969) );
  OAI21_X1 U5765 ( .B1(n6005), .B2(n6952), .A(n9754), .ZN(n6977) );
  INV_X1 U5766 ( .A(n4572), .ZN(n6970) );
  AND2_X1 U5767 ( .A1(n4572), .A2(n4571), .ZN(n6983) );
  NAND2_X1 U5768 ( .A1(n6950), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n4571) );
  NAND2_X1 U5769 ( .A1(n8359), .A2(n6937), .ZN(n8373) );
  NAND2_X1 U5770 ( .A1(n8373), .A2(n8374), .ZN(n8372) );
  NOR2_X1 U5771 ( .A1(n7017), .A2(n4570), .ZN(n7020) );
  AND2_X1 U5772 ( .A1(n7022), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n4570) );
  INV_X1 U5773 ( .A(n4569), .ZN(n7135) );
  NAND2_X1 U5774 ( .A1(n7142), .A2(n7143), .ZN(n7146) );
  AOI21_X1 U5775 ( .B1(n7334), .B2(n7179), .A(n7333), .ZN(n8381) );
  NOR2_X1 U5776 ( .A1(n7448), .A2(n7447), .ZN(n7450) );
  AND2_X1 U5777 ( .A1(n6117), .A2(n6133), .ZN(n7845) );
  NOR2_X1 U5778 ( .A1(n8430), .A2(n4474), .ZN(n8445) );
  XNOR2_X1 U5779 ( .A(n4478), .B(n8672), .ZN(n8453) );
  NAND2_X1 U5780 ( .A1(n8444), .A2(n8443), .ZN(n4478) );
  AND2_X1 U5781 ( .A1(n6941), .A2(n8464), .ZN(n10056) );
  NAND2_X1 U5782 ( .A1(n6303), .A2(n6302), .ZN(n8753) );
  OAI21_X1 U5783 ( .B1(n8507), .B2(n10089), .A(n8506), .ZN(n8760) );
  INV_X1 U5784 ( .A(n8779), .ZN(n8580) );
  INV_X1 U5785 ( .A(n8610), .ZN(n4939) );
  NAND2_X1 U5786 ( .A1(n4518), .A2(n4725), .ZN(n8622) );
  NAND2_X1 U5787 ( .A1(n8650), .A2(n6383), .ZN(n8636) );
  OAI21_X1 U5788 ( .B1(n8676), .B2(n4931), .A(n4929), .ZN(n8643) );
  AND2_X1 U5789 ( .A1(n4933), .A2(n4424), .ZN(n8659) );
  NAND2_X1 U5790 ( .A1(n8676), .A2(n8482), .ZN(n4933) );
  NAND2_X1 U5791 ( .A1(n6188), .A2(n6187), .ZN(n8811) );
  NAND2_X1 U5792 ( .A1(n4517), .A2(n4719), .ZN(n8735) );
  NAND2_X1 U5793 ( .A1(n8028), .A2(n4946), .ZN(n8476) );
  NAND2_X1 U5794 ( .A1(n6104), .A2(n6103), .ZN(n8026) );
  NAND2_X1 U5795 ( .A1(n7700), .A2(n7699), .ZN(n7703) );
  INV_X1 U5796 ( .A(n4733), .ZN(n4732) );
  NAND2_X1 U5797 ( .A1(n5960), .A2(n6245), .ZN(n4734) );
  OAI21_X1 U5798 ( .B1(n5964), .B2(n9581), .A(n5963), .ZN(n4733) );
  INV_X1 U5799 ( .A(n10147), .ZN(n10103) );
  NAND2_X1 U5800 ( .A1(n7891), .A2(n7237), .ZN(n7749) );
  INV_X1 U5801 ( .A(n10102), .ZN(n8703) );
  OR2_X1 U5802 ( .A1(n7229), .A2(n10110), .ZN(n10096) );
  AND2_X1 U5803 ( .A1(n10081), .A2(n7688), .ZN(n10102) );
  INV_X1 U5804 ( .A(n10085), .ZN(n8727) );
  INV_X2 U5805 ( .A(n10200), .ZN(n10202) );
  AND2_X1 U5806 ( .A1(n5849), .A2(n5851), .ZN(n4949) );
  INV_X1 U5807 ( .A(n5829), .ZN(n5850) );
  INV_X1 U5808 ( .A(n6429), .ZN(n7662) );
  INV_X1 U5809 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n9695) );
  NOR2_X1 U5810 ( .A1(n6086), .A2(n4830), .ZN(n6149) );
  INV_X1 U5811 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n9644) );
  INV_X1 U5812 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6918) );
  INV_X1 U5813 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6912) );
  INV_X1 U5814 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6906) );
  OR2_X1 U5815 ( .A1(n5962), .A2(n5909), .ZN(n6959) );
  INV_X1 U5816 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6898) );
  INV_X1 U5817 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n4974) );
  NAND2_X1 U5818 ( .A1(n5177), .A2(n5176), .ZN(n9341) );
  NAND2_X1 U5819 ( .A1(n7723), .A2(n6536), .ZN(n7984) );
  AND2_X1 U5820 ( .A1(n6696), .A2(n7117), .ZN(n8979) );
  NAND2_X1 U5821 ( .A1(n5211), .A2(n5210), .ZN(n9363) );
  NAND2_X1 U5822 ( .A1(n4773), .A2(n4774), .ZN(n8944) );
  NAND2_X1 U5823 ( .A1(n6526), .A2(n7575), .ZN(n7722) );
  INV_X1 U5824 ( .A(n4629), .ZN(n4628) );
  OAI22_X1 U5825 ( .A1(n6893), .A2(n5463), .B1(n5464), .B2(n4973), .ZN(n4629)
         );
  OR2_X1 U5826 ( .A1(n6697), .A2(n7117), .ZN(n8972) );
  NAND2_X1 U5827 ( .A1(n4531), .A2(n4530), .ZN(n4529) );
  NOR2_X1 U5828 ( .A1(n4751), .A2(n8978), .ZN(n4530) );
  NAND2_X1 U5829 ( .A1(n8935), .A2(n4754), .ZN(n4531) );
  NAND2_X1 U5830 ( .A1(n4753), .A2(n4752), .ZN(n4751) );
  AND2_X1 U5831 ( .A1(n4759), .A2(n4756), .ZN(n4755) );
  NAND2_X1 U5832 ( .A1(n9249), .A2(n6693), .ZN(n8997) );
  AND2_X1 U5833 ( .A1(n7368), .A2(n5802), .ZN(n7042) );
  NAND2_X1 U5834 ( .A1(n5395), .A2(n5394), .ZN(n9017) );
  NOR2_X1 U5835 ( .A1(n5393), .A2(n4951), .ZN(n5395) );
  INV_X1 U5836 ( .A(n4664), .ZN(n7032) );
  INV_X1 U5837 ( .A(n4662), .ZN(n7091) );
  OAI22_X1 U5838 ( .A1(n4662), .A2(n7093), .B1(P1_REG2_REG_7__SCAN_IN), .B2(
        n7092), .ZN(n9909) );
  INV_X1 U5839 ( .A(n4658), .ZN(n7305) );
  INV_X1 U5840 ( .A(n4656), .ZN(n7599) );
  INV_X1 U5841 ( .A(n4653), .ZN(n9031) );
  OAI21_X1 U5842 ( .B1(n7919), .B2(n4651), .A(n4650), .ZN(n9048) );
  NAND2_X1 U5843 ( .A1(n4654), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n4651) );
  NAND2_X1 U5844 ( .A1(n9032), .A2(n4654), .ZN(n4650) );
  INV_X1 U5845 ( .A(n9034), .ZN(n4654) );
  INV_X1 U5846 ( .A(n9032), .ZN(n4652) );
  XNOR2_X1 U5847 ( .A(n4647), .B(n4646), .ZN(n9085) );
  INV_X1 U5848 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n4646) );
  OR2_X1 U5849 ( .A1(n9078), .A2(n4648), .ZN(n4647) );
  AND2_X1 U5850 ( .A1(n9080), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n4648) );
  INV_X1 U5851 ( .A(n9902), .ZN(n9938) );
  AOI21_X1 U5852 ( .B1(n8849), .B2(n4613), .A(n5144), .ZN(n9099) );
  NAND2_X1 U5853 ( .A1(n4889), .A2(n4891), .ZN(n9107) );
  AND2_X1 U5854 ( .A1(n9158), .A2(n9157), .ZN(n9359) );
  AOI21_X1 U5855 ( .B1(n8108), .B2(n4907), .A(n4400), .ZN(n9147) );
  NAND2_X1 U5856 ( .A1(n8108), .A2(n8107), .ZN(n9162) );
  NAND2_X1 U5857 ( .A1(n8080), .A2(n8079), .ZN(n9186) );
  NAND2_X1 U5858 ( .A1(n4700), .A2(n8073), .ZN(n9234) );
  NAND2_X1 U5859 ( .A1(n9242), .A2(n9243), .ZN(n4700) );
  OR2_X1 U5860 ( .A1(n9255), .A2(n4403), .ZN(n4918) );
  AND2_X1 U5861 ( .A1(n4924), .A2(n4923), .ZN(n9241) );
  NAND2_X1 U5862 ( .A1(n4701), .A2(n8067), .ZN(n9295) );
  NAND2_X1 U5863 ( .A1(n4898), .A2(n4902), .ZN(n9313) );
  NAND2_X1 U5864 ( .A1(n7957), .A2(n4899), .ZN(n4898) );
  AND2_X1 U5865 ( .A1(n9825), .A2(n7960), .ZN(n7962) );
  NAND2_X1 U5866 ( .A1(n7957), .A2(n7956), .ZN(n8095) );
  NAND2_X1 U5867 ( .A1(n4577), .A2(n4581), .ZN(n4967) );
  NAND2_X1 U5868 ( .A1(n7877), .A2(n7876), .ZN(n9842) );
  NOR2_X1 U5869 ( .A1(n9321), .A2(n7369), .ZN(n9953) );
  CLKBUF_X2 U5870 ( .A(n5574), .Z(n7522) );
  INV_X1 U5871 ( .A(n9972), .ZN(n9848) );
  NAND2_X1 U5872 ( .A1(n7204), .A2(n7203), .ZN(n10053) );
  NAND2_X1 U5873 ( .A1(n9338), .A2(n4428), .ZN(n9422) );
  AND2_X2 U5874 ( .A1(n7204), .A2(n7364), .ZN(n10042) );
  AND2_X1 U5875 ( .A1(n6834), .A2(n6686), .ZN(n9988) );
  INV_X1 U5876 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n4697) );
  NAND2_X1 U5877 ( .A1(n9438), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4698) );
  INV_X1 U5878 ( .A(n5165), .ZN(n9447) );
  NAND2_X1 U5879 ( .A1(n4960), .A2(n5074), .ZN(n5235) );
  NAND2_X1 U5880 ( .A1(n5617), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5619) );
  INV_X1 U5881 ( .A(n6433), .ZN(n7573) );
  XNOR2_X1 U5882 ( .A(n5292), .B(n5291), .ZN(n9086) );
  INV_X1 U5883 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n9593) );
  NAND2_X1 U5884 ( .A1(n5475), .A2(n4785), .ZN(n5343) );
  AND2_X1 U5885 ( .A1(n5475), .A2(n4786), .ZN(n5357) );
  INV_X1 U5886 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6920) );
  INV_X1 U5887 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n6916) );
  INV_X1 U5888 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n6908) );
  INV_X1 U5889 ( .A(n5960), .ZN(n6899) );
  INV_X1 U5890 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6889) );
  XNOR2_X1 U5891 ( .A(n5448), .B(n5449), .ZN(n6897) );
  NAND2_X1 U5892 ( .A1(n5418), .A2(n4660), .ZN(n6887) );
  OR2_X1 U5893 ( .A1(n5420), .A2(n5419), .ZN(n4660) );
  NAND2_X1 U5894 ( .A1(n6357), .A2(n4536), .ZN(n4537) );
  AOI211_X1 U5895 ( .C1(n9952), .C2(n9347), .A(n9131), .B(n9130), .ZN(n9132)
         );
  NAND2_X1 U5896 ( .A1(n4584), .A2(n4582), .ZN(P1_U3520) );
  OR2_X1 U5897 ( .A1(n10042), .A2(n4583), .ZN(n4582) );
  NAND2_X1 U5898 ( .A1(n9422), .A2(n10042), .ZN(n4584) );
  INV_X1 U5899 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n4583) );
  AND2_X1 U5900 ( .A1(n8591), .A2(n4940), .ZN(n4398) );
  AND2_X1 U5901 ( .A1(n4409), .A2(n6407), .ZN(n4399) );
  NAND2_X1 U5902 ( .A1(n8626), .A2(n4735), .ZN(n4737) );
  INV_X1 U5903 ( .A(n7615), .ZN(n10019) );
  INV_X2 U5904 ( .A(n5488), .ZN(n5523) );
  NAND2_X1 U5905 ( .A1(n4878), .A2(n4427), .ZN(n6324) );
  AND2_X1 U5906 ( .A1(n9175), .A2(n8110), .ZN(n4400) );
  INV_X1 U5907 ( .A(n8909), .ZN(n4758) );
  AOI21_X1 U5908 ( .B1(n5133), .B2(n4975), .A(n5132), .ZN(n9091) );
  INV_X1 U5909 ( .A(n8029), .ZN(n4948) );
  OR2_X1 U5910 ( .A1(n6394), .A2(n4724), .ZN(n4401) );
  AND2_X1 U5911 ( .A1(n4638), .A2(n9808), .ZN(n4402) );
  OR2_X1 U5912 ( .A1(n8103), .A2(n9258), .ZN(n4403) );
  INV_X1 U5913 ( .A(n7996), .ZN(n4945) );
  AND2_X1 U5914 ( .A1(n4617), .A2(n4616), .ZN(n4404) );
  AND2_X1 U5915 ( .A1(n9408), .A2(n9005), .ZN(n4405) );
  INV_X1 U5916 ( .A(n8073), .ZN(n4699) );
  NAND2_X1 U5917 ( .A1(n8926), .A2(n8928), .ZN(n8927) );
  INV_X1 U5918 ( .A(n7521), .ZN(n7408) );
  AND2_X1 U5919 ( .A1(n4890), .A2(n4887), .ZN(n4406) );
  NAND2_X1 U5920 ( .A1(n5511), .A2(n5510), .ZN(n7991) );
  INV_X1 U5921 ( .A(n4807), .ZN(n4806) );
  OAI22_X1 U5922 ( .A1(n8311), .A2(n4808), .B1(n8163), .B2(n8164), .ZN(n4807)
         );
  NOR2_X1 U5923 ( .A1(n4730), .A2(n4729), .ZN(n8649) );
  NAND2_X1 U5924 ( .A1(n6089), .A2(n6088), .ZN(n8023) );
  AND2_X1 U5925 ( .A1(n5635), .A2(n5634), .ZN(n4407) );
  AND2_X1 U5926 ( .A1(n5734), .A2(n4423), .ZN(n4408) );
  AND2_X1 U5927 ( .A1(n6403), .A2(n8668), .ZN(n4409) );
  AND2_X1 U5928 ( .A1(n4718), .A2(n6367), .ZN(n4410) );
  NAND2_X1 U5929 ( .A1(n5232), .A2(n5231), .ZN(n9166) );
  AND2_X1 U5930 ( .A1(n6541), .A2(n6536), .ZN(n4411) );
  AND3_X1 U5931 ( .A1(n6041), .A2(n6040), .A3(n6039), .ZN(n10157) );
  INV_X1 U5932 ( .A(n6724), .ZN(n6739) );
  INV_X1 U5933 ( .A(n5999), .ZN(n5964) );
  OR2_X1 U5934 ( .A1(n6410), .A2(n10123), .ZN(n6726) );
  NAND2_X1 U5935 ( .A1(n6342), .A2(n6372), .ZN(n4412) );
  BUF_X1 U5936 ( .A(n5994), .Z(n6307) );
  NAND2_X1 U5937 ( .A1(n5983), .A2(n5808), .ZN(n5950) );
  NAND4_X1 U5938 ( .A1(n5998), .A2(n5997), .A3(n5996), .A4(n5995), .ZN(n6725)
         );
  NAND2_X1 U5939 ( .A1(n6645), .A2(n6644), .ZN(n4413) );
  AND2_X1 U5940 ( .A1(n8551), .A2(n4634), .ZN(n4414) );
  NAND2_X1 U5941 ( .A1(n5786), .A2(n5127), .ZN(n4415) );
  AND2_X1 U5942 ( .A1(n6225), .A2(n6387), .ZN(n8609) );
  AND3_X1 U5943 ( .A1(n5416), .A2(n5415), .A3(n5414), .ZN(n4416) );
  INV_X1 U5944 ( .A(n6336), .ZN(n7684) );
  AND2_X1 U5945 ( .A1(n7876), .A2(n7878), .ZN(n4417) );
  NAND2_X1 U5946 ( .A1(n6744), .A2(n6743), .ZN(n4418) );
  AND2_X1 U5947 ( .A1(n8651), .A2(n6382), .ZN(n4419) );
  INV_X1 U5948 ( .A(n6458), .ZN(n6473) );
  AND2_X1 U5949 ( .A1(n6340), .A2(n6367), .ZN(n7704) );
  INV_X1 U5950 ( .A(n7237), .ZN(n4935) );
  NAND2_X1 U5951 ( .A1(n4918), .A2(n4920), .ZN(n9226) );
  NAND2_X1 U5952 ( .A1(n6293), .A2(n6292), .ZN(n8470) );
  INV_X1 U5953 ( .A(n8470), .ZN(n9792) );
  XOR2_X1 U5954 ( .A(n6593), .B(n6547), .Z(n4420) );
  AND2_X1 U5955 ( .A1(n4666), .A2(n8059), .ZN(n4421) );
  AND2_X1 U5956 ( .A1(n4785), .A2(n4784), .ZN(n4422) );
  XNOR2_X1 U5957 ( .A(n5872), .B(P2_IR_REG_21__SCAN_IN), .ZN(n6819) );
  INV_X1 U5958 ( .A(n8237), .ZN(n4810) );
  XNOR2_X1 U5959 ( .A(n4950), .B(n5852), .ZN(n5856) );
  AND3_X1 U5960 ( .A1(n5733), .A2(n4602), .A3(n8086), .ZN(n4423) );
  AND3_X1 U5961 ( .A1(n4791), .A2(n4794), .A3(n4790), .ZN(n5919) );
  INV_X1 U5962 ( .A(n6378), .ZN(n4515) );
  NAND2_X1 U5963 ( .A1(n6265), .A2(n6264), .ZN(n8768) );
  INV_X1 U5964 ( .A(n9140), .ZN(n4598) );
  XNOR2_X1 U5965 ( .A(n9351), .B(n9126), .ZN(n9140) );
  NAND2_X1 U5966 ( .A1(n8681), .A2(n8698), .ZN(n4424) );
  NAND2_X1 U5968 ( .A1(n5275), .A2(n5274), .ZN(n9381) );
  NAND2_X1 U5969 ( .A1(n5190), .A2(n5189), .ZN(n9351) );
  INV_X1 U5970 ( .A(n9351), .ZN(n4618) );
  NAND2_X1 U5971 ( .A1(n6162), .A2(n6161), .ZN(n8822) );
  AND2_X1 U5972 ( .A1(n4516), .A2(n6378), .ZN(n4425) );
  AND2_X1 U5973 ( .A1(n6771), .A2(n6770), .ZN(n4426) );
  NAND2_X1 U5974 ( .A1(n5372), .A2(n5371), .ZN(n7979) );
  NAND2_X1 U5975 ( .A1(n6393), .A2(n6279), .ZN(n8494) );
  INV_X1 U5976 ( .A(n8494), .ZN(n8539) );
  AND3_X1 U5977 ( .A1(n5987), .A2(n5988), .A3(n5989), .ZN(n7265) );
  INV_X1 U5978 ( .A(n7265), .ZN(n4942) );
  NOR2_X1 U5979 ( .A1(n8544), .A2(n4877), .ZN(n4427) );
  INV_X1 U5980 ( .A(n9139), .ZN(n4599) );
  AND2_X1 U5981 ( .A1(n9339), .A2(n9337), .ZN(n4428) );
  AND2_X1 U5982 ( .A1(n8565), .A2(n4687), .ZN(n4429) );
  AND2_X1 U5983 ( .A1(n8626), .A2(n6385), .ZN(n4430) );
  NAND2_X1 U5984 ( .A1(n5253), .A2(n5252), .ZN(n9378) );
  AND2_X1 U5985 ( .A1(n6531), .A2(n7575), .ZN(n4431) );
  AND2_X1 U5986 ( .A1(n6385), .A2(n6327), .ZN(n8489) );
  AND2_X1 U5987 ( .A1(n5504), .A2(n4588), .ZN(n4432) );
  AND2_X1 U5988 ( .A1(n7704), .A2(n7684), .ZN(n4433) );
  INV_X1 U5989 ( .A(n4900), .ZN(n4899) );
  OR2_X1 U5990 ( .A1(n8094), .A2(n4901), .ZN(n4900) );
  AND2_X1 U5991 ( .A1(n6381), .A2(n4519), .ZN(n4434) );
  NAND2_X1 U5992 ( .A1(n4737), .A2(n6387), .ZN(n4435) );
  AND2_X1 U5993 ( .A1(n4725), .A2(n8489), .ZN(n4436) );
  AND2_X1 U5994 ( .A1(n4421), .A2(n6323), .ZN(n4437) );
  AND2_X1 U5995 ( .A1(n8757), .A2(n8338), .ZN(n6394) );
  NOR2_X1 U5996 ( .A1(n9849), .A2(n7989), .ZN(n4438) );
  NOR2_X1 U5997 ( .A1(n8475), .A2(n8474), .ZN(n4439) );
  NOR2_X1 U5998 ( .A1(n8783), .A2(n8599), .ZN(n4440) );
  INV_X1 U5999 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n9439) );
  NOR2_X1 U6000 ( .A1(n6632), .A2(n8956), .ZN(n8881) );
  INV_X1 U6001 ( .A(n8881), .ZN(n4746) );
  AND2_X1 U6002 ( .A1(n4665), .A2(n4437), .ZN(n4441) );
  NOR2_X1 U6003 ( .A1(n6386), .A2(n4542), .ZN(n4442) );
  NAND2_X1 U6004 ( .A1(n5223), .A2(n5222), .ZN(n9356) );
  NOR2_X1 U6005 ( .A1(n9381), .A2(n9003), .ZN(n4443) );
  NOR2_X1 U6006 ( .A1(n8485), .A2(n8484), .ZN(n4444) );
  NAND2_X1 U6007 ( .A1(n5679), .A2(n5677), .ZN(n4445) );
  NAND2_X1 U6008 ( .A1(n9341), .A2(n9002), .ZN(n4446) );
  AND2_X1 U6009 ( .A1(n4485), .A2(n8142), .ZN(n4447) );
  NAND2_X1 U6010 ( .A1(n6346), .A2(n6157), .ZN(n4448) );
  INV_X1 U6011 ( .A(n4947), .ZN(n4946) );
  NAND2_X1 U6012 ( .A1(n4948), .A2(n8027), .ZN(n4947) );
  INV_X1 U6013 ( .A(n4941), .ZN(n8794) );
  NAND2_X1 U6014 ( .A1(n4939), .A2(n6386), .ZN(n4941) );
  AND2_X1 U6015 ( .A1(n5016), .A2(SI_11_), .ZN(n4449) );
  INV_X1 U6016 ( .A(n4833), .ZN(n4832) );
  NAND2_X1 U6017 ( .A1(n4835), .A2(n4841), .ZN(n4833) );
  OR2_X1 U6018 ( .A1(n9011), .A2(n7647), .ZN(n4450) );
  NAND2_X1 U6019 ( .A1(n5798), .A2(n5794), .ZN(n4451) );
  AND2_X1 U6020 ( .A1(n9152), .A2(n5233), .ZN(n4452) );
  NAND2_X1 U6021 ( .A1(n5726), .A2(n5733), .ZN(n8113) );
  INV_X1 U6022 ( .A(n8113), .ZN(n4890) );
  OR2_X1 U6023 ( .A1(n4699), .A2(n8074), .ZN(n4453) );
  INV_X1 U6024 ( .A(n4932), .ZN(n4931) );
  AND2_X1 U6025 ( .A1(n8483), .A2(n4424), .ZN(n4932) );
  INV_X1 U6026 ( .A(n9108), .ZN(n9104) );
  AND2_X1 U6027 ( .A1(n5732), .A2(n8086), .ZN(n9108) );
  AND2_X1 U6028 ( .A1(n4893), .A2(n9296), .ZN(n4454) );
  AND2_X1 U6029 ( .A1(n4819), .A2(n4418), .ZN(n4455) );
  AND2_X1 U6030 ( .A1(n7635), .A2(n7495), .ZN(n4456) );
  AND2_X1 U6031 ( .A1(n8068), .A2(n8067), .ZN(n4457) );
  AND2_X1 U6032 ( .A1(n7701), .A2(n7699), .ZN(n4458) );
  AND2_X1 U6033 ( .A1(n4889), .A2(n4887), .ZN(n4459) );
  NAND2_X1 U6034 ( .A1(n6198), .A2(n6197), .ZN(n8805) );
  INV_X1 U6035 ( .A(n4750), .ZN(n4749) );
  NOR2_X1 U6036 ( .A1(n4758), .A2(n8936), .ZN(n4750) );
  AND2_X1 U6037 ( .A1(n6388), .A2(n6387), .ZN(n4460) );
  NAND2_X1 U6038 ( .A1(n6436), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n4461) );
  INV_X1 U6039 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5811) );
  INV_X1 U6040 ( .A(n7399), .ZN(n4602) );
  AND3_X1 U6041 ( .A1(n6008), .A2(n6007), .A3(n6006), .ZN(n10136) );
  XNOR2_X1 U6042 ( .A(n5116), .B(n5115), .ZN(n8845) );
  AND4_X1 U6043 ( .A1(n4527), .A2(n4526), .A3(n4525), .A4(n4696), .ZN(n5431)
         );
  AND2_X1 U6044 ( .A1(n7219), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n4462) );
  INV_X1 U6045 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n4694) );
  OAI21_X1 U6046 ( .B1(n6086), .B2(n4826), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n6172) );
  OAI21_X1 U6047 ( .B1(n7957), .B2(n4895), .A(n4894), .ZN(n9292) );
  NAND2_X1 U6048 ( .A1(n5239), .A2(n5238), .ZN(n9366) );
  INV_X1 U6049 ( .A(n9366), .ZN(n4623) );
  OR2_X1 U6050 ( .A1(n9277), .A2(n9269), .ZN(n4463) );
  NAND2_X1 U6051 ( .A1(n4761), .A2(n4760), .ZN(n8964) );
  NAND2_X1 U6052 ( .A1(n8919), .A2(n8915), .ZN(n8926) );
  NAND2_X1 U6053 ( .A1(n8662), .A2(n4419), .ZN(n8650) );
  INV_X1 U6054 ( .A(n8215), .ZN(n4811) );
  INV_X1 U6055 ( .A(n5452), .ZN(n5167) );
  AND2_X1 U6056 ( .A1(n5834), .A2(n5833), .ZN(n8757) );
  INV_X1 U6057 ( .A(n8757), .ZN(n4635) );
  OR2_X1 U6058 ( .A1(n8475), .A2(n8738), .ZN(n4464) );
  AND2_X1 U6059 ( .A1(n8028), .A2(n8027), .ZN(n4465) );
  NAND2_X1 U6060 ( .A1(n4773), .A2(n4771), .ZN(n8942) );
  INV_X1 U6061 ( .A(n8303), .ZN(n10151) );
  NAND2_X1 U6062 ( .A1(n4734), .A2(n4732), .ZN(n8303) );
  AND2_X1 U6063 ( .A1(n7998), .A2(n4722), .ZN(n4466) );
  NAND2_X1 U6064 ( .A1(n8699), .A2(n4640), .ZN(n4643) );
  AND2_X1 U6065 ( .A1(n4653), .A2(n4652), .ZN(n4467) );
  INV_X1 U6066 ( .A(n4619), .ZN(n9148) );
  NOR2_X1 U6067 ( .A1(n9195), .A2(n4620), .ZN(n4619) );
  AND2_X1 U6068 ( .A1(n8208), .A2(n8209), .ZN(n4468) );
  AND2_X1 U6069 ( .A1(n8371), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n4469) );
  NAND2_X1 U6070 ( .A1(n4422), .A2(n5475), .ZN(n4470) );
  OR2_X1 U6071 ( .A1(n6086), .A2(n4828), .ZN(n4471) );
  INV_X1 U6072 ( .A(n10165), .ZN(n7698) );
  AND2_X1 U6073 ( .A1(n5913), .A2(n5912), .ZN(n10165) );
  NAND2_X1 U6074 ( .A1(n7683), .A2(n4433), .ZN(n4717) );
  INV_X1 U6075 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n4784) );
  INV_X1 U6076 ( .A(n7736), .ZN(n4504) );
  NAND2_X1 U6077 ( .A1(n7683), .A2(n7684), .ZN(n7682) );
  NAND2_X1 U6078 ( .A1(n6119), .A2(n6118), .ZN(n8475) );
  INV_X1 U6079 ( .A(n8475), .ZN(n4637) );
  INV_X1 U6080 ( .A(n8915), .ZN(n4764) );
  NAND2_X1 U6081 ( .A1(n4916), .A2(n7497), .ZN(n7632) );
  INV_X1 U6082 ( .A(n8999), .ZN(n8976) );
  OR2_X1 U6083 ( .A1(n6698), .A2(n6695), .ZN(n8999) );
  NAND2_X1 U6084 ( .A1(n5347), .A2(n5346), .ZN(n9408) );
  INV_X1 U6085 ( .A(n9408), .ZN(n4615) );
  AND2_X1 U6086 ( .A1(n4717), .A2(n4410), .ZN(n4472) );
  NAND2_X1 U6087 ( .A1(n5360), .A2(n5359), .ZN(n9416) );
  INV_X1 U6088 ( .A(n9416), .ZN(n4616) );
  NAND2_X1 U6089 ( .A1(n4779), .A2(n4780), .ZN(n7584) );
  OR2_X1 U6090 ( .A1(n7845), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n4473) );
  INV_X1 U6091 ( .A(n8350), .ZN(n4692) );
  XNOR2_X1 U6092 ( .A(n5131), .B(n5130), .ZN(n5804) );
  INV_X1 U6093 ( .A(n6407), .ZN(n4496) );
  AND2_X1 U6094 ( .A1(n8432), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n4474) );
  AND2_X1 U6095 ( .A1(n6456), .A2(n6457), .ZN(n4475) );
  NAND2_X1 U6096 ( .A1(n7538), .A2(n7428), .ZN(n7611) );
  INV_X1 U6097 ( .A(n7611), .ZN(n4614) );
  NAND2_X1 U6098 ( .A1(n6921), .A2(n6819), .ZN(n4476) );
  INV_X1 U6099 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n6320) );
  INV_X1 U6100 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n4792) );
  INV_X1 U6101 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5869) );
  XNOR2_X1 U6102 ( .A(n5748), .B(n5749), .ZN(n7494) );
  XNOR2_X1 U6103 ( .A(n4698), .B(n4697), .ZN(n9442) );
  INV_X1 U6104 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n4528) );
  INV_X1 U6105 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n8441) );
  INV_X1 U6106 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n4715) );
  NAND2_X1 U6107 ( .A1(n8693), .A2(n8695), .ZN(n8692) );
  OAI22_X2 U6108 ( .A1(n8613), .A2(n8489), .B1(n8600), .B2(n8795), .ZN(n8610)
         );
  NAND2_X1 U6109 ( .A1(n7930), .A2(n7855), .ZN(n7995) );
  AOI21_X1 U6110 ( .B1(n8733), .B2(n8734), .A(n8478), .ZN(n8714) );
  AOI21_X1 U6111 ( .B1(n8517), .B2(n8522), .A(n8498), .ZN(n8500) );
  INV_X2 U6112 ( .A(n5832), .ZN(n6245) );
  NAND2_X2 U6113 ( .A1(n6360), .A2(n6020), .ZN(n7750) );
  OAI211_X1 U6114 ( .C1(n7893), .C2(n4935), .A(n4477), .B(n7750), .ZN(n4936)
         );
  OAI21_X2 U6115 ( .B1(n8685), .B2(n8822), .A(n8692), .ZN(n8676) );
  NAND2_X1 U6116 ( .A1(n4976), .A2(n5422), .ZN(n4979) );
  NAND2_X1 U6117 ( .A1(n7808), .A2(n7809), .ZN(n7853) );
  NAND2_X1 U6118 ( .A1(n7928), .A2(n7927), .ZN(n7930) );
  BUF_X1 U6119 ( .A(n5855), .Z(n8853) );
  AOI22_X2 U6120 ( .A1(n7766), .A2(n4942), .B1(n7768), .B2(n6718), .ZN(n7893)
         );
  INV_X1 U6121 ( .A(n6985), .ZN(n6956) );
  NAND2_X1 U6122 ( .A1(n6987), .A2(n6986), .ZN(n6985) );
  NAND2_X1 U6123 ( .A1(n7027), .A2(n7026), .ZN(n7142) );
  OAI21_X1 U6124 ( .B1(n8935), .B2(n8936), .A(n6639), .ZN(n8908) );
  OAI21_X1 U6125 ( .B1(n8919), .B2(n4765), .A(n4762), .ZN(n6596) );
  INV_X1 U6126 ( .A(n8916), .ZN(n4522) );
  AND2_X2 U6127 ( .A1(n8882), .A2(n8883), .ZN(n4532) );
  INV_X4 U6128 ( .A(n6665), .ZN(n6658) );
  OR2_X2 U6129 ( .A1(n7256), .A2(n7255), .ZN(n7276) );
  INV_X1 U6130 ( .A(n10123), .ZN(n7247) );
  NAND2_X1 U6131 ( .A1(n6717), .A2(n4490), .ZN(n4489) );
  NAND2_X1 U6132 ( .A1(n8187), .A2(n8155), .ZN(n4491) );
  NAND3_X1 U6133 ( .A1(n5820), .A2(n5922), .A3(n5811), .ZN(n5871) );
  NAND4_X1 U6134 ( .A1(n4493), .A2(n4495), .A3(n4492), .A4(n4494), .ZN(n4535)
         );
  NAND2_X1 U6135 ( .A1(n6405), .A2(n4399), .ZN(n4492) );
  OR4_X1 U6136 ( .A1(n6405), .A2(n6404), .A3(n4496), .A4(n8668), .ZN(n4493) );
  OAI21_X1 U6137 ( .B1(n8521), .B2(n4401), .A(n4510), .ZN(n6399) );
  INV_X1 U6138 ( .A(n8521), .ZN(n4509) );
  NAND2_X1 U6139 ( .A1(n7999), .A2(n4721), .ZN(n4517) );
  NAND2_X1 U6140 ( .A1(n5799), .A2(n5798), .ZN(n5801) );
  NAND2_X1 U6141 ( .A1(n5786), .A2(n4911), .ZN(n4520) );
  NAND3_X1 U6142 ( .A1(n7166), .A2(n4770), .A3(n4768), .ZN(n7164) );
  XNOR2_X1 U6143 ( .A(n6462), .B(n6464), .ZN(n7166) );
  NAND2_X2 U6144 ( .A1(n4522), .A2(n4521), .ZN(n8919) );
  NAND2_X1 U6145 ( .A1(n4524), .A2(n8987), .ZN(n8916) );
  OAI21_X1 U6146 ( .B1(n8870), .B2(n6573), .A(n4523), .ZN(n8987) );
  NAND2_X1 U6147 ( .A1(n8986), .A2(n8989), .ZN(n4524) );
  NAND2_X1 U6148 ( .A1(n7723), .A2(n4411), .ZN(n7982) );
  NAND3_X1 U6149 ( .A1(n8977), .A2(n8976), .A3(n4529), .ZN(n8984) );
  NOR2_X2 U6150 ( .A1(n4532), .A2(n8881), .ZN(n8935) );
  AND3_X1 U6151 ( .A1(n5287), .A2(n5288), .A3(n5286), .ZN(n4786) );
  NAND2_X2 U6152 ( .A1(n7416), .A2(n6435), .ZN(n6665) );
  NAND4_X1 U6153 ( .A1(n4534), .A2(n4537), .A3(n4533), .A4(n6432), .ZN(
        P2_U3244) );
  NAND2_X1 U6154 ( .A1(n4441), .A2(n7718), .ZN(n4533) );
  NAND2_X1 U6155 ( .A1(n4535), .A2(n7718), .ZN(n4534) );
  INV_X1 U6156 ( .A(n6356), .ZN(n4538) );
  OAI21_X1 U6157 ( .B1(n5029), .B2(n4547), .A(n4545), .ZN(n5331) );
  NAND2_X1 U6158 ( .A1(n5029), .A2(n5028), .ZN(n5356) );
  AOI21_X1 U6159 ( .B1(n8359), .B2(n4563), .A(n4561), .ZN(n6991) );
  OAI21_X1 U6160 ( .B1(n8359), .B2(n4565), .A(n4563), .ZN(n4567) );
  INV_X1 U6161 ( .A(n4567), .ZN(n6993) );
  INV_X1 U6162 ( .A(n6992), .ZN(n4566) );
  OAI21_X2 U6163 ( .B1(n9263), .B2(n4576), .A(n4574), .ZN(n9209) );
  NAND2_X1 U6164 ( .A1(n4703), .A2(n7499), .ZN(n9955) );
  OAI21_X1 U6165 ( .B1(n4605), .B2(n4445), .A(n5678), .ZN(n5684) );
  NOR2_X1 U6166 ( .A1(n4607), .A2(n9309), .ZN(n4606) );
  AOI21_X1 U6167 ( .B1(n4612), .B2(n4611), .A(n4610), .ZN(n4609) );
  NAND3_X1 U6168 ( .A1(n4404), .A2(n4615), .A3(n9850), .ZN(n9319) );
  INV_X1 U6169 ( .A(n9277), .ZN(n4624) );
  NAND2_X1 U6170 ( .A1(n4625), .A2(n4624), .ZN(n9216) );
  INV_X1 U6171 ( .A(n4643), .ZN(n8667) );
  XNOR2_X1 U6172 ( .A(n9030), .B(n9036), .ZN(n7919) );
  MUX2_X1 U6173 ( .A(n6841), .B(P1_REG2_REG_2__SCAN_IN), .S(n6887), .Z(n6878)
         );
  NAND2_X1 U6174 ( .A1(n6313), .A2(n4667), .ZN(n4665) );
  NAND2_X1 U6175 ( .A1(n4665), .A2(n4421), .ZN(n6357) );
  INV_X1 U6176 ( .A(n6321), .ZN(n4667) );
  NAND2_X1 U6177 ( .A1(n6158), .A2(n4673), .ZN(n4677) );
  INV_X1 U6178 ( .A(n4672), .ZN(n4676) );
  NAND3_X1 U6179 ( .A1(n4681), .A2(n4678), .A3(n4945), .ZN(n6131) );
  NAND2_X1 U6180 ( .A1(n4692), .A2(n7785), .ZN(n6364) );
  OAI211_X2 U6181 ( .C1(n6897), .C2(n5832), .A(n5925), .B(n5924), .ZN(n7785)
         );
  NAND2_X1 U6182 ( .A1(n4695), .A2(n5576), .ZN(n5577) );
  OAI21_X1 U6183 ( .B1(n4695), .B2(n5758), .A(n5757), .ZN(n5762) );
  XNOR2_X1 U6184 ( .A(n4695), .B(n7511), .ZN(n7518) );
  NAND2_X1 U6185 ( .A1(n4701), .A2(n4457), .ZN(n9293) );
  NAND2_X1 U6186 ( .A1(n8080), .A2(n4702), .ZN(n9184) );
  NAND2_X1 U6187 ( .A1(n9955), .A2(n7875), .ZN(n7877) );
  NAND2_X1 U6188 ( .A1(n7499), .A2(n7498), .ZN(n7638) );
  INV_X1 U6189 ( .A(n7498), .ZN(n4704) );
  NAND2_X1 U6190 ( .A1(n9825), .A2(n4705), .ZN(n8065) );
  INV_X1 U6191 ( .A(n9106), .ZN(n4707) );
  XNOR2_X1 U6192 ( .A(n4709), .B(n9108), .ZN(n4708) );
  NOR2_X1 U6193 ( .A1(n9123), .A2(n9103), .ZN(n4709) );
  NAND3_X1 U6194 ( .A1(n5285), .A2(n4952), .A3(n4909), .ZN(n5134) );
  NAND4_X1 U6195 ( .A1(n5285), .A2(n4909), .A3(n4710), .A4(n4952), .ZN(n5137)
         );
  XNOR2_X1 U6196 ( .A(n6440), .B(n9991), .ZN(n7363) );
  NAND2_X2 U6197 ( .A1(n4713), .A2(n4711), .ZN(n4975) );
  NAND3_X1 U6198 ( .A1(n4712), .A2(P1_ADDR_REG_19__SCAN_IN), .A3(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n4711) );
  NAND3_X1 U6199 ( .A1(n8441), .A2(n4715), .A3(n4714), .ZN(n4713) );
  MUX2_X1 U6200 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(P1_DATAO_REG_1__SCAN_IN), 
        .S(n5831), .Z(n5461) );
  NAND2_X1 U6201 ( .A1(n4737), .A2(n4460), .ZN(n8594) );
  AND2_X1 U6202 ( .A1(n4738), .A2(n4461), .ZN(n4740) );
  NAND3_X1 U6203 ( .A1(n7373), .A2(n6834), .A3(n7361), .ZN(n4738) );
  NAND3_X1 U6204 ( .A1(n6435), .A2(n7416), .A3(n7361), .ZN(n4741) );
  NAND2_X1 U6205 ( .A1(n6867), .A2(n6866), .ZN(n6865) );
  NAND2_X1 U6206 ( .A1(n4740), .A2(n4739), .ZN(n6866) );
  AND2_X1 U6207 ( .A1(n4742), .A2(n4741), .ZN(n6867) );
  AND2_X1 U6208 ( .A1(n6436), .A2(P1_IR_REG_0__SCAN_IN), .ZN(n4743) );
  NAND3_X1 U6209 ( .A1(n4745), .A2(n4755), .A3(n4744), .ZN(n8977) );
  NAND2_X1 U6210 ( .A1(n8881), .A2(n4750), .ZN(n4744) );
  NAND2_X1 U6211 ( .A1(n8882), .A2(n4747), .ZN(n4745) );
  NAND2_X1 U6212 ( .A1(n8919), .A2(n4762), .ZN(n4761) );
  AND2_X2 U6213 ( .A1(n5431), .A2(n4766), .ZN(n5285) );
  NAND2_X1 U6214 ( .A1(n6448), .A2(n7127), .ZN(n7151) );
  NAND2_X1 U6215 ( .A1(n4769), .A2(n6457), .ZN(n4768) );
  NAND3_X1 U6216 ( .A1(n6457), .A2(n6448), .A3(n7127), .ZN(n4770) );
  NAND2_X1 U6217 ( .A1(n7150), .A2(n6457), .ZN(n7165) );
  NAND2_X1 U6218 ( .A1(n7151), .A2(n4475), .ZN(n7150) );
  NAND2_X1 U6219 ( .A1(n7391), .A2(n4781), .ZN(n4779) );
  NAND2_X1 U6220 ( .A1(n8899), .A2(n6619), .ZN(n6624) );
  NAND4_X1 U6221 ( .A1(n4794), .A2(n5809), .A3(n5808), .A4(n4793), .ZN(n5937)
         );
  NAND2_X1 U6222 ( .A1(n8241), .A2(n4796), .ZN(n4795) );
  OAI211_X1 U6223 ( .C1(n8241), .C2(n4800), .A(n4797), .B(n4795), .ZN(n8222)
         );
  NAND2_X1 U6224 ( .A1(n8241), .A2(n4809), .ZN(n4802) );
  NAND2_X1 U6225 ( .A1(n4814), .A2(n4813), .ZN(n8290) );
  NAND2_X1 U6226 ( .A1(n4455), .A2(n7278), .ZN(n4815) );
  OAI21_X1 U6227 ( .B1(n7831), .B2(n7830), .A(n6768), .ZN(n7944) );
  NAND2_X1 U6228 ( .A1(n4842), .A2(n4843), .ZN(n5009) );
  NAND2_X1 U6229 ( .A1(n5501), .A2(n4846), .ZN(n4842) );
  NAND2_X1 U6230 ( .A1(n5304), .A2(n5051), .ZN(n4853) );
  OAI21_X1 U6231 ( .B1(n5304), .B2(n4856), .A(n4854), .ZN(n5273) );
  NAND2_X1 U6232 ( .A1(n4852), .A2(n4850), .ZN(n5064) );
  NAND2_X1 U6233 ( .A1(n5304), .A2(n4854), .ZN(n4852) );
  NAND2_X1 U6234 ( .A1(n5208), .A2(n4863), .ZN(n4861) );
  NAND2_X1 U6235 ( .A1(n5208), .A2(n4870), .ZN(n4862) );
  OR2_X1 U6236 ( .A1(n5208), .A2(n5084), .ZN(n4867) );
  NAND2_X1 U6237 ( .A1(n6393), .A2(n6324), .ZN(n6281) );
  NAND2_X1 U6238 ( .A1(n5831), .A2(n4970), .ZN(n5975) );
  OAI21_X1 U6239 ( .B1(n9117), .B2(n4883), .A(n4879), .ZN(n9334) );
  INV_X1 U6240 ( .A(n4887), .ZN(n4882) );
  OR2_X1 U6241 ( .A1(n9346), .A2(n9142), .ZN(n4891) );
  NAND2_X1 U6242 ( .A1(n7957), .A2(n4894), .ZN(n4892) );
  NAND2_X1 U6243 ( .A1(n4892), .A2(n4454), .ZN(n8098) );
  OR2_X1 U6244 ( .A1(n9416), .A2(n9006), .ZN(n4902) );
  NAND4_X1 U6245 ( .A1(n5117), .A2(n5396), .A3(n5419), .A4(n5118), .ZN(n5429)
         );
  NAND3_X1 U6246 ( .A1(n5396), .A2(n5117), .A3(n5419), .ZN(n5446) );
  NAND2_X1 U6247 ( .A1(n8108), .A2(n4905), .ZN(n4904) );
  AOI21_X1 U6248 ( .B1(n7496), .B2(n4456), .A(n4912), .ZN(n7637) );
  NAND2_X1 U6249 ( .A1(n9255), .A2(n4920), .ZN(n4917) );
  NAND2_X1 U6250 ( .A1(n4917), .A2(n4919), .ZN(n8104) );
  INV_X1 U6251 ( .A(n4924), .ZN(n9257) );
  NAND2_X1 U6252 ( .A1(n4936), .A2(n7238), .ZN(n10100) );
  NAND2_X1 U6253 ( .A1(n8610), .A2(n4398), .ZN(n4937) );
  NOR2_X1 U6254 ( .A1(n8794), .A2(n8491), .ZN(n8585) );
  OAI21_X2 U6255 ( .B1(n7997), .B2(n4947), .A(n4944), .ZN(n8733) );
  NAND2_X1 U6256 ( .A1(n7700), .A2(n4458), .ZN(n7807) );
  NAND2_X2 U6257 ( .A1(n7671), .A2(n6336), .ZN(n7700) );
  AND2_X1 U6258 ( .A1(n5921), .A2(n5811), .ZN(n5909) );
  NAND2_X1 U6259 ( .A1(n5850), .A2(n4949), .ZN(n8846) );
  OAI22_X2 U6260 ( .A1(n7733), .A2(n7668), .B1(n8303), .B2(n8349), .ZN(n10078)
         );
  OAI21_X2 U6261 ( .B1(n7665), .B2(n7664), .A(n7667), .ZN(n7733) );
  NAND2_X1 U6262 ( .A1(n5865), .A2(n5864), .ZN(n6086) );
  INV_X1 U6263 ( .A(n6050), .ZN(n5865) );
  AND2_X1 U6264 ( .A1(n6359), .A2(n6358), .ZN(n7894) );
  NAND2_X1 U6265 ( .A1(n7894), .A2(n7895), .ZN(n7754) );
  NAND2_X1 U6266 ( .A1(n6716), .A2(n6819), .ZN(n7680) );
  NAND2_X1 U6267 ( .A1(n6716), .A2(n8668), .ZN(n6410) );
  NAND2_X1 U6268 ( .A1(n5561), .A2(n5560), .ZN(n5617) );
  NAND2_X1 U6269 ( .A1(n5559), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5561) );
  NAND2_X1 U6270 ( .A1(n8864), .A2(n6660), .ZN(n6714) );
  XNOR2_X1 U6271 ( .A(n8088), .B(n4890), .ZN(n8093) );
  AND2_X1 U6272 ( .A1(n5909), .A2(n5862), .ZN(n5899) );
  NAND2_X1 U6273 ( .A1(n4397), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5415) );
  XNOR2_X1 U6274 ( .A(n8864), .B(n8863), .ZN(n8869) );
  NAND2_X1 U6275 ( .A1(n8977), .A2(n6654), .ZN(n8864) );
  NAND2_X1 U6276 ( .A1(n5542), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n5457) );
  AND2_X2 U6277 ( .A1(n5856), .A2(n8853), .ZN(n5991) );
  NAND2_X1 U6278 ( .A1(n5856), .A2(n5857), .ZN(n5994) );
  OR2_X1 U6279 ( .A1(n8716), .A2(n8715), .ZN(n8829) );
  OAI21_X1 U6280 ( .B1(n7322), .B2(n7324), .A(n7323), .ZN(n6500) );
  OR2_X1 U6281 ( .A1(n6928), .A2(n6005), .ZN(n6006) );
  OR2_X1 U6282 ( .A1(n4390), .A2(n6954), .ZN(n5989) );
  MUX2_X1 U6283 ( .A(P2_IR_REG_0__SCAN_IN), .B(n8860), .S(n6928), .Z(n7792) );
  OR2_X1 U6284 ( .A1(n5992), .A2(n6953), .ZN(n5978) );
  INV_X1 U6285 ( .A(n5856), .ZN(n8850) );
  AND2_X1 U6286 ( .A1(n5542), .A2(n5392), .ZN(n4951) );
  AND2_X1 U6287 ( .A1(n5186), .A2(n5185), .ZN(n9127) );
  AND2_X1 U6288 ( .A1(n8539), .A2(n8540), .ZN(n4953) );
  OR2_X1 U6289 ( .A1(n9232), .A2(n9246), .ZN(n4955) );
  AOI21_X1 U6290 ( .B1(n7754), .B2(n7751), .A(n7750), .ZN(n7755) );
  AND4_X1 U6291 ( .A1(n8516), .A2(n8493), .A3(n8539), .A4(n6350), .ZN(n4956)
         );
  AND3_X1 U6292 ( .A1(n8250), .A2(n8324), .A3(n8251), .ZN(n4957) );
  AND2_X1 U6293 ( .A1(n9199), .A2(n9215), .ZN(n4958) );
  AND3_X1 U6294 ( .A1(n5305), .A2(n5307), .A3(n5290), .ZN(n4959) );
  OR2_X1 U6295 ( .A1(n7118), .A2(n4393), .ZN(n9959) );
  OR2_X1 U6296 ( .A1(n4975), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n4961) );
  AND2_X1 U6297 ( .A1(n5014), .A2(n5013), .ZN(n4962) );
  AND2_X1 U6298 ( .A1(n5028), .A2(n5027), .ZN(n4963) );
  INV_X1 U6299 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n4980) );
  AND2_X1 U6300 ( .A1(n5008), .A2(n5007), .ZN(n4964) );
  NAND2_X1 U6301 ( .A1(n9099), .A2(n9001), .ZN(n4965) );
  INV_X1 U6302 ( .A(n9970), .ZN(n9836) );
  AND2_X1 U6303 ( .A1(n9015), .A2(n7462), .ZN(n4966) );
  NAND2_X1 U6304 ( .A1(n6608), .A2(n6609), .ZN(n4968) );
  OAI21_X2 U6305 ( .B1(n7973), .B2(n6554), .A(n6553), .ZN(n8870) );
  AND2_X1 U6306 ( .A1(n6081), .A2(n6288), .ZN(n6082) );
  AOI21_X1 U6307 ( .B1(n6083), .B2(n6315), .A(n6082), .ZN(n6084) );
  NAND2_X1 U6308 ( .A1(n4956), .A2(n8499), .ZN(n6351) );
  NAND2_X1 U6309 ( .A1(n9091), .A2(n5722), .ZN(n5720) );
  INV_X1 U6310 ( .A(n6400), .ZN(n6401) );
  NAND2_X1 U6311 ( .A1(n6401), .A2(n6353), .ZN(n6354) );
  INV_X1 U6312 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n5119) );
  NAND2_X1 U6313 ( .A1(n6450), .A2(n6449), .ZN(n6451) );
  INV_X1 U6314 ( .A(n9187), .ZN(n8081) );
  INV_X1 U6315 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n5127) );
  INV_X1 U6316 ( .A(n6200), .ZN(n5844) );
  AND2_X1 U6317 ( .A1(n6717), .A2(n10123), .ZN(n6323) );
  INV_X1 U6318 ( .A(n6212), .ZN(n5845) );
  NAND2_X1 U6319 ( .A1(n8567), .A2(n8565), .ZN(n8556) );
  NAND2_X1 U6320 ( .A1(n6322), .A2(n6429), .ZN(n6717) );
  INV_X1 U6321 ( .A(n6629), .ZN(n6630) );
  XNOR2_X1 U6322 ( .A(n6451), .B(n6547), .ZN(n6452) );
  INV_X1 U6323 ( .A(n5242), .ZN(n5162) );
  INV_X1 U6324 ( .A(n5541), .ZN(n5156) );
  NAND2_X1 U6325 ( .A1(n7514), .A2(n7566), .ZN(n5761) );
  INV_X1 U6326 ( .A(n5303), .ZN(n5051) );
  INV_X1 U6327 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n5286) );
  XNOR2_X1 U6328 ( .A(n6724), .B(n4942), .ZN(n6720) );
  OR2_X1 U6329 ( .A1(n6091), .A2(n6090), .ZN(n6106) );
  NAND2_X1 U6330 ( .A1(n5844), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n6210) );
  OR2_X1 U6331 ( .A1(n6139), .A2(n6138), .ZN(n6165) );
  NAND2_X1 U6332 ( .A1(n5845), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n5889) );
  OR2_X1 U6333 ( .A1(n6122), .A2(n6121), .ZN(n6139) );
  AND2_X1 U6334 ( .A1(n8789), .A2(n8490), .ZN(n8491) );
  NAND2_X1 U6335 ( .A1(n5840), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n6122) );
  INV_X1 U6336 ( .A(n7704), .ZN(n7701) );
  INV_X1 U6337 ( .A(n5350), .ZN(n5158) );
  NAND2_X1 U6338 ( .A1(n6631), .A2(n6630), .ZN(n6632) );
  INV_X1 U6339 ( .A(n7985), .ZN(n6541) );
  INV_X1 U6340 ( .A(n5325), .ZN(n5159) );
  OR2_X1 U6341 ( .A1(n5225), .A2(n5224), .ZN(n5227) );
  NAND2_X1 U6342 ( .A1(n5162), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n5225) );
  NAND2_X1 U6343 ( .A1(n5160), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n5278) );
  OR2_X1 U6344 ( .A1(n5487), .A2(n5468), .ZN(n5521) );
  NAND2_X1 U6345 ( .A1(n5388), .A2(n4961), .ZN(n5132) );
  OR2_X1 U6346 ( .A1(n5561), .A2(n5560), .ZN(n5562) );
  NAND2_X1 U6347 ( .A1(n5842), .A2(n5841), .ZN(n6175) );
  OR2_X1 U6348 ( .A1(n5882), .A2(n8267), .ZN(n6238) );
  AND2_X1 U6349 ( .A1(n6329), .A2(n6382), .ZN(n8663) );
  INV_X1 U6350 ( .A(n9142), .ZN(n6706) );
  OR2_X1 U6351 ( .A1(n5336), .A2(n8930), .ZN(n5325) );
  OR2_X1 U6352 ( .A1(n5263), .A2(n9669), .ZN(n5265) );
  INV_X1 U6353 ( .A(n7721), .ZN(n6531) );
  NAND2_X1 U6354 ( .A1(n5159), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n5314) );
  INV_X1 U6355 ( .A(n8979), .ZN(n8995) );
  AND2_X1 U6356 ( .A1(n5227), .A2(n5226), .ZN(n9150) );
  OR2_X1 U6357 ( .A1(n5314), .A2(n5295), .ZN(n5297) );
  INV_X1 U6358 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n7102) );
  INV_X1 U6359 ( .A(n9091), .ZN(n9095) );
  INV_X1 U6360 ( .A(n9363), .ZN(n9175) );
  AND2_X1 U6361 ( .A1(n5677), .A2(n8072), .ZN(n9258) );
  AND2_X1 U6362 ( .A1(n5660), .A2(n7960), .ZN(n9827) );
  AOI21_X1 U6363 ( .B1(n9840), .B2(n7872), .A(n7871), .ZN(n7873) );
  OR2_X1 U6364 ( .A1(n7118), .A2(n6668), .ZN(n7368) );
  INV_X1 U6365 ( .A(n9959), .ZN(n9287) );
  INV_X1 U6366 ( .A(n10032), .ZN(n10010) );
  INV_X1 U6367 ( .A(n9010), .ZN(n9961) );
  OR2_X1 U6368 ( .A1(n7118), .A2(n7117), .ZN(n9960) );
  AND2_X1 U6369 ( .A1(n7375), .A2(n7374), .ZN(n9966) );
  AND2_X1 U6370 ( .A1(n5044), .A2(n5043), .ZN(n5330) );
  XNOR2_X1 U6371 ( .A(n5031), .B(SI_14_), .ZN(n5355) );
  NAND2_X1 U6372 ( .A1(n5003), .A2(n5002), .ZN(n5480) );
  AND2_X1 U6373 ( .A1(n6829), .A2(n6828), .ZN(n8315) );
  INV_X1 U6374 ( .A(n8317), .ZN(n8334) );
  AND4_X1 U6375 ( .A1(n6170), .A2(n6169), .A3(n6168), .A4(n6167), .ZN(n8718)
         );
  AND2_X1 U6376 ( .A1(n6964), .A2(n8857), .ZN(n10057) );
  INV_X1 U6377 ( .A(n8489), .ZN(n8621) );
  INV_X1 U6378 ( .A(n10089), .ZN(n8722) );
  NAND2_X1 U6379 ( .A1(n7693), .A2(n10096), .ZN(n10081) );
  INV_X1 U6380 ( .A(n10104), .ZN(n8749) );
  NAND2_X1 U6381 ( .A1(n8059), .A2(n7247), .ZN(n10194) );
  INV_X1 U6382 ( .A(n10199), .ZN(n10130) );
  NAND2_X1 U6383 ( .A1(n8717), .A2(n9806), .ZN(n10199) );
  AND2_X1 U6384 ( .A1(n6799), .A2(n6798), .ZN(n10109) );
  OR2_X1 U6385 ( .A1(n7121), .A2(n6668), .ZN(n10032) );
  INV_X1 U6386 ( .A(n8972), .ZN(n8991) );
  OR2_X1 U6387 ( .A1(n9136), .A2(n5302), .ZN(n5196) );
  INV_X1 U6388 ( .A(n4397), .ZN(n5282) );
  AND2_X1 U6389 ( .A1(n7006), .A2(n6838), .ZN(n9941) );
  INV_X1 U6390 ( .A(n9941), .ZN(n9886) );
  INV_X1 U6391 ( .A(n8112), .ZN(n9125) );
  AND2_X1 U6392 ( .A1(n8084), .A2(n5706), .ZN(n9154) );
  NAND2_X1 U6393 ( .A1(n9836), .A2(n7371), .ZN(n9972) );
  AND2_X1 U6394 ( .A1(n7361), .A2(n7521), .ZN(n7362) );
  AND2_X1 U6395 ( .A1(n6685), .A2(n7113), .ZN(n7203) );
  OR2_X1 U6396 ( .A1(n7121), .A2(n7398), .ZN(n10034) );
  OR2_X1 U6397 ( .A1(n7399), .A2(n7398), .ZN(n10015) );
  INV_X1 U6398 ( .A(n10030), .ZN(n9418) );
  NAND2_X1 U6399 ( .A1(n9966), .A2(n10015), .ZN(n10030) );
  INV_X1 U6400 ( .A(n10015), .ZN(n10039) );
  XNOR2_X1 U6401 ( .A(n4989), .B(SI_5_), .ZN(n5449) );
  NOR2_X1 U6402 ( .A1(n9781), .A2(n10261), .ZN(n9782) );
  INV_X1 U6403 ( .A(n8460), .ZN(n10058) );
  INV_X1 U6404 ( .A(n8800), .ZN(n8634) );
  NAND2_X1 U6405 ( .A1(n6829), .A2(n6813), .ZN(n8321) );
  OR2_X1 U6406 ( .A1(n6925), .A2(n6822), .ZN(n8340) );
  INV_X1 U6407 ( .A(n10056), .ZN(n10060) );
  INV_X1 U6408 ( .A(n10081), .ZN(n10104) );
  INV_X1 U6409 ( .A(n10081), .ZN(n10108) );
  NAND2_X1 U6410 ( .A1(n8749), .A2(n7735), .ZN(n8751) );
  OR2_X1 U6411 ( .A1(n7250), .A2(n7674), .ZN(n10217) );
  INV_X2 U6412 ( .A(n10217), .ZN(n10219) );
  OR2_X1 U6413 ( .A1(n7250), .A2(n7232), .ZN(n10200) );
  INV_X1 U6414 ( .A(n10114), .ZN(n10117) );
  INV_X1 U6415 ( .A(n6819), .ZN(n7552) );
  INV_X1 U6416 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n7012) );
  INV_X1 U6417 ( .A(n8992), .ZN(n8981) );
  INV_X1 U6418 ( .A(n8997), .ZN(n8985) );
  INV_X1 U6419 ( .A(n9127), .ZN(n9002) );
  OR2_X1 U6420 ( .A1(P1_U3083), .A2(n6860), .ZN(n9945) );
  INV_X1 U6421 ( .A(n9109), .ZN(n9308) );
  AND2_X1 U6422 ( .A1(n9249), .A2(n7479), .ZN(n9970) );
  AND2_X1 U6423 ( .A1(n9862), .A2(n9861), .ZN(n9876) );
  INV_X1 U6424 ( .A(n10042), .ZN(n10040) );
  INV_X1 U6425 ( .A(n9984), .ZN(n9985) );
  INV_X1 U6426 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n9696) );
  INV_X1 U6427 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n6910) );
  INV_X1 U6428 ( .A(n9730), .ZN(n9449) );
  AND2_X1 U6429 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n4969) );
  NAND2_X1 U6430 ( .A1(n4975), .A2(n4969), .ZN(n5386) );
  AND2_X1 U6431 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n4970) );
  NAND2_X1 U6432 ( .A1(n5386), .A2(n5975), .ZN(n4971) );
  NAND2_X1 U6433 ( .A1(n4971), .A2(SI_1_), .ZN(n4972) );
  INV_X1 U6434 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n4973) );
  XNOR2_X1 U6435 ( .A(n4977), .B(SI_2_), .ZN(n5421) );
  INV_X1 U6436 ( .A(n5421), .ZN(n4976) );
  NAND2_X1 U6437 ( .A1(n4977), .A2(SI_2_), .ZN(n4978) );
  NAND2_X1 U6438 ( .A1(n4979), .A2(n4978), .ZN(n5400) );
  NAND2_X1 U6439 ( .A1(n5400), .A2(n4981), .ZN(n4984) );
  NAND2_X1 U6440 ( .A1(n4982), .A2(SI_3_), .ZN(n4983) );
  NAND2_X1 U6441 ( .A1(n4984), .A2(n4983), .ZN(n5411) );
  MUX2_X1 U6442 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .S(n4975), .Z(n4986) );
  NAND2_X1 U6443 ( .A1(n5411), .A2(n4985), .ZN(n4988) );
  NAND2_X1 U6444 ( .A1(n4986), .A2(SI_4_), .ZN(n4987) );
  NAND2_X1 U6445 ( .A1(n4988), .A2(n4987), .ZN(n5448) );
  MUX2_X1 U6446 ( .A(n6898), .B(n6889), .S(n6891), .Z(n4989) );
  NAND2_X1 U6447 ( .A1(n5448), .A2(n5449), .ZN(n4992) );
  INV_X1 U6448 ( .A(n4989), .ZN(n4990) );
  NAND2_X1 U6449 ( .A1(n4990), .A2(SI_5_), .ZN(n4991) );
  MUX2_X1 U6450 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n6891), .Z(n4994) );
  NAND2_X1 U6451 ( .A1(n5435), .A2(n4993), .ZN(n4996) );
  NAND2_X1 U6452 ( .A1(n4994), .A2(SI_6_), .ZN(n4995) );
  MUX2_X1 U6453 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n6891), .Z(n4998) );
  NAND2_X1 U6454 ( .A1(n4998), .A2(SI_7_), .ZN(n4999) );
  MUX2_X1 U6455 ( .A(n6906), .B(n6908), .S(n6891), .Z(n5000) );
  INV_X1 U6456 ( .A(n5000), .ZN(n5001) );
  NAND2_X1 U6457 ( .A1(n5001), .A2(SI_8_), .ZN(n5002) );
  MUX2_X1 U6458 ( .A(n6912), .B(n6910), .S(n6891), .Z(n5005) );
  INV_X1 U6459 ( .A(SI_9_), .ZN(n5004) );
  NAND2_X1 U6460 ( .A1(n5005), .A2(n5004), .ZN(n5008) );
  INV_X1 U6461 ( .A(n5005), .ZN(n5006) );
  NAND2_X1 U6462 ( .A1(n5006), .A2(SI_9_), .ZN(n5007) );
  MUX2_X1 U6463 ( .A(n6918), .B(n6916), .S(n6891), .Z(n5011) );
  INV_X1 U6464 ( .A(SI_10_), .ZN(n5010) );
  NAND2_X1 U6465 ( .A1(n5011), .A2(n5010), .ZN(n5014) );
  INV_X1 U6466 ( .A(n5011), .ZN(n5012) );
  NAND2_X1 U6467 ( .A1(n5012), .A2(SI_10_), .ZN(n5013) );
  MUX2_X1 U6468 ( .A(n9644), .B(n6920), .S(n6891), .Z(n5015) );
  XNOR2_X1 U6469 ( .A(n5015), .B(SI_11_), .ZN(n5528) );
  INV_X1 U6470 ( .A(n5528), .ZN(n5017) );
  INV_X1 U6471 ( .A(n5015), .ZN(n5016) );
  MUX2_X1 U6472 ( .A(n7012), .B(n9696), .S(n6891), .Z(n5019) );
  INV_X1 U6473 ( .A(SI_12_), .ZN(n5018) );
  INV_X1 U6474 ( .A(n5019), .ZN(n5020) );
  NAND2_X1 U6475 ( .A1(n5020), .A2(SI_12_), .ZN(n5021) );
  NAND2_X1 U6476 ( .A1(n5022), .A2(n5021), .ZN(n5506) );
  INV_X1 U6477 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n7041) );
  INV_X1 U6478 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n5023) );
  MUX2_X1 U6479 ( .A(n7041), .B(n5023), .S(n6891), .Z(n5025) );
  INV_X1 U6480 ( .A(SI_13_), .ZN(n5024) );
  NAND2_X1 U6481 ( .A1(n5025), .A2(n5024), .ZN(n5028) );
  INV_X1 U6482 ( .A(n5025), .ZN(n5026) );
  NAND2_X1 U6483 ( .A1(n5026), .A2(SI_13_), .ZN(n5027) );
  NAND2_X1 U6484 ( .A1(n5367), .A2(n4963), .ZN(n5029) );
  INV_X1 U6485 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n7125) );
  INV_X1 U6486 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n5030) );
  MUX2_X1 U6487 ( .A(n7125), .B(n5030), .S(n6891), .Z(n5031) );
  INV_X1 U6488 ( .A(n5031), .ZN(n5032) );
  NAND2_X1 U6489 ( .A1(n5032), .A2(SI_14_), .ZN(n5033) );
  INV_X1 U6490 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n7163) );
  INV_X1 U6491 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n7161) );
  MUX2_X1 U6492 ( .A(n7163), .B(n7161), .S(n6891), .Z(n5035) );
  INV_X1 U6493 ( .A(SI_15_), .ZN(n5034) );
  INV_X1 U6494 ( .A(n5035), .ZN(n5036) );
  NAND2_X1 U6495 ( .A1(n5036), .A2(SI_15_), .ZN(n5037) );
  INV_X1 U6496 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n5039) );
  MUX2_X1 U6497 ( .A(n5039), .B(n9593), .S(n6891), .Z(n5041) );
  INV_X1 U6498 ( .A(SI_16_), .ZN(n5040) );
  NAND2_X1 U6499 ( .A1(n5041), .A2(n5040), .ZN(n5044) );
  INV_X1 U6500 ( .A(n5041), .ZN(n5042) );
  NAND2_X1 U6501 ( .A1(n5042), .A2(SI_16_), .ZN(n5043) );
  NAND2_X1 U6502 ( .A1(n5045), .A2(n5044), .ZN(n5320) );
  INV_X1 U6503 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n5046) );
  MUX2_X1 U6504 ( .A(n9695), .B(n5046), .S(n6891), .Z(n5047) );
  XNOR2_X1 U6505 ( .A(n5047), .B(SI_17_), .ZN(n5319) );
  INV_X1 U6506 ( .A(n5047), .ZN(n5048) );
  NAND2_X1 U6507 ( .A1(n5048), .A2(SI_17_), .ZN(n5049) );
  OAI21_X1 U6508 ( .B1(n5320), .B2(n5050), .A(n5049), .ZN(n5304) );
  MUX2_X1 U6509 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n6891), .Z(n5052) );
  XNOR2_X1 U6510 ( .A(n5052), .B(SI_18_), .ZN(n5303) );
  NAND2_X1 U6511 ( .A1(n5052), .A2(SI_18_), .ZN(n5053) );
  INV_X1 U6512 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n8123) );
  INV_X1 U6513 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7350) );
  MUX2_X1 U6514 ( .A(n8123), .B(n7350), .S(n6891), .Z(n5055) );
  INV_X1 U6515 ( .A(SI_19_), .ZN(n5054) );
  NAND2_X1 U6516 ( .A1(n5055), .A2(n5054), .ZN(n5058) );
  INV_X1 U6517 ( .A(n5055), .ZN(n5056) );
  NAND2_X1 U6518 ( .A1(n5056), .A2(SI_19_), .ZN(n5057) );
  NAND2_X1 U6519 ( .A1(n5058), .A2(n5057), .ZN(n5283) );
  INV_X1 U6520 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n8061) );
  INV_X1 U6521 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n9604) );
  MUX2_X1 U6522 ( .A(n8061), .B(n9604), .S(n6891), .Z(n5060) );
  INV_X1 U6523 ( .A(SI_20_), .ZN(n5059) );
  NAND2_X1 U6524 ( .A1(n5060), .A2(n5059), .ZN(n5063) );
  INV_X1 U6525 ( .A(n5060), .ZN(n5061) );
  NAND2_X1 U6526 ( .A1(n5061), .A2(SI_20_), .ZN(n5062) );
  NAND2_X1 U6527 ( .A1(n5064), .A2(n5063), .ZN(n5251) );
  INV_X1 U6528 ( .A(n5251), .ZN(n5065) );
  INV_X1 U6529 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7553) );
  INV_X1 U6530 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n9556) );
  MUX2_X1 U6531 ( .A(n7553), .B(n9556), .S(n6891), .Z(n5066) );
  XNOR2_X1 U6532 ( .A(n5066), .B(SI_21_), .ZN(n5250) );
  NAND2_X1 U6533 ( .A1(n5065), .A2(n5250), .ZN(n5069) );
  INV_X1 U6534 ( .A(n5066), .ZN(n5067) );
  NAND2_X1 U6535 ( .A1(n5067), .A2(SI_21_), .ZN(n5068) );
  INV_X1 U6536 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7663) );
  INV_X1 U6537 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n8063) );
  MUX2_X1 U6538 ( .A(n7663), .B(n8063), .S(n6891), .Z(n5071) );
  INV_X1 U6539 ( .A(SI_22_), .ZN(n5070) );
  NAND2_X1 U6540 ( .A1(n5071), .A2(n5070), .ZN(n5074) );
  INV_X1 U6541 ( .A(n5071), .ZN(n5072) );
  NAND2_X1 U6542 ( .A1(n5072), .A2(SI_22_), .ZN(n5073) );
  NAND2_X1 U6543 ( .A1(n5074), .A2(n5073), .ZN(n5258) );
  INV_X1 U6544 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n5075) );
  INV_X1 U6545 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n7732) );
  MUX2_X1 U6546 ( .A(n5075), .B(n7732), .S(n6891), .Z(n5077) );
  INV_X1 U6547 ( .A(SI_23_), .ZN(n5076) );
  NAND2_X1 U6548 ( .A1(n5077), .A2(n5076), .ZN(n5080) );
  INV_X1 U6549 ( .A(n5077), .ZN(n5078) );
  NAND2_X1 U6550 ( .A1(n5078), .A2(SI_23_), .ZN(n5079) );
  INV_X1 U6551 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n9671) );
  INV_X1 U6552 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7942) );
  MUX2_X1 U6553 ( .A(n9671), .B(n7942), .S(n6891), .Z(n5081) );
  XNOR2_X1 U6554 ( .A(n5081), .B(SI_24_), .ZN(n5209) );
  INV_X1 U6555 ( .A(n5209), .ZN(n5084) );
  INV_X1 U6556 ( .A(n5081), .ZN(n5082) );
  NAND2_X1 U6557 ( .A1(n5082), .A2(SI_24_), .ZN(n5083) );
  INV_X1 U6558 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n8012) );
  INV_X1 U6559 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n9542) );
  MUX2_X1 U6560 ( .A(n8012), .B(n9542), .S(n6891), .Z(n5085) );
  INV_X1 U6561 ( .A(SI_25_), .ZN(n9622) );
  NAND2_X1 U6562 ( .A1(n5085), .A2(n9622), .ZN(n5088) );
  INV_X1 U6563 ( .A(n5085), .ZN(n5086) );
  NAND2_X1 U6564 ( .A1(n5086), .A2(SI_25_), .ZN(n5087) );
  NAND2_X1 U6565 ( .A1(n5088), .A2(n5087), .ZN(n5220) );
  INV_X1 U6566 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n8041) );
  INV_X1 U6567 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n8045) );
  MUX2_X1 U6568 ( .A(n8041), .B(n8045), .S(n6891), .Z(n5090) );
  INV_X1 U6569 ( .A(SI_26_), .ZN(n5089) );
  NAND2_X1 U6570 ( .A1(n5090), .A2(n5089), .ZN(n5093) );
  INV_X1 U6571 ( .A(n5090), .ZN(n5091) );
  NAND2_X1 U6572 ( .A1(n5091), .A2(SI_26_), .ZN(n5092) );
  INV_X1 U6573 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n9684) );
  INV_X1 U6574 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n5199) );
  MUX2_X1 U6575 ( .A(n9684), .B(n5199), .S(n6891), .Z(n5094) );
  INV_X1 U6576 ( .A(SI_27_), .ZN(n9553) );
  NAND2_X1 U6577 ( .A1(n5094), .A2(n9553), .ZN(n5097) );
  INV_X1 U6578 ( .A(n5094), .ZN(n5095) );
  NAND2_X1 U6579 ( .A1(n5095), .A2(SI_27_), .ZN(n5096) );
  AND2_X1 U6580 ( .A1(n5097), .A2(n5096), .ZN(n5198) );
  NAND2_X1 U6581 ( .A1(n5197), .A2(n5198), .ZN(n5098) );
  INV_X1 U6582 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n5099) );
  INV_X1 U6583 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n5175) );
  MUX2_X1 U6584 ( .A(n5099), .B(n5175), .S(n4975), .Z(n5101) );
  XNOR2_X1 U6585 ( .A(n5101), .B(SI_28_), .ZN(n5173) );
  NAND2_X1 U6586 ( .A1(n5174), .A2(n5173), .ZN(n5103) );
  INV_X1 U6587 ( .A(SI_28_), .ZN(n5100) );
  NAND2_X1 U6588 ( .A1(n5101), .A2(n5100), .ZN(n5102) );
  NAND2_X1 U6589 ( .A1(n5103), .A2(n5102), .ZN(n5150) );
  INV_X1 U6590 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n5104) );
  INV_X1 U6591 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n9448) );
  MUX2_X1 U6592 ( .A(n5104), .B(n9448), .S(n4975), .Z(n5148) );
  INV_X1 U6593 ( .A(SI_29_), .ZN(n5105) );
  AND2_X1 U6594 ( .A1(n5148), .A2(n5105), .ZN(n5108) );
  INV_X1 U6595 ( .A(n5148), .ZN(n5106) );
  NAND2_X1 U6596 ( .A1(n5106), .A2(SI_29_), .ZN(n5107) );
  OAI21_X1 U6597 ( .B1(n5150), .B2(n5108), .A(n5107), .ZN(n5110) );
  MUX2_X1 U6598 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(P2_DATAO_REG_30__SCAN_IN), 
        .S(n6891), .Z(n5111) );
  XNOR2_X1 U6599 ( .A(n5110), .B(n5111), .ZN(n5143) );
  INV_X1 U6600 ( .A(n5143), .ZN(n5109) );
  NAND2_X1 U6601 ( .A1(n5109), .A2(SI_30_), .ZN(n5113) );
  NAND2_X1 U6602 ( .A1(n5110), .A2(n5111), .ZN(n5112) );
  NAND2_X1 U6603 ( .A1(n5113), .A2(n5112), .ZN(n5116) );
  MUX2_X1 U6604 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .S(n4975), .Z(n5114) );
  XNOR2_X1 U6605 ( .A(n5114), .B(SI_31_), .ZN(n5115) );
  INV_X1 U6606 ( .A(n8845), .ZN(n5133) );
  NOR2_X1 U6607 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), .ZN(
        n5123) );
  NOR2_X1 U6608 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n5122) );
  NOR2_X1 U6609 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n5121) );
  NOR2_X1 U6610 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_IR_REG_20__SCAN_IN), .ZN(
        n5120) );
  NAND4_X1 U6611 ( .A1(n5123), .A2(n5122), .A3(n5121), .A4(n5120), .ZN(n5126)
         );
  NOR2_X1 U6612 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n5288) );
  NOR2_X1 U6613 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n5287) );
  NOR2_X1 U6614 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n5124) );
  NAND3_X1 U6615 ( .A1(n5288), .A2(n5287), .A3(n5124), .ZN(n5125) );
  NAND2_X1 U6616 ( .A1(n5134), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5131) );
  NAND2_X1 U6617 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), 
        .ZN(n5128) );
  NAND2_X1 U6618 ( .A1(n5131), .A2(n5128), .ZN(n5129) );
  INV_X1 U6619 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5130) );
  NAND2_X1 U6620 ( .A1(n5136), .A2(P1_IR_REG_29__SCAN_IN), .ZN(n5135) );
  INV_X1 U6621 ( .A(n5137), .ZN(n5139) );
  NOR2_X1 U6622 ( .A1(P1_IR_REG_27__SCAN_IN), .A2(P1_IR_REG_29__SCAN_IN), .ZN(
        n5138) );
  NAND2_X1 U6623 ( .A1(n5139), .A2(n5138), .ZN(n9438) );
  NAND2_X1 U6624 ( .A1(n4397), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n5142) );
  NAND2_X1 U6625 ( .A1(n5543), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n5141) );
  INV_X1 U6626 ( .A(n5453), .ZN(n5488) );
  NAND2_X1 U6627 ( .A1(n5453), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n5140) );
  AND3_X1 U6628 ( .A1(n5142), .A2(n5141), .A3(n5140), .ZN(n5722) );
  INV_X1 U6629 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n9571) );
  NOR2_X1 U6630 ( .A1(n5464), .A2(n9571), .ZN(n5144) );
  NAND2_X1 U6631 ( .A1(n4397), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n5147) );
  NAND2_X1 U6632 ( .A1(n5523), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n5146) );
  NAND2_X1 U6633 ( .A1(n5543), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n5145) );
  NAND3_X1 U6634 ( .A1(n5147), .A2(n5146), .A3(n5145), .ZN(n9001) );
  XNOR2_X1 U6635 ( .A(n5148), .B(SI_29_), .ZN(n5149) );
  NAND2_X1 U6636 ( .A1(n8852), .A2(n4613), .ZN(n5152) );
  OR2_X1 U6637 ( .A1(n5464), .A2(n9448), .ZN(n5151) );
  NAND2_X1 U6638 ( .A1(n5423), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5494) );
  INV_X1 U6639 ( .A(n5494), .ZN(n5153) );
  NAND2_X1 U6640 ( .A1(n5153), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5496) );
  INV_X1 U6641 ( .A(n5496), .ZN(n5154) );
  NAND2_X1 U6642 ( .A1(n5154), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n5487) );
  INV_X1 U6643 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n5373) );
  INV_X1 U6644 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n5348) );
  INV_X1 U6645 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n8930) );
  INV_X1 U6646 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n5295) );
  INV_X1 U6647 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n8903) );
  INV_X1 U6648 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n9669) );
  INV_X1 U6649 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n5224) );
  NAND2_X1 U6650 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(P1_REG3_REG_28__SCAN_IN), 
        .ZN(n5164) );
  NAND2_X1 U6651 ( .A1(n4397), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n5170) );
  NAND2_X1 U6652 ( .A1(n5523), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n5169) );
  INV_X2 U6653 ( .A(n5167), .ZN(n5543) );
  NAND2_X1 U6654 ( .A1(n5543), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n5168) );
  AND3_X1 U6655 ( .A1(n5170), .A2(n5169), .A3(n5168), .ZN(n5171) );
  OAI21_X1 U6656 ( .B1(n8115), .B2(n5302), .A(n5171), .ZN(n9105) );
  INV_X1 U6657 ( .A(n9105), .ZN(n5172) );
  NAND2_X1 U6658 ( .A1(n9336), .A2(n5172), .ZN(n5733) );
  NAND2_X1 U6659 ( .A1(n8855), .A2(n4613), .ZN(n5177) );
  OR2_X1 U6660 ( .A1(n5464), .A2(n5175), .ZN(n5176) );
  INV_X1 U6661 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n5179) );
  INV_X1 U6662 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n5178) );
  OAI21_X1 U6663 ( .B1(n5202), .B2(n5179), .A(n5178), .ZN(n5180) );
  NAND2_X1 U6664 ( .A1(n9111), .A2(n4391), .ZN(n5186) );
  INV_X1 U6665 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n5183) );
  NAND2_X1 U6666 ( .A1(n5523), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n5182) );
  NAND2_X1 U6667 ( .A1(n5543), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n5181) );
  OAI211_X1 U6668 ( .C1(n5183), .C2(n5282), .A(n5182), .B(n5181), .ZN(n5184)
         );
  INV_X1 U6669 ( .A(n5184), .ZN(n5185) );
  NAND2_X1 U6670 ( .A1(n9341), .A2(n9127), .ZN(n8086) );
  OR2_X1 U6671 ( .A1(n5464), .A2(n8045), .ZN(n5189) );
  INV_X1 U6672 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n9608) );
  NAND2_X1 U6673 ( .A1(n5227), .A2(n9608), .ZN(n5191) );
  NAND2_X1 U6674 ( .A1(n5202), .A2(n5191), .ZN(n9136) );
  INV_X1 U6675 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n9519) );
  NAND2_X1 U6676 ( .A1(n5543), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n5193) );
  NAND2_X1 U6677 ( .A1(n5453), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n5192) );
  OAI211_X1 U6678 ( .C1(n5282), .C2(n9519), .A(n5193), .B(n5192), .ZN(n5194)
         );
  INV_X1 U6679 ( .A(n5194), .ZN(n5195) );
  OR2_X1 U6680 ( .A1(n5464), .A2(n5199), .ZN(n5200) );
  XNOR2_X1 U6681 ( .A(n5202), .B(P1_REG3_REG_27__SCAN_IN), .ZN(n9120) );
  NAND2_X1 U6682 ( .A1(n9120), .A2(n5542), .ZN(n5207) );
  INV_X1 U6683 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n9634) );
  NAND2_X1 U6684 ( .A1(n5453), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n5204) );
  NAND2_X1 U6685 ( .A1(n5543), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n5203) );
  OAI211_X1 U6686 ( .C1(n5282), .C2(n9634), .A(n5204), .B(n5203), .ZN(n5205)
         );
  INV_X1 U6687 ( .A(n5205), .ZN(n5206) );
  NAND2_X1 U6688 ( .A1(n9346), .A2(n6706), .ZN(n5730) );
  NAND2_X1 U6689 ( .A1(n7938), .A2(n4613), .ZN(n5211) );
  OR2_X1 U6690 ( .A1(n5464), .A2(n7942), .ZN(n5210) );
  INV_X1 U6691 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n5212) );
  NAND2_X1 U6692 ( .A1(n5242), .A2(n5212), .ZN(n5213) );
  NAND2_X1 U6693 ( .A1(n5225), .A2(n5213), .ZN(n9171) );
  INV_X1 U6694 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n5216) );
  NAND2_X1 U6695 ( .A1(n5543), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n5215) );
  NAND2_X1 U6696 ( .A1(n5523), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n5214) );
  OAI211_X1 U6697 ( .C1(n5282), .C2(n5216), .A(n5215), .B(n5214), .ZN(n5217)
         );
  INV_X1 U6698 ( .A(n5217), .ZN(n5218) );
  NAND2_X1 U6699 ( .A1(n9363), .A2(n8110), .ZN(n5569) );
  NAND2_X1 U6700 ( .A1(n8010), .A2(n4613), .ZN(n5223) );
  OR2_X1 U6701 ( .A1(n5464), .A2(n9542), .ZN(n5222) );
  NAND2_X1 U6702 ( .A1(n5225), .A2(n5224), .ZN(n5226) );
  NAND2_X1 U6703 ( .A1(n9150), .A2(n4391), .ZN(n5232) );
  INV_X1 U6704 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n9673) );
  NAND2_X1 U6705 ( .A1(n5523), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n5229) );
  NAND2_X1 U6706 ( .A1(n5543), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n5228) );
  OAI211_X1 U6707 ( .C1(n9673), .C2(n5282), .A(n5229), .B(n5228), .ZN(n5230)
         );
  INV_X1 U6708 ( .A(n5230), .ZN(n5231) );
  INV_X1 U6709 ( .A(n9166), .ZN(n5233) );
  NAND2_X1 U6710 ( .A1(n9356), .A2(n5233), .ZN(n5706) );
  OR2_X1 U6711 ( .A1(n5235), .A2(n5234), .ZN(n5236) );
  NAND2_X1 U6712 ( .A1(n5237), .A2(n5236), .ZN(n7729) );
  NAND2_X1 U6713 ( .A1(n7729), .A2(n4613), .ZN(n5239) );
  OR2_X1 U6714 ( .A1(n5464), .A2(n7732), .ZN(n5238) );
  INV_X1 U6715 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n5240) );
  NAND2_X1 U6716 ( .A1(n5265), .A2(n5240), .ZN(n5241) );
  NAND2_X1 U6717 ( .A1(n5242), .A2(n5241), .ZN(n9180) );
  OR2_X1 U6718 ( .A1(n9180), .A2(n5302), .ZN(n5248) );
  INV_X1 U6719 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n5245) );
  NAND2_X1 U6720 ( .A1(n5543), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n5244) );
  NAND2_X1 U6721 ( .A1(n5523), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n5243) );
  OAI211_X1 U6722 ( .C1(n5282), .C2(n5245), .A(n5244), .B(n5243), .ZN(n5246)
         );
  INV_X1 U6723 ( .A(n5246), .ZN(n5247) );
  NAND2_X1 U6724 ( .A1(n5248), .A2(n5247), .ZN(n9203) );
  INV_X1 U6725 ( .A(n9203), .ZN(n5249) );
  NAND2_X1 U6726 ( .A1(n9366), .A2(n5249), .ZN(n5608) );
  NAND2_X1 U6727 ( .A1(n8082), .A2(n5608), .ZN(n9187) );
  XNOR2_X1 U6728 ( .A(n5251), .B(n5250), .ZN(n7551) );
  NAND2_X1 U6729 ( .A1(n7551), .A2(n4613), .ZN(n5253) );
  OR2_X1 U6730 ( .A1(n5464), .A2(n9556), .ZN(n5252) );
  INV_X1 U6731 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n5257) );
  NAND2_X1 U6732 ( .A1(n5278), .A2(n8903), .ZN(n5254) );
  NAND2_X1 U6733 ( .A1(n5263), .A2(n5254), .ZN(n9219) );
  OR2_X1 U6734 ( .A1(n9219), .A2(n5302), .ZN(n5256) );
  AOI22_X1 U6735 ( .A1(n4397), .A2(P1_REG1_REG_21__SCAN_IN), .B1(n5523), .B2(
        P1_REG2_REG_21__SCAN_IN), .ZN(n5255) );
  OAI211_X1 U6736 ( .C1(n5167), .C2(n5257), .A(n5256), .B(n5255), .ZN(n9236)
         );
  INV_X1 U6737 ( .A(n9236), .ZN(n8960) );
  NAND2_X1 U6738 ( .A1(n9378), .A2(n8960), .ZN(n8077) );
  NAND2_X1 U6739 ( .A1(n5690), .A2(n8077), .ZN(n9213) );
  NAND2_X1 U6740 ( .A1(n5259), .A2(n5258), .ZN(n5260) );
  NAND2_X1 U6741 ( .A1(n4960), .A2(n5260), .ZN(n7661) );
  NAND2_X1 U6742 ( .A1(n7661), .A2(n4613), .ZN(n5262) );
  OR2_X1 U6743 ( .A1(n5464), .A2(n8063), .ZN(n5261) );
  NAND2_X1 U6744 ( .A1(n5263), .A2(n9669), .ZN(n5264) );
  AND2_X1 U6745 ( .A1(n5265), .A2(n5264), .ZN(n9197) );
  NAND2_X1 U6746 ( .A1(n9197), .A2(n5542), .ZN(n5271) );
  INV_X1 U6747 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n5268) );
  NAND2_X1 U6748 ( .A1(n5543), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n5267) );
  NAND2_X1 U6749 ( .A1(n5523), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n5266) );
  OAI211_X1 U6750 ( .C1(n5282), .C2(n5268), .A(n5267), .B(n5266), .ZN(n5269)
         );
  INV_X1 U6751 ( .A(n5269), .ZN(n5270) );
  NAND2_X1 U6752 ( .A1(n5271), .A2(n5270), .ZN(n9190) );
  INV_X1 U6753 ( .A(n9190), .ZN(n9215) );
  NAND2_X1 U6754 ( .A1(n9371), .A2(n9215), .ZN(n8079) );
  NAND2_X1 U6755 ( .A1(n8078), .A2(n8079), .ZN(n9201) );
  XNOR2_X1 U6756 ( .A(n5273), .B(n5272), .ZN(n7493) );
  NAND2_X1 U6757 ( .A1(n7493), .A2(n4613), .ZN(n5275) );
  OR2_X1 U6758 ( .A1(n5464), .A2(n9604), .ZN(n5274) );
  INV_X1 U6759 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n5281) );
  INV_X1 U6760 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n5276) );
  NAND2_X1 U6761 ( .A1(n5297), .A2(n5276), .ZN(n5277) );
  NAND2_X1 U6762 ( .A1(n5278), .A2(n5277), .ZN(n9229) );
  OR2_X1 U6763 ( .A1(n9229), .A2(n5302), .ZN(n5280) );
  AOI22_X1 U6764 ( .A1(n5543), .A2(P1_REG0_REG_20__SCAN_IN), .B1(n5523), .B2(
        P1_REG2_REG_20__SCAN_IN), .ZN(n5279) );
  OAI211_X1 U6765 ( .C1(n5282), .C2(n5281), .A(n5280), .B(n5279), .ZN(n9003)
         );
  INV_X1 U6766 ( .A(n9003), .ZN(n9246) );
  AND2_X1 U6767 ( .A1(n9381), .A2(n9246), .ZN(n8074) );
  NOR2_X1 U6768 ( .A1(n9381), .A2(n9246), .ZN(n8075) );
  NOR2_X1 U6769 ( .A1(n8074), .A2(n8075), .ZN(n9233) );
  XNOR2_X1 U6770 ( .A(n5284), .B(n5283), .ZN(n7349) );
  NAND2_X1 U6771 ( .A1(n7349), .A2(n4613), .ZN(n5294) );
  INV_X1 U6772 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5289) );
  INV_X1 U6773 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n5305) );
  INV_X1 U6774 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5307) );
  INV_X1 U6775 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n5290) );
  NAND2_X1 U6776 ( .A1(n5558), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5292) );
  INV_X1 U6777 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5291) );
  AOI22_X1 U6778 ( .A1(n5535), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n9250), .B2(
        n5534), .ZN(n5293) );
  NAND2_X1 U6779 ( .A1(n5314), .A2(n5295), .ZN(n5296) );
  NAND2_X1 U6780 ( .A1(n5297), .A2(n5296), .ZN(n9248) );
  NAND2_X1 U6781 ( .A1(n5523), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n5299) );
  NAND2_X1 U6782 ( .A1(n5543), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n5298) );
  AND2_X1 U6783 ( .A1(n5299), .A2(n5298), .ZN(n5301) );
  NAND2_X1 U6784 ( .A1(n4397), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n5300) );
  OAI211_X1 U6785 ( .C1(n9248), .C2(n5302), .A(n5301), .B(n5300), .ZN(n9237)
         );
  INV_X1 U6786 ( .A(n9237), .ZN(n9264) );
  OR2_X1 U6787 ( .A1(n9388), .A2(n9264), .ZN(n5679) );
  NAND2_X1 U6788 ( .A1(n9388), .A2(n9264), .ZN(n8073) );
  XNOR2_X1 U6789 ( .A(n5304), .B(n5303), .ZN(n7296) );
  NAND2_X1 U6790 ( .A1(n7296), .A2(n4613), .ZN(n5311) );
  NAND2_X1 U6791 ( .A1(n4470), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5332) );
  NAND2_X1 U6792 ( .A1(n5332), .A2(n5305), .ZN(n5306) );
  NAND2_X1 U6793 ( .A1(n5306), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5321) );
  NAND2_X1 U6794 ( .A1(n5321), .A2(n5307), .ZN(n5308) );
  NAND2_X1 U6795 ( .A1(n5308), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5309) );
  XNOR2_X1 U6796 ( .A(n5309), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9080) );
  AOI22_X1 U6797 ( .A1(n5535), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n9080), .B2(
        n5534), .ZN(n5310) );
  INV_X1 U6798 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n5312) );
  NAND2_X1 U6799 ( .A1(n5325), .A2(n5312), .ZN(n5313) );
  AND2_X1 U6800 ( .A1(n5314), .A2(n5313), .ZN(n9268) );
  NAND2_X1 U6801 ( .A1(n4391), .A2(n9268), .ZN(n5318) );
  NAND2_X1 U6802 ( .A1(n4397), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n5317) );
  NAND2_X1 U6803 ( .A1(n5523), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n5316) );
  NAND2_X1 U6804 ( .A1(n5543), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n5315) );
  NAND4_X1 U6805 ( .A1(n5318), .A2(n5317), .A3(n5316), .A4(n5315), .ZN(n9286)
         );
  INV_X1 U6806 ( .A(n9286), .ZN(n9244) );
  OR2_X1 U6807 ( .A1(n9269), .A2(n9244), .ZN(n5677) );
  NAND2_X1 U6808 ( .A1(n9269), .A2(n9244), .ZN(n8072) );
  XNOR2_X1 U6809 ( .A(n5320), .B(n5319), .ZN(n7208) );
  NAND2_X1 U6810 ( .A1(n7208), .A2(n4613), .ZN(n5323) );
  XNOR2_X1 U6811 ( .A(n5321), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9069) );
  AOI22_X1 U6812 ( .A1(n5535), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n5534), .B2(
        n9069), .ZN(n5322) );
  NAND2_X1 U6813 ( .A1(n4397), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n5329) );
  NAND2_X1 U6814 ( .A1(n5336), .A2(n8930), .ZN(n5324) );
  AND2_X1 U6815 ( .A1(n5325), .A2(n5324), .ZN(n9279) );
  NAND2_X1 U6816 ( .A1(n4391), .A2(n9279), .ZN(n5328) );
  NAND2_X1 U6817 ( .A1(n5523), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n5327) );
  NAND2_X1 U6818 ( .A1(n5543), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n5326) );
  NAND4_X1 U6819 ( .A1(n5329), .A2(n5328), .A3(n5327), .A4(n5326), .ZN(n9004)
         );
  INV_X1 U6820 ( .A(n9004), .ZN(n9299) );
  OR2_X1 U6821 ( .A1(n9398), .A2(n9299), .ZN(n8070) );
  NAND2_X1 U6822 ( .A1(n9398), .A2(n9299), .ZN(n9260) );
  NAND2_X1 U6823 ( .A1(n8070), .A2(n9260), .ZN(n9275) );
  XNOR2_X1 U6824 ( .A(n5331), .B(n5330), .ZN(n7158) );
  NAND2_X1 U6825 ( .A1(n7158), .A2(n4613), .ZN(n5334) );
  XNOR2_X1 U6826 ( .A(n5332), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9053) );
  AOI22_X1 U6827 ( .A1(n5535), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n5534), .B2(
        n9053), .ZN(n5333) );
  NAND2_X1 U6828 ( .A1(n4397), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n5340) );
  INV_X1 U6829 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n8921) );
  NAND2_X1 U6830 ( .A1(n5350), .A2(n8921), .ZN(n5335) );
  AND2_X1 U6831 ( .A1(n5336), .A2(n5335), .ZN(n9302) );
  NAND2_X1 U6832 ( .A1(n4391), .A2(n9302), .ZN(n5339) );
  NAND2_X1 U6833 ( .A1(n5523), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n5338) );
  NAND2_X1 U6834 ( .A1(n5543), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n5337) );
  NAND4_X1 U6835 ( .A1(n5340), .A2(n5339), .A3(n5338), .A4(n5337), .ZN(n9288)
         );
  INV_X1 U6836 ( .A(n9288), .ZN(n9311) );
  OR2_X1 U6837 ( .A1(n9405), .A2(n9311), .ZN(n5668) );
  NAND2_X1 U6838 ( .A1(n9405), .A2(n9311), .ZN(n8069) );
  NAND2_X1 U6839 ( .A1(n5668), .A2(n8069), .ZN(n9296) );
  XNOR2_X1 U6840 ( .A(n5342), .B(n5341), .ZN(n7160) );
  NAND2_X1 U6841 ( .A1(n7160), .A2(n4613), .ZN(n5347) );
  NAND2_X1 U6842 ( .A1(n5343), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5344) );
  XNOR2_X1 U6843 ( .A(n5344), .B(n4784), .ZN(n9036) );
  INV_X1 U6844 ( .A(n9036), .ZN(n5345) );
  AOI22_X1 U6845 ( .A1(n5535), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n5534), .B2(
        n5345), .ZN(n5346) );
  NAND2_X1 U6846 ( .A1(n4397), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n5354) );
  NAND2_X1 U6847 ( .A1(n5362), .A2(n5348), .ZN(n5349) );
  AND2_X1 U6848 ( .A1(n5350), .A2(n5349), .ZN(n9320) );
  NAND2_X1 U6849 ( .A1(n5542), .A2(n9320), .ZN(n5353) );
  NAND2_X1 U6850 ( .A1(n5523), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n5352) );
  NAND2_X1 U6851 ( .A1(n5543), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n5351) );
  NAND4_X1 U6852 ( .A1(n5354), .A2(n5353), .A3(n5352), .A4(n5351), .ZN(n9005)
         );
  INV_X1 U6853 ( .A(n9005), .ZN(n9298) );
  OR2_X1 U6854 ( .A1(n9408), .A2(n9298), .ZN(n8067) );
  NAND2_X1 U6855 ( .A1(n9408), .A2(n9298), .ZN(n8066) );
  NAND2_X1 U6856 ( .A1(n8067), .A2(n8066), .ZN(n9309) );
  XNOR2_X1 U6857 ( .A(n5356), .B(n5355), .ZN(n9733) );
  NAND2_X1 U6858 ( .A1(n9733), .A2(n4613), .ZN(n5360) );
  OR2_X1 U6859 ( .A1(n5357), .A2(n9439), .ZN(n5358) );
  XNOR2_X1 U6860 ( .A(n5358), .B(P1_IR_REG_14__SCAN_IN), .ZN(n9731) );
  AOI22_X1 U6861 ( .A1(n5535), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n5534), .B2(
        n9731), .ZN(n5359) );
  NAND2_X1 U6862 ( .A1(n4397), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n5366) );
  INV_X1 U6863 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n7597) );
  NAND2_X1 U6864 ( .A1(n5375), .A2(n7597), .ZN(n5361) );
  AND2_X1 U6865 ( .A1(n5362), .A2(n5361), .ZN(n8874) );
  NAND2_X1 U6866 ( .A1(n4391), .A2(n8874), .ZN(n5365) );
  NAND2_X1 U6867 ( .A1(n5523), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n5364) );
  NAND2_X1 U6868 ( .A1(n5543), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5363) );
  NAND4_X1 U6869 ( .A1(n5366), .A2(n5365), .A3(n5364), .A4(n5363), .ZN(n9006)
         );
  INV_X1 U6870 ( .A(n9006), .ZN(n9828) );
  OR2_X1 U6871 ( .A1(n9416), .A2(n9828), .ZN(n8064) );
  NAND2_X1 U6872 ( .A1(n9416), .A2(n9828), .ZN(n5657) );
  XNOR2_X1 U6873 ( .A(n5367), .B(n4963), .ZN(n7014) );
  NAND2_X1 U6874 ( .A1(n7014), .A2(n4613), .ZN(n5372) );
  OR2_X1 U6875 ( .A1(n5368), .A2(n9439), .ZN(n5531) );
  OAI21_X1 U6876 ( .B1(P1_IR_REG_11__SCAN_IN), .B2(P1_IR_REG_10__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5369) );
  NAND2_X1 U6877 ( .A1(n5531), .A2(n5369), .ZN(n5509) );
  OAI21_X1 U6878 ( .B1(n5509), .B2(P1_IR_REG_12__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5370) );
  XNOR2_X1 U6879 ( .A(n5370), .B(P1_IR_REG_13__SCAN_IN), .ZN(n7600) );
  AOI22_X1 U6880 ( .A1(n5535), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n5534), .B2(
        n7600), .ZN(n5371) );
  NAND2_X1 U6881 ( .A1(n5513), .A2(n5373), .ZN(n5374) );
  AND2_X1 U6882 ( .A1(n5375), .A2(n5374), .ZN(n9833) );
  NAND2_X1 U6883 ( .A1(n5542), .A2(n9833), .ZN(n5379) );
  NAND2_X1 U6884 ( .A1(n4397), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n5378) );
  NAND2_X1 U6885 ( .A1(n5523), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n5377) );
  NAND2_X1 U6886 ( .A1(n5543), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n5376) );
  NAND4_X1 U6887 ( .A1(n5379), .A2(n5378), .A3(n5377), .A4(n5376), .ZN(n9007)
         );
  INV_X1 U6888 ( .A(n9007), .ZN(n6549) );
  OR2_X1 U6889 ( .A1(n7979), .A2(n6549), .ZN(n5660) );
  NAND2_X1 U6890 ( .A1(n7979), .A2(n6549), .ZN(n7960) );
  NAND2_X1 U6891 ( .A1(n4391), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n5383) );
  NAND2_X1 U6892 ( .A1(n5452), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5382) );
  NAND2_X1 U6893 ( .A1(n5453), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n5380) );
  NAND4_X2 U6894 ( .A1(n5383), .A2(n5382), .A3(n5381), .A4(n5380), .ZN(n7361)
         );
  NAND2_X1 U6895 ( .A1(n6891), .A2(SI_0_), .ZN(n5385) );
  INV_X1 U6896 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5384) );
  NAND2_X1 U6897 ( .A1(n5385), .A2(n5384), .ZN(n5387) );
  AND2_X1 U6898 ( .A1(n5387), .A2(n5386), .ZN(n9736) );
  MUX2_X1 U6899 ( .A(P1_IR_REG_0__SCAN_IN), .B(n9736), .S(n5388), .Z(n7521) );
  INV_X1 U6900 ( .A(n7377), .ZN(n5389) );
  NAND2_X1 U6901 ( .A1(n7361), .A2(n7408), .ZN(n5754) );
  NAND2_X1 U6902 ( .A1(n5389), .A2(n5754), .ZN(n7120) );
  NAND2_X1 U6903 ( .A1(n5452), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n5391) );
  NAND2_X1 U6904 ( .A1(n5453), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5390) );
  NAND2_X1 U6905 ( .A1(n5391), .A2(n5390), .ZN(n5393) );
  INV_X1 U6906 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n5392) );
  NAND2_X1 U6907 ( .A1(n4397), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n5394) );
  NAND2_X1 U6908 ( .A1(n5420), .A2(n5419), .ZN(n5418) );
  NAND2_X1 U6909 ( .A1(n5418), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5398) );
  INV_X1 U6910 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n5397) );
  XNOR2_X1 U6911 ( .A(n5398), .B(n5397), .ZN(n6888) );
  XNOR2_X1 U6912 ( .A(n5400), .B(n5399), .ZN(n5949) );
  INV_X1 U6913 ( .A(n5949), .ZN(n6892) );
  OR2_X1 U6914 ( .A1(n5464), .A2(n4694), .ZN(n5401) );
  OAI211_X1 U6915 ( .C1(n7005), .C2(n6888), .A(n5402), .B(n5401), .ZN(n7566)
         );
  NAND2_X1 U6916 ( .A1(n9017), .A2(n10003), .ZN(n5620) );
  NAND2_X1 U6917 ( .A1(n5761), .A2(n5620), .ZN(n7556) );
  NAND2_X1 U6918 ( .A1(n4397), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5407) );
  INV_X1 U6919 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n5403) );
  XNOR2_X1 U6920 ( .A(n5403), .B(P1_REG3_REG_3__SCAN_IN), .ZN(n7429) );
  NAND2_X1 U6921 ( .A1(n5542), .A2(n7429), .ZN(n5406) );
  NAND2_X1 U6922 ( .A1(n5523), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n5405) );
  NAND2_X1 U6923 ( .A1(n5543), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5404) );
  OAI21_X1 U6924 ( .B1(P1_IR_REG_2__SCAN_IN), .B2(P1_IR_REG_3__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5408) );
  NAND2_X1 U6925 ( .A1(n5420), .A2(n5408), .ZN(n5409) );
  XNOR2_X1 U6926 ( .A(n5409), .B(P1_IR_REG_4__SCAN_IN), .ZN(n9884) );
  XNOR2_X1 U6927 ( .A(n5411), .B(n5410), .ZN(n5936) );
  INV_X1 U6928 ( .A(n5936), .ZN(n6895) );
  OR2_X1 U6929 ( .A1(n5463), .A2(n6895), .ZN(n5413) );
  INV_X1 U6930 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n9713) );
  OR2_X1 U6931 ( .A1(n5464), .A2(n9713), .ZN(n5412) );
  OAI211_X1 U6932 ( .C1(n9884), .C2(n7005), .A(n5413), .B(n5412), .ZN(n10009)
         );
  NAND2_X1 U6933 ( .A1(n7558), .A2(n10009), .ZN(n5629) );
  INV_X1 U6934 ( .A(n10009), .ZN(n7431) );
  NAND2_X1 U6935 ( .A1(n9016), .A2(n7431), .ZN(n5627) );
  NAND2_X1 U6936 ( .A1(n5629), .A2(n5627), .ZN(n7422) );
  NAND2_X1 U6937 ( .A1(n5542), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n5417) );
  NAND2_X1 U6938 ( .A1(n5452), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5416) );
  NAND2_X1 U6939 ( .A1(n5453), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5414) );
  XNOR2_X1 U6940 ( .A(n5421), .B(n5422), .ZN(n6000) );
  INV_X1 U6941 ( .A(n6000), .ZN(n6893) );
  NAND2_X1 U6942 ( .A1(n9018), .A2(n9997), .ZN(n5757) );
  NOR4_X1 U6943 ( .A1(n7120), .A2(n7556), .A3(n7422), .A4(n7511), .ZN(n5467)
         );
  NAND2_X1 U6944 ( .A1(n4397), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n5428) );
  INV_X1 U6945 ( .A(n5423), .ZN(n5441) );
  INV_X1 U6946 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n9566) );
  NAND2_X1 U6947 ( .A1(n5441), .A2(n9566), .ZN(n5424) );
  AND2_X1 U6948 ( .A1(n5494), .A2(n5424), .ZN(n7614) );
  NAND2_X1 U6949 ( .A1(n5542), .A2(n7614), .ZN(n5427) );
  NAND2_X1 U6950 ( .A1(n5523), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n5426) );
  NAND2_X1 U6951 ( .A1(n5543), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5425) );
  NAND4_X1 U6952 ( .A1(n5428), .A2(n5427), .A3(n5426), .A4(n5425), .ZN(n9014)
         );
  INV_X1 U6953 ( .A(n9014), .ZN(n7477) );
  NAND2_X1 U6954 ( .A1(n5429), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5430) );
  MUX2_X1 U6955 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5430), .S(
        P1_IR_REG_6__SCAN_IN), .Z(n5433) );
  INV_X1 U6956 ( .A(n5431), .ZN(n5432) );
  NAND2_X1 U6957 ( .A1(n5433), .A2(n5432), .ZN(n7031) );
  INV_X1 U6958 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6890) );
  OR2_X1 U6959 ( .A1(n5464), .A2(n6890), .ZN(n5436) );
  OAI211_X1 U6960 ( .C1(n7005), .C2(n7031), .A(n5437), .B(n5436), .ZN(n7615)
         );
  NAND2_X1 U6961 ( .A1(n7477), .A2(n7615), .ZN(n5632) );
  NAND2_X1 U6962 ( .A1(n4397), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5445) );
  INV_X1 U6963 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n5439) );
  NAND2_X1 U6964 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n5438) );
  NAND2_X1 U6965 ( .A1(n5439), .A2(n5438), .ZN(n5440) );
  AND2_X1 U6966 ( .A1(n5441), .A2(n5440), .ZN(n7533) );
  NAND2_X1 U6967 ( .A1(n5542), .A2(n7533), .ZN(n5444) );
  NAND2_X1 U6968 ( .A1(n5523), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n5443) );
  NAND2_X1 U6969 ( .A1(n5543), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n5442) );
  NAND4_X1 U6970 ( .A1(n5445), .A2(n5444), .A3(n5443), .A4(n5442), .ZN(n9015)
         );
  INV_X1 U6971 ( .A(n9015), .ZN(n7622) );
  NAND2_X1 U6972 ( .A1(n5446), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5447) );
  XNOR2_X1 U6973 ( .A(n5447), .B(n5118), .ZN(n7062) );
  OR2_X1 U6974 ( .A1(n5463), .A2(n6897), .ZN(n5451) );
  OR2_X1 U6975 ( .A1(n5464), .A2(n6889), .ZN(n5450) );
  OAI211_X1 U6976 ( .C1(n5388), .C2(n7062), .A(n5451), .B(n5450), .ZN(n7462)
         );
  NAND2_X1 U6977 ( .A1(n7622), .A2(n7462), .ZN(n5630) );
  INV_X1 U6978 ( .A(n7462), .ZN(n7538) );
  NAND2_X1 U6979 ( .A1(n9015), .A2(n7538), .ZN(n5631) );
  NAND2_X1 U6980 ( .A1(n5452), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n5456) );
  NAND2_X1 U6981 ( .A1(n4396), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n5455) );
  NAND2_X1 U6982 ( .A1(n5453), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5454) );
  AND3_X1 U6983 ( .A1(n5456), .A2(n5455), .A3(n5454), .ZN(n5458) );
  INV_X1 U6984 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n5460) );
  NAND2_X1 U6985 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5459) );
  XNOR2_X1 U6986 ( .A(n5460), .B(n5459), .ZN(n6885) );
  XNOR2_X1 U6987 ( .A(n5462), .B(n5461), .ZN(n5986) );
  INV_X1 U6988 ( .A(n5986), .ZN(n6894) );
  OR2_X1 U6989 ( .A1(n5463), .A2(n6894), .ZN(n5466) );
  NAND2_X1 U6990 ( .A1(n4589), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n5465) );
  OAI211_X1 U6991 ( .C1(n7005), .C2(n6885), .A(n5466), .B(n5465), .ZN(n5574)
         );
  INV_X1 U6992 ( .A(n5574), .ZN(n9991) );
  INV_X1 U6993 ( .A(n7363), .ZN(n5573) );
  NAND4_X1 U6994 ( .A1(n5467), .A2(n7620), .A3(n7618), .A4(n5573), .ZN(n5505)
         );
  NAND2_X1 U6995 ( .A1(n5487), .A2(n5468), .ZN(n5469) );
  AND2_X1 U6996 ( .A1(n5521), .A2(n5469), .ZN(n9968) );
  NAND2_X1 U6997 ( .A1(n5542), .A2(n9968), .ZN(n5473) );
  NAND2_X1 U6998 ( .A1(n4397), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n5472) );
  NAND2_X1 U6999 ( .A1(n5523), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n5471) );
  NAND2_X1 U7000 ( .A1(n5543), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5470) );
  NAND4_X1 U7001 ( .A1(n5473), .A2(n5472), .A3(n5471), .A4(n5470), .ZN(n9011)
         );
  INV_X1 U7002 ( .A(n9011), .ZN(n7645) );
  XNOR2_X1 U7003 ( .A(n5474), .B(n4964), .ZN(n6909) );
  NAND2_X1 U7004 ( .A1(n6909), .A2(n4613), .ZN(n5479) );
  INV_X1 U7005 ( .A(n5475), .ZN(n5476) );
  NAND2_X1 U7006 ( .A1(n5476), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5477) );
  XNOR2_X1 U7007 ( .A(n5477), .B(P1_IR_REG_9__SCAN_IN), .ZN(n7095) );
  AOI22_X1 U7008 ( .A1(n5535), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n5534), .B2(
        n7095), .ZN(n5478) );
  NAND2_X1 U7009 ( .A1(n5479), .A2(n5478), .ZN(n7647) );
  OR2_X1 U7010 ( .A1(n7645), .A2(n7647), .ZN(n5643) );
  NAND2_X1 U7011 ( .A1(n7647), .A2(n7645), .ZN(n7640) );
  NAND2_X1 U7012 ( .A1(n5643), .A2(n7640), .ZN(n9956) );
  XNOR2_X1 U7013 ( .A(n5481), .B(n5480), .ZN(n6905) );
  NAND2_X1 U7014 ( .A1(n6905), .A2(n4613), .ZN(n5485) );
  NAND2_X1 U7015 ( .A1(n5482), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5483) );
  XNOR2_X1 U7016 ( .A(n5483), .B(P1_IR_REG_8__SCAN_IN), .ZN(n7090) );
  AOI22_X1 U7017 ( .A1(n5535), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n5534), .B2(
        n7090), .ZN(n5484) );
  NAND2_X1 U7018 ( .A1(n5485), .A2(n5484), .ZN(n7633) );
  INV_X1 U7019 ( .A(n7633), .ZN(n7546) );
  INV_X1 U7020 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n7392) );
  NAND2_X1 U7021 ( .A1(n5496), .A2(n7392), .ZN(n5486) );
  AND2_X1 U7022 ( .A1(n5487), .A2(n5486), .ZN(n7543) );
  NAND2_X1 U7023 ( .A1(n4391), .A2(n7543), .ZN(n5492) );
  NAND2_X1 U7024 ( .A1(n4397), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5491) );
  NAND2_X1 U7025 ( .A1(n5523), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n5490) );
  NAND2_X1 U7026 ( .A1(n5543), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n5489) );
  NAND4_X1 U7027 ( .A1(n5492), .A2(n5491), .A3(n5490), .A4(n5489), .ZN(n9012)
         );
  NAND2_X1 U7028 ( .A1(n7546), .A2(n9012), .ZN(n9954) );
  INV_X1 U7029 ( .A(n9012), .ZN(n9958) );
  NAND2_X1 U7030 ( .A1(n9958), .A2(n7633), .ZN(n5641) );
  AND2_X1 U7031 ( .A1(n9954), .A2(n5641), .ZN(n7631) );
  INV_X1 U7032 ( .A(n7631), .ZN(n7500) );
  INV_X1 U7033 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n5493) );
  NAND2_X1 U7034 ( .A1(n5494), .A2(n5493), .ZN(n5495) );
  AND2_X1 U7035 ( .A1(n5496), .A2(n5495), .ZN(n7480) );
  NAND2_X1 U7036 ( .A1(n5542), .A2(n7480), .ZN(n5500) );
  NAND2_X1 U7037 ( .A1(n4397), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n5499) );
  NAND2_X1 U7038 ( .A1(n5523), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n5498) );
  NAND2_X1 U7039 ( .A1(n5543), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5497) );
  NAND4_X1 U7040 ( .A1(n5500), .A2(n5499), .A3(n5498), .A4(n5497), .ZN(n9013)
         );
  INV_X1 U7041 ( .A(n9013), .ZN(n7623) );
  INV_X1 U7042 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n9712) );
  OR2_X1 U7043 ( .A1(n5431), .A2(n9439), .ZN(n5503) );
  XNOR2_X1 U7044 ( .A(n5503), .B(P1_IR_REG_7__SCAN_IN), .ZN(n7092) );
  NAND2_X1 U7045 ( .A1(n5534), .A2(n7092), .ZN(n5504) );
  NAND2_X1 U7046 ( .A1(n7623), .A2(n7481), .ZN(n7498) );
  INV_X1 U7047 ( .A(n7481), .ZN(n10026) );
  NAND2_X1 U7048 ( .A1(n9013), .A2(n10026), .ZN(n5634) );
  NOR4_X1 U7049 ( .A1(n5505), .A2(n9956), .A3(n7500), .A4(n7495), .ZN(n5549)
         );
  XNOR2_X1 U7050 ( .A(n5507), .B(n5506), .ZN(n7011) );
  NAND2_X1 U7051 ( .A1(n7011), .A2(n4613), .ZN(n5511) );
  INV_X1 U7052 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n5508) );
  XNOR2_X1 U7053 ( .A(n5509), .B(n5508), .ZN(n7306) );
  AOI22_X1 U7054 ( .A1(n5535), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n5534), .B2(
        n7306), .ZN(n5510) );
  INV_X1 U7055 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n9653) );
  NAND2_X1 U7056 ( .A1(n5541), .A2(n9653), .ZN(n5512) );
  AND2_X1 U7057 ( .A1(n5513), .A2(n5512), .ZN(n7986) );
  NAND2_X1 U7058 ( .A1(n4391), .A2(n7986), .ZN(n5517) );
  NAND2_X1 U7059 ( .A1(n4397), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n5516) );
  NAND2_X1 U7060 ( .A1(n5523), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n5515) );
  NAND2_X1 U7061 ( .A1(n5543), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5514) );
  NAND4_X1 U7062 ( .A1(n5517), .A2(n5516), .A3(n5515), .A4(n5514), .ZN(n9008)
         );
  NAND2_X1 U7063 ( .A1(n7991), .A2(n9845), .ZN(n5646) );
  NAND2_X1 U7064 ( .A1(n5653), .A2(n5646), .ZN(n7879) );
  INV_X1 U7065 ( .A(n7879), .ZN(n7880) );
  XNOR2_X1 U7066 ( .A(n5518), .B(n4962), .ZN(n6915) );
  NAND2_X1 U7067 ( .A1(n6915), .A2(n4613), .ZN(n5520) );
  XNOR2_X1 U7068 ( .A(n5531), .B(P1_IR_REG_10__SCAN_IN), .ZN(n7219) );
  AOI22_X1 U7069 ( .A1(n5535), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n5534), .B2(
        n7219), .ZN(n5519) );
  NAND2_X1 U7070 ( .A1(n5521), .A2(n7102), .ZN(n5522) );
  AND2_X1 U7071 ( .A1(n5539), .A2(n5522), .ZN(n7648) );
  NAND2_X1 U7072 ( .A1(n4391), .A2(n7648), .ZN(n5527) );
  NAND2_X1 U7073 ( .A1(n4397), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n5526) );
  NAND2_X1 U7074 ( .A1(n5523), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n5525) );
  NAND2_X1 U7075 ( .A1(n5543), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5524) );
  NAND4_X1 U7076 ( .A1(n5527), .A2(n5526), .A3(n5525), .A4(n5524), .ZN(n9010)
         );
  NAND2_X1 U7077 ( .A1(n7868), .A2(n9961), .ZN(n5645) );
  NAND2_X1 U7078 ( .A1(n6919), .A2(n4613), .ZN(n5537) );
  INV_X1 U7079 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n5530) );
  NAND2_X1 U7080 ( .A1(n5531), .A2(n5530), .ZN(n5532) );
  NAND2_X1 U7081 ( .A1(n5532), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5533) );
  XNOR2_X1 U7082 ( .A(n5533), .B(P1_IR_REG_11__SCAN_IN), .ZN(n9930) );
  AOI22_X1 U7083 ( .A1(n5535), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n5534), .B2(
        n9930), .ZN(n5536) );
  NAND2_X1 U7084 ( .A1(n4397), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n5547) );
  INV_X1 U7085 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n5538) );
  NAND2_X1 U7086 ( .A1(n5539), .A2(n5538), .ZN(n5540) );
  AND2_X1 U7087 ( .A1(n5541), .A2(n5540), .ZN(n9847) );
  NAND2_X1 U7088 ( .A1(n5542), .A2(n9847), .ZN(n5546) );
  NAND2_X1 U7089 ( .A1(n5523), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n5545) );
  NAND2_X1 U7090 ( .A1(n5543), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5544) );
  NAND4_X1 U7091 ( .A1(n5547), .A2(n5546), .A3(n5545), .A4(n5544), .ZN(n9009)
         );
  NOR2_X1 U7092 ( .A1(n9849), .A2(n9009), .ZN(n7871) );
  NAND2_X1 U7093 ( .A1(n9849), .A2(n9009), .ZN(n7872) );
  INV_X1 U7094 ( .A(n7872), .ZN(n5548) );
  OR2_X1 U7095 ( .A1(n7871), .A2(n5548), .ZN(n9841) );
  AND4_X1 U7096 ( .A1(n5549), .A2(n7880), .A3(n7643), .A4(n9841), .ZN(n5550)
         );
  NAND3_X1 U7097 ( .A1(n7961), .A2(n9827), .A3(n5550), .ZN(n5551) );
  NOR4_X1 U7098 ( .A1(n9275), .A2(n9296), .A3(n9309), .A4(n5551), .ZN(n5552)
         );
  NAND4_X1 U7099 ( .A1(n9233), .A2(n9243), .A3(n9258), .A4(n5552), .ZN(n5553)
         );
  NOR4_X1 U7100 ( .A1(n9187), .A2(n9213), .A3(n9201), .A4(n5553), .ZN(n5554)
         );
  NAND4_X1 U7101 ( .A1(n8112), .A2(n9164), .A3(n9154), .A4(n5554), .ZN(n5555)
         );
  NOR4_X1 U7102 ( .A1(n8113), .A2(n9104), .A3(n9140), .A4(n5555), .ZN(n5557)
         );
  INV_X1 U7103 ( .A(n5722), .ZN(n9093) );
  NAND2_X1 U7104 ( .A1(n9095), .A2(n9093), .ZN(n5781) );
  INV_X1 U7105 ( .A(n9099), .ZN(n9330) );
  INV_X1 U7106 ( .A(n9001), .ZN(n5556) );
  NAND2_X1 U7107 ( .A1(n9330), .A2(n5556), .ZN(n5779) );
  NAND4_X1 U7108 ( .A1(n5777), .A2(n5557), .A3(n5781), .A4(n5779), .ZN(n5563)
         );
  INV_X1 U7109 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5749) );
  NAND2_X1 U7110 ( .A1(n5748), .A2(n5749), .ZN(n5559) );
  INV_X1 U7111 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5560) );
  AND2_X2 U7112 ( .A1(n5617), .A2(n5562), .ZN(n6433) );
  NAND2_X1 U7113 ( .A1(n5726), .A2(n5732), .ZN(n5568) );
  INV_X1 U7114 ( .A(n5568), .ZN(n5566) );
  INV_X1 U7115 ( .A(n5731), .ZN(n9103) );
  NAND2_X1 U7116 ( .A1(n9351), .A2(n9126), .ZN(n8085) );
  AND2_X1 U7117 ( .A1(n8086), .A2(n5730), .ZN(n5714) );
  OAI21_X1 U7118 ( .B1(n9103), .B2(n8085), .A(n5714), .ZN(n5565) );
  INV_X1 U7119 ( .A(n5733), .ZN(n5564) );
  AOI21_X1 U7120 ( .B1(n5566), .B2(n5565), .A(n5564), .ZN(n5571) );
  INV_X1 U7121 ( .A(n8084), .ZN(n5708) );
  OR2_X1 U7122 ( .A1(n9351), .A2(n9126), .ZN(n5567) );
  NAND2_X1 U7123 ( .A1(n5731), .A2(n5567), .ZN(n5715) );
  OR3_X1 U7124 ( .A1(n5568), .A2(n5708), .A3(n5715), .ZN(n5611) );
  AND2_X1 U7125 ( .A1(n5706), .A2(n5569), .ZN(n5698) );
  OR2_X1 U7126 ( .A1(n5611), .A2(n5698), .ZN(n5570) );
  AND2_X1 U7127 ( .A1(n5571), .A2(n5570), .ZN(n5773) );
  NAND2_X1 U7128 ( .A1(n9093), .A2(n9001), .ZN(n5572) );
  AND2_X1 U7129 ( .A1(n9330), .A2(n5572), .ZN(n5719) );
  INV_X1 U7130 ( .A(n5719), .ZN(n5734) );
  NAND2_X1 U7131 ( .A1(n5573), .A2(n7377), .ZN(n7376) );
  INV_X1 U7132 ( .A(n6440), .ZN(n7513) );
  NAND2_X1 U7133 ( .A1(n7513), .A2(n7522), .ZN(n5575) );
  INV_X1 U7134 ( .A(n7511), .ZN(n5576) );
  NAND2_X1 U7135 ( .A1(n5577), .A2(n5756), .ZN(n7555) );
  AND2_X1 U7136 ( .A1(n5627), .A2(n5620), .ZN(n5759) );
  INV_X1 U7137 ( .A(n5631), .ZN(n5578) );
  NAND2_X1 U7138 ( .A1(n5632), .A2(n5578), .ZN(n5579) );
  AND2_X1 U7139 ( .A1(n5579), .A2(n5624), .ZN(n7471) );
  NAND3_X1 U7140 ( .A1(n7555), .A2(n5759), .A3(n7471), .ZN(n5597) );
  AND2_X1 U7141 ( .A1(n5631), .A2(n5627), .ZN(n5622) );
  INV_X1 U7142 ( .A(n5622), .ZN(n5580) );
  AOI21_X1 U7143 ( .B1(n5629), .B2(n5761), .A(n5580), .ZN(n5581) );
  NAND2_X1 U7144 ( .A1(n5632), .A2(n5630), .ZN(n5764) );
  OAI21_X1 U7145 ( .B1(n5581), .B2(n5764), .A(n5624), .ZN(n5596) );
  AND2_X1 U7146 ( .A1(n8079), .A2(n8077), .ZN(n5688) );
  NAND2_X1 U7147 ( .A1(n5690), .A2(n8074), .ZN(n5582) );
  AND2_X1 U7148 ( .A1(n5688), .A2(n5582), .ZN(n5691) );
  INV_X1 U7149 ( .A(n5691), .ZN(n5605) );
  INV_X1 U7150 ( .A(n8075), .ZN(n9208) );
  NAND2_X1 U7151 ( .A1(n5677), .A2(n8070), .ZN(n5674) );
  INV_X1 U7152 ( .A(n5674), .ZN(n5584) );
  AND2_X1 U7153 ( .A1(n8073), .A2(n8072), .ZN(n5683) );
  INV_X1 U7154 ( .A(n5683), .ZN(n5583) );
  OR2_X1 U7155 ( .A1(n5584), .A2(n5583), .ZN(n5585) );
  AND4_X1 U7156 ( .A1(n9208), .A2(n5690), .A3(n5585), .A4(n5679), .ZN(n5586)
         );
  OAI21_X1 U7157 ( .B1(n5605), .B2(n5586), .A(n8078), .ZN(n5607) );
  AND2_X1 U7158 ( .A1(n9260), .A2(n8069), .ZN(n5587) );
  NAND2_X1 U7159 ( .A1(n8072), .A2(n5587), .ZN(n5602) );
  NAND2_X1 U7160 ( .A1(n8064), .A2(n5660), .ZN(n5658) );
  INV_X1 U7161 ( .A(n9009), .ZN(n7989) );
  NAND2_X1 U7162 ( .A1(n5646), .A2(n4438), .ZN(n5588) );
  AND2_X1 U7163 ( .A1(n5588), .A2(n5653), .ZN(n7958) );
  AND2_X1 U7164 ( .A1(n5643), .A2(n9954), .ZN(n7642) );
  AND2_X1 U7165 ( .A1(n7642), .A2(n5644), .ZN(n7875) );
  NAND2_X1 U7166 ( .A1(n9849), .A2(n7989), .ZN(n7878) );
  NAND2_X1 U7167 ( .A1(n5646), .A2(n7878), .ZN(n5654) );
  NAND2_X1 U7168 ( .A1(n5645), .A2(n7640), .ZN(n5637) );
  NAND2_X1 U7169 ( .A1(n5637), .A2(n5644), .ZN(n7876) );
  INV_X1 U7170 ( .A(n7876), .ZN(n5589) );
  OR3_X1 U7171 ( .A1(n7875), .A2(n5654), .A3(n5589), .ZN(n5590) );
  NAND2_X1 U7172 ( .A1(n7958), .A2(n5590), .ZN(n5591) );
  AND2_X1 U7173 ( .A1(n5591), .A2(n7960), .ZN(n5592) );
  OAI211_X1 U7174 ( .C1(n5658), .C2(n5592), .A(n8066), .B(n5657), .ZN(n5593)
         );
  AND3_X1 U7175 ( .A1(n5668), .A2(n8067), .A3(n5593), .ZN(n5594) );
  OR2_X1 U7176 ( .A1(n5602), .A2(n5594), .ZN(n5600) );
  NAND2_X1 U7177 ( .A1(n5600), .A2(n5634), .ZN(n5595) );
  OR2_X1 U7178 ( .A1(n5607), .A2(n5595), .ZN(n5765) );
  AOI21_X1 U7179 ( .B1(n5597), .B2(n5596), .A(n5765), .ZN(n5612) );
  AND2_X1 U7180 ( .A1(n5657), .A2(n7960), .ZN(n5662) );
  NAND3_X1 U7181 ( .A1(n7876), .A2(n5641), .A3(n7498), .ZN(n5598) );
  NOR2_X1 U7182 ( .A1(n5654), .A2(n5598), .ZN(n5599) );
  NAND3_X1 U7183 ( .A1(n8066), .A2(n5662), .A3(n5599), .ZN(n5601) );
  OAI21_X1 U7184 ( .B1(n5602), .B2(n5601), .A(n5600), .ZN(n5603) );
  NAND2_X1 U7185 ( .A1(n5603), .A2(n8073), .ZN(n5604) );
  NOR2_X1 U7186 ( .A1(n5605), .A2(n5604), .ZN(n5606) );
  OR2_X1 U7187 ( .A1(n5607), .A2(n5606), .ZN(n5609) );
  NAND2_X1 U7188 ( .A1(n5609), .A2(n5608), .ZN(n5769) );
  INV_X1 U7189 ( .A(n8082), .ZN(n5610) );
  NOR2_X1 U7190 ( .A1(n5611), .A2(n5610), .ZN(n5776) );
  OAI211_X1 U7191 ( .C1(n5612), .C2(n5769), .A(n5776), .B(n8083), .ZN(n5613)
         );
  AND3_X1 U7192 ( .A1(n5773), .A2(n5734), .A3(n5613), .ZN(n5615) );
  NAND2_X1 U7193 ( .A1(n4965), .A2(n9093), .ZN(n5725) );
  NAND2_X1 U7194 ( .A1(n9091), .A2(n5725), .ZN(n5718) );
  INV_X1 U7195 ( .A(n5718), .ZN(n5614) );
  OAI211_X1 U7196 ( .C1(n5615), .C2(n5614), .A(n6433), .B(n5781), .ZN(n5616)
         );
  NAND2_X1 U7197 ( .A1(n5741), .A2(n5616), .ZN(n5745) );
  INV_X1 U7198 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5618) );
  XNOR2_X2 U7199 ( .A(n5619), .B(n5618), .ZN(n6434) );
  NAND2_X1 U7200 ( .A1(n6434), .A2(n9250), .ZN(n7399) );
  AND2_X1 U7201 ( .A1(n5726), .A2(n7399), .ZN(n5721) );
  NAND2_X1 U7202 ( .A1(n7555), .A2(n5620), .ZN(n5621) );
  NAND2_X1 U7203 ( .A1(n5621), .A2(n5761), .ZN(n5628) );
  INV_X1 U7204 ( .A(n5629), .ZN(n5763) );
  OAI21_X1 U7205 ( .B1(n5628), .B2(n5763), .A(n5622), .ZN(n5623) );
  NAND3_X1 U7206 ( .A1(n5623), .A2(n7620), .A3(n5630), .ZN(n5625) );
  NAND3_X1 U7207 ( .A1(n5625), .A2(n5634), .A3(n5624), .ZN(n5626) );
  NAND2_X1 U7208 ( .A1(n5626), .A2(n7498), .ZN(n5636) );
  NAND2_X1 U7209 ( .A1(n5628), .A2(n5627), .ZN(n7470) );
  NAND2_X1 U7210 ( .A1(n7470), .A2(n5629), .ZN(n7619) );
  INV_X1 U7211 ( .A(n5630), .ZN(n7617) );
  OAI211_X1 U7212 ( .C1(n7619), .C2(n7617), .A(n7620), .B(n5631), .ZN(n5633)
         );
  NAND3_X1 U7213 ( .A1(n5633), .A2(n5632), .A3(n7498), .ZN(n5635) );
  INV_X1 U7214 ( .A(n5641), .ZN(n7639) );
  INV_X1 U7215 ( .A(n5637), .ZN(n5639) );
  NAND2_X1 U7216 ( .A1(n5653), .A2(n5644), .ZN(n5638) );
  AOI21_X1 U7217 ( .B1(n5640), .B2(n5639), .A(n5638), .ZN(n5651) );
  INV_X1 U7218 ( .A(n9954), .ZN(n5642) );
  AND2_X1 U7219 ( .A1(n5644), .A2(n5643), .ZN(n5648) );
  NAND2_X1 U7220 ( .A1(n5646), .A2(n5645), .ZN(n5647) );
  AOI21_X1 U7221 ( .B1(n5649), .B2(n5648), .A(n5647), .ZN(n5650) );
  MUX2_X1 U7222 ( .A(n5651), .B(n5650), .S(n7399), .Z(n5652) );
  NAND2_X1 U7223 ( .A1(n5652), .A2(n9841), .ZN(n5661) );
  INV_X1 U7224 ( .A(n5662), .ZN(n5656) );
  AND2_X1 U7225 ( .A1(n5654), .A2(n5653), .ZN(n5655) );
  NOR2_X1 U7226 ( .A1(n5656), .A2(n5655), .ZN(n5659) );
  AOI22_X1 U7227 ( .A1(n5661), .A2(n5659), .B1(n5658), .B2(n5657), .ZN(n5664)
         );
  NAND3_X1 U7228 ( .A1(n5661), .A2(n7958), .A3(n5660), .ZN(n5663) );
  INV_X1 U7229 ( .A(n9309), .ZN(n9312) );
  INV_X1 U7230 ( .A(n8066), .ZN(n5666) );
  INV_X1 U7231 ( .A(n8067), .ZN(n5665) );
  MUX2_X1 U7232 ( .A(n5666), .B(n5665), .S(n7399), .Z(n5667) );
  NOR2_X1 U7233 ( .A1(n9296), .A2(n5667), .ZN(n5671) );
  INV_X1 U7234 ( .A(n9275), .ZN(n9282) );
  MUX2_X1 U7235 ( .A(n5668), .B(n8069), .S(n7399), .Z(n5669) );
  NAND2_X1 U7236 ( .A1(n9282), .A2(n5669), .ZN(n5670) );
  AOI21_X1 U7237 ( .B1(n5672), .B2(n5671), .A(n5670), .ZN(n5676) );
  NAND2_X1 U7238 ( .A1(n8072), .A2(n9260), .ZN(n5673) );
  MUX2_X1 U7239 ( .A(n5674), .B(n5673), .S(n4602), .Z(n5675) );
  NOR2_X1 U7240 ( .A1(n8074), .A2(n7399), .ZN(n5678) );
  INV_X1 U7241 ( .A(n5679), .ZN(n5680) );
  OR3_X1 U7242 ( .A1(n8075), .A2(n5680), .A3(n4602), .ZN(n5681) );
  NAND3_X1 U7243 ( .A1(n5684), .A2(n5683), .A3(n5682), .ZN(n5685) );
  NAND2_X1 U7244 ( .A1(n5686), .A2(n5685), .ZN(n5693) );
  NAND3_X1 U7245 ( .A1(n5693), .A2(n5690), .A3(n9208), .ZN(n5689) );
  INV_X1 U7246 ( .A(n8078), .ZN(n5687) );
  AOI21_X1 U7247 ( .B1(n5689), .B2(n5688), .A(n5687), .ZN(n5694) );
  INV_X1 U7248 ( .A(n5690), .ZN(n5692) );
  MUX2_X1 U7249 ( .A(n9366), .B(n9203), .S(n4602), .Z(n5696) );
  NAND2_X1 U7250 ( .A1(n9366), .A2(n9203), .ZN(n8107) );
  NAND2_X1 U7251 ( .A1(n5696), .A2(n8107), .ZN(n5695) );
  INV_X1 U7252 ( .A(n5696), .ZN(n5699) );
  NAND3_X1 U7253 ( .A1(n9164), .A2(n5699), .A3(n9366), .ZN(n5697) );
  NAND2_X1 U7254 ( .A1(n5698), .A2(n5697), .ZN(n5702) );
  NAND3_X1 U7255 ( .A1(n9164), .A2(n5699), .A3(n9203), .ZN(n5700) );
  NAND3_X1 U7256 ( .A1(n5700), .A2(n8084), .A3(n8083), .ZN(n5701) );
  MUX2_X1 U7257 ( .A(n5702), .B(n5701), .S(n7399), .Z(n5703) );
  INV_X1 U7258 ( .A(n5703), .ZN(n5704) );
  NAND2_X1 U7259 ( .A1(n5705), .A2(n5704), .ZN(n5711) );
  INV_X1 U7260 ( .A(n5706), .ZN(n5707) );
  MUX2_X1 U7261 ( .A(n5708), .B(n5707), .S(n7399), .Z(n5709) );
  NOR2_X1 U7262 ( .A1(n9140), .A2(n5709), .ZN(n5710) );
  NAND2_X1 U7263 ( .A1(n5711), .A2(n5710), .ZN(n5713) );
  OR2_X1 U7264 ( .A1(n8085), .A2(n7399), .ZN(n5712) );
  NAND2_X1 U7265 ( .A1(n5713), .A2(n5712), .ZN(n5729) );
  OAI21_X1 U7266 ( .B1(n5729), .B2(n5715), .A(n5714), .ZN(n5716) );
  NAND4_X1 U7267 ( .A1(n5718), .A2(n5721), .A3(n5732), .A4(n5716), .ZN(n5717)
         );
  OAI21_X1 U7268 ( .B1(n5718), .B2(n7399), .A(n5717), .ZN(n5740) );
  NAND3_X1 U7269 ( .A1(n5720), .A2(n5719), .A3(n7399), .ZN(n5738) );
  NAND2_X1 U7270 ( .A1(n5721), .A2(n8113), .ZN(n5723) );
  NAND2_X1 U7271 ( .A1(n5723), .A2(n5722), .ZN(n5724) );
  NAND2_X1 U7272 ( .A1(n9095), .A2(n5724), .ZN(n5737) );
  NAND2_X1 U7273 ( .A1(n5725), .A2(n7399), .ZN(n5728) );
  MUX2_X1 U7274 ( .A(n5733), .B(n5726), .S(n7399), .Z(n5727) );
  NAND4_X1 U7275 ( .A1(n5728), .A2(n5727), .A3(n5734), .A4(n8113), .ZN(n5736)
         );
  NAND2_X1 U7276 ( .A1(n5732), .A2(n5731), .ZN(n8087) );
  NAND4_X1 U7277 ( .A1(n5738), .A2(n5737), .A3(n5736), .A4(n5735), .ZN(n5739)
         );
  INV_X1 U7278 ( .A(n7118), .ZN(n5743) );
  INV_X1 U7279 ( .A(n5741), .ZN(n5742) );
  AOI21_X1 U7280 ( .B1(n5746), .B2(n5743), .A(n5742), .ZN(n5744) );
  MUX2_X1 U7281 ( .A(n5745), .B(n5744), .S(n9250), .Z(n5752) );
  INV_X1 U7282 ( .A(n5746), .ZN(n5747) );
  NAND4_X1 U7283 ( .A1(n5747), .A2(n6433), .A3(n6434), .A4(n5781), .ZN(n5750)
         );
  INV_X1 U7284 ( .A(n7494), .ZN(n7398) );
  NAND2_X1 U7285 ( .A1(n5752), .A2(n5751), .ZN(n5793) );
  NAND2_X1 U7286 ( .A1(n6440), .A2(n9991), .ZN(n5753) );
  NAND3_X1 U7287 ( .A1(n5754), .A2(n5753), .A3(n6433), .ZN(n5755) );
  NAND2_X1 U7288 ( .A1(n5756), .A2(n5755), .ZN(n5758) );
  INV_X1 U7289 ( .A(n5759), .ZN(n5760) );
  AOI21_X1 U7290 ( .B1(n5762), .B2(n5761), .A(n5760), .ZN(n5768) );
  NOR2_X1 U7291 ( .A1(n5764), .A2(n5763), .ZN(n7469) );
  INV_X1 U7292 ( .A(n7469), .ZN(n5767) );
  INV_X1 U7293 ( .A(n5765), .ZN(n5766) );
  OAI211_X1 U7294 ( .C1(n5768), .C2(n5767), .A(n5766), .B(n7471), .ZN(n5772)
         );
  INV_X1 U7295 ( .A(n5769), .ZN(n5771) );
  INV_X1 U7296 ( .A(n8083), .ZN(n5770) );
  AOI21_X1 U7297 ( .B1(n5772), .B2(n5771), .A(n5770), .ZN(n5775) );
  INV_X1 U7298 ( .A(n5773), .ZN(n5774) );
  AOI21_X1 U7299 ( .B1(n5776), .B2(n5775), .A(n5774), .ZN(n5780) );
  INV_X1 U7300 ( .A(n5777), .ZN(n5778) );
  INV_X1 U7301 ( .A(n5781), .ZN(n5782) );
  NOR2_X1 U7302 ( .A1(n5783), .A2(n5782), .ZN(n5784) );
  XNOR2_X1 U7303 ( .A(n5784), .B(n9086), .ZN(n5785) );
  NAND2_X1 U7304 ( .A1(n5785), .A2(n7494), .ZN(n5791) );
  INV_X1 U7305 ( .A(n5786), .ZN(n5787) );
  NAND2_X1 U7306 ( .A1(n5787), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5788) );
  MUX2_X1 U7307 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5788), .S(
        P1_IR_REG_23__SCAN_IN), .Z(n5789) );
  NAND2_X1 U7308 ( .A1(n5789), .A2(n4415), .ZN(n6835) );
  INV_X1 U7309 ( .A(n6835), .ZN(n6715) );
  NAND2_X1 U7310 ( .A1(n6715), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7730) );
  INV_X1 U7311 ( .A(n7730), .ZN(n5790) );
  NAND2_X1 U7312 ( .A1(n5793), .A2(n5792), .ZN(n5807) );
  INV_X1 U7313 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5798) );
  NAND2_X1 U7314 ( .A1(n5801), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5795) );
  INV_X1 U7315 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n5794) );
  XNOR2_X1 U7316 ( .A(n5795), .B(n5794), .ZN(n8044) );
  NAND2_X1 U7317 ( .A1(n4415), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5797) );
  XNOR2_X1 U7318 ( .A(n5797), .B(n5796), .ZN(n7941) );
  OR2_X1 U7319 ( .A1(n5799), .A2(n5798), .ZN(n5800) );
  NAND2_X1 U7320 ( .A1(n5801), .A2(n5800), .ZN(n8013) );
  OR3_X2 U7321 ( .A1(n8044), .A2(n7941), .A3(n8013), .ZN(n6834) );
  AND2_X1 U7322 ( .A1(n6834), .A2(n6835), .ZN(n5802) );
  NOR2_X1 U7323 ( .A1(n4394), .A2(P1_U3084), .ZN(n8056) );
  NAND3_X1 U7324 ( .A1(n7042), .A2(n9287), .A3(n8056), .ZN(n5805) );
  OAI211_X1 U7325 ( .C1(n6437), .C2(n7730), .A(n5805), .B(P1_B_REG_SCAN_IN), 
        .ZN(n5806) );
  NAND2_X1 U7326 ( .A1(n5807), .A2(n5806), .ZN(P1_U3240) );
  NOR2_X1 U7327 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n5815) );
  NOR2_X1 U7328 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_13__SCAN_IN), .ZN(
        n5814) );
  NAND4_X1 U7329 ( .A1(n5815), .A2(n5814), .A3(n5813), .A4(n5812), .ZN(n5818)
         );
  INV_X1 U7330 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n5816) );
  NAND4_X1 U7331 ( .A1(n6320), .A2(n5869), .A3(n6115), .A4(n5816), .ZN(n5817)
         );
  INV_X1 U7332 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n5821) );
  NAND4_X1 U7333 ( .A1(n5822), .A2(n6411), .A3(n6422), .A4(n5821), .ZN(n5824)
         );
  NAND2_X1 U7334 ( .A1(n6418), .A2(n6425), .ZN(n5823) );
  NAND2_X1 U7335 ( .A1(n5827), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5828) );
  INV_X1 U7336 ( .A(n6001), .ZN(n5832) );
  NAND2_X1 U7337 ( .A1(n8852), .A2(n6245), .ZN(n5834) );
  NAND2_X1 U7338 ( .A1(n6234), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n5833) );
  INV_X1 U7339 ( .A(n6030), .ZN(n5836) );
  AND2_X1 U7340 ( .A1(P2_REG3_REG_7__SCAN_IN), .A2(P2_REG3_REG_6__SCAN_IN), 
        .ZN(n5835) );
  NAND2_X1 U7341 ( .A1(n5836), .A2(n5835), .ZN(n6031) );
  INV_X1 U7342 ( .A(n6031), .ZN(n5837) );
  NAND2_X1 U7343 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_REG3_REG_9__SCAN_IN), 
        .ZN(n5838) );
  INV_X1 U7344 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n6090) );
  INV_X1 U7345 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n6121) );
  INV_X1 U7346 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n6138) );
  AND2_X1 U7347 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(P2_REG3_REG_17__SCAN_IN), 
        .ZN(n5841) );
  INV_X1 U7348 ( .A(n6175), .ZN(n5843) );
  NAND2_X1 U7349 ( .A1(n5843), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n6190) );
  INV_X1 U7350 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n6189) );
  INV_X1 U7351 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n8231) );
  INV_X1 U7352 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n8189) );
  INV_X1 U7353 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n8267) );
  INV_X1 U7354 ( .A(n6238), .ZN(n5846) );
  NAND2_X1 U7355 ( .A1(n5846), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n6249) );
  INV_X1 U7356 ( .A(n6249), .ZN(n5847) );
  NAND2_X1 U7357 ( .A1(n5847), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n6273) );
  NAND2_X1 U7358 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(P2_REG3_REG_28__SCAN_IN), 
        .ZN(n5848) );
  OR2_X1 U7359 ( .A1(n6273), .A2(n5848), .ZN(n8509) );
  INV_X1 U7360 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5851) );
  INV_X1 U7361 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n5852) );
  INV_X1 U7362 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n8510) );
  INV_X1 U7363 ( .A(n5855), .ZN(n5857) );
  NAND2_X1 U7364 ( .A1(n6304), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n5859) );
  NAND2_X1 U7365 ( .A1(n6294), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n5858) );
  OAI211_X1 U7366 ( .C1(n8510), .C2(n6305), .A(n5859), .B(n5858), .ZN(n5860)
         );
  INV_X1 U7367 ( .A(n5860), .ZN(n5861) );
  OAI21_X1 U7368 ( .B1(n8509), .B2(n6251), .A(n5861), .ZN(n8338) );
  INV_X1 U7369 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5863) );
  NAND2_X1 U7370 ( .A1(n5899), .A2(n5863), .ZN(n6050) );
  INV_X1 U7371 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n6112) );
  INV_X1 U7372 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n5866) );
  AND3_X1 U7373 ( .A1(n6115), .A2(n6112), .A3(n5866), .ZN(n5867) );
  INV_X1 U7374 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n5868) );
  NAND2_X1 U7375 ( .A1(n6172), .A2(n5869), .ZN(n5870) );
  INV_X1 U7376 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n6318) );
  XNOR2_X1 U7377 ( .A(n6408), .B(P2_IR_REG_22__SCAN_IN), .ZN(n6429) );
  NAND2_X1 U7378 ( .A1(n5871), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5872) );
  OR2_X1 U7379 ( .A1(n6429), .A2(n7552), .ZN(n5873) );
  NAND2_X1 U7380 ( .A1(n7938), .A2(n6245), .ZN(n5875) );
  NAND2_X1 U7381 ( .A1(n6234), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n5874) );
  NAND2_X1 U7382 ( .A1(n5882), .A2(n8267), .ZN(n5876) );
  NAND2_X1 U7383 ( .A1(n6238), .A2(n5876), .ZN(n8587) );
  AOI22_X1 U7384 ( .A1(n6304), .A2(P2_REG1_REG_24__SCAN_IN), .B1(n6294), .B2(
        P2_REG0_REG_24__SCAN_IN), .ZN(n5878) );
  NAND2_X1 U7385 ( .A1(n5890), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n5877) );
  OAI211_X1 U7386 ( .C1(n8587), .C2(n6251), .A(n5878), .B(n5877), .ZN(n8599)
         );
  INV_X1 U7387 ( .A(n8599), .ZN(n8263) );
  NAND2_X1 U7388 ( .A1(n7729), .A2(n6245), .ZN(n5880) );
  NAND2_X1 U7389 ( .A1(n6234), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n5879) );
  NAND2_X1 U7390 ( .A1(n5889), .A2(n8189), .ZN(n5881) );
  NAND2_X1 U7391 ( .A1(n5882), .A2(n5881), .ZN(n8604) );
  AOI22_X1 U7392 ( .A1(n6304), .A2(P2_REG1_REG_23__SCAN_IN), .B1(n6294), .B2(
        P2_REG0_REG_23__SCAN_IN), .ZN(n5884) );
  NAND2_X1 U7393 ( .A1(n5890), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n5883) );
  OAI211_X1 U7394 ( .C1(n8604), .C2(n6251), .A(n5884), .B(n5883), .ZN(n8490)
         );
  NAND2_X1 U7395 ( .A1(n8607), .A2(n8490), .ZN(n6225) );
  AND2_X1 U7396 ( .A1(n6389), .A2(n6225), .ZN(n6233) );
  NAND2_X1 U7397 ( .A1(n7661), .A2(n6245), .ZN(n5886) );
  NAND2_X1 U7398 ( .A1(n6234), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n5885) );
  INV_X1 U7399 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n5887) );
  NAND2_X1 U7400 ( .A1(n6212), .A2(n5887), .ZN(n5888) );
  NAND2_X1 U7401 ( .A1(n5889), .A2(n5888), .ZN(n8617) );
  OR2_X1 U7402 ( .A1(n8617), .A2(n6251), .ZN(n5894) );
  NAND2_X1 U7403 ( .A1(n6304), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n5893) );
  NAND2_X1 U7404 ( .A1(n6294), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n5892) );
  NAND2_X1 U7405 ( .A1(n5890), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n5891) );
  NAND2_X1 U7406 ( .A1(n8795), .A2(n8230), .ZN(n6327) );
  INV_X1 U7407 ( .A(n6327), .ZN(n6224) );
  NAND2_X1 U7408 ( .A1(n6294), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5898) );
  INV_X1 U7409 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n7018) );
  OR2_X1 U7410 ( .A1(n5931), .A2(n7018), .ZN(n5897) );
  INV_X1 U7411 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n6054) );
  XNOR2_X1 U7412 ( .A(n6055), .B(n6054), .ZN(n7824) );
  OR2_X1 U7413 ( .A1(n6251), .A2(n7824), .ZN(n5896) );
  INV_X1 U7414 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n7711) );
  OR2_X1 U7415 ( .A1(n6305), .A2(n7711), .ZN(n5895) );
  NAND2_X1 U7416 ( .A1(n6909), .A2(n6245), .ZN(n5902) );
  OR2_X1 U7417 ( .A1(n5899), .A2(n6416), .ZN(n5900) );
  XNOR2_X1 U7418 ( .A(n5900), .B(P2_IR_REG_9__SCAN_IN), .ZN(n7141) );
  AOI22_X1 U7419 ( .A1(n6234), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6186), .B2(
        n7141), .ZN(n5901) );
  NAND2_X1 U7420 ( .A1(n5902), .A2(n5901), .ZN(n7805) );
  OR2_X1 U7421 ( .A1(n7834), .A2(n7805), .ZN(n6340) );
  NAND2_X1 U7422 ( .A1(n6304), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5908) );
  INV_X1 U7423 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n5903) );
  OR2_X1 U7424 ( .A1(n6307), .A2(n5903), .ZN(n5907) );
  INV_X1 U7425 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n9686) );
  NAND2_X1 U7426 ( .A1(n6031), .A2(n9686), .ZN(n5904) );
  NAND2_X1 U7427 ( .A1(n6055), .A2(n5904), .ZN(n7689) );
  OR2_X1 U7428 ( .A1(n6251), .A2(n7689), .ZN(n5906) );
  INV_X1 U7429 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7690) );
  OR2_X1 U7430 ( .A1(n6305), .A2(n7690), .ZN(n5905) );
  NAND4_X1 U7431 ( .A1(n5908), .A2(n5907), .A3(n5906), .A4(n5905), .ZN(n8347)
         );
  NAND2_X1 U7432 ( .A1(n6905), .A2(n6245), .ZN(n5913) );
  INV_X1 U7433 ( .A(n5909), .ZN(n6037) );
  OR2_X1 U7434 ( .A1(n6037), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n5910) );
  NAND2_X1 U7435 ( .A1(n5910), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5911) );
  XNOR2_X1 U7436 ( .A(n5911), .B(P2_IR_REG_8__SCAN_IN), .ZN(n7022) );
  AOI22_X1 U7437 ( .A1(n6234), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n6186), .B2(
        n7022), .ZN(n5912) );
  NAND2_X1 U7438 ( .A1(n8347), .A2(n10165), .ZN(n6044) );
  AND2_X1 U7439 ( .A1(n6340), .A2(n6044), .ZN(n6048) );
  NAND2_X1 U7440 ( .A1(n6304), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n5918) );
  INV_X1 U7441 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n5914) );
  OR2_X1 U7442 ( .A1(n6307), .A2(n5914), .ZN(n5917) );
  OAI21_X1 U7443 ( .B1(n5926), .B2(P2_REG3_REG_5__SCAN_IN), .A(n6030), .ZN(
        n7782) );
  OR2_X1 U7444 ( .A1(n6251), .A2(n7782), .ZN(n5916) );
  INV_X1 U7445 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n7780) );
  OR2_X1 U7446 ( .A1(n6305), .A2(n7780), .ZN(n5915) );
  NAND4_X1 U7447 ( .A1(n5918), .A2(n5917), .A3(n5916), .A4(n5915), .ZN(n8350)
         );
  NAND2_X1 U7448 ( .A1(n6234), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n5925) );
  NOR2_X1 U7449 ( .A1(n5919), .A2(n6416), .ZN(n5920) );
  MUX2_X1 U7450 ( .A(n6416), .B(n5920), .S(P2_IR_REG_5__SCAN_IN), .Z(n5923) );
  OR2_X1 U7451 ( .A1(n5923), .A2(n5922), .ZN(n6958) );
  INV_X1 U7452 ( .A(n6958), .ZN(n8358) );
  NAND2_X1 U7453 ( .A1(n6186), .A2(n8358), .ZN(n5924) );
  NAND2_X1 U7454 ( .A1(n6294), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n5935) );
  INV_X1 U7455 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n6949) );
  OR2_X1 U7456 ( .A1(n5992), .A2(n6949), .ZN(n5934) );
  INV_X1 U7457 ( .A(n5926), .ZN(n5930) );
  INV_X1 U7458 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n5928) );
  INV_X1 U7459 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n5927) );
  NAND2_X1 U7460 ( .A1(n5928), .A2(n5927), .ZN(n5929) );
  NAND2_X1 U7461 ( .A1(n5930), .A2(n5929), .ZN(n10097) );
  OR2_X1 U7462 ( .A1(n6251), .A2(n10097), .ZN(n5933) );
  INV_X1 U7463 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n6934) );
  OR2_X1 U7464 ( .A1(n5931), .A2(n6934), .ZN(n5932) );
  NAND2_X1 U7465 ( .A1(n6245), .A2(n5936), .ZN(n5941) );
  NAND2_X1 U7466 ( .A1(n6234), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n5940) );
  NAND2_X1 U7467 ( .A1(n5937), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5938) );
  XNOR2_X1 U7468 ( .A(n5938), .B(P2_IR_REG_4__SCAN_IN), .ZN(n6957) );
  NAND2_X1 U7469 ( .A1(n6186), .A2(n6957), .ZN(n5939) );
  NAND2_X1 U7470 ( .A1(n6364), .A2(n6332), .ZN(n5943) );
  NAND2_X1 U7471 ( .A1(n8350), .A2(n6740), .ZN(n6333) );
  INV_X1 U7472 ( .A(n6363), .ZN(n5942) );
  INV_X1 U7473 ( .A(n6023), .ZN(n5966) );
  NAND2_X1 U7474 ( .A1(n5991), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5948) );
  INV_X1 U7475 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n5944) );
  OR2_X1 U7476 ( .A1(n6307), .A2(n5944), .ZN(n5947) );
  OR2_X1 U7477 ( .A1(n6202), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n5946) );
  INV_X1 U7478 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n6951) );
  OR2_X1 U7479 ( .A1(n5992), .A2(n6951), .ZN(n5945) );
  NAND2_X1 U7480 ( .A1(n5999), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n5954) );
  NAND2_X1 U7481 ( .A1(n6001), .A2(n5949), .ZN(n5953) );
  NAND2_X1 U7482 ( .A1(n5950), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5951) );
  XNOR2_X1 U7483 ( .A(n5951), .B(P2_IR_REG_3__SCAN_IN), .ZN(n6950) );
  NAND2_X1 U7484 ( .A1(n6186), .A2(n6950), .ZN(n5952) );
  NAND2_X1 U7485 ( .A1(n6360), .A2(n6332), .ZN(n5965) );
  INV_X1 U7486 ( .A(n6364), .ZN(n7737) );
  NAND2_X1 U7487 ( .A1(n6294), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5959) );
  INV_X1 U7488 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n5955) );
  OR2_X1 U7489 ( .A1(n5931), .A2(n5955), .ZN(n5958) );
  INV_X1 U7490 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n6029) );
  XNOR2_X1 U7491 ( .A(n6030), .B(n6029), .ZN(n8305) );
  OR2_X1 U7492 ( .A1(n6251), .A2(n8305), .ZN(n5957) );
  INV_X1 U7493 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n6948) );
  OR2_X1 U7494 ( .A1(n6305), .A2(n6948), .ZN(n5956) );
  INV_X1 U7495 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n9581) );
  NOR2_X1 U7496 ( .A1(n5922), .A2(n6416), .ZN(n5961) );
  MUX2_X1 U7497 ( .A(n6416), .B(n5961), .S(P2_IR_REG_6__SCAN_IN), .Z(n5962) );
  INV_X1 U7498 ( .A(n6959), .ZN(n8371) );
  NAND2_X1 U7499 ( .A1(n6186), .A2(n8371), .ZN(n5963) );
  NOR2_X1 U7500 ( .A1(n8349), .A2(n10151), .ZN(n10068) );
  AOI211_X1 U7501 ( .C1(n5966), .C2(n5965), .A(n7737), .B(n10068), .ZN(n6018)
         );
  NAND2_X1 U7502 ( .A1(n8352), .A2(n10141), .ZN(n6020) );
  NOR2_X1 U7503 ( .A1(n6023), .A2(n7750), .ZN(n6016) );
  NAND2_X1 U7504 ( .A1(n5991), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5972) );
  INV_X1 U7505 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n5967) );
  INV_X1 U7506 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n7790) );
  INV_X1 U7507 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n5968) );
  NAND2_X1 U7508 ( .A1(n5831), .A2(SI_0_), .ZN(n5974) );
  INV_X1 U7509 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5973) );
  NAND2_X1 U7510 ( .A1(n5974), .A2(n5973), .ZN(n5976) );
  AND2_X1 U7511 ( .A1(n5976), .A2(n5975), .ZN(n8860) );
  INV_X1 U7512 ( .A(n7792), .ZN(n10122) );
  NAND2_X1 U7513 ( .A1(n5990), .A2(n10122), .ZN(n6331) );
  AND2_X1 U7514 ( .A1(n6331), .A2(n6819), .ZN(n6009) );
  NAND2_X1 U7515 ( .A1(n5991), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5981) );
  INV_X1 U7516 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n5977) );
  INV_X1 U7517 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n7770) );
  INV_X1 U7518 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n6953) );
  NAND2_X1 U7519 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5982) );
  MUX2_X1 U7520 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5982), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n5985) );
  INV_X1 U7521 ( .A(n5983), .ZN(n5984) );
  NAND2_X1 U7522 ( .A1(n5985), .A2(n5984), .ZN(n6954) );
  NAND2_X1 U7523 ( .A1(n6001), .A2(n5986), .ZN(n5988) );
  NAND2_X1 U7524 ( .A1(n5999), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n5987) );
  NAND2_X1 U7525 ( .A1(n6334), .A2(n7772), .ZN(n6359) );
  NAND2_X1 U7526 ( .A1(n5991), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5998) );
  INV_X1 U7527 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n6952) );
  OR2_X1 U7528 ( .A1(n5992), .A2(n6952), .ZN(n5997) );
  INV_X1 U7529 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n7258) );
  OR2_X1 U7530 ( .A1(n6202), .A2(n7258), .ZN(n5996) );
  INV_X1 U7531 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n5993) );
  OR2_X1 U7532 ( .A1(n5994), .A2(n5993), .ZN(n5995) );
  NAND2_X1 U7533 ( .A1(n5999), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n6008) );
  NAND2_X1 U7534 ( .A1(n6001), .A2(n6000), .ZN(n6007) );
  NOR2_X1 U7535 ( .A1(n5983), .A2(n6416), .ZN(n6002) );
  MUX2_X1 U7536 ( .A(n6416), .B(n6002), .S(P2_IR_REG_2__SCAN_IN), .Z(n6004) );
  INV_X1 U7537 ( .A(n5950), .ZN(n6003) );
  INV_X1 U7538 ( .A(n9752), .ZN(n6005) );
  NAND2_X1 U7539 ( .A1(n6725), .A2(n10136), .ZN(n6330) );
  NAND2_X1 U7540 ( .A1(n6718), .A2(n7265), .ZN(n6358) );
  OAI211_X1 U7541 ( .C1(n6009), .C2(n6359), .A(n6330), .B(n6358), .ZN(n6010)
         );
  NAND2_X1 U7542 ( .A1(n6010), .A2(n7751), .ZN(n6014) );
  NAND2_X1 U7543 ( .A1(n6358), .A2(n6331), .ZN(n6011) );
  NAND3_X1 U7544 ( .A1(n6011), .A2(n7751), .A3(n6334), .ZN(n6012) );
  NAND2_X1 U7545 ( .A1(n6012), .A2(n6330), .ZN(n6013) );
  MUX2_X1 U7546 ( .A(n6014), .B(n6013), .S(n6288), .Z(n6015) );
  NAND2_X1 U7547 ( .A1(n6016), .A2(n6015), .ZN(n6017) );
  OAI21_X1 U7548 ( .B1(n6018), .B2(n6288), .A(n6017), .ZN(n6019) );
  NAND2_X1 U7549 ( .A1(n8349), .A2(n10151), .ZN(n6021) );
  NAND2_X1 U7550 ( .A1(n6019), .A2(n6021), .ZN(n6026) );
  AND2_X1 U7551 ( .A1(n7242), .A2(n6020), .ZN(n6022) );
  OAI211_X1 U7552 ( .C1(n6023), .C2(n6022), .A(n6021), .B(n6333), .ZN(n6024)
         );
  NAND2_X1 U7553 ( .A1(n6024), .A2(n6288), .ZN(n6025) );
  NAND2_X1 U7554 ( .A1(n6026), .A2(n6025), .ZN(n6043) );
  NAND2_X1 U7555 ( .A1(n6294), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n6036) );
  INV_X1 U7556 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n6027) );
  OR2_X1 U7557 ( .A1(n5931), .A2(n6027), .ZN(n6035) );
  INV_X1 U7558 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n6028) );
  OAI21_X1 U7559 ( .B1(n6030), .B2(n6029), .A(n6028), .ZN(n6032) );
  NAND2_X1 U7560 ( .A1(n6032), .A2(n6031), .ZN(n10080) );
  OR2_X1 U7561 ( .A1(n6251), .A2(n10080), .ZN(n6034) );
  INV_X1 U7562 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n6947) );
  OR2_X1 U7563 ( .A1(n6305), .A2(n6947), .ZN(n6033) );
  NAND4_X1 U7564 ( .A1(n6036), .A2(n6035), .A3(n6034), .A4(n6033), .ZN(n8348)
         );
  NAND2_X1 U7565 ( .A1(n6245), .A2(n6902), .ZN(n6041) );
  NAND2_X1 U7566 ( .A1(n6234), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n6040) );
  NAND2_X1 U7567 ( .A1(n6037), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6038) );
  XNOR2_X1 U7568 ( .A(n6038), .B(P2_IR_REG_7__SCAN_IN), .ZN(n6946) );
  NAND2_X1 U7569 ( .A1(n6186), .A2(n6946), .ZN(n6039) );
  OR2_X1 U7570 ( .A1(n8348), .A2(n10157), .ZN(n6065) );
  NAND2_X1 U7571 ( .A1(n8348), .A2(n10157), .ZN(n6045) );
  AOI21_X1 U7572 ( .B1(n6288), .B2(n10068), .A(n10077), .ZN(n6042) );
  NAND2_X1 U7573 ( .A1(n6043), .A2(n6042), .ZN(n6067) );
  OR2_X1 U7574 ( .A1(n8347), .A2(n10165), .ZN(n6366) );
  NAND2_X1 U7575 ( .A1(n6366), .A2(n6044), .ZN(n6336) );
  INV_X1 U7576 ( .A(n6045), .ZN(n6365) );
  NOR2_X1 U7577 ( .A1(n6336), .A2(n6365), .ZN(n6046) );
  INV_X1 U7578 ( .A(n6366), .ZN(n7705) );
  AOI21_X1 U7579 ( .B1(n6067), .B2(n6046), .A(n7705), .ZN(n6047) );
  MUX2_X1 U7580 ( .A(n6048), .B(n6047), .S(n6288), .Z(n6049) );
  NAND2_X1 U7581 ( .A1(n7834), .A2(n7805), .ZN(n6367) );
  NAND2_X1 U7582 ( .A1(n6049), .A2(n6367), .ZN(n6064) );
  INV_X1 U7583 ( .A(n6340), .ZN(n6062) );
  NAND2_X1 U7584 ( .A1(n6915), .A2(n6245), .ZN(n6052) );
  NAND2_X1 U7585 ( .A1(n6050), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6069) );
  XNOR2_X1 U7586 ( .A(n6069), .B(P2_IR_REG_10__SCAN_IN), .ZN(n7184) );
  AOI22_X1 U7587 ( .A1(n6234), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6186), .B2(
        n7184), .ZN(n6051) );
  NAND2_X1 U7588 ( .A1(n6294), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n6060) );
  INV_X1 U7589 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n7136) );
  OR2_X1 U7590 ( .A1(n5931), .A2(n7136), .ZN(n6059) );
  INV_X1 U7591 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n6053) );
  OAI21_X1 U7592 ( .B1(n6055), .B2(n6054), .A(n6053), .ZN(n6056) );
  NAND2_X1 U7593 ( .A1(n6056), .A2(n6074), .ZN(n7833) );
  OR2_X1 U7594 ( .A1(n6251), .A2(n7833), .ZN(n6058) );
  INV_X1 U7595 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7813) );
  OR2_X1 U7596 ( .A1(n6305), .A2(n7813), .ZN(n6057) );
  NAND2_X1 U7597 ( .A1(n10178), .A2(n7947), .ZN(n6338) );
  NAND2_X1 U7598 ( .A1(n6338), .A2(n6367), .ZN(n6061) );
  MUX2_X1 U7599 ( .A(n6062), .B(n6061), .S(n6315), .Z(n6063) );
  INV_X1 U7600 ( .A(n6339), .ZN(n6368) );
  NOR2_X1 U7601 ( .A1(n6063), .A2(n6368), .ZN(n6066) );
  NAND2_X1 U7602 ( .A1(n6064), .A2(n6066), .ZN(n6085) );
  NAND4_X1 U7603 ( .A1(n6067), .A2(n6066), .A3(n7684), .A4(n6065), .ZN(n6080)
         );
  NAND2_X1 U7604 ( .A1(n6919), .A2(n6245), .ZN(n6073) );
  INV_X1 U7605 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n6068) );
  NAND2_X1 U7606 ( .A1(n6069), .A2(n6068), .ZN(n6070) );
  NAND2_X1 U7607 ( .A1(n6070), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6071) );
  XNOR2_X1 U7608 ( .A(n6071), .B(P2_IR_REG_11__SCAN_IN), .ZN(n7339) );
  AOI22_X1 U7609 ( .A1(n6234), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n6186), .B2(
        n7339), .ZN(n6072) );
  NAND2_X1 U7610 ( .A1(n6294), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n6079) );
  INV_X1 U7611 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n7179) );
  OR2_X1 U7612 ( .A1(n6305), .A2(n7179), .ZN(n6078) );
  INV_X1 U7613 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n7945) );
  NAND2_X1 U7614 ( .A1(n6074), .A2(n7945), .ZN(n6075) );
  NAND2_X1 U7615 ( .A1(n6091), .A2(n6075), .ZN(n7946) );
  OR2_X1 U7616 ( .A1(n6251), .A2(n7946), .ZN(n6077) );
  INV_X1 U7617 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n7182) );
  OR2_X1 U7618 ( .A1(n5931), .A2(n7182), .ZN(n6076) );
  NAND3_X1 U7619 ( .A1(n6080), .A2(n6339), .A3(n7857), .ZN(n6083) );
  NAND2_X1 U7620 ( .A1(n7950), .A2(n8020), .ZN(n6370) );
  NAND2_X1 U7621 ( .A1(n6370), .A2(n6338), .ZN(n6081) );
  NAND2_X1 U7622 ( .A1(n7011), .A2(n6245), .ZN(n6089) );
  NAND2_X1 U7623 ( .A1(n6086), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6087) );
  XNOR2_X1 U7624 ( .A(n6087), .B(P2_IR_REG_12__SCAN_IN), .ZN(n8384) );
  AOI22_X1 U7625 ( .A1(n6234), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n6186), .B2(
        n8384), .ZN(n6088) );
  NAND2_X1 U7626 ( .A1(n6294), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n6096) );
  INV_X1 U7627 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n7340) );
  OR2_X1 U7628 ( .A1(n5931), .A2(n7340), .ZN(n6095) );
  NAND2_X1 U7629 ( .A1(n6091), .A2(n6090), .ZN(n6092) );
  NAND2_X1 U7630 ( .A1(n6106), .A2(n6092), .ZN(n8019) );
  OR2_X1 U7631 ( .A1(n6251), .A2(n8019), .ZN(n6094) );
  INV_X1 U7632 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n7332) );
  OR2_X1 U7633 ( .A1(n6305), .A2(n7332), .ZN(n6093) );
  NAND2_X1 U7634 ( .A1(n8023), .A2(n8049), .ZN(n6372) );
  AND2_X1 U7635 ( .A1(n6372), .A2(n6370), .ZN(n6098) );
  OR2_X1 U7636 ( .A1(n8023), .A2(n8049), .ZN(n6342) );
  INV_X1 U7637 ( .A(n6342), .ZN(n6097) );
  NAND2_X1 U7638 ( .A1(n6342), .A2(n7857), .ZN(n6373) );
  INV_X1 U7639 ( .A(n6373), .ZN(n6100) );
  INV_X1 U7640 ( .A(n6372), .ZN(n6099) );
  NAND2_X1 U7641 ( .A1(n7014), .A2(n6245), .ZN(n6104) );
  OR2_X1 U7642 ( .A1(n6102), .A2(n6416), .ZN(n6113) );
  XNOR2_X1 U7643 ( .A(n6113), .B(P2_IR_REG_13__SCAN_IN), .ZN(n7452) );
  AOI22_X1 U7644 ( .A1(n6234), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n6186), .B2(
        n7452), .ZN(n6103) );
  NAND2_X1 U7645 ( .A1(n6294), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n6111) );
  INV_X1 U7646 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n6105) );
  OR2_X1 U7647 ( .A1(n5931), .A2(n6105), .ZN(n6110) );
  INV_X1 U7648 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n9689) );
  NAND2_X1 U7649 ( .A1(n6106), .A2(n9689), .ZN(n6107) );
  NAND2_X1 U7650 ( .A1(n6122), .A2(n6107), .ZN(n8048) );
  OR2_X1 U7651 ( .A1(n6251), .A2(n8048), .ZN(n6109) );
  INV_X1 U7652 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n8003) );
  OR2_X1 U7653 ( .A1(n6305), .A2(n8003), .ZN(n6108) );
  OR2_X1 U7654 ( .A1(n8026), .A2(n8179), .ZN(n6129) );
  NAND2_X1 U7655 ( .A1(n8026), .A2(n8179), .ZN(n6374) );
  NAND2_X1 U7656 ( .A1(n6129), .A2(n6374), .ZN(n7996) );
  INV_X1 U7657 ( .A(n6131), .ZN(n6148) );
  NAND2_X1 U7658 ( .A1(n9733), .A2(n6245), .ZN(n6119) );
  NAND2_X1 U7659 ( .A1(n6113), .A2(n6112), .ZN(n6114) );
  NAND2_X1 U7660 ( .A1(n6114), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6116) );
  OR2_X1 U7661 ( .A1(n6116), .A2(n6115), .ZN(n6117) );
  NAND2_X1 U7662 ( .A1(n6116), .A2(n6115), .ZN(n6133) );
  AOI22_X1 U7663 ( .A1(n6234), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n7845), .B2(
        n6186), .ZN(n6118) );
  NAND2_X1 U7664 ( .A1(n6294), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n6128) );
  INV_X1 U7665 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n6120) );
  OR2_X1 U7666 ( .A1(n5931), .A2(n6120), .ZN(n6127) );
  NAND2_X1 U7667 ( .A1(n6122), .A2(n6121), .ZN(n6123) );
  NAND2_X1 U7668 ( .A1(n6139), .A2(n6123), .ZN(n8178) );
  OR2_X1 U7669 ( .A1(n6251), .A2(n8178), .ZN(n6126) );
  INV_X1 U7670 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n6124) );
  OR2_X1 U7671 ( .A1(n6305), .A2(n6124), .ZN(n6125) );
  NAND4_X1 U7672 ( .A1(n6128), .A2(n6127), .A3(n6126), .A4(n6125), .ZN(n8474)
         );
  XNOR2_X1 U7673 ( .A(n8475), .B(n8474), .ZN(n8029) );
  NAND3_X1 U7674 ( .A1(n8029), .A2(n6288), .A3(n6374), .ZN(n6147) );
  INV_X1 U7675 ( .A(n8474), .ZN(n8738) );
  AND2_X1 U7676 ( .A1(n8029), .A2(n6129), .ZN(n6130) );
  AOI22_X1 U7677 ( .A1(n6131), .A2(n6130), .B1(n8738), .B2(n8475), .ZN(n6132)
         );
  NAND2_X1 U7678 ( .A1(n7160), .A2(n6245), .ZN(n6136) );
  NAND2_X1 U7679 ( .A1(n6133), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6134) );
  XNOR2_X1 U7680 ( .A(n6134), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8404) );
  AOI22_X1 U7681 ( .A1(n8404), .A2(n6186), .B1(n6234), .B2(
        P1_DATAO_REG_15__SCAN_IN), .ZN(n6135) );
  NAND2_X1 U7682 ( .A1(n6304), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n6145) );
  INV_X1 U7683 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n6137) );
  OR2_X1 U7684 ( .A1(n6307), .A2(n6137), .ZN(n6144) );
  NAND2_X1 U7685 ( .A1(n6139), .A2(n6138), .ZN(n6140) );
  NAND2_X1 U7686 ( .A1(n6165), .A2(n6140), .ZN(n8329) );
  OR2_X1 U7687 ( .A1(n6251), .A2(n8329), .ZN(n6143) );
  INV_X1 U7688 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n6141) );
  OR2_X1 U7689 ( .A1(n6305), .A2(n6141), .ZN(n6142) );
  NAND2_X1 U7690 ( .A1(n8745), .A2(n8719), .ZN(n6375) );
  NAND2_X1 U7691 ( .A1(n6376), .A2(n6375), .ZN(n8734) );
  INV_X1 U7692 ( .A(n8734), .ZN(n6345) );
  OAI211_X1 U7693 ( .C1(n6148), .C2(n6147), .A(n6146), .B(n6345), .ZN(n6158)
         );
  NAND2_X1 U7694 ( .A1(n7158), .A2(n6245), .ZN(n6152) );
  OR2_X1 U7695 ( .A1(n6149), .A2(n6416), .ZN(n6150) );
  XNOR2_X1 U7696 ( .A(n6150), .B(P2_IR_REG_16__SCAN_IN), .ZN(n8420) );
  AOI22_X1 U7697 ( .A1(n6234), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n8420), .B2(
        n6186), .ZN(n6151) );
  NAND2_X1 U7698 ( .A1(n6294), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n6156) );
  INV_X1 U7699 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n8397) );
  OR2_X1 U7700 ( .A1(n5931), .A2(n8397), .ZN(n6155) );
  INV_X1 U7701 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n6164) );
  XNOR2_X1 U7702 ( .A(n6165), .B(n6164), .ZN(n8724) );
  OR2_X1 U7703 ( .A1(n6251), .A2(n8724), .ZN(n6154) );
  INV_X1 U7704 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8725) );
  OR2_X1 U7705 ( .A1(n6305), .A2(n8725), .ZN(n6153) );
  OR2_X1 U7706 ( .A1(n8825), .A2(n8737), .ZN(n6159) );
  NAND2_X1 U7707 ( .A1(n8825), .A2(n8737), .ZN(n6378) );
  NAND2_X1 U7708 ( .A1(n6159), .A2(n6378), .ZN(n8713) );
  INV_X1 U7709 ( .A(n8713), .ZN(n6346) );
  MUX2_X1 U7710 ( .A(n6375), .B(n6376), .S(n6315), .Z(n6157) );
  INV_X1 U7711 ( .A(n6159), .ZN(n6377) );
  MUX2_X1 U7712 ( .A(n6377), .B(n4515), .S(n6315), .Z(n6171) );
  NAND2_X1 U7713 ( .A1(n7208), .A2(n6245), .ZN(n6162) );
  NAND2_X1 U7714 ( .A1(n4471), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6160) );
  XNOR2_X1 U7715 ( .A(n6160), .B(P2_IR_REG_17__SCAN_IN), .ZN(n8432) );
  AOI22_X1 U7716 ( .A1(n8432), .A2(n6186), .B1(n6234), .B2(
        P1_DATAO_REG_17__SCAN_IN), .ZN(n6161) );
  NAND2_X1 U7717 ( .A1(n6294), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n6170) );
  INV_X1 U7718 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n9610) );
  OR2_X1 U7719 ( .A1(n5931), .A2(n9610), .ZN(n6169) );
  INV_X1 U7720 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n6163) );
  OAI21_X1 U7721 ( .B1(n6165), .B2(n6164), .A(n6163), .ZN(n6166) );
  NAND2_X1 U7722 ( .A1(n6175), .A2(n6166), .ZN(n8705) );
  OR2_X1 U7723 ( .A1(n6251), .A2(n8705), .ZN(n6168) );
  INV_X1 U7724 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8706) );
  OR2_X1 U7725 ( .A1(n6305), .A2(n8706), .ZN(n6167) );
  NAND2_X1 U7726 ( .A1(n8822), .A2(n8718), .ZN(n6182) );
  NAND2_X1 U7727 ( .A1(n6379), .A2(n6182), .ZN(n8695) );
  NOR2_X1 U7728 ( .A1(n6171), .A2(n8695), .ZN(n6185) );
  NAND2_X1 U7729 ( .A1(n7296), .A2(n6245), .ZN(n6174) );
  XNOR2_X1 U7730 ( .A(n6172), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8447) );
  AOI22_X1 U7731 ( .A1(n8447), .A2(n6186), .B1(n6234), .B2(
        P1_DATAO_REG_18__SCAN_IN), .ZN(n6173) );
  NAND2_X1 U7732 ( .A1(n6294), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n6181) );
  INV_X1 U7733 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8431) );
  OR2_X1 U7734 ( .A1(n5931), .A2(n8431), .ZN(n6180) );
  INV_X1 U7735 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n9520) );
  NAND2_X1 U7736 ( .A1(n6175), .A2(n9520), .ZN(n6176) );
  NAND2_X1 U7737 ( .A1(n6190), .A2(n6176), .ZN(n8295) );
  OR2_X1 U7738 ( .A1(n6251), .A2(n8295), .ZN(n6179) );
  INV_X1 U7739 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n6177) );
  OR2_X1 U7740 ( .A1(n6305), .A2(n6177), .ZN(n6178) );
  NAND4_X1 U7741 ( .A1(n6181), .A2(n6180), .A3(n6179), .A4(n6178), .ZN(n8481)
         );
  INV_X1 U7742 ( .A(n8481), .ZN(n8698) );
  INV_X1 U7743 ( .A(n6182), .ZN(n6183) );
  NAND2_X1 U7744 ( .A1(n8815), .A2(n8698), .ZN(n6380) );
  INV_X1 U7745 ( .A(n6380), .ZN(n6196) );
  NAND2_X1 U7746 ( .A1(n7349), .A2(n6245), .ZN(n6188) );
  AOI22_X1 U7747 ( .A1(n6322), .A2(n6186), .B1(n6234), .B2(
        P1_DATAO_REG_19__SCAN_IN), .ZN(n6187) );
  NAND2_X1 U7748 ( .A1(n6294), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n6195) );
  INV_X1 U7749 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n8450) );
  OR2_X1 U7750 ( .A1(n5931), .A2(n8450), .ZN(n6194) );
  NAND2_X1 U7751 ( .A1(n6190), .A2(n6189), .ZN(n6191) );
  NAND2_X1 U7752 ( .A1(n6200), .A2(n6191), .ZN(n8671) );
  OR2_X1 U7753 ( .A1(n6251), .A2(n8671), .ZN(n6193) );
  INV_X1 U7754 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n8672) );
  OR2_X1 U7755 ( .A1(n6305), .A2(n8672), .ZN(n6192) );
  NAND4_X1 U7756 ( .A1(n6195), .A2(n6194), .A3(n6193), .A4(n6192), .ZN(n8687)
         );
  INV_X1 U7757 ( .A(n8687), .ZN(n8484) );
  OR2_X1 U7758 ( .A1(n8811), .A2(n8484), .ZN(n6329) );
  NAND2_X1 U7759 ( .A1(n7493), .A2(n6245), .ZN(n6198) );
  NAND2_X1 U7760 ( .A1(n6234), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n6197) );
  NAND2_X1 U7761 ( .A1(n6304), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n6207) );
  INV_X1 U7762 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n9531) );
  OR2_X1 U7763 ( .A1(n6307), .A2(n9531), .ZN(n6206) );
  INV_X1 U7764 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n6199) );
  NAND2_X1 U7765 ( .A1(n6200), .A2(n6199), .ZN(n6201) );
  NAND2_X1 U7766 ( .A1(n6210), .A2(n6201), .ZN(n8645) );
  OR2_X1 U7767 ( .A1(n6202), .A2(n8645), .ZN(n6205) );
  INV_X1 U7768 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n6203) );
  OR2_X1 U7769 ( .A1(n6305), .A2(n6203), .ZN(n6204) );
  NAND2_X1 U7770 ( .A1(n8805), .A2(n8229), .ZN(n6328) );
  NAND2_X1 U7771 ( .A1(n8811), .A2(n8484), .ZN(n6382) );
  NAND2_X1 U7772 ( .A1(n7551), .A2(n6245), .ZN(n6209) );
  NAND2_X1 U7773 ( .A1(n6234), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n6208) );
  INV_X1 U7774 ( .A(n6251), .ZN(n6278) );
  NAND2_X1 U7775 ( .A1(n6210), .A2(n8231), .ZN(n6211) );
  AND2_X1 U7776 ( .A1(n6212), .A2(n6211), .ZN(n8632) );
  NAND2_X1 U7777 ( .A1(n6278), .A2(n8632), .ZN(n6219) );
  INV_X1 U7778 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n6213) );
  OR2_X1 U7779 ( .A1(n5931), .A2(n6213), .ZN(n6218) );
  INV_X1 U7780 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n6214) );
  OR2_X1 U7781 ( .A1(n6307), .A2(n6214), .ZN(n6217) );
  INV_X1 U7782 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n6215) );
  OR2_X1 U7783 ( .A1(n6305), .A2(n6215), .ZN(n6216) );
  NAND4_X1 U7784 ( .A1(n6219), .A2(n6218), .A3(n6217), .A4(n6216), .ZN(n8652)
         );
  INV_X1 U7785 ( .A(n8652), .ZN(n8623) );
  OR2_X1 U7786 ( .A1(n8800), .A2(n8623), .ZN(n6230) );
  NAND3_X1 U7787 ( .A1(n6220), .A2(n6383), .A3(n6230), .ZN(n6221) );
  NAND2_X1 U7788 ( .A1(n8800), .A2(n8623), .ZN(n6384) );
  NAND3_X1 U7789 ( .A1(n6221), .A2(n6327), .A3(n6384), .ZN(n6222) );
  NAND2_X1 U7790 ( .A1(n6222), .A2(n6385), .ZN(n6223) );
  INV_X1 U7791 ( .A(n8490), .ZN(n8624) );
  NAND2_X1 U7792 ( .A1(n8789), .A2(n8624), .ZN(n6387) );
  INV_X1 U7793 ( .A(n8609), .ZN(n6386) );
  INV_X1 U7794 ( .A(n8660), .ZN(n6226) );
  OAI211_X1 U7795 ( .C1(n6227), .C2(n6226), .A(n6380), .B(n6382), .ZN(n6228)
         );
  NAND3_X1 U7796 ( .A1(n6228), .A2(n6329), .A3(n6383), .ZN(n6229) );
  NAND3_X1 U7797 ( .A1(n6229), .A2(n6328), .A3(n6384), .ZN(n6231) );
  NAND4_X1 U7798 ( .A1(n6231), .A2(n6288), .A3(n6230), .A4(n6385), .ZN(n6232)
         );
  NAND2_X1 U7799 ( .A1(n8783), .A2(n8263), .ZN(n6326) );
  NAND2_X1 U7800 ( .A1(n8010), .A2(n6245), .ZN(n6236) );
  NAND2_X1 U7801 ( .A1(n6234), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n6235) );
  INV_X1 U7802 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n6237) );
  NAND2_X1 U7803 ( .A1(n6238), .A2(n6237), .ZN(n6239) );
  AND2_X1 U7804 ( .A1(n6249), .A2(n6239), .ZN(n8577) );
  NAND2_X1 U7805 ( .A1(n8577), .A2(n6278), .ZN(n6244) );
  INV_X1 U7806 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n8579) );
  NAND2_X1 U7807 ( .A1(n6294), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n6241) );
  NAND2_X1 U7808 ( .A1(n6304), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n6240) );
  OAI211_X1 U7809 ( .C1(n6305), .C2(n8579), .A(n6241), .B(n6240), .ZN(n6242)
         );
  INV_X1 U7810 ( .A(n6242), .ZN(n6243) );
  NAND2_X1 U7811 ( .A1(n8779), .A2(n8592), .ZN(n6259) );
  NAND2_X1 U7812 ( .A1(n6234), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n6246) );
  INV_X1 U7813 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n6248) );
  NAND2_X1 U7814 ( .A1(n6249), .A2(n6248), .ZN(n6250) );
  NAND2_X1 U7815 ( .A1(n6273), .A2(n6250), .ZN(n8552) );
  OR2_X1 U7816 ( .A1(n8552), .A2(n6251), .ZN(n6257) );
  INV_X1 U7817 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n6254) );
  NAND2_X1 U7818 ( .A1(n6304), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n6253) );
  NAND2_X1 U7819 ( .A1(n6294), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n6252) );
  OAI211_X1 U7820 ( .C1(n6254), .C2(n6305), .A(n6253), .B(n6252), .ZN(n6255)
         );
  INV_X1 U7821 ( .A(n6255), .ZN(n6256) );
  INV_X1 U7822 ( .A(n6263), .ZN(n6258) );
  NAND2_X1 U7823 ( .A1(n6258), .A2(n6390), .ZN(n6261) );
  NAND2_X1 U7824 ( .A1(n8493), .A2(n6259), .ZN(n6260) );
  MUX2_X1 U7825 ( .A(n6261), .B(n6260), .S(n6315), .Z(n6262) );
  MUX2_X1 U7826 ( .A(n6392), .B(n6263), .S(n6315), .Z(n6270) );
  NAND2_X1 U7827 ( .A1(n8055), .A2(n6245), .ZN(n6265) );
  NAND2_X1 U7828 ( .A1(n6234), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n6264) );
  XNOR2_X1 U7829 ( .A(n6273), .B(P2_REG3_REG_27__SCAN_IN), .ZN(n8534) );
  INV_X1 U7830 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n6268) );
  NAND2_X1 U7831 ( .A1(n6304), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n6267) );
  NAND2_X1 U7832 ( .A1(n6294), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n6266) );
  OAI211_X1 U7833 ( .C1(n6268), .C2(n6305), .A(n6267), .B(n6266), .ZN(n6269)
         );
  AOI21_X1 U7834 ( .B1(n8534), .B2(n6278), .A(n6269), .ZN(n8339) );
  NAND2_X1 U7835 ( .A1(n8768), .A2(n8339), .ZN(n6279) );
  NAND2_X1 U7836 ( .A1(n6234), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n6271) );
  INV_X1 U7837 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n8166) );
  INV_X1 U7838 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n6272) );
  OAI21_X1 U7839 ( .B1(n6273), .B2(n8166), .A(n6272), .ZN(n6274) );
  INV_X1 U7840 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n8518) );
  NAND2_X1 U7841 ( .A1(n6304), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n6276) );
  NAND2_X1 U7842 ( .A1(n6294), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n6275) );
  OAI211_X1 U7843 ( .C1(n8518), .C2(n6305), .A(n6276), .B(n6275), .ZN(n6277)
         );
  AOI21_X1 U7844 ( .B1(n8216), .B2(n6278), .A(n6277), .ZN(n8544) );
  NAND2_X1 U7845 ( .A1(n8763), .A2(n8544), .ZN(n6325) );
  INV_X1 U7846 ( .A(n6325), .ZN(n6283) );
  INV_X1 U7847 ( .A(n6279), .ZN(n6280) );
  MUX2_X1 U7848 ( .A(n6281), .B(n6280), .S(n6315), .Z(n6282) );
  INV_X1 U7849 ( .A(n8544), .ZN(n8505) );
  OAI21_X1 U7850 ( .B1(n6286), .B2(n8505), .A(n8499), .ZN(n6285) );
  OAI21_X1 U7851 ( .B1(n6394), .B2(n6315), .A(n6285), .ZN(n6291) );
  INV_X1 U7852 ( .A(n6286), .ZN(n6287) );
  OAI211_X1 U7853 ( .C1(n6288), .C2(n8763), .A(n6287), .B(n6325), .ZN(n6290)
         );
  MUX2_X1 U7854 ( .A(n6395), .B(n6394), .S(n6315), .Z(n6289) );
  AOI21_X1 U7855 ( .B1(n6291), .B2(n6290), .A(n6289), .ZN(n6301) );
  NAND2_X1 U7856 ( .A1(n8849), .A2(n6245), .ZN(n6293) );
  NAND2_X1 U7857 ( .A1(n6234), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n6292) );
  INV_X1 U7858 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n6297) );
  NAND2_X1 U7859 ( .A1(n6304), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n6296) );
  NAND2_X1 U7860 ( .A1(n6294), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n6295) );
  OAI211_X1 U7861 ( .C1(n6305), .C2(n6297), .A(n6296), .B(n6295), .ZN(n8503)
         );
  NAND2_X1 U7862 ( .A1(n9792), .A2(n8503), .ZN(n6398) );
  INV_X1 U7863 ( .A(n6398), .ZN(n6300) );
  INV_X1 U7864 ( .A(n8503), .ZN(n6298) );
  NAND2_X1 U7865 ( .A1(n8470), .A2(n6298), .ZN(n6311) );
  INV_X1 U7866 ( .A(n6311), .ZN(n6299) );
  NOR3_X1 U7867 ( .A1(n6301), .A2(n6300), .A3(n6299), .ZN(n6313) );
  NAND2_X1 U7868 ( .A1(n8845), .A2(n6245), .ZN(n6303) );
  NAND2_X1 U7869 ( .A1(n5999), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n6302) );
  NAND2_X1 U7870 ( .A1(n6304), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n6310) );
  INV_X1 U7871 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n8462) );
  OR2_X1 U7872 ( .A1(n6305), .A2(n8462), .ZN(n6309) );
  INV_X1 U7873 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n6306) );
  OR2_X1 U7874 ( .A1(n6307), .A2(n6306), .ZN(n6308) );
  AND3_X1 U7875 ( .A1(n6310), .A2(n6309), .A3(n6308), .ZN(n6921) );
  NAND2_X1 U7876 ( .A1(n6403), .A2(n6398), .ZN(n6352) );
  INV_X1 U7877 ( .A(n6403), .ZN(n6317) );
  INV_X1 U7878 ( .A(n6314), .ZN(n6316) );
  MUX2_X1 U7879 ( .A(n6317), .B(n6316), .S(n6315), .Z(n6321) );
  XNOR2_X1 U7880 ( .A(n8800), .B(n8623), .ZN(n8635) );
  NAND2_X1 U7881 ( .A1(n6383), .A2(n6328), .ZN(n8642) );
  INV_X1 U7882 ( .A(n8642), .ZN(n8651) );
  INV_X1 U7883 ( .A(n8663), .ZN(n8658) );
  NAND2_X1 U7884 ( .A1(n8660), .A2(n6380), .ZN(n8682) );
  AND2_X1 U7885 ( .A1(n7751), .A2(n6330), .ZN(n7895) );
  NAND2_X1 U7886 ( .A1(n7772), .A2(n6331), .ZN(n10125) );
  NOR4_X1 U7887 ( .A1(n7892), .A2(n10125), .A3(n7750), .A4(n8059), .ZN(n6335)
         );
  INV_X1 U7888 ( .A(n10101), .ZN(n6362) );
  NAND2_X1 U7889 ( .A1(n6364), .A2(n6333), .ZN(n7243) );
  INV_X1 U7890 ( .A(n7243), .ZN(n7666) );
  INV_X1 U7891 ( .A(n7773), .ZN(n7769) );
  NAND4_X1 U7892 ( .A1(n6335), .A2(n6362), .A3(n7666), .A4(n7769), .ZN(n6337)
         );
  XNOR2_X1 U7893 ( .A(n8349), .B(n10151), .ZN(n7736) );
  NOR4_X1 U7894 ( .A1(n6337), .A2(n7736), .A3(n6336), .A4(n10077), .ZN(n6341)
         );
  NAND2_X1 U7895 ( .A1(n6339), .A2(n6338), .ZN(n7809) );
  INV_X1 U7896 ( .A(n7809), .ZN(n6369) );
  NAND3_X1 U7897 ( .A1(n6341), .A2(n6369), .A3(n7704), .ZN(n6343) );
  NAND2_X1 U7898 ( .A1(n7857), .A2(n6370), .ZN(n7927) );
  NOR4_X1 U7899 ( .A1(n6343), .A2(n4412), .A3(n7996), .A4(n7927), .ZN(n6344)
         );
  NAND4_X1 U7900 ( .A1(n6346), .A2(n6345), .A3(n6344), .A4(n8029), .ZN(n6347)
         );
  NOR4_X1 U7901 ( .A1(n8658), .A2(n8695), .A3(n8682), .A4(n6347), .ZN(n6348)
         );
  NAND4_X1 U7902 ( .A1(n8609), .A2(n8489), .A3(n8651), .A4(n6348), .ZN(n6349)
         );
  NOR4_X1 U7903 ( .A1(n8569), .A2(n8635), .A3(n8591), .A4(n6349), .ZN(n6350)
         );
  INV_X1 U7904 ( .A(n8499), .ZN(n8501) );
  INV_X1 U7905 ( .A(n8059), .ZN(n6406) );
  OAI22_X1 U7906 ( .A1(n6355), .A2(n6819), .B1(n6406), .B2(n6717), .ZN(n6356)
         );
  INV_X1 U7907 ( .A(n6360), .ZN(n6361) );
  NAND2_X1 U7908 ( .A1(n10088), .A2(n6362), .ZN(n7241) );
  INV_X1 U7909 ( .A(n6370), .ZN(n6371) );
  OAI21_X1 U7910 ( .B1(n7859), .B2(n6373), .A(n6372), .ZN(n7999) );
  OAI21_X1 U7911 ( .B1(n8696), .B2(n8695), .A(n6379), .ZN(n8683) );
  NAND2_X1 U7912 ( .A1(n8683), .A2(n6380), .ZN(n8661) );
  INV_X1 U7913 ( .A(n8591), .ZN(n6388) );
  NAND2_X1 U7914 ( .A1(n8594), .A2(n6389), .ZN(n8567) );
  INV_X1 U7915 ( .A(n8493), .ZN(n8557) );
  INV_X1 U7916 ( .A(n6390), .ZN(n8558) );
  NOR2_X1 U7917 ( .A1(n8557), .A2(n8558), .ZN(n6391) );
  NAND2_X1 U7918 ( .A1(n8556), .A2(n6391), .ZN(n8538) );
  INV_X1 U7919 ( .A(n6392), .ZN(n8540) );
  NAND2_X1 U7920 ( .A1(n8538), .A2(n4953), .ZN(n8537) );
  NAND2_X1 U7921 ( .A1(n8537), .A2(n6393), .ZN(n8521) );
  INV_X1 U7922 ( .A(n6395), .ZN(n6396) );
  INV_X1 U7923 ( .A(n6397), .ZN(n6405) );
  NAND2_X1 U7924 ( .A1(n6399), .A2(n6398), .ZN(n6402) );
  NAND2_X1 U7925 ( .A1(n6406), .A2(n6819), .ZN(n7245) );
  NAND2_X1 U7926 ( .A1(n6726), .A2(n7245), .ZN(n6407) );
  NAND2_X1 U7927 ( .A1(n6408), .A2(n6411), .ZN(n6409) );
  NAND2_X1 U7928 ( .A1(n6409), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6423) );
  XNOR2_X1 U7929 ( .A(n6423), .B(P2_IR_REG_23__SCAN_IN), .ZN(n6822) );
  AND2_X1 U7930 ( .A1(n6822), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7718) );
  NAND3_X1 U7931 ( .A1(n6411), .A2(n6422), .A3(n6425), .ZN(n6412) );
  NOR2_X1 U7932 ( .A1(n6413), .A2(n6412), .ZN(n6417) );
  NAND2_X1 U7933 ( .A1(n6417), .A2(n6418), .ZN(n6420) );
  NAND2_X1 U7934 ( .A1(n6420), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6414) );
  MUX2_X1 U7935 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6414), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n6415) );
  NAND2_X1 U7936 ( .A1(n6415), .A2(n5827), .ZN(n8042) );
  OR2_X1 U7937 ( .A1(n6417), .A2(n6416), .ZN(n6419) );
  MUX2_X1 U7938 ( .A(n6419), .B(P2_IR_REG_31__SCAN_IN), .S(n6418), .Z(n6421)
         );
  NAND2_X1 U7939 ( .A1(n6421), .A2(n6420), .ZN(n8011) );
  NOR2_X1 U7940 ( .A1(n8042), .A2(n8011), .ZN(n6428) );
  NAND2_X1 U7941 ( .A1(n6423), .A2(n6422), .ZN(n6424) );
  NAND2_X1 U7942 ( .A1(n6424), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6426) );
  XNOR2_X1 U7943 ( .A(n6426), .B(n6425), .ZN(n7939) );
  INV_X1 U7944 ( .A(n7939), .ZN(n6427) );
  NAND2_X1 U7945 ( .A1(n6428), .A2(n6427), .ZN(n6824) );
  NOR2_X1 U7946 ( .A1(n6822), .A2(P2_U3152), .ZN(n10119) );
  NAND2_X1 U7947 ( .A1(n6824), .A2(n10119), .ZN(n10110) );
  INV_X1 U7948 ( .A(n6930), .ZN(n8857) );
  NOR4_X1 U7949 ( .A1(n6410), .A2(n8464), .A3(n10110), .A4(n10072), .ZN(n6431)
         );
  INV_X1 U7950 ( .A(n7718), .ZN(n6926) );
  OAI21_X1 U7951 ( .B1(n6926), .B2(n6429), .A(P2_B_REG_SCAN_IN), .ZN(n6430) );
  OR2_X1 U7952 ( .A1(n6431), .A2(n6430), .ZN(n6432) );
  INV_X1 U7953 ( .A(n6834), .ZN(n6436) );
  INV_X1 U7954 ( .A(n6866), .ZN(n6438) );
  NAND2_X1 U7955 ( .A1(n6437), .A2(n9086), .ZN(n7372) );
  NAND2_X1 U7956 ( .A1(n7372), .A2(n6694), .ZN(n6497) );
  NAND2_X1 U7957 ( .A1(n6438), .A2(n6497), .ZN(n6439) );
  NAND2_X1 U7958 ( .A1(n6865), .A2(n6439), .ZN(n6447) );
  INV_X1 U7959 ( .A(n6447), .ZN(n6445) );
  NAND2_X1 U7960 ( .A1(n6435), .A2(n7522), .ZN(n6442) );
  NAND2_X1 U7961 ( .A1(n6458), .A2(n6440), .ZN(n6441) );
  NAND2_X1 U7962 ( .A1(n6442), .A2(n6441), .ZN(n6443) );
  XNOR2_X1 U7963 ( .A(n6443), .B(n6547), .ZN(n6446) );
  INV_X1 U7964 ( .A(n6446), .ZN(n6444) );
  NAND2_X1 U7965 ( .A1(n6445), .A2(n6444), .ZN(n7126) );
  AOI22_X1 U7966 ( .A1(n6658), .A2(n6440), .B1(n6458), .B2(n7522), .ZN(n7128)
         );
  NAND2_X1 U7967 ( .A1(n7126), .A2(n7128), .ZN(n6448) );
  NAND2_X1 U7968 ( .A1(n6447), .A2(n6446), .ZN(n7127) );
  NAND2_X1 U7969 ( .A1(n6458), .A2(n9018), .ZN(n6450) );
  NAND2_X1 U7970 ( .A1(n6435), .A2(n7520), .ZN(n6449) );
  AOI22_X1 U7971 ( .A1(n6658), .A2(n9018), .B1(n6458), .B2(n7520), .ZN(n6453)
         );
  NAND2_X1 U7972 ( .A1(n6452), .A2(n6453), .ZN(n6457) );
  INV_X1 U7973 ( .A(n6452), .ZN(n6455) );
  INV_X1 U7974 ( .A(n6453), .ZN(n6454) );
  NAND2_X1 U7975 ( .A1(n6455), .A2(n6454), .ZN(n6456) );
  NAND2_X1 U7976 ( .A1(n6458), .A2(n9017), .ZN(n6460) );
  NAND2_X1 U7977 ( .A1(n6435), .A2(n7566), .ZN(n6459) );
  NAND2_X1 U7978 ( .A1(n6460), .A2(n6459), .ZN(n6461) );
  XNOR2_X1 U7979 ( .A(n6461), .B(n6547), .ZN(n6464) );
  OAI22_X1 U7980 ( .A1(n6665), .A2(n7514), .B1(n10003), .B2(n6473), .ZN(n6462)
         );
  INV_X1 U7981 ( .A(n6462), .ZN(n6463) );
  NAND2_X1 U7982 ( .A1(n6464), .A2(n6463), .ZN(n6465) );
  NAND2_X1 U7983 ( .A1(n4395), .A2(n9016), .ZN(n6467) );
  NAND2_X1 U7984 ( .A1(n6646), .A2(n10009), .ZN(n6466) );
  NAND2_X1 U7985 ( .A1(n6467), .A2(n6466), .ZN(n6468) );
  XNOR2_X1 U7986 ( .A(n6468), .B(n6547), .ZN(n6469) );
  AOI22_X1 U7987 ( .A1(n6658), .A2(n9016), .B1(n4395), .B2(n10009), .ZN(n6470)
         );
  AND2_X1 U7988 ( .A1(n6469), .A2(n6470), .ZN(n7194) );
  INV_X1 U7989 ( .A(n6469), .ZN(n6472) );
  INV_X1 U7990 ( .A(n6470), .ZN(n6471) );
  NAND2_X1 U7991 ( .A1(n6472), .A2(n6471), .ZN(n7195) );
  NAND2_X1 U7992 ( .A1(n4395), .A2(n9014), .ZN(n6475) );
  NAND2_X1 U7993 ( .A1(n6646), .A2(n7615), .ZN(n6474) );
  NAND2_X1 U7994 ( .A1(n6475), .A2(n6474), .ZN(n6476) );
  XNOR2_X1 U7995 ( .A(n6476), .B(n6547), .ZN(n7439) );
  NAND2_X1 U7996 ( .A1(n6658), .A2(n9014), .ZN(n6478) );
  NAND2_X1 U7997 ( .A1(n4395), .A2(n7615), .ZN(n6477) );
  AND2_X1 U7998 ( .A1(n6478), .A2(n6477), .ZN(n7438) );
  NAND2_X1 U7999 ( .A1(n7439), .A2(n7438), .ZN(n7437) );
  NAND2_X1 U8000 ( .A1(n6458), .A2(n9015), .ZN(n6480) );
  NAND2_X1 U8001 ( .A1(n6646), .A2(n7462), .ZN(n6479) );
  NAND2_X1 U8002 ( .A1(n6480), .A2(n6479), .ZN(n6481) );
  NAND2_X1 U8003 ( .A1(n6658), .A2(n9015), .ZN(n6483) );
  NAND2_X1 U8004 ( .A1(n4395), .A2(n7462), .ZN(n6482) );
  AND2_X1 U8005 ( .A1(n6483), .A2(n6482), .ZN(n7354) );
  NAND2_X1 U8006 ( .A1(n7352), .A2(n7354), .ZN(n6484) );
  AND2_X1 U8007 ( .A1(n7437), .A2(n6484), .ZN(n6485) );
  NAND2_X1 U8008 ( .A1(n7351), .A2(n6485), .ZN(n6492) );
  OAI21_X1 U8009 ( .B1(n7352), .B2(n7354), .A(n7438), .ZN(n6490) );
  INV_X1 U8010 ( .A(n7439), .ZN(n6489) );
  INV_X1 U8011 ( .A(n7354), .ZN(n6487) );
  INV_X1 U8012 ( .A(n7438), .ZN(n6486) );
  AND2_X1 U8013 ( .A1(n6487), .A2(n6486), .ZN(n6488) );
  INV_X1 U8014 ( .A(n7352), .ZN(n7436) );
  AOI22_X1 U8015 ( .A1(n6490), .A2(n6489), .B1(n6488), .B2(n7436), .ZN(n6491)
         );
  NAND2_X1 U8016 ( .A1(n6492), .A2(n6491), .ZN(n7322) );
  NAND2_X1 U8017 ( .A1(n6658), .A2(n9013), .ZN(n6494) );
  NAND2_X1 U8018 ( .A1(n4395), .A2(n7481), .ZN(n6493) );
  NAND2_X1 U8019 ( .A1(n6494), .A2(n6493), .ZN(n7324) );
  NAND2_X1 U8020 ( .A1(n4395), .A2(n9013), .ZN(n6496) );
  NAND2_X1 U8021 ( .A1(n6646), .A2(n7481), .ZN(n6495) );
  NAND2_X1 U8022 ( .A1(n6496), .A2(n6495), .ZN(n6498) );
  XNOR2_X1 U8023 ( .A(n6498), .B(n7466), .ZN(n7323) );
  NAND2_X1 U8024 ( .A1(n7322), .A2(n7324), .ZN(n6499) );
  NAND2_X1 U8025 ( .A1(n6500), .A2(n6499), .ZN(n7391) );
  NAND2_X1 U8026 ( .A1(n6658), .A2(n9012), .ZN(n6502) );
  NAND2_X1 U8027 ( .A1(n4395), .A2(n7633), .ZN(n6501) );
  NAND2_X1 U8028 ( .A1(n6502), .A2(n6501), .ZN(n7389) );
  NAND2_X1 U8029 ( .A1(n4395), .A2(n9012), .ZN(n6504) );
  NAND2_X1 U8030 ( .A1(n7633), .A2(n6646), .ZN(n6503) );
  NAND2_X1 U8031 ( .A1(n6504), .A2(n6503), .ZN(n6505) );
  XNOR2_X1 U8032 ( .A(n6505), .B(n7466), .ZN(n7388) );
  NAND2_X1 U8033 ( .A1(n7647), .A2(n6646), .ZN(n6507) );
  NAND2_X1 U8034 ( .A1(n4395), .A2(n9011), .ZN(n6506) );
  NAND2_X1 U8035 ( .A1(n6507), .A2(n6506), .ZN(n6508) );
  XNOR2_X1 U8036 ( .A(n6508), .B(n6547), .ZN(n6511) );
  NAND2_X1 U8037 ( .A1(n7647), .A2(n4395), .ZN(n6510) );
  NAND2_X1 U8038 ( .A1(n6658), .A2(n9011), .ZN(n6509) );
  AND2_X1 U8039 ( .A1(n6510), .A2(n6509), .ZN(n6512) );
  NAND2_X1 U8040 ( .A1(n6511), .A2(n6512), .ZN(n6516) );
  INV_X1 U8041 ( .A(n6511), .ZN(n6514) );
  INV_X1 U8042 ( .A(n6512), .ZN(n6513) );
  NAND2_X1 U8043 ( .A1(n6514), .A2(n6513), .ZN(n6515) );
  NAND2_X1 U8044 ( .A1(n6516), .A2(n6515), .ZN(n7587) );
  NAND2_X1 U8045 ( .A1(n7585), .A2(n6516), .ZN(n7574) );
  NAND2_X1 U8046 ( .A1(n7868), .A2(n6646), .ZN(n6518) );
  NAND2_X1 U8047 ( .A1(n4395), .A2(n9010), .ZN(n6517) );
  NAND2_X1 U8048 ( .A1(n6518), .A2(n6517), .ZN(n6519) );
  XNOR2_X1 U8049 ( .A(n6519), .B(n7466), .ZN(n6522) );
  NAND2_X1 U8050 ( .A1(n7868), .A2(n4395), .ZN(n6521) );
  NAND2_X1 U8051 ( .A1(n6658), .A2(n9010), .ZN(n6520) );
  NAND2_X1 U8052 ( .A1(n6521), .A2(n6520), .ZN(n6523) );
  NAND2_X1 U8053 ( .A1(n6522), .A2(n6523), .ZN(n7576) );
  INV_X1 U8054 ( .A(n6522), .ZN(n6525) );
  INV_X1 U8055 ( .A(n6523), .ZN(n6524) );
  NAND2_X1 U8056 ( .A1(n6525), .A2(n6524), .ZN(n7575) );
  NAND2_X1 U8057 ( .A1(n9849), .A2(n6646), .ZN(n6528) );
  NAND2_X1 U8058 ( .A1(n4395), .A2(n9009), .ZN(n6527) );
  NAND2_X1 U8059 ( .A1(n6528), .A2(n6527), .ZN(n6529) );
  XNOR2_X1 U8060 ( .A(n6529), .B(n6547), .ZN(n6532) );
  NOR2_X1 U8061 ( .A1(n6665), .A2(n7989), .ZN(n6530) );
  AOI21_X1 U8062 ( .B1(n9849), .B2(n4395), .A(n6530), .ZN(n6533) );
  XNOR2_X1 U8063 ( .A(n6532), .B(n6533), .ZN(n7721) );
  INV_X1 U8064 ( .A(n6532), .ZN(n6535) );
  INV_X1 U8065 ( .A(n6533), .ZN(n6534) );
  NAND2_X1 U8066 ( .A1(n6535), .A2(n6534), .ZN(n6536) );
  NAND2_X1 U8067 ( .A1(n7991), .A2(n6646), .ZN(n6538) );
  NAND2_X1 U8068 ( .A1(n4395), .A2(n9008), .ZN(n6537) );
  NAND2_X1 U8069 ( .A1(n6538), .A2(n6537), .ZN(n6539) );
  XNOR2_X1 U8070 ( .A(n6539), .B(n6547), .ZN(n6543) );
  NOR2_X1 U8071 ( .A1(n6665), .A2(n9845), .ZN(n6540) );
  AOI21_X1 U8072 ( .B1(n7991), .B2(n4395), .A(n6540), .ZN(n6542) );
  XNOR2_X1 U8073 ( .A(n6543), .B(n6542), .ZN(n7985) );
  NAND2_X1 U8074 ( .A1(n6543), .A2(n6542), .ZN(n6544) );
  NAND2_X1 U8075 ( .A1(n7982), .A2(n6544), .ZN(n7973) );
  NAND2_X1 U8076 ( .A1(n7979), .A2(n6646), .ZN(n6546) );
  NAND2_X1 U8077 ( .A1(n4395), .A2(n9007), .ZN(n6545) );
  NAND2_X1 U8078 ( .A1(n6546), .A2(n6545), .ZN(n6548) );
  XNOR2_X1 U8079 ( .A(n6548), .B(n6547), .ZN(n7971) );
  NOR2_X1 U8080 ( .A1(n6665), .A2(n6549), .ZN(n6550) );
  AOI21_X1 U8081 ( .B1(n7979), .B2(n4395), .A(n6550), .ZN(n7970) );
  AND2_X1 U8082 ( .A1(n7971), .A2(n7970), .ZN(n6554) );
  INV_X1 U8083 ( .A(n7971), .ZN(n6552) );
  INV_X1 U8084 ( .A(n7970), .ZN(n6551) );
  NAND2_X1 U8085 ( .A1(n6552), .A2(n6551), .ZN(n6553) );
  NAND2_X1 U8086 ( .A1(n9416), .A2(n6646), .ZN(n6556) );
  NAND2_X1 U8087 ( .A1(n4395), .A2(n9006), .ZN(n6555) );
  NAND2_X1 U8088 ( .A1(n6556), .A2(n6555), .ZN(n6557) );
  XNOR2_X1 U8089 ( .A(n6557), .B(n7466), .ZN(n8872) );
  INV_X1 U8090 ( .A(n8872), .ZN(n6560) );
  NAND2_X1 U8091 ( .A1(n9416), .A2(n4395), .ZN(n6559) );
  NAND2_X1 U8092 ( .A1(n6658), .A2(n9006), .ZN(n6558) );
  NAND2_X1 U8093 ( .A1(n6559), .A2(n6558), .ZN(n6564) );
  INV_X1 U8094 ( .A(n6564), .ZN(n8871) );
  NAND2_X1 U8095 ( .A1(n6560), .A2(n8871), .ZN(n6572) );
  NAND2_X1 U8096 ( .A1(n8870), .A2(n6572), .ZN(n6568) );
  NAND2_X1 U8097 ( .A1(n9408), .A2(n6646), .ZN(n6562) );
  NAND2_X1 U8098 ( .A1(n4395), .A2(n9005), .ZN(n6561) );
  NAND2_X1 U8099 ( .A1(n6562), .A2(n6561), .ZN(n6563) );
  XNOR2_X1 U8100 ( .A(n6563), .B(n7466), .ZN(n6571) );
  INV_X1 U8101 ( .A(n6571), .ZN(n6566) );
  AND2_X1 U8102 ( .A1(n8872), .A2(n6564), .ZN(n6573) );
  INV_X1 U8103 ( .A(n6573), .ZN(n6565) );
  AND2_X1 U8104 ( .A1(n6566), .A2(n6565), .ZN(n6567) );
  NAND2_X1 U8105 ( .A1(n6568), .A2(n6567), .ZN(n8986) );
  NAND2_X1 U8106 ( .A1(n9408), .A2(n4395), .ZN(n6570) );
  NAND2_X1 U8107 ( .A1(n6658), .A2(n9005), .ZN(n6569) );
  NAND2_X1 U8108 ( .A1(n6570), .A2(n6569), .ZN(n8989) );
  NAND2_X1 U8109 ( .A1(n9405), .A2(n6646), .ZN(n6575) );
  NAND2_X1 U8110 ( .A1(n4395), .A2(n9288), .ZN(n6574) );
  NAND2_X1 U8111 ( .A1(n6575), .A2(n6574), .ZN(n6576) );
  XNOR2_X1 U8112 ( .A(n6576), .B(n7466), .ZN(n6579) );
  NAND2_X1 U8113 ( .A1(n9405), .A2(n4395), .ZN(n6578) );
  NAND2_X1 U8114 ( .A1(n6658), .A2(n9288), .ZN(n6577) );
  NAND2_X1 U8115 ( .A1(n6578), .A2(n6577), .ZN(n6580) );
  AND2_X1 U8116 ( .A1(n6579), .A2(n6580), .ZN(n8917) );
  INV_X1 U8117 ( .A(n6579), .ZN(n6582) );
  INV_X1 U8118 ( .A(n6580), .ZN(n6581) );
  NAND2_X1 U8119 ( .A1(n6582), .A2(n6581), .ZN(n8915) );
  NAND2_X1 U8120 ( .A1(n9398), .A2(n6646), .ZN(n6584) );
  NAND2_X1 U8121 ( .A1(n4395), .A2(n9004), .ZN(n6583) );
  NAND2_X1 U8122 ( .A1(n6584), .A2(n6583), .ZN(n6585) );
  XNOR2_X1 U8123 ( .A(n6585), .B(n7466), .ZN(n6587) );
  NOR2_X1 U8124 ( .A1(n6665), .A2(n9299), .ZN(n6586) );
  AOI21_X1 U8125 ( .B1(n9398), .B2(n4395), .A(n6586), .ZN(n6588) );
  XNOR2_X1 U8126 ( .A(n6587), .B(n6588), .ZN(n8928) );
  INV_X1 U8127 ( .A(n6587), .ZN(n6589) );
  NAND2_X1 U8128 ( .A1(n6589), .A2(n6588), .ZN(n6590) );
  NAND2_X1 U8129 ( .A1(n9269), .A2(n6646), .ZN(n6592) );
  NAND2_X1 U8130 ( .A1(n4395), .A2(n9286), .ZN(n6591) );
  NAND2_X1 U8131 ( .A1(n6592), .A2(n6591), .ZN(n6593) );
  NAND2_X1 U8132 ( .A1(n9269), .A2(n4395), .ZN(n6595) );
  NAND2_X1 U8133 ( .A1(n6658), .A2(n9286), .ZN(n6594) );
  NAND2_X1 U8134 ( .A1(n6595), .A2(n6594), .ZN(n8965) );
  NAND2_X1 U8135 ( .A1(n8964), .A2(n8965), .ZN(n8969) );
  INV_X1 U8136 ( .A(n6596), .ZN(n6597) );
  NAND2_X1 U8137 ( .A1(n9388), .A2(n6646), .ZN(n6599) );
  NAND2_X1 U8138 ( .A1(n9237), .A2(n4395), .ZN(n6598) );
  NAND2_X1 U8139 ( .A1(n6599), .A2(n6598), .ZN(n6600) );
  XNOR2_X1 U8140 ( .A(n6600), .B(n7466), .ZN(n8890) );
  NAND2_X1 U8141 ( .A1(n9388), .A2(n4395), .ZN(n6602) );
  NAND2_X1 U8142 ( .A1(n6658), .A2(n9237), .ZN(n6601) );
  NAND2_X1 U8143 ( .A1(n6602), .A2(n6601), .ZN(n8891) );
  NAND2_X1 U8144 ( .A1(n9381), .A2(n6646), .ZN(n6604) );
  NAND2_X1 U8145 ( .A1(n9003), .A2(n4395), .ZN(n6603) );
  NAND2_X1 U8146 ( .A1(n6604), .A2(n6603), .ZN(n6605) );
  XNOR2_X1 U8147 ( .A(n6605), .B(n7466), .ZN(n6608) );
  NAND2_X1 U8148 ( .A1(n9381), .A2(n4395), .ZN(n6607) );
  NAND2_X1 U8149 ( .A1(n9003), .A2(n6658), .ZN(n6606) );
  NAND2_X1 U8150 ( .A1(n6607), .A2(n6606), .ZN(n6609) );
  INV_X1 U8151 ( .A(n6608), .ZN(n6611) );
  INV_X1 U8152 ( .A(n6609), .ZN(n6610) );
  NAND2_X1 U8153 ( .A1(n6611), .A2(n6610), .ZN(n8945) );
  NAND2_X1 U8154 ( .A1(n8942), .A2(n8945), .ZN(n8900) );
  NAND2_X1 U8155 ( .A1(n9378), .A2(n6646), .ZN(n6613) );
  NAND2_X1 U8156 ( .A1(n9236), .A2(n4395), .ZN(n6612) );
  NAND2_X1 U8157 ( .A1(n6613), .A2(n6612), .ZN(n6614) );
  XNOR2_X1 U8158 ( .A(n6614), .B(n7466), .ZN(n6616) );
  AND2_X1 U8159 ( .A1(n9236), .A2(n6658), .ZN(n6615) );
  AOI21_X1 U8160 ( .B1(n9378), .B2(n4395), .A(n6615), .ZN(n6617) );
  XNOR2_X1 U8161 ( .A(n6616), .B(n6617), .ZN(n8901) );
  INV_X1 U8162 ( .A(n6616), .ZN(n6618) );
  NAND2_X1 U8163 ( .A1(n6618), .A2(n6617), .ZN(n6619) );
  AND2_X1 U8164 ( .A1(n9190), .A2(n6658), .ZN(n6620) );
  AOI21_X1 U8165 ( .B1(n9371), .B2(n4395), .A(n6620), .ZN(n6625) );
  NAND2_X1 U8166 ( .A1(n6624), .A2(n6625), .ZN(n8953) );
  NAND2_X1 U8167 ( .A1(n9371), .A2(n6435), .ZN(n6622) );
  NAND2_X1 U8168 ( .A1(n9190), .A2(n4395), .ZN(n6621) );
  NAND2_X1 U8169 ( .A1(n6622), .A2(n6621), .ZN(n6623) );
  XNOR2_X1 U8170 ( .A(n6623), .B(n7466), .ZN(n8954) );
  AND2_X2 U8171 ( .A1(n8953), .A2(n8954), .ZN(n8956) );
  INV_X1 U8172 ( .A(n6631), .ZN(n8952) );
  NAND2_X1 U8173 ( .A1(n9366), .A2(n6646), .ZN(n6627) );
  NAND2_X1 U8174 ( .A1(n9203), .A2(n4395), .ZN(n6626) );
  NAND2_X1 U8175 ( .A1(n6627), .A2(n6626), .ZN(n6628) );
  XNOR2_X1 U8176 ( .A(n6628), .B(n7466), .ZN(n6629) );
  AOI22_X1 U8177 ( .A1(n9366), .A2(n4395), .B1(n6658), .B2(n9203), .ZN(n8883)
         );
  AOI22_X1 U8178 ( .A1(n9363), .A2(n4395), .B1(n6658), .B2(n9183), .ZN(n6636)
         );
  NAND2_X1 U8179 ( .A1(n9363), .A2(n6646), .ZN(n6634) );
  NAND2_X1 U8180 ( .A1(n9183), .A2(n4395), .ZN(n6633) );
  NAND2_X1 U8181 ( .A1(n6634), .A2(n6633), .ZN(n6635) );
  XNOR2_X1 U8182 ( .A(n6635), .B(n7466), .ZN(n6638) );
  XOR2_X1 U8183 ( .A(n6636), .B(n6638), .Z(n8936) );
  INV_X1 U8184 ( .A(n6636), .ZN(n6637) );
  NAND2_X1 U8185 ( .A1(n9356), .A2(n6435), .ZN(n6641) );
  NAND2_X1 U8186 ( .A1(n9166), .A2(n4395), .ZN(n6640) );
  NAND2_X1 U8187 ( .A1(n6641), .A2(n6640), .ZN(n6642) );
  XNOR2_X1 U8188 ( .A(n6642), .B(n7466), .ZN(n6643) );
  AOI22_X1 U8189 ( .A1(n9356), .A2(n4395), .B1(n6658), .B2(n9166), .ZN(n6644)
         );
  XNOR2_X1 U8190 ( .A(n6643), .B(n6644), .ZN(n8909) );
  INV_X1 U8191 ( .A(n6643), .ZN(n6645) );
  NAND2_X1 U8192 ( .A1(n9351), .A2(n6646), .ZN(n6648) );
  NAND2_X1 U8193 ( .A1(n9156), .A2(n4395), .ZN(n6647) );
  NAND2_X1 U8194 ( .A1(n6648), .A2(n6647), .ZN(n6649) );
  XNOR2_X1 U8195 ( .A(n6649), .B(n7466), .ZN(n6651) );
  AND2_X1 U8196 ( .A1(n9156), .A2(n6658), .ZN(n6650) );
  AOI21_X1 U8197 ( .B1(n9351), .B2(n4395), .A(n6650), .ZN(n6652) );
  XNOR2_X1 U8198 ( .A(n6651), .B(n6652), .ZN(n8978) );
  NAND2_X1 U8199 ( .A1(n9346), .A2(n6646), .ZN(n6656) );
  NAND2_X1 U8200 ( .A1(n9142), .A2(n4395), .ZN(n6655) );
  NAND2_X1 U8201 ( .A1(n6656), .A2(n6655), .ZN(n6657) );
  XNOR2_X1 U8202 ( .A(n6657), .B(n7466), .ZN(n8862) );
  AND2_X1 U8203 ( .A1(n9142), .A2(n6658), .ZN(n6659) );
  AOI21_X1 U8204 ( .B1(n9346), .B2(n4395), .A(n6659), .ZN(n8861) );
  INV_X1 U8205 ( .A(n8861), .ZN(n6688) );
  NAND2_X1 U8206 ( .A1(n9341), .A2(n6435), .ZN(n6662) );
  NAND2_X1 U8207 ( .A1(n9002), .A2(n4395), .ZN(n6661) );
  NAND2_X1 U8208 ( .A1(n6662), .A2(n6661), .ZN(n6663) );
  XNOR2_X1 U8209 ( .A(n6663), .B(n6547), .ZN(n6667) );
  NAND2_X1 U8210 ( .A1(n9341), .A2(n6458), .ZN(n6664) );
  OAI21_X1 U8211 ( .B1(n9127), .B2(n6665), .A(n6664), .ZN(n6666) );
  XNOR2_X1 U8212 ( .A(n6667), .B(n6666), .ZN(n6708) );
  INV_X1 U8213 ( .A(n6708), .ZN(n6687) );
  NAND2_X1 U8214 ( .A1(n6434), .A2(n7573), .ZN(n7121) );
  NAND2_X1 U8215 ( .A1(n10032), .A2(n7118), .ZN(n6698) );
  NAND2_X1 U8216 ( .A1(n8013), .A2(P1_B_REG_SCAN_IN), .ZN(n6669) );
  MUX2_X1 U8217 ( .A(P1_B_REG_SCAN_IN), .B(n6669), .S(n7941), .Z(n6671) );
  INV_X1 U8218 ( .A(n8044), .ZN(n6670) );
  INV_X1 U8219 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n9987) );
  NAND2_X1 U8220 ( .A1(n7112), .A2(n9987), .ZN(n6673) );
  NAND2_X1 U8221 ( .A1(n8044), .A2(n8013), .ZN(n6672) );
  NOR4_X1 U8222 ( .A1(P1_D_REG_12__SCAN_IN), .A2(P1_D_REG_13__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_16__SCAN_IN), .ZN(n6677) );
  NOR4_X1 U8223 ( .A1(P1_D_REG_9__SCAN_IN), .A2(P1_D_REG_6__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_10__SCAN_IN), .ZN(n6676) );
  NOR4_X1 U8224 ( .A1(P1_D_REG_25__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_27__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n6675) );
  NOR4_X1 U8225 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_21__SCAN_IN), .A3(
        P1_D_REG_22__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n6674) );
  NAND4_X1 U8226 ( .A1(n6677), .A2(n6676), .A3(n6675), .A4(n6674), .ZN(n6683)
         );
  NOR2_X1 U8227 ( .A1(P1_D_REG_7__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .ZN(
        n6681) );
  NOR4_X1 U8228 ( .A1(P1_D_REG_28__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_14__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n6680) );
  NOR4_X1 U8229 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_5__SCAN_IN), .ZN(n6679) );
  NOR4_X1 U8230 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_18__SCAN_IN), .A3(
        P1_D_REG_23__SCAN_IN), .A4(P1_D_REG_11__SCAN_IN), .ZN(n6678) );
  NAND4_X1 U8231 ( .A1(n6681), .A2(n6680), .A3(n6679), .A4(n6678), .ZN(n6682)
         );
  NOR2_X1 U8232 ( .A1(n6683), .A2(n6682), .ZN(n7110) );
  NAND2_X1 U8233 ( .A1(n7110), .A2(P1_D_REG_0__SCAN_IN), .ZN(n6684) );
  NAND2_X1 U8234 ( .A1(n7112), .A2(n6684), .ZN(n6685) );
  NAND2_X1 U8235 ( .A1(n8044), .A2(n7941), .ZN(n7113) );
  AND2_X1 U8236 ( .A1(n7365), .A2(n7203), .ZN(n6700) );
  AND2_X1 U8237 ( .A1(n6835), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6686) );
  NAND2_X1 U8238 ( .A1(n6700), .A2(n9988), .ZN(n6695) );
  NAND2_X1 U8239 ( .A1(n6687), .A2(n8976), .ZN(n6713) );
  NAND2_X1 U8240 ( .A1(n8862), .A2(n6688), .ZN(n6707) );
  INV_X1 U8241 ( .A(n6707), .ZN(n6689) );
  NOR2_X1 U8242 ( .A1(n6689), .A2(n8999), .ZN(n6690) );
  AND2_X1 U8243 ( .A1(n6708), .A2(n6690), .ZN(n6691) );
  NAND2_X1 U8244 ( .A1(n6714), .A2(n6691), .ZN(n6712) );
  NAND2_X1 U8245 ( .A1(n9988), .A2(n9250), .ZN(n6692) );
  OR2_X1 U8246 ( .A1(n7121), .A2(n7494), .ZN(n7370) );
  OR2_X1 U8247 ( .A1(n7370), .A2(n6695), .ZN(n6693) );
  OR2_X1 U8248 ( .A1(n7372), .A2(n6694), .ZN(n7467) );
  NOR2_X1 U8249 ( .A1(n7467), .A2(n6695), .ZN(n6696) );
  INV_X1 U8250 ( .A(n4393), .ZN(n7117) );
  INV_X1 U8251 ( .A(n6696), .ZN(n6697) );
  AOI22_X1 U8252 ( .A1(n9105), .A2(n8991), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3084), .ZN(n6705) );
  OAI21_X1 U8253 ( .B1(n6698), .B2(n6700), .A(n7042), .ZN(n6699) );
  NAND2_X1 U8254 ( .A1(n6699), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6703) );
  NAND2_X1 U8255 ( .A1(n7370), .A2(n7467), .ZN(n6702) );
  INV_X1 U8256 ( .A(n6700), .ZN(n7045) );
  AND2_X1 U8257 ( .A1(n7045), .A2(n9988), .ZN(n6701) );
  NAND2_X1 U8258 ( .A1(n6702), .A2(n6701), .ZN(n7043) );
  NAND2_X1 U8259 ( .A1(n9111), .A2(n8992), .ZN(n6704) );
  OAI211_X1 U8260 ( .C1(n6706), .C2(n8995), .A(n6705), .B(n6704), .ZN(n6710)
         );
  NOR3_X1 U8261 ( .A1(n6708), .A2(n8999), .A3(n6707), .ZN(n6709) );
  AOI211_X1 U8262 ( .C1(n9341), .C2(n8997), .A(n6710), .B(n6709), .ZN(n6711)
         );
  OAI211_X1 U8263 ( .C1(n6714), .C2(n6713), .A(n6712), .B(n6711), .ZN(P1_U3218) );
  NOR2_X1 U8264 ( .A1(n6834), .A2(n6715), .ZN(n6860) );
  OR2_X1 U8265 ( .A1(n6824), .A2(P2_U3152), .ZN(n6925) );
  INV_X2 U8266 ( .A(n8340), .ZN(P2_U3966) );
  NAND2_X1 U8267 ( .A1(n6726), .A2(n6718), .ZN(n6721) );
  XNOR2_X1 U8268 ( .A(n6720), .B(n6721), .ZN(n7263) );
  NAND2_X1 U8269 ( .A1(n5990), .A2(n7792), .ZN(n7236) );
  INV_X1 U8270 ( .A(n7236), .ZN(n7768) );
  NAND2_X1 U8271 ( .A1(n6726), .A2(n7768), .ZN(n7172) );
  OR2_X1 U8272 ( .A1(n6724), .A2(n7792), .ZN(n6719) );
  AND2_X1 U8273 ( .A1(n7172), .A2(n6719), .ZN(n7264) );
  NAND2_X1 U8274 ( .A1(n7263), .A2(n7264), .ZN(n7262) );
  INV_X1 U8275 ( .A(n6720), .ZN(n6722) );
  NAND2_X1 U8276 ( .A1(n6722), .A2(n6721), .ZN(n6723) );
  NAND2_X1 U8277 ( .A1(n7262), .A2(n6723), .ZN(n7256) );
  INV_X1 U8278 ( .A(n10136), .ZN(n7902) );
  XNOR2_X1 U8279 ( .A(n6724), .B(n7902), .ZN(n6727) );
  AND2_X1 U8280 ( .A1(n6726), .A2(n6725), .ZN(n6728) );
  NAND2_X1 U8281 ( .A1(n6727), .A2(n6728), .ZN(n6731) );
  INV_X1 U8282 ( .A(n6727), .ZN(n7277) );
  INV_X1 U8283 ( .A(n6728), .ZN(n6729) );
  NAND2_X1 U8284 ( .A1(n7277), .A2(n6729), .ZN(n6730) );
  NAND2_X1 U8285 ( .A1(n6731), .A2(n6730), .ZN(n7255) );
  INV_X1 U8286 ( .A(n10141), .ZN(n7762) );
  XNOR2_X1 U8287 ( .A(n6724), .B(n7762), .ZN(n6734) );
  NAND2_X1 U8288 ( .A1(n8212), .A2(n8352), .ZN(n6732) );
  XNOR2_X1 U8289 ( .A(n6734), .B(n6732), .ZN(n7274) );
  INV_X1 U8290 ( .A(n6732), .ZN(n6733) );
  NAND2_X1 U8291 ( .A1(n6734), .A2(n6733), .ZN(n6735) );
  XNOR2_X1 U8292 ( .A(n6724), .B(n10103), .ZN(n7291) );
  AND2_X1 U8293 ( .A1(n8212), .A2(n8351), .ZN(n6736) );
  AND2_X1 U8294 ( .A1(n7291), .A2(n6736), .ZN(n7283) );
  INV_X1 U8295 ( .A(n7291), .ZN(n6738) );
  INV_X1 U8296 ( .A(n6736), .ZN(n6737) );
  NAND2_X1 U8297 ( .A1(n6738), .A2(n6737), .ZN(n7285) );
  XNOR2_X1 U8298 ( .A(n6724), .B(n6740), .ZN(n6741) );
  NAND2_X1 U8299 ( .A1(n8212), .A2(n8350), .ZN(n6742) );
  XNOR2_X1 U8300 ( .A(n6741), .B(n6742), .ZN(n7315) );
  INV_X1 U8301 ( .A(n6741), .ZN(n6744) );
  INV_X1 U8302 ( .A(n6742), .ZN(n6743) );
  XNOR2_X1 U8303 ( .A(n6724), .B(n10151), .ZN(n6745) );
  NAND2_X1 U8304 ( .A1(n8212), .A2(n8349), .ZN(n6746) );
  NAND2_X1 U8305 ( .A1(n6745), .A2(n6746), .ZN(n6750) );
  INV_X1 U8306 ( .A(n6745), .ZN(n6748) );
  INV_X1 U8307 ( .A(n6746), .ZN(n6747) );
  NAND2_X1 U8308 ( .A1(n6748), .A2(n6747), .ZN(n6749) );
  AND2_X1 U8309 ( .A1(n6750), .A2(n6749), .ZN(n8301) );
  NAND2_X1 U8310 ( .A1(n8300), .A2(n8301), .ZN(n8299) );
  XNOR2_X1 U8311 ( .A(n6724), .B(n10157), .ZN(n6751) );
  NAND2_X1 U8312 ( .A1(n8212), .A2(n8348), .ZN(n6752) );
  XNOR2_X1 U8313 ( .A(n6751), .B(n6752), .ZN(n7487) );
  INV_X1 U8314 ( .A(n6751), .ZN(n6754) );
  INV_X1 U8315 ( .A(n6752), .ZN(n6753) );
  NAND2_X1 U8316 ( .A1(n6754), .A2(n6753), .ZN(n6755) );
  XNOR2_X1 U8317 ( .A(n6724), .B(n7698), .ZN(n6758) );
  NAND2_X1 U8318 ( .A1(n8212), .A2(n8347), .ZN(n6756) );
  XNOR2_X1 U8319 ( .A(n6758), .B(n6756), .ZN(n7654) );
  INV_X1 U8320 ( .A(n6756), .ZN(n6757) );
  AND2_X1 U8321 ( .A1(n6758), .A2(n6757), .ZN(n6759) );
  INV_X1 U8322 ( .A(n7805), .ZN(n10171) );
  XNOR2_X1 U8323 ( .A(n6724), .B(n10171), .ZN(n6760) );
  INV_X1 U8324 ( .A(n7834), .ZN(n8346) );
  NAND2_X1 U8325 ( .A1(n8212), .A2(n8346), .ZN(n6761) );
  NAND2_X1 U8326 ( .A1(n6760), .A2(n6761), .ZN(n6765) );
  INV_X1 U8327 ( .A(n6760), .ZN(n6763) );
  INV_X1 U8328 ( .A(n6761), .ZN(n6762) );
  NAND2_X1 U8329 ( .A1(n6763), .A2(n6762), .ZN(n6764) );
  AND2_X1 U8330 ( .A1(n6765), .A2(n6764), .ZN(n7821) );
  XNOR2_X1 U8331 ( .A(n10178), .B(n6724), .ZN(n6767) );
  INV_X1 U8332 ( .A(n7947), .ZN(n8345) );
  AND2_X1 U8333 ( .A1(n8212), .A2(n8345), .ZN(n6766) );
  XNOR2_X1 U8334 ( .A(n6767), .B(n6766), .ZN(n7830) );
  NAND2_X1 U8335 ( .A1(n6767), .A2(n6766), .ZN(n6768) );
  XNOR2_X1 U8336 ( .A(n7950), .B(n6724), .ZN(n6771) );
  INV_X1 U8337 ( .A(n8020), .ZN(n8344) );
  NAND2_X1 U8338 ( .A1(n8212), .A2(n8344), .ZN(n6769) );
  XNOR2_X1 U8339 ( .A(n6771), .B(n6769), .ZN(n7943) );
  INV_X1 U8340 ( .A(n6769), .ZN(n6770) );
  XNOR2_X1 U8341 ( .A(n8023), .B(n6739), .ZN(n6772) );
  INV_X1 U8342 ( .A(n8049), .ZN(n8343) );
  NAND2_X1 U8343 ( .A1(n6726), .A2(n8343), .ZN(n6773) );
  NAND2_X1 U8344 ( .A1(n6772), .A2(n6773), .ZN(n8015) );
  INV_X1 U8345 ( .A(n6772), .ZN(n6775) );
  INV_X1 U8346 ( .A(n6773), .ZN(n6774) );
  NAND2_X1 U8347 ( .A1(n6775), .A2(n6774), .ZN(n8016) );
  NAND2_X1 U8348 ( .A1(n6776), .A2(n8016), .ZN(n8046) );
  XNOR2_X1 U8349 ( .A(n8026), .B(n6724), .ZN(n6777) );
  INV_X1 U8350 ( .A(n8179), .ZN(n8342) );
  AND2_X1 U8351 ( .A1(n8212), .A2(n8342), .ZN(n6778) );
  NAND2_X1 U8352 ( .A1(n6777), .A2(n6778), .ZN(n6781) );
  INV_X1 U8353 ( .A(n6777), .ZN(n8173) );
  INV_X1 U8354 ( .A(n6778), .ZN(n6779) );
  NAND2_X1 U8355 ( .A1(n8173), .A2(n6779), .ZN(n6780) );
  AND2_X1 U8356 ( .A1(n6781), .A2(n6780), .ZN(n8047) );
  XNOR2_X1 U8357 ( .A(n8475), .B(n6724), .ZN(n6783) );
  NAND2_X1 U8358 ( .A1(n6726), .A2(n8474), .ZN(n6784) );
  XNOR2_X1 U8359 ( .A(n6783), .B(n6784), .ZN(n8185) );
  AND2_X1 U8360 ( .A1(n8185), .A2(n6781), .ZN(n6782) );
  INV_X1 U8361 ( .A(n6783), .ZN(n6785) );
  NAND2_X1 U8362 ( .A1(n6785), .A2(n6784), .ZN(n6786) );
  XNOR2_X1 U8363 ( .A(n8825), .B(n6724), .ZN(n8252) );
  INV_X1 U8364 ( .A(n8737), .ZN(n8479) );
  AND2_X1 U8365 ( .A1(n6726), .A2(n8479), .ZN(n6789) );
  INV_X1 U8366 ( .A(n8719), .ZN(n8477) );
  AND2_X1 U8367 ( .A1(n8212), .A2(n8477), .ZN(n6788) );
  XNOR2_X1 U8368 ( .A(n8745), .B(n6724), .ZN(n8248) );
  AOI22_X1 U8369 ( .A1(n8252), .A2(n6789), .B1(n6788), .B2(n8248), .ZN(n6787)
         );
  INV_X1 U8370 ( .A(n8252), .ZN(n6791) );
  OAI21_X1 U8371 ( .B1(n8248), .B2(n6788), .A(n6789), .ZN(n6790) );
  INV_X1 U8372 ( .A(n8248), .ZN(n8250) );
  INV_X1 U8373 ( .A(n6788), .ZN(n8324) );
  INV_X1 U8374 ( .A(n6789), .ZN(n8251) );
  AOI21_X1 U8375 ( .B1(n6791), .B2(n6790), .A(n4957), .ZN(n6792) );
  XNOR2_X1 U8376 ( .A(n8822), .B(n6724), .ZN(n6793) );
  INV_X1 U8377 ( .A(n8718), .ZN(n8685) );
  AND2_X1 U8378 ( .A1(n8212), .A2(n8685), .ZN(n6794) );
  NAND2_X1 U8379 ( .A1(n6793), .A2(n6794), .ZN(n8125) );
  INV_X1 U8380 ( .A(n6793), .ZN(n8292) );
  INV_X1 U8381 ( .A(n6794), .ZN(n6795) );
  NAND2_X1 U8382 ( .A1(n8292), .A2(n6795), .ZN(n6796) );
  NAND2_X1 U8383 ( .A1(n8125), .A2(n6796), .ZN(n6816) );
  INV_X1 U8384 ( .A(n8042), .ZN(n6799) );
  XNOR2_X1 U8385 ( .A(n7939), .B(P2_B_REG_SCAN_IN), .ZN(n6797) );
  NAND2_X1 U8386 ( .A1(n8011), .A2(n6797), .ZN(n6798) );
  INV_X1 U8387 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n10118) );
  AND2_X1 U8388 ( .A1(n8011), .A2(n8042), .ZN(n10120) );
  AOI21_X1 U8389 ( .B1(n10109), .B2(n10118), .A(n10120), .ZN(n7676) );
  NOR4_X1 U8390 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_16__SCAN_IN), .A3(
        P2_D_REG_17__SCAN_IN), .A4(P2_D_REG_19__SCAN_IN), .ZN(n6803) );
  NOR4_X1 U8391 ( .A1(P2_D_REG_13__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), .A3(
        P2_D_REG_12__SCAN_IN), .A4(P2_D_REG_14__SCAN_IN), .ZN(n6802) );
  NOR4_X1 U8392 ( .A1(P2_D_REG_25__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_27__SCAN_IN), .A4(P2_D_REG_30__SCAN_IN), .ZN(n6801) );
  NOR4_X1 U8393 ( .A1(P2_D_REG_21__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .A3(
        P2_D_REG_23__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n6800) );
  NAND4_X1 U8394 ( .A1(n6803), .A2(n6802), .A3(n6801), .A4(n6800), .ZN(n6809)
         );
  NOR2_X1 U8395 ( .A1(P2_D_REG_31__SCAN_IN), .A2(P2_D_REG_18__SCAN_IN), .ZN(
        n6807) );
  NOR4_X1 U8396 ( .A1(P2_D_REG_28__SCAN_IN), .A2(P2_D_REG_29__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n6806) );
  NOR4_X1 U8397 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_8__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_10__SCAN_IN), .ZN(n6805) );
  NOR4_X1 U8398 ( .A1(P2_D_REG_3__SCAN_IN), .A2(P2_D_REG_4__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_6__SCAN_IN), .ZN(n6804) );
  NAND4_X1 U8399 ( .A1(n6807), .A2(n6806), .A3(n6805), .A4(n6804), .ZN(n6808)
         );
  OAI21_X1 U8400 ( .B1(n6809), .B2(n6808), .A(n10109), .ZN(n7675) );
  INV_X1 U8401 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n10115) );
  NAND2_X1 U8402 ( .A1(n10109), .A2(n10115), .ZN(n6811) );
  AND2_X1 U8403 ( .A1(n7939), .A2(n8042), .ZN(n10116) );
  INV_X1 U8404 ( .A(n10116), .ZN(n6810) );
  NAND2_X1 U8405 ( .A1(n6811), .A2(n6810), .ZN(n7674) );
  INV_X1 U8406 ( .A(n7674), .ZN(n7232) );
  AND2_X1 U8407 ( .A1(n7675), .A2(n7232), .ZN(n6812) );
  NAND2_X1 U8408 ( .A1(n7676), .A2(n6812), .ZN(n6821) );
  NOR2_X1 U8409 ( .A1(n6821), .A2(n10110), .ZN(n6829) );
  INV_X1 U8410 ( .A(n6927), .ZN(n7233) );
  AND2_X1 U8411 ( .A1(n10192), .A2(n7233), .ZN(n6813) );
  INV_X1 U8412 ( .A(n6816), .ZN(n6814) );
  INV_X1 U8413 ( .A(n8290), .ZN(n6815) );
  AOI211_X1 U8414 ( .C1(n6817), .C2(n6816), .A(n8321), .B(n6815), .ZN(n6833)
         );
  INV_X1 U8415 ( .A(n8822), .ZN(n8704) );
  NOR2_X1 U8416 ( .A1(n8059), .A2(n10123), .ZN(n7688) );
  NAND2_X1 U8417 ( .A1(n6829), .A2(n7688), .ZN(n6820) );
  INV_X1 U8418 ( .A(n8319), .ZN(n8337) );
  NOR2_X1 U8419 ( .A1(n8704), .A2(n8337), .ZN(n6832) );
  NAND2_X1 U8420 ( .A1(n6821), .A2(n7229), .ZN(n6826) );
  INV_X1 U8421 ( .A(n6822), .ZN(n6823) );
  NAND2_X1 U8422 ( .A1(n6824), .A2(n6823), .ZN(n6825) );
  AOI21_X1 U8423 ( .B1(n6410), .B2(n6927), .A(n6825), .ZN(n7679) );
  NAND2_X1 U8424 ( .A1(n6826), .A2(n7679), .ZN(n6827) );
  OAI22_X1 U8425 ( .A1(n8317), .A2(n8705), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6163), .ZN(n6831) );
  INV_X1 U8426 ( .A(n6410), .ZN(n6828) );
  NAND2_X1 U8427 ( .A1(n8315), .A2(n8686), .ZN(n8331) );
  NAND2_X1 U8428 ( .A1(n8315), .A2(n8684), .ZN(n8330) );
  OAI22_X1 U8429 ( .A1(n8698), .A2(n8331), .B1(n8330), .B2(n8737), .ZN(n6830)
         );
  OR4_X1 U8430 ( .A1(n6833), .A2(n6832), .A3(n6831), .A4(n6830), .ZN(P2_U3230)
         );
  NAND2_X1 U8431 ( .A1(n7118), .A2(n6834), .ZN(n6836) );
  NAND2_X1 U8432 ( .A1(n6836), .A2(n6835), .ZN(n7006) );
  NAND2_X1 U8433 ( .A1(n7006), .A2(n5388), .ZN(n6837) );
  NAND2_X1 U8434 ( .A1(n6837), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U3083) );
  NOR2_X1 U8435 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n9566), .ZN(n7443) );
  AND2_X1 U8436 ( .A1(n8056), .A2(n7117), .ZN(n6838) );
  INV_X1 U8437 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n6843) );
  INV_X1 U8438 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n7427) );
  INV_X1 U8439 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n6842) );
  INV_X1 U8440 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n6841) );
  INV_X1 U8441 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n6839) );
  MUX2_X1 U8442 ( .A(n6839), .B(P1_REG2_REG_1__SCAN_IN), .S(n6885), .Z(n9022)
         );
  AND2_X1 U8443 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n9021) );
  NAND2_X1 U8444 ( .A1(n9022), .A2(n9021), .ZN(n9020) );
  INV_X1 U8445 ( .A(n6885), .ZN(n9019) );
  NAND2_X1 U8446 ( .A1(n9019), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6840) );
  NAND2_X1 U8447 ( .A1(n9020), .A2(n6840), .ZN(n6877) );
  OAI21_X1 U8448 ( .B1(n6887), .B2(n6841), .A(n6876), .ZN(n7054) );
  XNOR2_X1 U8449 ( .A(n6888), .B(P1_REG2_REG_3__SCAN_IN), .ZN(n7055) );
  NAND2_X1 U8450 ( .A1(n7054), .A2(n7055), .ZN(n7053) );
  OAI21_X1 U8451 ( .B1(n6888), .B2(n6842), .A(n7053), .ZN(n9882) );
  MUX2_X1 U8452 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n7427), .S(n9884), .Z(n9883)
         );
  NOR2_X1 U8453 ( .A1(n9882), .A2(n9883), .ZN(n9881) );
  AOI21_X1 U8454 ( .B1(n9884), .B2(n7427), .A(n9881), .ZN(n7065) );
  XOR2_X1 U8455 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n7062), .Z(n7064) );
  NOR2_X1 U8456 ( .A1(n7065), .A2(n7064), .ZN(n7063) );
  AOI21_X1 U8457 ( .B1(n6843), .B2(n7062), .A(n7063), .ZN(n6846) );
  INV_X1 U8458 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n6844) );
  MUX2_X1 U8459 ( .A(n6844), .B(P1_REG2_REG_6__SCAN_IN), .S(n7031), .Z(n6845)
         );
  NOR2_X1 U8460 ( .A1(n6846), .A2(n6845), .ZN(n6847) );
  NOR3_X1 U8461 ( .A1(n9886), .A2(n7032), .A3(n6847), .ZN(n6864) );
  OR2_X1 U8462 ( .A1(n4393), .A2(P1_U3084), .ZN(n9450) );
  INV_X1 U8463 ( .A(n4394), .ZN(n6868) );
  NOR2_X1 U8464 ( .A1(n9450), .A2(n6868), .ZN(n6848) );
  NAND2_X1 U8465 ( .A1(n7006), .A2(n6848), .ZN(n9902) );
  INV_X1 U8466 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n10045) );
  MUX2_X1 U8467 ( .A(n10045), .B(P1_REG1_REG_2__SCAN_IN), .S(n6887), .Z(n6875)
         );
  INV_X1 U8468 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n10043) );
  MUX2_X1 U8469 ( .A(n10043), .B(P1_REG1_REG_1__SCAN_IN), .S(n6885), .Z(n9025)
         );
  AND2_X1 U8470 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n9024) );
  NAND2_X1 U8471 ( .A1(n9025), .A2(n9024), .ZN(n9023) );
  NAND2_X1 U8472 ( .A1(n9019), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6849) );
  NAND2_X1 U8473 ( .A1(n9023), .A2(n6849), .ZN(n6874) );
  NAND2_X1 U8474 ( .A1(n6875), .A2(n6874), .ZN(n6873) );
  INV_X1 U8475 ( .A(n6887), .ZN(n6850) );
  NAND2_X1 U8476 ( .A1(n6850), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6851) );
  NAND2_X1 U8477 ( .A1(n6873), .A2(n6851), .ZN(n7051) );
  XNOR2_X1 U8478 ( .A(n6888), .B(P1_REG1_REG_3__SCAN_IN), .ZN(n7052) );
  NAND2_X1 U8479 ( .A1(n7051), .A2(n7052), .ZN(n7050) );
  INV_X1 U8480 ( .A(n6888), .ZN(n7059) );
  NAND2_X1 U8481 ( .A1(n7059), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6852) );
  NAND2_X1 U8482 ( .A1(n7050), .A2(n6852), .ZN(n9889) );
  INV_X1 U8483 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n10049) );
  MUX2_X1 U8484 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n10049), .S(n9884), .Z(n9888)
         );
  OR2_X1 U8485 ( .A1(n9889), .A2(n9888), .ZN(n9891) );
  NAND2_X1 U8486 ( .A1(n9884), .A2(n10049), .ZN(n6853) );
  AND2_X1 U8487 ( .A1(n9891), .A2(n6853), .ZN(n7067) );
  XNOR2_X1 U8488 ( .A(n7062), .B(P1_REG1_REG_5__SCAN_IN), .ZN(n7068) );
  NAND2_X1 U8489 ( .A1(n7067), .A2(n7068), .ZN(n7066) );
  INV_X1 U8490 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n6854) );
  OR2_X1 U8491 ( .A1(n7062), .A2(n6854), .ZN(n6855) );
  AND2_X1 U8492 ( .A1(n7066), .A2(n6855), .ZN(n6858) );
  INV_X1 U8493 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n6856) );
  MUX2_X1 U8494 ( .A(n6856), .B(P1_REG1_REG_6__SCAN_IN), .S(n7031), .Z(n6857)
         );
  NAND2_X1 U8495 ( .A1(n6858), .A2(n6857), .ZN(n7033) );
  OAI21_X1 U8496 ( .B1(n6858), .B2(n6857), .A(n7033), .ZN(n6859) );
  AND2_X1 U8497 ( .A1(n9938), .A2(n6859), .ZN(n6863) );
  INV_X1 U8498 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n9623) );
  AND2_X1 U8499 ( .A1(n8056), .A2(n4393), .ZN(n6861) );
  NAND2_X1 U8500 ( .A1(n7006), .A2(n6861), .ZN(n9922) );
  OAI22_X1 U8501 ( .A1(n9945), .A2(n9623), .B1(n7031), .B2(n9922), .ZN(n6862)
         );
  OR4_X1 U8502 ( .A1(n7443), .A2(n6864), .A3(n6863), .A4(n6862), .ZN(P1_U3247)
         );
  OAI21_X1 U8503 ( .B1(n6867), .B2(n6866), .A(n6865), .ZN(n7046) );
  MUX2_X1 U8504 ( .A(n7046), .B(n4528), .S(n6868), .Z(n6870) );
  NOR2_X1 U8505 ( .A1(n4394), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n6869) );
  NOR2_X1 U8506 ( .A1(n6869), .A2(n4393), .ZN(n7002) );
  MUX2_X1 U8507 ( .A(P1_IR_REG_0__SCAN_IN), .B(n6870), .S(n7002), .Z(n6871) );
  NAND2_X1 U8508 ( .A1(n6871), .A2(P1_U4006), .ZN(n9895) );
  INV_X1 U8509 ( .A(n9895), .ZN(n6884) );
  INV_X1 U8510 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n6872) );
  NOR2_X1 U8511 ( .A1(n9945), .A2(n6872), .ZN(n6883) );
  INV_X1 U8512 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n7156) );
  OAI22_X1 U8513 ( .A1(n9922), .A2(n6887), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n7156), .ZN(n6882) );
  OAI21_X1 U8514 ( .B1(n6875), .B2(n6874), .A(n6873), .ZN(n6880) );
  OAI211_X1 U8515 ( .C1(n6878), .C2(n6877), .A(n9941), .B(n6876), .ZN(n6879)
         );
  OAI21_X1 U8516 ( .B1(n9902), .B2(n6880), .A(n6879), .ZN(n6881) );
  OR4_X1 U8517 ( .A1(n6884), .A2(n6883), .A3(n6882), .A4(n6881), .ZN(P1_U3243)
         );
  NOR2_X1 U8518 ( .A1(n4975), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9730) );
  INV_X1 U8519 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6886) );
  NAND2_X1 U8520 ( .A1(n4975), .A2(P1_U3084), .ZN(n9452) );
  OAI222_X1 U8521 ( .A1(n9449), .A2(n6886), .B1(n9452), .B2(n6894), .C1(
        P1_U3084), .C2(n6885), .ZN(P1_U3352) );
  OAI222_X1 U8522 ( .A1(n9449), .A2(n4973), .B1(n9452), .B2(n6893), .C1(
        P1_U3084), .C2(n6887), .ZN(P1_U3351) );
  OAI222_X1 U8523 ( .A1(n9449), .A2(n4694), .B1(n9452), .B2(n6892), .C1(
        P1_U3084), .C2(n6888), .ZN(P1_U3350) );
  OAI222_X1 U8524 ( .A1(n9449), .A2(n9713), .B1(n9452), .B2(n6895), .C1(
        P1_U3084), .C2(n9884), .ZN(P1_U3349) );
  INV_X1 U8525 ( .A(n9452), .ZN(n9732) );
  INV_X1 U8526 ( .A(n9732), .ZN(n9445) );
  OAI222_X1 U8527 ( .A1(n9449), .A2(n6889), .B1(n9445), .B2(n6897), .C1(
        P1_U3084), .C2(n7062), .ZN(P1_U3348) );
  OAI222_X1 U8528 ( .A1(n9449), .A2(n6890), .B1(n9452), .B2(n6899), .C1(
        P1_U3084), .C2(n7031), .ZN(P1_U3347) );
  AND2_X1 U8529 ( .A1(n6891), .A2(P2_U3152), .ZN(n8856) );
  INV_X1 U8530 ( .A(n8856), .ZN(n8124) );
  INV_X1 U8531 ( .A(n6950), .ZN(n6980) );
  OAI222_X1 U8532 ( .A1(n8124), .A2(n4980), .B1(n8859), .B2(n6892), .C1(
        P2_U3152), .C2(n6980), .ZN(P2_U3355) );
  OAI222_X1 U8533 ( .A1(n8124), .A2(n4974), .B1(n8859), .B2(n6893), .C1(
        P2_U3152), .C2(n6005), .ZN(P2_U3356) );
  INV_X1 U8534 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n9710) );
  OAI222_X1 U8535 ( .A1(n8124), .A2(n9710), .B1(n8859), .B2(n6894), .C1(
        P2_U3152), .C2(n6954), .ZN(P2_U3357) );
  INV_X1 U8536 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6896) );
  INV_X1 U8537 ( .A(n6957), .ZN(n6990) );
  OAI222_X1 U8538 ( .A1(n8124), .A2(n6896), .B1(n8859), .B2(n6895), .C1(
        P2_U3152), .C2(n6990), .ZN(P2_U3354) );
  OAI222_X1 U8539 ( .A1(n8124), .A2(n6898), .B1(n8859), .B2(n6897), .C1(
        P2_U3152), .C2(n6958), .ZN(P2_U3353) );
  OAI222_X1 U8540 ( .A1(n8124), .A2(n9581), .B1(n8859), .B2(n6899), .C1(
        P2_U3152), .C2(n6959), .ZN(P2_U3352) );
  INV_X1 U8541 ( .A(n7112), .ZN(n6900) );
  AND2_X1 U8542 ( .A1(n9988), .A2(n6900), .ZN(n9984) );
  INV_X1 U8543 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n7109) );
  NAND2_X1 U8544 ( .A1(n9984), .A2(n7113), .ZN(n6901) );
  OAI21_X1 U8545 ( .B1(n9984), .B2(n7109), .A(n6901), .ZN(P1_U3440) );
  INV_X1 U8546 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6903) );
  INV_X1 U8547 ( .A(n6902), .ZN(n6904) );
  INV_X1 U8548 ( .A(n6946), .ZN(n7001) );
  OAI222_X1 U8549 ( .A1(n8124), .A2(n6903), .B1(n8859), .B2(n6904), .C1(
        P2_U3152), .C2(n7001), .ZN(P2_U3351) );
  INV_X1 U8550 ( .A(n7092), .ZN(n7079) );
  OAI222_X1 U8551 ( .A1(n9449), .A2(n9712), .B1(n9452), .B2(n6904), .C1(
        P1_U3084), .C2(n7079), .ZN(P1_U3346) );
  INV_X1 U8552 ( .A(n6905), .ZN(n6907) );
  INV_X1 U8553 ( .A(n7022), .ZN(n6969) );
  OAI222_X1 U8554 ( .A1(n8124), .A2(n6906), .B1(n8859), .B2(n6907), .C1(
        P2_U3152), .C2(n6969), .ZN(P2_U3350) );
  INV_X1 U8555 ( .A(n7090), .ZN(n9906) );
  OAI222_X1 U8556 ( .A1(n9449), .A2(n6908), .B1(n9452), .B2(n6907), .C1(
        P1_U3084), .C2(n9906), .ZN(P1_U3345) );
  INV_X1 U8557 ( .A(n6909), .ZN(n6911) );
  INV_X1 U8558 ( .A(n7095), .ZN(n9921) );
  OAI222_X1 U8559 ( .A1(n9445), .A2(n6911), .B1(n9921), .B2(P1_U3084), .C1(
        n6910), .C2(n9449), .ZN(P1_U3344) );
  INV_X1 U8560 ( .A(n7141), .ZN(n7030) );
  OAI222_X1 U8561 ( .A1(n8124), .A2(n6912), .B1(n8859), .B2(n6911), .C1(n7030), 
        .C2(P2_U3152), .ZN(P2_U3349) );
  OAI21_X1 U8562 ( .B1(n10110), .B2(n7233), .A(n6928), .ZN(n6914) );
  NAND2_X1 U8563 ( .A1(n10110), .A2(n6926), .ZN(n6913) );
  NAND2_X1 U8564 ( .A1(n6914), .A2(n6913), .ZN(n8460) );
  NOR2_X1 U8565 ( .A1(n10058), .A2(P2_U3966), .ZN(P2_U3151) );
  INV_X1 U8566 ( .A(n6915), .ZN(n6917) );
  INV_X1 U8567 ( .A(n7219), .ZN(n7085) );
  OAI222_X1 U8568 ( .A1(n9445), .A2(n6917), .B1(n7085), .B2(P1_U3084), .C1(
        n6916), .C2(n9449), .ZN(P1_U3343) );
  INV_X1 U8569 ( .A(n7184), .ZN(n7149) );
  OAI222_X1 U8570 ( .A1(n8124), .A2(n6918), .B1(n8859), .B2(n6917), .C1(n7149), 
        .C2(P2_U3152), .ZN(P2_U3348) );
  INV_X1 U8571 ( .A(n6919), .ZN(n6924) );
  INV_X1 U8572 ( .A(n9930), .ZN(n7217) );
  OAI222_X1 U8573 ( .A1(n9445), .A2(n6924), .B1(n7217), .B2(P1_U3084), .C1(
        n6920), .C2(n9449), .ZN(P1_U3342) );
  INV_X1 U8574 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n6923) );
  INV_X1 U8575 ( .A(n6921), .ZN(n8466) );
  NAND2_X1 U8576 ( .A1(n8466), .A2(P2_U3966), .ZN(n6922) );
  OAI21_X1 U8577 ( .B1(P2_U3966), .B2(n6923), .A(n6922), .ZN(P2_U3583) );
  INV_X1 U8578 ( .A(n7339), .ZN(n7334) );
  OAI222_X1 U8579 ( .A1(P2_U3152), .A2(n7334), .B1(n8859), .B2(n6924), .C1(
        n9644), .C2(n8124), .ZN(P2_U3347) );
  OAI211_X1 U8580 ( .C1(n10110), .C2(n6927), .A(n6926), .B(n6925), .ZN(n6929)
         );
  NAND2_X1 U8581 ( .A1(n6929), .A2(n6928), .ZN(n6940) );
  NAND2_X1 U8582 ( .A1(n8340), .A2(n6940), .ZN(n6963) );
  AND2_X1 U8583 ( .A1(n6963), .A2(n6930), .ZN(n9753) );
  INV_X1 U8584 ( .A(n9753), .ZN(n10059) );
  NAND2_X1 U8585 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3152), .ZN(n7656) );
  INV_X1 U8586 ( .A(n7656), .ZN(n6945) );
  MUX2_X1 U8587 ( .A(n5955), .B(P2_REG1_REG_6__SCAN_IN), .S(n6959), .Z(n8374)
         );
  XNOR2_X1 U8588 ( .A(n6958), .B(P2_REG1_REG_5__SCAN_IN), .ZN(n8361) );
  NAND2_X1 U8589 ( .A1(n6957), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n6936) );
  INV_X1 U8590 ( .A(n6954), .ZN(n9741) );
  NAND2_X1 U8591 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n9739) );
  INV_X1 U8592 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n6931) );
  MUX2_X1 U8593 ( .A(P2_REG1_REG_1__SCAN_IN), .B(n6931), .S(n6954), .Z(n9738)
         );
  NOR2_X1 U8594 ( .A1(n9739), .A2(n9738), .ZN(n9737) );
  AOI21_X1 U8595 ( .B1(n9741), .B2(P2_REG1_REG_1__SCAN_IN), .A(n9737), .ZN(
        n9750) );
  INV_X1 U8596 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n6932) );
  MUX2_X1 U8597 ( .A(n6932), .B(P2_REG1_REG_2__SCAN_IN), .S(n9752), .Z(n9749)
         );
  NAND2_X1 U8598 ( .A1(n6950), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6933) );
  OAI21_X1 U8599 ( .B1(n6950), .B2(P2_REG1_REG_3__SCAN_IN), .A(n6933), .ZN(
        n6971) );
  MUX2_X1 U8600 ( .A(n6934), .B(P2_REG1_REG_4__SCAN_IN), .S(n6957), .Z(n6982)
         );
  NOR2_X1 U8601 ( .A1(n6983), .A2(n6982), .ZN(n6981) );
  INV_X1 U8602 ( .A(n6981), .ZN(n6935) );
  NAND2_X1 U8603 ( .A1(n6936), .A2(n6935), .ZN(n8360) );
  NAND2_X1 U8604 ( .A1(n8361), .A2(n8360), .ZN(n8359) );
  NAND2_X1 U8605 ( .A1(n8358), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6937) );
  NAND2_X1 U8606 ( .A1(n6946), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6938) );
  OAI21_X1 U8607 ( .B1(n6946), .B2(P2_REG1_REG_7__SCAN_IN), .A(n6938), .ZN(
        n6992) );
  AOI21_X1 U8608 ( .B1(n6946), .B2(P2_REG1_REG_7__SCAN_IN), .A(n6991), .ZN(
        n6943) );
  NAND2_X1 U8609 ( .A1(n7022), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n6939) );
  OAI21_X1 U8610 ( .B1(n7022), .B2(P2_REG1_REG_8__SCAN_IN), .A(n6939), .ZN(
        n6942) );
  INV_X1 U8611 ( .A(n6940), .ZN(n6941) );
  AOI211_X1 U8612 ( .C1(n6943), .C2(n6942), .A(n7017), .B(n10060), .ZN(n6944)
         );
  AOI211_X1 U8613 ( .C1(n10058), .C2(P2_ADDR_REG_8__SCAN_IN), .A(n6945), .B(
        n6944), .ZN(n6968) );
  NAND2_X1 U8614 ( .A1(n6946), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n6960) );
  MUX2_X1 U8615 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n6947), .S(n6946), .Z(n6997)
         );
  MUX2_X1 U8616 ( .A(n6948), .B(P2_REG2_REG_6__SCAN_IN), .S(n6959), .Z(n8367)
         );
  MUX2_X1 U8617 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n7780), .S(n6958), .Z(n8354)
         );
  MUX2_X1 U8618 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n6949), .S(n6957), .Z(n6986)
         );
  NAND2_X1 U8619 ( .A1(n6950), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n6955) );
  MUX2_X1 U8620 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n6951), .S(n6950), .Z(n6976)
         );
  MUX2_X1 U8621 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n6952), .S(n9752), .Z(n9755)
         );
  MUX2_X1 U8622 ( .A(n6953), .B(P2_REG2_REG_1__SCAN_IN), .S(n6954), .Z(n9743)
         );
  NAND3_X1 U8623 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .A3(n9743), .ZN(n9742) );
  OAI21_X1 U8624 ( .B1(n6954), .B2(n6953), .A(n9742), .ZN(n9756) );
  NAND2_X1 U8625 ( .A1(n9755), .A2(n9756), .ZN(n9754) );
  NAND2_X1 U8626 ( .A1(n6976), .A2(n6977), .ZN(n6975) );
  NAND2_X1 U8627 ( .A1(n6955), .A2(n6975), .ZN(n6987) );
  AOI21_X1 U8628 ( .B1(n6957), .B2(P2_REG2_REG_4__SCAN_IN), .A(n6956), .ZN(
        n8353) );
  OAI21_X1 U8629 ( .B1(n7780), .B2(n6958), .A(n8356), .ZN(n8368) );
  NAND2_X1 U8630 ( .A1(n8367), .A2(n8368), .ZN(n8366) );
  NAND2_X1 U8631 ( .A1(n6997), .A2(n6998), .ZN(n6996) );
  NAND2_X1 U8632 ( .A1(n6960), .A2(n6996), .ZN(n6966) );
  MUX2_X1 U8633 ( .A(n7690), .B(P2_REG2_REG_8__SCAN_IN), .S(n7022), .Z(n6961)
         );
  INV_X1 U8634 ( .A(n6961), .ZN(n6965) );
  INV_X1 U8635 ( .A(n8464), .ZN(n6962) );
  NAND2_X1 U8636 ( .A1(n6963), .A2(n6962), .ZN(n10061) );
  INV_X1 U8637 ( .A(n10061), .ZN(n6964) );
  NAND2_X1 U8638 ( .A1(n6965), .A2(n6966), .ZN(n7023) );
  OAI211_X1 U8639 ( .C1(n6966), .C2(n6965), .A(n10057), .B(n7023), .ZN(n6967)
         );
  OAI211_X1 U8640 ( .C1(n10059), .C2(n6969), .A(n6968), .B(n6967), .ZN(
        P2_U3253) );
  NOR2_X1 U8641 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5928), .ZN(n6974) );
  AOI211_X1 U8642 ( .C1(n6972), .C2(n6971), .A(n6970), .B(n10060), .ZN(n6973)
         );
  AOI211_X1 U8643 ( .C1(n10058), .C2(P2_ADDR_REG_3__SCAN_IN), .A(n6974), .B(
        n6973), .ZN(n6979) );
  OAI211_X1 U8644 ( .C1(n6977), .C2(n6976), .A(n10057), .B(n6975), .ZN(n6978)
         );
  OAI211_X1 U8645 ( .C1(n10059), .C2(n6980), .A(n6979), .B(n6978), .ZN(
        P2_U3248) );
  AND2_X1 U8646 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3152), .ZN(n7290) );
  AOI211_X1 U8647 ( .C1(n6983), .C2(n6982), .A(n6981), .B(n10060), .ZN(n6984)
         );
  AOI211_X1 U8648 ( .C1(n10058), .C2(P2_ADDR_REG_4__SCAN_IN), .A(n7290), .B(
        n6984), .ZN(n6989) );
  OAI211_X1 U8649 ( .C1(n6987), .C2(n6986), .A(n10057), .B(n6985), .ZN(n6988)
         );
  OAI211_X1 U8650 ( .C1(n10059), .C2(n6990), .A(n6989), .B(n6988), .ZN(
        P2_U3249) );
  NOR2_X1 U8651 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6028), .ZN(n6995) );
  AOI211_X1 U8652 ( .C1(n6993), .C2(n6992), .A(n6991), .B(n10060), .ZN(n6994)
         );
  AOI211_X1 U8653 ( .C1(n10058), .C2(P2_ADDR_REG_7__SCAN_IN), .A(n6995), .B(
        n6994), .ZN(n7000) );
  OAI211_X1 U8654 ( .C1(n6998), .C2(n6997), .A(n10057), .B(n6996), .ZN(n6999)
         );
  OAI211_X1 U8655 ( .C1(n10059), .C2(n7001), .A(n7000), .B(n6999), .ZN(
        P2_U3252) );
  INV_X1 U8656 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n7010) );
  INV_X1 U8657 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n7207) );
  AOI21_X1 U8658 ( .B1(n4394), .B2(n7207), .A(P1_IR_REG_0__SCAN_IN), .ZN(n7003) );
  MUX2_X1 U8659 ( .A(P1_IR_REG_0__SCAN_IN), .B(n7003), .S(n7002), .Z(n7004) );
  AND4_X1 U8660 ( .A1(n7006), .A2(P1_STATE_REG_SCAN_IN), .A3(n7005), .A4(n7004), .ZN(n7008) );
  NOR3_X1 U8661 ( .A1(n9902), .A2(P1_REG1_REG_0__SCAN_IN), .A3(n4528), .ZN(
        n7007) );
  AOI211_X1 U8662 ( .C1(P1_REG3_REG_0__SCAN_IN), .C2(P1_U3084), .A(n7008), .B(
        n7007), .ZN(n7009) );
  OAI21_X1 U8663 ( .B1(n9945), .B2(n7010), .A(n7009), .ZN(P1_U3241) );
  INV_X1 U8664 ( .A(n7011), .ZN(n7013) );
  INV_X1 U8665 ( .A(n8384), .ZN(n7335) );
  OAI222_X1 U8666 ( .A1(n8124), .A2(n7012), .B1(n8859), .B2(n7013), .C1(
        P2_U3152), .C2(n7335), .ZN(P2_U3346) );
  INV_X1 U8667 ( .A(n7306), .ZN(n7216) );
  OAI222_X1 U8668 ( .A1(n9449), .A2(n9696), .B1(n9452), .B2(n7013), .C1(
        P1_U3084), .C2(n7216), .ZN(P1_U3341) );
  INV_X1 U8669 ( .A(n7014), .ZN(n7040) );
  AOI22_X1 U8670 ( .A1(n7600), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n9730), .ZN(n7015) );
  OAI21_X1 U8671 ( .B1(n7040), .B2(n9445), .A(n7015), .ZN(P1_U3340) );
  INV_X1 U8672 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n9591) );
  NAND2_X1 U8673 ( .A1(n9093), .A2(P1_U4006), .ZN(n7016) );
  OAI21_X1 U8674 ( .B1(P1_U4006), .B2(n9591), .A(n7016), .ZN(P1_U3586) );
  AND2_X1 U8675 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3152), .ZN(n7826) );
  MUX2_X1 U8676 ( .A(n7018), .B(P2_REG1_REG_9__SCAN_IN), .S(n7141), .Z(n7019)
         );
  AOI211_X1 U8677 ( .C1(n7020), .C2(n7019), .A(n7135), .B(n10060), .ZN(n7021)
         );
  AOI211_X1 U8678 ( .C1(n10058), .C2(P2_ADDR_REG_9__SCAN_IN), .A(n7826), .B(
        n7021), .ZN(n7029) );
  NAND2_X1 U8679 ( .A1(n7022), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n7024) );
  NAND2_X1 U8680 ( .A1(n7024), .A2(n7023), .ZN(n7027) );
  MUX2_X1 U8681 ( .A(n7711), .B(P2_REG2_REG_9__SCAN_IN), .S(n7141), .Z(n7025)
         );
  INV_X1 U8682 ( .A(n7025), .ZN(n7026) );
  OAI211_X1 U8683 ( .C1(n7027), .C2(n7026), .A(n10057), .B(n7142), .ZN(n7028)
         );
  OAI211_X1 U8684 ( .C1(n10059), .C2(n7030), .A(n7029), .B(n7028), .ZN(
        P2_U3254) );
  INV_X1 U8685 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n7039) );
  INV_X1 U8686 ( .A(n9922), .ZN(n9931) );
  AND2_X1 U8687 ( .A1(P1_U3084), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n7327) );
  XNOR2_X1 U8688 ( .A(n7092), .B(P1_REG2_REG_7__SCAN_IN), .ZN(n7093) );
  INV_X1 U8689 ( .A(n7031), .ZN(n7034) );
  XNOR2_X1 U8690 ( .A(n7093), .B(n7091), .ZN(n7036) );
  XNOR2_X1 U8691 ( .A(n7092), .B(P1_REG1_REG_7__SCAN_IN), .ZN(n7077) );
  OAI21_X1 U8692 ( .B1(n7034), .B2(P1_REG1_REG_6__SCAN_IN), .A(n7033), .ZN(
        n7075) );
  XNOR2_X1 U8693 ( .A(n7077), .B(n7075), .ZN(n7035) );
  OAI22_X1 U8694 ( .A1(n9886), .A2(n7036), .B1(n7035), .B2(n9902), .ZN(n7037)
         );
  AOI211_X1 U8695 ( .C1(n9931), .C2(n7092), .A(n7327), .B(n7037), .ZN(n7038)
         );
  OAI21_X1 U8696 ( .B1(n9945), .B2(n7039), .A(n7038), .ZN(P1_U3248) );
  INV_X1 U8697 ( .A(n7452), .ZN(n7344) );
  OAI222_X1 U8698 ( .A1(n8124), .A2(n7041), .B1(n8859), .B2(n7040), .C1(n7344), 
        .C2(P2_U3152), .ZN(P2_U3345) );
  NAND2_X1 U8699 ( .A1(n7042), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7108) );
  INV_X1 U8700 ( .A(n7043), .ZN(n7044) );
  AOI211_X1 U8701 ( .C1(n10032), .C2(n7045), .A(n7108), .B(n7044), .ZN(n7157)
         );
  INV_X1 U8702 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n7049) );
  AOI22_X1 U8703 ( .A1(n8991), .A2(n6440), .B1(n7521), .B2(n8997), .ZN(n7048)
         );
  NAND2_X1 U8704 ( .A1(n7046), .A2(n8976), .ZN(n7047) );
  OAI211_X1 U8705 ( .C1(n7157), .C2(n7049), .A(n7048), .B(n7047), .ZN(P1_U3230) );
  INV_X1 U8706 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n7061) );
  NOR2_X1 U8707 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n5392), .ZN(n7169) );
  OAI211_X1 U8708 ( .C1(n7052), .C2(n7051), .A(n9938), .B(n7050), .ZN(n7057)
         );
  OAI211_X1 U8709 ( .C1(n7055), .C2(n7054), .A(n9941), .B(n7053), .ZN(n7056)
         );
  NAND2_X1 U8710 ( .A1(n7057), .A2(n7056), .ZN(n7058) );
  AOI211_X1 U8711 ( .C1(n9931), .C2(n7059), .A(n7169), .B(n7058), .ZN(n7060)
         );
  OAI21_X1 U8712 ( .B1(n7061), .B2(n9945), .A(n7060), .ZN(P1_U3244) );
  INV_X1 U8713 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n7074) );
  INV_X1 U8714 ( .A(n7062), .ZN(n7072) );
  AND2_X1 U8715 ( .A1(P1_U3084), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n7357) );
  AOI21_X1 U8716 ( .B1(n7065), .B2(n7064), .A(n7063), .ZN(n7070) );
  OAI211_X1 U8717 ( .C1(n7068), .C2(n7067), .A(n9938), .B(n7066), .ZN(n7069)
         );
  OAI21_X1 U8718 ( .B1(n9886), .B2(n7070), .A(n7069), .ZN(n7071) );
  AOI211_X1 U8719 ( .C1(n9931), .C2(n7072), .A(n7357), .B(n7071), .ZN(n7073)
         );
  OAI21_X1 U8720 ( .B1(n9945), .B2(n7074), .A(n7073), .ZN(P1_U3246) );
  INV_X1 U8721 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n7105) );
  XNOR2_X1 U8722 ( .A(n7095), .B(P1_REG1_REG_9__SCAN_IN), .ZN(n9925) );
  INV_X1 U8723 ( .A(n7075), .ZN(n7076) );
  OR2_X1 U8724 ( .A1(n7077), .A2(n7076), .ZN(n7081) );
  INV_X1 U8725 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n7078) );
  NAND2_X1 U8726 ( .A1(n7079), .A2(n7078), .ZN(n7080) );
  NAND2_X1 U8727 ( .A1(n7081), .A2(n7080), .ZN(n9899) );
  OR2_X1 U8728 ( .A1(n7090), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n7083) );
  NAND2_X1 U8729 ( .A1(n7090), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n7082) );
  NAND2_X1 U8730 ( .A1(n7083), .A2(n7082), .ZN(n9898) );
  NOR2_X1 U8731 ( .A1(n9899), .A2(n9898), .ZN(n9901) );
  AOI21_X1 U8732 ( .B1(P1_REG1_REG_8__SCAN_IN), .B2(n7090), .A(n9901), .ZN(
        n7084) );
  INV_X1 U8733 ( .A(n7084), .ZN(n9924) );
  OAI22_X1 U8734 ( .A1(n9925), .A2(n9924), .B1(P1_REG1_REG_9__SCAN_IN), .B2(
        n7095), .ZN(n7087) );
  INV_X1 U8735 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n7804) );
  AOI22_X1 U8736 ( .A1(P1_REG1_REG_10__SCAN_IN), .A2(n7219), .B1(n7085), .B2(
        n7804), .ZN(n7086) );
  NAND2_X1 U8737 ( .A1(n7086), .A2(n7087), .ZN(n7210) );
  OAI21_X1 U8738 ( .B1(n7087), .B2(n7086), .A(n7210), .ZN(n7101) );
  INV_X1 U8739 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n7088) );
  XNOR2_X1 U8740 ( .A(n7095), .B(n7088), .ZN(n9917) );
  OR2_X1 U8741 ( .A1(n7090), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n7094) );
  NOR2_X1 U8742 ( .A1(n7090), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n7089) );
  AOI21_X1 U8743 ( .B1(P1_REG2_REG_8__SCAN_IN), .B2(n7090), .A(n7089), .ZN(
        n9910) );
  NAND2_X1 U8744 ( .A1(n9910), .A2(n9909), .ZN(n9908) );
  OR2_X1 U8745 ( .A1(n7219), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n7097) );
  NAND2_X1 U8746 ( .A1(P1_REG2_REG_10__SCAN_IN), .A2(n7219), .ZN(n7096) );
  NAND2_X1 U8747 ( .A1(n7097), .A2(n7096), .ZN(n7098) );
  AOI211_X1 U8748 ( .C1(n7099), .C2(n7098), .A(n7218), .B(n9886), .ZN(n7100)
         );
  AOI21_X1 U8749 ( .B1(n9938), .B2(n7101), .A(n7100), .ZN(n7104) );
  NOR2_X1 U8750 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7102), .ZN(n7578) );
  AOI21_X1 U8751 ( .B1(n9931), .B2(n7219), .A(n7578), .ZN(n7103) );
  OAI211_X1 U8752 ( .C1(n9945), .C2(n7105), .A(n7104), .B(n7103), .ZN(P1_U3251) );
  INV_X1 U8753 ( .A(n7365), .ZN(n7106) );
  OAI21_X1 U8754 ( .B1(n10034), .B2(n9086), .A(n7106), .ZN(n7107) );
  NAND2_X1 U8755 ( .A1(n7112), .A2(n7109), .ZN(n7114) );
  INV_X1 U8756 ( .A(n7110), .ZN(n7111) );
  AOI22_X1 U8757 ( .A1(n7114), .A2(n7113), .B1(n7112), .B2(n7111), .ZN(n7364)
         );
  INV_X1 U8758 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n7123) );
  INV_X1 U8759 ( .A(n7467), .ZN(n7116) );
  INV_X1 U8760 ( .A(n7121), .ZN(n7115) );
  NOR2_X1 U8761 ( .A1(n7116), .A2(n7115), .ZN(n7119) );
  AOI22_X1 U8762 ( .A1(n7120), .A2(n7119), .B1(n9285), .B2(n6440), .ZN(n7420)
         );
  OAI21_X1 U8763 ( .B1(n7408), .B2(n7121), .A(n7420), .ZN(n7205) );
  NAND2_X1 U8764 ( .A1(n7205), .A2(n10042), .ZN(n7122) );
  OAI21_X1 U8765 ( .B1(n10042), .B2(n7123), .A(n7122), .ZN(P1_U3454) );
  INV_X1 U8766 ( .A(n9733), .ZN(n7124) );
  INV_X1 U8767 ( .A(n7845), .ZN(n7840) );
  OAI222_X1 U8768 ( .A1(n8124), .A2(n7125), .B1(n8859), .B2(n7124), .C1(n7840), 
        .C2(P2_U3152), .ZN(P2_U3344) );
  NAND2_X1 U8769 ( .A1(n7126), .A2(n7127), .ZN(n7129) );
  XNOR2_X1 U8770 ( .A(n7129), .B(n7128), .ZN(n7134) );
  INV_X1 U8771 ( .A(n7157), .ZN(n7132) );
  AOI22_X1 U8772 ( .A1(n8991), .A2(n9018), .B1(n8979), .B2(n7361), .ZN(n7130)
         );
  OAI21_X1 U8773 ( .B1(n9991), .B2(n8985), .A(n7130), .ZN(n7131) );
  AOI21_X1 U8774 ( .B1(n7132), .B2(P1_REG3_REG_1__SCAN_IN), .A(n7131), .ZN(
        n7133) );
  OAI21_X1 U8775 ( .B1(n7134), .B2(n8999), .A(n7133), .ZN(P1_U3220) );
  NAND2_X1 U8776 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3152), .ZN(n7832) );
  INV_X1 U8777 ( .A(n7832), .ZN(n7140) );
  MUX2_X1 U8778 ( .A(n7136), .B(P2_REG1_REG_10__SCAN_IN), .S(n7184), .Z(n7137)
         );
  NOR2_X1 U8779 ( .A1(n7138), .A2(n7137), .ZN(n7183) );
  AOI211_X1 U8780 ( .C1(n7138), .C2(n7137), .A(n7183), .B(n10060), .ZN(n7139)
         );
  AOI211_X1 U8781 ( .C1(n10058), .C2(P2_ADDR_REG_10__SCAN_IN), .A(n7140), .B(
        n7139), .ZN(n7148) );
  NAND2_X1 U8782 ( .A1(n7141), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n7143) );
  MUX2_X1 U8783 ( .A(n7813), .B(P2_REG2_REG_10__SCAN_IN), .S(n7184), .Z(n7144)
         );
  INV_X1 U8784 ( .A(n7144), .ZN(n7145) );
  NAND2_X1 U8785 ( .A1(n7145), .A2(n7146), .ZN(n7177) );
  OAI211_X1 U8786 ( .C1(n7146), .C2(n7145), .A(n10057), .B(n7177), .ZN(n7147)
         );
  OAI211_X1 U8787 ( .C1(n10059), .C2(n7149), .A(n7148), .B(n7147), .ZN(
        P2_U3255) );
  OAI21_X1 U8788 ( .B1(n4475), .B2(n7151), .A(n7150), .ZN(n7152) );
  NAND2_X1 U8789 ( .A1(n7152), .A2(n8976), .ZN(n7155) );
  OAI22_X1 U8790 ( .A1(n8995), .A2(n7513), .B1(n7514), .B2(n8972), .ZN(n7153)
         );
  AOI21_X1 U8791 ( .B1(n7520), .B2(n8997), .A(n7153), .ZN(n7154) );
  OAI211_X1 U8792 ( .C1(n7157), .C2(n7156), .A(n7155), .B(n7154), .ZN(P1_U3235) );
  INV_X1 U8793 ( .A(n7158), .ZN(n7176) );
  AOI22_X1 U8794 ( .A1(n8420), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_16__SCAN_IN), .B2(n8856), .ZN(n7159) );
  OAI21_X1 U8795 ( .B1(n7176), .B2(n8859), .A(n7159), .ZN(P2_U3342) );
  INV_X1 U8796 ( .A(n7160), .ZN(n7162) );
  OAI222_X1 U8797 ( .A1(n9449), .A2(n7161), .B1(n9452), .B2(n7162), .C1(
        P1_U3084), .C2(n9036), .ZN(P1_U3338) );
  INV_X1 U8798 ( .A(n8404), .ZN(n8394) );
  OAI222_X1 U8799 ( .A1(n8124), .A2(n7163), .B1(n8859), .B2(n7162), .C1(
        P2_U3152), .C2(n8394), .ZN(P2_U3343) );
  OAI21_X1 U8800 ( .B1(n7166), .B2(n7165), .A(n7164), .ZN(n7167) );
  NAND2_X1 U8801 ( .A1(n7167), .A2(n8976), .ZN(n7171) );
  OAI22_X1 U8802 ( .A1(n10003), .A2(n8985), .B1(n8972), .B2(n7558), .ZN(n7168)
         );
  AOI211_X1 U8803 ( .C1(n8979), .C2(n9018), .A(n7169), .B(n7168), .ZN(n7170)
         );
  OAI211_X1 U8804 ( .C1(P1_REG3_REG_3__SCAN_IN), .C2(n8981), .A(n7171), .B(
        n7170), .ZN(P1_U3216) );
  NOR2_X1 U8805 ( .A1(n8334), .A2(P2_U3152), .ZN(n7267) );
  INV_X1 U8806 ( .A(n8331), .ZN(n8304) );
  AOI22_X1 U8807 ( .A1(n8304), .A2(n6718), .B1(n7792), .B2(n8319), .ZN(n7175)
         );
  OR2_X1 U8808 ( .A1(n8321), .A2(n8165), .ZN(n8291) );
  INV_X1 U8809 ( .A(n5990), .ZN(n7266) );
  OAI22_X1 U8810 ( .A1(n8291), .A2(n7266), .B1(n10122), .B2(n8321), .ZN(n7173)
         );
  NAND2_X1 U8811 ( .A1(n7173), .A2(n7172), .ZN(n7174) );
  OAI211_X1 U8812 ( .C1(n7267), .C2(n7790), .A(n7175), .B(n7174), .ZN(P2_U3234) );
  INV_X1 U8813 ( .A(n9053), .ZN(n9044) );
  OAI222_X1 U8814 ( .A1(n9445), .A2(n7176), .B1(n9044), .B2(P1_U3084), .C1(
        n9593), .C2(n9449), .ZN(P1_U3337) );
  NAND2_X1 U8815 ( .A1(n7184), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n7178) );
  NAND2_X1 U8816 ( .A1(n7178), .A2(n7177), .ZN(n7181) );
  MUX2_X1 U8817 ( .A(n7179), .B(P2_REG2_REG_11__SCAN_IN), .S(n7339), .Z(n7180)
         );
  NOR2_X1 U8818 ( .A1(n7181), .A2(n7180), .ZN(n7333) );
  AOI21_X1 U8819 ( .B1(n7181), .B2(n7180), .A(n7333), .ZN(n7193) );
  INV_X1 U8820 ( .A(n10057), .ZN(n7850) );
  MUX2_X1 U8821 ( .A(n7182), .B(P2_REG1_REG_11__SCAN_IN), .S(n7339), .Z(n7186)
         );
  AOI21_X1 U8822 ( .B1(n7184), .B2(P2_REG1_REG_10__SCAN_IN), .A(n7183), .ZN(
        n7185) );
  NOR2_X1 U8823 ( .A1(n7185), .A2(n7186), .ZN(n7338) );
  AOI21_X1 U8824 ( .B1(n7186), .B2(n7185), .A(n7338), .ZN(n7190) );
  INV_X1 U8825 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n7188) );
  OR2_X1 U8826 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7945), .ZN(n7187) );
  OAI21_X1 U8827 ( .B1(n8460), .B2(n7188), .A(n7187), .ZN(n7189) );
  AOI21_X1 U8828 ( .B1(n10056), .B2(n7190), .A(n7189), .ZN(n7192) );
  NAND2_X1 U8829 ( .A1(n9753), .A2(n7339), .ZN(n7191) );
  OAI211_X1 U8830 ( .C1(n7193), .C2(n7850), .A(n7192), .B(n7191), .ZN(P2_U3256) );
  INV_X1 U8831 ( .A(n7194), .ZN(n7196) );
  NAND2_X1 U8832 ( .A1(n7196), .A2(n7195), .ZN(n7197) );
  XNOR2_X1 U8833 ( .A(n7198), .B(n7197), .ZN(n7202) );
  NOR2_X1 U8834 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n5403), .ZN(n9893) );
  OAI22_X1 U8835 ( .A1(n8995), .A2(n7514), .B1(n7431), .B2(n8985), .ZN(n7199)
         );
  AOI211_X1 U8836 ( .C1(n8991), .C2(n9015), .A(n9893), .B(n7199), .ZN(n7201)
         );
  NAND2_X1 U8837 ( .A1(n8992), .A2(n7429), .ZN(n7200) );
  OAI211_X1 U8838 ( .C1(n7202), .C2(n8999), .A(n7201), .B(n7200), .ZN(P1_U3228) );
  NAND2_X1 U8839 ( .A1(n7205), .A2(n4392), .ZN(n7206) );
  OAI21_X1 U8840 ( .B1(n4392), .B2(n7207), .A(n7206), .ZN(P1_U3523) );
  INV_X1 U8841 ( .A(n7208), .ZN(n7228) );
  AOI22_X1 U8842 ( .A1(n9069), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n9730), .ZN(n7209) );
  OAI21_X1 U8843 ( .B1(n7228), .B2(n9452), .A(n7209), .ZN(P1_U3336) );
  INV_X1 U8844 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n9874) );
  AOI22_X1 U8845 ( .A1(n9930), .A2(P1_REG1_REG_11__SCAN_IN), .B1(n9874), .B2(
        n7217), .ZN(n9937) );
  OAI21_X1 U8846 ( .B1(P1_REG1_REG_10__SCAN_IN), .B2(n7219), .A(n7210), .ZN(
        n9936) );
  NAND2_X1 U8847 ( .A1(n9937), .A2(n9936), .ZN(n9935) );
  OAI21_X1 U8848 ( .B1(P1_REG1_REG_11__SCAN_IN), .B2(n9930), .A(n9935), .ZN(
        n7213) );
  INV_X1 U8849 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n7211) );
  MUX2_X1 U8850 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n7211), .S(n7306), .Z(n7212)
         );
  NAND2_X1 U8851 ( .A1(n7212), .A2(n7213), .ZN(n7301) );
  OAI21_X1 U8852 ( .B1(n7213), .B2(n7212), .A(n7301), .ZN(n7225) );
  INV_X1 U8853 ( .A(n9945), .ZN(n9894) );
  NAND2_X1 U8854 ( .A1(n9894), .A2(P1_ADDR_REG_12__SCAN_IN), .ZN(n7215) );
  NAND2_X1 U8855 ( .A1(P1_REG3_REG_12__SCAN_IN), .A2(P1_U3084), .ZN(n7214) );
  OAI211_X1 U8856 ( .C1(n7216), .C2(n9922), .A(n7215), .B(n7214), .ZN(n7224)
         );
  INV_X1 U8857 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n9551) );
  AOI22_X1 U8858 ( .A1(n9930), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n9551), .B2(
        n7217), .ZN(n9934) );
  OAI21_X1 U8859 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n9930), .A(n9932), .ZN(
        n7222) );
  NAND2_X1 U8860 ( .A1(P1_REG2_REG_12__SCAN_IN), .A2(n7306), .ZN(n7220) );
  OAI21_X1 U8861 ( .B1(n7306), .B2(P1_REG2_REG_12__SCAN_IN), .A(n7220), .ZN(
        n7221) );
  AOI211_X1 U8862 ( .C1(n7222), .C2(n7221), .A(n7305), .B(n9886), .ZN(n7223)
         );
  AOI211_X1 U8863 ( .C1(n9938), .C2(n7225), .A(n7224), .B(n7223), .ZN(n7226)
         );
  INV_X1 U8864 ( .A(n7226), .ZN(P1_U3253) );
  INV_X1 U8865 ( .A(n8432), .ZN(n7227) );
  OAI222_X1 U8866 ( .A1(n8124), .A2(n9695), .B1(n8859), .B2(n7228), .C1(n7227), 
        .C2(P2_U3152), .ZN(P2_U3341) );
  AND2_X1 U8867 ( .A1(n7675), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7231) );
  INV_X1 U8868 ( .A(n7676), .ZN(n7230) );
  NAND4_X1 U8869 ( .A1(n7679), .A2(n7231), .A3(n7230), .A4(n7229), .ZN(n7250)
         );
  NAND2_X1 U8870 ( .A1(n7680), .A2(n7662), .ZN(n7235) );
  AND2_X1 U8871 ( .A1(n8668), .A2(n7233), .ZN(n7234) );
  NAND2_X1 U8872 ( .A1(n7235), .A2(n7234), .ZN(n8717) );
  NAND2_X1 U8873 ( .A1(n7773), .A2(n7236), .ZN(n7766) );
  OR2_X1 U8874 ( .A1(n6725), .A2(n7902), .ZN(n7237) );
  INV_X1 U8875 ( .A(n8352), .ZN(n7257) );
  NAND2_X1 U8876 ( .A1(n7257), .A2(n10141), .ZN(n7238) );
  NAND2_X1 U8877 ( .A1(n10100), .A2(n10101), .ZN(n7240) );
  OR2_X1 U8878 ( .A1(n8351), .A2(n10103), .ZN(n7239) );
  XNOR2_X1 U8879 ( .A(n7665), .B(n7666), .ZN(n7788) );
  NAND2_X1 U8880 ( .A1(n7241), .A2(n7242), .ZN(n7244) );
  XNOR2_X1 U8881 ( .A(n7243), .B(n7244), .ZN(n7246) );
  INV_X1 U8882 ( .A(n8351), .ZN(n7759) );
  INV_X1 U8883 ( .A(n8349), .ZN(n10073) );
  OAI22_X1 U8884 ( .A1(n7759), .A2(n10072), .B1(n10073), .B2(n10070), .ZN(
        n7317) );
  AOI21_X1 U8885 ( .B1(n7246), .B2(n8722), .A(n7317), .ZN(n7779) );
  NAND2_X1 U8886 ( .A1(n7900), .A2(n10141), .ZN(n10093) );
  OR2_X1 U8887 ( .A1(n10093), .A2(n10103), .ZN(n10094) );
  AOI211_X1 U8888 ( .C1(n7785), .C2(n10094), .A(n10194), .B(n7743), .ZN(n7781)
         );
  AOI21_X1 U8889 ( .B1(n10128), .B2(n7785), .A(n7781), .ZN(n7248) );
  OAI211_X1 U8890 ( .C1(n10130), .C2(n7788), .A(n7779), .B(n7248), .ZN(n7251)
         );
  NAND2_X1 U8891 ( .A1(n7251), .A2(n10202), .ZN(n7249) );
  OAI21_X1 U8892 ( .B1(n10202), .B2(n5914), .A(n7249), .ZN(P2_U3466) );
  INV_X1 U8893 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n7253) );
  NAND2_X1 U8894 ( .A1(n7251), .A2(n10219), .ZN(n7252) );
  OAI21_X1 U8895 ( .B1(n10219), .B2(n7253), .A(n7252), .ZN(P2_U3525) );
  INV_X1 U8896 ( .A(n7276), .ZN(n7254) );
  AOI211_X1 U8897 ( .C1(n7256), .C2(n7255), .A(n8321), .B(n7254), .ZN(n7261)
         );
  OAI22_X1 U8898 ( .A1(n10136), .A2(n8337), .B1(n8331), .B2(n7257), .ZN(n7260)
         );
  OAI22_X1 U8899 ( .A1(n7267), .A2(n7258), .B1(n4943), .B2(n8330), .ZN(n7259)
         );
  OR3_X1 U8900 ( .A1(n7261), .A2(n7260), .A3(n7259), .ZN(P2_U3239) );
  OAI21_X1 U8901 ( .B1(n7264), .B2(n7263), .A(n7262), .ZN(n7270) );
  INV_X1 U8902 ( .A(n6725), .ZN(n7758) );
  OAI22_X1 U8903 ( .A1(n7265), .A2(n8337), .B1(n8331), .B2(n7758), .ZN(n7269)
         );
  OAI22_X1 U8904 ( .A1(n7267), .A2(n7770), .B1(n7266), .B2(n8330), .ZN(n7268)
         );
  AOI211_X1 U8905 ( .C1(n8325), .C2(n7270), .A(n7269), .B(n7268), .ZN(n7271)
         );
  INV_X1 U8906 ( .A(n7271), .ZN(P2_U3224) );
  INV_X1 U8907 ( .A(n8330), .ZN(n8307) );
  OAI22_X1 U8908 ( .A1(n8317), .A2(P2_REG3_REG_3__SCAN_IN), .B1(
        P2_STATE_REG_SCAN_IN), .B2(n5928), .ZN(n7273) );
  OAI22_X1 U8909 ( .A1(n10141), .A2(n8337), .B1(n8331), .B2(n7759), .ZN(n7272)
         );
  AOI211_X1 U8910 ( .C1(n8307), .C2(n6725), .A(n7273), .B(n7272), .ZN(n7282)
         );
  INV_X1 U8911 ( .A(n7274), .ZN(n7275) );
  AOI21_X1 U8912 ( .B1(n7276), .B2(n7275), .A(n8321), .ZN(n7280) );
  NOR3_X1 U8913 ( .A1(n8291), .A2(n7277), .A3(n7758), .ZN(n7279) );
  OAI21_X1 U8914 ( .B1(n7280), .B2(n7279), .A(n7278), .ZN(n7281) );
  NAND2_X1 U8915 ( .A1(n7282), .A2(n7281), .ZN(P2_U3220) );
  INV_X1 U8916 ( .A(n7283), .ZN(n7284) );
  NAND2_X1 U8917 ( .A1(n7284), .A2(n7285), .ZN(n7286) );
  MUX2_X1 U8918 ( .A(n7286), .B(n7285), .S(n7292), .Z(n7295) );
  NAND2_X1 U8919 ( .A1(n8352), .A2(n8684), .ZN(n7288) );
  NAND2_X1 U8920 ( .A1(n8350), .A2(n8686), .ZN(n7287) );
  NAND2_X1 U8921 ( .A1(n7288), .A2(n7287), .ZN(n10091) );
  OAI22_X1 U8922 ( .A1(n8337), .A2(n10147), .B1(n8317), .B2(n10097), .ZN(n7289) );
  AOI211_X1 U8923 ( .C1(n8315), .C2(n10091), .A(n7290), .B(n7289), .ZN(n7294)
         );
  INV_X1 U8924 ( .A(n8291), .ZN(n8323) );
  NAND4_X1 U8925 ( .A1(n7292), .A2(n8323), .A3(n7291), .A4(n8351), .ZN(n7293)
         );
  OAI211_X1 U8926 ( .C1(n7295), .C2(n8321), .A(n7294), .B(n7293), .ZN(P2_U3232) );
  INV_X1 U8927 ( .A(n7296), .ZN(n7299) );
  AOI22_X1 U8928 ( .A1(n8447), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_18__SCAN_IN), .B2(n8856), .ZN(n7297) );
  OAI21_X1 U8929 ( .B1(n7299), .B2(n8859), .A(n7297), .ZN(P2_U3340) );
  AOI22_X1 U8930 ( .A1(n9080), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n9730), .ZN(n7298) );
  OAI21_X1 U8931 ( .B1(n7299), .B2(n9445), .A(n7298), .ZN(P1_U3335) );
  INV_X1 U8932 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n7314) );
  INV_X1 U8933 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n7300) );
  MUX2_X1 U8934 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n7300), .S(n7600), .Z(n7303)
         );
  OAI21_X1 U8935 ( .B1(n7306), .B2(P1_REG1_REG_12__SCAN_IN), .A(n7301), .ZN(
        n7302) );
  NAND2_X1 U8936 ( .A1(n7303), .A2(n7302), .ZN(n7594) );
  OAI21_X1 U8937 ( .B1(n7303), .B2(n7302), .A(n7594), .ZN(n7312) );
  INV_X1 U8938 ( .A(n7600), .ZN(n7304) );
  NAND2_X1 U8939 ( .A1(P1_U3084), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n7974) );
  OAI21_X1 U8940 ( .B1(n9922), .B2(n7304), .A(n7974), .ZN(n7311) );
  NAND2_X1 U8941 ( .A1(P1_REG2_REG_13__SCAN_IN), .A2(n7600), .ZN(n7307) );
  OAI21_X1 U8942 ( .B1(n7600), .B2(P1_REG2_REG_13__SCAN_IN), .A(n7307), .ZN(
        n7308) );
  AOI211_X1 U8943 ( .C1(n7309), .C2(n7308), .A(n7599), .B(n9886), .ZN(n7310)
         );
  AOI211_X1 U8944 ( .C1(n9938), .C2(n7312), .A(n7311), .B(n7310), .ZN(n7313)
         );
  OAI21_X1 U8945 ( .B1(n9945), .B2(n7314), .A(n7313), .ZN(P1_U3254) );
  XNOR2_X1 U8946 ( .A(n7316), .B(n7315), .ZN(n7321) );
  AOI22_X1 U8947 ( .A1(n8315), .A2(n7317), .B1(P2_REG3_REG_5__SCAN_IN), .B2(
        P2_U3152), .ZN(n7320) );
  INV_X1 U8948 ( .A(n7782), .ZN(n7318) );
  AOI22_X1 U8949 ( .A1(n8319), .A2(n7785), .B1(n8334), .B2(n7318), .ZN(n7319)
         );
  OAI211_X1 U8950 ( .C1(n7321), .C2(n8321), .A(n7320), .B(n7319), .ZN(P2_U3229) );
  XOR2_X1 U8951 ( .A(n7324), .B(n7323), .Z(n7325) );
  XNOR2_X1 U8952 ( .A(n7322), .B(n7325), .ZN(n7331) );
  NOR2_X1 U8953 ( .A1(n8972), .A2(n9958), .ZN(n7326) );
  AOI211_X1 U8954 ( .C1(n8979), .C2(n9014), .A(n7327), .B(n7326), .ZN(n7328)
         );
  OAI21_X1 U8955 ( .B1(n10026), .B2(n8985), .A(n7328), .ZN(n7329) );
  AOI21_X1 U8956 ( .B1(n7480), .B2(n8992), .A(n7329), .ZN(n7330) );
  OAI21_X1 U8957 ( .B1(n7331), .B2(n8999), .A(n7330), .ZN(P1_U3211) );
  MUX2_X1 U8958 ( .A(P2_REG2_REG_12__SCAN_IN), .B(n7332), .S(n8384), .Z(n8380)
         );
  NAND2_X1 U8959 ( .A1(n8380), .A2(n8381), .ZN(n8379) );
  OAI21_X1 U8960 ( .B1(n7332), .B2(n7335), .A(n8379), .ZN(n7337) );
  AOI22_X1 U8961 ( .A1(n7452), .A2(n8003), .B1(P2_REG2_REG_13__SCAN_IN), .B2(
        n7344), .ZN(n7336) );
  NOR2_X1 U8962 ( .A1(n7337), .A2(n7336), .ZN(n7447) );
  AOI21_X1 U8963 ( .B1(n7337), .B2(n7336), .A(n7447), .ZN(n7348) );
  AOI22_X1 U8964 ( .A1(n7452), .A2(P2_REG1_REG_13__SCAN_IN), .B1(n6105), .B2(
        n7344), .ZN(n7342) );
  MUX2_X1 U8965 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n7340), .S(n8384), .Z(n8387)
         );
  OAI21_X1 U8966 ( .B1(n7342), .B2(n7341), .A(n7451), .ZN(n7343) );
  NAND2_X1 U8967 ( .A1(n7343), .A2(n10056), .ZN(n7347) );
  AND2_X1 U8968 ( .A1(P2_U3152), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n8051) );
  NOR2_X1 U8969 ( .A1(n10059), .A2(n7344), .ZN(n7345) );
  AOI211_X1 U8970 ( .C1(n10058), .C2(P2_ADDR_REG_13__SCAN_IN), .A(n8051), .B(
        n7345), .ZN(n7346) );
  OAI211_X1 U8971 ( .C1(n7348), .C2(n7850), .A(n7347), .B(n7346), .ZN(P2_U3258) );
  INV_X1 U8972 ( .A(n7349), .ZN(n8122) );
  OAI222_X1 U8973 ( .A1(n9449), .A2(n7350), .B1(n9445), .B2(n8122), .C1(n9086), 
        .C2(P1_U3084), .ZN(P1_U3334) );
  INV_X1 U8974 ( .A(n7533), .ZN(n7360) );
  XNOR2_X1 U8975 ( .A(n7351), .B(n7352), .ZN(n7353) );
  NAND2_X1 U8976 ( .A1(n7353), .A2(n7354), .ZN(n7435) );
  OAI21_X1 U8977 ( .B1(n7354), .B2(n7353), .A(n7435), .ZN(n7355) );
  NAND2_X1 U8978 ( .A1(n7355), .A2(n8976), .ZN(n7359) );
  OAI22_X1 U8979 ( .A1(n7538), .A2(n8985), .B1(n8972), .B2(n7477), .ZN(n7356)
         );
  AOI211_X1 U8980 ( .C1(n8979), .C2(n9016), .A(n7357), .B(n7356), .ZN(n7358)
         );
  OAI211_X1 U8981 ( .C1(n8981), .C2(n7360), .A(n7359), .B(n7358), .ZN(P1_U3225) );
  OAI21_X1 U8982 ( .B1(n7363), .B2(n7362), .A(n7401), .ZN(n9989) );
  INV_X1 U8983 ( .A(n7364), .ZN(n7366) );
  NAND2_X1 U8984 ( .A1(n7365), .A2(n9988), .ZN(n9986) );
  NOR2_X1 U8985 ( .A1(n7366), .A2(n9986), .ZN(n7367) );
  NAND2_X1 U8986 ( .A1(n7368), .A2(n7367), .ZN(n7479) );
  INV_X2 U8987 ( .A(n9836), .ZN(n9321) );
  NAND2_X1 U8988 ( .A1(n7373), .A2(n9250), .ZN(n7369) );
  INV_X1 U8989 ( .A(n9953), .ZN(n7890) );
  INV_X1 U8990 ( .A(n7370), .ZN(n7371) );
  AOI22_X1 U8991 ( .A1(n9848), .A2(n7522), .B1(n9970), .B2(
        P1_REG2_REG_1__SCAN_IN), .ZN(n7387) );
  OR2_X1 U8992 ( .A1(n7373), .A2(n7372), .ZN(n7375) );
  OR2_X1 U8993 ( .A1(n7416), .A2(n7573), .ZN(n7374) );
  AOI22_X1 U8994 ( .A1(n9287), .A2(n7361), .B1(n9285), .B2(n9018), .ZN(n7382)
         );
  OAI21_X1 U8995 ( .B1(n5573), .B2(n7377), .A(n7376), .ZN(n7380) );
  OR2_X1 U8996 ( .A1(n6434), .A2(n9086), .ZN(n7379) );
  NAND2_X1 U8997 ( .A1(n6433), .A2(n7398), .ZN(n7378) );
  NAND2_X1 U8998 ( .A1(n7380), .A2(n9963), .ZN(n7381) );
  OAI211_X1 U8999 ( .C1(n9989), .C2(n9966), .A(n7382), .B(n7381), .ZN(n9992)
         );
  INV_X1 U9000 ( .A(n10034), .ZN(n10011) );
  XNOR2_X1 U9001 ( .A(n7408), .B(n7522), .ZN(n7383) );
  NAND2_X1 U9002 ( .A1(n10011), .A2(n7383), .ZN(n9990) );
  INV_X1 U9003 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n7384) );
  OAI22_X1 U9004 ( .A1(n9990), .A2(n9250), .B1(n9249), .B2(n7384), .ZN(n7385)
         );
  OAI21_X1 U9005 ( .B1(n9992), .B2(n7385), .A(n9836), .ZN(n7386) );
  OAI211_X1 U9006 ( .C1(n9989), .C2(n7890), .A(n7387), .B(n7386), .ZN(P1_U3290) );
  XOR2_X1 U9007 ( .A(n7389), .B(n7388), .Z(n7390) );
  XNOR2_X1 U9008 ( .A(n7391), .B(n7390), .ZN(n7397) );
  NOR2_X1 U9009 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7392), .ZN(n9903) );
  AOI21_X1 U9010 ( .B1(n8991), .B2(n9011), .A(n9903), .ZN(n7394) );
  NAND2_X1 U9011 ( .A1(n8992), .A2(n7543), .ZN(n7393) );
  OAI211_X1 U9012 ( .C1(n7623), .C2(n8995), .A(n7394), .B(n7393), .ZN(n7395)
         );
  AOI21_X1 U9013 ( .B1(n7633), .B2(n8997), .A(n7395), .ZN(n7396) );
  OAI21_X1 U9014 ( .B1(n7397), .B2(n8999), .A(n7396), .ZN(P1_U3219) );
  INV_X1 U9015 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n9569) );
  NAND2_X1 U9016 ( .A1(n6440), .A2(n7522), .ZN(n7400) );
  NAND2_X1 U9017 ( .A1(n7512), .A2(n7511), .ZN(n7510) );
  NAND2_X1 U9018 ( .A1(n7557), .A2(n9997), .ZN(n7402) );
  NAND2_X1 U9019 ( .A1(n7510), .A2(n7402), .ZN(n7554) );
  NAND2_X1 U9020 ( .A1(n7554), .A2(n7556), .ZN(n7404) );
  NAND2_X1 U9021 ( .A1(n7514), .A2(n10003), .ZN(n7403) );
  NAND2_X1 U9022 ( .A1(n7404), .A2(n7403), .ZN(n7421) );
  NAND2_X1 U9023 ( .A1(n7421), .A2(n7422), .ZN(n7406) );
  NAND2_X1 U9024 ( .A1(n7558), .A2(n7431), .ZN(n7405) );
  NAND2_X1 U9025 ( .A1(n7406), .A2(n7405), .ZN(n7461) );
  XNOR2_X1 U9026 ( .A(n7461), .B(n7618), .ZN(n7537) );
  XNOR2_X1 U9027 ( .A(n7619), .B(n7618), .ZN(n7407) );
  AOI222_X1 U9028 ( .A1(n9016), .A2(n9287), .B1(n9014), .B2(n9285), .C1(n9963), 
        .C2(n7407), .ZN(n7536) );
  NAND3_X1 U9029 ( .A1(n9991), .A2(n9997), .A3(n7408), .ZN(n7563) );
  OR2_X1 U9030 ( .A1(n7563), .A2(n7566), .ZN(n7564) );
  INV_X1 U9031 ( .A(n7428), .ZN(n7409) );
  AOI211_X1 U9032 ( .C1(n7462), .C2(n7409), .A(n10034), .B(n4614), .ZN(n7534)
         );
  AOI21_X1 U9033 ( .B1(n10010), .B2(n7462), .A(n7534), .ZN(n7410) );
  OAI211_X1 U9034 ( .C1(n9418), .C2(n7537), .A(n7536), .B(n7410), .ZN(n7412)
         );
  NAND2_X1 U9035 ( .A1(n7412), .A2(n10042), .ZN(n7411) );
  OAI21_X1 U9036 ( .B1(n10042), .B2(n9569), .A(n7411), .ZN(P1_U3469) );
  NAND2_X1 U9037 ( .A1(n7412), .A2(n4392), .ZN(n7413) );
  OAI21_X1 U9038 ( .B1(n4392), .B2(n6854), .A(n7413), .ZN(P1_U3528) );
  INV_X2 U9039 ( .A(n9249), .ZN(n9969) );
  INV_X1 U9040 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n7414) );
  NOR2_X1 U9041 ( .A1(n9836), .A2(n7414), .ZN(n7415) );
  AOI21_X1 U9042 ( .B1(n9969), .B2(P1_REG3_REG_0__SCAN_IN), .A(n7415), .ZN(
        n7419) );
  OR2_X1 U9043 ( .A1(n7416), .A2(n6433), .ZN(n7417) );
  NOR2_X2 U9044 ( .A1(n9321), .A2(n7417), .ZN(n9952) );
  OAI21_X1 U9045 ( .B1(n9848), .B2(n9952), .A(n7521), .ZN(n7418) );
  OAI211_X1 U9046 ( .C1(n9970), .C2(n7420), .A(n7419), .B(n7418), .ZN(P1_U3291) );
  XNOR2_X1 U9047 ( .A(n7422), .B(n7421), .ZN(n7426) );
  INV_X1 U9048 ( .A(n7426), .ZN(n10016) );
  INV_X1 U9049 ( .A(n9966), .ZN(n9846) );
  XNOR2_X1 U9050 ( .A(n7422), .B(n5628), .ZN(n7424) );
  AOI22_X1 U9051 ( .A1(n9287), .A2(n9017), .B1(n9285), .B2(n9015), .ZN(n7423)
         );
  OAI21_X1 U9052 ( .B1(n7424), .B2(n9844), .A(n7423), .ZN(n7425) );
  AOI21_X1 U9053 ( .B1(n9846), .B2(n7426), .A(n7425), .ZN(n10014) );
  MUX2_X1 U9054 ( .A(n7427), .B(n10014), .S(n9836), .Z(n7434) );
  AOI21_X1 U9055 ( .B1(n10009), .B2(n7564), .A(n7428), .ZN(n10012) );
  INV_X1 U9056 ( .A(n7429), .ZN(n7430) );
  OAI22_X1 U9057 ( .A1(n9972), .A2(n7431), .B1(n7430), .B2(n9249), .ZN(n7432)
         );
  AOI21_X1 U9058 ( .B1(n9952), .B2(n10012), .A(n7432), .ZN(n7433) );
  OAI211_X1 U9059 ( .C1(n10016), .C2(n7890), .A(n7434), .B(n7433), .ZN(
        P1_U3287) );
  OAI21_X1 U9060 ( .B1(n7436), .B2(n7351), .A(n7435), .ZN(n7441) );
  OAI21_X1 U9061 ( .B1(n7439), .B2(n7438), .A(n7437), .ZN(n7440) );
  XNOR2_X1 U9062 ( .A(n7441), .B(n7440), .ZN(n7446) );
  OAI22_X1 U9063 ( .A1(n8995), .A2(n7622), .B1(n10019), .B2(n8985), .ZN(n7442)
         );
  AOI211_X1 U9064 ( .C1(n8991), .C2(n9013), .A(n7443), .B(n7442), .ZN(n7445)
         );
  NAND2_X1 U9065 ( .A1(n8992), .A2(n7614), .ZN(n7444) );
  OAI211_X1 U9066 ( .C1(n7446), .C2(n8999), .A(n7445), .B(n7444), .ZN(P1_U3237) );
  NOR2_X1 U9067 ( .A1(n7452), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n7448) );
  AOI22_X1 U9068 ( .A1(n7845), .A2(n6124), .B1(P2_REG2_REG_14__SCAN_IN), .B2(
        n7840), .ZN(n7449) );
  NOR2_X1 U9069 ( .A1(n7450), .A2(n7449), .ZN(n7839) );
  AOI21_X1 U9070 ( .B1(n7450), .B2(n7449), .A(n7839), .ZN(n7460) );
  AOI22_X1 U9071 ( .A1(n7845), .A2(P2_REG1_REG_14__SCAN_IN), .B1(n6120), .B2(
        n7840), .ZN(n7454) );
  OAI21_X1 U9072 ( .B1(n7452), .B2(P2_REG1_REG_13__SCAN_IN), .A(n7451), .ZN(
        n7453) );
  NAND2_X1 U9073 ( .A1(n7454), .A2(n7453), .ZN(n7844) );
  OAI21_X1 U9074 ( .B1(n7454), .B2(n7453), .A(n7844), .ZN(n7455) );
  NAND2_X1 U9075 ( .A1(n7455), .A2(n10056), .ZN(n7459) );
  INV_X1 U9076 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n7456) );
  NAND2_X1 U9077 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3152), .ZN(n8177) );
  OAI21_X1 U9078 ( .B1(n8460), .B2(n7456), .A(n8177), .ZN(n7457) );
  AOI21_X1 U9079 ( .B1(n9753), .B2(n7845), .A(n7457), .ZN(n7458) );
  OAI211_X1 U9080 ( .C1(n7460), .C2(n7850), .A(n7459), .B(n7458), .ZN(P2_U3259) );
  INV_X1 U9081 ( .A(n7461), .ZN(n7464) );
  INV_X1 U9082 ( .A(n7618), .ZN(n7463) );
  AOI21_X1 U9083 ( .B1(n7464), .B2(n7463), .A(n4966), .ZN(n7610) );
  NAND2_X1 U9084 ( .A1(n7610), .A2(n7609), .ZN(n7608) );
  NAND2_X1 U9085 ( .A1(n7477), .A2(n10019), .ZN(n7465) );
  NAND2_X1 U9086 ( .A1(n7608), .A2(n7465), .ZN(n7496) );
  XNOR2_X1 U9087 ( .A(n7496), .B(n7495), .ZN(n10029) );
  INV_X1 U9088 ( .A(n10029), .ZN(n7486) );
  NAND2_X1 U9089 ( .A1(n7467), .A2(n7466), .ZN(n7468) );
  NOR2_X1 U9090 ( .A1(n9321), .A2(n7468), .ZN(n9109) );
  NAND2_X1 U9091 ( .A1(n7470), .A2(n7469), .ZN(n7472) );
  NAND2_X1 U9092 ( .A1(n7472), .A2(n7471), .ZN(n7475) );
  INV_X1 U9093 ( .A(n7475), .ZN(n7473) );
  INV_X1 U9094 ( .A(n7499), .ZN(n7474) );
  AOI21_X1 U9095 ( .B1(n7495), .B2(n7475), .A(n7474), .ZN(n7476) );
  OAI222_X1 U9096 ( .A1(n9960), .A2(n9958), .B1(n9959), .B2(n7477), .C1(n9844), 
        .C2(n7476), .ZN(n10027) );
  INV_X1 U9097 ( .A(n7613), .ZN(n7478) );
  INV_X1 U9098 ( .A(n7504), .ZN(n7505) );
  OAI211_X1 U9099 ( .C1(n10026), .C2(n7478), .A(n7505), .B(n10011), .ZN(n10025) );
  NOR2_X1 U9100 ( .A1(n7479), .A2(n9250), .ZN(n9301) );
  INV_X1 U9101 ( .A(n9301), .ZN(n9272) );
  AOI22_X1 U9102 ( .A1(n9321), .A2(P1_REG2_REG_7__SCAN_IN), .B1(n9969), .B2(
        n7480), .ZN(n7483) );
  NAND2_X1 U9103 ( .A1(n9848), .A2(n7481), .ZN(n7482) );
  OAI211_X1 U9104 ( .C1(n10025), .C2(n9272), .A(n7483), .B(n7482), .ZN(n7484)
         );
  AOI21_X1 U9105 ( .B1(n10027), .B2(n9836), .A(n7484), .ZN(n7485) );
  OAI21_X1 U9106 ( .B1(n7486), .B2(n9308), .A(n7485), .ZN(P1_U3284) );
  XNOR2_X1 U9107 ( .A(n7488), .B(n7487), .ZN(n7492) );
  OAI22_X1 U9108 ( .A1(n8317), .A2(n10080), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6028), .ZN(n7490) );
  INV_X1 U9109 ( .A(n8347), .ZN(n10071) );
  OAI22_X1 U9110 ( .A1(n10157), .A2(n8337), .B1(n8331), .B2(n10071), .ZN(n7489) );
  AOI211_X1 U9111 ( .C1(n8307), .C2(n8349), .A(n7490), .B(n7489), .ZN(n7491)
         );
  OAI21_X1 U9112 ( .B1(n7492), .B2(n8321), .A(n7491), .ZN(P2_U3215) );
  INV_X1 U9113 ( .A(n7493), .ZN(n8060) );
  OAI222_X1 U9114 ( .A1(n9449), .A2(n9604), .B1(P1_U3084), .B2(n7494), .C1(
        n9445), .C2(n8060), .ZN(P1_U3333) );
  INV_X1 U9115 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n7509) );
  NAND2_X1 U9116 ( .A1(n7623), .A2(n10026), .ZN(n7497) );
  XNOR2_X1 U9117 ( .A(n7632), .B(n7500), .ZN(n7548) );
  INV_X1 U9118 ( .A(n7548), .ZN(n7507) );
  XNOR2_X1 U9119 ( .A(n7638), .B(n7500), .ZN(n7502) );
  AOI22_X1 U9120 ( .A1(n9287), .A2(n9013), .B1(n9285), .B2(n9011), .ZN(n7501)
         );
  OAI21_X1 U9121 ( .B1(n7502), .B2(n9844), .A(n7501), .ZN(n7503) );
  AOI21_X1 U9122 ( .B1(n7548), .B2(n9846), .A(n7503), .ZN(n7550) );
  AOI21_X1 U9123 ( .B1(n7633), .B2(n7505), .A(n9950), .ZN(n7542) );
  AOI22_X1 U9124 ( .A1(n7542), .A2(n10011), .B1(n10010), .B2(n7633), .ZN(n7506) );
  OAI211_X1 U9125 ( .C1(n7507), .C2(n10015), .A(n7550), .B(n7506), .ZN(n7530)
         );
  NAND2_X1 U9126 ( .A1(n7530), .A2(n10042), .ZN(n7508) );
  OAI21_X1 U9127 ( .B1(n10042), .B2(n7509), .A(n7508), .ZN(P1_U3478) );
  OAI21_X1 U9128 ( .B1(n7512), .B2(n7511), .A(n7510), .ZN(n10001) );
  NAND2_X1 U9129 ( .A1(n10001), .A2(n9846), .ZN(n7517) );
  OAI22_X1 U9130 ( .A1(n7514), .A2(n9960), .B1(n9959), .B2(n7513), .ZN(n7515)
         );
  INV_X1 U9131 ( .A(n7515), .ZN(n7516) );
  OAI211_X1 U9132 ( .C1(n9844), .C2(n7518), .A(n7517), .B(n7516), .ZN(n9999)
         );
  MUX2_X1 U9133 ( .A(n9999), .B(P1_REG2_REG_2__SCAN_IN), .S(n9970), .Z(n7519)
         );
  INV_X1 U9134 ( .A(n7519), .ZN(n7529) );
  AND2_X1 U9135 ( .A1(n10001), .A2(n9953), .ZN(n7527) );
  OAI21_X1 U9136 ( .B1(n7522), .B2(n7521), .A(n7520), .ZN(n7523) );
  AND2_X1 U9137 ( .A1(n7563), .A2(n7523), .ZN(n9996) );
  NAND2_X1 U9138 ( .A1(n9952), .A2(n9996), .ZN(n7525) );
  NAND2_X1 U9139 ( .A1(n9969), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n7524) );
  OAI211_X1 U9140 ( .C1(n9972), .C2(n9997), .A(n7525), .B(n7524), .ZN(n7526)
         );
  NOR2_X1 U9141 ( .A1(n7527), .A2(n7526), .ZN(n7528) );
  NAND2_X1 U9142 ( .A1(n7529), .A2(n7528), .ZN(P1_U3289) );
  INV_X1 U9143 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n7532) );
  NAND2_X1 U9144 ( .A1(n7530), .A2(n4392), .ZN(n7531) );
  OAI21_X1 U9145 ( .B1(n4392), .B2(n7532), .A(n7531), .ZN(P1_U3531) );
  AOI22_X1 U9146 ( .A1(n7534), .A2(n9086), .B1(n9969), .B2(n7533), .ZN(n7535)
         );
  AOI21_X1 U9147 ( .B1(n7536), .B2(n7535), .A(n9321), .ZN(n7541) );
  NOR2_X1 U9148 ( .A1(n7537), .A2(n9308), .ZN(n7540) );
  OAI22_X1 U9149 ( .A1(n9972), .A2(n7538), .B1(n6843), .B2(n9836), .ZN(n7539)
         );
  OR3_X1 U9150 ( .A1(n7541), .A2(n7540), .A3(n7539), .ZN(P1_U3286) );
  NAND2_X1 U9151 ( .A1(n7542), .A2(n9952), .ZN(n7545) );
  AOI22_X1 U9152 ( .A1(n9970), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n9969), .B2(
        n7543), .ZN(n7544) );
  OAI211_X1 U9153 ( .C1(n7546), .C2(n9972), .A(n7545), .B(n7544), .ZN(n7547)
         );
  AOI21_X1 U9154 ( .B1(n7548), .B2(n9953), .A(n7547), .ZN(n7549) );
  OAI21_X1 U9155 ( .B1(n7550), .B2(n9321), .A(n7549), .ZN(P1_U3283) );
  INV_X1 U9156 ( .A(n7551), .ZN(n7572) );
  OAI222_X1 U9157 ( .A1(n8124), .A2(n7553), .B1(n8859), .B2(n7572), .C1(n7552), 
        .C2(P2_U3152), .ZN(P2_U3337) );
  XOR2_X1 U9158 ( .A(n7556), .B(n7554), .Z(n7562) );
  XOR2_X1 U9159 ( .A(n7556), .B(n7555), .Z(n7560) );
  OAI22_X1 U9160 ( .A1(n7558), .A2(n9960), .B1(n9959), .B2(n7557), .ZN(n7559)
         );
  AOI21_X1 U9161 ( .B1(n7560), .B2(n9963), .A(n7559), .ZN(n7561) );
  OAI21_X1 U9162 ( .B1(n7562), .B2(n9966), .A(n7561), .ZN(n10005) );
  INV_X1 U9163 ( .A(n10005), .ZN(n7571) );
  INV_X1 U9164 ( .A(n7562), .ZN(n10007) );
  INV_X1 U9165 ( .A(n9952), .ZN(n9324) );
  INV_X1 U9166 ( .A(n7563), .ZN(n7565) );
  OAI21_X1 U9167 ( .B1(n7565), .B2(n10003), .A(n7564), .ZN(n10004) );
  AOI22_X1 U9168 ( .A1(n9321), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n9969), .B2(
        n5392), .ZN(n7568) );
  NAND2_X1 U9169 ( .A1(n9848), .A2(n7566), .ZN(n7567) );
  OAI211_X1 U9170 ( .C1(n9324), .C2(n10004), .A(n7568), .B(n7567), .ZN(n7569)
         );
  AOI21_X1 U9171 ( .B1(n10007), .B2(n9953), .A(n7569), .ZN(n7570) );
  OAI21_X1 U9172 ( .B1(n7571), .B2(n9321), .A(n7570), .ZN(P1_U3288) );
  OAI222_X1 U9173 ( .A1(n9449), .A2(n9556), .B1(P1_U3084), .B2(n7573), .C1(
        n9445), .C2(n7572), .ZN(P1_U3332) );
  NAND2_X1 U9174 ( .A1(n7576), .A2(n7575), .ZN(n7577) );
  XNOR2_X1 U9175 ( .A(n7574), .B(n7577), .ZN(n7583) );
  NAND2_X1 U9176 ( .A1(n8992), .A2(n7648), .ZN(n7580) );
  AOI21_X1 U9177 ( .B1(n8979), .B2(n9011), .A(n7578), .ZN(n7579) );
  OAI211_X1 U9178 ( .C1(n7989), .C2(n8972), .A(n7580), .B(n7579), .ZN(n7581)
         );
  AOI21_X1 U9179 ( .B1(n7868), .B2(n8997), .A(n7581), .ZN(n7582) );
  OAI21_X1 U9180 ( .B1(n7583), .B2(n8999), .A(n7582), .ZN(P1_U3215) );
  INV_X1 U9181 ( .A(n7585), .ZN(n7586) );
  AOI21_X1 U9182 ( .B1(n7587), .B2(n7584), .A(n7586), .ZN(n7592) );
  AND2_X1 U9183 ( .A1(P1_U3084), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n9918) );
  AOI21_X1 U9184 ( .B1(n8991), .B2(n9010), .A(n9918), .ZN(n7589) );
  NAND2_X1 U9185 ( .A1(n8992), .A2(n9968), .ZN(n7588) );
  OAI211_X1 U9186 ( .C1(n9958), .C2(n8995), .A(n7589), .B(n7588), .ZN(n7590)
         );
  AOI21_X1 U9187 ( .B1(n7647), .B2(n8997), .A(n7590), .ZN(n7591) );
  OAI21_X1 U9188 ( .B1(n7592), .B2(n8999), .A(n7591), .ZN(P1_U3229) );
  INV_X1 U9189 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n7607) );
  NOR2_X1 U9190 ( .A1(n9731), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n7593) );
  AOI21_X1 U9191 ( .B1(P1_REG1_REG_14__SCAN_IN), .B2(n9731), .A(n7593), .ZN(
        n7596) );
  OAI21_X1 U9192 ( .B1(n7600), .B2(P1_REG1_REG_13__SCAN_IN), .A(n7594), .ZN(
        n7595) );
  NAND2_X1 U9193 ( .A1(n7596), .A2(n7595), .ZN(n7907) );
  OAI21_X1 U9194 ( .B1(n7596), .B2(n7595), .A(n7907), .ZN(n7605) );
  INV_X1 U9195 ( .A(n9731), .ZN(n7914) );
  NOR2_X1 U9196 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7597), .ZN(n8875) );
  INV_X1 U9197 ( .A(n8875), .ZN(n7598) );
  OAI21_X1 U9198 ( .B1(n9922), .B2(n7914), .A(n7598), .ZN(n7604) );
  XNOR2_X1 U9199 ( .A(n7914), .B(n7915), .ZN(n7602) );
  INV_X1 U9200 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n7601) );
  NOR2_X1 U9201 ( .A1(n7601), .A2(n7602), .ZN(n7916) );
  AOI211_X1 U9202 ( .C1(n7602), .C2(n7601), .A(n7916), .B(n9886), .ZN(n7603)
         );
  AOI211_X1 U9203 ( .C1(n9938), .C2(n7605), .A(n7604), .B(n7603), .ZN(n7606)
         );
  OAI21_X1 U9204 ( .B1(n9945), .B2(n7607), .A(n7606), .ZN(P1_U3255) );
  OAI21_X1 U9205 ( .B1(n7610), .B2(n7609), .A(n7608), .ZN(n10023) );
  NAND2_X1 U9206 ( .A1(n7611), .A2(n7615), .ZN(n7612) );
  NAND2_X1 U9207 ( .A1(n7613), .A2(n7612), .ZN(n10020) );
  AOI22_X1 U9208 ( .A1(n9848), .A2(n7615), .B1(n7614), .B2(n9969), .ZN(n7616)
         );
  OAI21_X1 U9209 ( .B1(n9324), .B2(n10020), .A(n7616), .ZN(n7629) );
  AOI21_X1 U9210 ( .B1(n7619), .B2(n7618), .A(n7617), .ZN(n7621) );
  XNOR2_X1 U9211 ( .A(n7621), .B(n7620), .ZN(n7627) );
  NAND2_X1 U9212 ( .A1(n10023), .A2(n9846), .ZN(n7626) );
  OAI22_X1 U9213 ( .A1(n7623), .A2(n9960), .B1(n9959), .B2(n7622), .ZN(n7624)
         );
  INV_X1 U9214 ( .A(n7624), .ZN(n7625) );
  OAI211_X1 U9215 ( .C1(n9844), .C2(n7627), .A(n7626), .B(n7625), .ZN(n10021)
         );
  MUX2_X1 U9216 ( .A(n10021), .B(P1_REG2_REG_6__SCAN_IN), .S(n9970), .Z(n7628)
         );
  AOI211_X1 U9217 ( .C1(n9953), .C2(n10023), .A(n7629), .B(n7628), .ZN(n7630)
         );
  INV_X1 U9218 ( .A(n7630), .ZN(P1_U3285) );
  NAND2_X1 U9219 ( .A1(n9012), .A2(n7633), .ZN(n9946) );
  NAND2_X1 U9220 ( .A1(n7647), .A2(n9011), .ZN(n7634) );
  AND2_X1 U9221 ( .A1(n9946), .A2(n7634), .ZN(n7635) );
  INV_X1 U9222 ( .A(n7870), .ZN(n7636) );
  AOI21_X1 U9223 ( .B1(n7643), .B2(n7637), .A(n7636), .ZN(n7799) );
  INV_X1 U9224 ( .A(n7640), .ZN(n7641) );
  AOI21_X1 U9225 ( .B1(n9955), .B2(n7642), .A(n7641), .ZN(n7644) );
  XNOR2_X1 U9226 ( .A(n7644), .B(n7643), .ZN(n7646) );
  OAI222_X1 U9227 ( .A1(n9960), .A2(n7989), .B1(n7646), .B2(n9844), .C1(n9959), 
        .C2(n7645), .ZN(n7796) );
  INV_X1 U9228 ( .A(n7868), .ZN(n7651) );
  INV_X1 U9229 ( .A(n7647), .ZN(n10033) );
  NAND2_X1 U9230 ( .A1(n9950), .A2(n10033), .ZN(n9949) );
  INV_X1 U9231 ( .A(n7883), .ZN(n9852) );
  AOI211_X1 U9232 ( .C1(n7868), .C2(n9949), .A(n10034), .B(n9852), .ZN(n7797)
         );
  NAND2_X1 U9233 ( .A1(n7797), .A2(n9301), .ZN(n7650) );
  AOI22_X1 U9234 ( .A1(n9970), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n9969), .B2(
        n7648), .ZN(n7649) );
  OAI211_X1 U9235 ( .C1(n7651), .C2(n9972), .A(n7650), .B(n7649), .ZN(n7652)
         );
  AOI21_X1 U9236 ( .B1(n7796), .B2(n9836), .A(n7652), .ZN(n7653) );
  OAI21_X1 U9237 ( .B1(n7799), .B2(n9308), .A(n7653), .ZN(P1_U3281) );
  XNOR2_X1 U9238 ( .A(n7655), .B(n7654), .ZN(n7660) );
  OAI21_X1 U9239 ( .B1(n8317), .B2(n7689), .A(n7656), .ZN(n7658) );
  OAI22_X1 U9240 ( .A1(n10165), .A2(n8337), .B1(n8331), .B2(n7834), .ZN(n7657)
         );
  AOI211_X1 U9241 ( .C1(n8307), .C2(n8348), .A(n7658), .B(n7657), .ZN(n7659)
         );
  OAI21_X1 U9242 ( .B1(n7660), .B2(n8321), .A(n7659), .ZN(P2_U3223) );
  INV_X1 U9243 ( .A(n7661), .ZN(n8062) );
  OAI222_X1 U9244 ( .A1(n8124), .A2(n7663), .B1(n8859), .B2(n8062), .C1(
        P2_U3152), .C2(n7662), .ZN(P2_U3336) );
  NOR2_X1 U9245 ( .A1(n8350), .A2(n7785), .ZN(n7664) );
  NAND2_X1 U9246 ( .A1(n7666), .A2(n7785), .ZN(n7667) );
  AND2_X1 U9247 ( .A1(n8349), .A2(n8303), .ZN(n7668) );
  NAND2_X1 U9248 ( .A1(n10078), .A2(n10077), .ZN(n7670) );
  INV_X1 U9249 ( .A(n10157), .ZN(n10083) );
  OR2_X1 U9250 ( .A1(n8348), .A2(n10083), .ZN(n7669) );
  NAND2_X1 U9251 ( .A1(n7670), .A2(n7669), .ZN(n7672) );
  INV_X1 U9252 ( .A(n7672), .ZN(n7671) );
  NAND2_X1 U9253 ( .A1(n7672), .A2(n7684), .ZN(n7673) );
  NAND2_X1 U9254 ( .A1(n7700), .A2(n7673), .ZN(n10164) );
  AND3_X1 U9255 ( .A1(n7675), .A2(P2_STATE_REG_SCAN_IN), .A3(n7674), .ZN(n7677) );
  AND2_X1 U9256 ( .A1(n7677), .A2(n7676), .ZN(n7678) );
  NAND2_X1 U9257 ( .A1(n7679), .A2(n7678), .ZN(n7693) );
  OR2_X1 U9258 ( .A1(n7680), .A2(n8668), .ZN(n7734) );
  INV_X1 U9259 ( .A(n7734), .ZN(n7681) );
  NAND2_X1 U9260 ( .A1(n8749), .A2(n7681), .ZN(n8730) );
  OAI21_X1 U9261 ( .B1(n7684), .B2(n7683), .A(n7682), .ZN(n7685) );
  NAND2_X1 U9262 ( .A1(n7685), .A2(n8722), .ZN(n7687) );
  AOI22_X1 U9263 ( .A1(n8346), .A2(n8686), .B1(n8684), .B2(n8348), .ZN(n7686)
         );
  OAI211_X1 U9264 ( .C1(n10164), .C2(n8717), .A(n7687), .B(n7686), .ZN(n10167)
         );
  NAND2_X1 U9265 ( .A1(n10167), .A2(n8749), .ZN(n7697) );
  OAI22_X1 U9266 ( .A1(n10081), .A2(n7690), .B1(n7689), .B2(n10096), .ZN(n7695) );
  NAND2_X1 U9267 ( .A1(n7691), .A2(n7698), .ZN(n7692) );
  NAND2_X1 U9268 ( .A1(n7712), .A2(n7692), .ZN(n10166) );
  OR2_X1 U9269 ( .A1(n7693), .A2(n6322), .ZN(n10098) );
  INV_X1 U9270 ( .A(n10098), .ZN(n8709) );
  NAND2_X1 U9271 ( .A1(n8709), .A2(n10126), .ZN(n10085) );
  NOR2_X1 U9272 ( .A1(n10166), .A2(n10085), .ZN(n7694) );
  AOI211_X1 U9273 ( .C1(n10102), .C2(n7698), .A(n7695), .B(n7694), .ZN(n7696)
         );
  OAI211_X1 U9274 ( .C1(n10164), .C2(n8730), .A(n7697), .B(n7696), .ZN(
        P2_U3288) );
  NAND2_X1 U9275 ( .A1(n8347), .A2(n7698), .ZN(n7699) );
  INV_X1 U9276 ( .A(n7807), .ZN(n7702) );
  AOI21_X1 U9277 ( .B1(n7704), .B2(n7703), .A(n7702), .ZN(n10170) );
  AOI22_X1 U9278 ( .A1(n8345), .A2(n8686), .B1(n8684), .B2(n8347), .ZN(n7710)
         );
  INV_X1 U9279 ( .A(n7682), .ZN(n7706) );
  NOR3_X1 U9280 ( .A1(n7706), .A2(n7705), .A3(n7704), .ZN(n7708) );
  OAI21_X1 U9281 ( .B1(n7708), .B2(n7707), .A(n8722), .ZN(n7709) );
  OAI211_X1 U9282 ( .C1(n10170), .C2(n8717), .A(n7710), .B(n7709), .ZN(n10173)
         );
  NAND2_X1 U9283 ( .A1(n10173), .A2(n8749), .ZN(n7717) );
  OAI22_X1 U9284 ( .A1(n10081), .A2(n7711), .B1(n7824), .B2(n10096), .ZN(n7715) );
  NAND2_X1 U9285 ( .A1(n7712), .A2(n7805), .ZN(n7713) );
  NAND2_X1 U9286 ( .A1(n7814), .A2(n7713), .ZN(n10172) );
  NOR2_X1 U9287 ( .A1(n10172), .A2(n10085), .ZN(n7714) );
  AOI211_X1 U9288 ( .C1(n10102), .C2(n7805), .A(n7715), .B(n7714), .ZN(n7716)
         );
  OAI211_X1 U9289 ( .C1(n10170), .C2(n8730), .A(n7717), .B(n7716), .ZN(
        P2_U3287) );
  INV_X1 U9290 ( .A(n7729), .ZN(n7720) );
  AOI21_X1 U9291 ( .B1(P1_DATAO_REG_23__SCAN_IN), .B2(n8856), .A(n7718), .ZN(
        n7719) );
  OAI21_X1 U9292 ( .B1(n7720), .B2(n8859), .A(n7719), .ZN(P2_U3335) );
  INV_X1 U9293 ( .A(n9849), .ZN(n9869) );
  AOI21_X1 U9294 ( .B1(n7722), .B2(n7721), .A(n8999), .ZN(n7724) );
  NAND2_X1 U9295 ( .A1(n7724), .A2(n7723), .ZN(n7728) );
  NOR2_X1 U9296 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n5538), .ZN(n9929) );
  AOI21_X1 U9297 ( .B1(n8991), .B2(n9008), .A(n9929), .ZN(n7725) );
  OAI21_X1 U9298 ( .B1(n9961), .B2(n8995), .A(n7725), .ZN(n7726) );
  AOI21_X1 U9299 ( .B1(n9847), .B2(n8992), .A(n7726), .ZN(n7727) );
  OAI211_X1 U9300 ( .C1(n9869), .C2(n8985), .A(n7728), .B(n7727), .ZN(P1_U3234) );
  NAND2_X1 U9301 ( .A1(n7729), .A2(n9732), .ZN(n7731) );
  OAI211_X1 U9302 ( .C1(n7732), .C2(n9449), .A(n7731), .B(n7730), .ZN(P1_U3330) );
  XOR2_X1 U9303 ( .A(n7736), .B(n7733), .Z(n10155) );
  INV_X1 U9304 ( .A(n10155), .ZN(n7748) );
  NAND2_X1 U9305 ( .A1(n8717), .A2(n7734), .ZN(n7735) );
  INV_X1 U9306 ( .A(n8348), .ZN(n7741) );
  NOR2_X1 U9307 ( .A1(n4504), .A2(n7737), .ZN(n7739) );
  AOI21_X1 U9308 ( .B1(n7739), .B2(n7738), .A(n10069), .ZN(n7740) );
  OAI222_X1 U9309 ( .A1(n10070), .A2(n7741), .B1(n10072), .B2(n4692), .C1(
        n10089), .C2(n7740), .ZN(n10153) );
  NAND2_X1 U9310 ( .A1(n10153), .A2(n8749), .ZN(n7747) );
  OAI22_X1 U9311 ( .A1(n10096), .A2(n8305), .B1(n6948), .B2(n10081), .ZN(n7745) );
  INV_X1 U9312 ( .A(n10079), .ZN(n7742) );
  OAI21_X1 U9313 ( .B1(n10151), .B2(n7743), .A(n7742), .ZN(n10152) );
  NOR2_X1 U9314 ( .A1(n10152), .A2(n10085), .ZN(n7744) );
  AOI211_X1 U9315 ( .C1(n10102), .C2(n8303), .A(n7745), .B(n7744), .ZN(n7746)
         );
  OAI211_X1 U9316 ( .C1(n7748), .C2(n8751), .A(n7747), .B(n7746), .ZN(P2_U3290) );
  XNOR2_X1 U9317 ( .A(n7749), .B(n7750), .ZN(n10144) );
  INV_X1 U9318 ( .A(n10144), .ZN(n7765) );
  INV_X1 U9319 ( .A(n7750), .ZN(n7753) );
  INV_X1 U9320 ( .A(n7751), .ZN(n7752) );
  NOR2_X1 U9321 ( .A1(n7753), .A2(n7752), .ZN(n7756) );
  AOI21_X1 U9322 ( .B1(n7756), .B2(n7754), .A(n7755), .ZN(n7757) );
  OAI222_X1 U9323 ( .A1(n10070), .A2(n7759), .B1(n10072), .B2(n7758), .C1(
        n10089), .C2(n7757), .ZN(n10142) );
  NAND2_X1 U9324 ( .A1(n10142), .A2(n8749), .ZN(n7764) );
  NOR2_X1 U9325 ( .A1(n8749), .A2(n6951), .ZN(n7761) );
  OAI211_X1 U9326 ( .C1(n7900), .C2(n10141), .A(n10126), .B(n10093), .ZN(
        n10140) );
  OAI22_X1 U9327 ( .A1(n10098), .A2(n10140), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        n10096), .ZN(n7760) );
  AOI211_X1 U9328 ( .C1(n10102), .C2(n7762), .A(n7761), .B(n7760), .ZN(n7763)
         );
  OAI211_X1 U9329 ( .C1(n7765), .C2(n8751), .A(n7764), .B(n7763), .ZN(P2_U3293) );
  INV_X1 U9330 ( .A(n7766), .ZN(n7767) );
  AOI21_X1 U9331 ( .B1(n7769), .B2(n7768), .A(n7767), .ZN(n10131) );
  AOI21_X1 U9332 ( .B1(n7792), .B2(n4942), .A(n7899), .ZN(n10127) );
  OAI22_X1 U9333 ( .A1(n10081), .A2(n6953), .B1(n7770), .B2(n10096), .ZN(n7771) );
  AOI21_X1 U9334 ( .B1(n8727), .B2(n10127), .A(n7771), .ZN(n7778) );
  XNOR2_X1 U9335 ( .A(n7773), .B(n7772), .ZN(n7774) );
  NAND2_X1 U9336 ( .A1(n7774), .A2(n8722), .ZN(n7776) );
  AOI22_X1 U9337 ( .A1(n8684), .A2(n5990), .B1(n6725), .B2(n8686), .ZN(n7775)
         );
  NAND2_X1 U9338 ( .A1(n7776), .A2(n7775), .ZN(n10132) );
  AOI22_X1 U9339 ( .A1(n10102), .A2(n4942), .B1(n10081), .B2(n10132), .ZN(
        n7777) );
  OAI211_X1 U9340 ( .C1(n10131), .C2(n8751), .A(n7778), .B(n7777), .ZN(
        P2_U3295) );
  MUX2_X1 U9341 ( .A(n7780), .B(n7779), .S(n10081), .Z(n7787) );
  INV_X1 U9342 ( .A(n7781), .ZN(n7783) );
  OAI22_X1 U9343 ( .A1(n7783), .A2(n10098), .B1(n7782), .B2(n10096), .ZN(n7784) );
  AOI21_X1 U9344 ( .B1(n10102), .B2(n7785), .A(n7784), .ZN(n7786) );
  OAI211_X1 U9345 ( .C1(n7788), .C2(n8751), .A(n7787), .B(n7786), .ZN(P2_U3291) );
  INV_X1 U9346 ( .A(n10125), .ZN(n7795) );
  AND2_X1 U9347 ( .A1(n6718), .A2(n8686), .ZN(n7789) );
  AOI21_X1 U9348 ( .B1(n8722), .B2(n10125), .A(n7789), .ZN(n10121) );
  OAI22_X1 U9349 ( .A1(n10108), .A2(n10121), .B1(n7790), .B2(n10096), .ZN(
        n7791) );
  AOI21_X1 U9350 ( .B1(P2_REG2_REG_0__SCAN_IN), .B2(n10104), .A(n7791), .ZN(
        n7794) );
  OAI21_X1 U9351 ( .B1(n8727), .B2(n10102), .A(n7792), .ZN(n7793) );
  OAI211_X1 U9352 ( .C1(n7795), .C2(n8751), .A(n7794), .B(n7793), .ZN(P2_U3296) );
  INV_X1 U9353 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n7801) );
  AOI211_X1 U9354 ( .C1(n10010), .C2(n7868), .A(n7797), .B(n7796), .ZN(n7798)
         );
  OAI21_X1 U9355 ( .B1(n7799), .B2(n9418), .A(n7798), .ZN(n7802) );
  NAND2_X1 U9356 ( .A1(n7802), .A2(n10042), .ZN(n7800) );
  OAI21_X1 U9357 ( .B1(n10042), .B2(n7801), .A(n7800), .ZN(P1_U3484) );
  NAND2_X1 U9358 ( .A1(n7802), .A2(n4392), .ZN(n7803) );
  OAI21_X1 U9359 ( .B1(n4392), .B2(n7804), .A(n7803), .ZN(P1_U3533) );
  OR2_X1 U9360 ( .A1(n8346), .A2(n7805), .ZN(n7806) );
  OAI21_X1 U9361 ( .B1(n7808), .B2(n7809), .A(n7853), .ZN(n10177) );
  XNOR2_X1 U9362 ( .A(n4472), .B(n7809), .ZN(n7811) );
  OAI22_X1 U9363 ( .A1(n7834), .A2(n10072), .B1(n8020), .B2(n10070), .ZN(n7810) );
  AOI21_X1 U9364 ( .B1(n7811), .B2(n8722), .A(n7810), .ZN(n7812) );
  OAI21_X1 U9365 ( .B1(n8717), .B2(n10177), .A(n7812), .ZN(n10181) );
  NAND2_X1 U9366 ( .A1(n10181), .A2(n8749), .ZN(n7819) );
  OAI22_X1 U9367 ( .A1(n10081), .A2(n7813), .B1(n7833), .B2(n10096), .ZN(n7817) );
  AND2_X1 U9368 ( .A1(n7814), .A2(n10178), .ZN(n7815) );
  OR2_X1 U9369 ( .A1(n7815), .A2(n7931), .ZN(n10180) );
  NOR2_X1 U9370 ( .A1(n10180), .A2(n10085), .ZN(n7816) );
  AOI211_X1 U9371 ( .C1(n10102), .C2(n10178), .A(n7817), .B(n7816), .ZN(n7818)
         );
  OAI211_X1 U9372 ( .C1(n10177), .C2(n8730), .A(n7819), .B(n7818), .ZN(
        P2_U3286) );
  OAI21_X1 U9373 ( .B1(n7822), .B2(n7821), .A(n7820), .ZN(n7823) );
  NAND2_X1 U9374 ( .A1(n7823), .A2(n8325), .ZN(n7829) );
  INV_X1 U9375 ( .A(n7824), .ZN(n7827) );
  OAI22_X1 U9376 ( .A1(n10071), .A2(n8330), .B1(n8331), .B2(n7947), .ZN(n7825)
         );
  AOI211_X1 U9377 ( .C1(n7827), .C2(n8334), .A(n7826), .B(n7825), .ZN(n7828)
         );
  OAI211_X1 U9378 ( .C1(n10171), .C2(n8337), .A(n7829), .B(n7828), .ZN(
        P2_U3233) );
  XNOR2_X1 U9379 ( .A(n7831), .B(n7830), .ZN(n7838) );
  OAI21_X1 U9380 ( .B1(n8317), .B2(n7833), .A(n7832), .ZN(n7836) );
  OAI22_X1 U9381 ( .A1(n7834), .A2(n8330), .B1(n8331), .B2(n8020), .ZN(n7835)
         );
  AOI211_X1 U9382 ( .C1(n10178), .C2(n8319), .A(n7836), .B(n7835), .ZN(n7837)
         );
  OAI21_X1 U9383 ( .B1(n7838), .B2(n8321), .A(n7837), .ZN(P2_U3219) );
  AOI21_X1 U9384 ( .B1(n7840), .B2(n6124), .A(n7839), .ZN(n8403) );
  XNOR2_X1 U9385 ( .A(n8403), .B(n8404), .ZN(n7841) );
  NOR2_X1 U9386 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n7841), .ZN(n8405) );
  AOI21_X1 U9387 ( .B1(n7841), .B2(P2_REG2_REG_15__SCAN_IN), .A(n8405), .ZN(
        n7851) );
  INV_X1 U9388 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n7843) );
  AND2_X1 U9389 ( .A1(P2_REG3_REG_15__SCAN_IN), .A2(P2_U3152), .ZN(n8333) );
  INV_X1 U9390 ( .A(n8333), .ZN(n7842) );
  OAI21_X1 U9391 ( .B1(n8460), .B2(n7843), .A(n7842), .ZN(n7848) );
  INV_X1 U9392 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n9801) );
  AOI211_X1 U9393 ( .C1(n7846), .C2(n9801), .A(n8395), .B(n10060), .ZN(n7847)
         );
  AOI211_X1 U9394 ( .C1(n9753), .C2(n8404), .A(n7848), .B(n7847), .ZN(n7849)
         );
  OAI21_X1 U9395 ( .B1(n7851), .B2(n7850), .A(n7849), .ZN(P2_U3260) );
  NAND2_X1 U9396 ( .A1(n10178), .A2(n8345), .ZN(n7852) );
  NAND2_X1 U9397 ( .A1(n7853), .A2(n7852), .ZN(n7928) );
  NAND2_X1 U9398 ( .A1(n7950), .A2(n8344), .ZN(n7854) );
  AND2_X1 U9399 ( .A1(n7930), .A2(n7854), .ZN(n7856) );
  AND2_X1 U9400 ( .A1(n7854), .A2(n4412), .ZN(n7855) );
  OAI21_X1 U9401 ( .B1(n7856), .B2(n4412), .A(n7995), .ZN(n10198) );
  INV_X1 U9402 ( .A(n10198), .ZN(n7867) );
  INV_X1 U9403 ( .A(n7857), .ZN(n7858) );
  NOR2_X1 U9404 ( .A1(n7859), .A2(n7858), .ZN(n7860) );
  XNOR2_X1 U9405 ( .A(n7860), .B(n4412), .ZN(n7861) );
  OAI222_X1 U9406 ( .A1(n10072), .A2(n8020), .B1(n10070), .B2(n8179), .C1(
        n10089), .C2(n7861), .ZN(n10196) );
  INV_X1 U9407 ( .A(n8023), .ZN(n10193) );
  INV_X1 U9408 ( .A(n7950), .ZN(n10188) );
  INV_X1 U9409 ( .A(n8004), .ZN(n7862) );
  OAI21_X1 U9410 ( .B1(n10193), .B2(n7933), .A(n7862), .ZN(n10195) );
  OAI22_X1 U9411 ( .A1(n10081), .A2(n7332), .B1(n8019), .B2(n10096), .ZN(n7863) );
  AOI21_X1 U9412 ( .B1(n10102), .B2(n8023), .A(n7863), .ZN(n7864) );
  OAI21_X1 U9413 ( .B1(n10195), .B2(n10085), .A(n7864), .ZN(n7865) );
  AOI21_X1 U9414 ( .B1(n10196), .B2(n8749), .A(n7865), .ZN(n7866) );
  OAI21_X1 U9415 ( .B1(n7867), .B2(n8751), .A(n7866), .ZN(P2_U3284) );
  OR2_X1 U9416 ( .A1(n7868), .A2(n9010), .ZN(n7869) );
  NAND2_X1 U9417 ( .A1(n7873), .A2(n7879), .ZN(n7954) );
  OR2_X1 U9418 ( .A1(n7873), .A2(n7879), .ZN(n7874) );
  NAND2_X1 U9419 ( .A1(n7954), .A2(n7874), .ZN(n9863) );
  AOI22_X1 U9420 ( .A1(n9287), .A2(n9009), .B1(n9285), .B2(n9007), .ZN(n7882)
         );
  OAI211_X1 U9421 ( .C1(n4967), .C2(n7880), .A(n7959), .B(n9963), .ZN(n7881)
         );
  OAI211_X1 U9422 ( .C1(n9863), .C2(n9966), .A(n7882), .B(n7881), .ZN(n9866)
         );
  NAND2_X1 U9423 ( .A1(n9866), .A2(n9836), .ZN(n7889) );
  INV_X1 U9424 ( .A(n7991), .ZN(n9865) );
  NOR2_X2 U9425 ( .A1(n7883), .A2(n9849), .ZN(n9850) );
  INV_X1 U9426 ( .A(n9821), .ZN(n7884) );
  OAI211_X1 U9427 ( .C1(n9865), .C2(n9850), .A(n7884), .B(n10011), .ZN(n9864)
         );
  INV_X1 U9428 ( .A(n9864), .ZN(n7887) );
  AOI22_X1 U9429 ( .A1(n9970), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n9969), .B2(
        n7986), .ZN(n7885) );
  OAI21_X1 U9430 ( .B1(n9865), .B2(n9972), .A(n7885), .ZN(n7886) );
  AOI21_X1 U9431 ( .B1(n7887), .B2(n9301), .A(n7886), .ZN(n7888) );
  OAI211_X1 U9432 ( .C1(n9863), .C2(n7890), .A(n7889), .B(n7888), .ZN(P1_U3279) );
  INV_X1 U9433 ( .A(n8751), .ZN(n10105) );
  OAI21_X1 U9434 ( .B1(n7893), .B2(n7892), .A(n7891), .ZN(n10139) );
  OAI21_X1 U9435 ( .B1(n7895), .B2(n7894), .A(n7754), .ZN(n7896) );
  NAND2_X1 U9436 ( .A1(n7896), .A2(n8722), .ZN(n7898) );
  AOI22_X1 U9437 ( .A1(n8686), .A2(n8352), .B1(n6718), .B2(n8684), .ZN(n7897)
         );
  NAND2_X1 U9438 ( .A1(n7898), .A2(n7897), .ZN(n10138) );
  MUX2_X1 U9439 ( .A(n10138), .B(P2_REG2_REG_2__SCAN_IN), .S(n10108), .Z(n7905) );
  INV_X1 U9440 ( .A(n7899), .ZN(n7901) );
  AOI211_X1 U9441 ( .C1(n7902), .C2(n7901), .A(n10194), .B(n7900), .ZN(n10134)
         );
  INV_X1 U9442 ( .A(n10096), .ZN(n8743) );
  AOI22_X1 U9443 ( .A1(n10134), .A2(n8709), .B1(P2_REG3_REG_2__SCAN_IN), .B2(
        n8743), .ZN(n7903) );
  OAI21_X1 U9444 ( .B1(n8703), .B2(n10136), .A(n7903), .ZN(n7904) );
  AOI211_X1 U9445 ( .C1(n10105), .C2(n10139), .A(n7905), .B(n7904), .ZN(n7906)
         );
  INV_X1 U9446 ( .A(n7906), .ZN(P2_U3294) );
  OAI21_X1 U9447 ( .B1(n9731), .B2(P1_REG1_REG_14__SCAN_IN), .A(n7907), .ZN(
        n9035) );
  XNOR2_X1 U9448 ( .A(n9036), .B(n9035), .ZN(n7908) );
  INV_X1 U9449 ( .A(n7908), .ZN(n7911) );
  INV_X1 U9450 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n7909) );
  NOR2_X1 U9451 ( .A1(n7909), .A2(n7908), .ZN(n9037) );
  INV_X1 U9452 ( .A(n9037), .ZN(n7910) );
  OAI211_X1 U9453 ( .C1(P1_REG1_REG_15__SCAN_IN), .C2(n7911), .A(n9938), .B(
        n7910), .ZN(n7913) );
  NOR2_X1 U9454 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n5348), .ZN(n8990) );
  INV_X1 U9455 ( .A(n8990), .ZN(n7912) );
  OAI211_X1 U9456 ( .C1(n9922), .C2(n9036), .A(n7913), .B(n7912), .ZN(n7921)
         );
  NOR2_X1 U9457 ( .A1(n7915), .A2(n7914), .ZN(n7917) );
  NOR2_X1 U9458 ( .A1(n7917), .A2(n7916), .ZN(n9030) );
  INV_X1 U9459 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n7918) );
  AOI211_X1 U9460 ( .C1(n7919), .C2(n7918), .A(n9031), .B(n9886), .ZN(n7920)
         );
  AOI211_X1 U9461 ( .C1(n9894), .C2(P1_ADDR_REG_15__SCAN_IN), .A(n7921), .B(
        n7920), .ZN(n7922) );
  INV_X1 U9462 ( .A(n7922), .ZN(P1_U3256) );
  INV_X1 U9463 ( .A(n7946), .ZN(n7926) );
  XOR2_X1 U9464 ( .A(n7927), .B(n7923), .Z(n7924) );
  AOI222_X1 U9465 ( .A1(n8722), .A2(n7924), .B1(n8343), .B2(n8686), .C1(n8345), 
        .C2(n8684), .ZN(n10187) );
  INV_X1 U9466 ( .A(n10187), .ZN(n7925) );
  AOI21_X1 U9467 ( .B1(n7926), .B2(n8743), .A(n7925), .ZN(n7937) );
  OR2_X1 U9468 ( .A1(n7928), .A2(n7927), .ZN(n7929) );
  AND2_X1 U9469 ( .A1(n7930), .A2(n7929), .ZN(n10190) );
  OAI21_X1 U9470 ( .B1(n7931), .B2(n10188), .A(n10126), .ZN(n7932) );
  OR2_X1 U9471 ( .A1(n7933), .A2(n7932), .ZN(n10186) );
  AOI22_X1 U9472 ( .A1(n10102), .A2(n7950), .B1(n10108), .B2(
        P2_REG2_REG_11__SCAN_IN), .ZN(n7934) );
  OAI21_X1 U9473 ( .B1(n10186), .B2(n10098), .A(n7934), .ZN(n7935) );
  AOI21_X1 U9474 ( .B1(n10190), .B2(n10105), .A(n7935), .ZN(n7936) );
  OAI21_X1 U9475 ( .B1(n7937), .B2(n10108), .A(n7936), .ZN(P2_U3285) );
  INV_X1 U9476 ( .A(n7938), .ZN(n7940) );
  OAI222_X1 U9477 ( .A1(P2_U3152), .A2(n7939), .B1(n8859), .B2(n7940), .C1(
        n9671), .C2(n8124), .ZN(P2_U3334) );
  OAI222_X1 U9478 ( .A1(n9449), .A2(n7942), .B1(P1_U3084), .B2(n7941), .C1(
        n9445), .C2(n7940), .ZN(P1_U3329) );
  XNOR2_X1 U9479 ( .A(n7944), .B(n7943), .ZN(n7952) );
  OAI22_X1 U9480 ( .A1(n8317), .A2(n7946), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7945), .ZN(n7949) );
  OAI22_X1 U9481 ( .A1(n7947), .A2(n8330), .B1(n8331), .B2(n8049), .ZN(n7948)
         );
  AOI211_X1 U9482 ( .C1(n7950), .C2(n8319), .A(n7949), .B(n7948), .ZN(n7951)
         );
  OAI21_X1 U9483 ( .B1(n7952), .B2(n8321), .A(n7951), .ZN(P2_U3238) );
  NAND2_X1 U9484 ( .A1(n7991), .A2(n9008), .ZN(n7953) );
  NAND2_X1 U9485 ( .A1(n7954), .A2(n7953), .ZN(n9820) );
  OR2_X1 U9486 ( .A1(n7979), .A2(n9007), .ZN(n7955) );
  NAND2_X1 U9487 ( .A1(n9820), .A2(n7955), .ZN(n7957) );
  NAND2_X1 U9488 ( .A1(n7979), .A2(n9007), .ZN(n7956) );
  XOR2_X1 U9489 ( .A(n7961), .B(n8095), .Z(n9419) );
  OAI211_X1 U9490 ( .C1(n7962), .C2(n7961), .A(n8065), .B(n9963), .ZN(n7964)
         );
  AOI22_X1 U9491 ( .A1(n9287), .A2(n9007), .B1(n9285), .B2(n9005), .ZN(n7963)
         );
  NAND2_X1 U9492 ( .A1(n7964), .A2(n7963), .ZN(n9414) );
  INV_X1 U9493 ( .A(n7979), .ZN(n9857) );
  INV_X1 U9494 ( .A(n9317), .ZN(n7965) );
  AOI211_X1 U9495 ( .C1(n9416), .C2(n9823), .A(n10034), .B(n7965), .ZN(n9415)
         );
  NAND2_X1 U9496 ( .A1(n9415), .A2(n9301), .ZN(n7967) );
  AOI22_X1 U9497 ( .A1(n9970), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n9969), .B2(
        n8874), .ZN(n7966) );
  OAI211_X1 U9498 ( .C1(n4616), .C2(n9972), .A(n7967), .B(n7966), .ZN(n7968)
         );
  AOI21_X1 U9499 ( .B1(n9836), .B2(n9414), .A(n7968), .ZN(n7969) );
  OAI21_X1 U9500 ( .B1(n9419), .B2(n9308), .A(n7969), .ZN(P1_U3277) );
  XNOR2_X1 U9501 ( .A(n7971), .B(n7970), .ZN(n7972) );
  XNOR2_X1 U9502 ( .A(n7973), .B(n7972), .ZN(n7981) );
  INV_X1 U9503 ( .A(n7974), .ZN(n7975) );
  AOI21_X1 U9504 ( .B1(n8991), .B2(n9006), .A(n7975), .ZN(n7977) );
  NAND2_X1 U9505 ( .A1(n8992), .A2(n9833), .ZN(n7976) );
  OAI211_X1 U9506 ( .C1(n9845), .C2(n8995), .A(n7977), .B(n7976), .ZN(n7978)
         );
  AOI21_X1 U9507 ( .B1(n7979), .B2(n8997), .A(n7978), .ZN(n7980) );
  OAI21_X1 U9508 ( .B1(n7981), .B2(n8999), .A(n7980), .ZN(P1_U3232) );
  INV_X1 U9509 ( .A(n7982), .ZN(n7983) );
  AOI21_X1 U9510 ( .B1(n7985), .B2(n7984), .A(n7983), .ZN(n7993) );
  AOI22_X1 U9511 ( .A1(n8991), .A2(n9007), .B1(P1_REG3_REG_12__SCAN_IN), .B2(
        P1_U3084), .ZN(n7988) );
  NAND2_X1 U9512 ( .A1(n8992), .A2(n7986), .ZN(n7987) );
  OAI211_X1 U9513 ( .C1(n7989), .C2(n8995), .A(n7988), .B(n7987), .ZN(n7990)
         );
  AOI21_X1 U9514 ( .B1(n7991), .B2(n8997), .A(n7990), .ZN(n7992) );
  OAI21_X1 U9515 ( .B1(n7993), .B2(n8999), .A(n7992), .ZN(P1_U3222) );
  OR2_X1 U9516 ( .A1(n8023), .A2(n8343), .ZN(n7994) );
  AND2_X2 U9517 ( .A1(n7995), .A2(n7994), .ZN(n7997) );
  OAI21_X1 U9518 ( .B1(n7997), .B2(n7996), .A(n8028), .ZN(n9807) );
  OAI21_X1 U9519 ( .B1(n4945), .B2(n7999), .A(n7998), .ZN(n8001) );
  OAI22_X1 U9520 ( .A1(n8738), .A2(n10070), .B1(n8049), .B2(n10072), .ZN(n8000) );
  AOI21_X1 U9521 ( .B1(n8001), .B2(n8722), .A(n8000), .ZN(n8002) );
  OAI21_X1 U9522 ( .B1(n8717), .B2(n9807), .A(n8002), .ZN(n9810) );
  NAND2_X1 U9523 ( .A1(n9810), .A2(n8749), .ZN(n8009) );
  OAI22_X1 U9524 ( .A1(n10081), .A2(n8003), .B1(n8048), .B2(n10096), .ZN(n8007) );
  INV_X1 U9525 ( .A(n8026), .ZN(n9808) );
  OR2_X1 U9526 ( .A1(n8004), .A2(n9808), .ZN(n8005) );
  NAND2_X1 U9527 ( .A1(n8033), .A2(n8005), .ZN(n9809) );
  NOR2_X1 U9528 ( .A1(n9809), .A2(n10085), .ZN(n8006) );
  AOI211_X1 U9529 ( .C1(n10102), .C2(n8026), .A(n8007), .B(n8006), .ZN(n8008)
         );
  OAI211_X1 U9530 ( .C1(n9807), .C2(n8730), .A(n8009), .B(n8008), .ZN(P2_U3283) );
  INV_X1 U9531 ( .A(n8010), .ZN(n8014) );
  OAI222_X1 U9532 ( .A1(n8124), .A2(n8012), .B1(n8859), .B2(n8014), .C1(
        P2_U3152), .C2(n8011), .ZN(P2_U3333) );
  OAI222_X1 U9533 ( .A1(n9449), .A2(n9542), .B1(n9452), .B2(n8014), .C1(n8013), 
        .C2(P1_U3084), .ZN(P1_U3328) );
  NAND2_X1 U9534 ( .A1(n8016), .A2(n8015), .ZN(n8018) );
  XOR2_X1 U9535 ( .A(n8018), .B(n8017), .Z(n8025) );
  NAND2_X1 U9536 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3152), .ZN(n8382) );
  OAI21_X1 U9537 ( .B1(n8317), .B2(n8019), .A(n8382), .ZN(n8022) );
  OAI22_X1 U9538 ( .A1(n8179), .A2(n8331), .B1(n8330), .B2(n8020), .ZN(n8021)
         );
  AOI211_X1 U9539 ( .C1(n8023), .C2(n8319), .A(n8022), .B(n8021), .ZN(n8024)
         );
  OAI21_X1 U9540 ( .B1(n8025), .B2(n8321), .A(n8024), .ZN(P2_U3226) );
  NAND2_X1 U9541 ( .A1(n8026), .A2(n8342), .ZN(n8027) );
  OAI21_X1 U9542 ( .B1(n4465), .B2(n4948), .A(n8476), .ZN(n9805) );
  INV_X1 U9543 ( .A(n9805), .ZN(n8039) );
  AOI211_X1 U9544 ( .C1(n4948), .C2(n8030), .A(n10089), .B(n4466), .ZN(n8032)
         );
  OAI22_X1 U9545 ( .A1(n8719), .A2(n10070), .B1(n8179), .B2(n10072), .ZN(n8031) );
  OR2_X1 U9546 ( .A1(n8032), .A2(n8031), .ZN(n9803) );
  INV_X1 U9547 ( .A(n8033), .ZN(n8034) );
  OAI21_X1 U9548 ( .B1(n8034), .B2(n4637), .A(n8739), .ZN(n9802) );
  OAI22_X1 U9549 ( .A1(n10081), .A2(n6124), .B1(n8178), .B2(n10096), .ZN(n8035) );
  AOI21_X1 U9550 ( .B1(n8475), .B2(n10102), .A(n8035), .ZN(n8036) );
  OAI21_X1 U9551 ( .B1(n9802), .B2(n10085), .A(n8036), .ZN(n8037) );
  AOI21_X1 U9552 ( .B1(n9803), .B2(n8749), .A(n8037), .ZN(n8038) );
  OAI21_X1 U9553 ( .B1(n8039), .B2(n8751), .A(n8038), .ZN(P2_U3282) );
  INV_X1 U9554 ( .A(n8040), .ZN(n8043) );
  OAI222_X1 U9555 ( .A1(P2_U3152), .A2(n8042), .B1(n8859), .B2(n8043), .C1(
        n8041), .C2(n8124), .ZN(P2_U3332) );
  OAI222_X1 U9556 ( .A1(n9449), .A2(n8045), .B1(P1_U3084), .B2(n8044), .C1(
        n9445), .C2(n8043), .ZN(P1_U3327) );
  OAI211_X1 U9557 ( .C1(n8047), .C2(n8046), .A(n8172), .B(n8325), .ZN(n8054)
         );
  INV_X1 U9558 ( .A(n8048), .ZN(n8052) );
  OAI22_X1 U9559 ( .A1(n8049), .A2(n8330), .B1(n8331), .B2(n8738), .ZN(n8050)
         );
  AOI211_X1 U9560 ( .C1(n8334), .C2(n8052), .A(n8051), .B(n8050), .ZN(n8053)
         );
  OAI211_X1 U9561 ( .C1(n9808), .C2(n8337), .A(n8054), .B(n8053), .ZN(P2_U3236) );
  INV_X1 U9562 ( .A(n8055), .ZN(n8058) );
  AOI21_X1 U9563 ( .B1(P2_DATAO_REG_27__SCAN_IN), .B2(n9730), .A(n8056), .ZN(
        n8057) );
  OAI21_X1 U9564 ( .B1(n8058), .B2(n9452), .A(n8057), .ZN(P1_U3326) );
  OAI222_X1 U9565 ( .A1(n8124), .A2(n9684), .B1(n8859), .B2(n8058), .C1(n8464), 
        .C2(P2_U3152), .ZN(P2_U3331) );
  OAI222_X1 U9566 ( .A1(n8124), .A2(n8061), .B1(n8859), .B2(n8060), .C1(n8059), 
        .C2(P2_U3152), .ZN(P2_U3338) );
  OAI222_X1 U9567 ( .A1(n9449), .A2(n8063), .B1(n9452), .B2(n8062), .C1(n6434), 
        .C2(P1_U3084), .ZN(P1_U3331) );
  NAND2_X1 U9568 ( .A1(n8065), .A2(n8064), .ZN(n9310) );
  INV_X1 U9569 ( .A(n9296), .ZN(n8068) );
  NAND2_X1 U9570 ( .A1(n9293), .A2(n8069), .ZN(n9283) );
  NAND2_X1 U9571 ( .A1(n9283), .A2(n8070), .ZN(n9261) );
  NAND2_X1 U9572 ( .A1(n9261), .A2(n9260), .ZN(n8071) );
  NOR2_X1 U9573 ( .A1(n9213), .A2(n8075), .ZN(n8076) );
  NAND2_X1 U9574 ( .A1(n9209), .A2(n8076), .ZN(n9210) );
  NAND2_X1 U9575 ( .A1(n9210), .A2(n8077), .ZN(n9200) );
  NAND2_X1 U9576 ( .A1(n9200), .A2(n8078), .ZN(n8080) );
  NAND2_X1 U9577 ( .A1(n9165), .A2(n9164), .ZN(n9163) );
  NAND2_X1 U9578 ( .A1(n9163), .A2(n8083), .ZN(n9155) );
  NAND2_X1 U9579 ( .A1(n9155), .A2(n9154), .ZN(n9153) );
  NAND2_X1 U9580 ( .A1(n9153), .A2(n8084), .ZN(n9139) );
  INV_X1 U9581 ( .A(P1_B_REG_SCAN_IN), .ZN(n8089) );
  NOR2_X1 U9582 ( .A1(n4394), .A2(n8089), .ZN(n8090) );
  NOR2_X1 U9583 ( .A1(n9960), .A2(n8090), .ZN(n9094) );
  NAND2_X1 U9584 ( .A1(n9094), .A2(n9001), .ZN(n8091) );
  AND2_X1 U9585 ( .A1(n9416), .A2(n9006), .ZN(n8094) );
  NOR2_X1 U9586 ( .A1(n9408), .A2(n9005), .ZN(n8096) );
  NAND2_X1 U9587 ( .A1(n9405), .A2(n9288), .ZN(n8097) );
  NAND2_X1 U9588 ( .A1(n8098), .A2(n8097), .ZN(n9276) );
  AND2_X1 U9589 ( .A1(n9398), .A2(n9004), .ZN(n8099) );
  OR2_X1 U9590 ( .A1(n9398), .A2(n9004), .ZN(n8100) );
  NAND2_X1 U9591 ( .A1(n8101), .A2(n8100), .ZN(n9255) );
  NOR2_X1 U9592 ( .A1(n9388), .A2(n9237), .ZN(n8103) );
  INV_X1 U9593 ( .A(n9388), .ZN(n8102) );
  INV_X1 U9594 ( .A(n9381), .ZN(n9232) );
  NAND2_X1 U9595 ( .A1(n8104), .A2(n4955), .ZN(n9207) );
  AOI22_X1 U9596 ( .A1(n9207), .A2(n9213), .B1(n9378), .B2(n9236), .ZN(n9194)
         );
  NAND2_X1 U9597 ( .A1(n9371), .A2(n9190), .ZN(n8105) );
  INV_X1 U9598 ( .A(n9371), .ZN(n9199) );
  AOI21_X1 U9599 ( .B1(n9194), .B2(n8105), .A(n4958), .ZN(n9178) );
  NAND2_X1 U9600 ( .A1(n9178), .A2(n8106), .ZN(n8108) );
  NOR2_X1 U9601 ( .A1(n9351), .A2(n9156), .ZN(n8111) );
  OAI22_X1 U9602 ( .A1(n9133), .A2(n8111), .B1(n9126), .B2(n4618), .ZN(n9117)
         );
  NAND2_X1 U9603 ( .A1(n9334), .A2(n9109), .ZN(n8121) );
  INV_X1 U9604 ( .A(n9398), .ZN(n9281) );
  NAND2_X1 U9605 ( .A1(n9300), .A2(n9281), .ZN(n9277) );
  INV_X1 U9606 ( .A(n9378), .ZN(n9223) );
  INV_X1 U9607 ( .A(n9356), .ZN(n9152) );
  INV_X1 U9608 ( .A(n9110), .ZN(n8114) );
  INV_X1 U9609 ( .A(n9336), .ZN(n8118) );
  AOI211_X1 U9610 ( .C1(n9336), .C2(n8114), .A(n10034), .B(n9098), .ZN(n9335)
         );
  INV_X1 U9611 ( .A(n8115), .ZN(n8116) );
  AOI22_X1 U9612 ( .A1(n8116), .A2(n9969), .B1(P1_REG2_REG_29__SCAN_IN), .B2(
        n9321), .ZN(n8117) );
  OAI21_X1 U9613 ( .B1(n8118), .B2(n9972), .A(n8117), .ZN(n8119) );
  AOI21_X1 U9614 ( .B1(n9335), .B2(n9301), .A(n8119), .ZN(n8120) );
  OAI211_X1 U9615 ( .C1(n9338), .C2(n9321), .A(n8121), .B(n8120), .ZN(P1_U3355) );
  OAI222_X1 U9616 ( .A1(n8124), .A2(n8123), .B1(n8859), .B2(n8122), .C1(
        P2_U3152), .C2(n8668), .ZN(P2_U3339) );
  AND2_X1 U9617 ( .A1(n8599), .A2(n6726), .ZN(n8157) );
  XNOR2_X1 U9618 ( .A(n8783), .B(n6724), .ZN(n8156) );
  NAND2_X1 U9619 ( .A1(n8290), .A2(n8125), .ZN(n8130) );
  XNOR2_X1 U9620 ( .A(n8815), .B(n6724), .ZN(n8126) );
  AND2_X1 U9621 ( .A1(n8212), .A2(n8481), .ZN(n8127) );
  NAND2_X1 U9622 ( .A1(n8126), .A2(n8127), .ZN(n8131) );
  INV_X1 U9623 ( .A(n8126), .ZN(n8195) );
  INV_X1 U9624 ( .A(n8127), .ZN(n8128) );
  NAND2_X1 U9625 ( .A1(n8195), .A2(n8128), .ZN(n8129) );
  AND2_X1 U9626 ( .A1(n8131), .A2(n8129), .ZN(n8288) );
  NAND2_X1 U9627 ( .A1(n8130), .A2(n8288), .ZN(n8194) );
  XNOR2_X1 U9628 ( .A(n8811), .B(n6724), .ZN(n8133) );
  NAND2_X1 U9629 ( .A1(n8212), .A2(n8687), .ZN(n8134) );
  XNOR2_X1 U9630 ( .A(n8133), .B(n8134), .ZN(n8205) );
  AND2_X1 U9631 ( .A1(n8205), .A2(n8131), .ZN(n8132) );
  INV_X1 U9632 ( .A(n8133), .ZN(n8135) );
  NAND2_X1 U9633 ( .A1(n8135), .A2(n8134), .ZN(n8136) );
  XNOR2_X1 U9634 ( .A(n8805), .B(n6724), .ZN(n8137) );
  INV_X1 U9635 ( .A(n8229), .ZN(n8486) );
  AND2_X1 U9636 ( .A1(n6726), .A2(n8486), .ZN(n8138) );
  NAND2_X1 U9637 ( .A1(n8137), .A2(n8138), .ZN(n8142) );
  INV_X1 U9638 ( .A(n8137), .ZN(n8225) );
  INV_X1 U9639 ( .A(n8138), .ZN(n8139) );
  NAND2_X1 U9640 ( .A1(n8225), .A2(n8139), .ZN(n8140) );
  NAND2_X1 U9641 ( .A1(n8142), .A2(n8140), .ZN(n8272) );
  INV_X1 U9642 ( .A(n8272), .ZN(n8141) );
  XNOR2_X1 U9643 ( .A(n8800), .B(n6724), .ZN(n8145) );
  NAND2_X1 U9644 ( .A1(n8212), .A2(n8652), .ZN(n8143) );
  XNOR2_X1 U9645 ( .A(n8145), .B(n8143), .ZN(n8223) );
  INV_X1 U9646 ( .A(n8143), .ZN(n8144) );
  NAND2_X1 U9647 ( .A1(n8145), .A2(n8144), .ZN(n8146) );
  NAND2_X1 U9648 ( .A1(n8226), .A2(n8146), .ZN(n8149) );
  XNOR2_X1 U9649 ( .A(n8795), .B(n6739), .ZN(n8147) );
  XNOR2_X1 U9650 ( .A(n8149), .B(n8147), .ZN(n8281) );
  INV_X1 U9651 ( .A(n8230), .ZN(n8600) );
  NAND2_X1 U9652 ( .A1(n6726), .A2(n8600), .ZN(n8280) );
  INV_X1 U9653 ( .A(n8147), .ZN(n8148) );
  NOR2_X1 U9654 ( .A1(n8149), .A2(n8148), .ZN(n8150) );
  AOI21_X1 U9655 ( .B1(n8281), .B2(n8280), .A(n8150), .ZN(n8153) );
  XNOR2_X1 U9656 ( .A(n8607), .B(n6724), .ZN(n8152) );
  INV_X1 U9657 ( .A(n8152), .ZN(n8151) );
  AND2_X1 U9658 ( .A1(n8153), .A2(n8151), .ZN(n8259) );
  OAI21_X1 U9659 ( .B1(n8157), .B2(n8156), .A(n8259), .ZN(n8158) );
  XNOR2_X1 U9660 ( .A(n8153), .B(n8152), .ZN(n8187) );
  AND2_X1 U9661 ( .A1(n6726), .A2(n8490), .ZN(n8188) );
  INV_X1 U9662 ( .A(n8156), .ZN(n8261) );
  INV_X1 U9663 ( .A(n8157), .ZN(n8265) );
  XNOR2_X1 U9664 ( .A(n8779), .B(n6724), .ZN(n8159) );
  NOR2_X1 U9665 ( .A1(n8592), .A2(n8165), .ZN(n8160) );
  AND2_X1 U9666 ( .A1(n8159), .A2(n8160), .ZN(n8238) );
  INV_X1 U9667 ( .A(n8159), .ZN(n8239) );
  INV_X1 U9668 ( .A(n8160), .ZN(n8161) );
  NAND2_X1 U9669 ( .A1(n8239), .A2(n8161), .ZN(n8237) );
  INV_X1 U9670 ( .A(n8543), .ZN(n8492) );
  NAND2_X1 U9671 ( .A1(n8492), .A2(n8212), .ZN(n8163) );
  XNOR2_X1 U9672 ( .A(n8774), .B(n6724), .ZN(n8162) );
  XOR2_X1 U9673 ( .A(n8163), .B(n8162), .Z(n8311) );
  INV_X1 U9674 ( .A(n8162), .ZN(n8164) );
  INV_X1 U9675 ( .A(n8768), .ZN(n8536) );
  XNOR2_X1 U9676 ( .A(n8536), .B(n6724), .ZN(n8207) );
  NOR2_X1 U9677 ( .A1(n8339), .A2(n8165), .ZN(n8209) );
  XNOR2_X1 U9678 ( .A(n8207), .B(n8209), .ZN(n8210) );
  XNOR2_X1 U9679 ( .A(n8211), .B(n8210), .ZN(n8171) );
  INV_X1 U9680 ( .A(n8534), .ZN(n8167) );
  OAI22_X1 U9681 ( .A1(n8167), .A2(n8317), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8166), .ZN(n8169) );
  OAI22_X1 U9682 ( .A1(n8544), .A2(n8331), .B1(n8330), .B2(n8543), .ZN(n8168)
         );
  AOI211_X1 U9683 ( .C1(n8768), .C2(n8319), .A(n8169), .B(n8168), .ZN(n8170)
         );
  OAI21_X1 U9684 ( .B1(n8171), .B2(n8321), .A(n8170), .ZN(P2_U3216) );
  INV_X1 U9685 ( .A(n8172), .ZN(n8175) );
  NOR3_X1 U9686 ( .A1(n8173), .A2(n8179), .A3(n8291), .ZN(n8174) );
  AOI21_X1 U9687 ( .B1(n8175), .B2(n8325), .A(n8174), .ZN(n8186) );
  NOR2_X1 U9688 ( .A1(n8176), .A2(n8321), .ZN(n8183) );
  AND2_X1 U9689 ( .A1(n8475), .A2(n8319), .ZN(n8182) );
  OAI21_X1 U9690 ( .B1(n8317), .B2(n8178), .A(n8177), .ZN(n8181) );
  OAI22_X1 U9691 ( .A1(n8719), .A2(n8331), .B1(n8330), .B2(n8179), .ZN(n8180)
         );
  NOR4_X1 U9692 ( .A1(n8183), .A2(n8182), .A3(n8181), .A4(n8180), .ZN(n8184)
         );
  OAI21_X1 U9693 ( .B1(n8186), .B2(n8185), .A(n8184), .ZN(P2_U3217) );
  AOI22_X1 U9694 ( .A1(n8187), .A2(n8325), .B1(n8323), .B2(n8490), .ZN(n8193)
         );
  AND2_X1 U9695 ( .A1(n8187), .A2(n8188), .ZN(n8260) );
  OAI22_X1 U9696 ( .A1(n8317), .A2(n8604), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8189), .ZN(n8191) );
  OAI22_X1 U9697 ( .A1(n8263), .A2(n8331), .B1(n8330), .B2(n8230), .ZN(n8190)
         );
  AOI211_X1 U9698 ( .C1(n8789), .C2(n8319), .A(n8191), .B(n8190), .ZN(n8192)
         );
  OAI21_X1 U9699 ( .B1(n8193), .B2(n8260), .A(n8192), .ZN(P2_U3218) );
  INV_X1 U9700 ( .A(n8194), .ZN(n8197) );
  NOR3_X1 U9701 ( .A1(n8195), .A2(n8698), .A3(n8291), .ZN(n8196) );
  AOI21_X1 U9702 ( .B1(n8197), .B2(n8325), .A(n8196), .ZN(n8206) );
  OR2_X1 U9703 ( .A1(n8229), .A2(n10070), .ZN(n8199) );
  NAND2_X1 U9704 ( .A1(n8481), .A2(n8684), .ZN(n8198) );
  NAND2_X1 U9705 ( .A1(n8199), .A2(n8198), .ZN(n8665) );
  AOI22_X1 U9706 ( .A1(n8315), .A2(n8665), .B1(P2_REG3_REG_19__SCAN_IN), .B2(
        P2_U3152), .ZN(n8200) );
  OAI21_X1 U9707 ( .B1(n8671), .B2(n8317), .A(n8200), .ZN(n8203) );
  NOR2_X1 U9708 ( .A1(n8201), .A2(n8321), .ZN(n8202) );
  AOI211_X1 U9709 ( .C1(n8811), .C2(n8319), .A(n8203), .B(n8202), .ZN(n8204)
         );
  OAI21_X1 U9710 ( .B1(n8206), .B2(n8205), .A(n8204), .ZN(P2_U3221) );
  INV_X1 U9711 ( .A(n8207), .ZN(n8208) );
  NAND2_X1 U9712 ( .A1(n8505), .A2(n8212), .ZN(n8213) );
  XOR2_X1 U9713 ( .A(n6724), .B(n8213), .Z(n8214) );
  XNOR2_X1 U9714 ( .A(n8763), .B(n8214), .ZN(n8215) );
  INV_X1 U9715 ( .A(n8216), .ZN(n8526) );
  OR2_X1 U9716 ( .A1(n8339), .A2(n10072), .ZN(n8218) );
  NAND2_X1 U9717 ( .A1(n8338), .A2(n8686), .ZN(n8217) );
  NAND2_X1 U9718 ( .A1(n8218), .A2(n8217), .ZN(n8523) );
  AOI22_X1 U9719 ( .A1(n8523), .A2(n8315), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3152), .ZN(n8219) );
  OAI21_X1 U9720 ( .B1(n8526), .B2(n8317), .A(n8219), .ZN(n8220) );
  AOI21_X1 U9721 ( .B1(n8763), .B2(n8319), .A(n8220), .ZN(n8221) );
  OAI21_X1 U9722 ( .B1(n8222), .B2(n8321), .A(n8221), .ZN(P2_U3222) );
  INV_X1 U9723 ( .A(n8223), .ZN(n8224) );
  AOI21_X1 U9724 ( .B1(n8274), .B2(n8224), .A(n8321), .ZN(n8228) );
  NOR3_X1 U9725 ( .A1(n8225), .A2(n8229), .A3(n8291), .ZN(n8227) );
  OAI21_X1 U9726 ( .B1(n8228), .B2(n8227), .A(n8226), .ZN(n8236) );
  INV_X1 U9727 ( .A(n8315), .ZN(n8233) );
  OAI22_X1 U9728 ( .A1(n8230), .A2(n10070), .B1(n8229), .B2(n10072), .ZN(n8637) );
  INV_X1 U9729 ( .A(n8637), .ZN(n8232) );
  OAI22_X1 U9730 ( .A1(n8233), .A2(n8232), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8231), .ZN(n8234) );
  AOI21_X1 U9731 ( .B1(n8632), .B2(n8334), .A(n8234), .ZN(n8235) );
  OAI211_X1 U9732 ( .C1(n8634), .C2(n8337), .A(n8236), .B(n8235), .ZN(P2_U3225) );
  OR3_X1 U9733 ( .A1(n8238), .A2(n4810), .A3(n8321), .ZN(n8243) );
  NOR3_X1 U9734 ( .A1(n8239), .A2(n8592), .A3(n8291), .ZN(n8240) );
  AOI21_X1 U9735 ( .B1(n8325), .B2(n4810), .A(n8240), .ZN(n8242) );
  MUX2_X1 U9736 ( .A(n8243), .B(n8242), .S(n8241), .Z(n8247) );
  OAI22_X1 U9737 ( .A1(n8543), .A2(n10070), .B1(n8263), .B2(n10072), .ZN(n8571) );
  AOI22_X1 U9738 ( .A1(n8571), .A2(n8315), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3152), .ZN(n8246) );
  NAND2_X1 U9739 ( .A1(n8779), .A2(n8319), .ZN(n8245) );
  NAND2_X1 U9740 ( .A1(n8334), .A2(n8577), .ZN(n8244) );
  NAND4_X1 U9741 ( .A1(n8247), .A2(n8246), .A3(n8245), .A4(n8244), .ZN(
        P2_U3227) );
  XNOR2_X1 U9742 ( .A(n8249), .B(n8248), .ZN(n8326) );
  AOI22_X1 U9743 ( .A1(n8326), .A2(n8324), .B1(n8250), .B2(n8249), .ZN(n8254)
         );
  XNOR2_X1 U9744 ( .A(n8252), .B(n8251), .ZN(n8253) );
  XNOR2_X1 U9745 ( .A(n8254), .B(n8253), .ZN(n8258) );
  NAND2_X1 U9746 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(P2_U3152), .ZN(n8401) );
  OAI21_X1 U9747 ( .B1(n8317), .B2(n8724), .A(n8401), .ZN(n8256) );
  OAI22_X1 U9748 ( .A1(n8719), .A2(n8330), .B1(n8331), .B2(n8718), .ZN(n8255)
         );
  AOI211_X1 U9749 ( .C1(n8825), .C2(n8319), .A(n8256), .B(n8255), .ZN(n8257)
         );
  OAI21_X1 U9750 ( .B1(n8258), .B2(n8321), .A(n8257), .ZN(P2_U3228) );
  NOR2_X1 U9751 ( .A1(n8260), .A2(n8259), .ZN(n8262) );
  XNOR2_X1 U9752 ( .A(n8262), .B(n8261), .ZN(n8266) );
  OAI22_X1 U9753 ( .A1(n8266), .A2(n8321), .B1(n8263), .B2(n8291), .ZN(n8264)
         );
  OAI21_X1 U9754 ( .B1(n8266), .B2(n8265), .A(n8264), .ZN(n8271) );
  OAI22_X1 U9755 ( .A1(n8317), .A2(n8587), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8267), .ZN(n8269) );
  OAI22_X1 U9756 ( .A1(n8624), .A2(n8330), .B1(n8331), .B2(n8592), .ZN(n8268)
         );
  AOI211_X1 U9757 ( .C1(n8783), .C2(n8319), .A(n8269), .B(n8268), .ZN(n8270)
         );
  NAND2_X1 U9758 ( .A1(n8271), .A2(n8270), .ZN(P2_U3231) );
  INV_X1 U9759 ( .A(n8805), .ZN(n8648) );
  AOI21_X1 U9760 ( .B1(n8273), .B2(n8272), .A(n8321), .ZN(n8275) );
  NAND2_X1 U9761 ( .A1(n8275), .A2(n8274), .ZN(n8279) );
  NOR2_X1 U9762 ( .A1(n8317), .A2(n8645), .ZN(n8277) );
  OAI22_X1 U9763 ( .A1(n8623), .A2(n8331), .B1(n8330), .B2(n8484), .ZN(n8276)
         );
  AOI211_X1 U9764 ( .C1(P2_REG3_REG_20__SCAN_IN), .C2(P2_U3152), .A(n8277), 
        .B(n8276), .ZN(n8278) );
  OAI211_X1 U9765 ( .C1(n8648), .C2(n8337), .A(n8279), .B(n8278), .ZN(P2_U3235) );
  INV_X1 U9766 ( .A(n8795), .ZN(n8620) );
  NAND2_X1 U9767 ( .A1(n8323), .A2(n8600), .ZN(n8283) );
  NAND2_X1 U9768 ( .A1(n8325), .A2(n8280), .ZN(n8282) );
  MUX2_X1 U9769 ( .A(n8283), .B(n8282), .S(n8281), .Z(n8287) );
  NOR2_X1 U9770 ( .A1(n8317), .A2(n8617), .ZN(n8285) );
  OAI22_X1 U9771 ( .A1(n8624), .A2(n8331), .B1(n8330), .B2(n8623), .ZN(n8284)
         );
  AOI211_X1 U9772 ( .C1(P2_REG3_REG_22__SCAN_IN), .C2(P2_U3152), .A(n8285), 
        .B(n8284), .ZN(n8286) );
  OAI211_X1 U9773 ( .C1(n8620), .C2(n8337), .A(n8287), .B(n8286), .ZN(P2_U3237) );
  INV_X1 U9774 ( .A(n8815), .ZN(n8681) );
  INV_X1 U9775 ( .A(n8288), .ZN(n8289) );
  AOI21_X1 U9776 ( .B1(n8290), .B2(n8289), .A(n8321), .ZN(n8294) );
  NOR3_X1 U9777 ( .A1(n8292), .A2(n8718), .A3(n8291), .ZN(n8293) );
  OAI21_X1 U9778 ( .B1(n8294), .B2(n8293), .A(n8194), .ZN(n8298) );
  INV_X1 U9779 ( .A(n8295), .ZN(n8679) );
  AND2_X1 U9780 ( .A1(P2_U3152), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8437) );
  OAI22_X1 U9781 ( .A1(n8718), .A2(n8330), .B1(n8331), .B2(n8484), .ZN(n8296)
         );
  AOI211_X1 U9782 ( .C1(n8334), .C2(n8679), .A(n8437), .B(n8296), .ZN(n8297)
         );
  OAI211_X1 U9783 ( .C1(n8681), .C2(n8337), .A(n8298), .B(n8297), .ZN(P2_U3240) );
  OAI21_X1 U9784 ( .B1(n8301), .B2(n8300), .A(n8299), .ZN(n8302) );
  NAND2_X1 U9785 ( .A1(n8302), .A2(n8325), .ZN(n8310) );
  AOI22_X1 U9786 ( .A1(n8304), .A2(n8348), .B1(n8303), .B2(n8319), .ZN(n8309)
         );
  NAND2_X1 U9787 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3152), .ZN(n8369) );
  OAI21_X1 U9788 ( .B1(n8317), .B2(n8305), .A(n8369), .ZN(n8306) );
  AOI21_X1 U9789 ( .B1(n8307), .B2(n8350), .A(n8306), .ZN(n8308) );
  NAND3_X1 U9790 ( .A1(n8310), .A2(n8309), .A3(n8308), .ZN(P2_U3241) );
  XNOR2_X1 U9791 ( .A(n8312), .B(n8311), .ZN(n8322) );
  OR2_X1 U9792 ( .A1(n8339), .A2(n10070), .ZN(n8314) );
  INV_X1 U9793 ( .A(n8592), .ZN(n8341) );
  NAND2_X1 U9794 ( .A1(n8341), .A2(n8684), .ZN(n8313) );
  NAND2_X1 U9795 ( .A1(n8314), .A2(n8313), .ZN(n8560) );
  AOI22_X1 U9796 ( .A1(n8560), .A2(n8315), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3152), .ZN(n8316) );
  OAI21_X1 U9797 ( .B1(n8552), .B2(n8317), .A(n8316), .ZN(n8318) );
  AOI21_X1 U9798 ( .B1(n8774), .B2(n8319), .A(n8318), .ZN(n8320) );
  OAI21_X1 U9799 ( .B1(n8322), .B2(n8321), .A(n8320), .ZN(P2_U3242) );
  INV_X1 U9800 ( .A(n8745), .ZN(n9796) );
  NAND2_X1 U9801 ( .A1(n8323), .A2(n8477), .ZN(n8328) );
  NAND2_X1 U9802 ( .A1(n8325), .A2(n8324), .ZN(n8327) );
  MUX2_X1 U9803 ( .A(n8328), .B(n8327), .S(n8326), .Z(n8336) );
  INV_X1 U9804 ( .A(n8329), .ZN(n8744) );
  OAI22_X1 U9805 ( .A1(n8737), .A2(n8331), .B1(n8330), .B2(n8738), .ZN(n8332)
         );
  AOI211_X1 U9806 ( .C1(n8744), .C2(n8334), .A(n8333), .B(n8332), .ZN(n8335)
         );
  OAI211_X1 U9807 ( .C1(n9796), .C2(n8337), .A(n8336), .B(n8335), .ZN(P2_U3243) );
  MUX2_X1 U9808 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n8503), .S(P2_U3966), .Z(
        P2_U3582) );
  MUX2_X1 U9809 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n8338), .S(P2_U3966), .Z(
        P2_U3581) );
  MUX2_X1 U9810 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n8505), .S(P2_U3966), .Z(
        P2_U3580) );
  INV_X1 U9811 ( .A(n8339), .ZN(n8495) );
  MUX2_X1 U9812 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8495), .S(P2_U3966), .Z(
        P2_U3579) );
  MUX2_X1 U9813 ( .A(n8492), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8340), .Z(
        P2_U3578) );
  MUX2_X1 U9814 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n8341), .S(P2_U3966), .Z(
        P2_U3577) );
  MUX2_X1 U9815 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n8599), .S(P2_U3966), .Z(
        P2_U3576) );
  MUX2_X1 U9816 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(n8490), .S(P2_U3966), .Z(
        P2_U3575) );
  MUX2_X1 U9817 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8600), .S(P2_U3966), .Z(
        P2_U3574) );
  MUX2_X1 U9818 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n8652), .S(P2_U3966), .Z(
        P2_U3573) );
  MUX2_X1 U9819 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8486), .S(P2_U3966), .Z(
        P2_U3572) );
  MUX2_X1 U9820 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n8687), .S(P2_U3966), .Z(
        P2_U3571) );
  MUX2_X1 U9821 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n8481), .S(P2_U3966), .Z(
        P2_U3570) );
  MUX2_X1 U9822 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8685), .S(P2_U3966), .Z(
        P2_U3569) );
  MUX2_X1 U9823 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n8479), .S(P2_U3966), .Z(
        P2_U3568) );
  MUX2_X1 U9824 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n8477), .S(P2_U3966), .Z(
        P2_U3567) );
  MUX2_X1 U9825 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n8474), .S(P2_U3966), .Z(
        P2_U3566) );
  MUX2_X1 U9826 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n8342), .S(P2_U3966), .Z(
        P2_U3565) );
  MUX2_X1 U9827 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n8343), .S(P2_U3966), .Z(
        P2_U3564) );
  MUX2_X1 U9828 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n8344), .S(P2_U3966), .Z(
        P2_U3563) );
  MUX2_X1 U9829 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n8345), .S(P2_U3966), .Z(
        P2_U3562) );
  MUX2_X1 U9830 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n8346), .S(P2_U3966), .Z(
        P2_U3561) );
  MUX2_X1 U9831 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n8347), .S(P2_U3966), .Z(
        P2_U3560) );
  MUX2_X1 U9832 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n8348), .S(P2_U3966), .Z(
        P2_U3559) );
  MUX2_X1 U9833 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n8349), .S(P2_U3966), .Z(
        P2_U3558) );
  MUX2_X1 U9834 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(n8350), .S(P2_U3966), .Z(
        P2_U3557) );
  MUX2_X1 U9835 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n8351), .S(P2_U3966), .Z(
        P2_U3556) );
  MUX2_X1 U9836 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(n8352), .S(P2_U3966), .Z(
        P2_U3555) );
  MUX2_X1 U9837 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(n6725), .S(P2_U3966), .Z(
        P2_U3554) );
  MUX2_X1 U9838 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n6718), .S(P2_U3966), .Z(
        P2_U3553) );
  MUX2_X1 U9839 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(n5990), .S(P2_U3966), .Z(
        P2_U3552) );
  NAND2_X1 U9840 ( .A1(n8354), .A2(n8353), .ZN(n8355) );
  NAND3_X1 U9841 ( .A1(n10057), .A2(n8356), .A3(n8355), .ZN(n8365) );
  INV_X1 U9842 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n9683) );
  NOR2_X1 U9843 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9683), .ZN(n8357) );
  AOI21_X1 U9844 ( .B1(n10058), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n8357), .ZN(
        n8364) );
  NAND2_X1 U9845 ( .A1(n9753), .A2(n8358), .ZN(n8363) );
  OAI211_X1 U9846 ( .C1(n8361), .C2(n8360), .A(n10056), .B(n8359), .ZN(n8362)
         );
  NAND4_X1 U9847 ( .A1(n8365), .A2(n8364), .A3(n8363), .A4(n8362), .ZN(
        P2_U3250) );
  OAI211_X1 U9848 ( .C1(n8368), .C2(n8367), .A(n10057), .B(n8366), .ZN(n8378)
         );
  INV_X1 U9849 ( .A(n8369), .ZN(n8370) );
  AOI21_X1 U9850 ( .B1(n10058), .B2(P2_ADDR_REG_6__SCAN_IN), .A(n8370), .ZN(
        n8377) );
  NAND2_X1 U9851 ( .A1(n9753), .A2(n8371), .ZN(n8376) );
  OAI211_X1 U9852 ( .C1(n8374), .C2(n8373), .A(n10056), .B(n8372), .ZN(n8375)
         );
  NAND4_X1 U9853 ( .A1(n8378), .A2(n8377), .A3(n8376), .A4(n8375), .ZN(
        P2_U3251) );
  OAI211_X1 U9854 ( .C1(n8381), .C2(n8380), .A(n10057), .B(n8379), .ZN(n8392)
         );
  INV_X1 U9855 ( .A(n8382), .ZN(n8383) );
  AOI21_X1 U9856 ( .B1(n10058), .B2(P2_ADDR_REG_12__SCAN_IN), .A(n8383), .ZN(
        n8391) );
  NAND2_X1 U9857 ( .A1(n9753), .A2(n8384), .ZN(n8390) );
  OAI21_X1 U9858 ( .B1(n8387), .B2(n8386), .A(n8385), .ZN(n8388) );
  NAND2_X1 U9859 ( .A1(n10056), .A2(n8388), .ZN(n8389) );
  NAND4_X1 U9860 ( .A1(n8392), .A2(n8391), .A3(n8390), .A4(n8389), .ZN(
        P2_U3257) );
  NOR2_X1 U9861 ( .A1(n8394), .A2(n8393), .ZN(n8396) );
  XNOR2_X1 U9862 ( .A(n8420), .B(n8397), .ZN(n8398) );
  NAND2_X1 U9863 ( .A1(n8398), .A2(n8399), .ZN(n8421) );
  OAI21_X1 U9864 ( .B1(n8399), .B2(n8398), .A(n8421), .ZN(n8400) );
  NAND2_X1 U9865 ( .A1(n8400), .A2(n10056), .ZN(n8413) );
  INV_X1 U9866 ( .A(n8401), .ZN(n8402) );
  AOI21_X1 U9867 ( .B1(n10058), .B2(P2_ADDR_REG_16__SCAN_IN), .A(n8402), .ZN(
        n8412) );
  NOR2_X1 U9868 ( .A1(n8404), .A2(n8403), .ZN(n8406) );
  MUX2_X1 U9869 ( .A(n8725), .B(P2_REG2_REG_16__SCAN_IN), .S(n8420), .Z(n8407)
         );
  INV_X1 U9870 ( .A(n8407), .ZN(n8408) );
  NAND2_X1 U9871 ( .A1(n8408), .A2(n8409), .ZN(n8414) );
  OAI211_X1 U9872 ( .C1(n8409), .C2(n8408), .A(n10057), .B(n8414), .ZN(n8411)
         );
  NAND2_X1 U9873 ( .A1(n9753), .A2(n8420), .ZN(n8410) );
  NAND4_X1 U9874 ( .A1(n8413), .A2(n8412), .A3(n8411), .A4(n8410), .ZN(
        P2_U3261) );
  NAND2_X1 U9875 ( .A1(n8420), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n8415) );
  NAND2_X1 U9876 ( .A1(n8415), .A2(n8414), .ZN(n8418) );
  MUX2_X1 U9877 ( .A(n8706), .B(P2_REG2_REG_17__SCAN_IN), .S(n8432), .Z(n8416)
         );
  INV_X1 U9878 ( .A(n8416), .ZN(n8417) );
  NAND2_X1 U9879 ( .A1(n8417), .A2(n8418), .ZN(n8433) );
  OAI211_X1 U9880 ( .C1(n8418), .C2(n8417), .A(n10057), .B(n8433), .ZN(n8429)
         );
  NOR2_X1 U9881 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6163), .ZN(n8419) );
  AOI21_X1 U9882 ( .B1(n10058), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n8419), .ZN(
        n8428) );
  NAND2_X1 U9883 ( .A1(n9753), .A2(n8432), .ZN(n8427) );
  XNOR2_X1 U9884 ( .A(n8432), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n8424) );
  OR2_X1 U9885 ( .A1(n8420), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n8422) );
  AOI21_X1 U9886 ( .B1(n8424), .B2(n8423), .A(n8430), .ZN(n8425) );
  NAND2_X1 U9887 ( .A1(n10056), .A2(n8425), .ZN(n8426) );
  NAND4_X1 U9888 ( .A1(n8429), .A2(n8428), .A3(n8427), .A4(n8426), .ZN(
        P2_U3262) );
  XNOR2_X1 U9889 ( .A(n8447), .B(n8431), .ZN(n8446) );
  XOR2_X1 U9890 ( .A(n8445), .B(n8446), .Z(n8440) );
  NAND2_X1 U9891 ( .A1(n8432), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n8434) );
  NAND2_X1 U9892 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n8435), .ZN(n8444) );
  OAI211_X1 U9893 ( .C1(n8435), .C2(P2_REG2_REG_18__SCAN_IN), .A(n10057), .B(
        n8444), .ZN(n8439) );
  INV_X1 U9894 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n10256) );
  NOR2_X1 U9895 ( .A1(n8460), .A2(n10256), .ZN(n8436) );
  AOI211_X1 U9896 ( .C1(n9753), .C2(n8447), .A(n8437), .B(n8436), .ZN(n8438)
         );
  OAI211_X1 U9897 ( .C1(n8440), .C2(n10060), .A(n8439), .B(n8438), .ZN(
        P2_U3263) );
  NAND2_X1 U9898 ( .A1(n8442), .A2(n8447), .ZN(n8443) );
  OR2_X1 U9899 ( .A1(n8447), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n8448) );
  NAND2_X1 U9900 ( .A1(n8449), .A2(n8448), .ZN(n8451) );
  XNOR2_X1 U9901 ( .A(n8451), .B(n8450), .ZN(n8455) );
  INV_X1 U9902 ( .A(n8455), .ZN(n8452) );
  AOI22_X1 U9903 ( .A1(n8453), .A2(n10057), .B1(n8452), .B2(n10056), .ZN(n8457) );
  NOR2_X1 U9904 ( .A1(n8453), .A2(n10061), .ZN(n8454) );
  AOI211_X1 U9905 ( .C1(n10056), .C2(n8455), .A(n9753), .B(n8454), .ZN(n8456)
         );
  MUX2_X1 U9906 ( .A(n8457), .B(n8456), .S(n6322), .Z(n8459) );
  NAND2_X1 U9907 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(P2_U3152), .ZN(n8458) );
  OAI211_X1 U9908 ( .C1(n8441), .C2(n8460), .A(n8459), .B(n8458), .ZN(P2_U3264) );
  INV_X1 U9909 ( .A(n8825), .ZN(n8461) );
  NAND3_X1 U9910 ( .A1(n8644), .A2(n8634), .A3(n8620), .ZN(n8614) );
  NAND2_X1 U9911 ( .A1(n8573), .A2(n8580), .ZN(n8574) );
  XOR2_X1 U9912 ( .A(n8753), .B(n8469), .Z(n8755) );
  NOR2_X1 U9913 ( .A1(n8749), .A2(n8462), .ZN(n8467) );
  INV_X1 U9914 ( .A(P2_B_REG_SCAN_IN), .ZN(n8463) );
  NOR2_X1 U9915 ( .A1(n8464), .A2(n8463), .ZN(n8465) );
  NOR2_X1 U9916 ( .A1(n10070), .A2(n8465), .ZN(n8504) );
  NAND2_X1 U9917 ( .A1(n8466), .A2(n8504), .ZN(n9791) );
  NOR2_X1 U9918 ( .A1(n10104), .A2(n9791), .ZN(n8471) );
  AOI211_X1 U9919 ( .C1(n8753), .C2(n10102), .A(n8467), .B(n8471), .ZN(n8468)
         );
  OAI21_X1 U9920 ( .B1(n8755), .B2(n10085), .A(n8468), .ZN(P2_U3265) );
  AOI21_X1 U9921 ( .B1(n8470), .B2(n8508), .A(n8469), .ZN(n9794) );
  NAND2_X1 U9922 ( .A1(n9794), .A2(n8727), .ZN(n8473) );
  AOI21_X1 U9923 ( .B1(n10108), .B2(P2_REG2_REG_30__SCAN_IN), .A(n8471), .ZN(
        n8472) );
  OAI211_X1 U9924 ( .C1(n9792), .C2(n8703), .A(n8473), .B(n8472), .ZN(P2_U3266) );
  NOR2_X1 U9925 ( .A1(n8745), .A2(n8477), .ZN(n8478) );
  AND2_X2 U9926 ( .A1(n8714), .A2(n8713), .ZN(n8716) );
  NOR2_X2 U9927 ( .A1(n8716), .A2(n8480), .ZN(n8693) );
  NAND2_X1 U9928 ( .A1(n8815), .A2(n8481), .ZN(n8482) );
  INV_X1 U9929 ( .A(n8811), .ZN(n8485) );
  NAND2_X1 U9930 ( .A1(n8800), .A2(n8652), .ZN(n8488) );
  AOI21_X2 U9931 ( .B1(n8631), .B2(n8488), .A(n8487), .ZN(n8613) );
  OAI22_X2 U9932 ( .A1(n8550), .A2(n8493), .B1(n8774), .B2(n8492), .ZN(n8530)
         );
  NAND2_X1 U9933 ( .A1(n8530), .A2(n8494), .ZN(n8497) );
  NOR2_X1 U9934 ( .A1(n8763), .A2(n8505), .ZN(n8498) );
  XNOR2_X1 U9935 ( .A(n8500), .B(n8499), .ZN(n8756) );
  INV_X1 U9936 ( .A(n8756), .ZN(n8515) );
  XOR2_X1 U9937 ( .A(n8502), .B(n8501), .Z(n8507) );
  AOI22_X1 U9938 ( .A1(n8505), .A2(n8684), .B1(n8504), .B2(n8503), .ZN(n8506)
         );
  OAI21_X1 U9939 ( .B1(n4414), .B2(n8757), .A(n8508), .ZN(n8758) );
  OAI22_X1 U9940 ( .A1(n10081), .A2(n8510), .B1(n8509), .B2(n10096), .ZN(n8511) );
  AOI21_X1 U9941 ( .B1(n4635), .B2(n10102), .A(n8511), .ZN(n8512) );
  OAI21_X1 U9942 ( .B1(n8758), .B2(n10085), .A(n8512), .ZN(n8513) );
  AOI21_X1 U9943 ( .B1(n8760), .B2(n8749), .A(n8513), .ZN(n8514) );
  OAI21_X1 U9944 ( .B1(n8515), .B2(n8751), .A(n8514), .ZN(P2_U3267) );
  XNOR2_X1 U9945 ( .A(n8517), .B(n8516), .ZN(n8767) );
  AOI21_X1 U9946 ( .B1(n8763), .B2(n8531), .A(n4414), .ZN(n8764) );
  INV_X1 U9947 ( .A(n8763), .ZN(n8519) );
  OAI22_X1 U9948 ( .A1(n8519), .A2(n8703), .B1(n10081), .B2(n8518), .ZN(n8520)
         );
  AOI21_X1 U9949 ( .B1(n8764), .B2(n8727), .A(n8520), .ZN(n8529) );
  AOI21_X1 U9950 ( .B1(n4509), .B2(n8522), .A(n10089), .ZN(n8525) );
  AOI21_X1 U9951 ( .B1(n8525), .B2(n8524), .A(n8523), .ZN(n8766) );
  OAI21_X1 U9952 ( .B1(n8526), .B2(n10096), .A(n8766), .ZN(n8527) );
  NAND2_X1 U9953 ( .A1(n8527), .A2(n8749), .ZN(n8528) );
  OAI211_X1 U9954 ( .C1(n8767), .C2(n8751), .A(n8529), .B(n8528), .ZN(P2_U3268) );
  XNOR2_X1 U9955 ( .A(n8530), .B(n8539), .ZN(n8772) );
  INV_X1 U9956 ( .A(n8551), .ZN(n8533) );
  INV_X1 U9957 ( .A(n8531), .ZN(n8532) );
  AOI21_X1 U9958 ( .B1(n8768), .B2(n8533), .A(n8532), .ZN(n8769) );
  AOI22_X1 U9959 ( .A1(n10108), .A2(P2_REG2_REG_27__SCAN_IN), .B1(n8534), .B2(
        n8743), .ZN(n8535) );
  OAI21_X1 U9960 ( .B1(n8536), .B2(n8703), .A(n8535), .ZN(n8548) );
  INV_X1 U9961 ( .A(n8537), .ZN(n8542) );
  AOI21_X1 U9962 ( .B1(n8538), .B2(n8540), .A(n8539), .ZN(n8541) );
  NOR3_X1 U9963 ( .A1(n8542), .A2(n8541), .A3(n10089), .ZN(n8546) );
  OAI22_X1 U9964 ( .A1(n8544), .A2(n10070), .B1(n8543), .B2(n10072), .ZN(n8545) );
  NOR2_X1 U9965 ( .A1(n8546), .A2(n8545), .ZN(n8771) );
  NOR2_X1 U9966 ( .A1(n8771), .A2(n10108), .ZN(n8547) );
  AOI211_X1 U9967 ( .C1(n8727), .C2(n8769), .A(n8548), .B(n8547), .ZN(n8549)
         );
  OAI21_X1 U9968 ( .B1(n8772), .B2(n8751), .A(n8549), .ZN(P2_U3269) );
  XNOR2_X1 U9969 ( .A(n8550), .B(n8557), .ZN(n8777) );
  AOI211_X1 U9970 ( .C1(n8774), .C2(n8574), .A(n10194), .B(n8551), .ZN(n8773)
         );
  INV_X1 U9971 ( .A(n8774), .ZN(n8555) );
  INV_X1 U9972 ( .A(n8552), .ZN(n8553) );
  AOI22_X1 U9973 ( .A1(n10104), .A2(P2_REG2_REG_26__SCAN_IN), .B1(n8553), .B2(
        n8743), .ZN(n8554) );
  OAI21_X1 U9974 ( .B1(n8555), .B2(n8703), .A(n8554), .ZN(n8563) );
  INV_X1 U9975 ( .A(n8556), .ZN(n8568) );
  OAI21_X1 U9976 ( .B1(n8568), .B2(n8558), .A(n8557), .ZN(n8559) );
  AOI21_X1 U9977 ( .B1(n8559), .B2(n8538), .A(n10089), .ZN(n8561) );
  NOR2_X1 U9978 ( .A1(n8561), .A2(n8560), .ZN(n8776) );
  NOR2_X1 U9979 ( .A1(n8776), .A2(n10104), .ZN(n8562) );
  AOI211_X1 U9980 ( .C1(n8773), .C2(n8709), .A(n8563), .B(n8562), .ZN(n8564)
         );
  OAI21_X1 U9981 ( .B1(n8777), .B2(n8751), .A(n8564), .ZN(P2_U3270) );
  XNOR2_X1 U9982 ( .A(n8566), .B(n8565), .ZN(n8782) );
  INV_X1 U9983 ( .A(n8567), .ZN(n8570) );
  AOI211_X1 U9984 ( .C1(n8570), .C2(n8569), .A(n10089), .B(n8568), .ZN(n8572)
         );
  NOR2_X1 U9985 ( .A1(n8572), .A2(n8571), .ZN(n8781) );
  INV_X1 U9986 ( .A(n8573), .ZN(n8576) );
  INV_X1 U9987 ( .A(n8574), .ZN(n8575) );
  AOI211_X1 U9988 ( .C1(n8779), .C2(n8576), .A(n10194), .B(n8575), .ZN(n8778)
         );
  AOI22_X1 U9989 ( .A1(n8778), .A2(n8668), .B1(n8743), .B2(n8577), .ZN(n8578)
         );
  AOI21_X1 U9990 ( .B1(n8781), .B2(n8578), .A(n10104), .ZN(n8582) );
  OAI22_X1 U9991 ( .A1(n8580), .A2(n8703), .B1(n10081), .B2(n8579), .ZN(n8581)
         );
  NOR2_X1 U9992 ( .A1(n8582), .A2(n8581), .ZN(n8583) );
  OAI21_X1 U9993 ( .B1(n8782), .B2(n8751), .A(n8583), .ZN(P2_U3271) );
  OAI21_X1 U9994 ( .B1(n8585), .B2(n8591), .A(n8584), .ZN(n8586) );
  INV_X1 U9995 ( .A(n8586), .ZN(n8787) );
  XOR2_X1 U9996 ( .A(n8783), .B(n8602), .Z(n8784) );
  INV_X1 U9997 ( .A(n8783), .ZN(n8590) );
  INV_X1 U9998 ( .A(n8587), .ZN(n8588) );
  AOI22_X1 U9999 ( .A1(n10104), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n8588), .B2(
        n8743), .ZN(n8589) );
  OAI21_X1 U10000 ( .B1(n8590), .B2(n8703), .A(n8589), .ZN(n8597) );
  AOI21_X1 U10001 ( .B1(n4435), .B2(n8591), .A(n10089), .ZN(n8595) );
  OAI22_X1 U10002 ( .A1(n8592), .A2(n10070), .B1(n8624), .B2(n10072), .ZN(
        n8593) );
  AOI21_X1 U10003 ( .B1(n8595), .B2(n8594), .A(n8593), .ZN(n8786) );
  NOR2_X1 U10004 ( .A1(n8786), .A2(n10108), .ZN(n8596) );
  AOI211_X1 U10005 ( .C1(n8784), .C2(n8727), .A(n8597), .B(n8596), .ZN(n8598)
         );
  OAI21_X1 U10006 ( .B1(n8787), .B2(n8751), .A(n8598), .ZN(P2_U3272) );
  OAI21_X1 U10007 ( .B1(n4430), .B2(n8609), .A(n4737), .ZN(n8601) );
  AOI222_X1 U10008 ( .A1(n8722), .A2(n8601), .B1(n8600), .B2(n8684), .C1(n8599), .C2(n8686), .ZN(n8792) );
  INV_X1 U10009 ( .A(n8602), .ZN(n8603) );
  AOI21_X1 U10010 ( .B1(n8789), .B2(n8614), .A(n8603), .ZN(n8790) );
  INV_X1 U10011 ( .A(n8604), .ZN(n8605) );
  AOI22_X1 U10012 ( .A1(n10104), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n8605), 
        .B2(n8743), .ZN(n8606) );
  OAI21_X1 U10013 ( .B1(n8607), .B2(n8703), .A(n8606), .ZN(n8608) );
  AOI21_X1 U10014 ( .B1(n8790), .B2(n8727), .A(n8608), .ZN(n8612) );
  NAND2_X1 U10015 ( .A1(n8610), .A2(n8609), .ZN(n8788) );
  NAND3_X1 U10016 ( .A1(n4941), .A2(n10105), .A3(n8788), .ZN(n8611) );
  OAI211_X1 U10017 ( .C1(n8792), .C2(n10104), .A(n8612), .B(n8611), .ZN(
        P2_U3273) );
  XNOR2_X1 U10018 ( .A(n8613), .B(n8621), .ZN(n8799) );
  INV_X1 U10019 ( .A(n8614), .ZN(n8616) );
  AOI21_X1 U10020 ( .B1(n8644), .B2(n8634), .A(n8620), .ZN(n8615) );
  NOR2_X1 U10021 ( .A1(n8616), .A2(n8615), .ZN(n8796) );
  INV_X1 U10022 ( .A(n8617), .ZN(n8618) );
  AOI22_X1 U10023 ( .A1(n10104), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n8618), 
        .B2(n8743), .ZN(n8619) );
  OAI21_X1 U10024 ( .B1(n8620), .B2(n8703), .A(n8619), .ZN(n8629) );
  AOI21_X1 U10025 ( .B1(n8622), .B2(n8621), .A(n10089), .ZN(n8627) );
  OAI22_X1 U10026 ( .A1(n8624), .A2(n10070), .B1(n8623), .B2(n10072), .ZN(
        n8625) );
  AOI21_X1 U10027 ( .B1(n8627), .B2(n8626), .A(n8625), .ZN(n8798) );
  NOR2_X1 U10028 ( .A1(n8798), .A2(n10108), .ZN(n8628) );
  AOI211_X1 U10029 ( .C1(n8796), .C2(n8727), .A(n8629), .B(n8628), .ZN(n8630)
         );
  OAI21_X1 U10030 ( .B1(n8799), .B2(n8751), .A(n8630), .ZN(P2_U3274) );
  XOR2_X1 U10031 ( .A(n8635), .B(n8631), .Z(n8804) );
  XNOR2_X1 U10032 ( .A(n8644), .B(n8800), .ZN(n8801) );
  AOI22_X1 U10033 ( .A1(n10104), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n8632), 
        .B2(n8743), .ZN(n8633) );
  OAI21_X1 U10034 ( .B1(n8634), .B2(n8703), .A(n8633), .ZN(n8640) );
  XNOR2_X1 U10035 ( .A(n8636), .B(n8635), .ZN(n8638) );
  AOI21_X1 U10036 ( .B1(n8638), .B2(n8722), .A(n8637), .ZN(n8803) );
  NOR2_X1 U10037 ( .A1(n8803), .A2(n10108), .ZN(n8639) );
  AOI211_X1 U10038 ( .C1(n8801), .C2(n8727), .A(n8640), .B(n8639), .ZN(n8641)
         );
  OAI21_X1 U10039 ( .B1(n8804), .B2(n8751), .A(n8641), .ZN(P2_U3275) );
  XNOR2_X1 U10040 ( .A(n8643), .B(n8642), .ZN(n8809) );
  AOI21_X1 U10041 ( .B1(n8805), .B2(n4643), .A(n8644), .ZN(n8806) );
  INV_X1 U10042 ( .A(n8645), .ZN(n8646) );
  AOI22_X1 U10043 ( .A1(n10108), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n8646), 
        .B2(n8743), .ZN(n8647) );
  OAI21_X1 U10044 ( .B1(n8648), .B2(n8703), .A(n8647), .ZN(n8656) );
  OAI211_X1 U10045 ( .C1(n8649), .C2(n8651), .A(n8650), .B(n8722), .ZN(n8654)
         );
  AOI22_X1 U10046 ( .A1(n8686), .A2(n8652), .B1(n8687), .B2(n8684), .ZN(n8653)
         );
  AND2_X1 U10047 ( .A1(n8654), .A2(n8653), .ZN(n8808) );
  NOR2_X1 U10048 ( .A1(n8808), .A2(n10108), .ZN(n8655) );
  AOI211_X1 U10049 ( .C1(n8806), .C2(n8727), .A(n8656), .B(n8655), .ZN(n8657)
         );
  OAI21_X1 U10050 ( .B1(n8751), .B2(n8809), .A(n8657), .ZN(P2_U3276) );
  XNOR2_X1 U10051 ( .A(n8659), .B(n8658), .ZN(n8814) );
  AND2_X1 U10052 ( .A1(n8661), .A2(n8660), .ZN(n8664) );
  OAI21_X1 U10053 ( .B1(n8664), .B2(n8663), .A(n8662), .ZN(n8666) );
  AOI21_X1 U10054 ( .B1(n8666), .B2(n8722), .A(n8665), .ZN(n8813) );
  AOI211_X1 U10055 ( .C1(n8811), .C2(n8677), .A(n10194), .B(n8667), .ZN(n8810)
         );
  NAND2_X1 U10056 ( .A1(n8810), .A2(n8668), .ZN(n8669) );
  OAI211_X1 U10057 ( .C1(n8814), .C2(n8717), .A(n8813), .B(n8669), .ZN(n8670)
         );
  NAND2_X1 U10058 ( .A1(n8670), .A2(n8749), .ZN(n8675) );
  OAI22_X1 U10059 ( .A1(n8749), .A2(n8672), .B1(n8671), .B2(n10096), .ZN(n8673) );
  AOI21_X1 U10060 ( .B1(n8811), .B2(n10102), .A(n8673), .ZN(n8674) );
  OAI211_X1 U10061 ( .C1(n8814), .C2(n8730), .A(n8675), .B(n8674), .ZN(
        P2_U3277) );
  XOR2_X1 U10062 ( .A(n8676), .B(n8682), .Z(n8819) );
  INV_X1 U10063 ( .A(n8677), .ZN(n8678) );
  AOI21_X1 U10064 ( .B1(n8815), .B2(n8700), .A(n8678), .ZN(n8816) );
  AOI22_X1 U10065 ( .A1(n10108), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n8679), 
        .B2(n8743), .ZN(n8680) );
  OAI21_X1 U10066 ( .B1(n8681), .B2(n8703), .A(n8680), .ZN(n8690) );
  XNOR2_X1 U10067 ( .A(n8683), .B(n8682), .ZN(n8688) );
  AOI222_X1 U10068 ( .A1(n8722), .A2(n8688), .B1(n8687), .B2(n8686), .C1(n8685), .C2(n8684), .ZN(n8818) );
  NOR2_X1 U10069 ( .A1(n8818), .A2(n10108), .ZN(n8689) );
  AOI211_X1 U10070 ( .C1(n8816), .C2(n8727), .A(n8690), .B(n8689), .ZN(n8691)
         );
  OAI21_X1 U10071 ( .B1(n8819), .B2(n8751), .A(n8691), .ZN(P2_U3278) );
  OAI21_X1 U10072 ( .B1(n8693), .B2(n8695), .A(n8692), .ZN(n8694) );
  INV_X1 U10073 ( .A(n8694), .ZN(n8824) );
  XNOR2_X1 U10074 ( .A(n8696), .B(n8695), .ZN(n8697) );
  OAI222_X1 U10075 ( .A1(n10072), .A2(n8737), .B1(n10070), .B2(n8698), .C1(
        n10089), .C2(n8697), .ZN(n8820) );
  NAND2_X1 U10076 ( .A1(n8820), .A2(n8749), .ZN(n8711) );
  INV_X1 U10077 ( .A(n8699), .ZN(n8702) );
  INV_X1 U10078 ( .A(n8700), .ZN(n8701) );
  AOI211_X1 U10079 ( .C1(n8822), .C2(n8702), .A(n10194), .B(n8701), .ZN(n8821)
         );
  NOR2_X1 U10080 ( .A1(n8704), .A2(n8703), .ZN(n8708) );
  OAI22_X1 U10081 ( .A1(n8749), .A2(n8706), .B1(n8705), .B2(n10096), .ZN(n8707) );
  AOI211_X1 U10082 ( .C1(n8821), .C2(n8709), .A(n8708), .B(n8707), .ZN(n8710)
         );
  OAI211_X1 U10083 ( .C1(n8824), .C2(n8751), .A(n8711), .B(n8710), .ZN(
        P2_U3279) );
  XNOR2_X1 U10084 ( .A(n8712), .B(n8713), .ZN(n8723) );
  NOR2_X1 U10085 ( .A1(n8714), .A2(n8713), .ZN(n8715) );
  NOR2_X1 U10086 ( .A1(n8829), .A2(n8717), .ZN(n8721) );
  OAI22_X1 U10087 ( .A1(n8719), .A2(n10072), .B1(n8718), .B2(n10070), .ZN(
        n8720) );
  AOI211_X1 U10088 ( .C1(n8723), .C2(n8722), .A(n8721), .B(n8720), .ZN(n8828)
         );
  OAI22_X1 U10089 ( .A1(n10081), .A2(n8725), .B1(n8724), .B2(n10096), .ZN(
        n8726) );
  AOI21_X1 U10090 ( .B1(n8825), .B2(n10102), .A(n8726), .ZN(n8729) );
  XNOR2_X1 U10091 ( .A(n8740), .B(n8825), .ZN(n8826) );
  NAND2_X1 U10092 ( .A1(n8826), .A2(n8727), .ZN(n8728) );
  OAI211_X1 U10093 ( .C1(n8829), .C2(n8730), .A(n8729), .B(n8728), .ZN(n8731)
         );
  INV_X1 U10094 ( .A(n8731), .ZN(n8732) );
  OAI21_X1 U10095 ( .B1(n8828), .B2(n10108), .A(n8732), .ZN(P2_U3280) );
  XNOR2_X1 U10096 ( .A(n8733), .B(n8734), .ZN(n9800) );
  INV_X1 U10097 ( .A(n9800), .ZN(n8752) );
  XNOR2_X1 U10098 ( .A(n8735), .B(n8734), .ZN(n8736) );
  OAI222_X1 U10099 ( .A1(n10072), .A2(n8738), .B1(n10070), .B2(n8737), .C1(
        n10089), .C2(n8736), .ZN(n9798) );
  INV_X1 U10100 ( .A(n8739), .ZN(n8742) );
  INV_X1 U10101 ( .A(n8740), .ZN(n8741) );
  OAI21_X1 U10102 ( .B1(n9796), .B2(n8742), .A(n8741), .ZN(n9797) );
  AOI22_X1 U10103 ( .A1(n10108), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n8744), 
        .B2(n8743), .ZN(n8747) );
  NAND2_X1 U10104 ( .A1(n8745), .A2(n10102), .ZN(n8746) );
  OAI211_X1 U10105 ( .C1(n9797), .C2(n10085), .A(n8747), .B(n8746), .ZN(n8748)
         );
  AOI21_X1 U10106 ( .B1(n9798), .B2(n8749), .A(n8748), .ZN(n8750) );
  OAI21_X1 U10107 ( .B1(n8752), .B2(n8751), .A(n8750), .ZN(P2_U3281) );
  NAND2_X1 U10108 ( .A1(n8753), .A2(n10128), .ZN(n8754) );
  OAI211_X1 U10109 ( .C1(n8755), .C2(n10194), .A(n9791), .B(n8754), .ZN(n8830)
         );
  MUX2_X1 U10110 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n8830), .S(n10219), .Z(
        P2_U3551) );
  NAND2_X1 U10111 ( .A1(n8756), .A2(n10199), .ZN(n8762) );
  OAI22_X1 U10112 ( .A1(n8758), .A2(n10194), .B1(n8757), .B2(n10192), .ZN(
        n8759) );
  NOR2_X1 U10113 ( .A1(n8760), .A2(n8759), .ZN(n8761) );
  NAND2_X1 U10114 ( .A1(n8762), .A2(n8761), .ZN(n8831) );
  MUX2_X1 U10115 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n8831), .S(n10219), .Z(
        P2_U3549) );
  AOI22_X1 U10116 ( .A1(n8764), .A2(n10126), .B1(n10128), .B2(n8763), .ZN(
        n8765) );
  OAI211_X1 U10117 ( .C1(n8767), .C2(n10130), .A(n8766), .B(n8765), .ZN(n8832)
         );
  MUX2_X1 U10118 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n8832), .S(n10219), .Z(
        P2_U3548) );
  AOI22_X1 U10119 ( .A1(n8769), .A2(n10126), .B1(n10128), .B2(n8768), .ZN(
        n8770) );
  OAI211_X1 U10120 ( .C1(n8772), .C2(n10130), .A(n8771), .B(n8770), .ZN(n8833)
         );
  MUX2_X1 U10121 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n8833), .S(n10219), .Z(
        P2_U3547) );
  AOI21_X1 U10122 ( .B1(n10128), .B2(n8774), .A(n8773), .ZN(n8775) );
  OAI211_X1 U10123 ( .C1(n8777), .C2(n10130), .A(n8776), .B(n8775), .ZN(n8834)
         );
  MUX2_X1 U10124 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n8834), .S(n10219), .Z(
        P2_U3546) );
  AOI21_X1 U10125 ( .B1(n10128), .B2(n8779), .A(n8778), .ZN(n8780) );
  OAI211_X1 U10126 ( .C1(n10130), .C2(n8782), .A(n8781), .B(n8780), .ZN(n8835)
         );
  MUX2_X1 U10127 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n8835), .S(n10219), .Z(
        P2_U3545) );
  AOI22_X1 U10128 ( .A1(n8784), .A2(n10126), .B1(n10128), .B2(n8783), .ZN(
        n8785) );
  OAI211_X1 U10129 ( .C1(n8787), .C2(n10130), .A(n8786), .B(n8785), .ZN(n8836)
         );
  MUX2_X1 U10130 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n8836), .S(n10219), .Z(
        P2_U3544) );
  NAND2_X1 U10131 ( .A1(n8788), .A2(n10199), .ZN(n8793) );
  AOI22_X1 U10132 ( .A1(n8790), .A2(n10126), .B1(n10128), .B2(n8789), .ZN(
        n8791) );
  OAI211_X1 U10133 ( .C1(n8794), .C2(n8793), .A(n8792), .B(n8791), .ZN(n8837)
         );
  MUX2_X1 U10134 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n8837), .S(n10219), .Z(
        P2_U3543) );
  AOI22_X1 U10135 ( .A1(n8796), .A2(n10126), .B1(n10128), .B2(n8795), .ZN(
        n8797) );
  OAI211_X1 U10136 ( .C1(n10130), .C2(n8799), .A(n8798), .B(n8797), .ZN(n8838)
         );
  MUX2_X1 U10137 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n8838), .S(n10219), .Z(
        P2_U3542) );
  AOI22_X1 U10138 ( .A1(n8801), .A2(n10126), .B1(n10128), .B2(n8800), .ZN(
        n8802) );
  OAI211_X1 U10139 ( .C1(n8804), .C2(n10130), .A(n8803), .B(n8802), .ZN(n8839)
         );
  MUX2_X1 U10140 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n8839), .S(n10219), .Z(
        P2_U3541) );
  AOI22_X1 U10141 ( .A1(n8806), .A2(n10126), .B1(n10128), .B2(n8805), .ZN(
        n8807) );
  OAI211_X1 U10142 ( .C1(n10130), .C2(n8809), .A(n8808), .B(n8807), .ZN(n8840)
         );
  MUX2_X1 U10143 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n8840), .S(n10219), .Z(
        P2_U3540) );
  AOI21_X1 U10144 ( .B1(n10128), .B2(n8811), .A(n8810), .ZN(n8812) );
  OAI211_X1 U10145 ( .C1(n10130), .C2(n8814), .A(n8813), .B(n8812), .ZN(n8841)
         );
  MUX2_X1 U10146 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n8841), .S(n10219), .Z(
        P2_U3539) );
  AOI22_X1 U10147 ( .A1(n8816), .A2(n10126), .B1(n10128), .B2(n8815), .ZN(
        n8817) );
  OAI211_X1 U10148 ( .C1(n10130), .C2(n8819), .A(n8818), .B(n8817), .ZN(n8842)
         );
  MUX2_X1 U10149 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n8842), .S(n10219), .Z(
        P2_U3538) );
  AOI211_X1 U10150 ( .C1(n10128), .C2(n8822), .A(n8821), .B(n8820), .ZN(n8823)
         );
  OAI21_X1 U10151 ( .B1(n10130), .B2(n8824), .A(n8823), .ZN(n8843) );
  MUX2_X1 U10152 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n8843), .S(n10219), .Z(
        P2_U3537) );
  AOI22_X1 U10153 ( .A1(n8826), .A2(n10126), .B1(n10128), .B2(n8825), .ZN(
        n8827) );
  OAI211_X1 U10154 ( .C1(n9806), .C2(n8829), .A(n8828), .B(n8827), .ZN(n8844)
         );
  MUX2_X1 U10155 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n8844), .S(n10219), .Z(
        P2_U3536) );
  MUX2_X1 U10156 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n8830), .S(n10202), .Z(
        P2_U3519) );
  MUX2_X1 U10157 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n8831), .S(n10202), .Z(
        P2_U3517) );
  MUX2_X1 U10158 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n8832), .S(n10202), .Z(
        P2_U3516) );
  MUX2_X1 U10159 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n8833), .S(n10202), .Z(
        P2_U3515) );
  MUX2_X1 U10160 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n8834), .S(n10202), .Z(
        P2_U3514) );
  MUX2_X1 U10161 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n8835), .S(n10202), .Z(
        P2_U3513) );
  MUX2_X1 U10162 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n8836), .S(n10202), .Z(
        P2_U3512) );
  MUX2_X1 U10163 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n8837), .S(n10202), .Z(
        P2_U3511) );
  MUX2_X1 U10164 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n8838), .S(n10202), .Z(
        P2_U3510) );
  MUX2_X1 U10165 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n8839), .S(n10202), .Z(
        P2_U3509) );
  MUX2_X1 U10166 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n8840), .S(n10202), .Z(
        P2_U3508) );
  MUX2_X1 U10167 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n8841), .S(n10202), .Z(
        P2_U3507) );
  MUX2_X1 U10168 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n8842), .S(n10202), .Z(
        P2_U3505) );
  MUX2_X1 U10169 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n8843), .S(n10202), .Z(
        P2_U3502) );
  MUX2_X1 U10170 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n8844), .S(n10202), .Z(
        P2_U3499) );
  NOR4_X1 U10171 ( .A1(n8846), .A2(P2_IR_REG_30__SCAN_IN), .A3(n6416), .A4(
        P2_U3152), .ZN(n8847) );
  AOI21_X1 U10172 ( .B1(n8856), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n8847), .ZN(
        n8848) );
  OAI21_X1 U10173 ( .B1(n5133), .B2(n8859), .A(n8848), .ZN(P2_U3327) );
  INV_X1 U10174 ( .A(n8849), .ZN(n9444) );
  AOI22_X1 U10175 ( .A1(n8850), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n8856), .ZN(n8851) );
  OAI21_X1 U10176 ( .B1(n9444), .B2(n8859), .A(n8851), .ZN(P2_U3328) );
  INV_X1 U10177 ( .A(n8852), .ZN(n9446) );
  AOI22_X1 U10178 ( .A1(n8853), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_29__SCAN_IN), .B2(n8856), .ZN(n8854) );
  OAI21_X1 U10179 ( .B1(n9446), .B2(n8859), .A(n8854), .ZN(P2_U3329) );
  INV_X1 U10180 ( .A(n8855), .ZN(n9453) );
  AOI22_X1 U10181 ( .A1(n8857), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_28__SCAN_IN), .B2(n8856), .ZN(n8858) );
  OAI21_X1 U10182 ( .B1(n9453), .B2(n8859), .A(n8858), .ZN(P2_U3330) );
  MUX2_X1 U10183 ( .A(n8860), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3358) );
  XNOR2_X1 U10184 ( .A(n8862), .B(n8861), .ZN(n8863) );
  AOI22_X1 U10185 ( .A1(n9156), .A2(n8979), .B1(P1_REG3_REG_27__SCAN_IN), .B2(
        P1_U3084), .ZN(n8866) );
  NAND2_X1 U10186 ( .A1(n9120), .A2(n8992), .ZN(n8865) );
  OAI211_X1 U10187 ( .C1(n9127), .C2(n8972), .A(n8866), .B(n8865), .ZN(n8867)
         );
  AOI21_X1 U10188 ( .B1(n9346), .B2(n8997), .A(n8867), .ZN(n8868) );
  OAI21_X1 U10189 ( .B1(n8869), .B2(n8999), .A(n8868), .ZN(P1_U3212) );
  XNOR2_X1 U10190 ( .A(n8872), .B(n8871), .ZN(n8873) );
  XNOR2_X1 U10191 ( .A(n8870), .B(n8873), .ZN(n8880) );
  NAND2_X1 U10192 ( .A1(n8992), .A2(n8874), .ZN(n8877) );
  AOI21_X1 U10193 ( .B1(n8979), .B2(n9007), .A(n8875), .ZN(n8876) );
  OAI211_X1 U10194 ( .C1(n9298), .C2(n8972), .A(n8877), .B(n8876), .ZN(n8878)
         );
  AOI21_X1 U10195 ( .B1(n9416), .B2(n8997), .A(n8878), .ZN(n8879) );
  OAI21_X1 U10196 ( .B1(n8880), .B2(n8999), .A(n8879), .ZN(P1_U3213) );
  NAND2_X1 U10197 ( .A1(n4746), .A2(n8882), .ZN(n8884) );
  XNOR2_X1 U10198 ( .A(n8884), .B(n8883), .ZN(n8889) );
  AOI22_X1 U10199 ( .A1(n9183), .A2(n8991), .B1(P1_REG3_REG_23__SCAN_IN), .B2(
        P1_U3084), .ZN(n8886) );
  NAND2_X1 U10200 ( .A1(n8979), .A2(n9190), .ZN(n8885) );
  OAI211_X1 U10201 ( .C1(n8981), .C2(n9180), .A(n8886), .B(n8885), .ZN(n8887)
         );
  AOI21_X1 U10202 ( .B1(n9366), .B2(n8997), .A(n8887), .ZN(n8888) );
  OAI21_X1 U10203 ( .B1(n8889), .B2(n8999), .A(n8888), .ZN(P1_U3214) );
  XOR2_X1 U10204 ( .A(n8891), .B(n8890), .Z(n8892) );
  XNOR2_X1 U10205 ( .A(n8893), .B(n8892), .ZN(n8898) );
  NAND2_X1 U10206 ( .A1(P1_U3084), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9089) );
  OAI21_X1 U10207 ( .B1(n8995), .B2(n9244), .A(n9089), .ZN(n8894) );
  AOI21_X1 U10208 ( .B1(n8991), .B2(n9003), .A(n8894), .ZN(n8895) );
  OAI21_X1 U10209 ( .B1(n8981), .B2(n9248), .A(n8895), .ZN(n8896) );
  AOI21_X1 U10210 ( .B1(n9388), .B2(n8997), .A(n8896), .ZN(n8897) );
  OAI21_X1 U10211 ( .B1(n8898), .B2(n8999), .A(n8897), .ZN(P1_U3217) );
  OAI21_X1 U10212 ( .B1(n8901), .B2(n8900), .A(n8899), .ZN(n8902) );
  NAND2_X1 U10213 ( .A1(n8902), .A2(n8976), .ZN(n8907) );
  OAI22_X1 U10214 ( .A1(n9215), .A2(n8972), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8903), .ZN(n8905) );
  NOR2_X1 U10215 ( .A1(n8981), .A2(n9219), .ZN(n8904) );
  AOI211_X1 U10216 ( .C1(n8979), .C2(n9003), .A(n8905), .B(n8904), .ZN(n8906)
         );
  OAI211_X1 U10217 ( .C1(n9223), .C2(n8985), .A(n8907), .B(n8906), .ZN(
        P1_U3221) );
  XOR2_X1 U10218 ( .A(n8908), .B(n8909), .Z(n8914) );
  AOI22_X1 U10219 ( .A1(n9183), .A2(n8979), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3084), .ZN(n8911) );
  NAND2_X1 U10220 ( .A1(n9150), .A2(n8992), .ZN(n8910) );
  OAI211_X1 U10221 ( .C1(n9126), .C2(n8972), .A(n8911), .B(n8910), .ZN(n8912)
         );
  AOI21_X1 U10222 ( .B1(n9356), .B2(n8997), .A(n8912), .ZN(n8913) );
  OAI21_X1 U10223 ( .B1(n8914), .B2(n8999), .A(n8913), .ZN(P1_U3223) );
  INV_X1 U10224 ( .A(n9405), .ZN(n9305) );
  OAI21_X1 U10225 ( .B1(n8917), .B2(n4764), .A(n8916), .ZN(n8918) );
  OAI21_X1 U10226 ( .B1(n8919), .B2(n4764), .A(n8918), .ZN(n8920) );
  NAND2_X1 U10227 ( .A1(n8920), .A2(n8976), .ZN(n8925) );
  NOR2_X1 U10228 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n8921), .ZN(n9041) );
  AOI21_X1 U10229 ( .B1(n8991), .B2(n9004), .A(n9041), .ZN(n8922) );
  OAI21_X1 U10230 ( .B1(n9298), .B2(n8995), .A(n8922), .ZN(n8923) );
  AOI21_X1 U10231 ( .B1(n9302), .B2(n8992), .A(n8923), .ZN(n8924) );
  OAI211_X1 U10232 ( .C1(n9305), .C2(n8985), .A(n8925), .B(n8924), .ZN(
        P1_U3224) );
  OAI21_X1 U10233 ( .B1(n8928), .B2(n8926), .A(n8927), .ZN(n8929) );
  NAND2_X1 U10234 ( .A1(n8929), .A2(n8976), .ZN(n8934) );
  OAI22_X1 U10235 ( .A1(n8972), .A2(n9244), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8930), .ZN(n8932) );
  NOR2_X1 U10236 ( .A1(n8995), .A2(n9311), .ZN(n8931) );
  AOI211_X1 U10237 ( .C1(n9279), .C2(n8992), .A(n8932), .B(n8931), .ZN(n8933)
         );
  OAI211_X1 U10238 ( .C1(n9281), .C2(n8985), .A(n8934), .B(n8933), .ZN(
        P1_U3226) );
  XOR2_X1 U10239 ( .A(n8936), .B(n8935), .Z(n8941) );
  AOI22_X1 U10240 ( .A1(n9166), .A2(n8991), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3084), .ZN(n8938) );
  NAND2_X1 U10241 ( .A1(n9203), .A2(n8979), .ZN(n8937) );
  OAI211_X1 U10242 ( .C1(n8981), .C2(n9171), .A(n8938), .B(n8937), .ZN(n8939)
         );
  AOI21_X1 U10243 ( .B1(n9363), .B2(n8997), .A(n8939), .ZN(n8940) );
  OAI21_X1 U10244 ( .B1(n8941), .B2(n8999), .A(n8940), .ZN(P1_U3227) );
  INV_X1 U10245 ( .A(n8942), .ZN(n8946) );
  NAND2_X1 U10246 ( .A1(n4968), .A2(n8945), .ZN(n8943) );
  AOI22_X1 U10247 ( .A1(n8946), .A2(n8945), .B1(n8944), .B2(n8943), .ZN(n8951)
         );
  AOI22_X1 U10248 ( .A1(n8991), .A2(n9236), .B1(P1_REG3_REG_20__SCAN_IN), .B2(
        P1_U3084), .ZN(n8948) );
  NAND2_X1 U10249 ( .A1(n8979), .A2(n9237), .ZN(n8947) );
  OAI211_X1 U10250 ( .C1(n8981), .C2(n9229), .A(n8948), .B(n8947), .ZN(n8949)
         );
  AOI21_X1 U10251 ( .B1(n9381), .B2(n8997), .A(n8949), .ZN(n8950) );
  OAI21_X1 U10252 ( .B1(n8951), .B2(n8999), .A(n8950), .ZN(P1_U3231) );
  AOI21_X1 U10253 ( .B1(n6631), .B2(n8953), .A(n8954), .ZN(n8957) );
  INV_X1 U10254 ( .A(n8954), .ZN(n8955) );
  OAI22_X1 U10255 ( .A1(n8957), .A2(n8956), .B1(n8955), .B2(n6631), .ZN(n8958)
         );
  NAND2_X1 U10256 ( .A1(n8958), .A2(n8976), .ZN(n8963) );
  AOI22_X1 U10257 ( .A1(n9203), .A2(n8991), .B1(P1_REG3_REG_22__SCAN_IN), .B2(
        P1_U3084), .ZN(n8959) );
  OAI21_X1 U10258 ( .B1(n8960), .B2(n8995), .A(n8959), .ZN(n8961) );
  AOI21_X1 U10259 ( .B1(n9197), .B2(n8992), .A(n8961), .ZN(n8962) );
  OAI211_X1 U10260 ( .C1(n9199), .C2(n8985), .A(n8963), .B(n8962), .ZN(
        P1_U3233) );
  INV_X1 U10261 ( .A(n9269), .ZN(n9393) );
  INV_X1 U10262 ( .A(n8966), .ZN(n8970) );
  AOI21_X1 U10263 ( .B1(n8966), .B2(n8964), .A(n8965), .ZN(n8967) );
  NOR2_X1 U10264 ( .A1(n8967), .A2(n8999), .ZN(n8968) );
  OAI21_X1 U10265 ( .B1(n8970), .B2(n8969), .A(n8968), .ZN(n8975) );
  NAND2_X1 U10266 ( .A1(n8979), .A2(n9004), .ZN(n8971) );
  NAND2_X1 U10267 ( .A1(P1_U3084), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9066) );
  OAI211_X1 U10268 ( .C1(n9264), .C2(n8972), .A(n8971), .B(n9066), .ZN(n8973)
         );
  AOI21_X1 U10269 ( .B1(n9268), .B2(n8992), .A(n8973), .ZN(n8974) );
  OAI211_X1 U10270 ( .C1(n9393), .C2(n8985), .A(n8975), .B(n8974), .ZN(
        P1_U3236) );
  AOI22_X1 U10271 ( .A1(n9166), .A2(n8979), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3084), .ZN(n8980) );
  OAI21_X1 U10272 ( .B1(n8981), .B2(n9136), .A(n8980), .ZN(n8982) );
  AOI21_X1 U10273 ( .B1(n8991), .B2(n9142), .A(n8982), .ZN(n8983) );
  OAI211_X1 U10274 ( .C1(n4618), .C2(n8985), .A(n8984), .B(n8983), .ZN(
        P1_U3238) );
  NAND2_X1 U10275 ( .A1(n8987), .A2(n8986), .ZN(n8988) );
  XOR2_X1 U10276 ( .A(n8989), .B(n8988), .Z(n9000) );
  AOI21_X1 U10277 ( .B1(n8991), .B2(n9288), .A(n8990), .ZN(n8994) );
  NAND2_X1 U10278 ( .A1(n8992), .A2(n9320), .ZN(n8993) );
  OAI211_X1 U10279 ( .C1(n9828), .C2(n8995), .A(n8994), .B(n8993), .ZN(n8996)
         );
  AOI21_X1 U10280 ( .B1(n9408), .B2(n8997), .A(n8996), .ZN(n8998) );
  OAI21_X1 U10281 ( .B1(n9000), .B2(n8999), .A(n8998), .ZN(P1_U3239) );
  MUX2_X1 U10282 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9001), .S(P1_U4006), .Z(
        P1_U3585) );
  MUX2_X1 U10283 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n9105), .S(P1_U4006), .Z(
        P1_U3584) );
  MUX2_X1 U10284 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9002), .S(P1_U4006), .Z(
        P1_U3583) );
  MUX2_X1 U10285 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9142), .S(P1_U4006), .Z(
        P1_U3582) );
  MUX2_X1 U10286 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9156), .S(P1_U4006), .Z(
        P1_U3581) );
  MUX2_X1 U10287 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9166), .S(P1_U4006), .Z(
        P1_U3580) );
  MUX2_X1 U10288 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9183), .S(P1_U4006), .Z(
        P1_U3579) );
  MUX2_X1 U10289 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9203), .S(P1_U4006), .Z(
        P1_U3578) );
  MUX2_X1 U10290 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9190), .S(P1_U4006), .Z(
        P1_U3577) );
  MUX2_X1 U10291 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9236), .S(P1_U4006), .Z(
        P1_U3576) );
  MUX2_X1 U10292 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9003), .S(P1_U4006), .Z(
        P1_U3575) );
  MUX2_X1 U10293 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9237), .S(P1_U4006), .Z(
        P1_U3574) );
  MUX2_X1 U10294 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9286), .S(P1_U4006), .Z(
        P1_U3573) );
  MUX2_X1 U10295 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9004), .S(P1_U4006), .Z(
        P1_U3572) );
  MUX2_X1 U10296 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9288), .S(P1_U4006), .Z(
        P1_U3571) );
  MUX2_X1 U10297 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n9005), .S(P1_U4006), .Z(
        P1_U3570) );
  MUX2_X1 U10298 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n9006), .S(P1_U4006), .Z(
        P1_U3569) );
  MUX2_X1 U10299 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9007), .S(P1_U4006), .Z(
        P1_U3568) );
  MUX2_X1 U10300 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n9008), .S(P1_U4006), .Z(
        P1_U3567) );
  MUX2_X1 U10301 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n9009), .S(P1_U4006), .Z(
        P1_U3566) );
  MUX2_X1 U10302 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n9010), .S(P1_U4006), .Z(
        P1_U3565) );
  MUX2_X1 U10303 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n9011), .S(P1_U4006), .Z(
        P1_U3564) );
  MUX2_X1 U10304 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n9012), .S(P1_U4006), .Z(
        P1_U3563) );
  MUX2_X1 U10305 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n9013), .S(P1_U4006), .Z(
        P1_U3562) );
  MUX2_X1 U10306 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n9014), .S(P1_U4006), .Z(
        P1_U3561) );
  MUX2_X1 U10307 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n9015), .S(P1_U4006), .Z(
        P1_U3560) );
  MUX2_X1 U10308 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n9016), .S(P1_U4006), .Z(
        P1_U3559) );
  MUX2_X1 U10309 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n9017), .S(P1_U4006), .Z(
        P1_U3558) );
  MUX2_X1 U10310 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n9018), .S(P1_U4006), .Z(
        P1_U3557) );
  MUX2_X1 U10311 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n6440), .S(P1_U4006), .Z(
        P1_U3556) );
  MUX2_X1 U10312 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n7361), .S(P1_U4006), .Z(
        P1_U3555) );
  NAND2_X1 U10313 ( .A1(n9894), .A2(P1_ADDR_REG_1__SCAN_IN), .ZN(n9029) );
  AOI22_X1 U10314 ( .A1(n9931), .A2(n9019), .B1(P1_REG3_REG_1__SCAN_IN), .B2(
        P1_U3084), .ZN(n9028) );
  OAI211_X1 U10315 ( .C1(n9022), .C2(n9021), .A(n9941), .B(n9020), .ZN(n9027)
         );
  OAI211_X1 U10316 ( .C1(n9025), .C2(n9024), .A(n9938), .B(n9023), .ZN(n9026)
         );
  NAND4_X1 U10317 ( .A1(n9029), .A2(n9028), .A3(n9027), .A4(n9026), .ZN(
        P1_U3242) );
  NOR2_X1 U10318 ( .A1(n9030), .A2(n9036), .ZN(n9032) );
  NAND2_X1 U10319 ( .A1(P1_REG2_REG_16__SCAN_IN), .A2(n9053), .ZN(n9033) );
  OAI21_X1 U10320 ( .B1(n9053), .B2(P1_REG2_REG_16__SCAN_IN), .A(n9033), .ZN(
        n9034) );
  AOI211_X1 U10321 ( .C1(n4467), .C2(n9034), .A(n9048), .B(n9886), .ZN(n9047)
         );
  NOR2_X1 U10322 ( .A1(n9036), .A2(n9035), .ZN(n9038) );
  NOR2_X1 U10323 ( .A1(n9038), .A2(n9037), .ZN(n9040) );
  XNOR2_X1 U10324 ( .A(n9053), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n9039) );
  NOR2_X1 U10325 ( .A1(n9040), .A2(n9039), .ZN(n9052) );
  AOI211_X1 U10326 ( .C1(n9040), .C2(n9039), .A(n9052), .B(n9902), .ZN(n9046)
         );
  NAND2_X1 U10327 ( .A1(n9894), .A2(P1_ADDR_REG_16__SCAN_IN), .ZN(n9043) );
  INV_X1 U10328 ( .A(n9041), .ZN(n9042) );
  OAI211_X1 U10329 ( .C1(n9922), .C2(n9044), .A(n9043), .B(n9042), .ZN(n9045)
         );
  OR3_X1 U10330 ( .A1(n9047), .A2(n9046), .A3(n9045), .ZN(P1_U3257) );
  INV_X1 U10331 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n9062) );
  AOI21_X1 U10332 ( .B1(n9053), .B2(P1_REG2_REG_16__SCAN_IN), .A(n9048), .ZN(
        n9051) );
  NAND2_X1 U10333 ( .A1(P1_REG2_REG_17__SCAN_IN), .A2(n9069), .ZN(n9049) );
  OAI21_X1 U10334 ( .B1(n9069), .B2(P1_REG2_REG_17__SCAN_IN), .A(n9049), .ZN(
        n9050) );
  NOR2_X1 U10335 ( .A1(n9051), .A2(n9050), .ZN(n9068) );
  AOI211_X1 U10336 ( .C1(n9051), .C2(n9050), .A(n9068), .B(n9886), .ZN(n9060)
         );
  AOI21_X1 U10337 ( .B1(n9053), .B2(P1_REG1_REG_16__SCAN_IN), .A(n9052), .ZN(
        n9055) );
  XNOR2_X1 U10338 ( .A(n9069), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n9054) );
  NOR2_X1 U10339 ( .A1(n9055), .A2(n9054), .ZN(n9063) );
  AOI211_X1 U10340 ( .C1(n9055), .C2(n9054), .A(n9063), .B(n9902), .ZN(n9059)
         );
  INV_X1 U10341 ( .A(n9069), .ZN(n9057) );
  NAND2_X1 U10342 ( .A1(P1_REG3_REG_17__SCAN_IN), .A2(P1_U3084), .ZN(n9056) );
  OAI21_X1 U10343 ( .B1(n9922), .B2(n9057), .A(n9056), .ZN(n9058) );
  NOR3_X1 U10344 ( .A1(n9060), .A2(n9059), .A3(n9058), .ZN(n9061) );
  OAI21_X1 U10345 ( .B1(n9945), .B2(n9062), .A(n9061), .ZN(P1_U3258) );
  INV_X1 U10346 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n9077) );
  XOR2_X1 U10347 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9080), .Z(n9065) );
  AOI21_X1 U10348 ( .B1(n9069), .B2(P1_REG1_REG_17__SCAN_IN), .A(n9063), .ZN(
        n9064) );
  NAND2_X1 U10349 ( .A1(n9065), .A2(n9064), .ZN(n9079) );
  OAI21_X1 U10350 ( .B1(n9065), .B2(n9064), .A(n9079), .ZN(n9075) );
  INV_X1 U10351 ( .A(n9080), .ZN(n9067) );
  OAI21_X1 U10352 ( .B1(n9922), .B2(n9067), .A(n9066), .ZN(n9074) );
  NAND2_X1 U10353 ( .A1(n9080), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9070) );
  OAI21_X1 U10354 ( .B1(n9080), .B2(P1_REG2_REG_18__SCAN_IN), .A(n9070), .ZN(
        n9071) );
  AOI211_X1 U10355 ( .C1(n9072), .C2(n9071), .A(n9078), .B(n9886), .ZN(n9073)
         );
  AOI211_X1 U10356 ( .C1(n9938), .C2(n9075), .A(n9074), .B(n9073), .ZN(n9076)
         );
  OAI21_X1 U10357 ( .B1(n9945), .B2(n9077), .A(n9076), .ZN(P1_U3259) );
  INV_X1 U10358 ( .A(n9085), .ZN(n9083) );
  OAI21_X1 U10359 ( .B1(n9080), .B2(P1_REG1_REG_18__SCAN_IN), .A(n9079), .ZN(
        n9081) );
  XNOR2_X1 U10360 ( .A(n9081), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n9084) );
  OAI21_X1 U10361 ( .B1(n9084), .B2(n9902), .A(n9922), .ZN(n9082) );
  AOI21_X1 U10362 ( .B1(n9083), .B2(n9941), .A(n9082), .ZN(n9088) );
  AOI22_X1 U10363 ( .A1(n9085), .A2(n9941), .B1(n9938), .B2(n9084), .ZN(n9087)
         );
  MUX2_X1 U10364 ( .A(n9088), .B(n9087), .S(n9086), .Z(n9090) );
  OAI211_X1 U10365 ( .C1(n4715), .C2(n9945), .A(n9090), .B(n9089), .ZN(
        P1_U3260) );
  NAND2_X1 U10366 ( .A1(n9099), .A2(n9098), .ZN(n9092) );
  XNOR2_X1 U10367 ( .A(n9091), .B(n9092), .ZN(n9329) );
  NAND2_X1 U10368 ( .A1(n9094), .A2(n9093), .ZN(n9332) );
  NOR2_X1 U10369 ( .A1(n9332), .A2(n9321), .ZN(n9101) );
  NOR2_X1 U10370 ( .A1(n9095), .A2(n9972), .ZN(n9096) );
  AOI211_X1 U10371 ( .C1(n9970), .C2(P1_REG2_REG_31__SCAN_IN), .A(n9101), .B(
        n9096), .ZN(n9097) );
  OAI21_X1 U10372 ( .B1(n9329), .B2(n9324), .A(n9097), .ZN(P1_U3261) );
  XNOR2_X1 U10373 ( .A(n9099), .B(n9098), .ZN(n9333) );
  NOR2_X1 U10374 ( .A1(n9099), .A2(n9972), .ZN(n9100) );
  AOI211_X1 U10375 ( .C1(n9970), .C2(P1_REG2_REG_30__SCAN_IN), .A(n9101), .B(
        n9100), .ZN(n9102) );
  OAI21_X1 U10376 ( .B1(n9324), .B2(n9333), .A(n9102), .ZN(P1_U3262) );
  AOI22_X1 U10377 ( .A1(n9142), .A2(n9287), .B1(n9105), .B2(n9285), .ZN(n9106)
         );
  AOI21_X1 U10378 ( .B1(n9108), .B2(n9107), .A(n4459), .ZN(n9340) );
  NAND2_X1 U10379 ( .A1(n9340), .A2(n9109), .ZN(n9116) );
  AOI21_X1 U10380 ( .B1(n9341), .B2(n9118), .A(n9110), .ZN(n9342) );
  INV_X1 U10381 ( .A(n9341), .ZN(n9113) );
  AOI22_X1 U10382 ( .A1(n9111), .A2(n9969), .B1(P1_REG2_REG_28__SCAN_IN), .B2(
        n9321), .ZN(n9112) );
  OAI21_X1 U10383 ( .B1(n9113), .B2(n9972), .A(n9112), .ZN(n9114) );
  AOI21_X1 U10384 ( .B1(n9342), .B2(n9952), .A(n9114), .ZN(n9115) );
  OAI211_X1 U10385 ( .C1(n9970), .C2(n9344), .A(n9116), .B(n9115), .ZN(
        P1_U3263) );
  XNOR2_X1 U10386 ( .A(n9117), .B(n9125), .ZN(n9350) );
  INV_X1 U10387 ( .A(n9118), .ZN(n9119) );
  AOI21_X1 U10388 ( .B1(n9346), .B2(n9134), .A(n9119), .ZN(n9347) );
  INV_X1 U10389 ( .A(n9346), .ZN(n9122) );
  AOI22_X1 U10390 ( .A1(n9120), .A2(n9969), .B1(P1_REG2_REG_27__SCAN_IN), .B2(
        n9321), .ZN(n9121) );
  OAI21_X1 U10391 ( .B1(n9122), .B2(n9972), .A(n9121), .ZN(n9131) );
  AOI211_X1 U10392 ( .C1(n9125), .C2(n9124), .A(n9844), .B(n9123), .ZN(n9129)
         );
  OAI22_X1 U10393 ( .A1(n9127), .A2(n9960), .B1(n9126), .B2(n9959), .ZN(n9128)
         );
  NOR2_X1 U10394 ( .A1(n9129), .A2(n9128), .ZN(n9349) );
  NOR2_X1 U10395 ( .A1(n9349), .A2(n9321), .ZN(n9130) );
  OAI21_X1 U10396 ( .B1(n9350), .B2(n9308), .A(n9132), .ZN(P1_U3264) );
  XOR2_X1 U10397 ( .A(n9140), .B(n9133), .Z(n9355) );
  INV_X1 U10398 ( .A(n9134), .ZN(n9135) );
  AOI21_X1 U10399 ( .B1(n9351), .B2(n9148), .A(n9135), .ZN(n9352) );
  INV_X1 U10400 ( .A(n9136), .ZN(n9137) );
  AOI22_X1 U10401 ( .A1(n9137), .A2(n9969), .B1(P1_REG2_REG_26__SCAN_IN), .B2(
        n9321), .ZN(n9138) );
  OAI21_X1 U10402 ( .B1(n4618), .B2(n9972), .A(n9138), .ZN(n9145) );
  OAI21_X1 U10403 ( .B1(n4599), .B2(n4598), .A(n9141), .ZN(n9143) );
  AOI222_X1 U10404 ( .A1(n9963), .A2(n9143), .B1(n9142), .B2(n9285), .C1(n9166), .C2(n9287), .ZN(n9354) );
  NOR2_X1 U10405 ( .A1(n9354), .A2(n9321), .ZN(n9144) );
  AOI211_X1 U10406 ( .C1(n9352), .C2(n9952), .A(n9145), .B(n9144), .ZN(n9146)
         );
  OAI21_X1 U10407 ( .B1(n9355), .B2(n9308), .A(n9146), .ZN(P1_U3265) );
  XOR2_X1 U10408 ( .A(n9154), .B(n9147), .Z(n9360) );
  INV_X1 U10409 ( .A(n9169), .ZN(n9149) );
  AOI21_X1 U10410 ( .B1(n9356), .B2(n9149), .A(n4619), .ZN(n9357) );
  AOI22_X1 U10411 ( .A1(n9150), .A2(n9969), .B1(P1_REG2_REG_25__SCAN_IN), .B2(
        n9321), .ZN(n9151) );
  OAI21_X1 U10412 ( .B1(n9152), .B2(n9972), .A(n9151), .ZN(n9160) );
  OAI211_X1 U10413 ( .C1(n9155), .C2(n9154), .A(n9153), .B(n9963), .ZN(n9158)
         );
  AOI22_X1 U10414 ( .A1(n9156), .A2(n9285), .B1(n9287), .B2(n9183), .ZN(n9157)
         );
  NOR2_X1 U10415 ( .A1(n9359), .A2(n9321), .ZN(n9159) );
  AOI211_X1 U10416 ( .C1(n9357), .C2(n9952), .A(n9160), .B(n9159), .ZN(n9161)
         );
  OAI21_X1 U10417 ( .B1(n9360), .B2(n9308), .A(n9161), .ZN(P1_U3266) );
  XOR2_X1 U10418 ( .A(n9162), .B(n9164), .Z(n9365) );
  OAI211_X1 U10419 ( .C1(n9165), .C2(n9164), .A(n9163), .B(n9963), .ZN(n9168)
         );
  AOI22_X1 U10420 ( .A1(n9166), .A2(n9285), .B1(n9287), .B2(n9203), .ZN(n9167)
         );
  NAND2_X1 U10421 ( .A1(n9168), .A2(n9167), .ZN(n9361) );
  INV_X1 U10422 ( .A(n9179), .ZN(n9170) );
  AOI211_X1 U10423 ( .C1(n9363), .C2(n9170), .A(n10034), .B(n9169), .ZN(n9362)
         );
  NAND2_X1 U10424 ( .A1(n9362), .A2(n9301), .ZN(n9174) );
  INV_X1 U10425 ( .A(n9171), .ZN(n9172) );
  AOI22_X1 U10426 ( .A1(n9172), .A2(n9969), .B1(P1_REG2_REG_24__SCAN_IN), .B2(
        n9321), .ZN(n9173) );
  OAI211_X1 U10427 ( .C1(n9175), .C2(n9972), .A(n9174), .B(n9173), .ZN(n9176)
         );
  AOI21_X1 U10428 ( .B1(n9361), .B2(n9836), .A(n9176), .ZN(n9177) );
  OAI21_X1 U10429 ( .B1(n9365), .B2(n9308), .A(n9177), .ZN(P1_U3267) );
  XNOR2_X1 U10430 ( .A(n9178), .B(n9187), .ZN(n9370) );
  AOI21_X1 U10431 ( .B1(n9366), .B2(n9195), .A(n9179), .ZN(n9367) );
  INV_X1 U10432 ( .A(n9180), .ZN(n9181) );
  AOI22_X1 U10433 ( .A1(n9181), .A2(n9969), .B1(n9321), .B2(
        P1_REG2_REG_23__SCAN_IN), .ZN(n9182) );
  OAI21_X1 U10434 ( .B1(n4623), .B2(n9972), .A(n9182), .ZN(n9192) );
  AND2_X1 U10435 ( .A1(n9183), .A2(n9285), .ZN(n9189) );
  INV_X1 U10436 ( .A(n9184), .ZN(n9185) );
  AOI211_X1 U10437 ( .C1(n9187), .C2(n9186), .A(n9844), .B(n9185), .ZN(n9188)
         );
  AOI211_X1 U10438 ( .C1(n9287), .C2(n9190), .A(n9189), .B(n9188), .ZN(n9369)
         );
  NOR2_X1 U10439 ( .A1(n9369), .A2(n9321), .ZN(n9191) );
  AOI211_X1 U10440 ( .C1(n9367), .C2(n9952), .A(n9192), .B(n9191), .ZN(n9193)
         );
  OAI21_X1 U10441 ( .B1(n9370), .B2(n9308), .A(n9193), .ZN(P1_U3268) );
  XOR2_X1 U10442 ( .A(n9194), .B(n9201), .Z(n9375) );
  INV_X1 U10443 ( .A(n9195), .ZN(n9196) );
  AOI21_X1 U10444 ( .B1(n9371), .B2(n9216), .A(n9196), .ZN(n9372) );
  AOI22_X1 U10445 ( .A1(n9321), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n9969), .B2(
        n9197), .ZN(n9198) );
  OAI21_X1 U10446 ( .B1(n9199), .B2(n9972), .A(n9198), .ZN(n9205) );
  XOR2_X1 U10447 ( .A(n9201), .B(n9200), .Z(n9202) );
  AOI222_X1 U10448 ( .A1(n9236), .A2(n9287), .B1(n9203), .B2(n9285), .C1(n9963), .C2(n9202), .ZN(n9374) );
  NOR2_X1 U10449 ( .A1(n9374), .A2(n9321), .ZN(n9204) );
  AOI211_X1 U10450 ( .C1(n9372), .C2(n9952), .A(n9205), .B(n9204), .ZN(n9206)
         );
  OAI21_X1 U10451 ( .B1(n9375), .B2(n9308), .A(n9206), .ZN(P1_U3269) );
  XNOR2_X1 U10452 ( .A(n9207), .B(n9213), .ZN(n9380) );
  NAND2_X1 U10453 ( .A1(n9209), .A2(n9208), .ZN(n9212) );
  INV_X1 U10454 ( .A(n9210), .ZN(n9211) );
  AOI21_X1 U10455 ( .B1(n9213), .B2(n9212), .A(n9211), .ZN(n9214) );
  OAI222_X1 U10456 ( .A1(n9960), .A2(n9215), .B1(n9959), .B2(n9246), .C1(n9844), .C2(n9214), .ZN(n9376) );
  INV_X1 U10457 ( .A(n9227), .ZN(n9218) );
  INV_X1 U10458 ( .A(n9216), .ZN(n9217) );
  AOI211_X1 U10459 ( .C1(n9378), .C2(n9218), .A(n10034), .B(n9217), .ZN(n9377)
         );
  NAND2_X1 U10460 ( .A1(n9377), .A2(n9301), .ZN(n9222) );
  INV_X1 U10461 ( .A(n9219), .ZN(n9220) );
  AOI22_X1 U10462 ( .A1(n9321), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n9969), .B2(
        n9220), .ZN(n9221) );
  OAI211_X1 U10463 ( .C1(n9223), .C2(n9972), .A(n9222), .B(n9221), .ZN(n9224)
         );
  AOI21_X1 U10464 ( .B1(n9376), .B2(n9836), .A(n9224), .ZN(n9225) );
  OAI21_X1 U10465 ( .B1(n9380), .B2(n9308), .A(n9225), .ZN(P1_U3270) );
  XOR2_X1 U10466 ( .A(n9233), .B(n9226), .Z(n9385) );
  INV_X1 U10467 ( .A(n9247), .ZN(n9228) );
  AOI21_X1 U10468 ( .B1(n9381), .B2(n9228), .A(n9227), .ZN(n9382) );
  INV_X1 U10469 ( .A(n9229), .ZN(n9230) );
  AOI22_X1 U10470 ( .A1(n9321), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9969), .B2(
        n9230), .ZN(n9231) );
  OAI21_X1 U10471 ( .B1(n9232), .B2(n9972), .A(n9231), .ZN(n9239) );
  XNOR2_X1 U10472 ( .A(n9234), .B(n9233), .ZN(n9235) );
  AOI222_X1 U10473 ( .A1(n9237), .A2(n9287), .B1(n9236), .B2(n9285), .C1(n9963), .C2(n9235), .ZN(n9384) );
  NOR2_X1 U10474 ( .A1(n9384), .A2(n9321), .ZN(n9238) );
  AOI211_X1 U10475 ( .C1(n9382), .C2(n9952), .A(n9239), .B(n9238), .ZN(n9240)
         );
  OAI21_X1 U10476 ( .B1(n9308), .B2(n9385), .A(n9240), .ZN(P1_U3271) );
  XNOR2_X1 U10477 ( .A(n9241), .B(n9243), .ZN(n9390) );
  AOI22_X1 U10478 ( .A1(n9388), .A2(n9848), .B1(n9970), .B2(
        P1_REG2_REG_19__SCAN_IN), .ZN(n9254) );
  XOR2_X1 U10479 ( .A(n9243), .B(n9242), .Z(n9245) );
  OAI222_X1 U10480 ( .A1(n9960), .A2(n9246), .B1(n9245), .B2(n9844), .C1(n9959), .C2(n9244), .ZN(n9386) );
  AOI211_X1 U10481 ( .C1(n9388), .C2(n4463), .A(n10034), .B(n9247), .ZN(n9387)
         );
  INV_X1 U10482 ( .A(n9387), .ZN(n9251) );
  OAI22_X1 U10483 ( .A1(n9251), .A2(n9250), .B1(n9249), .B2(n9248), .ZN(n9252)
         );
  OAI21_X1 U10484 ( .B1(n9386), .B2(n9252), .A(n9836), .ZN(n9253) );
  OAI211_X1 U10485 ( .C1(n9390), .C2(n9308), .A(n9254), .B(n9253), .ZN(
        P1_U3272) );
  AND2_X1 U10486 ( .A1(n9255), .A2(n9258), .ZN(n9256) );
  OR2_X1 U10487 ( .A1(n9257), .A2(n9256), .ZN(n9391) );
  INV_X1 U10488 ( .A(n9258), .ZN(n9259) );
  NAND3_X1 U10489 ( .A1(n9261), .A2(n9260), .A3(n9259), .ZN(n9262) );
  AOI21_X1 U10490 ( .B1(n9263), .B2(n9262), .A(n9844), .ZN(n9266) );
  OAI22_X1 U10491 ( .A1(n9264), .A2(n9960), .B1(n9959), .B2(n9299), .ZN(n9265)
         );
  OR2_X1 U10492 ( .A1(n9266), .A2(n9265), .ZN(n9395) );
  AOI21_X1 U10493 ( .B1(n9277), .B2(n9269), .A(n10034), .ZN(n9267) );
  NAND2_X1 U10494 ( .A1(n9267), .A2(n4463), .ZN(n9392) );
  AOI22_X1 U10495 ( .A1(n9970), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9969), .B2(
        n9268), .ZN(n9271) );
  NAND2_X1 U10496 ( .A1(n9269), .A2(n9848), .ZN(n9270) );
  OAI211_X1 U10497 ( .C1(n9392), .C2(n9272), .A(n9271), .B(n9270), .ZN(n9273)
         );
  AOI21_X1 U10498 ( .B1(n9395), .B2(n9836), .A(n9273), .ZN(n9274) );
  OAI21_X1 U10499 ( .B1(n9391), .B2(n9308), .A(n9274), .ZN(P1_U3273) );
  XNOR2_X1 U10500 ( .A(n9276), .B(n9275), .ZN(n9402) );
  INV_X1 U10501 ( .A(n9300), .ZN(n9278) );
  AOI21_X1 U10502 ( .B1(n9398), .B2(n9278), .A(n4624), .ZN(n9399) );
  AOI22_X1 U10503 ( .A1(n9321), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9969), .B2(
        n9279), .ZN(n9280) );
  OAI21_X1 U10504 ( .B1(n9281), .B2(n9972), .A(n9280), .ZN(n9290) );
  XNOR2_X1 U10505 ( .A(n9283), .B(n9282), .ZN(n9284) );
  AOI222_X1 U10506 ( .A1(n9288), .A2(n9287), .B1(n9286), .B2(n9285), .C1(n9963), .C2(n9284), .ZN(n9401) );
  NOR2_X1 U10507 ( .A1(n9401), .A2(n9321), .ZN(n9289) );
  AOI211_X1 U10508 ( .C1(n9399), .C2(n9952), .A(n9290), .B(n9289), .ZN(n9291)
         );
  OAI21_X1 U10509 ( .B1(n9308), .B2(n9402), .A(n9291), .ZN(P1_U3274) );
  XNOR2_X1 U10510 ( .A(n9292), .B(n9296), .ZN(n9407) );
  INV_X1 U10511 ( .A(n9293), .ZN(n9294) );
  AOI21_X1 U10512 ( .B1(n9296), .B2(n9295), .A(n9294), .ZN(n9297) );
  OAI222_X1 U10513 ( .A1(n9960), .A2(n9299), .B1(n9959), .B2(n9298), .C1(n9844), .C2(n9297), .ZN(n9403) );
  AOI211_X1 U10514 ( .C1(n9405), .C2(n9319), .A(n10034), .B(n9300), .ZN(n9404)
         );
  NAND2_X1 U10515 ( .A1(n9404), .A2(n9301), .ZN(n9304) );
  AOI22_X1 U10516 ( .A1(n9321), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n9969), .B2(
        n9302), .ZN(n9303) );
  OAI211_X1 U10517 ( .C1(n9305), .C2(n9972), .A(n9304), .B(n9303), .ZN(n9306)
         );
  AOI21_X1 U10518 ( .B1(n9403), .B2(n9836), .A(n9306), .ZN(n9307) );
  OAI21_X1 U10519 ( .B1(n9308), .B2(n9407), .A(n9307), .ZN(P1_U3275) );
  XNOR2_X1 U10520 ( .A(n9310), .B(n9309), .ZN(n9316) );
  OAI22_X1 U10521 ( .A1(n9311), .A2(n9960), .B1(n9959), .B2(n9828), .ZN(n9315)
         );
  XNOR2_X1 U10522 ( .A(n9313), .B(n9312), .ZN(n9413) );
  NOR2_X1 U10523 ( .A1(n9413), .A2(n9966), .ZN(n9314) );
  AOI211_X1 U10524 ( .C1(n9963), .C2(n9316), .A(n9315), .B(n9314), .ZN(n9412)
         );
  INV_X1 U10525 ( .A(n9413), .ZN(n9326) );
  NAND2_X1 U10526 ( .A1(n9317), .A2(n9408), .ZN(n9318) );
  NAND2_X1 U10527 ( .A1(n9319), .A2(n9318), .ZN(n9409) );
  AOI22_X1 U10528 ( .A1(n9321), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n9969), .B2(
        n9320), .ZN(n9323) );
  NAND2_X1 U10529 ( .A1(n9408), .A2(n9848), .ZN(n9322) );
  OAI211_X1 U10530 ( .C1(n9409), .C2(n9324), .A(n9323), .B(n9322), .ZN(n9325)
         );
  AOI21_X1 U10531 ( .B1(n9326), .B2(n9953), .A(n9325), .ZN(n9327) );
  OAI21_X1 U10532 ( .B1(n9412), .B2(n9321), .A(n9327), .ZN(P1_U3276) );
  NAND2_X1 U10533 ( .A1(n9091), .A2(n10010), .ZN(n9328) );
  OAI211_X1 U10534 ( .C1(n9329), .C2(n10034), .A(n9328), .B(n9332), .ZN(n9420)
         );
  MUX2_X1 U10535 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n9420), .S(n4392), .Z(
        P1_U3554) );
  NAND2_X1 U10536 ( .A1(n9330), .A2(n10010), .ZN(n9331) );
  OAI211_X1 U10537 ( .C1(n9333), .C2(n10034), .A(n9332), .B(n9331), .ZN(n9421)
         );
  MUX2_X1 U10538 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n9421), .S(n4392), .Z(
        P1_U3553) );
  NAND2_X1 U10539 ( .A1(n9334), .A2(n10030), .ZN(n9339) );
  AOI21_X1 U10540 ( .B1(n10010), .B2(n9336), .A(n9335), .ZN(n9337) );
  MUX2_X1 U10541 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n9422), .S(n4392), .Z(
        P1_U3552) );
  NAND2_X1 U10542 ( .A1(n9340), .A2(n10030), .ZN(n9345) );
  AOI22_X1 U10543 ( .A1(n9342), .A2(n10011), .B1(n10010), .B2(n9341), .ZN(
        n9343) );
  NAND3_X1 U10544 ( .A1(n9345), .A2(n9344), .A3(n9343), .ZN(n9423) );
  MUX2_X1 U10545 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n9423), .S(n4392), .Z(
        P1_U3551) );
  AOI22_X1 U10546 ( .A1(n9347), .A2(n10011), .B1(n10010), .B2(n9346), .ZN(
        n9348) );
  OAI211_X1 U10547 ( .C1(n9350), .C2(n9418), .A(n9349), .B(n9348), .ZN(n9424)
         );
  MUX2_X1 U10548 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9424), .S(n4392), .Z(
        P1_U3550) );
  AOI22_X1 U10549 ( .A1(n9352), .A2(n10011), .B1(n10010), .B2(n9351), .ZN(
        n9353) );
  OAI211_X1 U10550 ( .C1(n9355), .C2(n9418), .A(n9354), .B(n9353), .ZN(n9425)
         );
  MUX2_X1 U10551 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9425), .S(n4392), .Z(
        P1_U3549) );
  AOI22_X1 U10552 ( .A1(n9357), .A2(n10011), .B1(n10010), .B2(n9356), .ZN(
        n9358) );
  OAI211_X1 U10553 ( .C1(n9360), .C2(n9418), .A(n9359), .B(n9358), .ZN(n9426)
         );
  MUX2_X1 U10554 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9426), .S(n4392), .Z(
        P1_U3548) );
  AOI211_X1 U10555 ( .C1(n10010), .C2(n9363), .A(n9362), .B(n9361), .ZN(n9364)
         );
  OAI21_X1 U10556 ( .B1(n9365), .B2(n9418), .A(n9364), .ZN(n9427) );
  MUX2_X1 U10557 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9427), .S(n4392), .Z(
        P1_U3547) );
  AOI22_X1 U10558 ( .A1(n9367), .A2(n10011), .B1(n10010), .B2(n9366), .ZN(
        n9368) );
  OAI211_X1 U10559 ( .C1(n9370), .C2(n9418), .A(n9369), .B(n9368), .ZN(n9428)
         );
  MUX2_X1 U10560 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9428), .S(n4392), .Z(
        P1_U3546) );
  AOI22_X1 U10561 ( .A1(n9372), .A2(n10011), .B1(n10010), .B2(n9371), .ZN(
        n9373) );
  OAI211_X1 U10562 ( .C1(n9375), .C2(n9418), .A(n9374), .B(n9373), .ZN(n9429)
         );
  MUX2_X1 U10563 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9429), .S(n4392), .Z(
        P1_U3545) );
  AOI211_X1 U10564 ( .C1(n10010), .C2(n9378), .A(n9377), .B(n9376), .ZN(n9379)
         );
  OAI21_X1 U10565 ( .B1(n9380), .B2(n9418), .A(n9379), .ZN(n9430) );
  MUX2_X1 U10566 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9430), .S(n4392), .Z(
        P1_U3544) );
  AOI22_X1 U10567 ( .A1(n9382), .A2(n10011), .B1(n10010), .B2(n9381), .ZN(
        n9383) );
  OAI211_X1 U10568 ( .C1(n9385), .C2(n9418), .A(n9384), .B(n9383), .ZN(n9431)
         );
  MUX2_X1 U10569 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9431), .S(n4392), .Z(
        P1_U3543) );
  AOI211_X1 U10570 ( .C1(n10010), .C2(n9388), .A(n9387), .B(n9386), .ZN(n9389)
         );
  OAI21_X1 U10571 ( .B1(n9390), .B2(n9418), .A(n9389), .ZN(n9432) );
  MUX2_X1 U10572 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9432), .S(n4392), .Z(
        P1_U3542) );
  OR2_X1 U10573 ( .A1(n9391), .A2(n9418), .ZN(n9397) );
  OAI21_X1 U10574 ( .B1(n9393), .B2(n10032), .A(n9392), .ZN(n9394) );
  NOR2_X1 U10575 ( .A1(n9395), .A2(n9394), .ZN(n9396) );
  NAND2_X1 U10576 ( .A1(n9397), .A2(n9396), .ZN(n9433) );
  MUX2_X1 U10577 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9433), .S(n4392), .Z(
        P1_U3541) );
  AOI22_X1 U10578 ( .A1(n9399), .A2(n10011), .B1(n10010), .B2(n9398), .ZN(
        n9400) );
  OAI211_X1 U10579 ( .C1(n9402), .C2(n9418), .A(n9401), .B(n9400), .ZN(n9434)
         );
  MUX2_X1 U10580 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9434), .S(n4392), .Z(
        P1_U3540) );
  AOI211_X1 U10581 ( .C1(n10010), .C2(n9405), .A(n9404), .B(n9403), .ZN(n9406)
         );
  OAI21_X1 U10582 ( .B1(n9418), .B2(n9407), .A(n9406), .ZN(n9435) );
  MUX2_X1 U10583 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9435), .S(n4392), .Z(
        P1_U3539) );
  OAI22_X1 U10584 ( .A1(n9409), .A2(n10034), .B1(n4615), .B2(n10032), .ZN(
        n9410) );
  INV_X1 U10585 ( .A(n9410), .ZN(n9411) );
  OAI211_X1 U10586 ( .C1(n9413), .C2(n10015), .A(n9412), .B(n9411), .ZN(n9436)
         );
  MUX2_X1 U10587 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n9436), .S(n4392), .Z(
        P1_U3538) );
  AOI211_X1 U10588 ( .C1(n10010), .C2(n9416), .A(n9415), .B(n9414), .ZN(n9417)
         );
  OAI21_X1 U10589 ( .B1(n9419), .B2(n9418), .A(n9417), .ZN(n9437) );
  MUX2_X1 U10590 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n9437), .S(n4392), .Z(
        P1_U3537) );
  MUX2_X1 U10591 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n9420), .S(n10042), .Z(
        P1_U3522) );
  MUX2_X1 U10592 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n9421), .S(n10042), .Z(
        P1_U3521) );
  MUX2_X1 U10593 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n9423), .S(n10042), .Z(
        P1_U3519) );
  MUX2_X1 U10594 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9424), .S(n10042), .Z(
        P1_U3518) );
  MUX2_X1 U10595 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9425), .S(n10042), .Z(
        P1_U3517) );
  MUX2_X1 U10596 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9426), .S(n10042), .Z(
        P1_U3516) );
  MUX2_X1 U10597 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9427), .S(n10042), .Z(
        P1_U3515) );
  MUX2_X1 U10598 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9428), .S(n10042), .Z(
        P1_U3514) );
  MUX2_X1 U10599 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9429), .S(n10042), .Z(
        P1_U3513) );
  MUX2_X1 U10600 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9430), .S(n10042), .Z(
        P1_U3512) );
  MUX2_X1 U10601 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9431), .S(n10042), .Z(
        P1_U3511) );
  MUX2_X1 U10602 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9432), .S(n10042), .Z(
        P1_U3510) );
  MUX2_X1 U10603 ( .A(n9433), .B(P1_REG0_REG_18__SCAN_IN), .S(n10040), .Z(
        P1_U3508) );
  MUX2_X1 U10604 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9434), .S(n10042), .Z(
        P1_U3505) );
  MUX2_X1 U10605 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n9435), .S(n10042), .Z(
        P1_U3502) );
  MUX2_X1 U10606 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n9436), .S(n10042), .Z(
        P1_U3499) );
  MUX2_X1 U10607 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n9437), .S(n10042), .Z(
        P1_U3496) );
  NOR4_X1 U10608 ( .A1(n9438), .A2(P1_IR_REG_30__SCAN_IN), .A3(P1_U3084), .A4(
        n9439), .ZN(n9440) );
  AOI21_X1 U10609 ( .B1(n9730), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9440), .ZN(
        n9441) );
  OAI21_X1 U10610 ( .B1(n5133), .B2(n9445), .A(n9441), .ZN(P1_U3322) );
  OAI222_X1 U10611 ( .A1(n9449), .A2(n9571), .B1(n9445), .B2(n9444), .C1(
        P1_U3084), .C2(n9442), .ZN(P1_U3323) );
  OAI222_X1 U10612 ( .A1(n9449), .A2(n9448), .B1(P1_U3084), .B2(n9447), .C1(
        n9446), .C2(n9445), .ZN(P1_U3324) );
  NAND2_X1 U10613 ( .A1(n9730), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n9451) );
  OAI211_X1 U10614 ( .C1(n9453), .C2(n9452), .A(n9451), .B(n9450), .ZN(
        P1_U3325) );
  NOR2_X1 U10615 ( .A1(keyinput63), .A2(keyinput67), .ZN(n9454) );
  NAND3_X1 U10616 ( .A1(keyinput25), .A2(keyinput127), .A3(n9454), .ZN(n9455)
         );
  NOR3_X1 U10617 ( .A1(keyinput53), .A2(keyinput76), .A3(n9455), .ZN(n9515) );
  NOR4_X1 U10618 ( .A1(keyinput45), .A2(keyinput17), .A3(keyinput115), .A4(
        keyinput71), .ZN(n9456) );
  NAND3_X1 U10619 ( .A1(keyinput32), .A2(keyinput35), .A3(n9456), .ZN(n9464)
         );
  NAND2_X1 U10620 ( .A1(keyinput95), .A2(keyinput3), .ZN(n9457) );
  NOR3_X1 U10621 ( .A1(keyinput9), .A2(keyinput56), .A3(n9457), .ZN(n9462) );
  NOR4_X1 U10622 ( .A1(keyinput34), .A2(keyinput30), .A3(keyinput27), .A4(
        keyinput117), .ZN(n9461) );
  INV_X1 U10623 ( .A(keyinput18), .ZN(n9458) );
  NOR4_X1 U10624 ( .A1(keyinput82), .A2(keyinput121), .A3(keyinput33), .A4(
        n9458), .ZN(n9460) );
  AND4_X1 U10625 ( .A1(keyinput99), .A2(keyinput105), .A3(keyinput123), .A4(
        keyinput122), .ZN(n9459) );
  NAND4_X1 U10626 ( .A1(n9462), .A2(n9461), .A3(n9460), .A4(n9459), .ZN(n9463)
         );
  NOR4_X1 U10627 ( .A1(keyinput109), .A2(keyinput42), .A3(n9464), .A4(n9463), 
        .ZN(n9514) );
  INV_X1 U10628 ( .A(keyinput39), .ZN(n9465) );
  NAND4_X1 U10629 ( .A1(keyinput44), .A2(keyinput2), .A3(keyinput23), .A4(
        n9465), .ZN(n9512) );
  NOR2_X1 U10630 ( .A1(keyinput37), .A2(keyinput78), .ZN(n9466) );
  NAND3_X1 U10631 ( .A1(keyinput94), .A2(keyinput116), .A3(n9466), .ZN(n9511)
         );
  NOR2_X1 U10632 ( .A1(keyinput114), .A2(keyinput0), .ZN(n9467) );
  NAND3_X1 U10633 ( .A1(keyinput80), .A2(keyinput40), .A3(n9467), .ZN(n9468)
         );
  NOR3_X1 U10634 ( .A1(keyinput61), .A2(keyinput41), .A3(n9468), .ZN(n9476) );
  NAND4_X1 U10635 ( .A1(keyinput73), .A2(keyinput58), .A3(keyinput108), .A4(
        keyinput1), .ZN(n9474) );
  NOR2_X1 U10636 ( .A1(keyinput14), .A2(keyinput87), .ZN(n9469) );
  NAND3_X1 U10637 ( .A1(keyinput103), .A2(keyinput46), .A3(n9469), .ZN(n9473)
         );
  OR4_X1 U10638 ( .A1(keyinput36), .A2(keyinput48), .A3(keyinput38), .A4(
        keyinput4), .ZN(n9472) );
  NOR2_X1 U10639 ( .A1(keyinput20), .A2(keyinput83), .ZN(n9470) );
  NAND3_X1 U10640 ( .A1(keyinput6), .A2(keyinput13), .A3(n9470), .ZN(n9471) );
  NOR4_X1 U10641 ( .A1(n9474), .A2(n9473), .A3(n9472), .A4(n9471), .ZN(n9475)
         );
  NAND4_X1 U10642 ( .A1(keyinput12), .A2(keyinput93), .A3(n9476), .A4(n9475), 
        .ZN(n9510) );
  NAND2_X1 U10643 ( .A1(keyinput120), .A2(keyinput15), .ZN(n9477) );
  NOR3_X1 U10644 ( .A1(keyinput10), .A2(keyinput88), .A3(n9477), .ZN(n9478) );
  NAND3_X1 U10645 ( .A1(keyinput84), .A2(keyinput29), .A3(n9478), .ZN(n9491)
         );
  NOR2_X1 U10646 ( .A1(keyinput59), .A2(keyinput112), .ZN(n9479) );
  NAND3_X1 U10647 ( .A1(keyinput85), .A2(keyinput81), .A3(n9479), .ZN(n9480)
         );
  NOR3_X1 U10648 ( .A1(keyinput19), .A2(keyinput26), .A3(n9480), .ZN(n9489) );
  INV_X1 U10649 ( .A(keyinput65), .ZN(n9481) );
  NAND4_X1 U10650 ( .A1(keyinput22), .A2(keyinput119), .A3(keyinput111), .A4(
        n9481), .ZN(n9487) );
  NOR2_X1 U10651 ( .A1(keyinput7), .A2(keyinput72), .ZN(n9482) );
  NAND3_X1 U10652 ( .A1(keyinput113), .A2(keyinput64), .A3(n9482), .ZN(n9486)
         );
  OR4_X1 U10653 ( .A1(keyinput55), .A2(keyinput49), .A3(keyinput96), .A4(
        keyinput75), .ZN(n9485) );
  INV_X1 U10654 ( .A(keyinput21), .ZN(n9483) );
  NAND4_X1 U10655 ( .A1(keyinput24), .A2(keyinput74), .A3(keyinput70), .A4(
        n9483), .ZN(n9484) );
  NOR4_X1 U10656 ( .A1(n9487), .A2(n9486), .A3(n9485), .A4(n9484), .ZN(n9488)
         );
  NAND4_X1 U10657 ( .A1(keyinput62), .A2(keyinput101), .A3(n9489), .A4(n9488), 
        .ZN(n9490) );
  NOR4_X1 U10658 ( .A1(keyinput69), .A2(keyinput31), .A3(n9491), .A4(n9490), 
        .ZN(n9508) );
  NAND2_X1 U10659 ( .A1(keyinput50), .A2(keyinput52), .ZN(n9492) );
  NOR3_X1 U10660 ( .A1(keyinput57), .A2(keyinput91), .A3(n9492), .ZN(n9507) );
  INV_X1 U10661 ( .A(keyinput106), .ZN(n9493) );
  NOR4_X1 U10662 ( .A1(keyinput79), .A2(keyinput104), .A3(keyinput89), .A4(
        n9493), .ZN(n9506) );
  NAND2_X1 U10663 ( .A1(keyinput11), .A2(keyinput51), .ZN(n9494) );
  NOR3_X1 U10664 ( .A1(keyinput8), .A2(keyinput97), .A3(n9494), .ZN(n9495) );
  NAND3_X1 U10665 ( .A1(keyinput47), .A2(keyinput66), .A3(n9495), .ZN(n9504)
         );
  NOR4_X1 U10666 ( .A1(keyinput118), .A2(keyinput92), .A3(keyinput16), .A4(
        keyinput98), .ZN(n9502) );
  NAND3_X1 U10667 ( .A1(keyinput90), .A2(keyinput100), .A3(keyinput43), .ZN(
        n9496) );
  NOR2_X1 U10668 ( .A1(keyinput5), .A2(n9496), .ZN(n9501) );
  NAND2_X1 U10669 ( .A1(keyinput125), .A2(keyinput28), .ZN(n9497) );
  NOR3_X1 U10670 ( .A1(keyinput54), .A2(keyinput102), .A3(n9497), .ZN(n9500)
         );
  INV_X1 U10671 ( .A(keyinput77), .ZN(n9498) );
  NOR4_X1 U10672 ( .A1(keyinput86), .A2(keyinput60), .A3(keyinput110), .A4(
        n9498), .ZN(n9499) );
  NAND4_X1 U10673 ( .A1(n9502), .A2(n9501), .A3(n9500), .A4(n9499), .ZN(n9503)
         );
  NOR4_X1 U10674 ( .A1(keyinput107), .A2(keyinput68), .A3(n9504), .A4(n9503), 
        .ZN(n9505) );
  NAND4_X1 U10675 ( .A1(n9508), .A2(n9507), .A3(n9506), .A4(n9505), .ZN(n9509)
         );
  NOR4_X1 U10676 ( .A1(n9512), .A2(n9511), .A3(n9510), .A4(n9509), .ZN(n9513)
         );
  NAND4_X1 U10677 ( .A1(keyinput124), .A2(n9515), .A3(n9514), .A4(n9513), .ZN(
        n9516) );
  AND2_X1 U10678 ( .A1(n9516), .A2(keyinput126), .ZN(n9729) );
  INV_X1 U10679 ( .A(P1_D_REG_20__SCAN_IN), .ZN(n9978) );
  AOI22_X1 U10680 ( .A1(n7074), .A2(keyinput7), .B1(n9978), .B2(keyinput64), 
        .ZN(n9517) );
  OAI221_X1 U10681 ( .B1(n7074), .B2(keyinput7), .C1(n9978), .C2(keyinput64), 
        .A(n9517), .ZN(n9526) );
  AOI22_X1 U10682 ( .A1(n9520), .A2(keyinput72), .B1(n9519), .B2(keyinput119), 
        .ZN(n9518) );
  OAI221_X1 U10683 ( .B1(n9520), .B2(keyinput72), .C1(n9519), .C2(keyinput119), 
        .A(n9518), .ZN(n9525) );
  AOI22_X1 U10684 ( .A1(n5749), .A2(keyinput22), .B1(keyinput111), .B2(n6203), 
        .ZN(n9521) );
  OAI221_X1 U10685 ( .B1(n5749), .B2(keyinput22), .C1(n6203), .C2(keyinput111), 
        .A(n9521), .ZN(n9524) );
  INV_X1 U10686 ( .A(P1_D_REG_29__SCAN_IN), .ZN(n9976) );
  AOI22_X1 U10687 ( .A1(n6948), .A2(keyinput65), .B1(n9976), .B2(keyinput21), 
        .ZN(n9522) );
  OAI221_X1 U10688 ( .B1(n6948), .B2(keyinput65), .C1(n9976), .C2(keyinput21), 
        .A(n9522), .ZN(n9523) );
  NOR4_X1 U10689 ( .A1(n9526), .A2(n9525), .A3(n9524), .A4(n9523), .ZN(n9564)
         );
  AOI22_X1 U10690 ( .A1(n7105), .A2(keyinput70), .B1(n5538), .B2(keyinput55), 
        .ZN(n9527) );
  OAI221_X1 U10691 ( .B1(n7105), .B2(keyinput70), .C1(n5538), .C2(keyinput55), 
        .A(n9527), .ZN(n9537) );
  INV_X1 U10692 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n9529) );
  INV_X1 U10693 ( .A(P1_D_REG_18__SCAN_IN), .ZN(n9980) );
  AOI22_X1 U10694 ( .A1(n9529), .A2(keyinput24), .B1(n9980), .B2(keyinput74), 
        .ZN(n9528) );
  OAI221_X1 U10695 ( .B1(n9529), .B2(keyinput24), .C1(n9980), .C2(keyinput74), 
        .A(n9528), .ZN(n9536) );
  AOI22_X1 U10696 ( .A1(n9531), .A2(keyinput75), .B1(n5852), .B2(keyinput15), 
        .ZN(n9530) );
  OAI221_X1 U10697 ( .B1(n9531), .B2(keyinput75), .C1(n5852), .C2(keyinput15), 
        .A(n9530), .ZN(n9535) );
  INV_X1 U10698 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n10224) );
  XOR2_X1 U10699 ( .A(n10224), .B(keyinput49), .Z(n9533) );
  XNOR2_X1 U10700 ( .A(P2_IR_REG_3__SCAN_IN), .B(keyinput96), .ZN(n9532) );
  NAND2_X1 U10701 ( .A1(n9533), .A2(n9532), .ZN(n9534) );
  NOR4_X1 U10702 ( .A1(n9537), .A2(n9536), .A3(n9535), .A4(n9534), .ZN(n9563)
         );
  AOI22_X1 U10703 ( .A1(n5927), .A2(keyinput31), .B1(n5869), .B2(keyinput85), 
        .ZN(n9538) );
  OAI221_X1 U10704 ( .B1(n5927), .B2(keyinput31), .C1(n5869), .C2(keyinput85), 
        .A(n9538), .ZN(n9548) );
  INV_X1 U10705 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n10201) );
  AOI22_X1 U10706 ( .A1(n9077), .A2(keyinput29), .B1(n10201), .B2(keyinput10), 
        .ZN(n9539) );
  OAI221_X1 U10707 ( .B1(n9077), .B2(keyinput29), .C1(n10201), .C2(keyinput10), 
        .A(n9539), .ZN(n9547) );
  INV_X1 U10708 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n9541) );
  AOI22_X1 U10709 ( .A1(n9542), .A2(keyinput88), .B1(keyinput84), .B2(n9541), 
        .ZN(n9540) );
  OAI221_X1 U10710 ( .B1(n9542), .B2(keyinput88), .C1(n9541), .C2(keyinput84), 
        .A(n9540), .ZN(n9546) );
  XNOR2_X1 U10711 ( .A(P1_IR_REG_28__SCAN_IN), .B(keyinput69), .ZN(n9544) );
  XNOR2_X1 U10712 ( .A(SI_4_), .B(keyinput120), .ZN(n9543) );
  NAND2_X1 U10713 ( .A1(n9544), .A2(n9543), .ZN(n9545) );
  NOR4_X1 U10714 ( .A1(n9548), .A2(n9547), .A3(n9546), .A4(n9545), .ZN(n9562)
         );
  INV_X1 U10715 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n9550) );
  AOI22_X1 U10716 ( .A1(n9551), .A2(keyinput59), .B1(n9550), .B2(keyinput81), 
        .ZN(n9549) );
  OAI221_X1 U10717 ( .B1(n9551), .B2(keyinput59), .C1(n9550), .C2(keyinput81), 
        .A(n9549), .ZN(n9560) );
  AOI22_X1 U10718 ( .A1(n9553), .A2(keyinput112), .B1(keyinput62), .B2(n5914), 
        .ZN(n9552) );
  OAI221_X1 U10719 ( .B1(n9553), .B2(keyinput112), .C1(n5914), .C2(keyinput62), 
        .A(n9552), .ZN(n9559) );
  INV_X1 U10720 ( .A(P2_D_REG_20__SCAN_IN), .ZN(n10112) );
  AOI22_X1 U10721 ( .A1(n10112), .A2(keyinput101), .B1(P2_U3152), .B2(
        keyinput19), .ZN(n9554) );
  OAI221_X1 U10722 ( .B1(n10112), .B2(keyinput101), .C1(P2_U3152), .C2(
        keyinput19), .A(n9554), .ZN(n9558) );
  INV_X1 U10723 ( .A(P1_D_REG_23__SCAN_IN), .ZN(n9977) );
  AOI22_X1 U10724 ( .A1(n9556), .A2(keyinput26), .B1(n9977), .B2(keyinput106), 
        .ZN(n9555) );
  OAI221_X1 U10725 ( .B1(n9556), .B2(keyinput26), .C1(n9977), .C2(keyinput106), 
        .A(n9555), .ZN(n9557) );
  NOR4_X1 U10726 ( .A1(n9560), .A2(n9559), .A3(n9558), .A4(n9557), .ZN(n9561)
         );
  NAND4_X1 U10727 ( .A1(n9564), .A2(n9563), .A3(n9562), .A4(n9561), .ZN(n9727)
         );
  INV_X1 U10728 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n9567) );
  AOI22_X1 U10729 ( .A1(n9567), .A2(keyinput104), .B1(n9566), .B2(keyinput79), 
        .ZN(n9565) );
  OAI221_X1 U10730 ( .B1(n9567), .B2(keyinput104), .C1(n9566), .C2(keyinput79), 
        .A(n9565), .ZN(n9577) );
  AOI22_X1 U10731 ( .A1(n9569), .A2(keyinput89), .B1(keyinput57), .B2(n6297), 
        .ZN(n9568) );
  OAI221_X1 U10732 ( .B1(n9569), .B2(keyinput89), .C1(n6297), .C2(keyinput57), 
        .A(n9568), .ZN(n9576) );
  AOI22_X1 U10733 ( .A1(n9571), .A2(keyinput52), .B1(n6856), .B2(keyinput91), 
        .ZN(n9570) );
  OAI221_X1 U10734 ( .B1(n9571), .B2(keyinput52), .C1(n6856), .C2(keyinput91), 
        .A(n9570), .ZN(n9575) );
  INV_X1 U10735 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n9573) );
  AOI22_X1 U10736 ( .A1(n9573), .A2(keyinput50), .B1(keyinput43), .B2(n6272), 
        .ZN(n9572) );
  OAI221_X1 U10737 ( .B1(n9573), .B2(keyinput50), .C1(n6272), .C2(keyinput43), 
        .A(n9572), .ZN(n9574) );
  NOR4_X1 U10738 ( .A1(n9577), .A2(n9576), .A3(n9575), .A4(n9574), .ZN(n9618)
         );
  INV_X1 U10739 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n9579) );
  INV_X1 U10740 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n10249) );
  AOI22_X1 U10741 ( .A1(n9579), .A2(keyinput90), .B1(keyinput16), .B2(n10249), 
        .ZN(n9578) );
  OAI221_X1 U10742 ( .B1(n9579), .B2(keyinput90), .C1(n10249), .C2(keyinput16), 
        .A(n9578), .ZN(n9588) );
  INV_X1 U10743 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n10002) );
  AOI22_X1 U10744 ( .A1(n10002), .A2(keyinput92), .B1(n9581), .B2(keyinput100), 
        .ZN(n9580) );
  OAI221_X1 U10745 ( .B1(n10002), .B2(keyinput92), .C1(n9581), .C2(keyinput100), .A(n9580), .ZN(n9587) );
  XOR2_X1 U10746 ( .A(n6843), .B(keyinput118), .Z(n9585) );
  XOR2_X1 U10747 ( .A(n7188), .B(keyinput47), .Z(n9584) );
  XNOR2_X1 U10748 ( .A(P1_IR_REG_23__SCAN_IN), .B(keyinput5), .ZN(n9583) );
  XNOR2_X1 U10749 ( .A(SI_0_), .B(keyinput98), .ZN(n9582) );
  NAND4_X1 U10750 ( .A1(n9585), .A2(n9584), .A3(n9583), .A4(n9582), .ZN(n9586)
         );
  NOR3_X1 U10751 ( .A1(n9588), .A2(n9587), .A3(n9586), .ZN(n9617) );
  INV_X1 U10752 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n9590) );
  AOI22_X1 U10753 ( .A1(n9591), .A2(keyinput66), .B1(keyinput107), .B2(n9590), 
        .ZN(n9589) );
  OAI221_X1 U10754 ( .B1(n9591), .B2(keyinput66), .C1(n9590), .C2(keyinput107), 
        .A(n9589), .ZN(n9602) );
  AOI22_X1 U10755 ( .A1(n6028), .A2(keyinput68), .B1(n9593), .B2(keyinput51), 
        .ZN(n9592) );
  OAI221_X1 U10756 ( .B1(n6028), .B2(keyinput68), .C1(n9593), .C2(keyinput51), 
        .A(n9592), .ZN(n9601) );
  INV_X1 U10757 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n9596) );
  INV_X1 U10758 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n9595) );
  AOI22_X1 U10759 ( .A1(n9596), .A2(keyinput8), .B1(n9595), .B2(keyinput11), 
        .ZN(n9594) );
  OAI221_X1 U10760 ( .B1(n9596), .B2(keyinput8), .C1(n9595), .C2(keyinput11), 
        .A(n9594), .ZN(n9600) );
  INV_X1 U10761 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n9598) );
  AOI22_X1 U10762 ( .A1(n5403), .A2(keyinput97), .B1(keyinput86), .B2(n9598), 
        .ZN(n9597) );
  OAI221_X1 U10763 ( .B1(n5403), .B2(keyinput97), .C1(n9598), .C2(keyinput86), 
        .A(n9597), .ZN(n9599) );
  NOR4_X1 U10764 ( .A1(n9602), .A2(n9601), .A3(n9600), .A4(n9599), .ZN(n9616)
         );
  INV_X1 U10765 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n9783) );
  AOI22_X1 U10766 ( .A1(n9783), .A2(keyinput60), .B1(n9604), .B2(keyinput110), 
        .ZN(n9603) );
  OAI221_X1 U10767 ( .B1(n9783), .B2(keyinput60), .C1(n9604), .C2(keyinput110), 
        .A(n9603), .ZN(n9614) );
  INV_X1 U10768 ( .A(SI_11_), .ZN(n9606) );
  AOI22_X1 U10769 ( .A1(n9606), .A2(keyinput77), .B1(keyinput54), .B2(n4792), 
        .ZN(n9605) );
  OAI221_X1 U10770 ( .B1(n9606), .B2(keyinput77), .C1(n4792), .C2(keyinput54), 
        .A(n9605), .ZN(n9613) );
  INV_X1 U10771 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n9877) );
  AOI22_X1 U10772 ( .A1(n9877), .A2(keyinput28), .B1(n9608), .B2(keyinput125), 
        .ZN(n9607) );
  OAI221_X1 U10773 ( .B1(n9877), .B2(keyinput28), .C1(n9608), .C2(keyinput125), 
        .A(n9607), .ZN(n9612) );
  INV_X1 U10774 ( .A(P1_D_REG_11__SCAN_IN), .ZN(n9982) );
  AOI22_X1 U10775 ( .A1(n9982), .A2(keyinput124), .B1(keyinput102), .B2(n9610), 
        .ZN(n9609) );
  OAI221_X1 U10776 ( .B1(n9982), .B2(keyinput124), .C1(n9610), .C2(keyinput102), .A(n9609), .ZN(n9611) );
  NOR4_X1 U10777 ( .A1(n9614), .A2(n9613), .A3(n9612), .A4(n9611), .ZN(n9615)
         );
  NAND4_X1 U10778 ( .A1(n9618), .A2(n9617), .A3(n9616), .A4(n9615), .ZN(n9726)
         );
  INV_X1 U10779 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n9620) );
  AOI22_X1 U10780 ( .A1(n6842), .A2(keyinput87), .B1(n9620), .B2(keyinput73), 
        .ZN(n9619) );
  OAI221_X1 U10781 ( .B1(n6842), .B2(keyinput87), .C1(n9620), .C2(keyinput73), 
        .A(n9619), .ZN(n9631) );
  AOI22_X1 U10782 ( .A1(n9623), .A2(keyinput103), .B1(n9622), .B2(keyinput46), 
        .ZN(n9621) );
  OAI221_X1 U10783 ( .B1(n9623), .B2(keyinput103), .C1(n9622), .C2(keyinput46), 
        .A(n9621), .ZN(n9630) );
  INV_X1 U10784 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n9626) );
  AOI22_X1 U10785 ( .A1(n9626), .A2(keyinput1), .B1(n9625), .B2(keyinput94), 
        .ZN(n9624) );
  OAI221_X1 U10786 ( .B1(n9626), .B2(keyinput1), .C1(n9625), .C2(keyinput94), 
        .A(n9624), .ZN(n9629) );
  AOI22_X1 U10787 ( .A1(n6237), .A2(keyinput58), .B1(keyinput108), .B2(n6215), 
        .ZN(n9627) );
  OAI221_X1 U10788 ( .B1(n6237), .B2(keyinput58), .C1(n6215), .C2(keyinput108), 
        .A(n9627), .ZN(n9628) );
  NOR4_X1 U10789 ( .A1(n9631), .A2(n9630), .A3(n9629), .A4(n9628), .ZN(n9667)
         );
  INV_X1 U10790 ( .A(SI_7_), .ZN(n9633) );
  AOI22_X1 U10791 ( .A1(n9634), .A2(keyinput0), .B1(n9633), .B2(keyinput12), 
        .ZN(n9632) );
  OAI221_X1 U10792 ( .B1(n9634), .B2(keyinput0), .C1(n9633), .C2(keyinput12), 
        .A(n9632), .ZN(n9641) );
  INV_X1 U10793 ( .A(P2_D_REG_31__SCAN_IN), .ZN(n10111) );
  AOI22_X1 U10794 ( .A1(n7018), .A2(keyinput80), .B1(n10111), .B2(keyinput40), 
        .ZN(n9635) );
  OAI221_X1 U10795 ( .B1(n7018), .B2(keyinput80), .C1(n10111), .C2(keyinput40), 
        .A(n9635), .ZN(n9640) );
  INV_X1 U10796 ( .A(P1_D_REG_7__SCAN_IN), .ZN(n9983) );
  INV_X1 U10797 ( .A(P1_D_REG_19__SCAN_IN), .ZN(n9979) );
  AOI22_X1 U10798 ( .A1(n9983), .A2(keyinput41), .B1(keyinput14), .B2(n9979), 
        .ZN(n9636) );
  OAI221_X1 U10799 ( .B1(n9983), .B2(keyinput41), .C1(n9979), .C2(keyinput14), 
        .A(n9636), .ZN(n9639) );
  INV_X1 U10800 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n9818) );
  AOI22_X1 U10801 ( .A1(n5240), .A2(keyinput93), .B1(keyinput61), .B2(n9818), 
        .ZN(n9637) );
  OAI221_X1 U10802 ( .B1(n5240), .B2(keyinput93), .C1(n9818), .C2(keyinput61), 
        .A(n9637), .ZN(n9638) );
  NOR4_X1 U10803 ( .A1(n9641), .A2(n9640), .A3(n9639), .A4(n9638), .ZN(n9666)
         );
  AOI22_X1 U10804 ( .A1(n5822), .A2(keyinput48), .B1(keyinput38), .B2(n8003), 
        .ZN(n9642) );
  OAI221_X1 U10805 ( .B1(n5822), .B2(keyinput48), .C1(n8003), .C2(keyinput38), 
        .A(n9642), .ZN(n9651) );
  INV_X1 U10806 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n10263) );
  AOI22_X1 U10807 ( .A1(n9644), .A2(keyinput83), .B1(keyinput36), .B2(n10263), 
        .ZN(n9643) );
  OAI221_X1 U10808 ( .B1(n9644), .B2(keyinput83), .C1(n10263), .C2(keyinput36), 
        .A(n9643), .ZN(n9650) );
  INV_X1 U10809 ( .A(P1_D_REG_14__SCAN_IN), .ZN(n9981) );
  AOI22_X1 U10810 ( .A1(n9981), .A2(keyinput4), .B1(keyinput113), .B2(n7607), 
        .ZN(n9645) );
  OAI221_X1 U10811 ( .B1(n9981), .B2(keyinput4), .C1(n7607), .C2(keyinput113), 
        .A(n9645), .ZN(n9649) );
  XNOR2_X1 U10812 ( .A(P2_IR_REG_31__SCAN_IN), .B(keyinput13), .ZN(n9647) );
  XNOR2_X1 U10813 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(keyinput20), .ZN(n9646)
         );
  NAND2_X1 U10814 ( .A1(n9647), .A2(n9646), .ZN(n9648) );
  NOR4_X1 U10815 ( .A1(n9651), .A2(n9650), .A3(n9649), .A4(n9648), .ZN(n9665)
         );
  INV_X1 U10816 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n9813) );
  AOI22_X1 U10817 ( .A1(n9813), .A2(keyinput44), .B1(n9653), .B2(keyinput23), 
        .ZN(n9652) );
  OAI221_X1 U10818 ( .B1(n9813), .B2(keyinput44), .C1(n9653), .C2(keyinput23), 
        .A(n9652), .ZN(n9654) );
  INV_X1 U10819 ( .A(n9654), .ZN(n9663) );
  XNOR2_X1 U10820 ( .A(P2_IR_REG_12__SCAN_IN), .B(keyinput116), .ZN(n9657) );
  XNOR2_X1 U10821 ( .A(P2_IR_REG_8__SCAN_IN), .B(keyinput78), .ZN(n9656) );
  XNOR2_X1 U10822 ( .A(keyinput37), .B(P2_REG1_REG_7__SCAN_IN), .ZN(n9655) );
  AND3_X1 U10823 ( .A1(n9657), .A2(n9656), .A3(n9655), .ZN(n9662) );
  INV_X1 U10824 ( .A(P2_D_REG_18__SCAN_IN), .ZN(n10113) );
  XNOR2_X1 U10825 ( .A(n10113), .B(n9465), .ZN(n9661) );
  XNOR2_X1 U10826 ( .A(P1_IR_REG_5__SCAN_IN), .B(keyinput6), .ZN(n9659) );
  XNOR2_X1 U10827 ( .A(keyinput2), .B(P1_REG2_REG_4__SCAN_IN), .ZN(n9658) );
  AND2_X1 U10828 ( .A1(n9659), .A2(n9658), .ZN(n9660) );
  AND4_X1 U10829 ( .A1(n9663), .A2(n9662), .A3(n9661), .A4(n9660), .ZN(n9664)
         );
  NAND4_X1 U10830 ( .A1(n9667), .A2(n9666), .A3(n9665), .A4(n9664), .ZN(n9725)
         );
  AOI22_X1 U10831 ( .A1(n9669), .A2(keyinput42), .B1(keyinput45), .B2(n10256), 
        .ZN(n9668) );
  OAI221_X1 U10832 ( .B1(n9669), .B2(keyinput42), .C1(n10256), .C2(keyinput45), 
        .A(n9668), .ZN(n9679) );
  AOI22_X1 U10833 ( .A1(n9671), .A2(keyinput35), .B1(keyinput115), .B2(n6931), 
        .ZN(n9670) );
  OAI221_X1 U10834 ( .B1(n9671), .B2(keyinput35), .C1(n6931), .C2(keyinput115), 
        .A(n9670), .ZN(n9678) );
  AOI22_X1 U10835 ( .A1(P1_U3084), .A2(keyinput71), .B1(keyinput34), .B2(n9673), .ZN(n9672) );
  OAI221_X1 U10836 ( .B1(P1_U3084), .B2(keyinput71), .C1(n9673), .C2(
        keyinput34), .A(n9672), .ZN(n9677) );
  INV_X1 U10837 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n10264) );
  XOR2_X1 U10838 ( .A(n10264), .B(keyinput17), .Z(n9675) );
  XNOR2_X1 U10839 ( .A(P1_IR_REG_19__SCAN_IN), .B(keyinput32), .ZN(n9674) );
  NAND2_X1 U10840 ( .A1(n9675), .A2(n9674), .ZN(n9676) );
  NOR4_X1 U10841 ( .A1(n9679), .A2(n9678), .A3(n9677), .A4(n9676), .ZN(n9723)
         );
  INV_X1 U10842 ( .A(keyinput126), .ZN(n9681) );
  XNOR2_X1 U10843 ( .A(P2_REG1_REG_21__SCAN_IN), .B(keyinput67), .ZN(n9680) );
  OAI21_X1 U10844 ( .B1(P1_IR_REG_15__SCAN_IN), .B2(n9681), .A(n9680), .ZN(
        n9693) );
  AOI22_X1 U10845 ( .A1(n9684), .A2(keyinput63), .B1(keyinput25), .B2(n9683), 
        .ZN(n9682) );
  OAI221_X1 U10846 ( .B1(n9684), .B2(keyinput63), .C1(n9683), .C2(keyinput25), 
        .A(n9682), .ZN(n9692) );
  INV_X1 U10847 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n10191) );
  AOI22_X1 U10848 ( .A1(n10191), .A2(keyinput76), .B1(n9686), .B2(keyinput109), 
        .ZN(n9685) );
  OAI221_X1 U10849 ( .B1(n10191), .B2(keyinput76), .C1(n9686), .C2(keyinput109), .A(n9685), .ZN(n9691) );
  INV_X1 U10850 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n9688) );
  AOI22_X1 U10851 ( .A1(n9689), .A2(keyinput127), .B1(n9688), .B2(keyinput53), 
        .ZN(n9687) );
  OAI221_X1 U10852 ( .B1(n9689), .B2(keyinput127), .C1(n9688), .C2(keyinput53), 
        .A(n9687), .ZN(n9690) );
  NOR4_X1 U10853 ( .A1(n9693), .A2(n9692), .A3(n9691), .A4(n9690), .ZN(n9722)
         );
  AOI22_X1 U10854 ( .A1(n9696), .A2(keyinput18), .B1(n9695), .B2(keyinput123), 
        .ZN(n9694) );
  OAI221_X1 U10855 ( .B1(n9696), .B2(keyinput18), .C1(n9695), .C2(keyinput123), 
        .A(n9694), .ZN(n9707) );
  INV_X1 U10856 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n9698) );
  AOI22_X1 U10857 ( .A1(n5348), .A2(keyinput105), .B1(keyinput82), .B2(n9698), 
        .ZN(n9697) );
  OAI221_X1 U10858 ( .B1(n5348), .B2(keyinput105), .C1(n9698), .C2(keyinput82), 
        .A(n9697), .ZN(n9706) );
  INV_X1 U10859 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n9700) );
  AOI22_X1 U10860 ( .A1(n5851), .A2(keyinput33), .B1(keyinput114), .B2(n9700), 
        .ZN(n9699) );
  OAI221_X1 U10861 ( .B1(n5851), .B2(keyinput33), .C1(n9700), .C2(keyinput114), 
        .A(n9699), .ZN(n9705) );
  INV_X1 U10862 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n9703) );
  INV_X1 U10863 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n9702) );
  AOI22_X1 U10864 ( .A1(n9703), .A2(keyinput122), .B1(keyinput121), .B2(n9702), 
        .ZN(n9701) );
  OAI221_X1 U10865 ( .B1(n9703), .B2(keyinput122), .C1(n9702), .C2(keyinput121), .A(n9701), .ZN(n9704) );
  NOR4_X1 U10866 ( .A1(n9707), .A2(n9706), .A3(n9705), .A4(n9704), .ZN(n9721)
         );
  AOI22_X1 U10867 ( .A1(n8579), .A2(keyinput56), .B1(keyinput99), .B2(n5967), 
        .ZN(n9708) );
  OAI221_X1 U10868 ( .B1(n8579), .B2(keyinput56), .C1(n5967), .C2(keyinput99), 
        .A(n9708), .ZN(n9719) );
  AOI22_X1 U10869 ( .A1(n6320), .A2(keyinput9), .B1(n9710), .B2(keyinput95), 
        .ZN(n9709) );
  OAI221_X1 U10870 ( .B1(n6320), .B2(keyinput9), .C1(n9710), .C2(keyinput95), 
        .A(n9709), .ZN(n9718) );
  AOI22_X1 U10871 ( .A1(n9713), .A2(keyinput30), .B1(n9712), .B2(keyinput27), 
        .ZN(n9711) );
  OAI221_X1 U10872 ( .B1(n9713), .B2(keyinput30), .C1(n9712), .C2(keyinput27), 
        .A(n9711), .ZN(n9717) );
  XNOR2_X1 U10873 ( .A(P1_IR_REG_24__SCAN_IN), .B(keyinput3), .ZN(n9715) );
  XNOR2_X1 U10874 ( .A(keyinput117), .B(P2_REG1_REG_12__SCAN_IN), .ZN(n9714)
         );
  NAND2_X1 U10875 ( .A1(n9715), .A2(n9714), .ZN(n9716) );
  NOR4_X1 U10876 ( .A1(n9719), .A2(n9718), .A3(n9717), .A4(n9716), .ZN(n9720)
         );
  NAND4_X1 U10877 ( .A1(n9723), .A2(n9722), .A3(n9721), .A4(n9720), .ZN(n9724)
         );
  NOR4_X1 U10878 ( .A1(n9727), .A2(n9726), .A3(n9725), .A4(n9724), .ZN(n9728)
         );
  OAI21_X1 U10879 ( .B1(n9729), .B2(n4784), .A(n9728), .ZN(n9735) );
  AOI222_X1 U10880 ( .A1(n9733), .A2(n9732), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9731), .C1(P2_DATAO_REG_14__SCAN_IN), .C2(n9730), .ZN(n9734) );
  XOR2_X1 U10881 ( .A(n9735), .B(n9734), .Z(P1_U3339) );
  MUX2_X1 U10882 ( .A(n9736), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3353) );
  AOI22_X1 U10883 ( .A1(n10058), .A2(P2_ADDR_REG_1__SCAN_IN), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(P2_U3152), .ZN(n9747) );
  AOI211_X1 U10884 ( .C1(n9739), .C2(n9738), .A(n9737), .B(n10060), .ZN(n9740)
         );
  AOI21_X1 U10885 ( .B1(n9753), .B2(n9741), .A(n9740), .ZN(n9746) );
  AND2_X1 U10886 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n9744) );
  OAI211_X1 U10887 ( .C1(n9744), .C2(n9743), .A(n10057), .B(n9742), .ZN(n9745)
         );
  NAND3_X1 U10888 ( .A1(n9747), .A2(n9746), .A3(n9745), .ZN(P2_U3246) );
  AOI22_X1 U10889 ( .A1(n10058), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3152), .ZN(n9759) );
  AOI211_X1 U10890 ( .C1(n9750), .C2(n9749), .A(n9748), .B(n10060), .ZN(n9751)
         );
  AOI21_X1 U10891 ( .B1(n9753), .B2(n9752), .A(n9751), .ZN(n9758) );
  OAI211_X1 U10892 ( .C1(n9756), .C2(n9755), .A(n10057), .B(n9754), .ZN(n9757)
         );
  NAND3_X1 U10893 ( .A1(n9759), .A2(n9758), .A3(n9757), .ZN(P2_U3247) );
  NOR2_X1 U10894 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n9760) );
  AOI21_X1 U10895 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n9760), .ZN(n10227) );
  NOR2_X1 U10896 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n9761) );
  AOI21_X1 U10897 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n9761), .ZN(n10230) );
  NOR2_X1 U10898 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n9762) );
  AOI21_X1 U10899 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n9762), .ZN(n10233) );
  NOR2_X1 U10900 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n9763) );
  AOI21_X1 U10901 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n9763), .ZN(n10236) );
  NOR2_X1 U10902 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n9764) );
  AOI21_X1 U10903 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n9764), .ZN(n10239) );
  NOR2_X1 U10904 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n9771) );
  XNOR2_X1 U10905 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10271) );
  NAND2_X1 U10906 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n9769) );
  XOR2_X1 U10907 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(P2_ADDR_REG_3__SCAN_IN), .Z(
        n10269) );
  NAND2_X1 U10908 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n9767) );
  XOR2_X1 U10909 ( .A(P2_ADDR_REG_2__SCAN_IN), .B(P1_ADDR_REG_2__SCAN_IN), .Z(
        n10267) );
  AOI21_X1 U10910 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10220) );
  INV_X1 U10911 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n9765) );
  NAND3_X1 U10912 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_1__SCAN_IN), .ZN(n10222) );
  OAI21_X1 U10913 ( .B1(n10220), .B2(n9765), .A(n10222), .ZN(n10266) );
  NAND2_X1 U10914 ( .A1(n10267), .A2(n10266), .ZN(n9766) );
  NAND2_X1 U10915 ( .A1(n9767), .A2(n9766), .ZN(n10268) );
  NAND2_X1 U10916 ( .A1(n10269), .A2(n10268), .ZN(n9768) );
  NAND2_X1 U10917 ( .A1(n9769), .A2(n9768), .ZN(n10270) );
  NOR2_X1 U10918 ( .A1(n10271), .A2(n10270), .ZN(n9770) );
  NOR2_X1 U10919 ( .A1(n9771), .A2(n9770), .ZN(n9772) );
  NOR2_X1 U10920 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n9772), .ZN(n10251) );
  AND2_X1 U10921 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n9772), .ZN(n10252) );
  NOR2_X1 U10922 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n10252), .ZN(n9773) );
  NOR2_X1 U10923 ( .A1(n10251), .A2(n9773), .ZN(n9774) );
  NAND2_X1 U10924 ( .A1(n9774), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n9776) );
  XOR2_X1 U10925 ( .A(n9774), .B(P1_ADDR_REG_6__SCAN_IN), .Z(n10250) );
  NAND2_X1 U10926 ( .A1(n10250), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n9775) );
  NAND2_X1 U10927 ( .A1(n9776), .A2(n9775), .ZN(n9777) );
  NAND2_X1 U10928 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n9777), .ZN(n9779) );
  XOR2_X1 U10929 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n9777), .Z(n10265) );
  NAND2_X1 U10930 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n10265), .ZN(n9778) );
  NAND2_X1 U10931 ( .A1(n9779), .A2(n9778), .ZN(n9780) );
  AND2_X1 U10932 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n9780), .ZN(n9781) );
  XNOR2_X1 U10933 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(n9780), .ZN(n10262) );
  NOR2_X1 U10934 ( .A1(n10263), .A2(n10262), .ZN(n10261) );
  NOR2_X1 U10935 ( .A1(n9782), .A2(n9783), .ZN(n9784) );
  INV_X1 U10936 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n10260) );
  XNOR2_X1 U10937 ( .A(n9783), .B(n9782), .ZN(n10259) );
  NOR2_X1 U10938 ( .A1(n10260), .A2(n10259), .ZN(n10258) );
  NOR2_X1 U10939 ( .A1(n9784), .A2(n10258), .ZN(n10248) );
  NAND2_X1 U10940 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n9785) );
  OAI21_X1 U10941 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n9785), .ZN(n10247) );
  NOR2_X1 U10942 ( .A1(n10248), .A2(n10247), .ZN(n10246) );
  AOI21_X1 U10943 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n10246), .ZN(n10245) );
  NAND2_X1 U10944 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n9786) );
  OAI21_X1 U10945 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n9786), .ZN(n10244) );
  NOR2_X1 U10946 ( .A1(n10245), .A2(n10244), .ZN(n10243) );
  AOI21_X1 U10947 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n10243), .ZN(n10242) );
  NOR2_X1 U10948 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n9787) );
  AOI21_X1 U10949 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n9787), .ZN(n10241) );
  NAND2_X1 U10950 ( .A1(n10242), .A2(n10241), .ZN(n10240) );
  OAI21_X1 U10951 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10240), .ZN(n10238) );
  NAND2_X1 U10952 ( .A1(n10239), .A2(n10238), .ZN(n10237) );
  OAI21_X1 U10953 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n10237), .ZN(n10235) );
  NAND2_X1 U10954 ( .A1(n10236), .A2(n10235), .ZN(n10234) );
  OAI21_X1 U10955 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10234), .ZN(n10232) );
  NAND2_X1 U10956 ( .A1(n10233), .A2(n10232), .ZN(n10231) );
  OAI21_X1 U10957 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n10231), .ZN(n10229) );
  NAND2_X1 U10958 ( .A1(n10230), .A2(n10229), .ZN(n10228) );
  OAI21_X1 U10959 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n10228), .ZN(n10226) );
  NAND2_X1 U10960 ( .A1(n10227), .A2(n10226), .ZN(n10225) );
  OAI21_X1 U10961 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10225), .ZN(n10255) );
  NOR2_X1 U10962 ( .A1(n10256), .A2(n10255), .ZN(n9788) );
  NAND2_X1 U10963 ( .A1(n10256), .A2(n10255), .ZN(n10254) );
  OAI21_X1 U10964 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n9788), .A(n10254), .ZN(
        n9790) );
  XOR2_X1 U10965 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(P1_ADDR_REG_19__SCAN_IN), 
        .Z(n9789) );
  XNOR2_X1 U10966 ( .A(n9790), .B(n9789), .ZN(ADD_1071_U4) );
  OAI21_X1 U10967 ( .B1(n9792), .B2(n10192), .A(n9791), .ZN(n9793) );
  AOI21_X1 U10968 ( .B1(n9794), .B2(n10126), .A(n9793), .ZN(n9814) );
  INV_X1 U10969 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n9795) );
  AOI22_X1 U10970 ( .A1(n10219), .A2(n9814), .B1(n9795), .B2(n10217), .ZN(
        P2_U3550) );
  OAI22_X1 U10971 ( .A1(n9797), .A2(n10194), .B1(n9796), .B2(n10192), .ZN(
        n9799) );
  AOI211_X1 U10972 ( .C1(n10199), .C2(n9800), .A(n9799), .B(n9798), .ZN(n9815)
         );
  AOI22_X1 U10973 ( .A1(n10219), .A2(n9815), .B1(n9801), .B2(n10217), .ZN(
        P2_U3535) );
  OAI22_X1 U10974 ( .A1(n9802), .A2(n10194), .B1(n4637), .B2(n10192), .ZN(
        n9804) );
  AOI211_X1 U10975 ( .C1(n10199), .C2(n9805), .A(n9804), .B(n9803), .ZN(n9817)
         );
  AOI22_X1 U10976 ( .A1(n10219), .A2(n9817), .B1(n6120), .B2(n10217), .ZN(
        P2_U3534) );
  INV_X1 U10977 ( .A(n9806), .ZN(n10184) );
  INV_X1 U10978 ( .A(n9807), .ZN(n9812) );
  OAI22_X1 U10979 ( .A1(n9809), .A2(n10194), .B1(n9808), .B2(n10192), .ZN(
        n9811) );
  AOI211_X1 U10980 ( .C1(n10184), .C2(n9812), .A(n9811), .B(n9810), .ZN(n9819)
         );
  AOI22_X1 U10981 ( .A1(n10219), .A2(n9819), .B1(n6105), .B2(n10217), .ZN(
        P2_U3533) );
  AOI22_X1 U10982 ( .A1(n10202), .A2(n9814), .B1(n9813), .B2(n10200), .ZN(
        P2_U3518) );
  AOI22_X1 U10983 ( .A1(n10202), .A2(n9815), .B1(n6137), .B2(n10200), .ZN(
        P2_U3496) );
  INV_X1 U10984 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n9816) );
  AOI22_X1 U10985 ( .A1(n10202), .A2(n9817), .B1(n9816), .B2(n10200), .ZN(
        P2_U3493) );
  AOI22_X1 U10986 ( .A1(n10202), .A2(n9819), .B1(n9818), .B2(n10200), .ZN(
        P2_U3490) );
  XNOR2_X1 U10987 ( .A(n9820), .B(n9827), .ZN(n9860) );
  OR2_X1 U10988 ( .A1(n9821), .A2(n9857), .ZN(n9822) );
  NAND2_X1 U10989 ( .A1(n9823), .A2(n9822), .ZN(n9858) );
  INV_X1 U10990 ( .A(n9858), .ZN(n9824) );
  AOI22_X1 U10991 ( .A1(n9860), .A2(n9953), .B1(n9952), .B2(n9824), .ZN(n9839)
         );
  NAND2_X1 U10992 ( .A1(n9860), .A2(n9846), .ZN(n9832) );
  OAI21_X1 U10993 ( .B1(n9827), .B2(n9826), .A(n9825), .ZN(n9830) );
  OAI22_X1 U10994 ( .A1(n9845), .A2(n9959), .B1(n9960), .B2(n9828), .ZN(n9829)
         );
  AOI21_X1 U10995 ( .B1(n9830), .B2(n9963), .A(n9829), .ZN(n9831) );
  AND2_X1 U10996 ( .A1(n9832), .A2(n9831), .ZN(n9862) );
  INV_X1 U10997 ( .A(n9862), .ZN(n9837) );
  AOI22_X1 U10998 ( .A1(n9970), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n9969), .B2(
        n9833), .ZN(n9834) );
  OAI21_X1 U10999 ( .B1(n9857), .B2(n9972), .A(n9834), .ZN(n9835) );
  AOI21_X1 U11000 ( .B1(n9837), .B2(n9836), .A(n9835), .ZN(n9838) );
  NAND2_X1 U11001 ( .A1(n9839), .A2(n9838), .ZN(P1_U3278) );
  XOR2_X1 U11002 ( .A(n9841), .B(n9840), .Z(n9873) );
  XOR2_X1 U11003 ( .A(n9842), .B(n9841), .Z(n9843) );
  OAI222_X1 U11004 ( .A1(n9960), .A2(n9845), .B1(n9959), .B2(n9961), .C1(n9844), .C2(n9843), .ZN(n9872) );
  AOI21_X1 U11005 ( .B1(n9873), .B2(n9846), .A(n9872), .ZN(n9856) );
  AOI222_X1 U11006 ( .A1(n9849), .A2(n9848), .B1(n9847), .B2(n9969), .C1(
        P1_REG2_REG_11__SCAN_IN), .C2(n9321), .ZN(n9855) );
  INV_X1 U11007 ( .A(n9850), .ZN(n9851) );
  OAI21_X1 U11008 ( .B1(n9869), .B2(n9852), .A(n9851), .ZN(n9870) );
  INV_X1 U11009 ( .A(n9870), .ZN(n9853) );
  AOI22_X1 U11010 ( .A1(n9873), .A2(n9953), .B1(n9952), .B2(n9853), .ZN(n9854)
         );
  OAI211_X1 U11011 ( .C1(n9970), .C2(n9856), .A(n9855), .B(n9854), .ZN(
        P1_U3280) );
  OAI22_X1 U11012 ( .A1(n9858), .A2(n10034), .B1(n9857), .B2(n10032), .ZN(
        n9859) );
  AOI21_X1 U11013 ( .B1(n9860), .B2(n10039), .A(n9859), .ZN(n9861) );
  AOI22_X1 U11014 ( .A1(n4392), .A2(n9876), .B1(n7300), .B2(n10053), .ZN(
        P1_U3536) );
  INV_X1 U11015 ( .A(n9863), .ZN(n9868) );
  OAI21_X1 U11016 ( .B1(n9865), .B2(n10032), .A(n9864), .ZN(n9867) );
  AOI211_X1 U11017 ( .C1(n10039), .C2(n9868), .A(n9867), .B(n9866), .ZN(n9878)
         );
  AOI22_X1 U11018 ( .A1(n4392), .A2(n9878), .B1(n7211), .B2(n10053), .ZN(
        P1_U3535) );
  OAI22_X1 U11019 ( .A1(n9870), .A2(n10034), .B1(n9869), .B2(n10032), .ZN(
        n9871) );
  AOI211_X1 U11020 ( .C1(n9873), .C2(n10030), .A(n9872), .B(n9871), .ZN(n9880)
         );
  AOI22_X1 U11021 ( .A1(n4392), .A2(n9880), .B1(n9874), .B2(n10053), .ZN(
        P1_U3534) );
  INV_X1 U11022 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n9875) );
  AOI22_X1 U11023 ( .A1(n10042), .A2(n9876), .B1(n9875), .B2(n10040), .ZN(
        P1_U3493) );
  AOI22_X1 U11024 ( .A1(n10042), .A2(n9878), .B1(n9877), .B2(n10040), .ZN(
        P1_U3490) );
  INV_X1 U11025 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n9879) );
  AOI22_X1 U11026 ( .A1(n10042), .A2(n9880), .B1(n9879), .B2(n10040), .ZN(
        P1_U3487) );
  XNOR2_X1 U11027 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U11028 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  AOI21_X1 U11029 ( .B1(n9883), .B2(n9882), .A(n9881), .ZN(n9885) );
  OAI22_X1 U11030 ( .A1(n9886), .A2(n9885), .B1(n9884), .B2(n9922), .ZN(n9887)
         );
  INV_X1 U11031 ( .A(n9887), .ZN(n9897) );
  NAND2_X1 U11032 ( .A1(n9889), .A2(n9888), .ZN(n9890) );
  AOI21_X1 U11033 ( .B1(n9891), .B2(n9890), .A(n9902), .ZN(n9892) );
  AOI211_X1 U11034 ( .C1(P1_ADDR_REG_4__SCAN_IN), .C2(n9894), .A(n9893), .B(
        n9892), .ZN(n9896) );
  NAND3_X1 U11035 ( .A1(n9897), .A2(n9896), .A3(n9895), .ZN(P1_U3245) );
  AND2_X1 U11036 ( .A1(n9899), .A2(n9898), .ZN(n9900) );
  OR3_X1 U11037 ( .A1(n9902), .A2(n9901), .A3(n9900), .ZN(n9905) );
  INV_X1 U11038 ( .A(n9903), .ZN(n9904) );
  OAI211_X1 U11039 ( .C1(n9922), .C2(n9906), .A(n9905), .B(n9904), .ZN(n9907)
         );
  INV_X1 U11040 ( .A(n9907), .ZN(n9913) );
  OAI21_X1 U11041 ( .B1(n9910), .B2(n9909), .A(n9908), .ZN(n9911) );
  NAND2_X1 U11042 ( .A1(n9941), .A2(n9911), .ZN(n9912) );
  OAI211_X1 U11043 ( .C1(n10263), .C2(n9945), .A(n9913), .B(n9912), .ZN(
        P1_U3249) );
  INV_X1 U11044 ( .A(n9914), .ZN(n9915) );
  OAI211_X1 U11045 ( .C1(n9917), .C2(n9916), .A(n9941), .B(n9915), .ZN(n9920)
         );
  INV_X1 U11046 ( .A(n9918), .ZN(n9919) );
  OAI211_X1 U11047 ( .C1(n9922), .C2(n9921), .A(n9920), .B(n9919), .ZN(n9923)
         );
  INV_X1 U11048 ( .A(n9923), .ZN(n9928) );
  XNOR2_X1 U11049 ( .A(n9925), .B(n9924), .ZN(n9926) );
  NAND2_X1 U11050 ( .A1(n9938), .A2(n9926), .ZN(n9927) );
  OAI211_X1 U11051 ( .C1(n10260), .C2(n9945), .A(n9928), .B(n9927), .ZN(
        P1_U3250) );
  INV_X1 U11052 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n9944) );
  AOI21_X1 U11053 ( .B1(n9931), .B2(n9930), .A(n9929), .ZN(n9943) );
  OAI21_X1 U11054 ( .B1(n9934), .B2(n9933), .A(n9932), .ZN(n9940) );
  OAI21_X1 U11055 ( .B1(n9937), .B2(n9936), .A(n9935), .ZN(n9939) );
  AOI22_X1 U11056 ( .A1(n9941), .A2(n9940), .B1(n9939), .B2(n9938), .ZN(n9942)
         );
  OAI211_X1 U11057 ( .C1(n9945), .C2(n9944), .A(n9943), .B(n9942), .ZN(
        P1_U3252) );
  NAND2_X1 U11058 ( .A1(n9947), .A2(n9946), .ZN(n9948) );
  XNOR2_X1 U11059 ( .A(n9948), .B(n9956), .ZN(n9967) );
  INV_X1 U11060 ( .A(n9967), .ZN(n10038) );
  OAI21_X1 U11061 ( .B1(n9950), .B2(n10033), .A(n9949), .ZN(n10035) );
  INV_X1 U11062 ( .A(n10035), .ZN(n9951) );
  AOI22_X1 U11063 ( .A1(n10038), .A2(n9953), .B1(n9952), .B2(n9951), .ZN(n9975) );
  NAND2_X1 U11064 ( .A1(n9955), .A2(n9954), .ZN(n9957) );
  XNOR2_X1 U11065 ( .A(n9957), .B(n9956), .ZN(n9964) );
  OAI22_X1 U11066 ( .A1(n9961), .A2(n9960), .B1(n9959), .B2(n9958), .ZN(n9962)
         );
  AOI21_X1 U11067 ( .B1(n9964), .B2(n9963), .A(n9962), .ZN(n9965) );
  OAI21_X1 U11068 ( .B1(n9967), .B2(n9966), .A(n9965), .ZN(n10036) );
  AOI22_X1 U11069 ( .A1(n9970), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n9969), .B2(
        n9968), .ZN(n9971) );
  OAI21_X1 U11070 ( .B1(n9972), .B2(n10033), .A(n9971), .ZN(n9973) );
  AOI21_X1 U11071 ( .B1(n10036), .B2(n9836), .A(n9973), .ZN(n9974) );
  NAND2_X1 U11072 ( .A1(n9975), .A2(n9974), .ZN(P1_U3282) );
  AND2_X1 U11073 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n9985), .ZN(P1_U3292) );
  AND2_X1 U11074 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n9985), .ZN(P1_U3293) );
  NOR2_X1 U11075 ( .A1(n9984), .A2(n9976), .ZN(P1_U3294) );
  AND2_X1 U11076 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n9985), .ZN(P1_U3295) );
  AND2_X1 U11077 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n9985), .ZN(P1_U3296) );
  AND2_X1 U11078 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n9985), .ZN(P1_U3297) );
  AND2_X1 U11079 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n9985), .ZN(P1_U3298) );
  AND2_X1 U11080 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n9985), .ZN(P1_U3299) );
  NOR2_X1 U11081 ( .A1(n9984), .A2(n9977), .ZN(P1_U3300) );
  AND2_X1 U11082 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n9985), .ZN(P1_U3301) );
  AND2_X1 U11083 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n9985), .ZN(P1_U3302) );
  NOR2_X1 U11084 ( .A1(n9984), .A2(n9978), .ZN(P1_U3303) );
  NOR2_X1 U11085 ( .A1(n9984), .A2(n9979), .ZN(P1_U3304) );
  NOR2_X1 U11086 ( .A1(n9984), .A2(n9980), .ZN(P1_U3305) );
  AND2_X1 U11087 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n9985), .ZN(P1_U3306) );
  AND2_X1 U11088 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n9985), .ZN(P1_U3307) );
  AND2_X1 U11089 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n9985), .ZN(P1_U3308) );
  NOR2_X1 U11090 ( .A1(n9984), .A2(n9981), .ZN(P1_U3309) );
  AND2_X1 U11091 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n9985), .ZN(P1_U3310) );
  AND2_X1 U11092 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n9985), .ZN(P1_U3311) );
  NOR2_X1 U11093 ( .A1(n9984), .A2(n9982), .ZN(P1_U3312) );
  AND2_X1 U11094 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n9985), .ZN(P1_U3313) );
  AND2_X1 U11095 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n9985), .ZN(P1_U3314) );
  AND2_X1 U11096 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n9985), .ZN(P1_U3315) );
  NOR2_X1 U11097 ( .A1(n9984), .A2(n9983), .ZN(P1_U3316) );
  AND2_X1 U11098 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n9985), .ZN(P1_U3317) );
  AND2_X1 U11099 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n9985), .ZN(P1_U3318) );
  AND2_X1 U11100 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n9985), .ZN(P1_U3319) );
  AND2_X1 U11101 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n9985), .ZN(P1_U3320) );
  AND2_X1 U11102 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n9985), .ZN(P1_U3321) );
  OAI21_X1 U11103 ( .B1(n9988), .B2(n9987), .A(n9986), .ZN(P1_U3441) );
  INV_X1 U11104 ( .A(n9989), .ZN(n9994) );
  OAI21_X1 U11105 ( .B1(n9991), .B2(n10032), .A(n9990), .ZN(n9993) );
  AOI211_X1 U11106 ( .C1(n10039), .C2(n9994), .A(n9993), .B(n9992), .ZN(n10044) );
  INV_X1 U11107 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n9995) );
  AOI22_X1 U11108 ( .A1(n10042), .A2(n10044), .B1(n9995), .B2(n10040), .ZN(
        P1_U3457) );
  INV_X1 U11109 ( .A(n9996), .ZN(n9998) );
  OAI22_X1 U11110 ( .A1(n9998), .A2(n10034), .B1(n9997), .B2(n10032), .ZN(
        n10000) );
  AOI211_X1 U11111 ( .C1(n10039), .C2(n10001), .A(n10000), .B(n9999), .ZN(
        n10046) );
  AOI22_X1 U11112 ( .A1(n10042), .A2(n10046), .B1(n10002), .B2(n10040), .ZN(
        P1_U3460) );
  OAI22_X1 U11113 ( .A1(n10004), .A2(n10034), .B1(n10003), .B2(n10032), .ZN(
        n10006) );
  AOI211_X1 U11114 ( .C1(n10039), .C2(n10007), .A(n10006), .B(n10005), .ZN(
        n10048) );
  INV_X1 U11115 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n10008) );
  AOI22_X1 U11116 ( .A1(n10042), .A2(n10048), .B1(n10008), .B2(n10040), .ZN(
        P1_U3463) );
  AOI22_X1 U11117 ( .A1(n10012), .A2(n10011), .B1(n10010), .B2(n10009), .ZN(
        n10013) );
  OAI211_X1 U11118 ( .C1(n10016), .C2(n10015), .A(n10014), .B(n10013), .ZN(
        n10017) );
  INV_X1 U11119 ( .A(n10017), .ZN(n10050) );
  INV_X1 U11120 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n10018) );
  AOI22_X1 U11121 ( .A1(n10042), .A2(n10050), .B1(n10018), .B2(n10040), .ZN(
        P1_U3466) );
  OAI22_X1 U11122 ( .A1(n10020), .A2(n10034), .B1(n10019), .B2(n10032), .ZN(
        n10022) );
  AOI211_X1 U11123 ( .C1(n10039), .C2(n10023), .A(n10022), .B(n10021), .ZN(
        n10051) );
  INV_X1 U11124 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n10024) );
  AOI22_X1 U11125 ( .A1(n10042), .A2(n10051), .B1(n10024), .B2(n10040), .ZN(
        P1_U3472) );
  OAI21_X1 U11126 ( .B1(n10026), .B2(n10032), .A(n10025), .ZN(n10028) );
  AOI211_X1 U11127 ( .C1(n10030), .C2(n10029), .A(n10028), .B(n10027), .ZN(
        n10052) );
  INV_X1 U11128 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n10031) );
  AOI22_X1 U11129 ( .A1(n10042), .A2(n10052), .B1(n10031), .B2(n10040), .ZN(
        P1_U3475) );
  OAI22_X1 U11130 ( .A1(n10035), .A2(n10034), .B1(n10033), .B2(n10032), .ZN(
        n10037) );
  AOI211_X1 U11131 ( .C1(n10039), .C2(n10038), .A(n10037), .B(n10036), .ZN(
        n10055) );
  INV_X1 U11132 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n10041) );
  AOI22_X1 U11133 ( .A1(n10042), .A2(n10055), .B1(n10041), .B2(n10040), .ZN(
        P1_U3481) );
  AOI22_X1 U11134 ( .A1(n4392), .A2(n10044), .B1(n10043), .B2(n10053), .ZN(
        P1_U3524) );
  AOI22_X1 U11135 ( .A1(n4392), .A2(n10046), .B1(n10045), .B2(n10053), .ZN(
        P1_U3525) );
  INV_X1 U11136 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n10047) );
  AOI22_X1 U11137 ( .A1(n4392), .A2(n10048), .B1(n10047), .B2(n10053), .ZN(
        P1_U3526) );
  AOI22_X1 U11138 ( .A1(n4392), .A2(n10050), .B1(n10049), .B2(n10053), .ZN(
        P1_U3527) );
  AOI22_X1 U11139 ( .A1(n4392), .A2(n10051), .B1(n6856), .B2(n10053), .ZN(
        P1_U3529) );
  AOI22_X1 U11140 ( .A1(n4392), .A2(n10052), .B1(n7078), .B2(n10053), .ZN(
        P1_U3530) );
  INV_X1 U11141 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n10054) );
  AOI22_X1 U11142 ( .A1(n4392), .A2(n10055), .B1(n10054), .B2(n10053), .ZN(
        P1_U3532) );
  AOI22_X1 U11143 ( .A1(n10057), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n10056), .ZN(n10066) );
  AOI22_X1 U11144 ( .A1(n10058), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3152), .ZN(n10065) );
  OAI21_X1 U11145 ( .B1(n10060), .B2(P2_REG1_REG_0__SCAN_IN), .A(n10059), .ZN(
        n10063) );
  NOR2_X1 U11146 ( .A1(n10061), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n10062) );
  OAI21_X1 U11147 ( .B1(n10063), .B2(n10062), .A(P2_IR_REG_0__SCAN_IN), .ZN(
        n10064) );
  OAI211_X1 U11148 ( .C1(P2_IR_REG_0__SCAN_IN), .C2(n10066), .A(n10065), .B(
        n10064), .ZN(P2_U3245) );
  NOR2_X1 U11149 ( .A1(n10067), .A2(n10089), .ZN(n10076) );
  OAI21_X1 U11150 ( .B1(n10069), .B2(n10068), .A(n10077), .ZN(n10075) );
  OAI22_X1 U11151 ( .A1(n10073), .A2(n10072), .B1(n10071), .B2(n10070), .ZN(
        n10074) );
  AOI21_X1 U11152 ( .B1(n10076), .B2(n10075), .A(n10074), .ZN(n10159) );
  XNOR2_X1 U11153 ( .A(n10078), .B(n10077), .ZN(n10162) );
  XNOR2_X1 U11154 ( .A(n10079), .B(n10157), .ZN(n10158) );
  OAI22_X1 U11155 ( .A1(n10081), .A2(n6947), .B1(n10080), .B2(n10096), .ZN(
        n10082) );
  AOI21_X1 U11156 ( .B1(n10102), .B2(n10083), .A(n10082), .ZN(n10084) );
  OAI21_X1 U11157 ( .B1(n10158), .B2(n10085), .A(n10084), .ZN(n10086) );
  AOI21_X1 U11158 ( .B1(n10162), .B2(n10105), .A(n10086), .ZN(n10087) );
  OAI21_X1 U11159 ( .B1(n10108), .B2(n10159), .A(n10087), .ZN(P2_U3289) );
  INV_X1 U11160 ( .A(n10088), .ZN(n10090) );
  AOI21_X1 U11161 ( .B1(n10090), .B2(n10101), .A(n10089), .ZN(n10092) );
  AOI21_X1 U11162 ( .B1(n10092), .B2(n7241), .A(n10091), .ZN(n10146) );
  AOI21_X1 U11163 ( .B1(n10093), .B2(n10103), .A(n10194), .ZN(n10095) );
  NAND2_X1 U11164 ( .A1(n10095), .A2(n10094), .ZN(n10145) );
  OAI22_X1 U11165 ( .A1(n10098), .A2(n10145), .B1(n10097), .B2(n10096), .ZN(
        n10099) );
  INV_X1 U11166 ( .A(n10099), .ZN(n10107) );
  XNOR2_X1 U11167 ( .A(n10101), .B(n10100), .ZN(n10149) );
  AOI222_X1 U11168 ( .A1(n10149), .A2(n10105), .B1(P2_REG2_REG_4__SCAN_IN), 
        .B2(n10104), .C1(n10103), .C2(n10102), .ZN(n10106) );
  OAI211_X1 U11169 ( .C1(n10108), .C2(n10146), .A(n10107), .B(n10106), .ZN(
        P2_U3292) );
  NOR2_X1 U11170 ( .A1(n10110), .A2(n10109), .ZN(n10114) );
  NOR2_X1 U11171 ( .A1(n10114), .A2(n10111), .ZN(P2_U3297) );
  AND2_X1 U11172 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n10117), .ZN(P2_U3298) );
  AND2_X1 U11173 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n10117), .ZN(P2_U3299) );
  AND2_X1 U11174 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n10117), .ZN(P2_U3300) );
  AND2_X1 U11175 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n10117), .ZN(P2_U3301) );
  AND2_X1 U11176 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n10117), .ZN(P2_U3302) );
  AND2_X1 U11177 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n10117), .ZN(P2_U3303) );
  AND2_X1 U11178 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n10117), .ZN(P2_U3304) );
  AND2_X1 U11179 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n10117), .ZN(P2_U3305) );
  AND2_X1 U11180 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n10117), .ZN(P2_U3306) );
  AND2_X1 U11181 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n10117), .ZN(P2_U3307) );
  NOR2_X1 U11182 ( .A1(n10114), .A2(n10112), .ZN(P2_U3308) );
  AND2_X1 U11183 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n10117), .ZN(P2_U3309) );
  NOR2_X1 U11184 ( .A1(n10114), .A2(n10113), .ZN(P2_U3310) );
  AND2_X1 U11185 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n10117), .ZN(P2_U3311) );
  AND2_X1 U11186 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n10117), .ZN(P2_U3312) );
  AND2_X1 U11187 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n10117), .ZN(P2_U3313) );
  AND2_X1 U11188 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n10117), .ZN(P2_U3314) );
  AND2_X1 U11189 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n10117), .ZN(P2_U3315) );
  AND2_X1 U11190 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n10117), .ZN(P2_U3316) );
  AND2_X1 U11191 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n10117), .ZN(P2_U3317) );
  AND2_X1 U11192 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n10117), .ZN(P2_U3318) );
  AND2_X1 U11193 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n10117), .ZN(P2_U3319) );
  AND2_X1 U11194 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n10117), .ZN(P2_U3320) );
  AND2_X1 U11195 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n10117), .ZN(P2_U3321) );
  AND2_X1 U11196 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n10117), .ZN(P2_U3322) );
  AND2_X1 U11197 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n10117), .ZN(P2_U3323) );
  AND2_X1 U11198 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n10117), .ZN(P2_U3324) );
  AND2_X1 U11199 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n10117), .ZN(P2_U3325) );
  AND2_X1 U11200 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n10117), .ZN(P2_U3326) );
  AOI22_X1 U11201 ( .A1(n10116), .A2(n10119), .B1(n10115), .B2(n10117), .ZN(
        P2_U3437) );
  AOI22_X1 U11202 ( .A1(n10120), .A2(n10119), .B1(n10118), .B2(n10117), .ZN(
        P2_U3438) );
  OAI21_X1 U11203 ( .B1(n10123), .B2(n10122), .A(n10121), .ZN(n10124) );
  AOI21_X1 U11204 ( .B1(n10125), .B2(n10199), .A(n10124), .ZN(n10204) );
  AOI22_X1 U11205 ( .A1(n10202), .A2(n10204), .B1(n5967), .B2(n10200), .ZN(
        P2_U3451) );
  AOI22_X1 U11206 ( .A1(n10128), .A2(n4942), .B1(n10127), .B2(n10126), .ZN(
        n10129) );
  OAI21_X1 U11207 ( .B1(n10131), .B2(n10130), .A(n10129), .ZN(n10133) );
  NOR2_X1 U11208 ( .A1(n10133), .A2(n10132), .ZN(n10205) );
  AOI22_X1 U11209 ( .A1(n10202), .A2(n10205), .B1(n5977), .B2(n10200), .ZN(
        P2_U3454) );
  INV_X1 U11210 ( .A(n10134), .ZN(n10135) );
  OAI21_X1 U11211 ( .B1(n10136), .B2(n10192), .A(n10135), .ZN(n10137) );
  AOI211_X1 U11212 ( .C1(n10199), .C2(n10139), .A(n10138), .B(n10137), .ZN(
        n10206) );
  AOI22_X1 U11213 ( .A1(n10202), .A2(n10206), .B1(n5993), .B2(n10200), .ZN(
        P2_U3457) );
  OAI21_X1 U11214 ( .B1(n10141), .B2(n10192), .A(n10140), .ZN(n10143) );
  AOI211_X1 U11215 ( .C1(n10199), .C2(n10144), .A(n10143), .B(n10142), .ZN(
        n10208) );
  AOI22_X1 U11216 ( .A1(n10202), .A2(n10208), .B1(n5944), .B2(n10200), .ZN(
        P2_U3460) );
  OAI211_X1 U11217 ( .C1(n10147), .C2(n10192), .A(n10146), .B(n10145), .ZN(
        n10148) );
  AOI21_X1 U11218 ( .B1(n10199), .B2(n10149), .A(n10148), .ZN(n10209) );
  INV_X1 U11219 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n10150) );
  AOI22_X1 U11220 ( .A1(n10202), .A2(n10209), .B1(n10150), .B2(n10200), .ZN(
        P2_U3463) );
  OAI22_X1 U11221 ( .A1(n10152), .A2(n10194), .B1(n10151), .B2(n10192), .ZN(
        n10154) );
  AOI211_X1 U11222 ( .C1(n10199), .C2(n10155), .A(n10154), .B(n10153), .ZN(
        n10210) );
  INV_X1 U11223 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10156) );
  AOI22_X1 U11224 ( .A1(n10202), .A2(n10210), .B1(n10156), .B2(n10200), .ZN(
        P2_U3469) );
  OAI22_X1 U11225 ( .A1(n10158), .A2(n10194), .B1(n10157), .B2(n10192), .ZN(
        n10161) );
  INV_X1 U11226 ( .A(n10159), .ZN(n10160) );
  AOI211_X1 U11227 ( .C1(n10199), .C2(n10162), .A(n10161), .B(n10160), .ZN(
        n10211) );
  INV_X1 U11228 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n10163) );
  AOI22_X1 U11229 ( .A1(n10202), .A2(n10211), .B1(n10163), .B2(n10200), .ZN(
        P2_U3472) );
  INV_X1 U11230 ( .A(n10164), .ZN(n10169) );
  OAI22_X1 U11231 ( .A1(n10166), .A2(n10194), .B1(n10165), .B2(n10192), .ZN(
        n10168) );
  AOI211_X1 U11232 ( .C1(n10184), .C2(n10169), .A(n10168), .B(n10167), .ZN(
        n10213) );
  AOI22_X1 U11233 ( .A1(n10202), .A2(n10213), .B1(n5903), .B2(n10200), .ZN(
        P2_U3475) );
  INV_X1 U11234 ( .A(n10170), .ZN(n10175) );
  OAI22_X1 U11235 ( .A1(n10172), .A2(n10194), .B1(n10171), .B2(n10192), .ZN(
        n10174) );
  AOI211_X1 U11236 ( .C1(n10184), .C2(n10175), .A(n10174), .B(n10173), .ZN(
        n10214) );
  INV_X1 U11237 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n10176) );
  AOI22_X1 U11238 ( .A1(n10202), .A2(n10214), .B1(n10176), .B2(n10200), .ZN(
        P2_U3478) );
  INV_X1 U11239 ( .A(n10177), .ZN(n10183) );
  INV_X1 U11240 ( .A(n10178), .ZN(n10179) );
  OAI22_X1 U11241 ( .A1(n10180), .A2(n10194), .B1(n10179), .B2(n10192), .ZN(
        n10182) );
  AOI211_X1 U11242 ( .C1(n10184), .C2(n10183), .A(n10182), .B(n10181), .ZN(
        n10215) );
  INV_X1 U11243 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n10185) );
  AOI22_X1 U11244 ( .A1(n10202), .A2(n10215), .B1(n10185), .B2(n10200), .ZN(
        P2_U3481) );
  OAI211_X1 U11245 ( .C1(n10188), .C2(n10192), .A(n10187), .B(n10186), .ZN(
        n10189) );
  AOI21_X1 U11246 ( .B1(n10190), .B2(n10199), .A(n10189), .ZN(n10216) );
  AOI22_X1 U11247 ( .A1(n10202), .A2(n10216), .B1(n10191), .B2(n10200), .ZN(
        P2_U3484) );
  OAI22_X1 U11248 ( .A1(n10195), .A2(n10194), .B1(n10193), .B2(n10192), .ZN(
        n10197) );
  AOI211_X1 U11249 ( .C1(n10199), .C2(n10198), .A(n10197), .B(n10196), .ZN(
        n10218) );
  AOI22_X1 U11250 ( .A1(n10202), .A2(n10218), .B1(n10201), .B2(n10200), .ZN(
        P2_U3487) );
  INV_X1 U11251 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n10203) );
  AOI22_X1 U11252 ( .A1(n10219), .A2(n10204), .B1(n10203), .B2(n10217), .ZN(
        P2_U3520) );
  AOI22_X1 U11253 ( .A1(n10219), .A2(n10205), .B1(n6931), .B2(n10217), .ZN(
        P2_U3521) );
  AOI22_X1 U11254 ( .A1(n10219), .A2(n10206), .B1(n6932), .B2(n10217), .ZN(
        P2_U3522) );
  INV_X1 U11255 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n10207) );
  AOI22_X1 U11256 ( .A1(n10219), .A2(n10208), .B1(n10207), .B2(n10217), .ZN(
        P2_U3523) );
  AOI22_X1 U11257 ( .A1(n10219), .A2(n10209), .B1(n6934), .B2(n10217), .ZN(
        P2_U3524) );
  AOI22_X1 U11258 ( .A1(n10219), .A2(n10210), .B1(n5955), .B2(n10217), .ZN(
        P2_U3526) );
  AOI22_X1 U11259 ( .A1(n10219), .A2(n10211), .B1(n6027), .B2(n10217), .ZN(
        P2_U3527) );
  INV_X1 U11260 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n10212) );
  AOI22_X1 U11261 ( .A1(n10219), .A2(n10213), .B1(n10212), .B2(n10217), .ZN(
        P2_U3528) );
  AOI22_X1 U11262 ( .A1(n10219), .A2(n10214), .B1(n7018), .B2(n10217), .ZN(
        P2_U3529) );
  AOI22_X1 U11263 ( .A1(n10219), .A2(n10215), .B1(n7136), .B2(n10217), .ZN(
        P2_U3530) );
  AOI22_X1 U11264 ( .A1(n10219), .A2(n10216), .B1(n7182), .B2(n10217), .ZN(
        P2_U3531) );
  AOI22_X1 U11265 ( .A1(n10219), .A2(n10218), .B1(n7340), .B2(n10217), .ZN(
        P2_U3532) );
  INV_X1 U11266 ( .A(n10220), .ZN(n10221) );
  NAND2_X1 U11267 ( .A1(n10222), .A2(n10221), .ZN(n10223) );
  XNOR2_X1 U11268 ( .A(P2_ADDR_REG_1__SCAN_IN), .B(n10223), .ZN(ADD_1071_U5)
         );
  AOI22_X1 U11269 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .B1(n10224), .B2(n7010), .ZN(ADD_1071_U46) );
  OAI21_X1 U11270 ( .B1(n10227), .B2(n10226), .A(n10225), .ZN(ADD_1071_U56) );
  OAI21_X1 U11271 ( .B1(n10230), .B2(n10229), .A(n10228), .ZN(ADD_1071_U57) );
  OAI21_X1 U11272 ( .B1(n10233), .B2(n10232), .A(n10231), .ZN(ADD_1071_U58) );
  OAI21_X1 U11273 ( .B1(n10236), .B2(n10235), .A(n10234), .ZN(ADD_1071_U59) );
  OAI21_X1 U11274 ( .B1(n10239), .B2(n10238), .A(n10237), .ZN(ADD_1071_U60) );
  OAI21_X1 U11275 ( .B1(n10242), .B2(n10241), .A(n10240), .ZN(ADD_1071_U61) );
  AOI21_X1 U11276 ( .B1(n10245), .B2(n10244), .A(n10243), .ZN(ADD_1071_U62) );
  AOI21_X1 U11277 ( .B1(n10248), .B2(n10247), .A(n10246), .ZN(ADD_1071_U63) );
  XNOR2_X1 U11278 ( .A(n10250), .B(n10249), .ZN(ADD_1071_U50) );
  NOR2_X1 U11279 ( .A1(n10252), .A2(n10251), .ZN(n10253) );
  XNOR2_X1 U11280 ( .A(n10253), .B(n7074), .ZN(ADD_1071_U51) );
  OAI21_X1 U11281 ( .B1(n10256), .B2(n10255), .A(n10254), .ZN(n10257) );
  XNOR2_X1 U11282 ( .A(n10257), .B(P1_ADDR_REG_18__SCAN_IN), .ZN(ADD_1071_U55)
         );
  AOI21_X1 U11283 ( .B1(n10260), .B2(n10259), .A(n10258), .ZN(ADD_1071_U47) );
  AOI21_X1 U11284 ( .B1(n10263), .B2(n10262), .A(n10261), .ZN(ADD_1071_U48) );
  XNOR2_X1 U11285 ( .A(n10265), .B(n10264), .ZN(ADD_1071_U49) );
  XOR2_X1 U11286 ( .A(n10267), .B(n10266), .Z(ADD_1071_U54) );
  XOR2_X1 U11287 ( .A(n10269), .B(n10268), .Z(ADD_1071_U53) );
  XNOR2_X1 U11288 ( .A(n10271), .B(n10270), .ZN(ADD_1071_U52) );
  CLKBUF_X1 U4910 ( .A(n5388), .Z(n7005) );
endmodule

