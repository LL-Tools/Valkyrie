

module b17_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, P1_MEMORYFETCH_REG_SCAN_IN, 
        DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, 
        DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, 
        DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, 
        DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, 
        DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, 
        DATAI_0_, HOLD, NA, BS16, READY1, READY2, P1_READREQUEST_REG_SCAN_IN, 
        P1_ADS_N_REG_SCAN_IN, P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, 
        P1_D_C_N_REG_SCAN_IN, P1_REQUESTPENDING_REG_SCAN_IN, 
        P1_STATEBS16_REG_SCAN_IN, P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, 
        P1_W_R_N_REG_SCAN_IN, P1_BYTEENABLE_REG_0__SCAN_IN, 
        P1_BYTEENABLE_REG_1__SCAN_IN, P1_BYTEENABLE_REG_2__SCAN_IN, 
        P1_BYTEENABLE_REG_3__SCAN_IN, P1_REIP_REG_31__SCAN_IN, 
        P1_REIP_REG_30__SCAN_IN, P1_REIP_REG_29__SCAN_IN, 
        P1_REIP_REG_28__SCAN_IN, P1_REIP_REG_27__SCAN_IN, 
        P1_REIP_REG_26__SCAN_IN, P1_REIP_REG_25__SCAN_IN, 
        P1_REIP_REG_24__SCAN_IN, P1_REIP_REG_23__SCAN_IN, 
        P1_REIP_REG_22__SCAN_IN, P1_REIP_REG_21__SCAN_IN, 
        P1_REIP_REG_20__SCAN_IN, P1_REIP_REG_19__SCAN_IN, 
        P1_REIP_REG_18__SCAN_IN, P1_REIP_REG_17__SCAN_IN, 
        P1_REIP_REG_16__SCAN_IN, P1_REIP_REG_15__SCAN_IN, 
        P1_REIP_REG_14__SCAN_IN, P1_REIP_REG_13__SCAN_IN, 
        P1_REIP_REG_12__SCAN_IN, P1_REIP_REG_11__SCAN_IN, 
        P1_REIP_REG_10__SCAN_IN, P1_REIP_REG_9__SCAN_IN, 
        P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN, 
        P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, P1_REIP_REG_3__SCAN_IN, 
        P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN, 
        P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, P1_EBX_REG_29__SCAN_IN, 
        P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN, 
        P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, P1_EBX_REG_23__SCAN_IN, 
        P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN, 
        P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, P1_EBX_REG_17__SCAN_IN, 
        P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN, 
        P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, P1_EBX_REG_11__SCAN_IN, 
        P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, P1_EBX_REG_8__SCAN_IN, 
        P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, P1_EBX_REG_5__SCAN_IN, 
        P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, P1_EBX_REG_2__SCAN_IN, 
        P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, P1_EAX_REG_31__SCAN_IN, 
        P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN, 
        P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, P1_EAX_REG_25__SCAN_IN, 
        P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN, 
        P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, P1_EAX_REG_19__SCAN_IN, 
        P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN, 
        P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, P1_EAX_REG_13__SCAN_IN, 
        P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, 
        P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, 
        P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, 
        P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, 
        P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, U355, 
        U356, U357, U358, U359, U360, U361, U362, U363, U364, U366, U367, U368, 
        U369, U370, U371, U372, U373, U374, U375, U347, U348, U349, U350, U351, 
        U352, U353, U354, U365, U376, U247, U246, U245, U244, U243, U242, U241, 
        U240, U239, U238, U237, U236, U235, U234, U233, U232, U231, U230, U229, 
        U228, U227, U226, U225, U224, U223, U222, U221, U220, U219, U218, U217, 
        U216, U251, U252, U253, U254, U255, U256, U257, U258, U259, U260, U261, 
        U262, U263, U264, U265, U266, U267, U268, U269, U270, U271, U272, U273, 
        U274, U275, U276, U277, U278, U279, U280, U281, U282, U212, U215, U213, 
        U214, P3_U3274, P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, 
        P3_U3059, P3_U3058, P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, 
        P3_U3052, P3_U3051, P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, 
        P3_U3045, P3_U3044, P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, 
        P3_U3038, P3_U3037, P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, 
        P3_U3031, P3_U3030, P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, 
        P3_U3026, P3_U3025, P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, 
        P3_U3019, P3_U3018, P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, 
        P3_U3012, P3_U3011, P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, 
        P3_U3005, P3_U3004, P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, 
        P3_U3282, P3_U2998, P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, 
        P3_U2992, P3_U2991, P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, 
        P3_U2985, P3_U2984, P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, 
        P3_U2978, P3_U2977, P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, 
        P3_U2971, P3_U2970, P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, 
        P3_U2964, P3_U2963, P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, 
        P3_U2957, P3_U2956, P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, 
        P3_U2950, P3_U2949, P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, 
        P3_U2943, P3_U2942, P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, 
        P3_U2936, P3_U2935, P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, 
        P3_U2929, P3_U2928, P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, 
        P3_U2922, P3_U2921, P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, 
        P3_U2915, P3_U2914, P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, 
        P3_U2908, P3_U2907, P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, 
        P3_U2901, P3_U2900, P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, 
        P3_U2894, P3_U2893, P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, 
        P3_U2887, P3_U2886, P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, 
        P3_U2880, P3_U2879, P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, 
        P3_U2873, P3_U2872, P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, 
        P3_U3285, P3_U3288, P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, 
        P3_U2864, P3_U2863, P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, 
        P3_U2857, P3_U2856, P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, 
        P3_U2850, P3_U2849, P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, 
        P3_U2843, P3_U2842, P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, 
        P3_U2836, P3_U2835, P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, 
        P3_U2829, P3_U2828, P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, 
        P3_U2822, P3_U2821, P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, 
        P3_U2815, P3_U2814, P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, 
        P3_U2808, P3_U2807, P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, 
        P3_U2801, P3_U2800, P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, 
        P3_U2794, P3_U2793, P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, 
        P3_U2787, P3_U2786, P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, 
        P3_U2780, P3_U2779, P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, 
        P3_U2773, P3_U2772, P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, 
        P3_U2766, P3_U2765, P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, 
        P3_U2759, P3_U2758, P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, 
        P3_U2752, P3_U2751, P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, 
        P3_U2745, P3_U2744, P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, 
        P3_U2738, P3_U2737, P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, 
        P3_U2731, P3_U2730, P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, 
        P3_U2724, P3_U2723, P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, 
        P3_U2717, P3_U2716, P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, 
        P3_U2710, P3_U2709, P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, 
        P3_U2703, P3_U2702, P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, 
        P3_U2696, P3_U2695, P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, 
        P3_U2689, P3_U2688, P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, 
        P3_U2682, P3_U2681, P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, 
        P3_U2675, P3_U2674, P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, 
        P3_U2668, P3_U2667, P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, 
        P3_U2661, P3_U2660, P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, 
        P3_U2654, P3_U2653, P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, 
        P3_U2647, P3_U2646, P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, 
        P3_U2640, P3_U2639, P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, 
        P3_U3295, P3_U2636, P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, 
        P3_U3298, P3_U3299, P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, 
        P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, 
        P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, 
        P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, 
        P2_U3179, P2_U3593, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, 
        P2_U3173, P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, 
        P2_U3166, P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, 
        P2_U3159, P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, 
        P2_U3152, P2_U3151, P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, 
        P2_U3145, P2_U3144, P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, 
        P2_U3138, P2_U3137, P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, 
        P2_U3131, P2_U3130, P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, 
        P2_U3124, P2_U3123, P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, 
        P2_U3117, P2_U3116, P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, 
        P2_U3110, P2_U3109, P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, 
        P2_U3103, P2_U3102, P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, 
        P2_U3096, P2_U3095, P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, 
        P2_U3089, P2_U3088, P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, 
        P2_U3082, P2_U3081, P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, 
        P2_U3075, P2_U3074, P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, 
        P2_U3068, P2_U3067, P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, 
        P2_U3061, P2_U3060, P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, 
        P2_U3054, P2_U3053, P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, 
        P2_U3595, P2_U3596, P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, 
        P2_U3603, P2_U3604, P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, 
        P2_U3042, P2_U3041, P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, 
        P2_U3035, P2_U3034, P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, 
        P2_U3028, P2_U3027, P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, 
        P2_U3021, P2_U3020, P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, 
        P2_U3014, P2_U3013, P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, 
        P2_U3007, P2_U3006, P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, 
        P2_U3000, P2_U2999, P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, 
        P2_U2993, P2_U2992, P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, 
        P2_U2986, P2_U2985, P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, 
        P2_U2979, P2_U2978, P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, 
        P2_U2972, P2_U2971, P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, 
        P2_U2965, P2_U2964, P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, 
        P2_U2958, P2_U2957, P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, 
        P2_U2951, P2_U2950, P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, 
        P2_U2944, P2_U2943, P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, 
        P2_U2937, P2_U2936, P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, 
        P2_U2930, P2_U2929, P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, 
        P2_U2923, P2_U2922, P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, 
        P2_U2916, P2_U2915, P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, 
        P2_U2909, P2_U2908, P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, 
        P2_U2902, P2_U2901, P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, 
        P2_U2895, P2_U2894, P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, 
        P2_U2888, P2_U2887, P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, 
        P2_U2881, P2_U2880, P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, 
        P2_U2874, P2_U2873, P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, 
        P2_U2867, P2_U2866, P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, 
        P2_U2860, P2_U2859, P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, 
        P2_U2853, P2_U2852, P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, 
        P2_U2846, P2_U2845, P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, 
        P2_U2839, P2_U2838, P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, 
        P2_U2832, P2_U2831, P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, 
        P2_U2825, P2_U2824, P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, 
        P2_U2819, P2_U3609, P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, 
        P2_U2815, P2_U3612, P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, 
        P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, 
        P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, 
        P1_U3212, P1_U3211, P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, 
        P1_U3205, P1_U3204, P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, 
        P1_U3198, P1_U3197, P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, 
        P1_U3193, P1_U3192, P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, 
        P1_U3186, P1_U3185, P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, 
        P1_U3179, P1_U3178, P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, 
        P1_U3172, P1_U3171, P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, 
        P1_U3165, P1_U3164, P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, 
        P1_U3159, P1_U3158, P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, 
        P1_U3152, P1_U3151, P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, 
        P1_U3145, P1_U3144, P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, 
        P1_U3138, P1_U3137, P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, 
        P1_U3131, P1_U3130, P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, 
        P1_U3124, P1_U3123, P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, 
        P1_U3117, P1_U3116, P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, 
        P1_U3110, P1_U3109, P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, 
        P1_U3103, P1_U3102, P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, 
        P1_U3096, P1_U3095, P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, 
        P1_U3089, P1_U3088, P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, 
        P1_U3082, P1_U3081, P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, 
        P1_U3075, P1_U3074, P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, 
        P1_U3068, P1_U3067, P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, 
        P1_U3061, P1_U3060, P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, 
        P1_U3054, P1_U3053, P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, 
        P1_U3047, P1_U3046, P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, 
        P1_U3040, P1_U3039, P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, 
        P1_U3033, P1_U3468, P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, 
        P1_U3475, P1_U3476, P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, 
        P1_U3028, P1_U3027, P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, 
        P1_U3021, P1_U3020, P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, 
        P1_U3014, P1_U3013, P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, 
        P1_U3007, P1_U3006, P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, 
        P1_U3000, P1_U2999, P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, 
        P1_U2993, P1_U2992, P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, 
        P1_U2986, P1_U2985, P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, 
        P1_U2979, P1_U2978, P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, 
        P1_U2972, P1_U2971, P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, 
        P1_U2965, P1_U2964, P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, 
        P1_U2958, P1_U2957, P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, 
        P1_U2951, P1_U2950, P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, 
        P1_U2944, P1_U2943, P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, 
        P1_U2937, P1_U2936, P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, 
        P1_U2930, P1_U2929, P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, 
        P1_U2923, P1_U2922, P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, 
        P1_U2916, P1_U2915, P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, 
        P1_U2909, P1_U2908, P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, 
        P1_U2902, P1_U2901, P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, 
        P1_U2895, P1_U2894, P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, 
        P1_U2888, P1_U2887, P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, 
        P1_U2881, P1_U2880, P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, 
        P1_U2874, P1_U2873, P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, 
        P1_U2867, P1_U2866, P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, 
        P1_U2860, P1_U2859, P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, 
        P1_U2853, P1_U2852, P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, 
        P1_U2846, P1_U2845, P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, 
        P1_U2839, P1_U2838, P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, 
        P1_U2832, P1_U2831, P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, 
        P1_U2825, P1_U2824, P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, 
        P1_U2818, P1_U2817, P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, 
        P1_U2811, P1_U2810, P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, 
        P1_U3483, P1_U2806, P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, 
        P1_U2803, P1_U2802, P1_U3487, P1_U2801 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_,
         DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_,
         DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_,
         DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_,
         DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_,
         DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_,
         HOLD, NA, BS16, READY1, READY2, P1_READREQUEST_REG_SCAN_IN,
         P1_ADS_N_REG_SCAN_IN, P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN,
         P1_D_C_N_REG_SCAN_IN, P1_REQUESTPENDING_REG_SCAN_IN,
         P1_STATEBS16_REG_SCAN_IN, P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN,
         P1_W_R_N_REG_SCAN_IN, P1_BYTEENABLE_REG_0__SCAN_IN,
         P1_BYTEENABLE_REG_1__SCAN_IN, P1_BYTEENABLE_REG_2__SCAN_IN,
         P1_BYTEENABLE_REG_3__SCAN_IN, P1_REIP_REG_31__SCAN_IN,
         P1_REIP_REG_30__SCAN_IN, P1_REIP_REG_29__SCAN_IN,
         P1_REIP_REG_28__SCAN_IN, P1_REIP_REG_27__SCAN_IN,
         P1_REIP_REG_26__SCAN_IN, P1_REIP_REG_25__SCAN_IN,
         P1_REIP_REG_24__SCAN_IN, P1_REIP_REG_23__SCAN_IN,
         P1_REIP_REG_22__SCAN_IN, P1_REIP_REG_21__SCAN_IN,
         P1_REIP_REG_20__SCAN_IN, P1_REIP_REG_19__SCAN_IN,
         P1_REIP_REG_18__SCAN_IN, P1_REIP_REG_17__SCAN_IN,
         P1_REIP_REG_16__SCAN_IN, P1_REIP_REG_15__SCAN_IN,
         P1_REIP_REG_14__SCAN_IN, P1_REIP_REG_13__SCAN_IN,
         P1_REIP_REG_12__SCAN_IN, P1_REIP_REG_11__SCAN_IN,
         P1_REIP_REG_10__SCAN_IN, P1_REIP_REG_9__SCAN_IN,
         P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN,
         P1_REIP_REG_6__SCAN_IN, P1_REIP_REG_5__SCAN_IN,
         P1_REIP_REG_4__SCAN_IN, P1_REIP_REG_3__SCAN_IN,
         P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN,
         P1_REIP_REG_0__SCAN_IN, P1_EBX_REG_31__SCAN_IN,
         P1_EBX_REG_30__SCAN_IN, P1_EBX_REG_29__SCAN_IN,
         P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN,
         P1_EBX_REG_26__SCAN_IN, P1_EBX_REG_25__SCAN_IN,
         P1_EBX_REG_24__SCAN_IN, P1_EBX_REG_23__SCAN_IN,
         P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN,
         P1_EBX_REG_20__SCAN_IN, P1_EBX_REG_19__SCAN_IN,
         P1_EBX_REG_18__SCAN_IN, P1_EBX_REG_17__SCAN_IN,
         P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN,
         P1_EBX_REG_14__SCAN_IN, P1_EBX_REG_13__SCAN_IN,
         P1_EBX_REG_12__SCAN_IN, P1_EBX_REG_11__SCAN_IN,
         P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, P1_EBX_REG_8__SCAN_IN,
         P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, P1_EBX_REG_5__SCAN_IN,
         P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, P1_EBX_REG_2__SCAN_IN,
         P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, P1_EAX_REG_31__SCAN_IN,
         P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN,
         P1_EAX_REG_28__SCAN_IN, P1_EAX_REG_27__SCAN_IN,
         P1_EAX_REG_26__SCAN_IN, P1_EAX_REG_25__SCAN_IN,
         P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN,
         P1_EAX_REG_22__SCAN_IN, P1_EAX_REG_21__SCAN_IN,
         P1_EAX_REG_20__SCAN_IN, P1_EAX_REG_19__SCAN_IN,
         P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN,
         P1_EAX_REG_16__SCAN_IN, P1_EAX_REG_15__SCAN_IN,
         P1_EAX_REG_14__SCAN_IN, P1_EAX_REG_13__SCAN_IN,
         P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN,
         P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN,
         P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN,
         P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN,
         P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n10949, n10950, n10951, n10952, n10953, n10954, n10955, n10956,
         n10957, n10958, n10959, n10960, n10961, n10962, n10963, n10964,
         n10965, n10966, n10967, n10968, n10970, n10971, n10972, n10973,
         n10974, n10975, n10976, n10977, n10978, n10979, n10980, n10981,
         n10982, n10983, n10984, n10985, n10986, n10987, n10988, n10989,
         n10990, n10991, n10992, n10993, n10994, n10995, n10996, n10997,
         n10998, n10999, n11000, n11001, n11002, n11003, n11004, n11005,
         n11006, n11007, n11008, n11009, n11010, n11011, n11012, n11013,
         n11014, n11015, n11016, n11017, n11018, n11019, n11020, n11021,
         n11022, n11023, n11024, n11025, n11026, n11027, n11028, n11029,
         n11030, n11031, n11032, n11033, n11034, n11035, n11036, n11037,
         n11038, n11039, n11040, n11041, n11042, n11043, n11044, n11045,
         n11046, n11047, n11048, n11049, n11050, n11051, n11052, n11053,
         n11054, n11055, n11056, n11057, n11058, n11059, n11060, n11061,
         n11062, n11063, n11064, n11065, n11066, n11067, n11068, n11069,
         n11070, n11071, n11072, n11073, n11074, n11075, n11076, n11077,
         n11078, n11079, n11080, n11081, n11082, n11083, n11084, n11085,
         n11086, n11087, n11088, n11089, n11090, n11091, n11092, n11093,
         n11094, n11095, n11096, n11097, n11098, n11099, n11100, n11101,
         n11102, n11103, n11104, n11105, n11106, n11107, n11108, n11109,
         n11110, n11111, n11112, n11113, n11114, n11115, n11116, n11117,
         n11118, n11119, n11120, n11121, n11122, n11123, n11124, n11125,
         n11126, n11127, n11128, n11129, n11130, n11131, n11132, n11133,
         n11134, n11135, n11136, n11137, n11138, n11139, n11140, n11141,
         n11142, n11143, n11144, n11145, n11146, n11147, n11148, n11149,
         n11150, n11151, n11152, n11153, n11154, n11155, n11156, n11157,
         n11158, n11159, n11160, n11161, n11162, n11163, n11164, n11165,
         n11166, n11167, n11168, n11169, n11170, n11171, n11172, n11173,
         n11174, n11175, n11176, n11177, n11178, n11179, n11180, n11181,
         n11182, n11183, n11184, n11185, n11186, n11187, n11188, n11189,
         n11190, n11191, n11192, n11193, n11194, n11195, n11196, n11197,
         n11198, n11199, n11200, n11201, n11202, n11203, n11204, n11205,
         n11206, n11207, n11208, n11209, n11210, n11211, n11212, n11213,
         n11214, n11215, n11216, n11217, n11218, n11219, n11220, n11221,
         n11222, n11223, n11224, n11225, n11226, n11227, n11228, n11229,
         n11230, n11231, n11232, n11233, n11234, n11235, n11236, n11237,
         n11238, n11239, n11240, n11241, n11242, n11243, n11244, n11245,
         n11246, n11247, n11248, n11249, n11250, n11251, n11252, n11253,
         n11254, n11255, n11256, n11257, n11258, n11259, n11260, n11261,
         n11262, n11263, n11264, n11265, n11266, n11267, n11268, n11269,
         n11270, n11271, n11272, n11273, n11274, n11275, n11276, n11277,
         n11278, n11279, n11280, n11281, n11282, n11283, n11284, n11285,
         n11286, n11287, n11288, n11289, n11290, n11291, n11292, n11293,
         n11294, n11295, n11296, n11297, n11298, n11299, n11300, n11301,
         n11302, n11303, n11304, n11305, n11306, n11307, n11308, n11309,
         n11310, n11311, n11312, n11313, n11314, n11315, n11316, n11317,
         n11318, n11319, n11320, n11321, n11322, n11323, n11324, n11325,
         n11326, n11327, n11328, n11329, n11330, n11331, n11332, n11333,
         n11334, n11335, n11336, n11337, n11338, n11339, n11340, n11341,
         n11342, n11343, n11344, n11345, n11346, n11347, n11348, n11349,
         n11350, n11351, n11352, n11353, n11354, n11355, n11356, n11357,
         n11358, n11359, n11360, n11361, n11362, n11363, n11364, n11365,
         n11366, n11367, n11368, n11369, n11370, n11371, n11372, n11373,
         n11374, n11375, n11376, n11377, n11378, n11379, n11380, n11381,
         n11382, n11383, n11384, n11385, n11386, n11387, n11388, n11389,
         n11390, n11391, n11392, n11393, n11394, n11395, n11396, n11397,
         n11398, n11399, n11400, n11401, n11402, n11403, n11404, n11405,
         n11406, n11407, n11408, n11409, n11410, n11411, n11412, n11413,
         n11414, n11415, n11416, n11417, n11418, n11419, n11420, n11421,
         n11422, n11423, n11424, n11425, n11426, n11427, n11428, n11429,
         n11430, n11431, n11432, n11433, n11434, n11435, n11436, n11437,
         n11438, n11439, n11440, n11441, n11442, n11443, n11444, n11445,
         n11446, n11447, n11448, n11449, n11450, n11451, n11452, n11453,
         n11454, n11455, n11456, n11457, n11458, n11459, n11460, n11461,
         n11462, n11463, n11464, n11465, n11466, n11467, n11468, n11469,
         n11470, n11471, n11472, n11473, n11474, n11475, n11476, n11477,
         n11478, n11479, n11480, n11481, n11482, n11483, n11484, n11485,
         n11486, n11487, n11488, n11489, n11490, n11491, n11492, n11493,
         n11494, n11495, n11496, n11497, n11498, n11499, n11500, n11501,
         n11502, n11503, n11504, n11505, n11506, n11507, n11508, n11509,
         n11510, n11511, n11512, n11513, n11514, n11515, n11516, n11517,
         n11518, n11519, n11520, n11521, n11522, n11523, n11524, n11525,
         n11526, n11527, n11528, n11529, n11530, n11531, n11532, n11533,
         n11534, n11535, n11536, n11537, n11538, n11539, n11540, n11541,
         n11542, n11543, n11544, n11545, n11546, n11547, n11548, n11549,
         n11550, n11551, n11552, n11553, n11554, n11555, n11556, n11557,
         n11558, n11559, n11560, n11561, n11562, n11563, n11564, n11565,
         n11566, n11567, n11568, n11569, n11570, n11571, n11572, n11573,
         n11574, n11575, n11576, n11577, n11578, n11579, n11580, n11581,
         n11582, n11583, n11584, n11585, n11586, n11587, n11588, n11589,
         n11590, n11591, n11592, n11593, n11594, n11595, n11596, n11597,
         n11598, n11599, n11600, n11601, n11602, n11603, n11604, n11605,
         n11606, n11607, n11608, n11609, n11610, n11611, n11612, n11613,
         n11614, n11615, n11616, n11617, n11618, n11619, n11620, n11621,
         n11622, n11623, n11624, n11625, n11626, n11627, n11628, n11629,
         n11630, n11631, n11632, n11633, n11634, n11635, n11636, n11637,
         n11638, n11639, n11640, n11641, n11642, n11643, n11644, n11645,
         n11646, n11647, n11648, n11649, n11650, n11651, n11652, n11653,
         n11654, n11655, n11656, n11657, n11658, n11659, n11660, n11661,
         n11662, n11663, n11664, n11665, n11666, n11667, n11668, n11669,
         n11670, n11671, n11672, n11673, n11674, n11675, n11676, n11677,
         n11678, n11679, n11680, n11681, n11682, n11683, n11684, n11685,
         n11686, n11687, n11688, n11689, n11690, n11691, n11692, n11693,
         n11694, n11695, n11696, n11697, n11698, n11699, n11700, n11701,
         n11702, n11703, n11704, n11705, n11706, n11707, n11708, n11709,
         n11710, n11711, n11712, n11713, n11714, n11715, n11716, n11717,
         n11718, n11719, n11720, n11721, n11722, n11723, n11724, n11725,
         n11726, n11727, n11728, n11729, n11730, n11731, n11732, n11733,
         n11734, n11735, n11736, n11737, n11738, n11739, n11740, n11741,
         n11742, n11743, n11744, n11745, n11746, n11747, n11748, n11749,
         n11750, n11751, n11752, n11753, n11754, n11755, n11756, n11757,
         n11758, n11759, n11760, n11761, n11762, n11763, n11764, n11765,
         n11766, n11767, n11768, n11769, n11770, n11771, n11772, n11773,
         n11774, n11775, n11776, n11777, n11778, n11779, n11780, n11781,
         n11782, n11783, n11784, n11785, n11786, n11787, n11788, n11789,
         n11790, n11791, n11792, n11793, n11794, n11795, n11796, n11797,
         n11798, n11799, n11800, n11801, n11802, n11803, n11804, n11805,
         n11806, n11807, n11808, n11809, n11810, n11811, n11812, n11813,
         n11814, n11815, n11816, n11817, n11818, n11819, n11820, n11821,
         n11822, n11823, n11824, n11825, n11826, n11827, n11828, n11829,
         n11830, n11831, n11832, n11833, n11834, n11835, n11836, n11837,
         n11838, n11839, n11840, n11841, n11842, n11843, n11844, n11845,
         n11846, n11847, n11848, n11849, n11850, n11851, n11852, n11853,
         n11854, n11855, n11856, n11857, n11858, n11859, n11860, n11861,
         n11862, n11863, n11864, n11865, n11866, n11867, n11868, n11869,
         n11870, n11871, n11872, n11873, n11874, n11875, n11876, n11877,
         n11878, n11879, n11880, n11881, n11882, n11883, n11884, n11885,
         n11886, n11887, n11888, n11889, n11890, n11891, n11892, n11893,
         n11894, n11895, n11896, n11897, n11898, n11899, n11900, n11901,
         n11902, n11903, n11904, n11905, n11906, n11907, n11908, n11909,
         n11910, n11911, n11912, n11913, n11914, n11915, n11916, n11917,
         n11918, n11919, n11920, n11921, n11922, n11923, n11924, n11925,
         n11926, n11927, n11928, n11929, n11930, n11931, n11932, n11933,
         n11934, n11935, n11936, n11937, n11938, n11939, n11940, n11941,
         n11942, n11943, n11944, n11945, n11946, n11947, n11948, n11949,
         n11950, n11951, n11952, n11953, n11954, n11955, n11956, n11957,
         n11958, n11959, n11960, n11961, n11962, n11963, n11964, n11965,
         n11966, n11967, n11968, n11969, n11970, n11971, n11972, n11973,
         n11974, n11975, n11976, n11977, n11978, n11979, n11980, n11981,
         n11982, n11983, n11984, n11985, n11986, n11987, n11988, n11989,
         n11990, n11991, n11992, n11993, n11994, n11995, n11996, n11997,
         n11998, n11999, n12000, n12001, n12002, n12003, n12004, n12005,
         n12006, n12007, n12008, n12009, n12010, n12011, n12012, n12013,
         n12014, n12015, n12016, n12017, n12018, n12019, n12020, n12021,
         n12022, n12023, n12024, n12025, n12026, n12027, n12028, n12029,
         n12030, n12031, n12032, n12033, n12034, n12035, n12036, n12037,
         n12038, n12039, n12040, n12041, n12042, n12043, n12044, n12045,
         n12046, n12047, n12048, n12049, n12050, n12051, n12052, n12053,
         n12054, n12055, n12056, n12057, n12058, n12059, n12060, n12061,
         n12062, n12063, n12064, n12065, n12066, n12067, n12068, n12069,
         n12070, n12071, n12072, n12073, n12074, n12075, n12076, n12077,
         n12078, n12079, n12080, n12081, n12082, n12083, n12084, n12085,
         n12086, n12087, n12088, n12089, n12090, n12091, n12092, n12093,
         n12094, n12095, n12096, n12097, n12098, n12099, n12100, n12101,
         n12102, n12103, n12104, n12105, n12106, n12107, n12108, n12109,
         n12110, n12111, n12112, n12113, n12114, n12115, n12116, n12117,
         n12118, n12119, n12120, n12121, n12122, n12123, n12124, n12125,
         n12126, n12127, n12128, n12129, n12130, n12131, n12132, n12133,
         n12134, n12135, n12136, n12137, n12138, n12139, n12140, n12141,
         n12142, n12143, n12144, n12145, n12146, n12147, n12148, n12149,
         n12150, n12151, n12152, n12153, n12154, n12155, n12156, n12157,
         n12158, n12159, n12160, n12161, n12162, n12163, n12164, n12165,
         n12166, n12167, n12168, n12169, n12170, n12171, n12172, n12173,
         n12174, n12175, n12176, n12177, n12178, n12179, n12180, n12181,
         n12182, n12183, n12184, n12185, n12186, n12187, n12188, n12189,
         n12190, n12191, n12192, n12193, n12194, n12195, n12196, n12197,
         n12198, n12199, n12200, n12201, n12202, n12203, n12204, n12205,
         n12206, n12207, n12208, n12209, n12210, n12211, n12212, n12213,
         n12214, n12215, n12216, n12217, n12218, n12219, n12220, n12221,
         n12222, n12223, n12224, n12225, n12226, n12227, n12228, n12229,
         n12230, n12231, n12232, n12233, n12234, n12235, n12236, n12237,
         n12238, n12239, n12240, n12241, n12242, n12243, n12244, n12245,
         n12246, n12247, n12248, n12249, n12250, n12251, n12252, n12253,
         n12254, n12255, n12256, n12257, n12258, n12259, n12260, n12261,
         n12262, n12263, n12264, n12265, n12266, n12267, n12268, n12269,
         n12270, n12271, n12273, n12274, n12275, n12276, n12277, n12278,
         n12279, n12280, n12281, n12282, n12283, n12284, n12285, n12286,
         n12287, n12288, n12289, n12290, n12291, n12292, n12293, n12294,
         n12295, n12296, n12297, n12298, n12299, n12300, n12301, n12302,
         n12303, n12304, n12305, n12306, n12307, n12308, n12309, n12310,
         n12311, n12312, n12313, n12314, n12315, n12316, n12317, n12318,
         n12319, n12320, n12321, n12322, n12323, n12324, n12325, n12326,
         n12327, n12328, n12329, n12330, n12331, n12332, n12333, n12334,
         n12335, n12336, n12337, n12338, n12339, n12340, n12341, n12342,
         n12343, n12344, n12345, n12346, n12347, n12348, n12349, n12350,
         n12351, n12352, n12353, n12354, n12355, n12356, n12357, n12358,
         n12359, n12360, n12361, n12362, n12363, n12364, n12365, n12366,
         n12367, n12368, n12369, n12370, n12371, n12372, n12373, n12374,
         n12375, n12376, n12377, n12378, n12379, n12380, n12381, n12382,
         n12383, n12384, n12385, n12386, n12387, n12388, n12389, n12390,
         n12391, n12392, n12393, n12394, n12395, n12396, n12397, n12398,
         n12399, n12400, n12401, n12402, n12403, n12404, n12405, n12406,
         n12407, n12408, n12409, n12410, n12411, n12412, n12413, n12414,
         n12415, n12416, n12417, n12418, n12419, n12420, n12421, n12422,
         n12423, n12424, n12425, n12426, n12427, n12428, n12429, n12430,
         n12431, n12432, n12433, n12434, n12435, n12436, n12437, n12438,
         n12439, n12440, n12441, n12442, n12443, n12444, n12445, n12446,
         n12447, n12448, n12449, n12450, n12451, n12452, n12453, n12454,
         n12455, n12456, n12457, n12458, n12459, n12460, n12461, n12462,
         n12463, n12464, n12465, n12466, n12467, n12468, n12469, n12470,
         n12471, n12472, n12473, n12474, n12475, n12476, n12477, n12478,
         n12479, n12480, n12481, n12482, n12483, n12484, n12485, n12486,
         n12487, n12488, n12489, n12490, n12491, n12492, n12493, n12494,
         n12495, n12496, n12497, n12498, n12499, n12500, n12501, n12502,
         n12503, n12504, n12505, n12506, n12507, n12508, n12509, n12510,
         n12511, n12512, n12513, n12514, n12515, n12516, n12517, n12518,
         n12519, n12520, n12521, n12522, n12523, n12524, n12525, n12526,
         n12527, n12528, n12529, n12530, n12531, n12532, n12533, n12534,
         n12535, n12536, n12537, n12538, n12539, n12540, n12541, n12542,
         n12543, n12544, n12545, n12546, n12547, n12548, n12549, n12550,
         n12551, n12552, n12553, n12554, n12555, n12556, n12557, n12558,
         n12559, n12560, n12561, n12562, n12563, n12564, n12565, n12566,
         n12567, n12568, n12569, n12570, n12571, n12572, n12573, n12574,
         n12575, n12576, n12577, n12578, n12579, n12580, n12581, n12582,
         n12583, n12584, n12585, n12586, n12587, n12588, n12589, n12590,
         n12591, n12592, n12593, n12594, n12595, n12596, n12597, n12598,
         n12599, n12600, n12601, n12602, n12603, n12604, n12605, n12606,
         n12607, n12608, n12609, n12610, n12611, n12612, n12613, n12614,
         n12615, n12616, n12617, n12618, n12619, n12620, n12621, n12622,
         n12623, n12624, n12625, n12626, n12627, n12628, n12629, n12630,
         n12631, n12632, n12633, n12634, n12635, n12636, n12637, n12638,
         n12639, n12640, n12641, n12642, n12643, n12644, n12645, n12646,
         n12647, n12648, n12649, n12650, n12651, n12652, n12653, n12654,
         n12655, n12656, n12657, n12658, n12659, n12660, n12661, n12662,
         n12663, n12664, n12665, n12666, n12667, n12668, n12669, n12670,
         n12671, n12672, n12673, n12674, n12675, n12676, n12677, n12678,
         n12679, n12680, n12681, n12682, n12683, n12684, n12685, n12686,
         n12687, n12688, n12689, n12690, n12691, n12692, n12693, n12694,
         n12695, n12696, n12697, n12698, n12699, n12700, n12701, n12702,
         n12703, n12704, n12705, n12706, n12707, n12708, n12709, n12710,
         n12711, n12712, n12713, n12714, n12715, n12716, n12717, n12718,
         n12719, n12720, n12721, n12722, n12723, n12724, n12725, n12726,
         n12727, n12728, n12729, n12730, n12731, n12732, n12733, n12734,
         n12735, n12736, n12737, n12738, n12739, n12740, n12741, n12742,
         n12743, n12744, n12745, n12746, n12747, n12748, n12749, n12750,
         n12751, n12752, n12753, n12754, n12755, n12756, n12757, n12758,
         n12759, n12760, n12761, n12762, n12763, n12764, n12765, n12766,
         n12767, n12768, n12769, n12770, n12771, n12772, n12773, n12774,
         n12775, n12776, n12777, n12778, n12779, n12780, n12781, n12782,
         n12783, n12784, n12785, n12786, n12787, n12788, n12789, n12790,
         n12791, n12792, n12793, n12794, n12795, n12796, n12797, n12798,
         n12799, n12800, n12801, n12802, n12803, n12804, n12805, n12806,
         n12807, n12808, n12809, n12810, n12811, n12812, n12813, n12814,
         n12815, n12816, n12817, n12818, n12819, n12820, n12821, n12822,
         n12823, n12824, n12825, n12826, n12827, n12828, n12829, n12830,
         n12831, n12832, n12833, n12834, n12835, n12836, n12837, n12838,
         n12839, n12840, n12841, n12842, n12843, n12844, n12845, n12846,
         n12847, n12848, n12849, n12850, n12851, n12852, n12853, n12854,
         n12855, n12856, n12857, n12858, n12859, n12860, n12861, n12862,
         n12863, n12864, n12865, n12866, n12867, n12868, n12869, n12870,
         n12871, n12872, n12873, n12874, n12875, n12876, n12877, n12878,
         n12879, n12880, n12881, n12882, n12883, n12884, n12885, n12886,
         n12887, n12888, n12889, n12890, n12891, n12892, n12893, n12894,
         n12895, n12896, n12897, n12898, n12899, n12900, n12901, n12902,
         n12903, n12904, n12905, n12906, n12907, n12908, n12909, n12910,
         n12911, n12912, n12913, n12914, n12915, n12916, n12917, n12918,
         n12919, n12920, n12921, n12922, n12923, n12924, n12925, n12926,
         n12927, n12928, n12929, n12930, n12931, n12932, n12933, n12934,
         n12935, n12936, n12937, n12938, n12939, n12940, n12941, n12942,
         n12943, n12944, n12945, n12946, n12947, n12948, n12949, n12950,
         n12951, n12952, n12953, n12954, n12955, n12956, n12957, n12958,
         n12959, n12960, n12961, n12962, n12963, n12964, n12965, n12966,
         n12967, n12968, n12969, n12970, n12971, n12972, n12973, n12974,
         n12975, n12976, n12977, n12978, n12979, n12980, n12981, n12982,
         n12983, n12984, n12985, n12986, n12987, n12988, n12989, n12990,
         n12991, n12992, n12993, n12994, n12995, n12996, n12997, n12998,
         n12999, n13000, n13001, n13002, n13003, n13004, n13005, n13006,
         n13007, n13008, n13009, n13010, n13011, n13012, n13013, n13014,
         n13015, n13016, n13017, n13018, n13019, n13020, n13021, n13022,
         n13023, n13024, n13025, n13026, n13027, n13028, n13029, n13030,
         n13031, n13032, n13033, n13034, n13035, n13036, n13037, n13038,
         n13039, n13040, n13041, n13042, n13043, n13044, n13045, n13046,
         n13047, n13048, n13049, n13050, n13051, n13052, n13053, n13054,
         n13055, n13056, n13057, n13058, n13059, n13060, n13061, n13062,
         n13063, n13064, n13065, n13066, n13067, n13068, n13069, n13070,
         n13071, n13072, n13073, n13074, n13075, n13076, n13077, n13078,
         n13079, n13080, n13081, n13082, n13083, n13084, n13085, n13086,
         n13087, n13088, n13089, n13090, n13091, n13092, n13093, n13094,
         n13095, n13096, n13097, n13098, n13099, n13100, n13101, n13102,
         n13103, n13104, n13105, n13106, n13107, n13108, n13109, n13110,
         n13111, n13112, n13113, n13114, n13115, n13116, n13117, n13118,
         n13119, n13120, n13121, n13122, n13123, n13124, n13125, n13126,
         n13127, n13128, n13129, n13130, n13131, n13132, n13133, n13134,
         n13135, n13136, n13137, n13138, n13139, n13140, n13141, n13142,
         n13143, n13144, n13145, n13146, n13147, n13148, n13149, n13150,
         n13151, n13152, n13153, n13154, n13155, n13156, n13157, n13158,
         n13159, n13160, n13161, n13162, n13163, n13164, n13165, n13166,
         n13167, n13168, n13169, n13170, n13171, n13172, n13173, n13174,
         n13175, n13176, n13177, n13178, n13179, n13180, n13181, n13182,
         n13183, n13184, n13185, n13186, n13187, n13188, n13189, n13190,
         n13191, n13192, n13193, n13194, n13195, n13196, n13197, n13198,
         n13199, n13200, n13201, n13202, n13203, n13204, n13205, n13206,
         n13207, n13208, n13209, n13210, n13211, n13212, n13213, n13214,
         n13215, n13216, n13217, n13218, n13219, n13220, n13221, n13222,
         n13223, n13224, n13225, n13226, n13227, n13228, n13229, n13230,
         n13231, n13232, n13233, n13234, n13235, n13236, n13237, n13238,
         n13239, n13240, n13241, n13242, n13243, n13244, n13245, n13246,
         n13247, n13248, n13249, n13250, n13251, n13252, n13253, n13254,
         n13255, n13256, n13257, n13258, n13259, n13260, n13261, n13262,
         n13263, n13264, n13265, n13266, n13267, n13268, n13269, n13270,
         n13271, n13272, n13273, n13274, n13275, n13276, n13277, n13278,
         n13279, n13280, n13281, n13282, n13283, n13284, n13285, n13286,
         n13287, n13288, n13289, n13290, n13291, n13292, n13293, n13294,
         n13295, n13296, n13297, n13298, n13299, n13300, n13301, n13302,
         n13303, n13304, n13305, n13306, n13307, n13308, n13309, n13310,
         n13311, n13312, n13313, n13314, n13315, n13316, n13317, n13318,
         n13319, n13320, n13321, n13322, n13323, n13324, n13325, n13326,
         n13327, n13328, n13329, n13330, n13331, n13332, n13333, n13334,
         n13335, n13336, n13337, n13338, n13339, n13340, n13341, n13342,
         n13343, n13344, n13345, n13346, n13347, n13348, n13349, n13350,
         n13351, n13352, n13353, n13354, n13355, n13356, n13357, n13358,
         n13359, n13360, n13361, n13362, n13363, n13364, n13365, n13366,
         n13367, n13368, n13369, n13370, n13371, n13372, n13373, n13374,
         n13375, n13376, n13377, n13378, n13379, n13380, n13381, n13382,
         n13383, n13384, n13385, n13386, n13387, n13388, n13389, n13390,
         n13391, n13392, n13393, n13394, n13395, n13396, n13397, n13398,
         n13399, n13400, n13401, n13402, n13403, n13404, n13405, n13406,
         n13407, n13408, n13409, n13410, n13411, n13412, n13413, n13414,
         n13415, n13416, n13417, n13418, n13419, n13420, n13421, n13422,
         n13423, n13424, n13425, n13426, n13427, n13428, n13429, n13430,
         n13431, n13432, n13433, n13434, n13435, n13436, n13437, n13438,
         n13439, n13440, n13441, n13442, n13443, n13444, n13445, n13446,
         n13447, n13448, n13449, n13450, n13451, n13452, n13453, n13454,
         n13455, n13456, n13457, n13458, n13459, n13460, n13461, n13462,
         n13463, n13464, n13465, n13466, n13467, n13468, n13469, n13470,
         n13471, n13472, n13473, n13474, n13475, n13476, n13477, n13478,
         n13479, n13480, n13481, n13482, n13483, n13484, n13485, n13486,
         n13487, n13488, n13489, n13490, n13491, n13492, n13493, n13494,
         n13495, n13496, n13497, n13498, n13499, n13500, n13501, n13502,
         n13503, n13504, n13505, n13506, n13507, n13508, n13509, n13510,
         n13511, n13512, n13513, n13514, n13515, n13516, n13517, n13518,
         n13519, n13520, n13521, n13522, n13523, n13524, n13525, n13526,
         n13527, n13528, n13529, n13530, n13531, n13532, n13533, n13534,
         n13535, n13536, n13537, n13538, n13539, n13540, n13541, n13542,
         n13543, n13544, n13545, n13546, n13547, n13548, n13549, n13550,
         n13551, n13552, n13553, n13554, n13555, n13556, n13557, n13558,
         n13559, n13560, n13561, n13562, n13563, n13564, n13565, n13566,
         n13567, n13568, n13569, n13570, n13571, n13572, n13573, n13574,
         n13575, n13576, n13577, n13578, n13579, n13580, n13581, n13582,
         n13583, n13584, n13585, n13586, n13587, n13588, n13589, n13590,
         n13591, n13592, n13593, n13594, n13595, n13596, n13597, n13598,
         n13599, n13600, n13601, n13602, n13603, n13604, n13605, n13606,
         n13607, n13608, n13609, n13610, n13611, n13612, n13613, n13614,
         n13615, n13616, n13617, n13618, n13619, n13620, n13621, n13622,
         n13623, n13624, n13625, n13626, n13627, n13628, n13629, n13630,
         n13631, n13632, n13633, n13634, n13635, n13636, n13637, n13638,
         n13639, n13640, n13641, n13642, n13643, n13644, n13645, n13646,
         n13647, n13648, n13649, n13650, n13651, n13652, n13653, n13654,
         n13655, n13656, n13657, n13658, n13659, n13660, n13661, n13662,
         n13663, n13664, n13665, n13666, n13667, n13668, n13669, n13670,
         n13671, n13672, n13673, n13674, n13675, n13676, n13677, n13678,
         n13679, n13680, n13681, n13682, n13683, n13684, n13685, n13686,
         n13687, n13688, n13689, n13690, n13691, n13692, n13693, n13694,
         n13695, n13696, n13697, n13698, n13699, n13700, n13701, n13702,
         n13703, n13704, n13705, n13706, n13707, n13708, n13709, n13710,
         n13711, n13712, n13713, n13714, n13715, n13716, n13717, n13718,
         n13719, n13720, n13721, n13722, n13723, n13724, n13725, n13726,
         n13727, n13728, n13729, n13730, n13731, n13732, n13733, n13734,
         n13735, n13736, n13737, n13738, n13739, n13740, n13741, n13742,
         n13743, n13744, n13745, n13746, n13747, n13748, n13749, n13750,
         n13751, n13752, n13753, n13754, n13755, n13756, n13757, n13758,
         n13759, n13760, n13761, n13762, n13763, n13764, n13765, n13766,
         n13767, n13768, n13769, n13770, n13771, n13772, n13773, n13774,
         n13775, n13776, n13777, n13778, n13779, n13780, n13781, n13782,
         n13783, n13784, n13785, n13786, n13787, n13788, n13789, n13790,
         n13791, n13792, n13793, n13794, n13795, n13796, n13797, n13798,
         n13799, n13800, n13801, n13802, n13803, n13804, n13805, n13806,
         n13807, n13808, n13809, n13810, n13811, n13812, n13813, n13814,
         n13815, n13816, n13817, n13818, n13819, n13820, n13821, n13822,
         n13823, n13824, n13825, n13826, n13827, n13828, n13829, n13830,
         n13831, n13832, n13833, n13834, n13835, n13836, n13837, n13838,
         n13839, n13840, n13841, n13842, n13843, n13844, n13845, n13846,
         n13847, n13848, n13849, n13850, n13851, n13852, n13853, n13854,
         n13855, n13856, n13857, n13858, n13859, n13860, n13861, n13862,
         n13863, n13864, n13865, n13866, n13867, n13868, n13869, n13870,
         n13871, n13872, n13873, n13874, n13875, n13876, n13877, n13878,
         n13879, n13880, n13881, n13882, n13883, n13884, n13885, n13886,
         n13887, n13888, n13889, n13890, n13891, n13892, n13893, n13894,
         n13895, n13896, n13897, n13898, n13899, n13900, n13901, n13902,
         n13903, n13904, n13905, n13906, n13907, n13908, n13909, n13910,
         n13911, n13912, n13913, n13914, n13915, n13916, n13917, n13918,
         n13919, n13920, n13921, n13922, n13923, n13924, n13925, n13926,
         n13927, n13928, n13929, n13930, n13931, n13932, n13933, n13934,
         n13935, n13936, n13937, n13938, n13939, n13940, n13941, n13942,
         n13943, n13944, n13945, n13946, n13947, n13948, n13949, n13950,
         n13951, n13952, n13953, n13954, n13955, n13956, n13957, n13958,
         n13959, n13960, n13961, n13962, n13963, n13964, n13965, n13966,
         n13967, n13968, n13969, n13970, n13971, n13972, n13973, n13974,
         n13975, n13976, n13977, n13978, n13979, n13980, n13981, n13982,
         n13983, n13984, n13985, n13986, n13987, n13988, n13989, n13990,
         n13991, n13992, n13993, n13994, n13995, n13996, n13997, n13998,
         n13999, n14000, n14001, n14002, n14003, n14004, n14005, n14006,
         n14007, n14008, n14009, n14010, n14011, n14012, n14013, n14014,
         n14015, n14016, n14017, n14018, n14019, n14020, n14021, n14022,
         n14023, n14024, n14025, n14026, n14027, n14028, n14029, n14030,
         n14031, n14032, n14033, n14034, n14035, n14036, n14037, n14038,
         n14039, n14040, n14041, n14042, n14043, n14044, n14045, n14046,
         n14047, n14048, n14049, n14050, n14051, n14052, n14053, n14054,
         n14055, n14056, n14057, n14058, n14059, n14060, n14061, n14062,
         n14063, n14064, n14065, n14066, n14067, n14068, n14069, n14070,
         n14071, n14072, n14073, n14074, n14075, n14076, n14077, n14078,
         n14079, n14080, n14081, n14082, n14083, n14084, n14085, n14086,
         n14087, n14088, n14089, n14090, n14091, n14092, n14093, n14094,
         n14095, n14096, n14097, n14098, n14099, n14100, n14101, n14102,
         n14103, n14104, n14105, n14106, n14107, n14108, n14109, n14110,
         n14111, n14112, n14113, n14114, n14115, n14116, n14117, n14118,
         n14119, n14120, n14121, n14122, n14123, n14124, n14125, n14126,
         n14127, n14128, n14129, n14130, n14131, n14132, n14133, n14134,
         n14135, n14136, n14137, n14138, n14139, n14140, n14141, n14142,
         n14143, n14144, n14145, n14146, n14147, n14148, n14149, n14150,
         n14151, n14152, n14153, n14154, n14155, n14156, n14157, n14158,
         n14159, n14160, n14161, n14162, n14163, n14164, n14165, n14166,
         n14167, n14168, n14169, n14170, n14171, n14172, n14173, n14174,
         n14175, n14176, n14177, n14178, n14179, n14180, n14181, n14182,
         n14183, n14184, n14185, n14186, n14187, n14188, n14189, n14190,
         n14191, n14192, n14193, n14194, n14195, n14196, n14197, n14198,
         n14199, n14200, n14201, n14202, n14203, n14204, n14205, n14206,
         n14207, n14208, n14209, n14210, n14211, n14212, n14213, n14214,
         n14215, n14216, n14217, n14218, n14219, n14220, n14221, n14222,
         n14223, n14224, n14225, n14226, n14227, n14228, n14229, n14230,
         n14231, n14232, n14233, n14234, n14235, n14236, n14237, n14238,
         n14239, n14240, n14241, n14242, n14243, n14244, n14245, n14246,
         n14247, n14248, n14249, n14250, n14251, n14252, n14253, n14254,
         n14255, n14256, n14257, n14258, n14259, n14260, n14261, n14262,
         n14263, n14264, n14265, n14266, n14267, n14268, n14269, n14270,
         n14271, n14272, n14273, n14274, n14275, n14276, n14277, n14278,
         n14279, n14280, n14281, n14282, n14283, n14284, n14285, n14286,
         n14287, n14288, n14289, n14290, n14291, n14292, n14293, n14294,
         n14295, n14296, n14297, n14298, n14299, n14300, n14301, n14302,
         n14303, n14304, n14305, n14306, n14307, n14308, n14309, n14310,
         n14311, n14312, n14313, n14314, n14315, n14316, n14317, n14318,
         n14319, n14320, n14321, n14322, n14323, n14324, n14325, n14326,
         n14327, n14328, n14329, n14330, n14331, n14332, n14333, n14334,
         n14335, n14336, n14337, n14338, n14339, n14340, n14341, n14342,
         n14343, n14344, n14345, n14346, n14347, n14348, n14349, n14350,
         n14351, n14352, n14353, n14354, n14355, n14356, n14357, n14358,
         n14359, n14360, n14361, n14362, n14363, n14364, n14365, n14366,
         n14367, n14368, n14369, n14370, n14371, n14372, n14373, n14374,
         n14375, n14376, n14377, n14378, n14379, n14380, n14381, n14382,
         n14383, n14384, n14385, n14386, n14387, n14388, n14389, n14390,
         n14391, n14392, n14393, n14394, n14395, n14396, n14397, n14398,
         n14399, n14400, n14401, n14402, n14403, n14404, n14405, n14406,
         n14407, n14408, n14409, n14410, n14411, n14412, n14413, n14414,
         n14415, n14416, n14417, n14418, n14419, n14420, n14421, n14422,
         n14423, n14424, n14425, n14426, n14427, n14428, n14429, n14430,
         n14431, n14432, n14433, n14434, n14435, n14436, n14437, n14438,
         n14439, n14440, n14441, n14442, n14443, n14444, n14445, n14446,
         n14447, n14448, n14449, n14450, n14451, n14452, n14453, n14454,
         n14455, n14456, n14457, n14458, n14459, n14460, n14461, n14462,
         n14463, n14464, n14465, n14466, n14467, n14468, n14469, n14470,
         n14471, n14472, n14473, n14474, n14475, n14476, n14477, n14478,
         n14479, n14480, n14481, n14482, n14483, n14484, n14485, n14486,
         n14487, n14488, n14489, n14490, n14491, n14492, n14493, n14494,
         n14495, n14496, n14497, n14498, n14499, n14500, n14501, n14502,
         n14503, n14504, n14505, n14506, n14507, n14508, n14509, n14510,
         n14511, n14512, n14513, n14514, n14515, n14516, n14517, n14518,
         n14519, n14520, n14521, n14522, n14523, n14524, n14525, n14526,
         n14527, n14528, n14529, n14530, n14531, n14532, n14533, n14534,
         n14535, n14536, n14537, n14538, n14539, n14540, n14541, n14542,
         n14543, n14544, n14545, n14546, n14547, n14548, n14549, n14550,
         n14551, n14552, n14553, n14554, n14555, n14556, n14557, n14558,
         n14559, n14560, n14561, n14562, n14563, n14564, n14565, n14566,
         n14567, n14568, n14569, n14570, n14571, n14572, n14573, n14574,
         n14575, n14576, n14577, n14578, n14579, n14580, n14581, n14582,
         n14583, n14584, n14585, n14586, n14587, n14588, n14589, n14590,
         n14591, n14592, n14593, n14594, n14595, n14596, n14597, n14598,
         n14599, n14600, n14601, n14602, n14603, n14604, n14605, n14606,
         n14607, n14608, n14609, n14610, n14611, n14612, n14613, n14614,
         n14615, n14616, n14617, n14618, n14619, n14620, n14621, n14622,
         n14623, n14624, n14625, n14626, n14627, n14628, n14629, n14630,
         n14631, n14632, n14633, n14634, n14635, n14636, n14637, n14638,
         n14639, n14640, n14641, n14642, n14643, n14644, n14645, n14646,
         n14647, n14648, n14649, n14650, n14651, n14652, n14653, n14654,
         n14655, n14656, n14657, n14658, n14659, n14660, n14661, n14662,
         n14663, n14664, n14665, n14666, n14667, n14668, n14669, n14670,
         n14671, n14672, n14673, n14674, n14675, n14676, n14677, n14678,
         n14679, n14680, n14681, n14682, n14683, n14684, n14685, n14686,
         n14687, n14688, n14689, n14690, n14691, n14692, n14693, n14694,
         n14695, n14696, n14697, n14698, n14699, n14700, n14701, n14702,
         n14703, n14704, n14705, n14706, n14707, n14708, n14709, n14710,
         n14711, n14712, n14713, n14714, n14715, n14716, n14717, n14718,
         n14719, n14720, n14721, n14722, n14723, n14724, n14725, n14726,
         n14727, n14728, n14729, n14730, n14731, n14732, n14733, n14734,
         n14735, n14736, n14737, n14738, n14739, n14740, n14741, n14742,
         n14743, n14744, n14745, n14746, n14747, n14748, n14749, n14750,
         n14751, n14752, n14753, n14754, n14755, n14756, n14757, n14758,
         n14759, n14760, n14761, n14762, n14763, n14764, n14765, n14766,
         n14767, n14768, n14769, n14770, n14771, n14772, n14773, n14774,
         n14775, n14776, n14777, n14778, n14779, n14780, n14781, n14782,
         n14783, n14784, n14785, n14786, n14787, n14788, n14789, n14790,
         n14791, n14792, n14793, n14794, n14795, n14796, n14797, n14798,
         n14799, n14800, n14801, n14802, n14803, n14804, n14805, n14806,
         n14807, n14808, n14809, n14810, n14811, n14812, n14813, n14814,
         n14815, n14816, n14817, n14818, n14819, n14820, n14821, n14822,
         n14823, n14824, n14825, n14826, n14827, n14828, n14829, n14830,
         n14831, n14832, n14833, n14834, n14835, n14836, n14837, n14838,
         n14839, n14840, n14841, n14842, n14843, n14844, n14845, n14846,
         n14847, n14848, n14849, n14850, n14851, n14852, n14853, n14854,
         n14855, n14856, n14857, n14858, n14859, n14860, n14861, n14862,
         n14863, n14864, n14865, n14866, n14867, n14868, n14869, n14870,
         n14871, n14872, n14873, n14874, n14875, n14876, n14877, n14878,
         n14879, n14880, n14881, n14882, n14883, n14884, n14885, n14886,
         n14887, n14888, n14889, n14890, n14891, n14892, n14893, n14894,
         n14895, n14896, n14897, n14898, n14899, n14900, n14901, n14902,
         n14903, n14904, n14905, n14906, n14907, n14908, n14909, n14910,
         n14911, n14912, n14913, n14914, n14915, n14916, n14917, n14918,
         n14919, n14920, n14921, n14922, n14923, n14924, n14925, n14926,
         n14927, n14928, n14929, n14930, n14931, n14932, n14933, n14934,
         n14935, n14936, n14937, n14938, n14939, n14940, n14941, n14942,
         n14943, n14944, n14945, n14946, n14947, n14948, n14949, n14950,
         n14951, n14952, n14953, n14954, n14955, n14956, n14957, n14958,
         n14959, n14960, n14961, n14962, n14963, n14964, n14965, n14966,
         n14967, n14968, n14969, n14970, n14971, n14972, n14973, n14974,
         n14975, n14976, n14977, n14978, n14979, n14980, n14981, n14982,
         n14983, n14984, n14985, n14986, n14987, n14988, n14989, n14990,
         n14991, n14992, n14993, n14994, n14995, n14996, n14997, n14998,
         n14999, n15000, n15001, n15002, n15003, n15004, n15005, n15006,
         n15007, n15008, n15009, n15010, n15011, n15012, n15013, n15014,
         n15015, n15016, n15017, n15018, n15019, n15020, n15021, n15022,
         n15023, n15024, n15025, n15026, n15027, n15028, n15029, n15030,
         n15031, n15032, n15033, n15034, n15035, n15036, n15037, n15038,
         n15039, n15040, n15041, n15042, n15043, n15044, n15045, n15046,
         n15047, n15048, n15049, n15050, n15051, n15052, n15053, n15054,
         n15055, n15056, n15057, n15058, n15059, n15060, n15061, n15062,
         n15063, n15064, n15065, n15066, n15067, n15068, n15069, n15070,
         n15071, n15072, n15073, n15074, n15075, n15076, n15077, n15078,
         n15079, n15080, n15081, n15082, n15083, n15084, n15085, n15086,
         n15087, n15088, n15089, n15090, n15091, n15092, n15093, n15094,
         n15095, n15096, n15097, n15098, n15099, n15100, n15101, n15102,
         n15103, n15104, n15105, n15106, n15107, n15108, n15109, n15110,
         n15111, n15112, n15113, n15114, n15115, n15116, n15117, n15118,
         n15119, n15120, n15121, n15122, n15123, n15124, n15125, n15126,
         n15127, n15128, n15129, n15130, n15131, n15132, n15133, n15134,
         n15135, n15136, n15137, n15138, n15139, n15140, n15141, n15142,
         n15143, n15144, n15145, n15146, n15147, n15148, n15149, n15150,
         n15151, n15152, n15153, n15154, n15155, n15156, n15157, n15158,
         n15159, n15160, n15161, n15162, n15163, n15164, n15165, n15166,
         n15167, n15168, n15169, n15170, n15171, n15172, n15173, n15174,
         n15175, n15176, n15177, n15178, n15179, n15180, n15181, n15182,
         n15183, n15184, n15185, n15186, n15187, n15188, n15189, n15190,
         n15191, n15192, n15193, n15194, n15195, n15196, n15197, n15198,
         n15199, n15200, n15201, n15202, n15203, n15204, n15205, n15206,
         n15207, n15208, n15209, n15210, n15211, n15212, n15213, n15214,
         n15215, n15216, n15217, n15218, n15219, n15220, n15221, n15222,
         n15223, n15224, n15225, n15226, n15227, n15228, n15229, n15230,
         n15231, n15232, n15233, n15234, n15235, n15236, n15237, n15238,
         n15239, n15240, n15241, n15242, n15243, n15244, n15245, n15246,
         n15247, n15248, n15249, n15250, n15251, n15252, n15253, n15254,
         n15255, n15256, n15257, n15258, n15259, n15260, n15261, n15262,
         n15263, n15264, n15265, n15266, n15267, n15268, n15269, n15270,
         n15271, n15272, n15273, n15274, n15275, n15276, n15277, n15278,
         n15279, n15280, n15281, n15282, n15283, n15284, n15285, n15286,
         n15287, n15288, n15289, n15290, n15291, n15292, n15293, n15294,
         n15295, n15296, n15297, n15298, n15299, n15300, n15301, n15302,
         n15303, n15304, n15305, n15306, n15307, n15308, n15309, n15310,
         n15311, n15312, n15313, n15314, n15315, n15316, n15317, n15318,
         n15319, n15320, n15321, n15322, n15323, n15324, n15325, n15326,
         n15327, n15328, n15329, n15330, n15331, n15332, n15333, n15334,
         n15335, n15336, n15337, n15338, n15339, n15340, n15341, n15342,
         n15343, n15344, n15345, n15346, n15347, n15348, n15349, n15350,
         n15351, n15352, n15353, n15354, n15355, n15356, n15357, n15358,
         n15359, n15360, n15361, n15362, n15363, n15364, n15365, n15366,
         n15367, n15368, n15369, n15370, n15371, n15372, n15373, n15374,
         n15375, n15376, n15377, n15378, n15379, n15380, n15381, n15382,
         n15383, n15384, n15385, n15386, n15387, n15388, n15389, n15390,
         n15391, n15392, n15393, n15394, n15395, n15396, n15397, n15398,
         n15399, n15400, n15401, n15402, n15403, n15404, n15405, n15406,
         n15407, n15408, n15409, n15410, n15411, n15412, n15413, n15414,
         n15416, n15417, n15418, n15419, n15420, n15421, n15422, n15423,
         n15424, n15425, n15426, n15427, n15428, n15429, n15430, n15431,
         n15432, n15433, n15434, n15435, n15436, n15437, n15438, n15439,
         n15440, n15441, n15442, n15443, n15444, n15445, n15446, n15447,
         n15448, n15449, n15450, n15451, n15452, n15453, n15454, n15455,
         n15456, n15457, n15458, n15459, n15460, n15461, n15462, n15463,
         n15464, n15465, n15466, n15467, n15468, n15469, n15470, n15471,
         n15472, n15473, n15474, n15475, n15476, n15477, n15478, n15479,
         n15480, n15481, n15482, n15483, n15484, n15485, n15486, n15487,
         n15488, n15489, n15490, n15491, n15492, n15493, n15494, n15495,
         n15496, n15497, n15498, n15499, n15500, n15501, n15502, n15503,
         n15504, n15505, n15506, n15507, n15508, n15509, n15510, n15511,
         n15512, n15513, n15514, n15515, n15516, n15517, n15518, n15519,
         n15520, n15521, n15522, n15523, n15524, n15525, n15526, n15527,
         n15528, n15529, n15530, n15531, n15532, n15533, n15534, n15535,
         n15536, n15537, n15538, n15539, n15540, n15541, n15542, n15543,
         n15544, n15545, n15546, n15547, n15548, n15549, n15550, n15551,
         n15552, n15553, n15554, n15555, n15556, n15557, n15558, n15559,
         n15560, n15561, n15562, n15563, n15564, n15565, n15566, n15567,
         n15568, n15569, n15570, n15571, n15572, n15573, n15574, n15575,
         n15576, n15577, n15578, n15579, n15580, n15581, n15582, n15583,
         n15584, n15585, n15586, n15587, n15588, n15589, n15590, n15591,
         n15592, n15593, n15594, n15595, n15596, n15597, n15598, n15599,
         n15600, n15601, n15602, n15603, n15604, n15605, n15606, n15607,
         n15608, n15609, n15610, n15611, n15612, n15613, n15614, n15615,
         n15616, n15617, n15618, n15619, n15620, n15621, n15622, n15623,
         n15624, n15625, n15626, n15627, n15628, n15629, n15630, n15631,
         n15632, n15633, n15634, n15635, n15636, n15637, n15638, n15639,
         n15640, n15641, n15642, n15643, n15644, n15645, n15646, n15647,
         n15648, n15649, n15650, n15651, n15652, n15653, n15654, n15655,
         n15656, n15657, n15658, n15659, n15660, n15661, n15662, n15663,
         n15664, n15665, n15666, n15667, n15668, n15669, n15670, n15671,
         n15672, n15673, n15674, n15675, n15676, n15677, n15678, n15679,
         n15680, n15681, n15682, n15683, n15684, n15685, n15686, n15687,
         n15688, n15689, n15690, n15691, n15692, n15693, n15694, n15695,
         n15696, n15697, n15698, n15699, n15700, n15701, n15702, n15703,
         n15704, n15705, n15706, n15707, n15708, n15709, n15710, n15711,
         n15712, n15713, n15714, n15715, n15716, n15717, n15718, n15719,
         n15720, n15721, n15722, n15723, n15724, n15725, n15726, n15727,
         n15728, n15729, n15730, n15731, n15732, n15733, n15734, n15735,
         n15736, n15737, n15738, n15739, n15740, n15741, n15742, n15743,
         n15744, n15745, n15746, n15747, n15748, n15749, n15750, n15751,
         n15752, n15753, n15754, n15755, n15756, n15757, n15758, n15759,
         n15760, n15761, n15762, n15763, n15764, n15765, n15766, n15767,
         n15768, n15769, n15770, n15771, n15772, n15773, n15774, n15775,
         n15776, n15777, n15778, n15779, n15780, n15781, n15782, n15783,
         n15784, n15785, n15786, n15787, n15788, n15789, n15790, n15791,
         n15792, n15793, n15794, n15795, n15796, n15797, n15798, n15799,
         n15800, n15801, n15802, n15803, n15804, n15805, n15806, n15807,
         n15808, n15809, n15810, n15811, n15812, n15813, n15814, n15815,
         n15816, n15817, n15818, n15819, n15820, n15821, n15822, n15823,
         n15824, n15825, n15826, n15827, n15828, n15829, n15830, n15831,
         n15832, n15833, n15834, n15835, n15836, n15837, n15838, n15839,
         n15840, n15841, n15842, n15843, n15844, n15845, n15846, n15847,
         n15848, n15849, n15850, n15851, n15852, n15853, n15854, n15855,
         n15856, n15857, n15858, n15859, n15860, n15861, n15862, n15863,
         n15864, n15865, n15866, n15867, n15868, n15869, n15870, n15871,
         n15872, n15873, n15874, n15875, n15876, n15877, n15878, n15879,
         n15880, n15881, n15882, n15883, n15884, n15885, n15886, n15887,
         n15888, n15889, n15890, n15891, n15892, n15893, n15894, n15895,
         n15896, n15897, n15898, n15899, n15900, n15901, n15902, n15903,
         n15904, n15905, n15906, n15907, n15908, n15909, n15910, n15911,
         n15912, n15913, n15914, n15915, n15916, n15917, n15918, n15919,
         n15920, n15921, n15922, n15923, n15924, n15925, n15926, n15927,
         n15928, n15929, n15930, n15931, n15932, n15933, n15934, n15935,
         n15936, n15937, n15938, n15939, n15940, n15941, n15942, n15943,
         n15944, n15945, n15946, n15947, n15948, n15949, n15950, n15951,
         n15952, n15953, n15954, n15955, n15956, n15957, n15958, n15959,
         n15960, n15961, n15962, n15963, n15964, n15965, n15966, n15967,
         n15968, n15969, n15970, n15971, n15972, n15973, n15974, n15975,
         n15976, n15977, n15978, n15979, n15980, n15981, n15982, n15983,
         n15984, n15985, n15986, n15987, n15988, n15989, n15990, n15991,
         n15992, n15993, n15994, n15995, n15996, n15997, n15998, n15999,
         n16000, n16001, n16002, n16003, n16004, n16005, n16006, n16007,
         n16008, n16009, n16010, n16011, n16012, n16013, n16014, n16015,
         n16016, n16017, n16018, n16019, n16020, n16021, n16022, n16023,
         n16024, n16025, n16026, n16027, n16028, n16029, n16030, n16031,
         n16032, n16033, n16034, n16035, n16036, n16037, n16038, n16039,
         n16040, n16041, n16042, n16043, n16044, n16045, n16046, n16047,
         n16048, n16049, n16050, n16051, n16052, n16053, n16054, n16055,
         n16056, n16057, n16058, n16059, n16060, n16061, n16062, n16063,
         n16064, n16065, n16066, n16067, n16068, n16069, n16070, n16071,
         n16072, n16073, n16074, n16075, n16076, n16077, n16078, n16079,
         n16080, n16081, n16082, n16083, n16084, n16085, n16086, n16087,
         n16088, n16089, n16090, n16091, n16092, n16093, n16094, n16095,
         n16096, n16097, n16098, n16099, n16100, n16101, n16102, n16103,
         n16104, n16105, n16106, n16107, n16108, n16109, n16110, n16111,
         n16112, n16113, n16114, n16115, n16116, n16117, n16118, n16119,
         n16120, n16121, n16122, n16123, n16124, n16125, n16126, n16127,
         n16128, n16129, n16130, n16131, n16132, n16133, n16134, n16135,
         n16136, n16137, n16138, n16139, n16140, n16141, n16142, n16143,
         n16144, n16145, n16146, n16147, n16148, n16149, n16150, n16151,
         n16152, n16153, n16154, n16155, n16156, n16157, n16158, n16159,
         n16160, n16161, n16162, n16163, n16164, n16165, n16166, n16167,
         n16168, n16169, n16170, n16171, n16172, n16173, n16174, n16175,
         n16176, n16177, n16178, n16179, n16180, n16181, n16182, n16183,
         n16184, n16185, n16186, n16187, n16188, n16189, n16190, n16191,
         n16192, n16193, n16194, n16195, n16196, n16197, n16198, n16199,
         n16200, n16201, n16202, n16203, n16204, n16205, n16206, n16207,
         n16208, n16209, n16210, n16211, n16212, n16213, n16214, n16215,
         n16216, n16217, n16218, n16219, n16220, n16221, n16222, n16223,
         n16224, n16225, n16226, n16227, n16228, n16229, n16230, n16231,
         n16232, n16233, n16234, n16235, n16236, n16237, n16238, n16239,
         n16240, n16241, n16242, n16243, n16244, n16245, n16246, n16247,
         n16248, n16249, n16250, n16251, n16252, n16253, n16254, n16255,
         n16256, n16257, n16258, n16259, n16260, n16261, n16262, n16263,
         n16264, n16265, n16266, n16267, n16268, n16269, n16270, n16271,
         n16272, n16273, n16274, n16275, n16276, n16277, n16278, n16279,
         n16280, n16281, n16282, n16283, n16284, n16285, n16286, n16287,
         n16288, n16289, n16290, n16291, n16292, n16293, n16294, n16295,
         n16296, n16297, n16298, n16299, n16300, n16301, n16302, n16303,
         n16304, n16305, n16306, n16307, n16308, n16309, n16310, n16311,
         n16312, n16313, n16314, n16315, n16316, n16317, n16318, n16319,
         n16320, n16321, n16322, n16323, n16324, n16325, n16326, n16327,
         n16328, n16329, n16330, n16331, n16332, n16333, n16334, n16335,
         n16336, n16337, n16338, n16339, n16340, n16341, n16342, n16343,
         n16344, n16345, n16346, n16347, n16348, n16349, n16350, n16351,
         n16352, n16353, n16354, n16355, n16356, n16357, n16358, n16359,
         n16360, n16361, n16362, n16363, n16364, n16365, n16366, n16367,
         n16368, n16369, n16370, n16371, n16372, n16373, n16374, n16375,
         n16376, n16377, n16378, n16379, n16380, n16381, n16382, n16383,
         n16384, n16385, n16386, n16387, n16388, n16389, n16390, n16391,
         n16392, n16393, n16394, n16395, n16396, n16397, n16398, n16399,
         n16400, n16401, n16402, n16403, n16404, n16405, n16406, n16407,
         n16408, n16409, n16410, n16411, n16412, n16413, n16414, n16415,
         n16416, n16417, n16418, n16419, n16420, n16421, n16422, n16423,
         n16424, n16425, n16426, n16427, n16428, n16429, n16430, n16431,
         n16432, n16433, n16434, n16435, n16436, n16437, n16438, n16439,
         n16440, n16441, n16442, n16443, n16444, n16445, n16446, n16447,
         n16448, n16449, n16450, n16451, n16452, n16453, n16454, n16455,
         n16456, n16457, n16458, n16459, n16460, n16461, n16462, n16463,
         n16464, n16465, n16466, n16467, n16468, n16469, n16470, n16471,
         n16472, n16473, n16474, n16475, n16476, n16477, n16478, n16479,
         n16480, n16481, n16482, n16483, n16484, n16485, n16486, n16487,
         n16488, n16489, n16490, n16491, n16492, n16493, n16494, n16495,
         n16496, n16497, n16498, n16499, n16500, n16501, n16502, n16503,
         n16504, n16505, n16506, n16507, n16508, n16509, n16510, n16511,
         n16512, n16513, n16514, n16515, n16516, n16517, n16518, n16519,
         n16520, n16521, n16522, n16523, n16524, n16525, n16526, n16527,
         n16528, n16529, n16530, n16531, n16532, n16533, n16534, n16535,
         n16536, n16537, n16538, n16539, n16540, n16541, n16542, n16543,
         n16544, n16545, n16546, n16547, n16548, n16549, n16550, n16551,
         n16552, n16553, n16554, n16555, n16556, n16557, n16558, n16559,
         n16560, n16561, n16562, n16563, n16564, n16565, n16566, n16567,
         n16568, n16569, n16570, n16571, n16572, n16573, n16574, n16575,
         n16576, n16577, n16578, n16579, n16580, n16581, n16582, n16583,
         n16584, n16585, n16586, n16587, n16588, n16589, n16590, n16591,
         n16592, n16593, n16594, n16595, n16596, n16597, n16598, n16599,
         n16600, n16601, n16602, n16603, n16604, n16605, n16606, n16607,
         n16608, n16609, n16610, n16611, n16612, n16613, n16614, n16615,
         n16616, n16617, n16618, n16619, n16620, n16621, n16622, n16623,
         n16624, n16625, n16626, n16627, n16628, n16629, n16630, n16631,
         n16632, n16633, n16634, n16635, n16636, n16637, n16638, n16639,
         n16640, n16641, n16642, n16643, n16644, n16645, n16646, n16647,
         n16648, n16649, n16650, n16651, n16652, n16653, n16654, n16655,
         n16656, n16657, n16658, n16659, n16660, n16661, n16662, n16663,
         n16664, n16665, n16666, n16667, n16668, n16669, n16670, n16671,
         n16672, n16673, n16674, n16675, n16676, n16677, n16678, n16679,
         n16680, n16681, n16682, n16683, n16684, n16685, n16686, n16687,
         n16688, n16689, n16690, n16691, n16692, n16693, n16694, n16695,
         n16696, n16697, n16698, n16699, n16700, n16701, n16702, n16703,
         n16704, n16705, n16706, n16707, n16708, n16709, n16710, n16711,
         n16712, n16713, n16714, n16715, n16716, n16717, n16718, n16719,
         n16720, n16721, n16722, n16723, n16724, n16725, n16726, n16727,
         n16728, n16729, n16730, n16731, n16732, n16733, n16734, n16735,
         n16736, n16737, n16738, n16739, n16740, n16741, n16742, n16743,
         n16744, n16745, n16746, n16747, n16748, n16749, n16750, n16751,
         n16752, n16753, n16754, n16755, n16756, n16757, n16758, n16759,
         n16760, n16761, n16762, n16763, n16764, n16765, n16766, n16767,
         n16768, n16769, n16770, n16771, n16772, n16773, n16774, n16775,
         n16776, n16777, n16778, n16779, n16780, n16781, n16782, n16783,
         n16784, n16785, n16786, n16787, n16788, n16789, n16790, n16791,
         n16792, n16793, n16794, n16795, n16796, n16797, n16798, n16799,
         n16800, n16801, n16802, n16803, n16804, n16805, n16806, n16807,
         n16808, n16809, n16810, n16811, n16812, n16813, n16814, n16815,
         n16816, n16817, n16818, n16819, n16820, n16821, n16822, n16823,
         n16824, n16825, n16826, n16827, n16828, n16829, n16830, n16831,
         n16832, n16833, n16834, n16835, n16836, n16837, n16838, n16839,
         n16840, n16841, n16842, n16843, n16844, n16845, n16846, n16847,
         n16848, n16849, n16850, n16851, n16852, n16853, n16854, n16855,
         n16856, n16857, n16858, n16859, n16860, n16861, n16862, n16863,
         n16864, n16865, n16866, n16867, n16868, n16869, n16870, n16871,
         n16872, n16873, n16874, n16875, n16876, n16877, n16878, n16879,
         n16880, n16881, n16882, n16883, n16884, n16885, n16886, n16887,
         n16888, n16889, n16890, n16891, n16892, n16893, n16894, n16895,
         n16896, n16897, n16898, n16899, n16900, n16901, n16902, n16903,
         n16904, n16905, n16906, n16907, n16908, n16909, n16910, n16911,
         n16912, n16913, n16914, n16915, n16916, n16917, n16918, n16919,
         n16920, n16921, n16922, n16923, n16924, n16925, n16926, n16927,
         n16928, n16929, n16930, n16931, n16932, n16933, n16934, n16935,
         n16936, n16937, n16938, n16939, n16940, n16941, n16942, n16943,
         n16944, n16945, n16946, n16947, n16948, n16949, n16950, n16951,
         n16952, n16953, n16954, n16955, n16956, n16957, n16958, n16959,
         n16960, n16961, n16962, n16963, n16964, n16965, n16966, n16967,
         n16968, n16969, n16970, n16971, n16972, n16973, n16974, n16975,
         n16976, n16977, n16978, n16979, n16980, n16981, n16982, n16983,
         n16984, n16985, n16986, n16987, n16988, n16989, n16990, n16991,
         n16992, n16993, n16994, n16995, n16996, n16997, n16998, n16999,
         n17000, n17001, n17002, n17003, n17004, n17005, n17006, n17007,
         n17008, n17009, n17010, n17011, n17012, n17013, n17014, n17015,
         n17016, n17017, n17018, n17019, n17020, n17021, n17022, n17023,
         n17024, n17025, n17026, n17027, n17028, n17029, n17030, n17031,
         n17032, n17033, n17034, n17035, n17036, n17037, n17038, n17039,
         n17040, n17041, n17042, n17043, n17044, n17045, n17046, n17047,
         n17048, n17049, n17050, n17051, n17052, n17053, n17054, n17055,
         n17056, n17057, n17058, n17059, n17060, n17061, n17062, n17063,
         n17064, n17065, n17066, n17067, n17068, n17069, n17070, n17071,
         n17072, n17073, n17074, n17075, n17076, n17077, n17078, n17079,
         n17080, n17081, n17082, n17083, n17084, n17085, n17086, n17087,
         n17088, n17089, n17090, n17091, n17092, n17093, n17094, n17095,
         n17096, n17097, n17098, n17099, n17100, n17101, n17102, n17103,
         n17104, n17105, n17106, n17107, n17108, n17109, n17110, n17111,
         n17112, n17113, n17114, n17115, n17116, n17117, n17118, n17119,
         n17120, n17121, n17122, n17123, n17124, n17125, n17126, n17127,
         n17128, n17129, n17130, n17131, n17132, n17133, n17134, n17135,
         n17136, n17137, n17138, n17139, n17140, n17141, n17142, n17143,
         n17144, n17145, n17146, n17147, n17148, n17149, n17150, n17151,
         n17152, n17153, n17154, n17155, n17156, n17157, n17158, n17159,
         n17160, n17161, n17162, n17163, n17164, n17165, n17166, n17167,
         n17168, n17169, n17170, n17171, n17172, n17173, n17174, n17175,
         n17176, n17177, n17178, n17179, n17180, n17181, n17182, n17183,
         n17184, n17185, n17186, n17187, n17188, n17189, n17190, n17191,
         n17192, n17193, n17194, n17195, n17196, n17197, n17198, n17199,
         n17200, n17201, n17202, n17203, n17204, n17205, n17206, n17207,
         n17208, n17209, n17210, n17211, n17212, n17213, n17214, n17215,
         n17216, n17217, n17218, n17219, n17220, n17221, n17222, n17223,
         n17224, n17225, n17226, n17227, n17228, n17229, n17230, n17231,
         n17232, n17233, n17234, n17235, n17236, n17237, n17238, n17239,
         n17240, n17241, n17242, n17243, n17244, n17245, n17246, n17247,
         n17248, n17249, n17250, n17251, n17252, n17253, n17254, n17255,
         n17256, n17257, n17258, n17259, n17260, n17261, n17262, n17263,
         n17264, n17265, n17266, n17267, n17268, n17269, n17270, n17271,
         n17272, n17273, n17274, n17275, n17276, n17277, n17278, n17279,
         n17280, n17281, n17282, n17283, n17284, n17285, n17286, n17287,
         n17288, n17289, n17290, n17291, n17292, n17293, n17294, n17295,
         n17296, n17297, n17298, n17299, n17300, n17301, n17302, n17303,
         n17304, n17305, n17306, n17307, n17308, n17309, n17310, n17311,
         n17312, n17313, n17314, n17315, n17316, n17317, n17318, n17319,
         n17320, n17321, n17322, n17323, n17324, n17325, n17326, n17327,
         n17328, n17329, n17330, n17331, n17332, n17333, n17334, n17335,
         n17336, n17337, n17338, n17339, n17340, n17341, n17342, n17343,
         n17344, n17345, n17346, n17347, n17348, n17349, n17350, n17351,
         n17352, n17353, n17354, n17355, n17356, n17357, n17358, n17359,
         n17360, n17361, n17362, n17363, n17364, n17365, n17366, n17367,
         n17368, n17369, n17370, n17371, n17372, n17373, n17374, n17375,
         n17376, n17377, n17378, n17379, n17380, n17381, n17382, n17383,
         n17384, n17385, n17386, n17387, n17388, n17389, n17390, n17391,
         n17392, n17393, n17394, n17395, n17396, n17397, n17398, n17399,
         n17400, n17401, n17402, n17403, n17404, n17405, n17406, n17407,
         n17408, n17409, n17410, n17411, n17412, n17413, n17414, n17415,
         n17416, n17417, n17418, n17419, n17420, n17421, n17422, n17423,
         n17424, n17425, n17426, n17427, n17428, n17429, n17430, n17431,
         n17432, n17433, n17434, n17435, n17436, n17437, n17438, n17439,
         n17440, n17441, n17442, n17443, n17444, n17445, n17446, n17447,
         n17448, n17449, n17450, n17451, n17452, n17453, n17454, n17455,
         n17456, n17457, n17458, n17459, n17460, n17461, n17462, n17463,
         n17464, n17465, n17466, n17467, n17468, n17469, n17470, n17471,
         n17472, n17473, n17474, n17475, n17476, n17477, n17478, n17479,
         n17480, n17481, n17482, n17483, n17484, n17485, n17486, n17487,
         n17488, n17489, n17490, n17491, n17492, n17493, n17494, n17495,
         n17496, n17497, n17498, n17499, n17500, n17501, n17502, n17503,
         n17504, n17505, n17506, n17507, n17508, n17509, n17510, n17511,
         n17512, n17513, n17514, n17515, n17516, n17517, n17518, n17519,
         n17520, n17521, n17522, n17523, n17524, n17525, n17526, n17527,
         n17528, n17529, n17530, n17531, n17532, n17533, n17534, n17535,
         n17536, n17537, n17538, n17539, n17540, n17541, n17542, n17543,
         n17544, n17545, n17546, n17547, n17548, n17549, n17550, n17551,
         n17552, n17553, n17554, n17555, n17556, n17557, n17558, n17559,
         n17560, n17561, n17562, n17563, n17564, n17565, n17566, n17567,
         n17568, n17569, n17570, n17571, n17572, n17573, n17574, n17575,
         n17576, n17577, n17578, n17579, n17580, n17581, n17582, n17583,
         n17584, n17585, n17586, n17587, n17588, n17589, n17590, n17591,
         n17592, n17593, n17594, n17595, n17596, n17597, n17598, n17599,
         n17600, n17601, n17602, n17603, n17604, n17605, n17606, n17607,
         n17608, n17609, n17610, n17611, n17612, n17613, n17614, n17615,
         n17616, n17617, n17618, n17619, n17620, n17621, n17622, n17623,
         n17624, n17625, n17626, n17627, n17628, n17629, n17630, n17631,
         n17632, n17633, n17634, n17635, n17636, n17637, n17638, n17639,
         n17640, n17641, n17642, n17643, n17644, n17645, n17646, n17647,
         n17648, n17649, n17650, n17651, n17652, n17653, n17654, n17655,
         n17656, n17657, n17658, n17659, n17660, n17661, n17662, n17663,
         n17664, n17665, n17666, n17667, n17668, n17669, n17670, n17671,
         n17672, n17673, n17674, n17675, n17676, n17677, n17678, n17679,
         n17680, n17681, n17682, n17683, n17684, n17685, n17686, n17687,
         n17688, n17689, n17690, n17691, n17692, n17693, n17694, n17695,
         n17696, n17697, n17698, n17699, n17700, n17701, n17702, n17703,
         n17704, n17705, n17706, n17707, n17708, n17709, n17710, n17711,
         n17712, n17713, n17714, n17715, n17716, n17717, n17718, n17719,
         n17720, n17721, n17722, n17723, n17724, n17725, n17726, n17727,
         n17728, n17729, n17730, n17731, n17732, n17733, n17734, n17735,
         n17736, n17737, n17738, n17739, n17740, n17741, n17742, n17743,
         n17744, n17745, n17746, n17747, n17748, n17749, n17750, n17751,
         n17752, n17753, n17754, n17755, n17756, n17757, n17758, n17759,
         n17760, n17761, n17762, n17763, n17764, n17765, n17766, n17767,
         n17768, n17769, n17770, n17771, n17772, n17773, n17774, n17775,
         n17776, n17777, n17778, n17779, n17780, n17781, n17782, n17783,
         n17784, n17785, n17786, n17787, n17788, n17789, n17790, n17791,
         n17792, n17793, n17794, n17795, n17796, n17797, n17798, n17799,
         n17800, n17801, n17802, n17803, n17804, n17805, n17806, n17807,
         n17808, n17809, n17810, n17811, n17812, n17813, n17814, n17815,
         n17816, n17817, n17818, n17819, n17820, n17821, n17822, n17823,
         n17824, n17825, n17826, n17827, n17828, n17829, n17830, n17831,
         n17832, n17833, n17834, n17835, n17836, n17837, n17838, n17839,
         n17840, n17841, n17842, n17843, n17844, n17845, n17846, n17847,
         n17848, n17849, n17850, n17851, n17852, n17853, n17854, n17855,
         n17856, n17857, n17858, n17859, n17860, n17861, n17862, n17863,
         n17864, n17865, n17866, n17867, n17868, n17869, n17870, n17871,
         n17872, n17873, n17874, n17875, n17876, n17877, n17878, n17879,
         n17880, n17881, n17882, n17883, n17884, n17885, n17886, n17887,
         n17888, n17889, n17890, n17891, n17892, n17893, n17894, n17895,
         n17896, n17897, n17898, n17899, n17900, n17901, n17902, n17903,
         n17904, n17905, n17906, n17907, n17908, n17909, n17910, n17911,
         n17912, n17913, n17914, n17915, n17916, n17917, n17918, n17919,
         n17920, n17921, n17922, n17923, n17924, n17925, n17926, n17927,
         n17928, n17929, n17930, n17931, n17932, n17933, n17934, n17935,
         n17936, n17937, n17938, n17939, n17940, n17941, n17942, n17943,
         n17944, n17945, n17946, n17947, n17948, n17949, n17950, n17951,
         n17952, n17953, n17954, n17955, n17956, n17957, n17958, n17959,
         n17960, n17961, n17962, n17963, n17964, n17965, n17966, n17967,
         n17968, n17969, n17970, n17971, n17972, n17973, n17974, n17975,
         n17976, n17977, n17978, n17979, n17980, n17981, n17982, n17983,
         n17984, n17985, n17986, n17987, n17988, n17989, n17990, n17991,
         n17992, n17993, n17994, n17995, n17996, n17997, n17998, n17999,
         n18000, n18001, n18002, n18003, n18004, n18005, n18006, n18007,
         n18008, n18009, n18010, n18011, n18012, n18013, n18014, n18015,
         n18016, n18017, n18018, n18019, n18020, n18021, n18022, n18023,
         n18024, n18025, n18026, n18027, n18028, n18029, n18030, n18031,
         n18032, n18033, n18034, n18035, n18036, n18037, n18038, n18039,
         n18040, n18041, n18042, n18043, n18044, n18045, n18046, n18047,
         n18048, n18049, n18050, n18051, n18052, n18053, n18054, n18055,
         n18056, n18057, n18058, n18059, n18060, n18061, n18062, n18063,
         n18064, n18065, n18066, n18067, n18068, n18069, n18070, n18071,
         n18072, n18073, n18074, n18075, n18076, n18077, n18078, n18079,
         n18080, n18081, n18082, n18083, n18084, n18085, n18086, n18087,
         n18088, n18089, n18090, n18091, n18092, n18093, n18094, n18095,
         n18096, n18097, n18098, n18099, n18100, n18101, n18102, n18103,
         n18104, n18105, n18106, n18107, n18108, n18109, n18110, n18111,
         n18112, n18113, n18114, n18115, n18116, n18117, n18118, n18119,
         n18120, n18121, n18122, n18123, n18124, n18125, n18126, n18127,
         n18128, n18129, n18130, n18131, n18132, n18133, n18134, n18135,
         n18136, n18137, n18138, n18139, n18140, n18141, n18142, n18143,
         n18144, n18145, n18146, n18147, n18148, n18149, n18150, n18151,
         n18152, n18153, n18154, n18155, n18156, n18157, n18158, n18159,
         n18160, n18161, n18162, n18163, n18164, n18165, n18166, n18167,
         n18168, n18169, n18170, n18171, n18172, n18173, n18174, n18175,
         n18176, n18177, n18178, n18179, n18180, n18181, n18182, n18183,
         n18184, n18185, n18186, n18187, n18188, n18189, n18190, n18191,
         n18192, n18193, n18194, n18195, n18196, n18197, n18198, n18199,
         n18200, n18201, n18202, n18203, n18204, n18205, n18206, n18207,
         n18208, n18209, n18210, n18211, n18212, n18213, n18214, n18215,
         n18216, n18217, n18218, n18219, n18220, n18221, n18222, n18223,
         n18224, n18225, n18226, n18227, n18228, n18229, n18230, n18231,
         n18232, n18233, n18234, n18235, n18236, n18237, n18238, n18239,
         n18240, n18241, n18242, n18243, n18244, n18245, n18246, n18247,
         n18248, n18249, n18250, n18251, n18252, n18253, n18254, n18255,
         n18256, n18257, n18258, n18259, n18260, n18261, n18262, n18263,
         n18264, n18265, n18266, n18267, n18268, n18269, n18270, n18271,
         n18272, n18273, n18274, n18275, n18276, n18277, n18278, n18279,
         n18280, n18281, n18282, n18283, n18284, n18285, n18286, n18287,
         n18288, n18289, n18290, n18291, n18292, n18293, n18294, n18295,
         n18296, n18297, n18298, n18299, n18300, n18301, n18302, n18303,
         n18304, n18305, n18306, n18307, n18308, n18309, n18310, n18311,
         n18312, n18313, n18314, n18315, n18316, n18317, n18318, n18319,
         n18320, n18321, n18322, n18323, n18324, n18325, n18326, n18327,
         n18328, n18329, n18330, n18331, n18332, n18333, n18334, n18335,
         n18336, n18337, n18338, n18339, n18340, n18341, n18342, n18343,
         n18344, n18345, n18346, n18347, n18348, n18349, n18350, n18351,
         n18352, n18353, n18354, n18355, n18356, n18357, n18358, n18359,
         n18360, n18361, n18362, n18363, n18364, n18365, n18366, n18367,
         n18368, n18369, n18370, n18371, n18372, n18373, n18374, n18375,
         n18376, n18377, n18378, n18379, n18380, n18381, n18382, n18383,
         n18384, n18385, n18386, n18387, n18388, n18389, n18390, n18391,
         n18392, n18393, n18394, n18395, n18396, n18397, n18398, n18399,
         n18400, n18401, n18402, n18403, n18404, n18405, n18406, n18407,
         n18408, n18409, n18410, n18411, n18412, n18413, n18414, n18415,
         n18416, n18417, n18418, n18419, n18420, n18421, n18422, n18423,
         n18424, n18425, n18426, n18427, n18428, n18429, n18430, n18431,
         n18432, n18433, n18434, n18435, n18436, n18437, n18438, n18439,
         n18440, n18441, n18442, n18443, n18444, n18445, n18446, n18447,
         n18448, n18449, n18450, n18451, n18452, n18453, n18454, n18455,
         n18456, n18457, n18458, n18459, n18460, n18461, n18462, n18463,
         n18464, n18465, n18466, n18467, n18468, n18469, n18470, n18471,
         n18472, n18473, n18474, n18475, n18476, n18477, n18478, n18479,
         n18480, n18481, n18482, n18483, n18484, n18485, n18486, n18487,
         n18488, n18489, n18490, n18491, n18492, n18493, n18494, n18495,
         n18496, n18497, n18498, n18499, n18500, n18501, n18502, n18503,
         n18504, n18505, n18506, n18507, n18508, n18509, n18510, n18511,
         n18512, n18513, n18514, n18515, n18516, n18517, n18518, n18519,
         n18520, n18521, n18522, n18523, n18524, n18525, n18526, n18527,
         n18528, n18529, n18530, n18531, n18532, n18533, n18534, n18535,
         n18536, n18537, n18538, n18539, n18540, n18541, n18542, n18543,
         n18544, n18545, n18546, n18547, n18548, n18549, n18550, n18551,
         n18552, n18553, n18554, n18555, n18556, n18557, n18558, n18559,
         n18560, n18561, n18562, n18563, n18564, n18565, n18566, n18567,
         n18568, n18569, n18570, n18571, n18572, n18573, n18574, n18575,
         n18576, n18577, n18578, n18579, n18580, n18581, n18582, n18583,
         n18584, n18585, n18586, n18587, n18588, n18589, n18590, n18591,
         n18592, n18593, n18594, n18595, n18596, n18597, n18598, n18599,
         n18600, n18601, n18602, n18603, n18604, n18605, n18606, n18607,
         n18608, n18609, n18610, n18611, n18612, n18613, n18614, n18615,
         n18616, n18617, n18618, n18619, n18620, n18621, n18622, n18623,
         n18624, n18625, n18626, n18627, n18628, n18629, n18630, n18631,
         n18632, n18633, n18634, n18635, n18636, n18637, n18638, n18639,
         n18640, n18641, n18642, n18643, n18644, n18645, n18646, n18647,
         n18648, n18649, n18650, n18651, n18652, n18653, n18654, n18655,
         n18656, n18657, n18658, n18659, n18660, n18661, n18662, n18663,
         n18664, n18665, n18666, n18667, n18668, n18669, n18670, n18671,
         n18672, n18673, n18674, n18675, n18676, n18677, n18678, n18679,
         n18680, n18681, n18682, n18683, n18684, n18685, n18686, n18687,
         n18688, n18689, n18690, n18691, n18692, n18693, n18694, n18695,
         n18696, n18697, n18698, n18699, n18700, n18701, n18702, n18703,
         n18704, n18705, n18706, n18707, n18708, n18709, n18710, n18711,
         n18712, n18713, n18714, n18715, n18716, n18717, n18718, n18719,
         n18720, n18721, n18722, n18723, n18724, n18725, n18726, n18727,
         n18728, n18729, n18730, n18731, n18732, n18733, n18734, n18735,
         n18736, n18737, n18738, n18739, n18740, n18741, n18742, n18743,
         n18744, n18745, n18746, n18747, n18748, n18749, n18750, n18751,
         n18752, n18753, n18754, n18755, n18756, n18757, n18758, n18759,
         n18760, n18761, n18762, n18763, n18764, n18765, n18766, n18767,
         n18768, n18769, n18770, n18771, n18772, n18773, n18774, n18775,
         n18776, n18777, n18778, n18779, n18780, n18781, n18782, n18783,
         n18784, n18785, n18786, n18787, n18788, n18789, n18790, n18791,
         n18792, n18793, n18794, n18795, n18796, n18797, n18798, n18799,
         n18800, n18801, n18802, n18803, n18804, n18805, n18806, n18807,
         n18808, n18809, n18810, n18811, n18812, n18813, n18814, n18815,
         n18816, n18817, n18818, n18819, n18820, n18821, n18822, n18823,
         n18824, n18825, n18826, n18827, n18828, n18829, n18830, n18831,
         n18832, n18833, n18834, n18835, n18836, n18837, n18838, n18839,
         n18840, n18841, n18842, n18843, n18844, n18845, n18846, n18847,
         n18848, n18849, n18850, n18851, n18852, n18853, n18854, n18855,
         n18856, n18857, n18858, n18859, n18860, n18861, n18862, n18863,
         n18864, n18865, n18866, n18867, n18868, n18869, n18870, n18871,
         n18872, n18873, n18874, n18875, n18876, n18877, n18878, n18879,
         n18880, n18881, n18882, n18883, n18884, n18885, n18886, n18887,
         n18888, n18889, n18890, n18891, n18892, n18893, n18894, n18895,
         n18896, n18897, n18898, n18899, n18900, n18901, n18902, n18903,
         n18904, n18905, n18906, n18907, n18908, n18909, n18910, n18911,
         n18912, n18913, n18914, n18915, n18916, n18917, n18918, n18919,
         n18920, n18921, n18922, n18923, n18924, n18925, n18926, n18927,
         n18928, n18929, n18930, n18931, n18932, n18933, n18934, n18935,
         n18936, n18937, n18938, n18939, n18940, n18941, n18942, n18943,
         n18944, n18945, n18946, n18947, n18948, n18949, n18950, n18951,
         n18952, n18953, n18954, n18955, n18956, n18957, n18958, n18959,
         n18960, n18961, n18962, n18963, n18964, n18965, n18966, n18967,
         n18968, n18969, n18970, n18971, n18972, n18973, n18974, n18975,
         n18976, n18977, n18978, n18979, n18980, n18981, n18982, n18983,
         n18984, n18985, n18986, n18987, n18988, n18989, n18990, n18991,
         n18992, n18993, n18994, n18995, n18996, n18997, n18998, n18999,
         n19000, n19001, n19002, n19003, n19004, n19005, n19006, n19007,
         n19008, n19009, n19010, n19011, n19012, n19013, n19014, n19015,
         n19016, n19017, n19018, n19019, n19020, n19021, n19022, n19023,
         n19024, n19025, n19026, n19027, n19028, n19029, n19030, n19031,
         n19032, n19033, n19034, n19035, n19036, n19037, n19038, n19039,
         n19040, n19041, n19042, n19043, n19044, n19045, n19046, n19047,
         n19048, n19049, n19050, n19051, n19052, n19053, n19054, n19055,
         n19056, n19057, n19058, n19059, n19060, n19061, n19062, n19063,
         n19064, n19065, n19066, n19067, n19068, n19069, n19070, n19071,
         n19072, n19073, n19074, n19075, n19076, n19077, n19078, n19079,
         n19080, n19081, n19082, n19083, n19084, n19085, n19086, n19087,
         n19088, n19089, n19090, n19091, n19092, n19093, n19094, n19095,
         n19096, n19097, n19098, n19099, n19100, n19101, n19102, n19103,
         n19104, n19105, n19106, n19107, n19108, n19109, n19110, n19111,
         n19112, n19113, n19114, n19115, n19116, n19117, n19118, n19119,
         n19120, n19121, n19122, n19123, n19124, n19125, n19126, n19127,
         n19128, n19129, n19130, n19131, n19132, n19133, n19134, n19135,
         n19136, n19137, n19138, n19139, n19140, n19141, n19142, n19143,
         n19144, n19145, n19146, n19147, n19148, n19149, n19150, n19151,
         n19152, n19153, n19154, n19155, n19156, n19157, n19158, n19159,
         n19160, n19161, n19162, n19163, n19164, n19165, n19166, n19167,
         n19168, n19169, n19170, n19171, n19172, n19173, n19174, n19175,
         n19176, n19177, n19178, n19179, n19180, n19181, n19182, n19183,
         n19184, n19185, n19186, n19187, n19188, n19189, n19190, n19191,
         n19192, n19193, n19194, n19195, n19196, n19197, n19198, n19199,
         n19200, n19201, n19202, n19203, n19204, n19205, n19206, n19207,
         n19208, n19209, n19210, n19211, n19212, n19213, n19214, n19215,
         n19216, n19217, n19218, n19219, n19220, n19221, n19222, n19223,
         n19224, n19225, n19227, n19228, n19229, n19230, n19231, n19232,
         n19233, n19234, n19235, n19236, n19237, n19238, n19239, n19240,
         n19241, n19242, n19243, n19244, n19245, n19246, n19247, n19248,
         n19249, n19250, n19251, n19252, n19253, n19254, n19255, n19256,
         n19257, n19258, n19259, n19260, n19261, n19262, n19263, n19264,
         n19265, n19266, n19267, n19268, n19269, n19270, n19271, n19272,
         n19273, n19274, n19275, n19276, n19277, n19278, n19279, n19280,
         n19281, n19282, n19283, n19284, n19285, n19286, n19287, n19288,
         n19289, n19290, n19291, n19292, n19293, n19294, n19295, n19296,
         n19297, n19298, n19299, n19300, n19301, n19302, n19303, n19304,
         n19305, n19306, n19307, n19308, n19309, n19310, n19311, n19312,
         n19313, n19314, n19315, n19316, n19317, n19318, n19319, n19320,
         n19321, n19322, n19323, n19324, n19325, n19326, n19327, n19328,
         n19329, n19330, n19331, n19332, n19333, n19334, n19335, n19336,
         n19337, n19338, n19339, n19340, n19341, n19342, n19343, n19344,
         n19345, n19346, n19347, n19348, n19349, n19350, n19351, n19352,
         n19353, n19354, n19355, n19356, n19357, n19358, n19359, n19360,
         n19361, n19362, n19363, n19364, n19365, n19366, n19367, n19368,
         n19369, n19370, n19371, n19372, n19373, n19374, n19375, n19376,
         n19377, n19378, n19379, n19380, n19381, n19382, n19383, n19384,
         n19385, n19386, n19387, n19388, n19389, n19390, n19391, n19392,
         n19393, n19394, n19395, n19396, n19397, n19398, n19399, n19400,
         n19401, n19402, n19403, n19404, n19405, n19406, n19407, n19408,
         n19409, n19410, n19411, n19412, n19413, n19414, n19415, n19416,
         n19417, n19418, n19419, n19420, n19421, n19422, n19423, n19424,
         n19425, n19426, n19427, n19428, n19429, n19430, n19431, n19432,
         n19433, n19434, n19435, n19436, n19437, n19438, n19439, n19440,
         n19441, n19442, n19443, n19444, n19445, n19446, n19447, n19448,
         n19449, n19450, n19451, n19452, n19453, n19454, n19455, n19456,
         n19457, n19458, n19459, n19460, n19461, n19462, n19463, n19464,
         n19465, n19466, n19467, n19468, n19469, n19470, n19471, n19472,
         n19473, n19474, n19475, n19476, n19477, n19478, n19479, n19480,
         n19481, n19482, n19483, n19484, n19485, n19486, n19487, n19488,
         n19489, n19490, n19491, n19492, n19493, n19494, n19495, n19496,
         n19497, n19498, n19499, n19500, n19501, n19502, n19503, n19504,
         n19505, n19506, n19507, n19508, n19509, n19510, n19511, n19512,
         n19513, n19514, n19515, n19516, n19517, n19518, n19519, n19520,
         n19521, n19522, n19523, n19524, n19525, n19526, n19527, n19528,
         n19529, n19530, n19531, n19532, n19533, n19534, n19535, n19536,
         n19537, n19538, n19539, n19540, n19541, n19542, n19543, n19544,
         n19545, n19546, n19547, n19548, n19549, n19550, n19551, n19552,
         n19553, n19554, n19555, n19556, n19557, n19558, n19559, n19560,
         n19561, n19562, n19563, n19564, n19565, n19566, n19567, n19568,
         n19569, n19570, n19571, n19572, n19573, n19574, n19575, n19576,
         n19577, n19578, n19579, n19580, n19581, n19582, n19583, n19584,
         n19585, n19586, n19587, n19588, n19589, n19590, n19591, n19592,
         n19593, n19594, n19595, n19596, n19597, n19598, n19599, n19600,
         n19601, n19602, n19603, n19604, n19605, n19606, n19607, n19608,
         n19609, n19610, n19611, n19612, n19613, n19614, n19615, n19616,
         n19617, n19618, n19619, n19620, n19621, n19622, n19623, n19624,
         n19625, n19626, n19627, n19628, n19629, n19630, n19631, n19632,
         n19633, n19634, n19635, n19636, n19637, n19638, n19639, n19640,
         n19641, n19642, n19643, n19644, n19645, n19646, n19647, n19648,
         n19649, n19650, n19651, n19652, n19653, n19654, n19655, n19656,
         n19657, n19658, n19659, n19660, n19661, n19662, n19663, n19664,
         n19665, n19666, n19667, n19668, n19669, n19670, n19671, n19672,
         n19673, n19674, n19675, n19676, n19677, n19678, n19679, n19680,
         n19681, n19682, n19683, n19684, n19685, n19686, n19687, n19688,
         n19689, n19690, n19691, n19692, n19693, n19694, n19695, n19696,
         n19697, n19698, n19699, n19700, n19701, n19702, n19703, n19704,
         n19705, n19706, n19707, n19708, n19709, n19710, n19711, n19712,
         n19713, n19714, n19715, n19716, n19717, n19718, n19719, n19720,
         n19721, n19722, n19723, n19724, n19725, n19726, n19727, n19728,
         n19729, n19730, n19731, n19732, n19733, n19734, n19735, n19736,
         n19737, n19738, n19739, n19740, n19741, n19742, n19743, n19744,
         n19745, n19746, n19747, n19748, n19749, n19750, n19751, n19752,
         n19753, n19754, n19755, n19756, n19757, n19758, n19759, n19760,
         n19761, n19762, n19763, n19764, n19765, n19766, n19767, n19768,
         n19769, n19770, n19771, n19772, n19773, n19774, n19775, n19776,
         n19777, n19778, n19779, n19780, n19781, n19782, n19783, n19784,
         n19785, n19786, n19787, n19788, n19789, n19790, n19791, n19792,
         n19793, n19794, n19795, n19796, n19797, n19798, n19799, n19800,
         n19801, n19802, n19803, n19804, n19805, n19806, n19807, n19808,
         n19809, n19810, n19811, n19812, n19813, n19814, n19815, n19816,
         n19817, n19818, n19819, n19820, n19821, n19822, n19823, n19824,
         n19825, n19826, n19827, n19828, n19829, n19830, n19831, n19832,
         n19833, n19834, n19835, n19836, n19837, n19838, n19839, n19840,
         n19841, n19842, n19843, n19844, n19845, n19846, n19847, n19848,
         n19849, n19850, n19851, n19852, n19853, n19854, n19855, n19856,
         n19857, n19858, n19859, n19860, n19861, n19862, n19863, n19864,
         n19865, n19866, n19867, n19868, n19869, n19870, n19871, n19872,
         n19873, n19874, n19875, n19876, n19877, n19878, n19879, n19880,
         n19881, n19882, n19883, n19884, n19885, n19886, n19887, n19888,
         n19889, n19890, n19891, n19892, n19893, n19894, n19895, n19896,
         n19897, n19898, n19899, n19900, n19901, n19902, n19903, n19904,
         n19905, n19906, n19907, n19908, n19909, n19910, n19911, n19912,
         n19913, n19914, n19915, n19916, n19917, n19918, n19919, n19920,
         n19921, n19922, n19923, n19924, n19925, n19926, n19927, n19928,
         n19929, n19930, n19931, n19932, n19933, n19934, n19935, n19936,
         n19937, n19938, n19939, n19940, n19941, n19942, n19943, n19944,
         n19945, n19946, n19947, n19948, n19949, n19950, n19951, n19952,
         n19953, n19954, n19955, n19956, n19957, n19958, n19959, n19960,
         n19961, n19962, n19963, n19964, n19965, n19966, n19967, n19968,
         n19969, n19970, n19971, n19972, n19973, n19974, n19975, n19976,
         n19977, n19978, n19979, n19980, n19981, n19982, n19983, n19984,
         n19985, n19986, n19987, n19988, n19989, n19990, n19991, n19992,
         n19993, n19994, n19995, n19996, n19997, n19998, n19999, n20000,
         n20001, n20002, n20003, n20004, n20005, n20006, n20007, n20008,
         n20009, n20010, n20011, n20012, n20013, n20014, n20015, n20016,
         n20017, n20018, n20019, n20020, n20021, n20022, n20023, n20024,
         n20025, n20026, n20027, n20028, n20029, n20030, n20031, n20032,
         n20033, n20034, n20035, n20036, n20037, n20038, n20039, n20040,
         n20041, n20042, n20043, n20044, n20045, n20046, n20047, n20048,
         n20049, n20050, n20051, n20052, n20053, n20054, n20055, n20056,
         n20057, n20058, n20059, n20060, n20061, n20062, n20063, n20064,
         n20065, n20066, n20067, n20068, n20069, n20070, n20071, n20072,
         n20073, n20074, n20075, n20076, n20077, n20078, n20079, n20080,
         n20081, n20082, n20083, n20084, n20085, n20086, n20087, n20088,
         n20089, n20090, n20091, n20092, n20093, n20094, n20095, n20096,
         n20097, n20098, n20099, n20100, n20101, n20102, n20103, n20104,
         n20105, n20106, n20107, n20108, n20109, n20110, n20111, n20112,
         n20113, n20114, n20115, n20116, n20117, n20118, n20119, n20120,
         n20121, n20122, n20123, n20124, n20125, n20126, n20127, n20128,
         n20129, n20130, n20131, n20132, n20133, n20134, n20135, n20136,
         n20137, n20138, n20139, n20140, n20141, n20142, n20143, n20144,
         n20145, n20146, n20147, n20148, n20149, n20150, n20151, n20152,
         n20153, n20154, n20155, n20156, n20157, n20158, n20159, n20160,
         n20161, n20162, n20163, n20164, n20165, n20166, n20167, n20168,
         n20169, n20170, n20171, n20172, n20173, n20174, n20175, n20176,
         n20177, n20178, n20179, n20180, n20181, n20182, n20183, n20184,
         n20185, n20186, n20187, n20188, n20189, n20190, n20191, n20192,
         n20193, n20194, n20195, n20196, n20197, n20198, n20199, n20200,
         n20201, n20202, n20203, n20204, n20205, n20206, n20207, n20208,
         n20209, n20210, n20211, n20212, n20213, n20214, n20215, n20216,
         n20217, n20218, n20219, n20220, n20221, n20222, n20223, n20224,
         n20225, n20226, n20227, n20228, n20229, n20230, n20231, n20232,
         n20233, n20234, n20235, n20236, n20237, n20238, n20239, n20240,
         n20241, n20242, n20243, n20244, n20245, n20246, n20247, n20248,
         n20249, n20250, n20251, n20252, n20253, n20254, n20255, n20256,
         n20257, n20258, n20259, n20260, n20261, n20262, n20263, n20264,
         n20265, n20266, n20267, n20268, n20269, n20270, n20271, n20272,
         n20273, n20274, n20275, n20276, n20277, n20278, n20279, n20280,
         n20281, n20282, n20283, n20284, n20285, n20286, n20287, n20288,
         n20289, n20290, n20291, n20292, n20293, n20294, n20295, n20296,
         n20297, n20298, n20299, n20300, n20301, n20302, n20303, n20304,
         n20305, n20306, n20307, n20308, n20309, n20310, n20311, n20312,
         n20313, n20314, n20315, n20316, n20317, n20318, n20319, n20320,
         n20321, n20322, n20323, n20324, n20325, n20326, n20327, n20328,
         n20329, n20330, n20331, n20332, n20333, n20334, n20335, n20336,
         n20337, n20338, n20339, n20340, n20341, n20342, n20343, n20344,
         n20345, n20346, n20347, n20348, n20349, n20350, n20351, n20352,
         n20353, n20354, n20355, n20356, n20357, n20358, n20359, n20360,
         n20361, n20362, n20363, n20364, n20365, n20366, n20367, n20368,
         n20369, n20370, n20371, n20372, n20373, n20374, n20375, n20376,
         n20377, n20378, n20379, n20380, n20381, n20382, n20383, n20384,
         n20385, n20386, n20387, n20388, n20389, n20390, n20391, n20392,
         n20393, n20394, n20395, n20396, n20397, n20398, n20399, n20400,
         n20401, n20402, n20403, n20404, n20405, n20406, n20407, n20408,
         n20409, n20410, n20411, n20412, n20413, n20414, n20415, n20416,
         n20417, n20418, n20419, n20420, n20421, n20422, n20423, n20424,
         n20425, n20426, n20427, n20428, n20429, n20430, n20431, n20432,
         n20433, n20434, n20435, n20436, n20437, n20438, n20439, n20440,
         n20441, n20442, n20443, n20444, n20445, n20446, n20447, n20448,
         n20449, n20450, n20451, n20452, n20453, n20454, n20455, n20456,
         n20457, n20458, n20459, n20460, n20461, n20462, n20463, n20464,
         n20465, n20466, n20467, n20468, n20469, n20470, n20471, n20472,
         n20473, n20474, n20475, n20476, n20477, n20478, n20479, n20480,
         n20481, n20482, n20483, n20484, n20485, n20486, n20487, n20488,
         n20489, n20490, n20491, n20492, n20493, n20494, n20495, n20496,
         n20497, n20498, n20499, n20500, n20501, n20502, n20503, n20504,
         n20505, n20506, n20507, n20508, n20509, n20510, n20511, n20512,
         n20513, n20514, n20515, n20516, n20517, n20518, n20519, n20520,
         n20521, n20522, n20523, n20524, n20525, n20526, n20527, n20528,
         n20529, n20530, n20531, n20532, n20533, n20534, n20535, n20536,
         n20537, n20538, n20539, n20540, n20541, n20542, n20543, n20544,
         n20545, n20546, n20547, n20548, n20549, n20550, n20551, n20552,
         n20553, n20554, n20555, n20556, n20557, n20558, n20559, n20560,
         n20561, n20562, n20563, n20564, n20565, n20566, n20567, n20568,
         n20569, n20570, n20571, n20572, n20573, n20574, n20575, n20576,
         n20577, n20578, n20579, n20580, n20581, n20582, n20583, n20584,
         n20585, n20586, n20587, n20588, n20589, n20590, n20591, n20592,
         n20593, n20594, n20595, n20596, n20597, n20598, n20599, n20600,
         n20601, n20602, n20603, n20604, n20605, n20606, n20607, n20608,
         n20609, n20610, n20611, n20612, n20613, n20614, n20615, n20616,
         n20617, n20618, n20619, n20620, n20621, n20622, n20623, n20624,
         n20625, n20626, n20627, n20628, n20629, n20630, n20631, n20632,
         n20633, n20634, n20635, n20636, n20637, n20638, n20639, n20640,
         n20641, n20642, n20643, n20644, n20645, n20646, n20647, n20648,
         n20649, n20650, n20651, n20652, n20653, n20654, n20655, n20656,
         n20657, n20658, n20659, n20660, n20661, n20662, n20663, n20664,
         n20665, n20666, n20667, n20668, n20669, n20670, n20671, n20672,
         n20673, n20674, n20675, n20676, n20677, n20678, n20679, n20680,
         n20681, n20682, n20683, n20684, n20685, n20686, n20687, n20688,
         n20689, n20690, n20691, n20692, n20693, n20694, n20695, n20696,
         n20697, n20698, n20699, n20700, n20701, n20702, n20703, n20704,
         n20705, n20706, n20707, n20708, n20709, n20710, n20711, n20712,
         n20713, n20714, n20715, n20716, n20717, n20718, n20719, n20720,
         n20721, n20722, n20723, n20724, n20725, n20726, n20727, n20728,
         n20729, n20730, n20731, n20732, n20733, n20734, n20735, n20736,
         n20737, n20738, n20739, n20740, n20741, n20742, n20743, n20744,
         n20745, n20746, n20747, n20748, n20749, n20750, n20751, n20752,
         n20753, n20754, n20755, n20756, n20757, n20758, n20759, n20760,
         n20761, n20762, n20763, n20764, n20765, n20766, n20767, n20768,
         n20769, n20770, n20771, n20772, n20773, n20774, n20775, n20776,
         n20777, n20778, n20779, n20780, n20781, n20782, n20783, n20784,
         n20785, n20786, n20787, n20788, n20789, n20790, n20791, n20792,
         n20793, n20794, n20795, n20796, n20797, n20798, n20799, n20800,
         n20801, n20802, n20803, n20804, n20805, n20806, n20807, n20808,
         n20809, n20810, n20811, n20812, n20813, n20814, n20815, n20816,
         n20817, n20818, n20819, n20820, n20821, n20822, n20823, n20824,
         n20825, n20826, n20827, n20828, n20829, n20830, n20831, n20832,
         n20833, n20834, n20835, n20836, n20837, n20838, n20839, n20840,
         n20841, n20842, n20843, n20844, n20845, n20846, n20847, n20848,
         n20849, n20850, n20851, n20852, n20853, n20854, n20855, n20856,
         n20857, n20858, n20859, n20860, n20861, n20862, n20863, n20864,
         n20865, n20866, n20867, n20868, n20869, n20870, n20871, n20872,
         n20873, n20874, n20875, n20876, n20877, n20878, n20879, n20880,
         n20881, n20882, n20883, n20884, n20885, n20886, n20887, n20888,
         n20889, n20890, n20891, n20892, n20893, n20894, n20895, n20896,
         n20897, n20898, n20899, n20900, n20901, n20902, n20903, n20904,
         n20905, n20906, n20907, n20908, n20909, n20910, n20911, n20912,
         n20913, n20914, n20915, n20916, n20917, n20918, n20919, n20920,
         n20921, n20922, n20923, n20924, n20925, n20926, n20927, n20928,
         n20929, n20930, n20931, n20932, n20933, n20934, n20935, n20936,
         n20937, n20938, n20939, n20940, n20941, n20942, n20943, n20944,
         n20945, n20946, n20947, n20948, n20949, n20950, n20951, n20952,
         n20953, n20954, n20955, n20956, n20957, n20958, n20959, n20960,
         n20961, n20962, n20963, n20964, n20965, n20966, n20967, n20968,
         n20969, n20970, n20971, n20972, n20973, n20974, n20975, n20976,
         n20977, n20978, n20979, n20980, n20981, n20982, n20983, n20984,
         n20985, n20986, n20987, n20988, n20989, n20990, n20991, n20992,
         n20993, n20994, n20995, n20996, n20997, n20998, n20999, n21000,
         n21001, n21002, n21003, n21004, n21005, n21006, n21007, n21008,
         n21009, n21010, n21011, n21012, n21013, n21014, n21015, n21016,
         n21017, n21018, n21019, n21020, n21021, n21022, n21023, n21024,
         n21025, n21026, n21027, n21028, n21029, n21030, n21031, n21032,
         n21033, n21034, n21035, n21036, n21037, n21038, n21039, n21040,
         n21041, n21042, n21043, n21044, n21045, n21046, n21047, n21048,
         n21049, n21050, n21051, n21052, n21053, n21054, n21055, n21056,
         n21057, n21058, n21059, n21060, n21061, n21062, n21063, n21064,
         n21065, n21066, n21067, n21068, n21069, n21070, n21071, n21072,
         n21073, n21074, n21075, n21076, n21077, n21078, n21079, n21080,
         n21081, n21082, n21083, n21084, n21085, n21086, n21087, n21088,
         n21089, n21090, n21091, n21092, n21093, n21094, n21095, n21096,
         n21097, n21098, n21099, n21100, n21101, n21102, n21103, n21104,
         n21105, n21106, n21107, n21108, n21109, n21110, n21111, n21112,
         n21113, n21114, n21115, n21116, n21117, n21118, n21119, n21120,
         n21121, n21122, n21123, n21124, n21125, n21126, n21127, n21128,
         n21129, n21130, n21131, n21132, n21133, n21134, n21135, n21136,
         n21137, n21138, n21139, n21140, n21141, n21142, n21143, n21144,
         n21145, n21146, n21147, n21148, n21149, n21150, n21151, n21152,
         n21153, n21154, n21155, n21156, n21157, n21158, n21159, n21160,
         n21161, n21162, n21163, n21164, n21165, n21166, n21167, n21168,
         n21169, n21170, n21171, n21172, n21173, n21174, n21175, n21176,
         n21177, n21178, n21179, n21180, n21181, n21182, n21183, n21184,
         n21185, n21186, n21187, n21188, n21189, n21190, n21191, n21192,
         n21193, n21194, n21195, n21196, n21197, n21198, n21199, n21200,
         n21201, n21202, n21203, n21204, n21205, n21206, n21207, n21208,
         n21209, n21210, n21211, n21212, n21213, n21214, n21215, n21216,
         n21217, n21218, n21219, n21220, n21221, n21222, n21223, n21224,
         n21225, n21226, n21227, n21228, n21229, n21230, n21231, n21232,
         n21233, n21234, n21235, n21236, n21237, n21238, n21239, n21240,
         n21241, n21242, n21243, n21244, n21245, n21246, n21247, n21248,
         n21249, n21250, n21251, n21252, n21253, n21254, n21255, n21256,
         n21257, n21258, n21259, n21260, n21261, n21262, n21263, n21264,
         n21265, n21266, n21267, n21268, n21269, n21270, n21271, n21272,
         n21273, n21274, n21275, n21276, n21277, n21278, n21279, n21280,
         n21281, n21282, n21283, n21284, n21285, n21286, n21287, n21288,
         n21289, n21290, n21291, n21292, n21293, n21294, n21295, n21296,
         n21297, n21298, n21299, n21300, n21301, n21302, n21303, n21304,
         n21305, n21306, n21307, n21308, n21309, n21310, n21311, n21312,
         n21313, n21314, n21315, n21316, n21317, n21318, n21319, n21320,
         n21321, n21322, n21323, n21324, n21325, n21326, n21327, n21328,
         n21329, n21330, n21331, n21332, n21333, n21334, n21335, n21336,
         n21337, n21338, n21339, n21340, n21341, n21342, n21343, n21344,
         n21345, n21346, n21347, n21348, n21349, n21350, n21351, n21352,
         n21353, n21354, n21355, n21356, n21357, n21358, n21359, n21360,
         n21361, n21362, n21363, n21364, n21365, n21366, n21367, n21368,
         n21369, n21370, n21371, n21372, n21373, n21374, n21375, n21376,
         n21377, n21378, n21379, n21380, n21381, n21382, n21383, n21384,
         n21385, n21386, n21387, n21388, n21389, n21390, n21391, n21392,
         n21393, n21394, n21395, n21396, n21397, n21398, n21399, n21400,
         n21401, n21402, n21403, n21404, n21405, n21406, n21407, n21408,
         n21409, n21410, n21411, n21412, n21413, n21414, n21415, n21416,
         n21417, n21418, n21419, n21420, n21421, n21422, n21423, n21424,
         n21425, n21426, n21427, n21428, n21429, n21430, n21431, n21432,
         n21433, n21434, n21435, n21436, n21437, n21438, n21439, n21440,
         n21441, n21442, n21443, n21444, n21445, n21446, n21447, n21448,
         n21449, n21450, n21451, n21452, n21453, n21454, n21455, n21456,
         n21457, n21458, n21459, n21460, n21461, n21462, n21463, n21464,
         n21465, n21466, n21467, n21468, n21469, n21470, n21471, n21472,
         n21473, n21474, n21475, n21476, n21477, n21478, n21479, n21480,
         n21481, n21482, n21483, n21484, n21485, n21486, n21487, n21488,
         n21489, n21490, n21491, n21492, n21493, n21494, n21495, n21496,
         n21497, n21498, n21499, n21500, n21501, n21502, n21503, n21504,
         n21505, n21506, n21507, n21508, n21509, n21510, n21511, n21512,
         n21513, n21514, n21515, n21516, n21517, n21518, n21519, n21520,
         n21521, n21522, n21523, n21524, n21525, n21526, n21527, n21528,
         n21529, n21530, n21531, n21532, n21533, n21534, n21535, n21536,
         n21537, n21538, n21539, n21540, n21541, n21542, n21543, n21544,
         n21545, n21546, n21547, n21548, n21549, n21550, n21551, n21552,
         n21553, n21554, n21555, n21556, n21557, n21558, n21559, n21560,
         n21561, n21562, n21563, n21564, n21565, n21566, n21567, n21568,
         n21569, n21570, n21571, n21572, n21573, n21574, n21575, n21576,
         n21577, n21578, n21579, n21580, n21581, n21582, n21583, n21584,
         n21585, n21586, n21587, n21588, n21589, n21590, n21591, n21592,
         n21593, n21594, n21595, n21596, n21597, n21598, n21599, n21600,
         n21601, n21602, n21603, n21604, n21605, n21606, n21607, n21608,
         n21609, n21610, n21611, n21612, n21613, n21614, n21615, n21616,
         n21617, n21618, n21619, n21620, n21621, n21622, n21623, n21624,
         n21625, n21626, n21627, n21628, n21629, n21630, n21631, n21632,
         n21633, n21634, n21635, n21636, n21637, n21638, n21639, n21640,
         n21641, n21642, n21643, n21644, n21645, n21646, n21647, n21648,
         n21649, n21650, n21651, n21652, n21653, n21654, n21655, n21656,
         n21657, n21658, n21659, n21660, n21661, n21662, n21663, n21664,
         n21665, n21666, n21667, n21668, n21669, n21670, n21671, n21672,
         n21673, n21674, n21675, n21676, n21677, n21678, n21679, n21680,
         n21681, n21682, n21683, n21684, n21685, n21686, n21687, n21688,
         n21689, n21690, n21691, n21692, n21693, n21694, n21695, n21696,
         n21697, n21698, n21699, n21700, n21701, n21702, n21703, n21704,
         n21705, n21706, n21707, n21708, n21709, n21710, n21711, n21712,
         n21713, n21714, n21715, n21716, n21717, n21718, n21719, n21720,
         n21721, n21722, n21723, n21724, n21725, n21726, n21727, n21728,
         n21729, n21730, n21731, n21732, n21733, n21734, n21735, n21736,
         n21737, n21738, n21739, n21740, n21741, n21742, n21743, n21744,
         n21745, n21746, n21747, n21748, n21749, n21750, n21751, n21752,
         n21753, n21754, n21755, n21756, n21757, n21758, n21759, n21760,
         n21761, n21762, n21763, n21764, n21765, n21766, n21767, n21768,
         n21769, n21770, n21771, n21772, n21773, n21774, n21775, n21776,
         n21777, n21778, n21779, n21780, n21781, n21782, n21783, n21784,
         n21785, n21786, n21787, n21788, n21789, n21790, n21791, n21792,
         n21793, n21794, n21795, n21796, n21797, n21798, n21799, n21800,
         n21801, n21802, n21803, n21804, n21805, n21806, n21807, n21808,
         n21809, n21810, n21811, n21812, n21813, n21814, n21815, n21816,
         n21817, n21818, n21819, n21820, n21821, n21822, n21823, n21824,
         n21825, n21826, n21827, n21828, n21829, n21830, n21831, n21832,
         n21833, n21834, n21835, n21836, n21837, n21838, n21839, n21840,
         n21841, n21842, n21843, n21844, n21845, n21846, n21847, n21848,
         n21849, n21850, n21851, n21852, n21853, n21854, n21855, n21856,
         n21857, n21858, n21859, n21860, n21861, n21862, n21863, n21864,
         n21865, n21866, n21867, n21868, n21869, n21870, n21871, n21872,
         n21873, n21874, n21875, n21876, n21877, n21878, n21879, n21880,
         n21881, n21882, n21883, n21884, n21885, n21886, n21887, n21888,
         n21889, n21890, n21891, n21892, n21893, n21894, n21895, n21896,
         n21897, n21898, n21899, n21900, n21901, n21902, n21903, n21904,
         n21905, n21906, n21907, n21908, n21909, n21910, n21911, n21912,
         n21913, n21914, n21915, n21916, n21917, n21918, n21919, n21920,
         n21921, n21922, n21923, n21924, n21925, n21926, n21927, n21928,
         n21929, n21930, n21931, n21932, n21933, n21934, n21935, n21936,
         n21937, n21938, n21939, n21940, n21941, n21942, n21943, n21944,
         n21945, n21946, n21947, n21948, n21949, n21950, n21951, n21952,
         n21953, n21954, n21955, n21956, n21957, n21958, n21959, n21960,
         n21961, n21962, n21963, n21964, n21965, n21966, n21967, n21968,
         n21969, n21970, n21971, n21972, n21973, n21974, n21975, n21976,
         n21977, n21978, n21979, n21980, n21981, n21982, n21983, n21984,
         n21985, n21986, n21987, n21988, n21989, n21990, n21991, n21992,
         n21993, n21994, n21995, n21996, n21997, n21998, n21999, n22000,
         n22001, n22002, n22003, n22004, n22005, n22006, n22007, n22008,
         n22009, n22010, n22011, n22012, n22013, n22014, n22015, n22016,
         n22017, n22018, n22019, n22020, n22021, n22022, n22023, n22024,
         n22025, n22026, n22027, n22028, n22029, n22030, n22031, n22032,
         n22033, n22034, n22035, n22036, n22037, n22038, n22039, n22040,
         n22041, n22042, n22043, n22044, n22045, n22046, n22047, n22048,
         n22049, n22050, n22051, n22052, n22053, n22054, n22055, n22056,
         n22057, n22058, n22059, n22060, n22061, n22062, n22063, n22064,
         n22065, n22066, n22067, n22068, n22069, n22070, n22071, n22072,
         n22073, n22074, n22075, n22076, n22077, n22078, n22079, n22080,
         n22081, n22082, n22083, n22084, n22085, n22086, n22087, n22088,
         n22089, n22090, n22091, n22092, n22093, n22094, n22095, n22096,
         n22097, n22098, n22099, n22100, n22101, n22102, n22103, n22104,
         n22105, n22106, n22107, n22108, n22109, n22110, n22111, n22112,
         n22113, n22114, n22115, n22116, n22117, n22118, n22119, n22120,
         n22121, n22122, n22123, n22124, n22125, n22126, n22127, n22128,
         n22129, n22130, n22131, n22132, n22133, n22134, n22135, n22136,
         n22137, n22138, n22139, n22140, n22141, n22142, n22143, n22144,
         n22145, n22146, n22147, n22148, n22149, n22150, n22151, n22152,
         n22153, n22154, n22155, n22156, n22157, n22158, n22159, n22160,
         n22161, n22162, n22163, n22164, n22165, n22166, n22167, n22168,
         n22169, n22170, n22171, n22172, n22173, n22174, n22175, n22176,
         n22177, n22178, n22179, n22180, n22181, n22182, n22183, n22184,
         n22185, n22186, n22187, n22188, n22189, n22190, n22191, n22192,
         n22193, n22194, n22195, n22196, n22197, n22198, n22199, n22200,
         n22201, n22202, n22203, n22204, n22205, n22206, n22207, n22208,
         n22209, n22210, n22211, n22212, n22213, n22214, n22215, n22216,
         n22217, n22218, n22219, n22220, n22221;

  INV_X1 U11055 ( .A(n20391), .ZN(n20577) );
  INV_X2 U11056 ( .A(n20171), .ZN(n14680) );
  AND3_X1 U11057 ( .A1(n13305), .A2(n16684), .A3(n13058), .ZN(n13323) );
  CLKBUF_X1 U11058 ( .A(n11963), .Z(n12101) );
  INV_X1 U11059 ( .A(n13058), .ZN(n18090) );
  BUF_X2 U11060 ( .A(n12763), .Z(n15131) );
  NOR2_X1 U11061 ( .A1(n14555), .A2(n14554), .ZN(n20687) );
  AND2_X1 U11062 ( .A1(n16058), .A2(n12681), .ZN(n13366) );
  CLKBUF_X1 U11063 ( .A(n13367), .Z(n13343) );
  AND2_X1 U11064 ( .A1(n13107), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12898) );
  AND2_X1 U11065 ( .A1(n12873), .A2(n13041), .ZN(n12903) );
  AND2_X1 U11066 ( .A1(n13482), .A2(n13211), .ZN(n13354) );
  NOR2_X1 U11067 ( .A1(n18804), .A2(n14624), .ZN(n14661) );
  CLKBUF_X2 U11068 ( .A(n11540), .Z(n12263) );
  BUF_X2 U11069 ( .A(n10965), .Z(n10975) );
  CLKBUF_X1 U11070 ( .A(n14561), .Z(n17286) );
  CLKBUF_X2 U11071 ( .A(n10960), .Z(n17545) );
  CLKBUF_X2 U11072 ( .A(n10965), .Z(n10976) );
  CLKBUF_X2 U11073 ( .A(n14549), .Z(n10966) );
  CLKBUF_X1 U11074 ( .A(n10960), .Z(n10977) );
  BUF_X2 U11075 ( .A(n14682), .Z(n17540) );
  AND2_X1 U11076 ( .A1(n14298), .A2(n13747), .ZN(n21319) );
  CLKBUF_X1 U11077 ( .A(n14601), .Z(n10961) );
  CLKBUF_X2 U11078 ( .A(n14594), .Z(n10960) );
  NAND2_X1 U11079 ( .A1(n12384), .A2(n13732), .ZN(n12532) );
  CLKBUF_X3 U11080 ( .A(n14604), .Z(n10967) );
  INV_X2 U11081 ( .A(n14684), .ZN(n10965) );
  NAND2_X1 U11082 ( .A1(n14298), .A2(n13905), .ZN(n11180) );
  CLKBUF_X3 U11083 ( .A(n14681), .Z(n10968) );
  INV_X2 U11084 ( .A(n13732), .ZN(n14298) );
  INV_X1 U11086 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n21260) );
  AND2_X4 U11087 ( .A1(n13977), .A2(n13587), .ZN(n11585) );
  INV_X1 U11088 ( .A(n10950), .ZN(n10951) );
  INV_X1 U11089 ( .A(n10950), .ZN(n10954) );
  INV_X1 U11090 ( .A(n10950), .ZN(n10953) );
  INV_X1 U11091 ( .A(n13142), .ZN(n16067) );
  OAI22_X2 U11092 ( .A1(n20095), .A2(n14243), .B1(n16787), .B2(n13898), .ZN(
        n22089) );
  NAND2_X2 U11093 ( .A1(n20009), .A2(n14376), .ZN(n13898) );
  AOI21_X1 U11094 ( .B1(n12810), .B2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A(
        n12817), .ZN(n12819) );
  NOR2_X1 U11095 ( .A1(n20816), .A2(n21260), .ZN(n14682) );
  OR3_X1 U11096 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n20163), .ZN(n17208) );
  NAND2_X1 U11097 ( .A1(n14173), .A2(n11611), .ZN(n13570) );
  NAND2_X1 U11098 ( .A1(n13443), .A2(n11477), .ZN(n15436) );
  OAI211_X1 U11099 ( .C1(n11123), .C2(n16098), .A(n16095), .B(n11120), .ZN(
        n13172) );
  INV_X1 U11100 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12681) );
  AND2_X1 U11101 ( .A1(n14811), .A2(n14817), .ZN(n19204) );
  CLKBUF_X2 U11102 ( .A(n14601), .Z(n17505) );
  INV_X1 U11104 ( .A(n11640), .ZN(n14173) );
  AND2_X1 U11105 ( .A1(n15303), .A2(n15302), .ZN(n15306) );
  NOR2_X1 U11106 ( .A1(n16110), .A2(n16109), .ZN(n16108) );
  NOR3_X1 U11107 ( .A1(P3_STATEBS16_REG_SCAN_IN), .A2(n17954), .A3(n20798), 
        .ZN(n17802) );
  NAND2_X1 U11108 ( .A1(n17894), .A2(n17573), .ZN(n17883) );
  AND2_X1 U11109 ( .A1(n14678), .A2(n20807), .ZN(n16698) );
  INV_X1 U11110 ( .A(n11012), .ZN(n17205) );
  AND2_X1 U11111 ( .A1(n15596), .A2(n15595), .ZN(n10987) );
  NAND2_X1 U11112 ( .A1(n11136), .A2(n11135), .ZN(n15055) );
  NAND2_X1 U11113 ( .A1(n16131), .A2(n16132), .ZN(n16126) );
  INV_X1 U11114 ( .A(n18090), .ZN(n19605) );
  NAND2_X1 U11115 ( .A1(n11130), .A2(n12807), .ZN(n12838) );
  INV_X2 U11116 ( .A(n14730), .ZN(n20216) );
  NAND2_X1 U11117 ( .A1(n20769), .A2(P3_EAX_REG_16__SCAN_IN), .ZN(n20760) );
  NAND2_X1 U11118 ( .A1(n20638), .A2(P3_EAX_REG_7__SCAN_IN), .ZN(n20778) );
  INV_X2 U11119 ( .A(n20687), .ZN(n20711) );
  OR3_X1 U11120 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n14524), .ZN(n10949) );
  NAND2_X1 U11121 ( .A1(n11190), .A2(n13615), .ZN(n10950) );
  INV_X1 U11122 ( .A(n10950), .ZN(n10952) );
  NOR2_X2 U11123 ( .A1(n17706), .A2(n20990), .ZN(n20856) );
  NOR2_X2 U11124 ( .A1(n15134), .A2(n15133), .ZN(n15143) );
  XNOR2_X2 U11125 ( .A(n14897), .B(n14853), .ZN(n14893) );
  NAND2_X2 U11126 ( .A1(n14833), .A2(n14832), .ZN(n14897) );
  XNOR2_X2 U11127 ( .A(n11794), .B(n11146), .ZN(n12388) );
  NOR2_X1 U11128 ( .A1(n18804), .A2(n14622), .ZN(n20795) );
  AND2_X2 U11129 ( .A1(n12645), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n14026) );
  BUF_X4 U11130 ( .A(n11930), .Z(n10955) );
  BUF_X4 U11131 ( .A(n11930), .Z(n10956) );
  INV_X2 U11133 ( .A(n16061), .ZN(n10957) );
  NAND2_X2 U11134 ( .A1(n12875), .A2(n14027), .ZN(n16061) );
  NAND2_X2 U11135 ( .A1(n12822), .A2(n12821), .ZN(n13815) );
  INV_X4 U11136 ( .A(n10949), .ZN(n10958) );
  INV_X4 U11137 ( .A(n10949), .ZN(n10959) );
  NOR2_X1 U11138 ( .A1(n20163), .A2(n14522), .ZN(n14594) );
  NOR2_X1 U11139 ( .A1(n14523), .A2(n20824), .ZN(n14601) );
  NOR2_X2 U11140 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11500) );
  NAND2_X1 U11142 ( .A1(n13443), .A2(n11477), .ZN(n10963) );
  NOR2_X1 U11143 ( .A1(n16599), .A2(n16583), .ZN(n16582) );
  OAI21_X1 U11144 ( .B1(n15376), .B2(n15325), .A(n15374), .ZN(n11114) );
  NOR2_X1 U11145 ( .A1(n12378), .A2(n15513), .ZN(n15512) );
  OAI21_X1 U11146 ( .B1(n15897), .B2(n15881), .A(n10992), .ZN(n11212) );
  NAND2_X1 U11147 ( .A1(n11416), .A2(n11414), .ZN(n16304) );
  NAND2_X1 U11148 ( .A1(n14923), .A2(n14922), .ZN(n15996) );
  INV_X4 U11149 ( .A(n15994), .ZN(n15881) );
  INV_X2 U11151 ( .A(n12469), .ZN(n15994) );
  AND2_X1 U11152 ( .A1(n14811), .A2(n14818), .ZN(n14967) );
  AND2_X1 U11153 ( .A1(n14811), .A2(n14819), .ZN(n19235) );
  NAND2_X1 U11154 ( .A1(n21222), .A2(n21006), .ZN(n21141) );
  OR2_X1 U11155 ( .A1(n15102), .A2(n15101), .ZN(n15104) );
  BUF_X4 U11156 ( .A(n18403), .Z(n10964) );
  NAND2_X1 U11158 ( .A1(n14628), .A2(n14627), .ZN(n14679) );
  NOR2_X2 U11159 ( .A1(n21106), .A2(n17568), .ZN(n17774) );
  OR2_X1 U11160 ( .A1(n13725), .A2(n11444), .ZN(n11447) );
  NOR2_X1 U11161 ( .A1(n20104), .A2(n17148), .ZN(n21256) );
  INV_X4 U11162 ( .A(n12787), .ZN(n15227) );
  BUF_X2 U11163 ( .A(n13323), .Z(n15456) );
  NOR4_X1 U11164 ( .A1(n14615), .A2(n14623), .A3(n14632), .A4(n14658), .ZN(
        n14678) );
  AND3_X1 U11165 ( .A1(n13241), .A2(n14002), .A3(n13498), .ZN(n13647) );
  INV_X2 U11166 ( .A(n15131), .ZN(n16684) );
  INV_X4 U11167 ( .A(n15139), .ZN(n15420) );
  INV_X1 U11168 ( .A(n12384), .ZN(n12523) );
  NAND4_X1 U11169 ( .A1(n11536), .A2(n11535), .A3(n11534), .A4(n11533), .ZN(
        n11640) );
  NAND2_X1 U11170 ( .A1(n11095), .A2(n11093), .ZN(n12751) );
  NAND2_X1 U11171 ( .A1(n12730), .A2(n12729), .ZN(n14994) );
  CLKBUF_X2 U11172 ( .A(n11653), .Z(n12247) );
  CLKBUF_X2 U11173 ( .A(n11676), .Z(n12127) );
  BUF_X2 U11174 ( .A(n14549), .Z(n10971) );
  BUF_X2 U11175 ( .A(n11554), .Z(n12264) );
  CLKBUF_X2 U11176 ( .A(n11641), .Z(n12269) );
  INV_X4 U11177 ( .A(n13142), .ZN(n16058) );
  CLKBUF_X2 U11178 ( .A(n11834), .Z(n12270) );
  AND2_X4 U11179 ( .A1(n14026), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n16064) );
  BUF_X2 U11180 ( .A(n11584), .Z(n12218) );
  NAND2_X1 U11181 ( .A1(n20180), .A2(n20822), .ZN(n20816) );
  INV_X1 U11182 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13211) );
  NAND2_X1 U11183 ( .A1(n16332), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n16466) );
  NAND2_X1 U11184 ( .A1(n11450), .A2(n12506), .ZN(n15833) );
  NOR2_X1 U11185 ( .A1(n16319), .A2(n11161), .ZN(n16332) );
  AND2_X1 U11186 ( .A1(n16317), .A2(n16318), .ZN(n11161) );
  AND2_X1 U11187 ( .A1(n11429), .A2(n11091), .ZN(n15373) );
  AOI211_X1 U11188 ( .C1(n20005), .C2(n15739), .A(n15738), .B(n15737), .ZN(
        n15740) );
  NAND2_X1 U11189 ( .A1(n11092), .A2(n15283), .ZN(n11429) );
  XNOR2_X1 U11190 ( .A(n15512), .B(n12295), .ZN(n12519) );
  NAND2_X1 U11191 ( .A1(n11430), .A2(n15283), .ZN(n16600) );
  AOI21_X1 U11192 ( .B1(n15513), .B2(n12378), .A(n15512), .ZN(n15721) );
  NAND2_X1 U11193 ( .A1(n10983), .A2(n15541), .ZN(n15736) );
  OR2_X1 U11194 ( .A1(n15583), .A2(n11028), .ZN(n21603) );
  OR2_X1 U11195 ( .A1(n15641), .A2(n15539), .ZN(n21649) );
  XNOR2_X1 U11196 ( .A(n13117), .B(n11484), .ZN(n16110) );
  OR2_X1 U11197 ( .A1(n16304), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n16306) );
  INV_X1 U11198 ( .A(n20731), .ZN(n20727) );
  NOR2_X1 U11199 ( .A1(n15551), .A2(n15576), .ZN(n15572) );
  AND2_X1 U11200 ( .A1(n15602), .A2(n15604), .ZN(n15596) );
  OAI211_X1 U11201 ( .C1(n15268), .C2(n15272), .A(n11439), .B(n15271), .ZN(
        n16404) );
  NOR2_X2 U11202 ( .A1(n15377), .A2(n15319), .ZN(n16107) );
  NAND2_X1 U11203 ( .A1(n20712), .A2(P3_EAX_REG_25__SCAN_IN), .ZN(n20719) );
  NOR2_X1 U11204 ( .A1(n14460), .A2(n11054), .ZN(n11923) );
  AND2_X1 U11205 ( .A1(n12467), .A2(n12468), .ZN(n11457) );
  NAND2_X1 U11206 ( .A1(n14991), .A2(n14990), .ZN(n15266) );
  AND2_X1 U11207 ( .A1(n15784), .A2(n11034), .ZN(n11459) );
  AND2_X1 U11208 ( .A1(n15960), .A2(n12460), .ZN(n15784) );
  AND2_X1 U11209 ( .A1(n15795), .A2(n15797), .ZN(n15930) );
  AND2_X1 U11210 ( .A1(n15800), .A2(n15798), .ZN(n15960) );
  INV_X1 U11211 ( .A(n14940), .ZN(n11136) );
  NAND2_X1 U11212 ( .A1(n17815), .A2(n21115), .ZN(n17710) );
  CLKBUF_X1 U11213 ( .A(n17872), .Z(n10978) );
  AND2_X1 U11214 ( .A1(n11456), .A2(n12421), .ZN(n11024) );
  NAND2_X1 U11215 ( .A1(n14512), .A2(n14494), .ZN(n14794) );
  NAND2_X1 U11216 ( .A1(n17816), .A2(n21191), .ZN(n17815) );
  OAI21_X1 U11217 ( .B1(n17829), .B2(n21176), .A(n11277), .ZN(n17872) );
  NAND2_X1 U11218 ( .A1(n13775), .A2(n11813), .ZN(n13914) );
  XNOR2_X1 U11219 ( .A(n12414), .B(n12406), .ZN(n13873) );
  INV_X1 U11220 ( .A(n17966), .ZN(n17954) );
  XNOR2_X1 U11221 ( .A(n12431), .B(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n14313) );
  AND2_X1 U11222 ( .A1(n14981), .A2(n14980), .ZN(n14984) );
  AND2_X1 U11223 ( .A1(n11267), .A2(n11356), .ZN(n17816) );
  XNOR2_X1 U11224 ( .A(n12433), .B(n11854), .ZN(n12441) );
  OR2_X1 U11225 ( .A1(n11405), .A2(n16269), .ZN(n11402) );
  NAND2_X1 U11226 ( .A1(n12433), .A2(n12452), .ZN(n12469) );
  NOR2_X2 U11227 ( .A1(n21106), .A2(n20929), .ZN(n21203) );
  NAND2_X1 U11228 ( .A1(n17630), .A2(n17578), .ZN(n17849) );
  AND4_X1 U11229 ( .A1(n14815), .A2(n14814), .A3(n14813), .A4(n14812), .ZN(
        n14829) );
  AND4_X1 U11230 ( .A1(n14827), .A2(n14826), .A3(n14825), .A4(n14824), .ZN(
        n14828) );
  AND4_X1 U11231 ( .A1(n14837), .A2(n14836), .A3(n14835), .A4(n14834), .ZN(
        n14848) );
  NOR2_X1 U11232 ( .A1(n19335), .A2(n14840), .ZN(n14841) );
  NAND2_X1 U11233 ( .A1(n11783), .A2(n11787), .ZN(n14157) );
  NAND2_X1 U11234 ( .A1(n12404), .A2(n12403), .ZN(n13762) );
  NAND2_X1 U11235 ( .A1(n17883), .A2(n17884), .ZN(n17630) );
  NAND2_X1 U11236 ( .A1(n11804), .A2(n11805), .ZN(n11207) );
  NOR2_X2 U11237 ( .A1(n14821), .A2(n11250), .ZN(n15112) );
  INV_X1 U11238 ( .A(n11805), .ZN(n11802) );
  OAI21_X1 U11239 ( .B1(n17892), .B2(n17891), .A(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n17563) );
  AND2_X1 U11240 ( .A1(n14811), .A2(n14822), .ZN(n19214) );
  NAND2_X1 U11241 ( .A1(n20711), .A2(n20686), .ZN(n20785) );
  CLKBUF_X1 U11242 ( .A(n12371), .Z(n15694) );
  NAND2_X1 U11243 ( .A1(n11691), .A2(n11184), .ZN(n11805) );
  XNOR2_X1 U11244 ( .A(n19971), .B(n12401), .ZN(n13695) );
  NAND2_X1 U11245 ( .A1(n11668), .A2(n11784), .ZN(n11184) );
  NAND2_X1 U11246 ( .A1(n11737), .A2(n11736), .ZN(n13897) );
  NOR2_X2 U11247 ( .A1(n21457), .A2(n21463), .ZN(n21488) );
  NOR2_X2 U11248 ( .A1(n14244), .A2(n13905), .ZN(n21913) );
  NOR3_X2 U11249 ( .A1(n15707), .A2(n11611), .A3(n15506), .ZN(n15684) );
  AND2_X1 U11250 ( .A1(n15301), .A2(n15300), .ZN(n15303) );
  NAND2_X1 U11251 ( .A1(n19970), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n19971) );
  OR2_X1 U11252 ( .A1(n12394), .A2(n11667), .ZN(n11691) );
  NAND2_X1 U11253 ( .A1(n12852), .A2(n12851), .ZN(n18526) );
  NAND2_X1 U11254 ( .A1(n12393), .A2(n12392), .ZN(n19970) );
  NAND2_X1 U11255 ( .A1(n17909), .A2(n14776), .ZN(n17557) );
  OAI21_X1 U11256 ( .B1(n14112), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n11652), 
        .ZN(n12394) );
  AND2_X1 U11257 ( .A1(n12821), .A2(n11128), .ZN(n12839) );
  NOR2_X2 U11258 ( .A1(n19462), .A2(n19673), .ZN(n19463) );
  NOR2_X1 U11259 ( .A1(n14872), .A2(n14873), .ZN(n14953) );
  OR2_X1 U11260 ( .A1(n11010), .A2(n15218), .ZN(n15225) );
  NOR2_X2 U11261 ( .A1(n19509), .A2(n19673), .ZN(n16677) );
  XNOR2_X1 U11262 ( .A(n13819), .B(n13818), .ZN(n13816) );
  AOI21_X1 U11263 ( .B1(n11794), .B2(n11793), .A(n12450), .ZN(n11784) );
  NAND2_X1 U11264 ( .A1(n11119), .A2(n12785), .ZN(n11130) );
  OR2_X1 U11265 ( .A1(n14499), .A2(n14498), .ZN(n14872) );
  NAND2_X1 U11266 ( .A1(n12848), .A2(n12847), .ZN(n11119) );
  NAND2_X1 U11267 ( .A1(n11147), .A2(n11686), .ZN(n11794) );
  CLKBUF_X1 U11268 ( .A(n18507), .Z(n18473) );
  NOR2_X1 U11269 ( .A1(n21238), .A2(n21117), .ZN(n21133) );
  AOI21_X1 U11270 ( .B1(n12808), .B2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n12809), .ZN(n12818) );
  INV_X1 U11271 ( .A(n11639), .ZN(n13900) );
  NAND2_X1 U11272 ( .A1(n12549), .A2(n12548), .ZN(n14258) );
  AND2_X1 U11273 ( .A1(n11026), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11693) );
  OAI211_X1 U11274 ( .C1(n13822), .C2(n18602), .A(n12827), .B(n12826), .ZN(
        n13818) );
  NOR2_X1 U11275 ( .A1(n15163), .A2(n15162), .ZN(n15182) );
  OR2_X1 U11276 ( .A1(n15161), .A2(n15160), .ZN(n15163) );
  OR3_X1 U11277 ( .A1(n20673), .A2(n14621), .A3(n14631), .ZN(n14625) );
  AOI21_X1 U11278 ( .B1(n14012), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n11132), 
        .ZN(n12766) );
  NAND2_X1 U11279 ( .A1(n11017), .A2(n11447), .ZN(n11141) );
  NAND2_X1 U11280 ( .A1(n17949), .A2(n14754), .ZN(n17939) );
  NAND2_X1 U11281 ( .A1(n10980), .A2(n11133), .ZN(n14012) );
  OR2_X1 U11282 ( .A1(n11628), .A2(n13747), .ZN(n11137) );
  AND2_X1 U11283 ( .A1(n10988), .A2(n11067), .ZN(n10990) );
  NAND2_X1 U11284 ( .A1(n11571), .A2(n13662), .ZN(n13725) );
  OAI211_X1 U11285 ( .C1(n12787), .C2(n12777), .A(n11397), .B(n12778), .ZN(
        n12780) );
  AND2_X1 U11286 ( .A1(n15142), .A2(n11282), .ZN(n10988) );
  INV_X1 U11287 ( .A(n15436), .ZN(n15440) );
  OR2_X1 U11288 ( .A1(n14612), .A2(n20795), .ZN(n14662) );
  NOR2_X1 U11289 ( .A1(n20661), .A2(n14766), .ZN(n14741) );
  AND2_X1 U11290 ( .A1(n11609), .A2(n11608), .ZN(n11610) );
  AND2_X1 U11291 ( .A1(n19013), .A2(n18925), .ZN(n14612) );
  NAND2_X1 U11292 ( .A1(n12592), .A2(n12613), .ZN(n13680) );
  AND2_X1 U11293 ( .A1(n14002), .A2(n12772), .ZN(n13242) );
  NOR2_X1 U11294 ( .A1(n20687), .A2(n18885), .ZN(n14666) );
  OR2_X1 U11295 ( .A1(n13570), .A2(n12532), .ZN(n13748) );
  NAND3_X1 U11296 ( .A1(n14543), .A2(n14542), .A3(n14541), .ZN(n20166) );
  INV_X1 U11297 ( .A(n13184), .ZN(n13498) );
  NOR2_X2 U11298 ( .A1(n14588), .A2(n14587), .ZN(n18925) );
  INV_X2 U11299 ( .A(n19009), .ZN(n18884) );
  INV_X1 U11300 ( .A(n12751), .ZN(n19464) );
  NOR2_X1 U11301 ( .A1(n14994), .A2(n13265), .ZN(n12772) );
  AOI211_X1 U11302 ( .C1(n17547), .C2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A(
        n14540), .B(n14539), .ZN(n14541) );
  INV_X1 U11303 ( .A(n14999), .ZN(n19559) );
  INV_X1 U11304 ( .A(n12357), .ZN(n11631) );
  INV_X1 U11305 ( .A(n14008), .ZN(n12702) );
  INV_X1 U11306 ( .A(n14994), .ZN(n19676) );
  NOR2_X1 U11307 ( .A1(n12751), .A2(n14999), .ZN(n12755) );
  OR2_X1 U11308 ( .A1(n11560), .A2(n11559), .ZN(n12384) );
  OR2_X2 U11309 ( .A1(n11603), .A2(n11602), .ZN(n13732) );
  NAND2_X2 U11310 ( .A1(U214), .A2(n20037), .ZN(n20100) );
  INV_X2 U11311 ( .A(U214), .ZN(n20089) );
  NAND2_X1 U11312 ( .A1(n12745), .A2(n12744), .ZN(n14999) );
  NAND2_X1 U11313 ( .A1(n12701), .A2(n12700), .ZN(n14008) );
  NAND2_X1 U11314 ( .A1(n12728), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12729) );
  AND4_X1 U11315 ( .A1(n11504), .A2(n11503), .A3(n11502), .A4(n11501), .ZN(
        n11505) );
  AND4_X1 U11316 ( .A1(n11520), .A2(n11519), .A3(n11518), .A4(n11517), .ZN(
        n11536) );
  AND4_X1 U11317 ( .A1(n11528), .A2(n11527), .A3(n11526), .A4(n11525), .ZN(
        n11534) );
  AND4_X1 U11318 ( .A1(n11532), .A2(n11531), .A3(n11530), .A4(n11529), .ZN(
        n11533) );
  AND4_X1 U11319 ( .A1(n11575), .A2(n11574), .A3(n11573), .A4(n11572), .ZN(
        n11593) );
  AND4_X1 U11320 ( .A1(n11579), .A2(n11578), .A3(n11577), .A4(n11576), .ZN(
        n11592) );
  AND4_X1 U11321 ( .A1(n11583), .A2(n11582), .A3(n11581), .A4(n11580), .ZN(
        n11591) );
  AND4_X1 U11322 ( .A1(n11589), .A2(n11588), .A3(n11587), .A4(n11586), .ZN(
        n11590) );
  AND4_X1 U11323 ( .A1(n11498), .A2(n11497), .A3(n11496), .A4(n11495), .ZN(
        n11506) );
  AND4_X1 U11324 ( .A1(n11524), .A2(n11523), .A3(n11522), .A4(n11521), .ZN(
        n11535) );
  NOR2_X1 U11325 ( .A1(n16978), .A2(n18167), .ZN(n16407) );
  INV_X2 U11326 ( .A(n19008), .ZN(U215) );
  CLKBUF_X3 U11327 ( .A(n14572), .Z(n17539) );
  INV_X2 U11328 ( .A(n13625), .ZN(n11878) );
  NAND2_X2 U11329 ( .A1(n22219), .A2(n16774), .ZN(n16736) );
  CLKBUF_X2 U11330 ( .A(n14556), .Z(n17548) );
  BUF_X2 U11331 ( .A(n11537), .Z(n11962) );
  INV_X2 U11332 ( .A(n17208), .ZN(n17538) );
  CLKBUF_X1 U11333 ( .A(n16226), .Z(n16678) );
  BUF_X2 U11334 ( .A(n12866), .Z(n16062) );
  NAND2_X2 U11335 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(n21734), .ZN(n17137) );
  AND2_X2 U11336 ( .A1(n10957), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12885) );
  CLKBUF_X2 U11337 ( .A(n18030), .Z(n21248) );
  INV_X2 U11338 ( .A(n17208), .ZN(n10972) );
  INV_X2 U11339 ( .A(n21386), .ZN(n10970) );
  NOR3_X1 U11340 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n14523), .ZN(n14561) );
  NAND2_X1 U11341 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n20181), .ZN(
        n14730) );
  AND2_X1 U11342 ( .A1(n13614), .A2(n16011), .ZN(n11653) );
  NOR2_X1 U11343 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n20816), .ZN(
        n14681) );
  NOR2_X1 U11344 ( .A1(n20163), .A2(n20824), .ZN(n14556) );
  NOR2_X1 U11345 ( .A1(n20798), .A2(n17967), .ZN(n18030) );
  AND2_X2 U11346 ( .A1(n14026), .A2(n13211), .ZN(n12866) );
  OR2_X1 U11347 ( .A1(n14523), .A2(n16689), .ZN(n11012) );
  NAND2_X1 U11348 ( .A1(n20829), .A2(n20825), .ZN(n20163) );
  AND2_X1 U11349 ( .A1(n16011), .A2(n13977), .ZN(n11834) );
  NAND2_X2 U11350 ( .A1(n12875), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13142) );
  AND2_X2 U11351 ( .A1(n11493), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11190) );
  NAND2_X1 U11352 ( .A1(n20822), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n14522) );
  NOR2_X1 U11353 ( .A1(n11493), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11499) );
  NAND2_X1 U11354 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n21260), .ZN(
        n20824) );
  NOR2_X2 U11355 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n16011) );
  INV_X1 U11356 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n12647) );
  INV_X1 U11357 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n12646) );
  NOR2_X2 U11358 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n12873) );
  INV_X1 U11359 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n14027) );
  AND2_X1 U11360 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14013) );
  AND2_X1 U11361 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13977) );
  AND2_X1 U11362 ( .A1(n11492), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13614) );
  AND2_X1 U11363 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13613) );
  NAND2_X1 U11364 ( .A1(n11458), .A2(n12467), .ZN(n15777) );
  NAND2_X1 U11365 ( .A1(n13900), .A2(n11637), .ZN(n11696) );
  NAND3_X1 U11366 ( .A1(n11802), .A2(n11476), .A3(n13897), .ZN(n11763) );
  NAND2_X2 U11367 ( .A1(n14467), .A2(n12439), .ZN(n14876) );
  NAND2_X1 U11368 ( .A1(n11696), .A2(n14151), .ZN(n14112) );
  NAND3_X2 U11369 ( .A1(n11619), .A2(n11612), .A3(n14298), .ZN(n12348) );
  AND2_X1 U11370 ( .A1(n11499), .A2(n13977), .ZN(n11540) );
  NOR2_X1 U11371 ( .A1(n14524), .A2(n20824), .ZN(n14549) );
  AND2_X1 U11372 ( .A1(n11500), .A2(n13587), .ZN(n10974) );
  AND2_X1 U11373 ( .A1(n11500), .A2(n13587), .ZN(n11584) );
  NAND2_X2 U11374 ( .A1(n11611), .A2(n11631), .ZN(n13634) );
  AND2_X1 U11375 ( .A1(n11499), .A2(n11500), .ZN(n11554) );
  XNOR2_X2 U11376 ( .A(n19995), .B(n21347), .ZN(n21339) );
  OAI21_X2 U11377 ( .B1(n20186), .B2(n17760), .A(n19009), .ZN(n17768) );
  NOR2_X2 U11378 ( .A1(n15715), .A2(n15714), .ZN(n15716) );
  AOI211_X2 U11379 ( .C1(n20022), .C2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .A(
        n21341), .B(n19996), .ZN(n19997) );
  AND2_X2 U11380 ( .A1(n15088), .A2(n15704), .ZN(n15697) );
  AOI21_X4 U11381 ( .B1(n15085), .B2(n11960), .A(n11959), .ZN(n15088) );
  AOI22_X2 U11382 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n16018), .B1(n16017), 
        .B2(n13554), .ZN(n18403) );
  NAND2_X1 U11383 ( .A1(n15540), .A2(n11475), .ZN(n11474) );
  INV_X1 U11384 ( .A(n15640), .ZN(n11475) );
  INV_X1 U11385 ( .A(n16995), .ZN(n11092) );
  AND4_X1 U11386 ( .A1(n13359), .A2(n13358), .A3(n13357), .A4(n13356), .ZN(
        n13383) );
  AND2_X1 U11387 ( .A1(n12852), .A2(n11032), .ZN(n14819) );
  NAND2_X1 U11388 ( .A1(n11275), .A2(n11273), .ZN(n14628) );
  INV_X1 U11389 ( .A(n21281), .ZN(n11275) );
  NAND2_X1 U11390 ( .A1(n20113), .A2(n14629), .ZN(n11273) );
  NAND2_X1 U11391 ( .A1(n15747), .A2(n11220), .ZN(n11460) );
  NAND2_X1 U11392 ( .A1(n11607), .A2(n13747), .ZN(n11444) );
  BUF_X1 U11393 ( .A(n11545), .Z(n12271) );
  NAND2_X1 U11394 ( .A1(n14001), .A2(n12702), .ZN(n12705) );
  INV_X1 U11395 ( .A(n16352), .ZN(n11252) );
  INV_X1 U11396 ( .A(n16341), .ZN(n11251) );
  NAND2_X1 U11397 ( .A1(n16522), .A2(n11155), .ZN(n11154) );
  NAND2_X1 U11398 ( .A1(n15130), .A2(n15129), .ZN(n15275) );
  INV_X1 U11399 ( .A(n15269), .ZN(n15129) );
  INV_X1 U11400 ( .A(n11245), .ZN(n15130) );
  AND3_X1 U11401 ( .A1(n12756), .A2(n12757), .A3(n12755), .ZN(n12765) );
  INV_X1 U11402 ( .A(n21458), .ZN(n11380) );
  AND2_X1 U11403 ( .A1(n11465), .A2(n15604), .ZN(n11187) );
  AND2_X1 U11404 ( .A1(n11466), .A2(n15552), .ZN(n11465) );
  INV_X1 U11405 ( .A(n12287), .ZN(n12256) );
  NOR2_X2 U11406 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n12291) );
  NAND2_X1 U11407 ( .A1(n15994), .A2(n11216), .ZN(n11215) );
  NAND2_X1 U11408 ( .A1(n11220), .A2(n15994), .ZN(n11217) );
  INV_X1 U11409 ( .A(n11082), .ZN(n11216) );
  NAND2_X1 U11410 ( .A1(n16743), .A2(n21321), .ZN(n11147) );
  OR2_X1 U11411 ( .A1(n13349), .A2(n13348), .ZN(n15017) );
  INV_X1 U11412 ( .A(n15280), .ZN(n15282) );
  AND2_X1 U11413 ( .A1(n11431), .A2(n11081), .ZN(n11428) );
  INV_X1 U11414 ( .A(n15220), .ZN(n16318) );
  INV_X1 U11415 ( .A(n16525), .ZN(n11354) );
  NAND2_X1 U11416 ( .A1(n15270), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11237) );
  INV_X1 U11417 ( .A(n13408), .ZN(n13394) );
  OR2_X1 U11418 ( .A1(n15266), .A2(n15264), .ZN(n11236) );
  AND2_X1 U11419 ( .A1(n12702), .A2(n19559), .ZN(n14002) );
  NAND2_X1 U11420 ( .A1(n11117), .A2(n11235), .ZN(n13995) );
  AND2_X1 U11421 ( .A1(n14807), .A2(n14816), .ZN(n11112) );
  NOR2_X1 U11422 ( .A1(n14816), .A2(n14807), .ZN(n14823) );
  INV_X1 U11423 ( .A(n13265), .ZN(n13058) );
  NAND2_X1 U11424 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n20825), .ZN(
        n14523) );
  AND3_X1 U11425 ( .A1(n11255), .A2(n11260), .A3(n11259), .ZN(n17738) );
  NOR2_X1 U11426 ( .A1(n17711), .A2(n17712), .ZN(n11258) );
  NOR2_X1 U11427 ( .A1(n17849), .A2(n11378), .ZN(n17579) );
  NAND2_X1 U11428 ( .A1(n17536), .A2(n11379), .ZN(n11378) );
  NAND2_X1 U11429 ( .A1(n20788), .A2(n20783), .ZN(n11310) );
  INV_X1 U11430 ( .A(n14645), .ZN(n14654) );
  AOI21_X1 U11431 ( .B1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n16711), .A(
        n14649), .ZN(n14655) );
  NAND2_X1 U11432 ( .A1(n14620), .A2(n14619), .ZN(n14631) );
  OR2_X1 U11433 ( .A1(n14618), .A2(n14617), .ZN(n14619) );
  NOR2_X1 U11434 ( .A1(n14622), .A2(n18844), .ZN(n20809) );
  OR2_X1 U11435 ( .A1(n13724), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n12637) );
  NAND2_X1 U11436 ( .A1(n11473), .A2(n15527), .ZN(n11472) );
  INV_X1 U11437 ( .A(n11474), .ZN(n11473) );
  NAND2_X1 U11438 ( .A1(n11145), .A2(n11052), .ZN(n12508) );
  NAND2_X1 U11439 ( .A1(n12422), .A2(n11024), .ZN(n11454) );
  INV_X1 U11440 ( .A(n14313), .ZN(n11456) );
  AND2_X1 U11441 ( .A1(n13735), .A2(n13468), .ZN(n16758) );
  AND2_X1 U11442 ( .A1(n10990), .A2(n15152), .ZN(n11281) );
  XNOR2_X1 U11443 ( .A(n16645), .B(n12857), .ZN(n13646) );
  AND2_X1 U11444 ( .A1(n11062), .A2(n12883), .ZN(n11425) );
  INV_X1 U11445 ( .A(n16029), .ZN(n13449) );
  NAND2_X1 U11446 ( .A1(n15279), .A2(n15278), .ZN(n16995) );
  NAND2_X1 U11447 ( .A1(n16286), .A2(n15479), .ZN(n16260) );
  NAND2_X1 U11448 ( .A1(n11102), .A2(n11101), .ZN(n15475) );
  NAND2_X1 U11449 ( .A1(n11398), .A2(n11403), .ZN(n11101) );
  NAND2_X1 U11450 ( .A1(n16270), .A2(n11103), .ZN(n11102) );
  AND2_X1 U11451 ( .A1(n11398), .A2(n16271), .ZN(n11103) );
  AND2_X1 U11452 ( .A1(n16187), .A2(n16175), .ZN(n16176) );
  NOR2_X2 U11453 ( .A1(n16090), .A2(n16081), .ZN(n16082) );
  OR2_X1 U11454 ( .A1(n16398), .A2(n15150), .ZN(n11418) );
  NAND2_X1 U11455 ( .A1(n19331), .A2(n19316), .ZN(n19252) );
  BUF_X1 U11456 ( .A(n12753), .Z(n12828) );
  INV_X1 U11457 ( .A(n19331), .ZN(n19673) );
  INV_X1 U11458 ( .A(n18804), .ZN(n20673) );
  XNOR2_X1 U11459 ( .A(n20783), .B(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n17959) );
  AOI22_X1 U11460 ( .A1(n17205), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n10958), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n14532) );
  AOI211_X1 U11461 ( .C1(n17546), .C2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A(
        n14530), .B(n14529), .ZN(n14531) );
  INV_X1 U11462 ( .A(n21271), .ZN(n21269) );
  AND2_X1 U11463 ( .A1(n19987), .A2(n19974), .ZN(n20005) );
  NAND2_X1 U11464 ( .A1(n18508), .A2(n17019), .ZN(n15452) );
  OR2_X1 U11465 ( .A1(n12848), .A2(n12847), .ZN(n12849) );
  INV_X1 U11466 ( .A(n12343), .ZN(n12320) );
  AOI21_X1 U11467 ( .B1(n11968), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A(
        n11164), .ZN(n11739) );
  AND2_X1 U11468 ( .A1(n11585), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n11164) );
  AOI21_X1 U11469 ( .B1(n12270), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .A(
        n11173), .ZN(n11646) );
  AND2_X1 U11470 ( .A1(n11585), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11173) );
  AOI21_X1 U11471 ( .B1(n11968), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .A(
        n11163), .ZN(n11654) );
  AND2_X1 U11472 ( .A1(n11585), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n11163) );
  AND2_X1 U11473 ( .A1(n11477), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n11396) );
  AND2_X1 U11474 ( .A1(n12338), .A2(n12331), .ZN(n12334) );
  AND2_X1 U11475 ( .A1(n11585), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n11176) );
  INV_X1 U11476 ( .A(n14951), .ZN(n11463) );
  CLKBUF_X1 U11477 ( .A(n11997), .Z(n11968) );
  AND2_X1 U11478 ( .A1(n11585), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(
        n11162) );
  AND2_X1 U11479 ( .A1(n11585), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n11175) );
  OR2_X2 U11480 ( .A1(n11763), .A2(n11762), .ZN(n11848) );
  AOI21_X1 U11481 ( .B1(n10956), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .A(
        n11168), .ZN(n11726) );
  AND2_X1 U11482 ( .A1(n11585), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n11168) );
  INV_X1 U11483 ( .A(n12302), .ZN(n12333) );
  AND2_X1 U11484 ( .A1(n11620), .A2(n13662), .ZN(n12482) );
  NOR2_X1 U11485 ( .A1(n18627), .A2(n19296), .ZN(n11132) );
  NAND2_X1 U11486 ( .A1(n12798), .A2(n13995), .ZN(n11098) );
  INV_X1 U11487 ( .A(n12765), .ZN(n12758) );
  NAND2_X1 U11488 ( .A1(n12746), .A2(n12751), .ZN(n12771) );
  NAND2_X1 U11489 ( .A1(n12769), .A2(n13058), .ZN(n14003) );
  INV_X1 U11490 ( .A(n14002), .ZN(n14000) );
  NAND2_X1 U11491 ( .A1(n13231), .A2(n11124), .ZN(n13232) );
  NAND2_X1 U11492 ( .A1(n12768), .A2(n12748), .ZN(n13231) );
  NOR2_X1 U11493 ( .A1(n20646), .A2(n14740), .ZN(n17567) );
  NAND2_X1 U11494 ( .A1(n11310), .A2(n20666), .ZN(n14765) );
  NOR2_X1 U11495 ( .A1(n11270), .A2(n11269), .ZN(n11268) );
  INV_X1 U11496 ( .A(n14610), .ZN(n11269) );
  AND3_X1 U11497 ( .A1(n14173), .A2(n11631), .A3(n11148), .ZN(n11149) );
  INV_X1 U11498 ( .A(n11447), .ZN(n11139) );
  NAND2_X1 U11499 ( .A1(n13739), .A2(n12348), .ZN(n11143) );
  AND2_X1 U11500 ( .A1(n12522), .A2(n13747), .ZN(n11381) );
  AOI21_X1 U11501 ( .B1(n12247), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .A(
        n11174), .ZN(n12048) );
  OR2_X1 U11502 ( .A1(n15561), .A2(n15619), .ZN(n11470) );
  NAND2_X1 U11503 ( .A1(n11861), .A2(n11462), .ZN(n15077) );
  NOR2_X1 U11504 ( .A1(n11221), .A2(n15741), .ZN(n11220) );
  NAND2_X1 U11505 ( .A1(n15597), .A2(n11299), .ZN(n11298) );
  INV_X1 U11506 ( .A(n15611), .ZN(n11299) );
  OR2_X1 U11507 ( .A1(n15881), .A2(n14934), .ZN(n12459) );
  NAND2_X1 U11508 ( .A1(n13663), .A2(n12613), .ZN(n12614) );
  AND2_X1 U11509 ( .A1(n14309), .A2(n11295), .ZN(n11294) );
  INV_X1 U11510 ( .A(n14257), .ZN(n11295) );
  INV_X1 U11511 ( .A(n14258), .ZN(n11293) );
  OAI21_X1 U11512 ( .B1(n14295), .B2(n12397), .A(n11053), .ZN(n12398) );
  INV_X1 U11513 ( .A(n12489), .ZN(n11723) );
  AND2_X1 U11514 ( .A1(n11003), .A2(n11285), .ZN(n11284) );
  INV_X1 U11515 ( .A(n15402), .ZN(n11285) );
  NOR2_X1 U11516 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13041) );
  INV_X1 U11517 ( .A(n11121), .ZN(n11120) );
  OAI21_X1 U11518 ( .B1(n11122), .B2(n16098), .A(n16088), .ZN(n11121) );
  NOR2_X1 U11519 ( .A1(n11353), .A2(n11079), .ZN(n11352) );
  INV_X1 U11520 ( .A(n16227), .ZN(n11353) );
  INV_X1 U11521 ( .A(n16140), .ZN(n11419) );
  OR2_X1 U11522 ( .A1(n13328), .A2(n11336), .ZN(n11335) );
  INV_X1 U11523 ( .A(n14137), .ZN(n11336) );
  INV_X1 U11524 ( .A(n14001), .ZN(n13241) );
  NOR2_X1 U11525 ( .A1(n16146), .A2(n11325), .ZN(n11324) );
  INV_X1 U11526 ( .A(n16155), .ZN(n11325) );
  NOR2_X1 U11527 ( .A1(n14516), .A2(n14219), .ZN(n11320) );
  NAND2_X1 U11528 ( .A1(n14859), .A2(n14858), .ZN(n15015) );
  NAND2_X1 U11529 ( .A1(n13443), .A2(n13058), .ZN(n11440) );
  AND2_X1 U11530 ( .A1(n11402), .A2(n11399), .ZN(n11398) );
  INV_X1 U11531 ( .A(n16257), .ZN(n11399) );
  NOR2_X1 U11532 ( .A1(n16101), .A2(n11328), .ZN(n11327) );
  INV_X1 U11533 ( .A(n16106), .ZN(n11328) );
  AND2_X1 U11534 ( .A1(n15343), .A2(n11412), .ZN(n11409) );
  NAND2_X1 U11535 ( .A1(n15297), .A2(n15298), .ZN(n11412) );
  NOR2_X1 U11536 ( .A1(n15297), .A2(n15298), .ZN(n11411) );
  NAND2_X1 U11537 ( .A1(n11154), .A2(n11153), .ZN(n16316) );
  AOI21_X1 U11538 ( .B1(n11155), .B2(n11157), .A(n11055), .ZN(n11153) );
  INV_X1 U11539 ( .A(n11432), .ZN(n11431) );
  OAI21_X1 U11540 ( .B1(n16996), .B2(n11433), .A(n16532), .ZN(n11432) );
  AND2_X1 U11541 ( .A1(n11415), .A2(n15158), .ZN(n11414) );
  NAND2_X1 U11542 ( .A1(n11046), .A2(n15150), .ZN(n11415) );
  AND2_X1 U11543 ( .A1(n11344), .A2(n11341), .ZN(n11340) );
  INV_X1 U11544 ( .A(n13686), .ZN(n11341) );
  AOI21_X1 U11545 ( .B1(n13681), .B2(n11037), .A(n11345), .ZN(n11344) );
  INV_X1 U11546 ( .A(n13684), .ZN(n11345) );
  INV_X1 U11547 ( .A(n13846), .ZN(n11309) );
  NAND2_X1 U11548 ( .A1(n15128), .A2(n15127), .ZN(n15269) );
  OR2_X1 U11549 ( .A1(n15126), .A2(n15125), .ZN(n15128) );
  NAND2_X1 U11550 ( .A1(n14985), .A2(n14984), .ZN(n11245) );
  INV_X1 U11551 ( .A(n14454), .ZN(n11333) );
  NAND2_X1 U11552 ( .A1(n14852), .A2(n14851), .ZN(n14853) );
  OR2_X1 U11553 ( .A1(n13290), .A2(n13289), .ZN(n13499) );
  NAND2_X1 U11554 ( .A1(n15131), .A2(n13266), .ZN(n13408) );
  AOI21_X1 U11555 ( .B1(n13689), .B2(n13310), .A(n13309), .ZN(n13327) );
  INV_X1 U11556 ( .A(n11335), .ZN(n11334) );
  AND2_X1 U11557 ( .A1(n18526), .A2(n18108), .ZN(n14817) );
  NAND2_X1 U11558 ( .A1(n12694), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12701) );
  AND2_X1 U11559 ( .A1(n18521), .A2(n14805), .ZN(n14818) );
  INV_X1 U11560 ( .A(n14810), .ZN(n14805) );
  NOR2_X1 U11561 ( .A1(n13180), .A2(n13206), .ZN(n13181) );
  NAND2_X1 U11562 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n20829), .ZN(
        n14524) );
  INV_X1 U11563 ( .A(n14719), .ZN(n11369) );
  NAND2_X1 U11564 ( .A1(n10961), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(
        n11372) );
  NAND2_X1 U11565 ( .A1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n11226), .ZN(
        n11225) );
  NOR2_X1 U11566 ( .A1(n20413), .A2(n11227), .ZN(n11226) );
  INV_X1 U11567 ( .A(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n11227) );
  NOR2_X1 U11568 ( .A1(n17774), .A2(n17883), .ZN(n17602) );
  XNOR2_X1 U11569 ( .A(n17600), .B(n11261), .ZN(n17895) );
  INV_X1 U11570 ( .A(n17572), .ZN(n11261) );
  NAND2_X1 U11571 ( .A1(n17914), .A2(n14758), .ZN(n14759) );
  NAND2_X1 U11572 ( .A1(n17933), .A2(n14772), .ZN(n14773) );
  OR2_X1 U11573 ( .A1(n21324), .A2(n12517), .ZN(n12521) );
  NOR2_X1 U11574 ( .A1(n14258), .A2(n14257), .ZN(n14310) );
  NAND2_X1 U11575 ( .A1(n12343), .A2(n12352), .ZN(n12344) );
  NAND2_X1 U11576 ( .A1(n11357), .A2(n11023), .ZN(n12345) );
  NAND2_X1 U11577 ( .A1(n11613), .A2(n11148), .ZN(n13657) );
  AOI21_X1 U11578 ( .B1(n12262), .B2(n12261), .A(n12260), .ZN(n12380) );
  NOR2_X1 U11579 ( .A1(n13657), .A2(n11180), .ZN(n13584) );
  NOR2_X1 U11580 ( .A1(n13662), .A2(n21910), .ZN(n11772) );
  AND2_X1 U11581 ( .A1(n12291), .A2(n15739), .ZN(n12213) );
  AND2_X1 U11582 ( .A1(n11187), .A2(n11059), .ZN(n11186) );
  INV_X1 U11583 ( .A(n15576), .ZN(n11188) );
  NAND2_X1 U11584 ( .A1(n15897), .A2(n11082), .ZN(n11219) );
  NAND2_X1 U11585 ( .A1(n12473), .A2(n15881), .ZN(n15747) );
  NAND2_X1 U11586 ( .A1(n11144), .A2(n12415), .ZN(n14098) );
  NAND2_X1 U11587 ( .A1(n13873), .A2(n13872), .ZN(n11144) );
  NAND2_X1 U11588 ( .A1(n12388), .A2(n12440), .ZN(n12393) );
  INV_X1 U11589 ( .A(n16740), .ZN(n16006) );
  OR2_X1 U11590 ( .A1(n14401), .A2(n13897), .ZN(n14158) );
  NOR2_X1 U11591 ( .A1(n21845), .A2(n21771), .ZN(n21898) );
  OR2_X1 U11592 ( .A1(n14401), .A2(n14107), .ZN(n21885) );
  OR2_X1 U11593 ( .A1(n14157), .A2(n21671), .ZN(n21884) );
  INV_X1 U11594 ( .A(n21885), .ZN(n21889) );
  NAND2_X1 U11595 ( .A1(n21321), .A2(n13904), .ZN(n21771) );
  AOI21_X1 U11596 ( .B1(n21877), .B2(P1_STATE2_REG_3__SCAN_IN), .A(n21771), 
        .ZN(n21918) );
  AND2_X1 U11597 ( .A1(n16772), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n16766) );
  AND2_X1 U11598 ( .A1(n15306), .A2(n11283), .ZN(n15411) );
  AND2_X1 U11599 ( .A1(n11284), .A2(n15404), .ZN(n11283) );
  AND2_X1 U11600 ( .A1(n13264), .A2(n13263), .ZN(n16525) );
  AND2_X1 U11601 ( .A1(n14789), .A2(n14449), .ZN(n11355) );
  NAND2_X1 U11602 ( .A1(n15014), .A2(n11278), .ZN(n15134) );
  AND3_X1 U11603 ( .A1(n14858), .A2(n13526), .A3(n11280), .ZN(n11278) );
  INV_X1 U11604 ( .A(n14807), .ZN(n16046) );
  OR2_X1 U11605 ( .A1(n15347), .A2(n15379), .ZN(n15377) );
  AND2_X1 U11606 ( .A1(n12882), .A2(n13891), .ZN(n12883) );
  NAND2_X1 U11607 ( .A1(n15383), .A2(n15323), .ZN(n16198) );
  NOR2_X1 U11608 ( .A1(n11314), .A2(n11313), .ZN(n11312) );
  INV_X1 U11609 ( .A(n14286), .ZN(n11313) );
  NAND2_X1 U11610 ( .A1(n11384), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n17000) );
  INV_X1 U11611 ( .A(n16987), .ZN(n11384) );
  NAND2_X1 U11612 ( .A1(n16407), .A2(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16987) );
  NOR2_X1 U11613 ( .A1(n13881), .A2(n13960), .ZN(n13961) );
  INV_X1 U11614 ( .A(n11130), .ZN(n11129) );
  NAND2_X1 U11615 ( .A1(n14810), .A2(n11151), .ZN(n12852) );
  INV_X1 U11616 ( .A(n11119), .ZN(n11151) );
  NOR2_X1 U11617 ( .A1(n15424), .A2(n11436), .ZN(n11435) );
  NAND2_X1 U11618 ( .A1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n11436) );
  NAND2_X1 U11619 ( .A1(n16107), .A2(n16106), .ZN(n16105) );
  NOR2_X1 U11620 ( .A1(n15424), .A2(n15325), .ZN(n11434) );
  NAND2_X1 U11621 ( .A1(n11114), .A2(n11113), .ZN(n16291) );
  NAND2_X1 U11622 ( .A1(n15376), .A2(n15325), .ZN(n11113) );
  AOI21_X1 U11623 ( .B1(n15221), .B2(n15220), .A(n11015), .ZN(n15222) );
  NAND2_X1 U11624 ( .A1(n11429), .A2(n11428), .ZN(n16327) );
  OR2_X1 U11625 ( .A1(n17033), .A2(n11241), .ZN(n16339) );
  NAND2_X1 U11626 ( .A1(n11242), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n11241) );
  INV_X1 U11627 ( .A(n11243), .ZN(n11242) );
  AND2_X1 U11628 ( .A1(n14450), .A2(n11045), .ZN(n16523) );
  NAND2_X1 U11629 ( .A1(n16522), .A2(n16521), .ZN(n16520) );
  AND2_X1 U11630 ( .A1(n14292), .A2(n14293), .ZN(n14450) );
  NOR2_X1 U11631 ( .A1(n13861), .A2(n14087), .ZN(n14292) );
  INV_X1 U11632 ( .A(n16609), .ZN(n11417) );
  NAND2_X1 U11633 ( .A1(n16406), .A2(n16405), .ZN(n11249) );
  NAND2_X1 U11634 ( .A1(n11438), .A2(n15274), .ZN(n16397) );
  NAND2_X1 U11635 ( .A1(n16404), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11438) );
  NAND2_X1 U11636 ( .A1(n11236), .A2(n11237), .ZN(n15273) );
  OR2_X1 U11637 ( .A1(n16645), .A2(n12858), .ZN(n12859) );
  OAI21_X2 U11638 ( .B1(n16669), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n16668), 
        .ZN(n19331) );
  AOI21_X1 U11639 ( .B1(n20577), .B2(n11198), .A(n11197), .ZN(n11196) );
  INV_X1 U11640 ( .A(n20548), .ZN(n11198) );
  AOI21_X1 U11641 ( .B1(n20577), .B2(n11206), .A(n11205), .ZN(n11204) );
  INV_X1 U11642 ( .A(n20525), .ZN(n11205) );
  INV_X1 U11643 ( .A(n20503), .ZN(n11206) );
  AOI21_X1 U11644 ( .B1(n20577), .B2(n11211), .A(n11210), .ZN(n11209) );
  INV_X1 U11645 ( .A(n20452), .ZN(n11211) );
  NAND2_X1 U11646 ( .A1(n20451), .A2(n20452), .ZN(n20460) );
  NOR2_X1 U11647 ( .A1(n20264), .A2(n11231), .ZN(n11230) );
  NAND2_X1 U11648 ( .A1(n20166), .A2(n20165), .ZN(n20169) );
  INV_X1 U11649 ( .A(n14726), .ZN(n11265) );
  NAND2_X1 U11650 ( .A1(n14589), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n11264) );
  INV_X1 U11651 ( .A(n14728), .ZN(n11266) );
  AOI21_X1 U11652 ( .B1(n20613), .B2(n20612), .A(n20611), .ZN(n20615) );
  NOR2_X1 U11653 ( .A1(n11038), .A2(n20485), .ZN(n17701) );
  XNOR2_X1 U11654 ( .A(n14773), .B(n20914), .ZN(n17922) );
  NAND2_X1 U11655 ( .A1(n17965), .A2(n17959), .ZN(n17956) );
  NAND2_X1 U11656 ( .A1(n11257), .A2(n11258), .ZN(n11255) );
  AOI22_X1 U11657 ( .A1(n17581), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B1(
        n21198), .B2(n17774), .ZN(n11356) );
  INV_X1 U11658 ( .A(n17583), .ZN(n11267) );
  NAND2_X1 U11659 ( .A1(n11254), .A2(n17937), .ZN(n17926) );
  OAI21_X1 U11660 ( .B1(n17939), .B2(n17938), .A(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n11254) );
  NAND2_X1 U11661 ( .A1(n17939), .A2(n17938), .ZN(n17937) );
  INV_X1 U11662 ( .A(n11310), .ZN(n14769) );
  NOR3_X1 U11663 ( .A1(n16696), .A2(n16695), .A3(n16694), .ZN(n21271) );
  NAND2_X1 U11664 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n21290), .ZN(n21310) );
  INV_X1 U11665 ( .A(n14625), .ZN(n11274) );
  NAND2_X1 U11666 ( .A1(n12639), .A2(n12640), .ZN(n11304) );
  AND2_X1 U11667 ( .A1(n12636), .A2(n12635), .ZN(n21633) );
  INV_X1 U11668 ( .A(n21648), .ZN(n21611) );
  INV_X1 U11669 ( .A(n21633), .ZN(n21646) );
  OR2_X1 U11670 ( .A1(n12521), .A2(n10970), .ZN(n21422) );
  AND2_X1 U11671 ( .A1(n19969), .A2(n15506), .ZN(n19961) );
  XNOR2_X1 U11672 ( .A(n12496), .B(n12495), .ZN(n13952) );
  NAND2_X1 U11673 ( .A1(n21655), .A2(n12486), .ZN(n19987) );
  INV_X1 U11674 ( .A(n11451), .ZN(n11450) );
  INV_X1 U11675 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n21877) );
  OR2_X1 U11676 ( .A1(n15004), .A2(n13444), .ZN(n16029) );
  AND2_X1 U11677 ( .A1(n14043), .A2(n18099), .ZN(n18653) );
  AND2_X1 U11678 ( .A1(n15484), .A2(n15483), .ZN(n18491) );
  XNOR2_X1 U11679 ( .A(n13646), .B(n13645), .ZN(n19168) );
  NAND2_X1 U11680 ( .A1(n16102), .A2(n11124), .ZN(n16167) );
  INV_X1 U11681 ( .A(n17055), .ZN(n17046) );
  NAND2_X1 U11682 ( .A1(n18653), .A2(n18090), .ZN(n17058) );
  AOI21_X1 U11683 ( .B1(n19113), .B2(n18622), .A(n15468), .ZN(n15469) );
  OAI211_X1 U11684 ( .C1(n15488), .C2(n16018), .A(n11479), .B(n15467), .ZN(
        n15468) );
  XNOR2_X1 U11685 ( .A(n15445), .B(n15444), .ZN(n18508) );
  AOI21_X1 U11686 ( .B1(n15475), .B2(n15476), .A(n11104), .ZN(n15423) );
  AOI21_X1 U11687 ( .B1(n16420), .B2(n18568), .A(n11349), .ZN(n11348) );
  OR2_X1 U11688 ( .A1(n16418), .A2(n16419), .ZN(n11349) );
  OR2_X1 U11689 ( .A1(n16083), .A2(n16082), .ZN(n18474) );
  NAND2_X1 U11690 ( .A1(n11400), .A2(n11402), .ZN(n16258) );
  NAND2_X1 U11691 ( .A1(n11100), .A2(n11401), .ZN(n11400) );
  AND2_X1 U11692 ( .A1(n15049), .A2(n15013), .ZN(n18568) );
  INV_X1 U11693 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19323) );
  OR2_X1 U11694 ( .A1(n16645), .A2(n13652), .ZN(n19147) );
  CLKBUF_X1 U11695 ( .A(n19316), .Z(n19332) );
  INV_X1 U11696 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n19203) );
  INV_X1 U11697 ( .A(n19168), .ZN(n19152) );
  NAND2_X1 U11698 ( .A1(n16640), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n16669) );
  NAND2_X1 U11699 ( .A1(n11193), .A2(n11196), .ZN(n20576) );
  OR2_X1 U11700 ( .A1(n20549), .A2(n20391), .ZN(n11193) );
  NAND2_X1 U11701 ( .A1(n20549), .A2(n20548), .ZN(n20565) );
  NAND2_X1 U11702 ( .A1(n11201), .A2(n11204), .ZN(n20534) );
  OR2_X1 U11703 ( .A1(n20502), .A2(n20391), .ZN(n11201) );
  NAND2_X1 U11704 ( .A1(n20502), .A2(n20503), .ZN(n20523) );
  CLKBUF_X1 U11705 ( .A(n20450), .Z(n20579) );
  NOR2_X1 U11706 ( .A1(n17781), .A2(n21057), .ZN(n21108) );
  NOR2_X1 U11707 ( .A1(n11611), .A2(n21321), .ZN(n12305) );
  NAND2_X1 U11708 ( .A1(n14298), .A2(n11611), .ZN(n12308) );
  NOR2_X1 U11709 ( .A1(n12320), .A2(n12319), .ZN(n12324) );
  AOI21_X1 U11710 ( .B1(n12263), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .A(
        n11169), .ZN(n12243) );
  AND2_X1 U11711 ( .A1(n11585), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(
        n11169) );
  AOI21_X1 U11712 ( .B1(n10956), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .A(
        n11172), .ZN(n12219) );
  AND2_X1 U11713 ( .A1(n11585), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n11172) );
  AOI21_X1 U11714 ( .B1(n11997), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .A(
        n11167), .ZN(n12159) );
  AND2_X1 U11715 ( .A1(n11585), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(
        n11167) );
  AOI21_X1 U11716 ( .B1(n11968), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A(
        n11165), .ZN(n12114) );
  AND2_X1 U11717 ( .A1(n11585), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n11165) );
  NAND2_X1 U11718 ( .A1(n11620), .A2(n11192), .ZN(n11621) );
  AND2_X1 U11719 ( .A1(n14173), .A2(n13662), .ZN(n11192) );
  AND2_X1 U11720 ( .A1(n13945), .A2(n13571), .ZN(n11445) );
  AND2_X1 U11721 ( .A1(n12348), .A2(n11142), .ZN(n11138) );
  NAND2_X1 U11722 ( .A1(n11616), .A2(n13747), .ZN(n11142) );
  NAND2_X1 U11723 ( .A1(n10959), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n11271) );
  OR2_X1 U11724 ( .A1(n13747), .A2(n21321), .ZN(n11707) );
  NAND2_X1 U11725 ( .A1(n11364), .A2(n11362), .ZN(n11361) );
  AOI21_X1 U11726 ( .B1(n12323), .B2(n12324), .A(n11363), .ZN(n11362) );
  NAND2_X1 U11727 ( .A1(n12326), .A2(n12325), .ZN(n11364) );
  NOR2_X1 U11728 ( .A1(n12341), .A2(n12327), .ZN(n11363) );
  AOI21_X1 U11729 ( .B1(n10956), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .A(
        n11171), .ZN(n12182) );
  AND2_X1 U11730 ( .A1(n11585), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(
        n11171) );
  AND2_X1 U11731 ( .A1(n11585), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n11174) );
  AOI21_X1 U11732 ( .B1(n12271), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A(
        n11177), .ZN(n12002) );
  AND2_X1 U11733 ( .A1(n11585), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n11177) );
  AOI21_X1 U11734 ( .B1(n11968), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .A(
        n11166), .ZN(n11970) );
  AND2_X1 U11735 ( .A1(n11585), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n11166) );
  AOI21_X1 U11736 ( .B1(n10956), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .A(
        n11170), .ZN(n11931) );
  AND2_X1 U11737 ( .A1(n11585), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n11170) );
  OR2_X1 U11738 ( .A1(n11640), .A2(n21321), .ZN(n11708) );
  OR2_X1 U11739 ( .A1(n11759), .A2(n11758), .ZN(n12427) );
  OR2_X1 U11740 ( .A1(n11747), .A2(n11746), .ZN(n12424) );
  OR2_X1 U11741 ( .A1(n11651), .A2(n11650), .ZN(n12396) );
  OR2_X1 U11742 ( .A1(n11663), .A2(n11662), .ZN(n12453) );
  OR2_X1 U11743 ( .A1(n11718), .A2(n11717), .ZN(n12383) );
  NAND2_X1 U11744 ( .A1(n11191), .A2(n13634), .ZN(n13581) );
  INV_X1 U11745 ( .A(n11621), .ZN(n11191) );
  NAND2_X1 U11746 ( .A1(n21319), .A2(n11621), .ZN(n11446) );
  AND3_X1 U11747 ( .A1(n11640), .A2(n13747), .A3(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n12302) );
  NAND2_X1 U11748 ( .A1(n13443), .A2(n11396), .ZN(n11397) );
  AND2_X1 U11749 ( .A1(n11118), .A2(n14001), .ZN(n12798) );
  INV_X1 U11750 ( .A(n14003), .ZN(n11118) );
  INV_X1 U11751 ( .A(n12787), .ZN(n12811) );
  NOR2_X1 U11752 ( .A1(n16314), .A2(n11159), .ZN(n11158) );
  INV_X1 U11753 ( .A(n16313), .ZN(n11159) );
  CLKBUF_X1 U11754 ( .A(n15275), .Z(n15280) );
  INV_X1 U11755 ( .A(n14853), .ZN(n11099) );
  OR2_X1 U11756 ( .A1(n13195), .A2(n13194), .ZN(n13335) );
  INV_X1 U11757 ( .A(n11127), .ZN(n11126) );
  OAI21_X1 U11758 ( .B1(n11124), .B2(n13675), .A(n19203), .ZN(n11127) );
  INV_X1 U11759 ( .A(n19464), .ZN(n14993) );
  OR2_X1 U11760 ( .A1(n13304), .A2(n13303), .ZN(n13518) );
  OR2_X1 U11761 ( .A1(n13205), .A2(n13204), .ZN(n14831) );
  NAND2_X1 U11762 ( .A1(n13236), .A2(n12746), .ZN(n13998) );
  NAND2_X1 U11763 ( .A1(n10967), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n11374) );
  NAND2_X1 U11764 ( .A1(n10968), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(
        n11373) );
  INV_X1 U11765 ( .A(n14765), .ZN(n14764) );
  AOI21_X1 U11766 ( .B1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n21263), .A(
        n14638), .ZN(n14644) );
  INV_X1 U11767 ( .A(n14669), .ZN(n14614) );
  INV_X1 U11768 ( .A(n20809), .ZN(n14613) );
  INV_X1 U11769 ( .A(n14661), .ZN(n14616) );
  OR2_X1 U11770 ( .A1(n12332), .A2(n12334), .ZN(n12349) );
  NAND2_X1 U11771 ( .A1(n11708), .A2(n11707), .ZN(n12343) );
  INV_X1 U11772 ( .A(n12342), .ZN(n12352) );
  NAND2_X1 U11773 ( .A1(n12302), .A2(n12440), .ZN(n12341) );
  NAND2_X1 U11774 ( .A1(n11360), .A2(n11358), .ZN(n11357) );
  AOI21_X1 U11775 ( .B1(n12335), .B2(n12334), .A(n11359), .ZN(n11358) );
  NAND2_X1 U11776 ( .A1(n11361), .A2(n12336), .ZN(n11360) );
  AND2_X1 U11777 ( .A1(n21321), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n11359) );
  AOI22_X1 U11778 ( .A1(n11979), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12197), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11510) );
  AND2_X1 U11779 ( .A1(n11467), .A2(n12112), .ZN(n11466) );
  NOR2_X1 U11780 ( .A1(n15590), .A2(n11468), .ZN(n11467) );
  AOI21_X1 U11781 ( .B1(n12264), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .A(
        n11176), .ZN(n12017) );
  NAND2_X1 U11782 ( .A1(n11189), .A2(n11911), .ZN(n15085) );
  INV_X1 U11783 ( .A(n15077), .ZN(n11189) );
  AOI21_X1 U11784 ( .B1(n11962), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A(
        n11162), .ZN(n11896) );
  NOR2_X1 U11785 ( .A1(n11902), .A2(n21480), .ZN(n11906) );
  AOI21_X1 U11786 ( .B1(n12264), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A(
        n11175), .ZN(n11862) );
  NOR2_X1 U11787 ( .A1(n15574), .A2(n11291), .ZN(n11290) );
  INV_X1 U11788 ( .A(n15578), .ZN(n11291) );
  NAND2_X1 U11789 ( .A1(n15995), .A2(n11459), .ZN(n11458) );
  NAND2_X1 U11790 ( .A1(n11449), .A2(n12405), .ZN(n12414) );
  OAI21_X1 U11791 ( .B1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n13762), .A(
        n13761), .ZN(n11449) );
  OR2_X1 U11792 ( .A1(n11735), .A2(n11734), .ZN(n12411) );
  OR2_X1 U11793 ( .A1(n11682), .A2(n11681), .ZN(n12395) );
  INV_X1 U11794 ( .A(n11626), .ZN(n11627) );
  NAND2_X1 U11795 ( .A1(n13582), .A2(n11178), .ZN(n13750) );
  INV_X1 U11796 ( .A(n11179), .ZN(n11178) );
  INV_X1 U11797 ( .A(n13469), .ZN(n11571) );
  AND2_X1 U11798 ( .A1(n21905), .A2(n11699), .ZN(n14408) );
  NAND2_X1 U11799 ( .A1(n11288), .A2(n15195), .ZN(n11287) );
  NOR2_X1 U11800 ( .A1(n11289), .A2(n15171), .ZN(n11288) );
  INV_X1 U11801 ( .A(n15198), .ZN(n11289) );
  NOR2_X1 U11802 ( .A1(n15179), .A2(n15171), .ZN(n15199) );
  OR2_X1 U11803 ( .A1(n15190), .A2(n15177), .ZN(n15179) );
  NAND2_X1 U11804 ( .A1(n16114), .A2(n11485), .ZN(n13117) );
  AND2_X1 U11805 ( .A1(n11421), .A2(n16145), .ZN(n11420) );
  AND2_X1 U11806 ( .A1(n16159), .A2(n11422), .ZN(n11421) );
  INV_X1 U11807 ( .A(n16152), .ZN(n11422) );
  INV_X1 U11808 ( .A(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n11392) );
  NAND2_X1 U11809 ( .A1(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n11393) );
  OR2_X1 U11810 ( .A1(n15390), .A2(n15335), .ZN(n15447) );
  NOR2_X1 U11811 ( .A1(n16345), .A2(n11387), .ZN(n11386) );
  INV_X1 U11812 ( .A(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n11387) );
  NOR2_X1 U11813 ( .A1(n18265), .A2(n11390), .ZN(n11389) );
  INV_X1 U11814 ( .A(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n11390) );
  NAND2_X1 U11815 ( .A1(n13855), .A2(n11315), .ZN(n11314) );
  INV_X1 U11816 ( .A(n13925), .ZN(n11315) );
  NAND2_X1 U11817 ( .A1(n12807), .A2(n12785), .ZN(n14810) );
  OR2_X1 U11818 ( .A1(n12811), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12788) );
  NAND2_X1 U11819 ( .A1(n12801), .A2(n11097), .ZN(n12749) );
  NAND2_X1 U11820 ( .A1(n12800), .A2(n13498), .ZN(n11097) );
  OR2_X1 U11821 ( .A1(n15413), .A2(n15412), .ZN(n15417) );
  INV_X1 U11822 ( .A(n16199), .ZN(n11339) );
  AND2_X1 U11823 ( .A1(n18413), .A2(n15420), .ZN(n15307) );
  AND2_X1 U11824 ( .A1(n18349), .A2(n15420), .ZN(n15220) );
  NAND2_X1 U11825 ( .A1(n11416), .A2(n11110), .ZN(n15221) );
  NOR2_X1 U11826 ( .A1(n11111), .A2(n15165), .ZN(n11110) );
  INV_X1 U11827 ( .A(n11414), .ZN(n11111) );
  AOI21_X1 U11828 ( .B1(n11158), .B2(n16312), .A(n11156), .ZN(n11155) );
  INV_X1 U11829 ( .A(n16363), .ZN(n11156) );
  INV_X1 U11830 ( .A(n11158), .ZN(n11157) );
  OR2_X1 U11831 ( .A1(n11244), .A2(n16326), .ZN(n11243) );
  NAND2_X1 U11832 ( .A1(n16304), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n16305) );
  NAND2_X1 U11833 ( .A1(n11116), .A2(n18155), .ZN(n15137) );
  OR2_X1 U11834 ( .A1(n13320), .A2(n13319), .ZN(n13513) );
  OAI21_X1 U11835 ( .B1(n19605), .B2(n12758), .A(n11437), .ZN(n15000) );
  NAND2_X1 U11836 ( .A1(n19605), .A2(n14999), .ZN(n11437) );
  OAI21_X1 U11837 ( .B1(n14807), .B2(n14078), .A(n12844), .ZN(n12846) );
  AND2_X2 U11838 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n12875) );
  NAND2_X1 U11839 ( .A1(n13242), .A2(n11442), .ZN(n11441) );
  AND2_X1 U11840 ( .A1(n11021), .A2(n12754), .ZN(n11442) );
  NAND2_X1 U11841 ( .A1(n12846), .A2(n12845), .ZN(n12861) );
  AND2_X1 U11842 ( .A1(n18521), .A2(n14810), .ZN(n14822) );
  NAND2_X1 U11843 ( .A1(n11096), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11095) );
  NAND2_X1 U11844 ( .A1(n11094), .A2(n12681), .ZN(n11093) );
  AND2_X1 U11845 ( .A1(n17064), .A2(n18644), .ZN(n16667) );
  AND2_X1 U11846 ( .A1(n19323), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13213) );
  NAND2_X1 U11847 ( .A1(n13179), .A2(n13178), .ZN(n13207) );
  XNOR2_X1 U11848 ( .A(n12681), .B(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n13206) );
  AOI221_X1 U11849 ( .B1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(n13183), 
        .C1(n14054), .C2(n13183), .A(n13182), .ZN(n13489) );
  INV_X1 U11850 ( .A(n14628), .ZN(n16713) );
  INV_X1 U11851 ( .A(n20462), .ZN(n11210) );
  OR2_X1 U11852 ( .A1(n16689), .A2(n20163), .ZN(n17391) );
  NAND2_X1 U11853 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n11200) );
  NAND2_X1 U11854 ( .A1(n17701), .A2(n11004), .ZN(n17729) );
  AND2_X1 U11855 ( .A1(n20245), .A2(n11229), .ZN(n20310) );
  AND2_X1 U11856 ( .A1(n10995), .A2(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n11229) );
  INV_X1 U11857 ( .A(n17563), .ZN(n17561) );
  NAND2_X1 U11858 ( .A1(n17570), .A2(n17571), .ZN(n17600) );
  NAND2_X1 U11859 ( .A1(n17559), .A2(n17560), .ZN(n17892) );
  NAND2_X1 U11860 ( .A1(n14759), .A2(n14760), .ZN(n17570) );
  INV_X1 U11861 ( .A(n18925), .ZN(n14624) );
  NOR2_X1 U11862 ( .A1(n20673), .A2(n20674), .ZN(n14669) );
  AND2_X1 U11863 ( .A1(n14669), .A2(n20808), .ZN(n17146) );
  NAND2_X1 U11864 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n20192) );
  NAND2_X1 U11865 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n16689) );
  INV_X1 U11866 ( .A(n14609), .ZN(n11272) );
  NOR2_X1 U11867 ( .A1(n19925), .A2(n19924), .ZN(n11383) );
  NAND2_X1 U11868 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(P1_REIP_REG_22__SCAN_IN), 
        .ZN(n11377) );
  INV_X1 U11869 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n21543) );
  NAND2_X1 U11870 ( .A1(P1_REIP_REG_13__SCAN_IN), .A2(P1_REIP_REG_14__SCAN_IN), 
        .ZN(n11367) );
  INV_X1 U11871 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n21480) );
  NAND2_X1 U11872 ( .A1(n12633), .A2(n11000), .ZN(n21457) );
  NAND2_X1 U11873 ( .A1(n12633), .A2(n11381), .ZN(n21439) );
  AND2_X1 U11874 ( .A1(n13562), .A2(n13561), .ZN(n19854) );
  AND2_X1 U11875 ( .A1(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n12235), .ZN(
        n12236) );
  NAND2_X1 U11876 ( .A1(n12236), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12289) );
  NAND2_X1 U11877 ( .A1(n12178), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12234) );
  AND2_X1 U11878 ( .A1(n15761), .A2(n12291), .ZN(n12136) );
  NOR2_X1 U11879 ( .A1(n12093), .A2(n21593), .ZN(n12094) );
  NAND2_X1 U11880 ( .A1(n12060), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12093) );
  AND2_X1 U11881 ( .A1(n12058), .A2(n12057), .ZN(n15604) );
  NOR2_X1 U11882 ( .A1(n12027), .A2(n12022), .ZN(n12028) );
  NAND2_X1 U11883 ( .A1(n12028), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n12059) );
  OR2_X1 U11884 ( .A1(n11470), .A2(n15609), .ZN(n11469) );
  NOR2_X1 U11885 ( .A1(n11994), .A2(n21543), .ZN(n11995) );
  NAND2_X1 U11886 ( .A1(n11995), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12027) );
  NAND2_X1 U11887 ( .A1(n11978), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11994) );
  AND2_X1 U11888 ( .A1(n11961), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n11978) );
  NOR2_X1 U11889 ( .A1(n11953), .A2(n11924), .ZN(n11961) );
  NAND2_X1 U11890 ( .A1(n11907), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n11953) );
  AND2_X1 U11891 ( .A1(n11855), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11877) );
  OAI211_X1 U11892 ( .C1(n11822), .C2(n11847), .A(n11846), .B(n11845), .ZN(
        n14307) );
  AND2_X1 U11893 ( .A1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n11765), .ZN(
        n11817) );
  NAND2_X1 U11894 ( .A1(n13914), .A2(n13913), .ZN(n14204) );
  INV_X1 U11895 ( .A(n13778), .ZN(n11811) );
  OAI21_X1 U11896 ( .B1(n12508), .B2(n12507), .A(n12505), .ZN(n11451) );
  NOR2_X1 U11897 ( .A1(n11220), .A2(n15994), .ZN(n11218) );
  NAND2_X1 U11898 ( .A1(n15579), .A2(n11072), .ZN(n15531) );
  NAND2_X1 U11899 ( .A1(n15579), .A2(n11290), .ZN(n15871) );
  NAND2_X1 U11900 ( .A1(n15579), .A2(n15578), .ZN(n15577) );
  OR2_X1 U11901 ( .A1(n15592), .A2(n15584), .ZN(n15586) );
  NAND2_X1 U11902 ( .A1(n11150), .A2(n15881), .ZN(n15896) );
  NAND2_X1 U11903 ( .A1(n15777), .A2(n15909), .ZN(n11150) );
  NAND2_X1 U11904 ( .A1(n15605), .A2(n11297), .ZN(n11296) );
  NOR2_X1 U11905 ( .A1(n15593), .A2(n11298), .ZN(n11297) );
  NOR3_X1 U11906 ( .A1(n15612), .A2(n11301), .A3(n15611), .ZN(n15607) );
  NOR2_X1 U11907 ( .A1(n15612), .A2(n15611), .ZN(n15613) );
  OR2_X1 U11908 ( .A1(n15881), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15933) );
  NAND2_X1 U11909 ( .A1(n15995), .A2(n15784), .ZN(n15931) );
  INV_X1 U11910 ( .A(n21416), .ZN(n15967) );
  NAND2_X1 U11911 ( .A1(n15081), .A2(n15080), .ZN(n15102) );
  AND2_X1 U11912 ( .A1(n14953), .A2(n14952), .ZN(n15081) );
  AOI21_X1 U11913 ( .B1(n14906), .B2(n14907), .A(n12458), .ZN(n14923) );
  INV_X1 U11914 ( .A(n14463), .ZN(n11292) );
  AND2_X1 U11915 ( .A1(n12564), .A2(n12563), .ZN(n14498) );
  NAND2_X1 U11916 ( .A1(n11293), .A2(n11294), .ZN(n14464) );
  INV_X1 U11917 ( .A(n14099), .ZN(n12548) );
  INV_X1 U11918 ( .A(n14100), .ZN(n12549) );
  NOR2_X1 U11919 ( .A1(n13745), .A2(n13744), .ZN(n15987) );
  AND2_X1 U11920 ( .A1(n13768), .A2(n13767), .ZN(n13875) );
  INV_X1 U11921 ( .A(n15903), .ZN(n15982) );
  INV_X1 U11922 ( .A(n11793), .ZN(n11146) );
  INV_X1 U11923 ( .A(n11184), .ZN(n11183) );
  NAND2_X1 U11924 ( .A1(n11725), .A2(n11724), .ZN(n13978) );
  NOR2_X1 U11925 ( .A1(n12511), .A2(n14298), .ZN(n16744) );
  OR2_X1 U11926 ( .A1(n12407), .A2(n11056), .ZN(n21836) );
  INV_X1 U11927 ( .A(n11617), .ZN(n14182) );
  INV_X1 U11928 ( .A(n13735), .ZN(n13593) );
  NAND2_X1 U11929 ( .A1(n15411), .A2(n15410), .ZN(n15413) );
  OR2_X1 U11930 ( .A1(n15411), .A2(n15405), .ZN(n18441) );
  AND2_X1 U11931 ( .A1(n11352), .A2(n11351), .ZN(n11350) );
  INV_X1 U11932 ( .A(n15351), .ZN(n11351) );
  NAND2_X1 U11933 ( .A1(n16366), .A2(n11385), .ZN(n16322) );
  AND2_X1 U11934 ( .A1(n10996), .A2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n11385) );
  AND2_X1 U11935 ( .A1(n13413), .A2(n13412), .ZN(n16238) );
  NOR2_X1 U11936 ( .A1(n15179), .A2(n11286), .ZN(n15201) );
  INV_X1 U11937 ( .A(n11288), .ZN(n11286) );
  NOR2_X1 U11938 ( .A1(n16367), .A2(n17049), .ZN(n16366) );
  AND2_X1 U11939 ( .A1(n15182), .A2(n15181), .ZN(n15188) );
  NAND2_X1 U11940 ( .A1(n15188), .A2(n15187), .ZN(n15190) );
  NAND2_X1 U11941 ( .A1(n15143), .A2(n10988), .ZN(n15151) );
  NAND2_X1 U11942 ( .A1(n15143), .A2(n15142), .ZN(n15419) );
  NOR2_X1 U11943 ( .A1(n15016), .A2(n15015), .ZN(n15019) );
  NAND2_X1 U11944 ( .A1(n16163), .A2(n11324), .ZN(n16148) );
  OR2_X1 U11945 ( .A1(n12929), .A2(n12928), .ZN(n13397) );
  OR2_X1 U11946 ( .A1(n12909), .A2(n12908), .ZN(n13391) );
  NAND2_X1 U11947 ( .A1(n11123), .A2(n11122), .ZN(n16096) );
  NAND2_X1 U11948 ( .A1(n16478), .A2(n11352), .ZN(n15352) );
  NAND2_X1 U11949 ( .A1(n16478), .A2(n16227), .ZN(n16228) );
  CLKBUF_X1 U11950 ( .A(n16131), .Z(n16139) );
  NAND2_X1 U11951 ( .A1(n16160), .A2(n11420), .ZN(n16144) );
  NOR2_X1 U11952 ( .A1(n11008), .A2(n16238), .ZN(n16477) );
  AND2_X1 U11953 ( .A1(n16477), .A2(n16476), .ZN(n16478) );
  INV_X1 U11954 ( .A(n14939), .ZN(n11135) );
  NOR2_X1 U11955 ( .A1(n11335), .A2(n11332), .ZN(n11331) );
  NAND2_X1 U11956 ( .A1(n15042), .A2(n11333), .ZN(n11332) );
  INV_X1 U11957 ( .A(n13228), .ZN(n12760) );
  AND2_X1 U11958 ( .A1(n13641), .A2(n21735), .ZN(n17095) );
  NOR2_X1 U11959 ( .A1(n15447), .A2(n11391), .ZN(n16263) );
  OR3_X1 U11960 ( .A1(n11393), .A2(n11392), .A3(n16264), .ZN(n11391) );
  NOR2_X1 U11961 ( .A1(n15447), .A2(n11393), .ZN(n16283) );
  NAND2_X1 U11962 ( .A1(n15391), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15390) );
  AND2_X1 U11963 ( .A1(n15364), .A2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15391) );
  NOR2_X1 U11964 ( .A1(n16322), .A2(n15288), .ZN(n15364) );
  AND2_X1 U11965 ( .A1(n16163), .A2(n11058), .ZN(n16137) );
  INV_X1 U11966 ( .A(n16136), .ZN(n11323) );
  AND2_X1 U11967 ( .A1(n16137), .A2(n15241), .ZN(n15349) );
  NAND2_X1 U11968 ( .A1(n16366), .A2(n10996), .ZN(n16334) );
  NAND2_X1 U11969 ( .A1(n16163), .A2(n16155), .ZN(n16154) );
  INV_X1 U11970 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n16345) );
  NAND2_X1 U11971 ( .A1(n16366), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n16357) );
  NAND2_X1 U11972 ( .A1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n11006), .ZN(
        n11244) );
  AND2_X1 U11973 ( .A1(n17025), .A2(n11388), .ZN(n17050) );
  AND2_X1 U11974 ( .A1(n10997), .A2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n11388) );
  NAND2_X1 U11975 ( .A1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n17050), .ZN(
        n17049) );
  AND2_X1 U11976 ( .A1(n14220), .A2(n10989), .ZN(n14801) );
  NAND2_X1 U11977 ( .A1(n17025), .A2(n10997), .ZN(n17031) );
  NAND2_X1 U11978 ( .A1(n17025), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n17024) );
  NOR2_X1 U11979 ( .A1(n13857), .A2(n11314), .ZN(n14287) );
  NOR2_X1 U11980 ( .A1(n17023), .A2(n17014), .ZN(n17025) );
  NAND2_X1 U11981 ( .A1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n17008), .ZN(
        n17014) );
  NAND2_X1 U11982 ( .A1(n11311), .A2(n13855), .ZN(n13926) );
  NOR2_X1 U11983 ( .A1(n17007), .A2(n17000), .ZN(n17008) );
  NAND2_X1 U11984 ( .A1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n16979), .ZN(
        n16978) );
  NAND2_X1 U11985 ( .A1(n14865), .A2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n14900) );
  NOR2_X1 U11986 ( .A1(n14900), .A2(n18124), .ZN(n16979) );
  NAND2_X1 U11987 ( .A1(n11131), .A2(n12820), .ZN(n11128) );
  AND2_X1 U11988 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n14865) );
  INV_X1 U11989 ( .A(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n16041) );
  NAND2_X1 U11990 ( .A1(n10985), .A2(n11105), .ZN(n11104) );
  INV_X1 U11991 ( .A(n16256), .ZN(n11105) );
  NAND2_X1 U11992 ( .A1(n15407), .A2(n16427), .ZN(n11405) );
  AND3_X1 U11993 ( .A1(n18472), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n15420), .ZN(n16256) );
  NAND2_X1 U11994 ( .A1(n16107), .A2(n11069), .ZN(n16090) );
  INV_X1 U11995 ( .A(n16092), .ZN(n11326) );
  AND2_X1 U11996 ( .A1(n18458), .A2(n15420), .ZN(n16273) );
  AND2_X1 U11997 ( .A1(n15383), .A2(n11337), .ZN(n16187) );
  AND2_X1 U11998 ( .A1(n11066), .A2(n11338), .ZN(n11337) );
  INV_X1 U11999 ( .A(n16186), .ZN(n11338) );
  NAND2_X1 U12000 ( .A1(n15383), .A2(n11066), .ZN(n16196) );
  NAND2_X1 U12001 ( .A1(n16107), .A2(n11327), .ZN(n16099) );
  NOR2_X1 U12002 ( .A1(n11408), .A2(n15345), .ZN(n11407) );
  NAND2_X1 U12003 ( .A1(n11413), .A2(n11409), .ZN(n11115) );
  AND2_X1 U12004 ( .A1(n15343), .A2(n11411), .ZN(n11408) );
  AND2_X1 U12005 ( .A1(n11428), .A2(n15321), .ZN(n11091) );
  NAND2_X1 U12006 ( .A1(n11413), .A2(n11412), .ZN(n11406) );
  INV_X1 U12007 ( .A(n11411), .ZN(n11410) );
  AND2_X1 U12008 ( .A1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n15258), .ZN(
        n16474) );
  OR2_X1 U12009 ( .A1(n18330), .A2(n15214), .ZN(n16341) );
  NOR2_X1 U12010 ( .A1(n16162), .A2(n16161), .ZN(n16163) );
  NAND2_X1 U12011 ( .A1(n11152), .A2(n11155), .ZN(n16354) );
  OR2_X1 U12012 ( .A1(n16522), .A2(n11157), .ZN(n11152) );
  OR2_X1 U12013 ( .A1(n15208), .A2(n15207), .ZN(n16352) );
  OR2_X1 U12014 ( .A1(n15070), .A2(n15071), .ZN(n16162) );
  AND2_X1 U12015 ( .A1(n18547), .A2(n15257), .ZN(n16514) );
  AND2_X1 U12016 ( .A1(n10989), .A2(n14800), .ZN(n11319) );
  OR2_X1 U12017 ( .A1(n14946), .A2(n14947), .ZN(n15070) );
  AND2_X1 U12018 ( .A1(n14450), .A2(n14449), .ZN(n14791) );
  NAND2_X1 U12019 ( .A1(n16307), .A2(n16306), .ZN(n11253) );
  INV_X1 U12020 ( .A(n14289), .ZN(n14220) );
  NOR2_X1 U12021 ( .A1(n13721), .A2(n16590), .ZN(n13863) );
  NAND2_X1 U12022 ( .A1(n16995), .A2(n16996), .ZN(n11430) );
  AND3_X1 U12023 ( .A1(n13388), .A2(n13387), .A3(n13386), .ZN(n13686) );
  AND2_X1 U12024 ( .A1(n11342), .A2(n11340), .ZN(n13723) );
  NOR2_X1 U12025 ( .A1(n13888), .A2(n11027), .ZN(n13880) );
  NOR2_X1 U12026 ( .A1(n11027), .A2(n11308), .ZN(n11307) );
  INV_X1 U12027 ( .A(n13879), .ZN(n11308) );
  NAND2_X1 U12028 ( .A1(n11236), .A2(n10991), .ZN(n11439) );
  NAND2_X1 U12029 ( .A1(n11334), .A2(n11333), .ZN(n11330) );
  NAND2_X1 U12030 ( .A1(n11306), .A2(n13827), .ZN(n13890) );
  NAND2_X1 U12031 ( .A1(n15049), .A2(n15030), .ZN(n18608) );
  OAI211_X1 U12032 ( .C1(n13507), .C2(n13408), .A(n13321), .B(n13291), .ZN(
        n13669) );
  AND2_X1 U12033 ( .A1(n13669), .A2(n13670), .ZN(n13668) );
  OAI21_X1 U12034 ( .B1(n12846), .B2(n12845), .A(n12861), .ZN(n13666) );
  AND2_X1 U12035 ( .A1(n14011), .A2(n14010), .ZN(n15032) );
  INV_X1 U12036 ( .A(n14817), .ZN(n14806) );
  INV_X1 U12037 ( .A(n14818), .ZN(n11250) );
  NOR3_X2 U12038 ( .A1(n16679), .A2(n21695), .A3(n19252), .ZN(n19671) );
  NOR3_X2 U12039 ( .A1(n21695), .A2(n16678), .A3(n19252), .ZN(n19672) );
  NAND2_X1 U12040 ( .A1(n19168), .A2(n19151), .ZN(n19278) );
  NAND2_X1 U12041 ( .A1(n19168), .A2(n19147), .ZN(n19293) );
  INV_X1 U12042 ( .A(n19671), .ZN(n19679) );
  INV_X1 U12043 ( .A(n19672), .ZN(n19681) );
  INV_X1 U12044 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n14054) );
  NOR2_X1 U12045 ( .A1(n20171), .A2(n20166), .ZN(n20609) );
  NOR2_X1 U12046 ( .A1(n16713), .A2(n20613), .ZN(n21249) );
  CLKBUF_X1 U12047 ( .A(n20507), .Z(n20530) );
  NOR2_X1 U12048 ( .A1(n16689), .A2(n14524), .ZN(n14544) );
  NOR2_X1 U12049 ( .A1(n14524), .A2(n14522), .ZN(n14572) );
  NAND2_X1 U12050 ( .A1(n20662), .A2(n11483), .ZN(n20641) );
  NOR2_X1 U12051 ( .A1(n11370), .A2(n11369), .ZN(n11368) );
  INV_X1 U12052 ( .A(n20615), .ZN(n20686) );
  NOR2_X1 U12053 ( .A1(n14680), .A2(n14625), .ZN(n20111) );
  NOR2_X1 U12054 ( .A1(n17797), .A2(n20559), .ZN(n17769) );
  NOR2_X1 U12055 ( .A1(n17797), .A2(n11200), .ZN(n17785) );
  NAND2_X1 U12056 ( .A1(n17731), .A2(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n17797) );
  INV_X1 U12057 ( .A(n17729), .ZN(n17731) );
  NOR2_X1 U12058 ( .A1(n21125), .A2(n21032), .ZN(n17735) );
  NAND2_X1 U12059 ( .A1(n11224), .A2(n11073), .ZN(n11223) );
  INV_X1 U12060 ( .A(n11225), .ZN(n11224) );
  NOR2_X1 U12061 ( .A1(n17574), .A2(n11225), .ZN(n17649) );
  NOR3_X1 U12062 ( .A1(n17574), .A2(n11228), .A3(n20413), .ZN(n17672) );
  NOR2_X1 U12063 ( .A1(n17574), .A2(n20413), .ZN(n17588) );
  NAND2_X1 U12064 ( .A1(n17810), .A2(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n17574) );
  NOR2_X1 U12065 ( .A1(n17598), .A2(n17612), .ZN(n17810) );
  NAND2_X1 U12066 ( .A1(n17821), .A2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n17598) );
  NAND2_X1 U12067 ( .A1(n20310), .A2(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n17623) );
  NAND2_X1 U12068 ( .A1(n20245), .A2(n10995), .ZN(n17853) );
  XNOR2_X1 U12069 ( .A(n17557), .B(n11305), .ZN(n14778) );
  INV_X1 U12070 ( .A(n17558), .ZN(n11305) );
  INV_X1 U12071 ( .A(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n17928) );
  NOR2_X1 U12072 ( .A1(n14680), .A2(n21315), .ZN(n17577) );
  INV_X1 U12073 ( .A(n21119), .ZN(n17792) );
  INV_X1 U12074 ( .A(n17737), .ZN(n11259) );
  INV_X1 U12075 ( .A(n11260), .ZN(n17753) );
  INV_X1 U12076 ( .A(n17721), .ZN(n11256) );
  NAND2_X1 U12077 ( .A1(n17709), .A2(n17710), .ZN(n17722) );
  NOR2_X1 U12078 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17722), .ZN(
        n17721) );
  NAND2_X1 U12079 ( .A1(n17824), .A2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n21174) );
  AND2_X1 U12080 ( .A1(n20950), .A2(n20975), .ZN(n17828) );
  NOR2_X1 U12081 ( .A1(n20974), .A2(n17825), .ZN(n17824) );
  INV_X1 U12082 ( .A(n17576), .ZN(n20952) );
  INV_X1 U12083 ( .A(n21184), .ZN(n21229) );
  NAND2_X1 U12084 ( .A1(n17920), .A2(n14775), .ZN(n17910) );
  NAND2_X1 U12085 ( .A1(n17910), .A2(n17911), .ZN(n17909) );
  NAND2_X1 U12086 ( .A1(n17926), .A2(n17927), .ZN(n17925) );
  NAND2_X1 U12087 ( .A1(n17945), .A2(n14771), .ZN(n17934) );
  NAND2_X1 U12088 ( .A1(n17934), .A2(n17935), .ZN(n17933) );
  OAI21_X1 U12089 ( .B1(n14650), .B2(n14654), .A(n14655), .ZN(n21280) );
  OAI211_X1 U12090 ( .C1(n14657), .C2(n14656), .A(n14655), .B(n14654), .ZN(
        n21255) );
  NOR2_X1 U12091 ( .A1(n21141), .A2(n14680), .ZN(n21104) );
  INV_X1 U12092 ( .A(n21147), .ZN(n21254) );
  AND2_X1 U12093 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n20180) );
  INV_X1 U12094 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n21262) );
  NOR2_X1 U12095 ( .A1(n14567), .A2(n14566), .ZN(n18885) );
  NOR2_X2 U12096 ( .A1(n14600), .A2(n14599), .ZN(n18844) );
  NOR2_X1 U12097 ( .A1(n14578), .A2(n14577), .ZN(n18804) );
  NAND2_X1 U12098 ( .A1(n21309), .A2(n18684), .ZN(n19010) );
  INV_X1 U12099 ( .A(n14622), .ZN(n20674) );
  OAI22_X1 U12100 ( .A1(n21255), .A2(n21147), .B1(n17566), .B2(n21251), .ZN(
        n21257) );
  NAND2_X2 U12101 ( .A1(n12370), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n14376)
         );
  NAND2_X1 U12102 ( .A1(n15550), .A2(n11383), .ZN(n15511) );
  AND2_X1 U12103 ( .A1(n21654), .A2(P1_REIP_REG_27__SCAN_IN), .ZN(n15550) );
  AND2_X1 U12104 ( .A1(n21638), .A2(P1_REIP_REG_26__SCAN_IN), .ZN(n21654) );
  NAND2_X1 U12105 ( .A1(P1_REIP_REG_23__SCAN_IN), .A2(P1_REIP_REG_24__SCAN_IN), 
        .ZN(n11376) );
  INV_X1 U12106 ( .A(n21639), .ZN(n21523) );
  NOR3_X1 U12107 ( .A1(n21600), .A2(n11377), .A3(n19913), .ZN(n21617) );
  NAND2_X1 U12108 ( .A1(n21587), .A2(P1_REIP_REG_20__SCAN_IN), .ZN(n21600) );
  NOR2_X1 U12109 ( .A1(n21574), .A2(n21582), .ZN(n21587) );
  INV_X1 U12110 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n21573) );
  NAND2_X1 U12111 ( .A1(P1_REIP_REG_15__SCAN_IN), .A2(P1_REIP_REG_16__SCAN_IN), 
        .ZN(n11365) );
  NOR3_X1 U12112 ( .A1(n21532), .A2(n11367), .A3(n19904), .ZN(n21555) );
  NOR2_X1 U12113 ( .A1(n21532), .A2(n21522), .ZN(n21536) );
  NOR2_X1 U12114 ( .A1(n21507), .A2(n21509), .ZN(n21515) );
  NAND2_X1 U12115 ( .A1(n21422), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n21636) );
  INV_X1 U12116 ( .A(n21626), .ZN(n21640) );
  AND2_X1 U12117 ( .A1(n12638), .A2(n12637), .ZN(n21626) );
  AND2_X1 U12118 ( .A1(n13952), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13953) );
  NAND2_X1 U12119 ( .A1(n21648), .A2(n11070), .ZN(n21449) );
  INV_X1 U12120 ( .A(n21642), .ZN(n21627) );
  INV_X1 U12121 ( .A(n21636), .ZN(n21645) );
  INV_X1 U12122 ( .A(n15628), .ZN(n19962) );
  OAI21_X2 U12123 ( .B1(n13735), .B2(n13661), .A(n13660), .ZN(n19969) );
  INV_X1 U12124 ( .A(n19961), .ZN(n19965) );
  OR2_X1 U12125 ( .A1(n12379), .A2(n12380), .ZN(n12381) );
  INV_X1 U12126 ( .A(n15689), .ZN(n15682) );
  NOR2_X1 U12127 ( .A1(n15707), .A2(n13635), .ZN(n15709) );
  NAND2_X2 U12128 ( .A1(n12359), .A2(n12358), .ZN(n15703) );
  NAND2_X1 U12129 ( .A1(n13606), .A2(n20029), .ZN(n12359) );
  INV_X1 U12130 ( .A(n15709), .ZN(n15701) );
  OR2_X1 U12131 ( .A1(n15539), .A2(n15540), .ZN(n15541) );
  OAI21_X1 U12132 ( .B1(n15572), .B2(n11489), .A(n10982), .ZN(n21630) );
  NAND2_X1 U12133 ( .A1(n11145), .A2(n12477), .ZN(n12479) );
  NAND2_X1 U12134 ( .A1(n12476), .A2(n12475), .ZN(n15742) );
  AND2_X1 U12135 ( .A1(n15747), .A2(n15723), .ZN(n12475) );
  NOR2_X1 U12136 ( .A1(n11452), .A2(n11455), .ZN(n14469) );
  INV_X1 U12137 ( .A(n11454), .ZN(n11452) );
  NAND2_X1 U12138 ( .A1(n12422), .A2(n12421), .ZN(n14314) );
  NAND2_X1 U12139 ( .A1(n13753), .A2(n13752), .ZN(n21352) );
  INV_X1 U12140 ( .A(n21353), .ZN(n21410) );
  INV_X1 U12141 ( .A(n21352), .ZN(n21409) );
  INV_X1 U12142 ( .A(n21683), .ZN(n16010) );
  NAND2_X1 U12143 ( .A1(n21889), .A2(n21766), .ZN(n22134) );
  INV_X1 U12144 ( .A(n21806), .ZN(n22156) );
  NOR2_X1 U12145 ( .A1(n14158), .A2(n21884), .ZN(n22161) );
  OAI211_X1 U12146 ( .C1(n22167), .C2(n21868), .A(n21829), .B(n21852), .ZN(
        n22170) );
  NOR2_X2 U12147 ( .A1(n21836), .A2(n21884), .ZN(n22181) );
  INV_X1 U12148 ( .A(n22189), .ZN(n14269) );
  OAI21_X1 U12149 ( .B1(n21873), .B2(n21872), .A(n21871), .ZN(n22190) );
  AOI22_X1 U12150 ( .A1(n21863), .A2(n21872), .B1(n21862), .B2(n21861), .ZN(
        n22194) );
  OAI211_X1 U12151 ( .C1(n22201), .C2(n21899), .A(n21898), .B(n21897), .ZN(
        n22205) );
  NOR2_X1 U12152 ( .A1(n21771), .A2(n15690), .ZN(n21914) );
  NOR2_X1 U12153 ( .A1(n21771), .A2(n14344), .ZN(n21954) );
  NOR2_X1 U12154 ( .A1(n21771), .A2(n15677), .ZN(n21989) );
  NOR2_X1 U12155 ( .A1(n21771), .A2(n14334), .ZN(n22023) );
  NOR2_X1 U12156 ( .A1(n21771), .A2(n15668), .ZN(n22058) );
  NOR2_X1 U12157 ( .A1(n21771), .A2(n14367), .ZN(n22094) );
  NOR2_X1 U12158 ( .A1(n21771), .A2(n15660), .ZN(n22128) );
  NOR2_X1 U12159 ( .A1(n21771), .A2(n14787), .ZN(n22211) );
  NAND2_X1 U12160 ( .A1(n16766), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n21689) );
  NOR2_X1 U12161 ( .A1(n13593), .A2(n21868), .ZN(n21683) );
  INV_X1 U12162 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n16772) );
  INV_X2 U12163 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n21910) );
  INV_X1 U12164 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n21725) );
  AND3_X1 U12165 ( .A1(n16719), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(
        P2_STATE2_REG_2__SCAN_IN), .ZN(n18099) );
  INV_X1 U12166 ( .A(n16412), .ZN(n18475) );
  NAND2_X1 U12167 ( .A1(n14450), .A2(n11355), .ZN(n16524) );
  OR2_X1 U12168 ( .A1(n18095), .A2(n16024), .ZN(n18502) );
  AND2_X1 U12169 ( .A1(n15143), .A2(n10990), .ZN(n15153) );
  NOR2_X1 U12170 ( .A1(n16029), .A2(n16028), .ZN(n18457) );
  INV_X1 U12171 ( .A(n18453), .ZN(n18510) );
  INV_X1 U12172 ( .A(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n18167) );
  INV_X1 U12173 ( .A(n18507), .ZN(n18486) );
  INV_X1 U12174 ( .A(n18634), .ZN(n18493) );
  INV_X1 U12175 ( .A(n18499), .ZN(n18509) );
  OR2_X1 U12176 ( .A1(n19670), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n18499) );
  INV_X1 U12177 ( .A(n19147), .ZN(n19151) );
  NAND2_X1 U12178 ( .A1(n13839), .A2(n11425), .ZN(n14285) );
  OR2_X1 U12179 ( .A1(n12897), .A2(n12896), .ZN(n13928) );
  OR2_X1 U12180 ( .A1(n12881), .A2(n12880), .ZN(n13842) );
  NAND2_X1 U12181 ( .A1(n13839), .A2(n12883), .ZN(n13931) );
  AOI21_X1 U12182 ( .B1(n16054), .B2(n16053), .A(n16052), .ZN(n16078) );
  NAND2_X1 U12183 ( .A1(n16684), .A2(n11124), .ZN(n13251) );
  NAND2_X1 U12184 ( .A1(n19401), .A2(n11080), .ZN(n19403) );
  INV_X1 U12185 ( .A(n19658), .ZN(n19548) );
  NAND2_X1 U12186 ( .A1(n19401), .A2(n13233), .ZN(n19658) );
  INV_X2 U12188 ( .A(n16026), .ZN(n19667) );
  AND2_X1 U12189 ( .A1(n18090), .A2(n21729), .ZN(n13448) );
  OR2_X1 U12190 ( .A1(n17033), .A2(n11244), .ZN(n16370) );
  INV_X1 U12191 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n17007) );
  INV_X1 U12192 ( .A(n17000), .ZN(n16986) );
  INV_X1 U12193 ( .A(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n18124) );
  INV_X1 U12194 ( .A(n17058), .ZN(n17039) );
  INV_X1 U12195 ( .A(n17047), .ZN(n17042) );
  INV_X1 U12196 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n18120) );
  AND2_X1 U12197 ( .A1(n17022), .A2(n16718), .ZN(n17019) );
  INV_X1 U12198 ( .A(n17022), .ZN(n17052) );
  INV_X1 U12199 ( .A(n17019), .ZN(n17062) );
  NAND2_X1 U12200 ( .A1(n15491), .A2(n15490), .ZN(n15492) );
  NAND2_X1 U12201 ( .A1(n18491), .A2(n18622), .ZN(n15491) );
  XNOR2_X1 U12202 ( .A(n16082), .B(n15481), .ZN(n18498) );
  OAI21_X1 U12203 ( .B1(n16298), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n16297), .ZN(n16454) );
  NOR2_X1 U12204 ( .A1(n16455), .A2(n11089), .ZN(n11088) );
  NOR2_X1 U12205 ( .A1(n16294), .A2(n18605), .ZN(n11089) );
  INV_X1 U12206 ( .A(n11413), .ZN(n15299) );
  INV_X1 U12207 ( .A(n16321), .ZN(n18363) );
  NAND2_X1 U12208 ( .A1(n16328), .A2(n16327), .ZN(n16463) );
  XNOR2_X1 U12209 ( .A(n11160), .B(n11047), .ZN(n16465) );
  NAND2_X1 U12210 ( .A1(n16466), .A2(n16320), .ZN(n11160) );
  NAND2_X1 U12211 ( .A1(n16520), .A2(n16313), .ZN(n16365) );
  XNOR2_X1 U12212 ( .A(n16304), .B(n16570), .ZN(n17015) );
  AND2_X1 U12213 ( .A1(n11418), .A2(n11044), .ZN(n16585) );
  NAND2_X1 U12214 ( .A1(n11418), .A2(n15149), .ZN(n16612) );
  NAND2_X1 U12215 ( .A1(n11343), .A2(n11037), .ZN(n13685) );
  OR2_X1 U12216 ( .A1(n13682), .A2(n13681), .ZN(n11343) );
  NAND2_X1 U12217 ( .A1(n11239), .A2(n11238), .ZN(n15267) );
  NAND2_X1 U12218 ( .A1(n15266), .A2(n15020), .ZN(n11239) );
  OR2_X1 U12219 ( .A1(n15266), .A2(n15020), .ZN(n11238) );
  INV_X1 U12220 ( .A(n18108), .ZN(n18521) );
  INV_X1 U12221 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19296) );
  INV_X1 U12222 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19200) );
  NOR2_X1 U12223 ( .A1(n13329), .A2(n13328), .ZN(n14138) );
  OAI21_X1 U12224 ( .B1(n18108), .B2(n14078), .A(n12850), .ZN(n16645) );
  INV_X1 U12225 ( .A(n19219), .ZN(n17077) );
  OAI21_X1 U12226 ( .B1(n16676), .B2(n16675), .A(n16674), .ZN(n19781) );
  NOR2_X1 U12227 ( .A1(n19315), .A2(n19293), .ZN(n19494) );
  OAI22_X1 U12228 ( .A1(n19290), .A2(n19287), .B1(n19286), .B2(n19285), .ZN(
        n19752) );
  OAI21_X1 U12229 ( .B1(n19274), .B2(n19273), .A(n19272), .ZN(n19744) );
  AOI211_X1 U12230 ( .C1(P2_STATE2_REG_2__SCAN_IN), .C2(n11394), .A(n19233), 
        .B(P2_STATE2_REG_3__SCAN_IN), .ZN(n19234) );
  INV_X1 U12231 ( .A(n19235), .ZN(n11394) );
  OAI21_X1 U12232 ( .B1(n19238), .B2(n19237), .A(n19236), .ZN(n19725) );
  OAI22_X1 U12233 ( .A1(n19210), .A2(n19224), .B1(n19209), .B2(n19208), .ZN(
        n19713) );
  INV_X1 U12234 ( .A(n19701), .ZN(n19698) );
  INV_X1 U12235 ( .A(n19591), .ZN(n19596) );
  INV_X1 U12236 ( .A(n19540), .ZN(n19542) );
  INV_X1 U12237 ( .A(n19431), .ZN(n19449) );
  AND2_X1 U12238 ( .A1(n19160), .A2(n19159), .ZN(n19691) );
  OAI22_X1 U12239 ( .A1(n20091), .A2(n19681), .B1(n18660), .B2(n19679), .ZN(
        n19537) );
  INV_X1 U12240 ( .A(n19500), .ZN(n19503) );
  INV_X1 U12241 ( .A(n19486), .ZN(n19502) );
  OAI22_X1 U12242 ( .A1(n20095), .A2(n19681), .B1(n18657), .B2(n19679), .ZN(
        n19437) );
  INV_X1 U12243 ( .A(n19562), .ZN(n19784) );
  OR2_X1 U12244 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(n21728), .ZN(n17143) );
  NOR2_X1 U12245 ( .A1(n20609), .A2(n17149), .ZN(n20104) );
  NOR2_X1 U12246 ( .A1(n21249), .A2(n20112), .ZN(n20165) );
  AND2_X1 U12247 ( .A1(n14667), .A2(n14625), .ZN(n21281) );
  NAND2_X1 U12248 ( .A1(n21305), .A2(n21250), .ZN(n20112) );
  NAND2_X1 U12249 ( .A1(n21257), .A2(n21305), .ZN(n21315) );
  NAND2_X1 U12250 ( .A1(n11195), .A2(n11194), .ZN(n20591) );
  AOI21_X1 U12251 ( .B1(n11196), .B2(n20391), .A(n20391), .ZN(n11194) );
  NAND2_X1 U12252 ( .A1(n11203), .A2(n11202), .ZN(n20535) );
  AOI21_X1 U12253 ( .B1(n11204), .B2(n20391), .A(n20391), .ZN(n11202) );
  NAND2_X1 U12254 ( .A1(n20460), .A2(n20577), .ZN(n20461) );
  AND2_X1 U12255 ( .A1(n20245), .A2(n11230), .ZN(n17866) );
  NOR2_X1 U12256 ( .A1(n21293), .A2(n20391), .ZN(n20593) );
  INV_X1 U12257 ( .A(n20554), .ZN(n20603) );
  NOR2_X1 U12258 ( .A1(n20488), .A2(n17439), .ZN(n17444) );
  INV_X1 U12259 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n17523) );
  INV_X1 U12260 ( .A(n17525), .ZN(n17524) );
  NOR2_X2 U12261 ( .A1(n20719), .A2(n20720), .ZN(n20743) );
  INV_X1 U12262 ( .A(n20748), .ZN(n20712) );
  NOR2_X1 U12263 ( .A1(n20753), .A2(n20711), .ZN(n20749) );
  NAND2_X1 U12264 ( .A1(n20749), .A2(P3_EAX_REG_24__SCAN_IN), .ZN(n20748) );
  NOR3_X1 U12265 ( .A1(n20711), .A2(n20760), .A3(n20672), .ZN(n20703) );
  NOR2_X2 U12266 ( .A1(n17554), .A2(n17553), .ZN(n21106) );
  NOR2_X1 U12267 ( .A1(n14703), .A2(n14702), .ZN(n20646) );
  NOR2_X1 U12268 ( .A1(n14713), .A2(n14712), .ZN(n20661) );
  NOR2_X1 U12269 ( .A1(n11266), .A2(n11263), .ZN(n11262) );
  INV_X1 U12270 ( .A(n20781), .ZN(n20789) );
  INV_X1 U12271 ( .A(n20656), .ZN(n20790) );
  NOR2_X2 U12272 ( .A1(n20113), .A2(n20112), .ZN(n20152) );
  XNOR2_X1 U12273 ( .A(n11321), .B(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n21092) );
  NAND2_X1 U12274 ( .A1(n21108), .A2(n11322), .ZN(n11321) );
  INV_X1 U12275 ( .A(n21089), .ZN(n11322) );
  NAND2_X1 U12276 ( .A1(n17701), .A2(n11001), .ZN(n17756) );
  NAND2_X1 U12277 ( .A1(n20858), .A2(n21030), .ZN(n21125) );
  OR2_X1 U12278 ( .A1(n21172), .A2(n20994), .ZN(n20990) );
  INV_X1 U12279 ( .A(n17971), .ZN(n17840) );
  NOR2_X1 U12280 ( .A1(n17623), .A2(n17635), .ZN(n17821) );
  INV_X1 U12281 ( .A(n10962), .ZN(n17809) );
  OR2_X1 U12282 ( .A1(n17971), .A2(n20952), .ZN(n11277) );
  INV_X1 U12283 ( .A(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n20264) );
  NAND2_X1 U12284 ( .A1(n20245), .A2(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n17880) );
  INV_X1 U12285 ( .A(n17829), .ZN(n17885) );
  NOR2_X2 U12286 ( .A1(n21106), .A2(n17970), .ZN(n17886) );
  NOR2_X1 U12287 ( .A1(n17903), .A2(n20233), .ZN(n20245) );
  NAND2_X1 U12288 ( .A1(n17913), .A2(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n17903) );
  INV_X1 U12289 ( .A(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n20233) );
  NOR2_X1 U12290 ( .A1(n17923), .A2(n17928), .ZN(n17913) );
  NAND2_X1 U12291 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17923) );
  INV_X1 U12292 ( .A(n17961), .ZN(n17952) );
  NAND2_X1 U12293 ( .A1(n17760), .A2(n17809), .ZN(n17961) );
  OAI21_X1 U12294 ( .B1(n20108), .B2(P3_STATE2_REG_0__SCAN_IN), .A(n21315), 
        .ZN(n17966) );
  INV_X1 U12295 ( .A(n21108), .ZN(n21061) );
  NOR2_X1 U12296 ( .A1(n14637), .A2(n20836), .ZN(n21184) );
  NAND2_X1 U12297 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n17828), .ZN(
        n20994) );
  AOI21_X1 U12298 ( .B1(n14635), .B2(n14637), .A(n20828), .ZN(n21006) );
  AND2_X1 U12299 ( .A1(n21219), .A2(n11276), .ZN(n21222) );
  INV_X1 U12300 ( .A(n21219), .ZN(n21237) );
  NOR2_X1 U12301 ( .A1(n20968), .A2(n21234), .ZN(n21242) );
  INV_X1 U12302 ( .A(n21149), .ZN(n21177) );
  INV_X1 U12303 ( .A(n21141), .ZN(n21201) );
  INV_X1 U12304 ( .A(n21104), .ZN(n21251) );
  NAND2_X1 U12305 ( .A1(n14680), .A2(n21201), .ZN(n21147) );
  NAND2_X1 U12306 ( .A1(n21117), .A2(n21104), .ZN(n20929) );
  NAND2_X1 U12307 ( .A1(n21117), .A2(n21254), .ZN(n21048) );
  NOR2_X1 U12308 ( .A1(n14679), .A2(n16698), .ZN(n21219) );
  INV_X1 U12309 ( .A(n21117), .ZN(n21234) );
  NOR3_X1 U12310 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(P3_STATE2_REG_3__SCAN_IN), .A3(n21700), .ZN(n18703) );
  INV_X1 U12311 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n16711) );
  AOI211_X1 U12312 ( .C1(n21305), .C2(n21269), .A(n18685), .B(n16697), .ZN(
        n20843) );
  INV_X1 U12313 ( .A(n20843), .ZN(n20841) );
  INV_X1 U12314 ( .A(n21310), .ZN(n21305) );
  INV_X1 U12315 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n20798) );
  INV_X1 U12316 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n21296) );
  INV_X1 U12317 ( .A(n20113), .ZN(n21286) );
  INV_X1 U12318 ( .A(n18071), .ZN(n18077) );
  INV_X1 U12319 ( .A(n14376), .ZN(n14301) );
  OAI21_X1 U12321 ( .B1(n15806), .B2(n21646), .A(n11302), .ZN(P1_U2809) );
  AOI21_X1 U12322 ( .B1(n12519), .B2(n21611), .A(n11029), .ZN(n11302) );
  AOI21_X1 U12323 ( .B1(n12641), .B2(n19929), .A(n11304), .ZN(n11303) );
  OAI21_X1 U12324 ( .B1(n15833), .B2(n21655), .A(n12509), .ZN(P1_U2968) );
  INV_X1 U12325 ( .A(n18526), .ZN(n14808) );
  NAND2_X1 U12326 ( .A1(n15452), .A2(n15451), .ZN(n15453) );
  NAND2_X1 U12327 ( .A1(n15470), .A2(n15469), .ZN(n15471) );
  OAI21_X1 U12328 ( .B1(n16255), .B2(n18606), .A(n11316), .ZN(P2_U3016) );
  AND2_X1 U12329 ( .A1(n11318), .A2(n11317), .ZN(n11316) );
  OR2_X1 U12330 ( .A1(n18498), .A2(n18605), .ZN(n11318) );
  AOI21_X1 U12331 ( .B1(n16253), .B2(n18568), .A(n15492), .ZN(n11317) );
  INV_X1 U12332 ( .A(n11346), .ZN(n16421) );
  OAI211_X1 U12333 ( .C1(n18474), .C2(n18605), .A(n11348), .B(n11347), .ZN(
        n11346) );
  OR2_X1 U12334 ( .A1(n16412), .A2(n18594), .ZN(n11347) );
  NAND2_X1 U12335 ( .A1(n11090), .A2(n11086), .ZN(P2_U3020) );
  OR2_X1 U12336 ( .A1(n16454), .A2(n18617), .ZN(n11090) );
  INV_X1 U12337 ( .A(n11087), .ZN(n11086) );
  OAI21_X1 U12338 ( .B1(n16456), .B2(n18606), .A(n11088), .ZN(n11087) );
  OAI211_X1 U12339 ( .C1(n16465), .C2(n18606), .A(n11233), .B(n11232), .ZN(
        P2_U3025) );
  NOR2_X1 U12340 ( .A1(n16464), .A2(n11234), .ZN(n11233) );
  OR2_X1 U12341 ( .A1(n16463), .A2(n18617), .ZN(n11232) );
  AND2_X1 U12342 ( .A1(n18363), .A2(n18591), .ZN(n11234) );
  NAND2_X1 U12343 ( .A1(n20565), .A2(n20577), .ZN(n20566) );
  NAND2_X1 U12344 ( .A1(n20523), .A2(n20577), .ZN(n20524) );
  OR2_X1 U12345 ( .A1(n15620), .A2(n15619), .ZN(n15559) );
  AND2_X1 U12346 ( .A1(n11441), .A2(n13230), .ZN(n10980) );
  AND2_X1 U12347 ( .A1(n11425), .A2(n11050), .ZN(n10981) );
  INV_X1 U12348 ( .A(n12810), .ZN(n13822) );
  AND2_X2 U12349 ( .A1(n13041), .A2(n12874), .ZN(n12890) );
  NAND2_X1 U12350 ( .A1(n15602), .A2(n11186), .ZN(n10982) );
  OR2_X1 U12351 ( .A1(n10982), .A2(n11474), .ZN(n10983) );
  NOR2_X1 U12352 ( .A1(n14460), .A2(n11074), .ZN(n10984) );
  OR3_X1 U12353 ( .A1(n18488), .A2(n15139), .A3(n15487), .ZN(n10985) );
  NAND2_X1 U12354 ( .A1(n15602), .A2(n11187), .ZN(n15551) );
  NAND2_X1 U12355 ( .A1(n11258), .A2(n11256), .ZN(n10986) );
  AND2_X1 U12356 ( .A1(n11320), .A2(n14492), .ZN(n10989) );
  NAND2_X2 U12357 ( .A1(n13647), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12787) );
  AND2_X1 U12358 ( .A1(n16063), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13367) );
  AND2_X1 U12359 ( .A1(n11237), .A2(n15272), .ZN(n10991) );
  AND2_X1 U12360 ( .A1(n11217), .A2(n11215), .ZN(n10992) );
  AND2_X1 U12361 ( .A1(n11340), .A2(n13722), .ZN(n10993) );
  NAND2_X1 U12362 ( .A1(n16160), .A2(n16159), .ZN(n16151) );
  NOR2_X1 U12363 ( .A1(n11065), .A2(n21523), .ZN(n10994) );
  AND2_X1 U12364 ( .A1(n11230), .A2(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n10995) );
  AND2_X1 U12365 ( .A1(n11386), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n10996) );
  AND2_X1 U12366 ( .A1(n11389), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n10997) );
  AND2_X1 U12367 ( .A1(n11381), .A2(n11380), .ZN(n10998) );
  OR3_X1 U12368 ( .A1(n15612), .A2(n11301), .A3(n11298), .ZN(n10999) );
  AND2_X1 U12369 ( .A1(n10998), .A2(P1_REIP_REG_5__SCAN_IN), .ZN(n11000) );
  NAND2_X1 U12370 ( .A1(n11329), .A2(n11334), .ZN(n14139) );
  AND2_X1 U12371 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n11001) );
  AND2_X1 U12372 ( .A1(n11001), .A2(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11002) );
  AND2_X1 U12373 ( .A1(n15305), .A2(n11078), .ZN(n11003) );
  AND2_X1 U12374 ( .A1(n11002), .A2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n11004) );
  AND2_X1 U12375 ( .A1(n11290), .A2(n11071), .ZN(n11005) );
  AND2_X1 U12376 ( .A1(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n11006) );
  AND2_X1 U12377 ( .A1(n11383), .A2(P1_REIP_REG_30__SCAN_IN), .ZN(n11007) );
  NAND2_X2 U12378 ( .A1(n12523), .A2(n13747), .ZN(n12592) );
  INV_X2 U12379 ( .A(n20193), .ZN(n14589) );
  NAND2_X1 U12380 ( .A1(n11129), .A2(n12807), .ZN(n12851) );
  OR2_X1 U12381 ( .A1(n16503), .A2(n16502), .ZN(n11008) );
  OR3_X1 U12382 ( .A1(n21532), .A2(n11367), .A3(n11365), .ZN(n11009) );
  OR3_X1 U12383 ( .A1(n15179), .A2(n11287), .A3(n15168), .ZN(n11010) );
  OR2_X1 U12384 ( .A1(n15531), .A2(n15494), .ZN(n11011) );
  NAND2_X1 U12385 ( .A1(n14986), .A2(n11245), .ZN(n15020) );
  INV_X1 U12386 ( .A(n14013), .ZN(n12867) );
  NOR2_X1 U12387 ( .A1(n14523), .A2(n14522), .ZN(n14604) );
  BUF_X1 U12388 ( .A(n14556), .Z(n14603) );
  NOR2_X1 U12389 ( .A1(n17033), .A2(n16531), .ZN(n11013) );
  INV_X1 U12390 ( .A(n11625), .ZN(n11697) );
  NOR3_X1 U12391 ( .A1(n21600), .A2(n11377), .A3(n11376), .ZN(n11375) );
  AND3_X1 U12392 ( .A1(n12757), .A2(n12755), .A3(n14994), .ZN(n11014) );
  INV_X1 U12393 ( .A(n14544), .ZN(n14684) );
  NOR2_X1 U12394 ( .A1(n16318), .A2(n16475), .ZN(n11015) );
  NAND2_X1 U12395 ( .A1(n11183), .A2(n11691), .ZN(n11783) );
  OR2_X1 U12396 ( .A1(n15493), .A2(n20018), .ZN(n11016) );
  AND3_X1 U12397 ( .A1(n11446), .A2(n13748), .A3(n11445), .ZN(n11017) );
  NAND2_X1 U12398 ( .A1(n15596), .A2(n11467), .ZN(n11018) );
  NAND2_X1 U12399 ( .A1(n11490), .A2(n11491), .ZN(n11617) );
  NAND2_X1 U12400 ( .A1(n12379), .A2(n12380), .ZN(n12378) );
  AND2_X1 U12401 ( .A1(n14819), .A2(n14823), .ZN(n14970) );
  INV_X1 U12402 ( .A(n14968), .ZN(n15119) );
  NAND2_X1 U12403 ( .A1(n11406), .A2(n11410), .ZN(n15342) );
  AND2_X1 U12404 ( .A1(n15579), .A2(n11005), .ZN(n11019) );
  INV_X1 U12405 ( .A(n11611), .ZN(n11148) );
  AND4_X1 U12406 ( .A1(n14725), .A2(n14724), .A3(n14723), .A4(n14722), .ZN(
        n11020) );
  NAND2_X1 U12407 ( .A1(n11098), .A2(n19676), .ZN(n12801) );
  AND2_X1 U12408 ( .A1(n12862), .A2(n12746), .ZN(n11021) );
  AND2_X1 U12409 ( .A1(n15306), .A2(n11284), .ZN(n11022) );
  OR2_X1 U12410 ( .A1(n17721), .A2(n17774), .ZN(n11260) );
  INV_X1 U12411 ( .A(n15283), .ZN(n11433) );
  INV_X1 U12412 ( .A(n13662), .ZN(n15506) );
  OR2_X2 U12413 ( .A1(n11570), .A2(n11569), .ZN(n13662) );
  INV_X1 U12414 ( .A(n11125), .ZN(n13305) );
  NAND2_X1 U12415 ( .A1(n11124), .A2(n19203), .ZN(n11125) );
  OR2_X1 U12416 ( .A1(n12341), .A2(n12342), .ZN(n11023) );
  AND2_X1 U12417 ( .A1(n13292), .A2(n11126), .ZN(n11025) );
  OR2_X1 U12418 ( .A1(n11143), .A2(n11139), .ZN(n11026) );
  INV_X1 U12419 ( .A(n11240), .ZN(n16350) );
  OR2_X1 U12420 ( .A1(n17033), .A2(n11243), .ZN(n11240) );
  NOR2_X1 U12421 ( .A1(n10982), .A2(n11472), .ZN(n12379) );
  AND2_X1 U12422 ( .A1(n15275), .A2(n11395), .ZN(n15272) );
  INV_X1 U12423 ( .A(n11403), .ZN(n11401) );
  NAND2_X1 U12424 ( .A1(n15408), .A2(n11404), .ZN(n11403) );
  NAND2_X1 U12425 ( .A1(n13827), .A2(n11309), .ZN(n11027) );
  NAND2_X1 U12426 ( .A1(n12523), .A2(n14182), .ZN(n13571) );
  INV_X1 U12427 ( .A(n13571), .ZN(n11613) );
  AND2_X1 U12428 ( .A1(n15596), .A2(n11466), .ZN(n11028) );
  NAND2_X1 U12429 ( .A1(n12643), .A2(n11303), .ZN(n11029) );
  INV_X1 U12430 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n12645) );
  INV_X1 U12431 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n12648) );
  OR2_X1 U12432 ( .A1(n15179), .A2(n11287), .ZN(n11030) );
  AND3_X1 U12433 ( .A1(n14715), .A2(n14720), .A3(n14716), .ZN(n11031) );
  AND2_X1 U12434 ( .A1(n12851), .A2(n18108), .ZN(n11032) );
  AND2_X2 U12435 ( .A1(n16068), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13368) );
  NAND2_X1 U12436 ( .A1(n14897), .A2(n11099), .ZN(n14959) );
  OR2_X1 U12437 ( .A1(n15620), .A2(n11470), .ZN(n11471) );
  AND2_X1 U12438 ( .A1(n11016), .A2(n12491), .ZN(n11033) );
  INV_X1 U12439 ( .A(n16269), .ZN(n11404) );
  NAND2_X1 U12440 ( .A1(n15933), .A2(n12461), .ZN(n11034) );
  AND2_X1 U12441 ( .A1(n11294), .A2(n11292), .ZN(n11035) );
  INV_X1 U12442 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13622) );
  NAND2_X1 U12443 ( .A1(n12860), .A2(n12859), .ZN(n13665) );
  NAND2_X1 U12444 ( .A1(n13581), .A2(n16740), .ZN(n11036) );
  INV_X1 U12445 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n16719) );
  NAND2_X1 U12446 ( .A1(n11619), .A2(n11612), .ZN(n12511) );
  NOR2_X1 U12447 ( .A1(n13725), .A2(n13905), .ZN(n12510) );
  OR2_X1 U12448 ( .A1(n15139), .A2(n13408), .ZN(n11037) );
  OR2_X1 U12449 ( .A1(n17574), .A2(n11223), .ZN(n11038) );
  NAND2_X1 U12450 ( .A1(n13682), .A2(n11037), .ZN(n11342) );
  NAND2_X1 U12451 ( .A1(n12773), .A2(n13184), .ZN(n13247) );
  OR3_X1 U12452 ( .A1(n17797), .A2(n11200), .A3(n11199), .ZN(n11039) );
  INV_X1 U12453 ( .A(n11443), .ZN(n12440) );
  NAND2_X1 U12454 ( .A1(n13732), .A2(n11611), .ZN(n11443) );
  NAND2_X1 U12455 ( .A1(n11342), .A2(n11344), .ZN(n13683) );
  INV_X1 U12456 ( .A(n11861), .ZN(n14460) );
  AND2_X1 U12457 ( .A1(n16160), .A2(n11421), .ZN(n11040) );
  INV_X1 U12458 ( .A(n12388), .ZN(n21671) );
  AND2_X1 U12459 ( .A1(n16366), .A2(n11386), .ZN(n11041) );
  AND2_X1 U12460 ( .A1(n17025), .A2(n11389), .ZN(n11042) );
  INV_X1 U12461 ( .A(n12746), .ZN(n13233) );
  NAND2_X1 U12462 ( .A1(n14220), .A2(n14221), .ZN(n14489) );
  AND2_X1 U12463 ( .A1(n14220), .A2(n11320), .ZN(n11043) );
  OR2_X1 U12464 ( .A1(n11181), .A2(n11829), .ZN(n14306) );
  XNOR2_X1 U12465 ( .A(n15137), .B(n15243), .ZN(n16405) );
  INV_X1 U12466 ( .A(n21256), .ZN(n11276) );
  NOR2_X1 U12467 ( .A1(n17967), .A2(n17954), .ZN(n17759) );
  INV_X1 U12468 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11493) );
  AND2_X1 U12469 ( .A1(n15149), .A2(n11417), .ZN(n11044) );
  AND2_X1 U12470 ( .A1(n11355), .A2(n11354), .ZN(n11045) );
  NOR2_X1 U12471 ( .A1(n11829), .A2(n14204), .ZN(n14255) );
  AND2_X1 U12472 ( .A1(n11044), .A2(n16586), .ZN(n11046) );
  NAND2_X1 U12473 ( .A1(n13701), .A2(n12865), .ZN(n13839) );
  AND2_X1 U12474 ( .A1(n16303), .A2(n16302), .ZN(n11047) );
  NOR2_X1 U12475 ( .A1(n14460), .A2(n11876), .ZN(n11048) );
  AND2_X2 U12476 ( .A1(n12756), .A2(n11014), .ZN(n13443) );
  INV_X1 U12477 ( .A(n13443), .ZN(n11133) );
  NAND2_X1 U12478 ( .A1(n12633), .A2(n13747), .ZN(n11049) );
  INV_X1 U12479 ( .A(n11462), .ZN(n11461) );
  NOR3_X1 U12480 ( .A1(n11876), .A2(n11464), .A3(n11463), .ZN(n11462) );
  AND2_X1 U12481 ( .A1(n14222), .A2(n13397), .ZN(n11050) );
  OR2_X1 U12482 ( .A1(n21600), .A2(n21601), .ZN(n11051) );
  AND2_X1 U12483 ( .A1(n12478), .A2(n12477), .ZN(n11052) );
  AND2_X1 U12484 ( .A1(n11615), .A2(n11611), .ZN(n11053) );
  NOR2_X1 U12485 ( .A1(n15612), .A2(n11296), .ZN(n11300) );
  OR2_X1 U12486 ( .A1(n11461), .A2(n15083), .ZN(n11054) );
  INV_X1 U12487 ( .A(n11366), .ZN(n21541) );
  NOR2_X1 U12488 ( .A1(n21532), .A2(n11367), .ZN(n11366) );
  INV_X1 U12489 ( .A(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n16999) );
  INV_X1 U12490 ( .A(n11279), .ZN(n14859) );
  INV_X1 U12491 ( .A(n11424), .ZN(n11423) );
  NAND2_X1 U12492 ( .A1(n10981), .A2(n14514), .ZN(n11424) );
  OR2_X1 U12493 ( .A1(n11252), .A2(n11251), .ZN(n11055) );
  AND2_X1 U12494 ( .A1(n11207), .A2(n11814), .ZN(n11056) );
  OR2_X1 U12495 ( .A1(n15881), .A2(n15858), .ZN(n11057) );
  AND2_X1 U12496 ( .A1(n11324), .A2(n11323), .ZN(n11058) );
  AND2_X1 U12497 ( .A1(n11489), .A2(n11188), .ZN(n11059) );
  OR2_X1 U12498 ( .A1(n21600), .A2(n11377), .ZN(n11060) );
  INV_X1 U12499 ( .A(n15723), .ZN(n11221) );
  AND2_X1 U12500 ( .A1(n11045), .A2(n15058), .ZN(n11061) );
  AND2_X1 U12501 ( .A1(n13928), .A2(n13391), .ZN(n11062) );
  NAND2_X1 U12502 ( .A1(n13614), .A2(n13587), .ZN(n13625) );
  AND2_X1 U12503 ( .A1(n17701), .A2(n11002), .ZN(n11063) );
  INV_X1 U12504 ( .A(n15595), .ZN(n11468) );
  AND2_X1 U12505 ( .A1(n15049), .A2(n15048), .ZN(n18591) );
  AND2_X1 U12506 ( .A1(n15049), .A2(n15046), .ZN(n18622) );
  NOR2_X1 U12507 ( .A1(n13329), .A2(n11330), .ZN(n14453) );
  BUF_X1 U12508 ( .A(n12738), .Z(n16057) );
  OR2_X1 U12509 ( .A1(n15447), .A2(n15446), .ZN(n11064) );
  NAND2_X2 U12510 ( .A1(n16758), .A2(n20029), .ZN(n21655) );
  AND2_X1 U12511 ( .A1(n12633), .A2(n10998), .ZN(n11065) );
  AND2_X1 U12512 ( .A1(n11339), .A2(n15323), .ZN(n11066) );
  INV_X1 U12513 ( .A(n17774), .ZN(n21115) );
  OR2_X1 U12514 ( .A1(n15131), .A2(n18197), .ZN(n11067) );
  OR3_X1 U12515 ( .A1(n15447), .A2(n11393), .A3(n11392), .ZN(n11068) );
  NAND2_X1 U12516 ( .A1(n13961), .A2(n13838), .ZN(n13857) );
  AND2_X1 U12517 ( .A1(n11327), .A2(n11326), .ZN(n11069) );
  OR2_X1 U12518 ( .A1(n12939), .A2(n12938), .ZN(n14514) );
  INV_X1 U12519 ( .A(n14514), .ZN(n11426) );
  OR2_X1 U12520 ( .A1(n13944), .A2(n11180), .ZN(n11070) );
  AND2_X1 U12521 ( .A1(n15543), .A2(n15869), .ZN(n11071) );
  AND2_X1 U12522 ( .A1(n11005), .A2(n15529), .ZN(n11072) );
  AND2_X1 U12523 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n11073) );
  INV_X1 U12524 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11448) );
  NAND2_X1 U12525 ( .A1(n13839), .A2(n10981), .ZN(n11427) );
  NAND2_X1 U12526 ( .A1(n11631), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n11958) );
  INV_X1 U12527 ( .A(n11958), .ZN(n11991) );
  OR2_X1 U12528 ( .A1(n11876), .A2(n11464), .ZN(n11074) );
  AND2_X1 U12529 ( .A1(n12513), .A2(n13464), .ZN(n11075) );
  AND2_X1 U12530 ( .A1(n11420), .A2(n11419), .ZN(n11076) );
  AND2_X1 U12531 ( .A1(n11259), .A2(n21046), .ZN(n11077) );
  AND2_X2 U12532 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13587) );
  INV_X1 U12533 ( .A(n20567), .ZN(n11197) );
  OR2_X1 U12534 ( .A1(n15131), .A2(n18411), .ZN(n11078) );
  AND2_X1 U12535 ( .A1(n13419), .A2(n13418), .ZN(n11079) );
  NAND2_X1 U12536 ( .A1(n12382), .A2(n21881), .ZN(n20018) );
  INV_X1 U12537 ( .A(P1_REIP_REG_5__SCAN_IN), .ZN(n11382) );
  AND2_X1 U12538 ( .A1(n12769), .A2(n11124), .ZN(n11080) );
  AND3_X1 U12539 ( .A1(n15248), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        n15247), .ZN(n11081) );
  INV_X1 U12540 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n11379) );
  INV_X1 U12541 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n11231) );
  AND3_X1 U12542 ( .A1(n15885), .A2(n15889), .A3(n21398), .ZN(n11082) );
  INV_X1 U12543 ( .A(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n11228) );
  INV_X1 U12544 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n11199) );
  INV_X1 U12545 ( .A(n18261), .ZN(n18634) );
  OAI21_X2 U12546 ( .B1(n13703), .B2(n13702), .A(n13701), .ZN(n19328) );
  OAI21_X1 U12547 ( .B1(n13666), .B2(n13665), .A(n12861), .ZN(n13703) );
  NAND2_X1 U12548 ( .A1(n13702), .A2(n13703), .ZN(n13701) );
  NOR2_X1 U12549 ( .A1(n21758), .A2(n21756), .ZN(n18071) );
  NOR2_X2 U12550 ( .A1(n14244), .A2(n14173), .ZN(n22057) );
  NAND3_X1 U12551 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n21321), .A3(n13904), 
        .ZN(n14244) );
  OAI22_X2 U12552 ( .A1(n20086), .A2(n14243), .B1(n14242), .B2(n13898), .ZN(
        n21949) );
  NAND2_X1 U12553 ( .A1(n20009), .A2(n14301), .ZN(n14243) );
  INV_X1 U12554 ( .A(n22203), .ZN(n11083) );
  INV_X1 U12555 ( .A(n11083), .ZN(n11084) );
  OR2_X1 U12556 ( .A1(n19328), .A2(n19219), .ZN(n19169) );
  NAND2_X1 U12557 ( .A1(n19328), .A2(n19219), .ZN(n19315) );
  NAND2_X1 U12558 ( .A1(n19328), .A2(n17077), .ZN(n19267) );
  NOR2_X2 U12559 ( .A1(n18682), .A2(n19009), .ZN(n18757) );
  NAND2_X1 U12560 ( .A1(n18703), .A2(n18968), .ZN(n19009) );
  OAI22_X2 U12561 ( .A1(n20091), .A2(n14243), .B1(n16882), .B2(n13898), .ZN(
        n22018) );
  OAI22_X2 U12562 ( .A1(n20097), .A2(n14243), .B1(n16879), .B2(n13898), .ZN(
        n22123) );
  INV_X1 U12563 ( .A(n15703), .ZN(n15707) );
  CLKBUF_X1 U12564 ( .A(n19719), .Z(n11085) );
  XNOR2_X2 U12565 ( .A(n13815), .B(n13816), .ZN(n14816) );
  NAND2_X1 U12566 ( .A1(n15373), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15425) );
  NAND4_X1 U12567 ( .A1(n12680), .A2(n12677), .A3(n12679), .A4(n12678), .ZN(
        n11094) );
  NAND4_X1 U12568 ( .A1(n12673), .A2(n12676), .A3(n12675), .A4(n12674), .ZN(
        n11096) );
  NAND3_X1 U12569 ( .A1(n12705), .A2(n12706), .A3(n12704), .ZN(n12800) );
  NOR2_X2 U12570 ( .A1(n14959), .A2(n14958), .ZN(n14985) );
  NAND2_X1 U12571 ( .A1(n16270), .A2(n16271), .ZN(n11100) );
  NAND2_X2 U12572 ( .A1(n11108), .A2(n11106), .ZN(n12746) );
  NAND2_X1 U12573 ( .A1(n11107), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11106) );
  NAND4_X1 U12574 ( .A1(n12684), .A2(n12685), .A3(n12682), .A4(n12683), .ZN(
        n11107) );
  NAND2_X1 U12575 ( .A1(n11109), .A2(n12681), .ZN(n11108) );
  NAND4_X1 U12576 ( .A1(n12687), .A2(n12686), .A3(n12689), .A4(n12688), .ZN(
        n11109) );
  AND2_X2 U12577 ( .A1(n11112), .A2(n14817), .ZN(n19310) );
  AND2_X2 U12578 ( .A1(n11112), .A2(n14818), .ZN(n19301) );
  AND2_X2 U12579 ( .A1(n11112), .A2(n14822), .ZN(n19324) );
  AND2_X2 U12580 ( .A1(n11112), .A2(n14819), .ZN(n16673) );
  NAND3_X1 U12582 ( .A1(n15275), .A2(n11395), .A3(n15139), .ZN(n11116) );
  NAND4_X1 U12583 ( .A1(n12731), .A2(n12748), .A3(n12732), .A4(n19559), .ZN(
        n11117) );
  NAND4_X1 U12584 ( .A1(n13233), .A2(n12754), .A3(n19464), .A4(n12862), .ZN(
        n14001) );
  NAND2_X1 U12585 ( .A1(n12849), .A2(n11119), .ZN(n18108) );
  INV_X1 U12586 ( .A(n13155), .ZN(n11122) );
  INV_X1 U12587 ( .A(n13156), .ZN(n11123) );
  CLKBUF_X1 U12588 ( .A(n12746), .Z(n11124) );
  NOR2_X2 U12589 ( .A1(n11124), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n13277) );
  NAND2_X1 U12590 ( .A1(n12839), .A2(n12838), .ZN(n12822) );
  INV_X1 U12591 ( .A(n12819), .ZN(n11131) );
  OAI21_X2 U12592 ( .B1(n12865), .B2(n11424), .A(n11134), .ZN(n14512) );
  NAND3_X1 U12593 ( .A1(n13702), .A2(n13703), .A3(n11423), .ZN(n11134) );
  AND2_X2 U12594 ( .A1(n12837), .A2(n12864), .ZN(n13702) );
  AND2_X2 U12595 ( .A1(n16160), .A2(n11076), .ZN(n16131) );
  NOR2_X4 U12596 ( .A1(n15055), .A2(n15056), .ZN(n16160) );
  NAND4_X1 U12597 ( .A1(n11036), .A2(n13739), .A3(n11138), .A4(n11137), .ZN(
        n11140) );
  OAI21_X2 U12598 ( .B1(n11140), .B2(n11141), .A(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n11625) );
  OAI21_X2 U12599 ( .B1(n11625), .B2(n11448), .A(n11627), .ZN(n11671) );
  NAND2_X1 U12600 ( .A1(n12492), .A2(n11033), .ZN(P1_U2970) );
  NAND2_X1 U12601 ( .A1(n13695), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n12404) );
  NAND3_X1 U12602 ( .A1(n11460), .A2(n11057), .A3(n12476), .ZN(n11145) );
  NAND2_X1 U12603 ( .A1(n11149), .A2(n11615), .ZN(n13469) );
  NAND2_X2 U12604 ( .A1(n15996), .A2(n12459), .ZN(n15995) );
  NAND2_X2 U12605 ( .A1(n15896), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n12473) );
  NAND3_X1 U12606 ( .A1(n12768), .A2(n12748), .A3(n19464), .ZN(n13236) );
  NAND2_X1 U12607 ( .A1(n11585), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n11586) );
  INV_X1 U12608 ( .A(n11180), .ZN(n13460) );
  AND2_X1 U12609 ( .A1(n12308), .A2(n11180), .ZN(n12322) );
  OAI21_X1 U12610 ( .B1(n11628), .B2(n11180), .A(n13599), .ZN(n11179) );
  AOI21_X1 U12611 ( .B1(n13593), .B2(n11180), .A(n11075), .ZN(n20030) );
  NAND3_X1 U12612 ( .A1(n13914), .A2(n13913), .A3(n14307), .ZN(n11181) );
  XNOR2_X2 U12613 ( .A(n11182), .B(n11693), .ZN(n11639) );
  OAI21_X2 U12614 ( .B1(n11625), .B2(n11493), .A(n11624), .ZN(n11182) );
  NAND2_X1 U12615 ( .A1(n12394), .A2(n11667), .ZN(n11668) );
  NAND3_X1 U12616 ( .A1(n11207), .A2(n11991), .A3(n11814), .ZN(n11185) );
  NAND2_X1 U12617 ( .A1(n11185), .A2(n11809), .ZN(n11810) );
  INV_X1 U12618 ( .A(n11056), .ZN(n14401) );
  AND2_X4 U12619 ( .A1(n11190), .A2(n13977), .ZN(n11979) );
  AND2_X4 U12620 ( .A1(n11190), .A2(n11500), .ZN(n11537) );
  AND2_X1 U12621 ( .A1(n13614), .A2(n11190), .ZN(n11676) );
  NAND2_X1 U12622 ( .A1(n20549), .A2(n11196), .ZN(n11195) );
  INV_X1 U12623 ( .A(n17785), .ZN(n17800) );
  NAND2_X1 U12624 ( .A1(n20502), .A2(n11204), .ZN(n11203) );
  NAND2_X1 U12625 ( .A1(n11802), .A2(n11803), .ZN(n11814) );
  NAND3_X1 U12626 ( .A1(n11207), .A2(n11814), .A3(n12440), .ZN(n12387) );
  NAND2_X1 U12627 ( .A1(n11208), .A2(n11209), .ZN(n20480) );
  NAND2_X1 U12629 ( .A1(n20449), .A2(n20577), .ZN(n20451) );
  INV_X1 U12630 ( .A(n12473), .ZN(n11213) );
  INV_X1 U12631 ( .A(n11212), .ZN(n11214) );
  OAI21_X1 U12632 ( .B1(n11219), .B2(n11213), .A(n15994), .ZN(n12476) );
  OAI21_X2 U12633 ( .B1(n12473), .B2(n11218), .A(n11214), .ZN(n15734) );
  NAND2_X2 U12634 ( .A1(n12473), .A2(n15897), .ZN(n15882) );
  INV_X1 U12635 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n11222) );
  INV_X1 U12636 ( .A(n11235), .ZN(n12764) );
  NAND4_X1 U12637 ( .A1(n12731), .A2(n12747), .A3(n12750), .A4(n12732), .ZN(
        n11235) );
  AND2_X1 U12638 ( .A1(n14008), .A2(n12746), .ZN(n12757) );
  AND2_X1 U12639 ( .A1(n12828), .A2(n12754), .ZN(n12756) );
  NAND2_X1 U12640 ( .A1(n11245), .A2(n15269), .ZN(n11395) );
  NAND2_X1 U12641 ( .A1(n11246), .A2(n15138), .ZN(n11247) );
  INV_X1 U12642 ( .A(n16405), .ZN(n11246) );
  NAND3_X1 U12643 ( .A1(n11248), .A2(n11046), .A3(n11247), .ZN(n11416) );
  NAND3_X1 U12644 ( .A1(n15110), .A2(n15138), .A3(n15109), .ZN(n11248) );
  NAND2_X1 U12645 ( .A1(n15110), .A2(n15109), .ZN(n16406) );
  NAND2_X1 U12646 ( .A1(n11249), .A2(n15138), .ZN(n16398) );
  NAND2_X2 U12647 ( .A1(n16046), .A2(n14816), .ZN(n14821) );
  NAND3_X1 U12648 ( .A1(n16307), .A2(n16306), .A3(n16308), .ZN(n16311) );
  NAND2_X1 U12649 ( .A1(n11253), .A2(n16558), .ZN(n16375) );
  XNOR2_X1 U12650 ( .A(n11253), .B(n16559), .ZN(n17026) );
  NAND3_X1 U12651 ( .A1(n11255), .A2(n11260), .A3(n11077), .ZN(n21119) );
  NOR2_X1 U12652 ( .A1(n17721), .A2(n21042), .ZN(n11257) );
  NAND2_X2 U12653 ( .A1(n11020), .A2(n11262), .ZN(n20783) );
  NAND3_X1 U12654 ( .A1(n14727), .A2(n11265), .A3(n11264), .ZN(n11263) );
  NAND4_X1 U12655 ( .A1(n11272), .A2(n14608), .A3(n14606), .A4(n11268), .ZN(
        n14622) );
  NAND4_X1 U12656 ( .A1(n11271), .A2(n14611), .A3(n14607), .A4(n14605), .ZN(
        n11270) );
  NAND2_X2 U12657 ( .A1(n11274), .A2(n14680), .ZN(n20113) );
  INV_X2 U12658 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n20829) );
  INV_X2 U12659 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n20825) );
  OR2_X2 U12660 ( .A1(n21315), .A2(n20171), .ZN(n17971) );
  AND2_X4 U12661 ( .A1(n14013), .A2(n13211), .ZN(n12738) );
  AND2_X1 U12662 ( .A1(n15018), .A2(n13525), .ZN(n11280) );
  NAND2_X1 U12663 ( .A1(n13526), .A2(n13525), .ZN(n11279) );
  NAND2_X1 U12664 ( .A1(n15143), .A2(n11281), .ZN(n15161) );
  INV_X1 U12665 ( .A(n15140), .ZN(n11282) );
  NAND2_X1 U12666 ( .A1(n15306), .A2(n11003), .ZN(n15403) );
  NAND2_X1 U12667 ( .A1(n15306), .A2(n15305), .ZN(n15399) );
  NAND2_X1 U12668 ( .A1(n11293), .A2(n11035), .ZN(n14499) );
  INV_X1 U12669 ( .A(n11300), .ZN(n15592) );
  INV_X1 U12670 ( .A(n15605), .ZN(n11301) );
  INV_X1 U12671 ( .A(n13888), .ZN(n11306) );
  NAND2_X1 U12672 ( .A1(n11306), .A2(n11307), .ZN(n13881) );
  NOR2_X2 U12673 ( .A1(n21174), .A2(n17706), .ZN(n20858) );
  INV_X1 U12674 ( .A(n13857), .ZN(n11311) );
  NAND2_X1 U12675 ( .A1(n11311), .A2(n11312), .ZN(n14289) );
  NAND2_X1 U12676 ( .A1(n14220), .A2(n11319), .ZN(n14946) );
  INV_X1 U12677 ( .A(n13329), .ZN(n11329) );
  NAND2_X1 U12678 ( .A1(n11331), .A2(n11329), .ZN(n15041) );
  NAND2_X1 U12679 ( .A1(n11342), .A2(n10993), .ZN(n13721) );
  NAND2_X1 U12680 ( .A1(n16478), .A2(n11350), .ZN(n15381) );
  NAND2_X1 U12681 ( .A1(n14450), .A2(n11061), .ZN(n16503) );
  NAND3_X1 U12682 ( .A1(n11368), .A2(n11031), .A3(n14717), .ZN(n14761) );
  OR2_X1 U12683 ( .A1(n14718), .A2(n11371), .ZN(n11370) );
  NAND3_X1 U12684 ( .A1(n11374), .A2(n11373), .A3(n11372), .ZN(n11371) );
  INV_X1 U12685 ( .A(n11375), .ZN(n21616) );
  NAND2_X1 U12686 ( .A1(n15550), .A2(n11007), .ZN(n12642) );
  NAND2_X1 U12687 ( .A1(n15550), .A2(P1_REIP_REG_28__SCAN_IN), .ZN(n15533) );
  INV_X1 U12688 ( .A(n12642), .ZN(n12641) );
  INV_X2 U12689 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n20822) );
  NAND2_X1 U12690 ( .A1(n15223), .A2(n15222), .ZN(n11413) );
  INV_X1 U12691 ( .A(n11427), .ZN(n14515) );
  NAND2_X1 U12692 ( .A1(n11429), .A2(n11431), .ZN(n17033) );
  NAND2_X1 U12693 ( .A1(n15373), .A2(n11434), .ZN(n16297) );
  AND2_X2 U12694 ( .A1(n15373), .A2(n11435), .ZN(n16286) );
  NAND2_X1 U12695 ( .A1(n14992), .A2(n12765), .ZN(n13544) );
  NOR2_X2 U12696 ( .A1(n16046), .A2(n14816), .ZN(n14811) );
  NAND3_X1 U12697 ( .A1(n10980), .A2(n12790), .A3(n11440), .ZN(n12776) );
  NAND2_X1 U12698 ( .A1(n13550), .A2(n14002), .ZN(n12790) );
  AND3_X2 U12699 ( .A1(n12775), .A2(n13247), .A3(n12774), .ZN(n13550) );
  NAND2_X1 U12700 ( .A1(n12764), .A2(n19676), .ZN(n13230) );
  AND3_X1 U12701 ( .A1(n11446), .A2(n13748), .A3(n13945), .ZN(n11636) );
  XNOR2_X2 U12702 ( .A(n11671), .B(n11670), .ZN(n16743) );
  NAND2_X1 U12703 ( .A1(n11454), .A2(n11453), .ZN(n14467) );
  AND2_X1 U12704 ( .A1(n14468), .A2(n12432), .ZN(n11453) );
  INV_X1 U12705 ( .A(n12432), .ZN(n11455) );
  NAND2_X1 U12706 ( .A1(n11458), .A2(n11457), .ZN(n12470) );
  INV_X1 U12707 ( .A(n14870), .ZN(n11464) );
  NOR2_X2 U12708 ( .A1(n15620), .A2(n11469), .ZN(n15602) );
  INV_X1 U12709 ( .A(n11471), .ZN(n15560) );
  NOR2_X1 U12710 ( .A1(n10982), .A2(n15640), .ZN(n15539) );
  NAND2_X1 U12711 ( .A1(n11691), .A2(n11668), .ZN(n11786) );
  NAND3_X1 U12713 ( .A1(n11802), .A2(n13897), .A3(n11803), .ZN(n11816) );
  INV_X1 U12714 ( .A(n10964), .ZN(n16641) );
  OAI21_X1 U12715 ( .B1(n16017), .B2(n17046), .A(n15449), .ZN(n15450) );
  XOR2_X1 U12716 ( .A(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .B(n15448), .Z(
        n16017) );
  NAND2_X1 U12717 ( .A1(n16263), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15448) );
  NAND2_X1 U12718 ( .A1(n12699), .A2(n12681), .ZN(n12700) );
  OAI21_X2 U12719 ( .B1(n15020), .B2(n15420), .A(n18141), .ZN(n15108) );
  OR2_X1 U12720 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n12300), .ZN(
        n12329) );
  NOR2_X1 U12721 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11494) );
  INV_X1 U12722 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11492) );
  NAND2_X1 U12723 ( .A1(n12357), .A2(n13662), .ZN(n11614) );
  BUF_X4 U12724 ( .A(n11641), .Z(n12096) );
  OAI21_X1 U12725 ( .B1(n12808), .B2(n12789), .A(n12788), .ZN(n12793) );
  MUX2_X1 U12726 ( .A(n12770), .B(n13250), .S(n14008), .Z(n12775) );
  NAND2_X1 U12727 ( .A1(n12769), .A2(n14008), .ZN(n12732) );
  NAND2_X1 U12728 ( .A1(n16122), .A2(n16121), .ZN(n16120) );
  NOR3_X2 U12729 ( .A1(n16291), .A2(n16289), .A3(n16293), .ZN(n16270) );
  NAND2_X1 U12730 ( .A1(n14157), .A2(n21671), .ZN(n21786) );
  AND2_X1 U12731 ( .A1(n14823), .A2(n14822), .ZN(n14961) );
  AND2_X1 U12732 ( .A1(n14823), .A2(n14818), .ZN(n14968) );
  AND2_X1 U12733 ( .A1(n14823), .A2(n14817), .ZN(n14960) );
  INV_X1 U12734 ( .A(n11923), .ZN(n11960) );
  NAND2_X1 U12735 ( .A1(n12519), .A2(n12360), .ZN(n12377) );
  INV_X1 U12736 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n13554) );
  AND2_X1 U12737 ( .A1(n13265), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11477) );
  INV_X1 U12738 ( .A(n13277), .ZN(n13384) );
  AND2_X1 U12739 ( .A1(n16022), .A2(n16025), .ZN(n18250) );
  OR3_X1 U12740 ( .A1(n16416), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n15485), .ZN(n11478) );
  OR3_X1 U12741 ( .A1(n16416), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n15465), .ZN(n11479) );
  INV_X1 U12742 ( .A(n18885), .ZN(n14615) );
  AND2_X1 U12743 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(n21706), .ZN(n21710) );
  OR2_X1 U12744 ( .A1(n13680), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n11480) );
  OR2_X1 U12745 ( .A1(n13680), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n11481) );
  OR2_X1 U12746 ( .A1(n13680), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n11482) );
  INV_X1 U12747 ( .A(n21881), .ZN(n21915) );
  OR2_X1 U12748 ( .A1(n20037), .A2(n20089), .ZN(U212) );
  AND3_X1 U12749 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(P3_EAX_REG_3__SCAN_IN), 
        .A3(P3_EAX_REG_4__SCAN_IN), .ZN(n11483) );
  INV_X1 U12750 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n21695) );
  AND2_X1 U12751 ( .A1(n13116), .A2(n13136), .ZN(n11484) );
  OR2_X1 U12752 ( .A1(n16120), .A2(n13100), .ZN(n11485) );
  AND2_X1 U12753 ( .A1(n13117), .A2(n11484), .ZN(n11486) );
  AND4_X1 U12754 ( .A1(n14978), .A2(n14977), .A3(n14976), .A4(n14975), .ZN(
        n11487) );
  AND4_X1 U12755 ( .A1(n14965), .A2(n14964), .A3(n14963), .A4(n14962), .ZN(
        n11488) );
  AND2_X1 U12756 ( .A1(n12176), .A2(n12175), .ZN(n11489) );
  AND4_X1 U12757 ( .A1(n11544), .A2(n11543), .A3(n11542), .A4(n11541), .ZN(
        n11490) );
  AND4_X1 U12758 ( .A1(n11549), .A2(n11548), .A3(n11547), .A4(n11546), .ZN(
        n11491) );
  INV_X1 U12759 ( .A(n12520), .ZN(n11606) );
  NAND2_X1 U12760 ( .A1(n14298), .A2(n11606), .ZN(n11607) );
  NAND2_X1 U12761 ( .A1(n12703), .A2(n14993), .ZN(n12704) );
  INV_X1 U12762 ( .A(n12814), .ZN(n12815) );
  NAND2_X1 U12763 ( .A1(n21877), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12307) );
  OAI21_X1 U12764 ( .B1(n12297), .B2(n12307), .A(n12296), .ZN(n12318) );
  NAND2_X1 U12765 ( .A1(n12299), .A2(n12298), .ZN(n12330) );
  INV_X1 U12766 ( .A(n11849), .ZN(n11850) );
  BUF_X1 U12767 ( .A(n11878), .Z(n12223) );
  AND2_X1 U12768 ( .A1(n13746), .A2(n11632), .ZN(n11633) );
  AND2_X1 U12769 ( .A1(n19464), .A2(n14999), .ZN(n12747) );
  OAI21_X1 U12770 ( .B1(n14839), .B2(n14838), .A(n18090), .ZN(n14842) );
  NAND2_X1 U12771 ( .A1(n11488), .A2(n11487), .ZN(n14981) );
  AOI22_X1 U12772 ( .A1(n16064), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12866), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12736) );
  OR2_X1 U12773 ( .A1(n14643), .A2(n14644), .ZN(n14639) );
  AOI21_X1 U12774 ( .B1(n12330), .B2(n12329), .A(n12328), .ZN(n12338) );
  AND2_X1 U12775 ( .A1(n11761), .A2(n11760), .ZN(n11762) );
  INV_X1 U12776 ( .A(n12294), .ZN(n12023) );
  OR2_X1 U12777 ( .A1(n11840), .A2(n11839), .ZN(n12443) );
  AND2_X1 U12778 ( .A1(n11842), .A2(n11841), .ZN(n11849) );
  INV_X1 U12779 ( .A(n11614), .ZN(n13568) );
  INV_X1 U12780 ( .A(n13207), .ZN(n13180) );
  AND2_X1 U12781 ( .A1(n12653), .A2(n12681), .ZN(n12657) );
  AOI22_X1 U12782 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n16673), .B1(
        n19235), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n14845) );
  NOR2_X1 U12783 ( .A1(n14646), .A2(n14651), .ZN(n14638) );
  NAND2_X1 U12784 ( .A1(n13905), .A2(n13732), .ZN(n13945) );
  NAND2_X1 U12785 ( .A1(n12340), .A2(n12339), .ZN(n12342) );
  INV_X1 U12786 ( .A(n11772), .ZN(n11822) );
  AND2_X1 U12787 ( .A1(n15929), .A2(n12464), .ZN(n15782) );
  NAND2_X1 U12788 ( .A1(n11877), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11902) );
  OR2_X1 U12789 ( .A1(n13634), .A2(n11622), .ZN(n16740) );
  NAND2_X1 U12790 ( .A1(n21769), .A2(n21321), .ZN(n11737) );
  NAND2_X1 U12791 ( .A1(n12825), .A2(n12824), .ZN(n13819) );
  AND4_X1 U12792 ( .A1(n13365), .A2(n13364), .A3(n13363), .A4(n13362), .ZN(
        n13382) );
  INV_X1 U12793 ( .A(n15466), .ZN(n15467) );
  AND2_X1 U12794 ( .A1(n15205), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15217) );
  INV_X1 U12795 ( .A(n13384), .ZN(n15461) );
  INV_X1 U12796 ( .A(n12753), .ZN(n12862) );
  NAND2_X1 U12797 ( .A1(n12737), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12745) );
  AOI22_X1 U12798 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B1(n21263), .B2(n20825), .ZN(
        n14651) );
  NOR2_X1 U12799 ( .A1(n14624), .A2(n14615), .ZN(n20808) );
  AOI21_X1 U12800 ( .B1(n14626), .B2(n17146), .A(n20111), .ZN(n14627) );
  AOI21_X1 U12801 ( .B1(n12354), .B2(n12353), .A(n12352), .ZN(n13729) );
  INV_X1 U12802 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n11924) );
  NAND2_X1 U12803 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n11818) );
  AND2_X1 U12804 ( .A1(n12596), .A2(n12595), .ZN(n15611) );
  INV_X1 U12805 ( .A(n12617), .ZN(n12627) );
  INV_X1 U12806 ( .A(n11822), .ZN(n12285) );
  NAND2_X1 U12807 ( .A1(n16006), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12287) );
  INV_X1 U12808 ( .A(n13777), .ZN(n11812) );
  INV_X1 U12809 ( .A(n21319), .ZN(n14295) );
  AND2_X1 U12810 ( .A1(n21910), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n12294) );
  NOR2_X1 U12811 ( .A1(n12177), .A2(n21637), .ZN(n12178) );
  AND2_X1 U12812 ( .A1(n11906), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n11907) );
  NOR2_X1 U12813 ( .A1(n11777), .A2(n19982), .ZN(n11843) );
  AND2_X1 U12814 ( .A1(n11615), .A2(n13663), .ZN(n13471) );
  INV_X1 U12815 ( .A(n15823), .ZN(n15981) );
  NAND2_X1 U12816 ( .A1(n11703), .A2(n11702), .ZN(n11704) );
  OR2_X1 U12817 ( .A1(n11705), .A2(n11704), .ZN(n11706) );
  INV_X1 U12818 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n21864) );
  AOI21_X1 U12819 ( .B1(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n19200), .A(
        n13181), .ZN(n13183) );
  AND2_X1 U12820 ( .A1(n12864), .A2(n12863), .ZN(n12865) );
  OR2_X1 U12821 ( .A1(n13063), .A2(n19651), .ZN(n12857) );
  AND2_X1 U12822 ( .A1(n13411), .A2(n13410), .ZN(n16502) );
  INV_X1 U12823 ( .A(n13856), .ZN(n13855) );
  AND2_X1 U12824 ( .A1(n18548), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n16532) );
  OAI21_X1 U12825 ( .B1(n12828), .B2(n13554), .A(n19203), .ZN(n12853) );
  NAND2_X1 U12826 ( .A1(n16640), .A2(n18090), .ZN(n15011) );
  NAND2_X1 U12827 ( .A1(n17567), .A2(n20642), .ZN(n17568) );
  OR2_X1 U12828 ( .A1(n20808), .A2(n20806), .ZN(n14637) );
  NAND2_X1 U12829 ( .A1(n21563), .A2(P1_REIP_REG_18__SCAN_IN), .ZN(n21574) );
  AND2_X1 U12830 ( .A1(n11843), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11855) );
  NAND2_X1 U12831 ( .A1(n11812), .A2(n11811), .ZN(n13775) );
  NOR2_X1 U12832 ( .A1(n12139), .A2(n15757), .ZN(n12140) );
  NOR2_X1 U12833 ( .A1(n12059), .A2(n21573), .ZN(n12060) );
  AND2_X1 U12834 ( .A1(n12026), .A2(n12025), .ZN(n15561) );
  NAND2_X1 U12835 ( .A1(n15967), .A2(n21412), .ZN(n15938) );
  INV_X1 U12836 ( .A(n15970), .ZN(n21412) );
  OAI21_X1 U12837 ( .B1(n21684), .B2(n13902), .A(n16010), .ZN(n13904) );
  INV_X1 U12838 ( .A(n14407), .ZN(n14444) );
  INV_X1 U12839 ( .A(n22161), .ZN(n14248) );
  INV_X1 U12840 ( .A(n13901), .ZN(n14279) );
  NOR2_X1 U12841 ( .A1(n21862), .A2(n21771), .ZN(n21852) );
  NAND2_X1 U12842 ( .A1(n14157), .A2(n12388), .ZN(n14402) );
  AND2_X1 U12843 ( .A1(n13247), .A2(n21729), .ZN(n14039) );
  INV_X1 U12844 ( .A(n13924), .ZN(n15443) );
  OR2_X1 U12845 ( .A1(n12919), .A2(n12918), .ZN(n14222) );
  INV_X1 U12846 ( .A(n13887), .ZN(n13827) );
  AOI21_X1 U12847 ( .B1(n18526), .B2(n12856), .A(n12855), .ZN(n13645) );
  INV_X1 U12848 ( .A(n13100), .ZN(n13097) );
  INV_X1 U12849 ( .A(n13323), .ZN(n15463) );
  INV_X1 U12850 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n18282) );
  INV_X1 U12851 ( .A(n15489), .ZN(n15490) );
  OR2_X1 U12852 ( .A1(n15308), .A2(n16448), .ZN(n16290) );
  AND3_X1 U12853 ( .A1(n13338), .A2(n13337), .A3(n13336), .ZN(n14454) );
  INV_X1 U12854 ( .A(n18622), .ZN(n18594) );
  INV_X1 U12855 ( .A(n16667), .ZN(n16668) );
  OR2_X1 U12856 ( .A1(n14995), .A2(n13229), .ZN(n16640) );
  AND2_X1 U12857 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19232) );
  OR2_X1 U12858 ( .A1(n19328), .A2(n17077), .ZN(n19217) );
  NAND2_X1 U12859 ( .A1(n19152), .A2(n19151), .ZN(n19306) );
  NAND2_X1 U12860 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19331), .ZN(n19675) );
  INV_X1 U12861 ( .A(n21280), .ZN(n21250) );
  AOI22_X1 U12862 ( .A1(n10977), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n17505), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n14533) );
  INV_X1 U12863 ( .A(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n20293) );
  AOI221_X1 U12864 ( .B1(n17148), .B2(n17147), .C1(n21255), .C2(n17147), .A(
        n21310), .ZN(n20610) );
  AND2_X1 U12865 ( .A1(n20610), .A2(n20609), .ZN(n20611) );
  INV_X1 U12866 ( .A(n20950), .ZN(n21176) );
  INV_X1 U12867 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n21263) );
  OAI21_X1 U12868 ( .B1(n21301), .B2(n17531), .A(n16690), .ZN(n18684) );
  INV_X1 U12869 ( .A(n12532), .ZN(n15514) );
  OR2_X1 U12870 ( .A1(n15525), .A2(n19929), .ZN(n12643) );
  INV_X1 U12871 ( .A(n21571), .ZN(n21562) );
  NAND2_X1 U12872 ( .A1(n11817), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11777) );
  NAND2_X1 U12873 ( .A1(n21422), .A2(n21439), .ZN(n21639) );
  INV_X1 U12874 ( .A(n19969), .ZN(n15617) );
  NAND2_X1 U12875 ( .A1(n12378), .A2(n12381), .ZN(n15493) );
  INV_X1 U12876 ( .A(n14302), .ZN(n14395) );
  NAND2_X1 U12877 ( .A1(n14297), .A2(n14296), .ZN(n14398) );
  NAND2_X1 U12878 ( .A1(n12140), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n12177) );
  NAND2_X1 U12879 ( .A1(n12094), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n12139) );
  AND2_X1 U12880 ( .A1(n15099), .A2(n15098), .ZN(n19998) );
  INV_X1 U12881 ( .A(n21689), .ZN(n20029) );
  NOR2_X1 U12882 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n21881) );
  INV_X1 U12883 ( .A(n12503), .ZN(n15714) );
  OR2_X1 U12884 ( .A1(n21666), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12489) );
  AND2_X1 U12885 ( .A1(n13753), .A2(n13751), .ZN(n15970) );
  AOI21_X1 U12886 ( .B1(n13738), .B2(n13737), .A(n21689), .ZN(n13753) );
  AND2_X1 U12887 ( .A1(n13753), .A2(n16744), .ZN(n21416) );
  AND2_X1 U12888 ( .A1(n21787), .A2(n21855), .ZN(n22142) );
  AND2_X1 U12889 ( .A1(n12407), .A2(n14401), .ZN(n21787) );
  OAI211_X1 U12890 ( .C1(n21793), .C2(n21792), .A(n21852), .B(n21791), .ZN(
        n22149) );
  AND2_X1 U12891 ( .A1(n21787), .A2(n21888), .ZN(n22154) );
  AND2_X1 U12892 ( .A1(n21787), .A2(n21766), .ZN(n22155) );
  NOR2_X1 U12893 ( .A1(n14158), .A2(n14156), .ZN(n14407) );
  NOR2_X1 U12894 ( .A1(n14158), .A2(n21786), .ZN(n22162) );
  NOR2_X2 U12895 ( .A1(n14158), .A2(n14402), .ZN(n22169) );
  INV_X1 U12896 ( .A(n21836), .ZN(n21822) );
  NOR2_X2 U12897 ( .A1(n21836), .A2(n21786), .ZN(n22180) );
  NOR2_X1 U12898 ( .A1(n21836), .A2(n14402), .ZN(n22189) );
  NOR2_X1 U12899 ( .A1(n14157), .A2(n12388), .ZN(n21855) );
  NOR2_X2 U12900 ( .A1(n21885), .A2(n21884), .ZN(n22204) );
  INV_X1 U12901 ( .A(n22134), .ZN(n22213) );
  INV_X1 U12902 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n21321) );
  INV_X1 U12903 ( .A(n21675), .ZN(n21712) );
  AND2_X1 U12904 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n22221), .ZN(n19920) );
  AND2_X1 U12905 ( .A1(n13545), .A2(n13240), .ZN(n15030) );
  INV_X1 U12906 ( .A(n18502), .ZN(n18331) );
  CLKBUF_X1 U12907 ( .A(n18457), .Z(n18471) );
  NOR2_X1 U12908 ( .A1(n18331), .A2(n19203), .ZN(n18507) );
  OR2_X1 U12909 ( .A1(n12949), .A2(n12948), .ZN(n14494) );
  INV_X1 U12910 ( .A(n16167), .ZN(n16141) );
  XNOR2_X1 U12911 ( .A(n16120), .B(n13097), .ZN(n16116) );
  AND2_X1 U12912 ( .A1(n13249), .A2(n13248), .ZN(n19652) );
  INV_X1 U12913 ( .A(n19116), .ZN(n19668) );
  INV_X1 U12914 ( .A(n19116), .ZN(n19556) );
  INV_X1 U12915 ( .A(n16226), .ZN(n16679) );
  AND2_X1 U12916 ( .A1(n17022), .A2(n13506), .ZN(n17055) );
  AND2_X1 U12917 ( .A1(n18653), .A2(n19605), .ZN(n17047) );
  INV_X1 U12918 ( .A(n16117), .ZN(n18416) );
  INV_X1 U12919 ( .A(n18591), .ZN(n18605) );
  OR2_X1 U12920 ( .A1(n15256), .A2(n15255), .ZN(n18547) );
  AND2_X1 U12921 ( .A1(n15012), .A2(n18099), .ZN(n15049) );
  INV_X1 U12922 ( .A(n18606), .ZN(n18598) );
  INV_X1 U12923 ( .A(n19775), .ZN(n19779) );
  OR2_X1 U12924 ( .A1(n19168), .A2(n19151), .ZN(n19266) );
  INV_X1 U12925 ( .A(n19755), .ZN(n19757) );
  OAI21_X1 U12926 ( .B1(n19290), .B2(n19289), .A(n19288), .ZN(n19751) );
  NOR2_X2 U12927 ( .A1(n19267), .A2(n19266), .ZN(n19750) );
  NOR2_X1 U12928 ( .A1(n19267), .A2(n19293), .ZN(n19731) );
  INV_X1 U12929 ( .A(n19735), .ZN(n19625) );
  NOR2_X2 U12930 ( .A1(n19217), .A2(n19266), .ZN(n19724) );
  INV_X1 U12931 ( .A(n19422), .ZN(n19707) );
  NOR2_X1 U12932 ( .A1(n19278), .A2(n19217), .ZN(n19368) );
  NOR2_X1 U12933 ( .A1(n19169), .A2(n19266), .ZN(n19701) );
  INV_X1 U12934 ( .A(n19594), .ZN(n19598) );
  NAND2_X1 U12935 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_STATE2_REG_2__SCAN_IN), .ZN(n17064) );
  INV_X1 U12936 ( .A(P2_STATE_REG_1__SCAN_IN), .ZN(n21728) );
  INV_X1 U12937 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n21758) );
  AND2_X1 U12938 ( .A1(n20581), .A2(n20580), .ZN(n20595) );
  NAND3_X1 U12939 ( .A1(n14533), .A2(n14532), .A3(n14531), .ZN(n20171) );
  INV_X1 U12940 ( .A(n20507), .ZN(n20600) );
  NOR2_X1 U12941 ( .A1(n20167), .A2(n20169), .ZN(n20507) );
  NOR2_X2 U12942 ( .A1(n20513), .A2(n21296), .ZN(n20585) );
  NOR2_X1 U12943 ( .A1(n20711), .A2(n17415), .ZN(n17445) );
  AND2_X1 U12944 ( .A1(n17524), .A2(n17516), .ZN(n17489) );
  OR2_X1 U12945 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), .ZN(
        n20179) );
  NOR2_X1 U12946 ( .A1(n20694), .A2(n20699), .ZN(n20693) );
  NOR2_X1 U12947 ( .A1(n20112), .A2(n16712), .ZN(n18019) );
  NOR2_X1 U12948 ( .A1(n21707), .A2(n20112), .ZN(n20612) );
  INV_X1 U12949 ( .A(n20154), .ZN(n20159) );
  NOR2_X1 U12950 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n21296), .ZN(
        n21300) );
  INV_X1 U12951 ( .A(n19063), .ZN(n19076) );
  INV_X1 U12952 ( .A(n19045), .ZN(n19059) );
  INV_X1 U12953 ( .A(n19039), .ZN(n19053) );
  INV_X1 U12954 ( .A(n19027), .ZN(n19041) );
  INV_X1 U12955 ( .A(n19021), .ZN(n19035) );
  INV_X1 U12956 ( .A(n18998), .ZN(n19002) );
  NOR2_X1 U12957 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n21309), .ZN(n21290) );
  INV_X1 U12958 ( .A(n21755), .ZN(n21707) );
  INV_X1 U12959 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n21706) );
  OAI21_X1 U12960 ( .B1(n13260), .B2(n13259), .A(P2_ADDRESS_REG_29__SCAN_IN), 
        .ZN(n16226) );
  AND2_X1 U12961 ( .A1(n13735), .A2(n13451), .ZN(n14297) );
  NAND2_X1 U12962 ( .A1(n21490), .A2(n21488), .ZN(n21507) );
  NAND2_X1 U12963 ( .A1(n21422), .A2(n12518), .ZN(n21648) );
  NAND2_X1 U12964 ( .A1(n21422), .A2(n13953), .ZN(n21642) );
  NAND2_X1 U12965 ( .A1(n19969), .A2(n13662), .ZN(n15628) );
  INV_X1 U12966 ( .A(n19962), .ZN(n19966) );
  INV_X1 U12967 ( .A(n19998), .ZN(n21519) );
  INV_X1 U12968 ( .A(n19854), .ZN(n19885) );
  INV_X1 U12969 ( .A(n14398), .ZN(n14302) );
  NAND2_X1 U12970 ( .A1(n12485), .A2(n20024), .ZN(n12492) );
  INV_X1 U12971 ( .A(n20005), .ZN(n20028) );
  INV_X1 U12972 ( .A(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n19982) );
  OR2_X1 U12973 ( .A1(n12489), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n21386) );
  NAND2_X1 U12974 ( .A1(n13753), .A2(n13743), .ZN(n21353) );
  INV_X1 U12975 ( .A(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n16773) );
  INV_X1 U12976 ( .A(n21661), .ZN(n21663) );
  AOI22_X1 U12977 ( .A1(n21774), .A2(n21772), .B1(n21776), .B2(n21845), .ZN(
        n22139) );
  NAND2_X1 U12978 ( .A1(n21787), .A2(n21779), .ZN(n22146) );
  AOI22_X1 U12979 ( .A1(n21790), .A2(n21792), .B1(n21812), .B2(n21845), .ZN(
        n22152) );
  INV_X1 U12980 ( .A(n21799), .ZN(n22159) );
  NOR2_X1 U12981 ( .A1(n14406), .A2(n21814), .ZN(n14448) );
  INV_X1 U12982 ( .A(n14155), .ZN(n14252) );
  AOI22_X1 U12983 ( .A1(n21813), .A2(n21818), .B1(n21862), .B2(n21812), .ZN(
        n22166) );
  INV_X1 U12984 ( .A(n22162), .ZN(n14283) );
  NAND2_X1 U12985 ( .A1(n21822), .A2(n21855), .ZN(n22178) );
  AOI22_X1 U12986 ( .A1(n21850), .A2(n21847), .B1(n21845), .B2(n21844), .ZN(
        n22185) );
  NOR2_X1 U12987 ( .A1(n14123), .A2(n14122), .ZN(n14273) );
  INV_X1 U12988 ( .A(n22058), .ZN(n22050) );
  NAND2_X1 U12989 ( .A1(n21889), .A2(n21855), .ZN(n22200) );
  NAND2_X1 U12990 ( .A1(n21889), .A2(n21888), .ZN(n22218) );
  INV_X1 U12991 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n21868) );
  INV_X1 U12992 ( .A(n19917), .ZN(n19928) );
  NOR2_X1 U12993 ( .A1(n14040), .A2(n18649), .ZN(n18095) );
  OR2_X1 U12994 ( .A1(n16026), .A2(n16025), .ZN(n18453) );
  INV_X1 U12995 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n18265) );
  INV_X1 U12996 ( .A(n16102), .ZN(n16157) );
  AND2_X1 U12997 ( .A1(n13649), .A2(n18099), .ZN(n16102) );
  XNOR2_X1 U12998 ( .A(n13666), .B(n13665), .ZN(n19219) );
  INV_X2 U12999 ( .A(n19652), .ZN(n19401) );
  AND2_X1 U13000 ( .A1(n19659), .A2(n19658), .ZN(n19410) );
  NAND2_X1 U13001 ( .A1(n19401), .A2(n13250), .ZN(n19659) );
  NAND2_X1 U13002 ( .A1(n17095), .A2(n12760), .ZN(n13808) );
  INV_X1 U13003 ( .A(n17095), .ZN(n17128) );
  NAND2_X1 U13004 ( .A1(n13449), .A2(n19605), .ZN(n16026) );
  NAND2_X2 U13005 ( .A1(n13449), .A2(n13448), .ZN(n19670) );
  INV_X1 U13006 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n17023) );
  OR2_X1 U13007 ( .A1(n18653), .A2(n13495), .ZN(n17022) );
  NAND2_X1 U13008 ( .A1(n15049), .A2(n15029), .ZN(n18606) );
  INV_X1 U13009 ( .A(n18568), .ZN(n18617) );
  INV_X1 U13010 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19231) );
  AOI21_X1 U13011 ( .B1(n16672), .B2(n16671), .A(n19673), .ZN(n19788) );
  OR2_X1 U13012 ( .A1(n19315), .A2(n19266), .ZN(n19775) );
  INV_X1 U13013 ( .A(n19494), .ZN(n19767) );
  OR2_X1 U13014 ( .A1(n19315), .A2(n19278), .ZN(n19755) );
  AOI21_X1 U13015 ( .B1(n19269), .B2(n19273), .A(n19265), .ZN(n19748) );
  AND2_X1 U13016 ( .A1(n19256), .A2(n19255), .ZN(n19631) );
  INV_X1 U13017 ( .A(n19731), .ZN(n19741) );
  INV_X1 U13018 ( .A(n19724), .ZN(n19577) );
  OR2_X1 U13019 ( .A1(n19267), .A2(n19278), .ZN(n19735) );
  NOR2_X1 U13020 ( .A1(n19216), .A2(n19215), .ZN(n19722) );
  AOI21_X1 U13021 ( .B1(n19207), .B2(n19209), .A(n19202), .ZN(n19716) );
  AND2_X1 U13022 ( .A1(n19192), .A2(n19191), .ZN(n19422) );
  INV_X1 U13023 ( .A(n19368), .ZN(n19710) );
  INV_X1 U13024 ( .A(n19437), .ZN(n19452) );
  INV_X1 U13025 ( .A(n16677), .ZN(n19532) );
  NAND2_X1 U13026 ( .A1(n16664), .A2(n16663), .ZN(n19562) );
  AND2_X1 U13027 ( .A1(n19144), .A2(n19143), .ZN(n19610) );
  INV_X1 U13028 ( .A(n21698), .ZN(n17093) );
  INV_X2 U13029 ( .A(n17143), .ZN(n21734) );
  INV_X1 U13030 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n21700) );
  NAND4_X1 U13031 ( .A1(n20172), .A2(P3_EBX_REG_31__SCAN_IN), .A3(n20171), 
        .A4(n20170), .ZN(n20554) );
  INV_X1 U13032 ( .A(n20585), .ZN(n20558) );
  INV_X1 U13033 ( .A(n20604), .ZN(n20561) );
  NOR2_X1 U13034 ( .A1(n20515), .A2(n17429), .ZN(n17434) );
  INV_X1 U13035 ( .A(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17453) );
  AND2_X1 U13036 ( .A1(n17524), .A2(n20711), .ZN(n17526) );
  NOR2_X1 U13037 ( .A1(n20668), .A2(n20632), .ZN(n20636) );
  INV_X1 U13038 ( .A(n20785), .ZN(n20776) );
  NAND2_X1 U13039 ( .A1(n20795), .A2(n20686), .ZN(n20781) );
  INV_X1 U13040 ( .A(n18019), .ZN(n18018) );
  NAND2_X1 U13041 ( .A1(n20111), .A2(n20612), .ZN(n20154) );
  INV_X1 U13042 ( .A(n20152), .ZN(n20161) );
  INV_X1 U13043 ( .A(n17886), .ZN(n17876) );
  INV_X1 U13044 ( .A(n17577), .ZN(n17970) );
  INV_X1 U13045 ( .A(n21203), .ZN(n21246) );
  INV_X1 U13046 ( .A(n21133), .ZN(n21220) );
  INV_X1 U13047 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18692) );
  INV_X1 U13048 ( .A(n19090), .ZN(n19080) );
  INV_X1 U13049 ( .A(n19081), .ZN(n19111) );
  INV_X1 U13050 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n21309) );
  INV_X1 U13051 ( .A(n21703), .ZN(n16707) );
  INV_X1 U13052 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n20250) );
  NOR2_X1 U13053 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n13442), .ZN(n18966)
         );
  INV_X1 U13054 ( .A(n19850), .ZN(n19839) );
  AND2_X2 U13055 ( .A1(n13622), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13615) );
  AOI22_X1 U13056 ( .A1(n10951), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11676), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11498) );
  AND2_X2 U13057 ( .A1(n13615), .A2(n16011), .ZN(n11641) );
  AOI22_X1 U13058 ( .A1(n11641), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11540), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11497) );
  AND2_X2 U13059 ( .A1(n13613), .A2(n11494), .ZN(n11997) );
  AOI22_X1 U13060 ( .A1(n11584), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n11997), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11496) );
  AOI22_X1 U13061 ( .A1(n10955), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11585), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11495) );
  AOI22_X1 U13062 ( .A1(n11979), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11878), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11504) );
  BUF_X4 U13063 ( .A(n11537), .Z(n12197) );
  AOI22_X1 U13064 ( .A1(n12197), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n11554), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11503) );
  AOI22_X1 U13065 ( .A1(n11653), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n11834), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11502) );
  AND2_X2 U13066 ( .A1(n13615), .A2(n13587), .ZN(n11545) );
  AND2_X2 U13067 ( .A1(n11500), .A2(n16011), .ZN(n11963) );
  AOI22_X1 U13068 ( .A1(n11545), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11963), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11501) );
  NAND2_X2 U13069 ( .A1(n11506), .A2(n11505), .ZN(n12357) );
  AOI22_X1 U13070 ( .A1(n11653), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11554), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11509) );
  AOI22_X1 U13071 ( .A1(n11834), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11997), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11508) );
  AOI22_X1 U13072 ( .A1(n11878), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11963), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11507) );
  NAND4_X1 U13073 ( .A1(n11510), .A2(n11509), .A3(n11508), .A4(n11507), .ZN(
        n11516) );
  AOI22_X1 U13074 ( .A1(n12096), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11540), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11514) );
  AOI22_X1 U13075 ( .A1(n10955), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11585), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11513) );
  AOI22_X1 U13076 ( .A1(n11545), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11584), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11512) );
  AOI22_X1 U13077 ( .A1(n10954), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11676), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11511) );
  NAND4_X1 U13078 ( .A1(n11514), .A2(n11513), .A3(n11512), .A4(n11511), .ZN(
        n11515) );
  OR2_X2 U13079 ( .A1(n11516), .A2(n11515), .ZN(n11611) );
  NAND2_X1 U13080 ( .A1(n11878), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n11520) );
  NAND2_X1 U13081 ( .A1(n11676), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n11519) );
  NAND2_X1 U13082 ( .A1(n10956), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n11518) );
  NAND2_X1 U13083 ( .A1(n11653), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n11517) );
  NAND2_X1 U13084 ( .A1(n10953), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n11524) );
  NAND2_X1 U13085 ( .A1(n11979), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n11523) );
  NAND2_X1 U13086 ( .A1(n11540), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n11522) );
  NAND2_X1 U13087 ( .A1(n11834), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n11521) );
  NAND2_X1 U13088 ( .A1(n12197), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n11528) );
  NAND2_X1 U13089 ( .A1(n11545), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n11527) );
  NAND2_X1 U13090 ( .A1(n11554), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n11526) );
  NAND2_X1 U13091 ( .A1(n11963), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n11525) );
  NAND2_X1 U13092 ( .A1(n12269), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n11532) );
  NAND2_X1 U13093 ( .A1(n11585), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n11531) );
  NAND2_X1 U13094 ( .A1(n11997), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n11530) );
  NAND2_X1 U13095 ( .A1(n11584), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n11529) );
  AOI22_X1 U13096 ( .A1(n11878), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11963), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11544) );
  NAND2_X1 U13097 ( .A1(n11962), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(
        n11539) );
  NAND2_X1 U13098 ( .A1(n11554), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n11538) );
  AND2_X1 U13099 ( .A1(n11539), .A2(n11538), .ZN(n11543) );
  AOI22_X1 U13100 ( .A1(n11979), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11585), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11542) );
  AOI22_X1 U13101 ( .A1(n11653), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n11540), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11541) );
  AOI22_X1 U13102 ( .A1(n11676), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11834), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11549) );
  AOI22_X1 U13103 ( .A1(n12096), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11545), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11548) );
  AOI22_X1 U13104 ( .A1(n10951), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n10956), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11547) );
  AOI22_X1 U13105 ( .A1(n11584), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n11997), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11546) );
  AOI22_X1 U13106 ( .A1(n10952), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11676), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11553) );
  AOI22_X1 U13107 ( .A1(n12096), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11540), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11552) );
  AOI22_X1 U13108 ( .A1(n11584), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n11997), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11551) );
  AOI22_X1 U13109 ( .A1(n10955), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11585), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11550) );
  NAND4_X1 U13110 ( .A1(n11553), .A2(n11552), .A3(n11551), .A4(n11550), .ZN(
        n11560) );
  AOI22_X1 U13111 ( .A1(n11979), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11878), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11558) );
  AOI22_X1 U13112 ( .A1(n11962), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n11554), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11557) );
  AOI22_X1 U13113 ( .A1(n11653), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n11834), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11556) );
  AOI22_X1 U13114 ( .A1(n11545), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11963), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11555) );
  NAND4_X1 U13115 ( .A1(n11558), .A2(n11557), .A3(n11556), .A4(n11555), .ZN(
        n11559) );
  AND2_X2 U13116 ( .A1(n14182), .A2(n12384), .ZN(n11615) );
  AOI22_X1 U13117 ( .A1(n11962), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n11540), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11564) );
  AOI22_X1 U13118 ( .A1(n10951), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n10956), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11563) );
  AOI22_X1 U13119 ( .A1(n11545), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n10974), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11562) );
  AOI22_X1 U13120 ( .A1(n12096), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11585), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11561) );
  NAND4_X1 U13121 ( .A1(n11564), .A2(n11563), .A3(n11562), .A4(n11561), .ZN(
        n11570) );
  AOI22_X1 U13122 ( .A1(n11676), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n11554), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11568) );
  AOI22_X1 U13123 ( .A1(n11878), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n11963), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11567) );
  AOI22_X1 U13124 ( .A1(n11979), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11834), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11566) );
  AOI22_X1 U13125 ( .A1(n11653), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n11997), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11565) );
  NAND4_X1 U13126 ( .A1(n11568), .A2(n11567), .A3(n11566), .A4(n11565), .ZN(
        n11569) );
  NAND2_X1 U13127 ( .A1(n11676), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n11575) );
  NAND2_X1 U13128 ( .A1(n10954), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n11574) );
  NAND2_X1 U13129 ( .A1(n12269), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n11573) );
  NAND2_X1 U13130 ( .A1(n11540), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n11572) );
  NAND2_X1 U13131 ( .A1(n11979), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n11579) );
  NAND2_X1 U13132 ( .A1(n11878), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n11578) );
  NAND2_X1 U13133 ( .A1(n11545), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n11577) );
  NAND2_X1 U13134 ( .A1(n11963), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n11576) );
  NAND2_X1 U13135 ( .A1(n11653), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n11583) );
  NAND2_X1 U13136 ( .A1(n12197), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n11582) );
  NAND2_X1 U13137 ( .A1(n11554), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n11581) );
  NAND2_X1 U13138 ( .A1(n11834), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n11580) );
  NAND2_X1 U13139 ( .A1(n10955), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n11589) );
  NAND2_X1 U13140 ( .A1(n11584), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n11588) );
  NAND2_X1 U13141 ( .A1(n11997), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n11587) );
  NAND4_X4 U13142 ( .A1(n11593), .A2(n11592), .A3(n11591), .A4(n11590), .ZN(
        n13747) );
  AOI22_X1 U13143 ( .A1(n10952), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n10956), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11597) );
  AOI22_X1 U13144 ( .A1(n11979), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11545), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11596) );
  AOI22_X1 U13145 ( .A1(n11878), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n11584), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11595) );
  AOI22_X1 U13146 ( .A1(n11676), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n11834), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11594) );
  NAND4_X1 U13147 ( .A1(n11597), .A2(n11596), .A3(n11595), .A4(n11594), .ZN(
        n11603) );
  AOI22_X1 U13148 ( .A1(n11540), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11554), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11601) );
  AOI22_X1 U13149 ( .A1(n11962), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n11963), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11600) );
  AOI22_X1 U13150 ( .A1(n12096), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n11997), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11599) );
  AOI22_X1 U13151 ( .A1(n11653), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n11585), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11598) );
  NAND4_X1 U13152 ( .A1(n11601), .A2(n11600), .A3(n11599), .A4(n11598), .ZN(
        n11602) );
  NAND2_X1 U13153 ( .A1(n21725), .A2(P1_STATE_REG_1__SCAN_IN), .ZN(n21711) );
  INV_X1 U13154 ( .A(P1_STATE_REG_1__SCAN_IN), .ZN(n11604) );
  NAND2_X1 U13155 ( .A1(n11604), .A2(P1_STATE_REG_2__SCAN_IN), .ZN(n11605) );
  NAND2_X1 U13156 ( .A1(n21711), .A2(n11605), .ZN(n12520) );
  NAND2_X1 U13157 ( .A1(n13662), .A2(n11640), .ZN(n11622) );
  NAND2_X1 U13158 ( .A1(n11614), .A2(n11622), .ZN(n11609) );
  NAND3_X1 U13159 ( .A1(n14182), .A2(n11611), .A3(n12357), .ZN(n11608) );
  NAND2_X1 U13160 ( .A1(n13634), .A2(n12384), .ZN(n11630) );
  AND2_X2 U13161 ( .A1(n11610), .A2(n11630), .ZN(n11619) );
  NOR2_X1 U13162 ( .A1(n13570), .A2(n13747), .ZN(n11612) );
  NAND2_X1 U13163 ( .A1(n13584), .A2(n13568), .ZN(n13739) );
  INV_X1 U13164 ( .A(n11615), .ZN(n11616) );
  NAND2_X1 U13165 ( .A1(n13570), .A2(n11617), .ZN(n11618) );
  AND2_X2 U13166 ( .A1(n11619), .A2(n11618), .ZN(n11628) );
  NAND2_X1 U13167 ( .A1(n11148), .A2(n12357), .ZN(n11620) );
  INV_X1 U13168 ( .A(n13634), .ZN(n13579) );
  NAND2_X1 U13169 ( .A1(n16772), .A2(n21868), .ZN(n21666) );
  XNOR2_X1 U13170 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n21823) );
  OR2_X1 U13171 ( .A1(n16766), .A2(n21864), .ZN(n11692) );
  OAI21_X1 U13172 ( .B1(n12489), .B2(n21823), .A(n11692), .ZN(n11623) );
  INV_X1 U13173 ( .A(n11623), .ZN(n11624) );
  INV_X1 U13174 ( .A(n16766), .ZN(n11722) );
  MUX2_X1 U13175 ( .A(n11722), .B(n11723), .S(n21877), .Z(n11626) );
  NAND3_X1 U13176 ( .A1(n13581), .A2(n13732), .A3(n16740), .ZN(n11635) );
  INV_X1 U13177 ( .A(n11628), .ZN(n11629) );
  OAI21_X1 U13178 ( .B1(n13460), .B2(n11630), .A(n11629), .ZN(n11634) );
  NAND2_X1 U13179 ( .A1(n11613), .A2(n11631), .ZN(n13746) );
  OR2_X1 U13180 ( .A1(n21666), .A2(n21321), .ZN(n20033) );
  AOI21_X1 U13181 ( .B1(n11617), .B2(n13747), .A(n20033), .ZN(n11632) );
  NAND4_X1 U13182 ( .A1(n11636), .A2(n11635), .A3(n11634), .A4(n11633), .ZN(
        n11669) );
  NAND2_X1 U13183 ( .A1(n11671), .A2(n11669), .ZN(n11638) );
  INV_X1 U13184 ( .A(n11638), .ZN(n11637) );
  NAND2_X1 U13185 ( .A1(n11639), .A2(n11638), .ZN(n14151) );
  INV_X1 U13186 ( .A(n11708), .ZN(n11684) );
  AOI22_X1 U13187 ( .A1(n10955), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12096), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11645) );
  AOI22_X1 U13188 ( .A1(n11878), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12197), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11644) );
  AOI22_X1 U13189 ( .A1(n10953), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12264), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11643) );
  AOI22_X1 U13190 ( .A1(n11979), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11963), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11642) );
  NAND4_X1 U13191 ( .A1(n11645), .A2(n11644), .A3(n11643), .A4(n11642), .ZN(
        n11651) );
  AOI22_X1 U13192 ( .A1(n12247), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n11545), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11649) );
  AOI22_X1 U13193 ( .A1(n12127), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n11968), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11648) );
  AOI22_X1 U13194 ( .A1(n12263), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n12218), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11647) );
  NAND4_X1 U13195 ( .A1(n11649), .A2(n11648), .A3(n11647), .A4(n11646), .ZN(
        n11650) );
  NAND2_X1 U13196 ( .A1(n11684), .A2(n12396), .ZN(n11652) );
  AOI22_X1 U13197 ( .A1(n10953), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12223), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11657) );
  AOI22_X1 U13198 ( .A1(n12247), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n11545), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11656) );
  AOI22_X1 U13199 ( .A1(n12127), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12263), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11655) );
  NAND4_X1 U13200 ( .A1(n11657), .A2(n11656), .A3(n11655), .A4(n11654), .ZN(
        n11663) );
  AOI22_X1 U13201 ( .A1(n10955), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12096), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11661) );
  AOI22_X1 U13202 ( .A1(n11979), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12218), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11660) );
  AOI22_X1 U13203 ( .A1(n12264), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n11963), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11659) );
  AOI22_X1 U13204 ( .A1(n11962), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n12270), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11658) );
  NAND4_X1 U13205 ( .A1(n11661), .A2(n11660), .A3(n11659), .A4(n11658), .ZN(
        n11662) );
  NAND2_X1 U13206 ( .A1(n12302), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11666) );
  INV_X1 U13207 ( .A(n11707), .ZN(n11664) );
  NAND2_X1 U13208 ( .A1(n11664), .A2(n12396), .ZN(n11665) );
  OAI211_X1 U13209 ( .C1(n11708), .C2(n12453), .A(n11666), .B(n11665), .ZN(
        n11667) );
  INV_X1 U13210 ( .A(n11669), .ZN(n11670) );
  AOI22_X1 U13211 ( .A1(n10956), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12247), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11675) );
  AOI22_X1 U13212 ( .A1(n11979), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12197), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11674) );
  AOI22_X1 U13213 ( .A1(n12264), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n12218), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11673) );
  AOI22_X1 U13214 ( .A1(n12271), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11963), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11672) );
  NAND4_X1 U13215 ( .A1(n11675), .A2(n11674), .A3(n11673), .A4(n11672), .ZN(
        n11682) );
  AOI22_X1 U13216 ( .A1(n12127), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12096), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11680) );
  AOI22_X1 U13217 ( .A1(n11878), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12263), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11679) );
  AOI22_X1 U13218 ( .A1(n11585), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n11968), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11678) );
  AOI22_X1 U13219 ( .A1(n10953), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12270), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11677) );
  NAND4_X1 U13220 ( .A1(n11680), .A2(n11679), .A3(n11678), .A4(n11677), .ZN(
        n11681) );
  INV_X1 U13221 ( .A(n12395), .ZN(n11683) );
  XNOR2_X1 U13222 ( .A(n11683), .B(n12453), .ZN(n11685) );
  NAND2_X1 U13223 ( .A1(n11685), .A2(n11684), .ZN(n11686) );
  INV_X1 U13224 ( .A(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11689) );
  AOI21_X1 U13225 ( .B1(n14173), .B2(n12453), .A(n21321), .ZN(n11688) );
  NAND2_X1 U13226 ( .A1(n13905), .A2(n12395), .ZN(n11687) );
  OAI211_X1 U13227 ( .C1(n12333), .C2(n11689), .A(n11688), .B(n11687), .ZN(
        n11793) );
  INV_X1 U13228 ( .A(n12453), .ZN(n11690) );
  NOR2_X1 U13229 ( .A1(n11690), .A2(n11708), .ZN(n12450) );
  INV_X1 U13230 ( .A(n11692), .ZN(n11694) );
  OAI21_X1 U13231 ( .B1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n11694), .A(
        n11693), .ZN(n11695) );
  NAND2_X1 U13232 ( .A1(n11696), .A2(n11695), .ZN(n11705) );
  NAND2_X1 U13233 ( .A1(n11697), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11703) );
  NAND2_X1 U13234 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n21916) );
  INV_X1 U13235 ( .A(n21916), .ZN(n21909) );
  NAND2_X1 U13236 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21909), .ZN(
        n21905) );
  INV_X1 U13237 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n11700) );
  OR2_X1 U13238 ( .A1(n21864), .A2(n21877), .ZN(n11698) );
  NAND2_X1 U13239 ( .A1(n11700), .A2(n11698), .ZN(n11699) );
  NOR2_X1 U13240 ( .A1(n16766), .A2(n11700), .ZN(n11701) );
  AOI21_X1 U13241 ( .B1(n14408), .B2(n11723), .A(n11701), .ZN(n11702) );
  NAND2_X2 U13242 ( .A1(n11705), .A2(n11704), .ZN(n13979) );
  OR2_X2 U13244 ( .A1(n21860), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11720) );
  AOI22_X1 U13245 ( .A1(n10954), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11545), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11712) );
  AOI22_X1 U13246 ( .A1(n10956), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12269), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11711) );
  AOI22_X1 U13247 ( .A1(n11979), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12223), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11710) );
  AOI22_X1 U13248 ( .A1(n12263), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n12270), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11709) );
  NAND4_X1 U13249 ( .A1(n11712), .A2(n11711), .A3(n11710), .A4(n11709), .ZN(
        n11718) );
  AOI22_X1 U13250 ( .A1(n11962), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n11963), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11716) );
  AOI22_X1 U13251 ( .A1(n12247), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12218), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11715) );
  AOI22_X1 U13252 ( .A1(n12127), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n11968), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11714) );
  AOI22_X1 U13253 ( .A1(n12264), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n11585), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11713) );
  NAND4_X1 U13254 ( .A1(n11716), .A2(n11715), .A3(n11714), .A4(n11713), .ZN(
        n11717) );
  AOI22_X1 U13255 ( .A1(n12343), .A2(n12383), .B1(n12302), .B2(
        P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11719) );
  NAND2_X2 U13256 ( .A1(n11720), .A2(n11719), .ZN(n11803) );
  NAND2_X1 U13257 ( .A1(n11697), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11725) );
  NAND2_X1 U13258 ( .A1(n21905), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n11721) );
  NOR2_X1 U13259 ( .A1(n21905), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n13901) );
  NAND2_X1 U13260 ( .A1(n11721), .A2(n14279), .ZN(n21824) );
  AOI22_X1 U13261 ( .A1(n21824), .A2(n11723), .B1(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n11722), .ZN(n11724) );
  XNOR2_X2 U13262 ( .A(n13979), .B(n13978), .ZN(n21769) );
  AOI22_X1 U13263 ( .A1(n10951), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12127), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11729) );
  AOI22_X1 U13264 ( .A1(n12096), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12263), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11728) );
  AOI22_X1 U13265 ( .A1(n12218), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n11968), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11727) );
  NAND4_X1 U13266 ( .A1(n11729), .A2(n11728), .A3(n11727), .A4(n11726), .ZN(
        n11735) );
  AOI22_X1 U13267 ( .A1(n11979), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12223), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11733) );
  AOI22_X1 U13268 ( .A1(n11962), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n12264), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11732) );
  AOI22_X1 U13269 ( .A1(n12247), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12270), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11731) );
  AOI22_X1 U13270 ( .A1(n12271), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12101), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11730) );
  NAND4_X1 U13271 ( .A1(n11733), .A2(n11732), .A3(n11731), .A4(n11730), .ZN(
        n11734) );
  AOI22_X1 U13272 ( .A1(n12343), .A2(n12411), .B1(n12302), .B2(
        P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11736) );
  AOI22_X1 U13273 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n12127), .B1(
        n12269), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11741) );
  AOI22_X1 U13274 ( .A1(n10952), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12247), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11740) );
  AOI22_X1 U13275 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n12263), .B1(
        n12101), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11738) );
  NAND4_X1 U13276 ( .A1(n11741), .A2(n11740), .A3(n11739), .A4(n11738), .ZN(
        n11747) );
  AOI22_X1 U13277 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n12223), .B1(
        n11545), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11745) );
  AOI22_X1 U13278 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n12197), .B1(
        n12264), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11744) );
  AOI22_X1 U13279 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n11979), .B1(
        n12218), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11743) );
  AOI22_X1 U13280 ( .A1(n10955), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12270), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11742) );
  NAND4_X1 U13281 ( .A1(n11745), .A2(n11744), .A3(n11743), .A4(n11742), .ZN(
        n11746) );
  NAND2_X1 U13282 ( .A1(n12343), .A2(n12424), .ZN(n11749) );
  NAND2_X1 U13283 ( .A1(n12302), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n11748) );
  NAND2_X1 U13284 ( .A1(n11749), .A2(n11748), .ZN(n11771) );
  AOI22_X1 U13285 ( .A1(n10953), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12127), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11753) );
  AOI22_X1 U13286 ( .A1(n12096), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12263), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11752) );
  AOI22_X1 U13287 ( .A1(n12218), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11968), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11751) );
  AOI22_X1 U13288 ( .A1(n10955), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11585), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11750) );
  NAND4_X1 U13289 ( .A1(n11753), .A2(n11752), .A3(n11751), .A4(n11750), .ZN(
        n11759) );
  AOI22_X1 U13290 ( .A1(n11979), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11878), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11757) );
  AOI22_X1 U13291 ( .A1(n11962), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n12264), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11756) );
  AOI22_X1 U13292 ( .A1(n12247), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12270), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11755) );
  AOI22_X1 U13293 ( .A1(n12271), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12101), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11754) );
  NAND4_X1 U13294 ( .A1(n11757), .A2(n11756), .A3(n11755), .A4(n11754), .ZN(
        n11758) );
  NAND2_X1 U13295 ( .A1(n12343), .A2(n12427), .ZN(n11761) );
  NAND2_X1 U13296 ( .A1(n12302), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n11760) );
  NAND2_X1 U13297 ( .A1(n11763), .A2(n11762), .ZN(n11764) );
  AND2_X2 U13298 ( .A1(n11848), .A2(n11764), .ZN(n12423) );
  INV_X1 U13299 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n11769) );
  INV_X1 U13300 ( .A(n11818), .ZN(n11765) );
  AND2_X1 U13301 ( .A1(n11777), .A2(n19982), .ZN(n11766) );
  OR2_X1 U13302 ( .A1(n11766), .A2(n11843), .ZN(n21447) );
  NOR2_X1 U13303 ( .A1(n12023), .A2(n19982), .ZN(n11767) );
  AOI21_X1 U13304 ( .B1(n21447), .B2(n12291), .A(n11767), .ZN(n11768) );
  OAI21_X1 U13305 ( .B1(n11822), .B2(n11769), .A(n11768), .ZN(n11770) );
  AOI21_X1 U13306 ( .B1(n12423), .B2(n11991), .A(n11770), .ZN(n14254) );
  INV_X1 U13307 ( .A(n14254), .ZN(n11782) );
  XNOR2_X1 U13308 ( .A(n11816), .B(n11771), .ZN(n12416) );
  NAND2_X1 U13309 ( .A1(n13568), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n11825) );
  INV_X1 U13310 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n11775) );
  NAND2_X1 U13311 ( .A1(n21910), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11774) );
  NAND2_X1 U13312 ( .A1(n12285), .A2(P1_EAX_REG_4__SCAN_IN), .ZN(n11773) );
  OAI211_X1 U13313 ( .C1(n11825), .C2(n11775), .A(n11774), .B(n11773), .ZN(
        n11776) );
  INV_X1 U13314 ( .A(n12291), .ZN(n11799) );
  NAND2_X1 U13315 ( .A1(n11776), .A2(n11799), .ZN(n11779) );
  OAI21_X1 U13316 ( .B1(n11817), .B2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n11777), .ZN(n21444) );
  NAND2_X1 U13317 ( .A1(n21444), .A2(n12291), .ZN(n11778) );
  NAND2_X1 U13318 ( .A1(n11779), .A2(n11778), .ZN(n11780) );
  AOI21_X1 U13319 ( .B1(n12416), .B2(n11991), .A(n11780), .ZN(n14205) );
  INV_X1 U13320 ( .A(n14205), .ZN(n11781) );
  NAND2_X1 U13321 ( .A1(n11782), .A2(n11781), .ZN(n11829) );
  INV_X1 U13322 ( .A(n11784), .ZN(n11785) );
  NAND2_X1 U13323 ( .A1(n11786), .A2(n11785), .ZN(n11787) );
  NAND2_X1 U13324 ( .A1(n14157), .A2(n11991), .ZN(n11792) );
  AOI22_X1 U13325 ( .A1(n11772), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n21910), .ZN(n11790) );
  INV_X1 U13326 ( .A(n11825), .ZN(n11788) );
  NAND2_X1 U13327 ( .A1(n11788), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11789) );
  AND2_X1 U13328 ( .A1(n11790), .A2(n11789), .ZN(n11791) );
  NAND2_X1 U13329 ( .A1(n11792), .A2(n11791), .ZN(n13656) );
  NAND2_X1 U13330 ( .A1(n21671), .A2(n11631), .ZN(n11795) );
  NAND2_X1 U13331 ( .A1(n11795), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13637) );
  NAND2_X1 U13332 ( .A1(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n21910), .ZN(
        n11797) );
  NAND2_X1 U13333 ( .A1(n11772), .A2(P1_EAX_REG_0__SCAN_IN), .ZN(n11796) );
  OAI211_X1 U13334 ( .C1(n11825), .C2(n11448), .A(n11797), .B(n11796), .ZN(
        n11798) );
  AOI21_X1 U13335 ( .B1(n16743), .B2(n11991), .A(n11798), .ZN(n13636) );
  OR2_X1 U13336 ( .A1(n13637), .A2(n13636), .ZN(n13639) );
  INV_X1 U13337 ( .A(n13636), .ZN(n11800) );
  OR2_X1 U13338 ( .A1(n11800), .A2(n11799), .ZN(n11801) );
  NAND2_X1 U13339 ( .A1(n13639), .A2(n11801), .ZN(n13654) );
  NAND2_X1 U13340 ( .A1(n13656), .A2(n13654), .ZN(n13777) );
  INV_X1 U13341 ( .A(n11803), .ZN(n11804) );
  XNOR2_X1 U13342 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13954) );
  AOI21_X1 U13343 ( .B1(n12291), .B2(n13954), .A(n12294), .ZN(n11807) );
  NAND2_X1 U13344 ( .A1(n11772), .A2(P1_EAX_REG_2__SCAN_IN), .ZN(n11806) );
  OAI211_X1 U13345 ( .C1(n11825), .C2(n13622), .A(n11807), .B(n11806), .ZN(
        n11808) );
  INV_X1 U13346 ( .A(n11808), .ZN(n11809) );
  NAND2_X1 U13347 ( .A1(n12294), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11813) );
  NAND2_X1 U13348 ( .A1(n11810), .A2(n11813), .ZN(n13778) );
  INV_X1 U13349 ( .A(n13897), .ZN(n14107) );
  NAND2_X1 U13350 ( .A1(n11814), .A2(n14107), .ZN(n11815) );
  NAND2_X1 U13351 ( .A1(n11816), .A2(n11815), .ZN(n12407) );
  OR2_X1 U13352 ( .A1(n12407), .A2(n11958), .ZN(n11828) );
  INV_X1 U13353 ( .A(n11817), .ZN(n11821) );
  INV_X1 U13354 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n11819) );
  NAND2_X1 U13355 ( .A1(n11819), .A2(n11818), .ZN(n11820) );
  NAND2_X1 U13356 ( .A1(n11821), .A2(n11820), .ZN(n14092) );
  AOI22_X1 U13357 ( .A1(n14092), .A2(n12291), .B1(n12294), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n11824) );
  NAND2_X1 U13358 ( .A1(n12285), .A2(P1_EAX_REG_3__SCAN_IN), .ZN(n11823) );
  OAI211_X1 U13359 ( .C1(n11825), .C2(n11492), .A(n11824), .B(n11823), .ZN(
        n11826) );
  INV_X1 U13360 ( .A(n11826), .ZN(n11827) );
  NAND2_X1 U13361 ( .A1(n11828), .A2(n11827), .ZN(n13913) );
  INV_X1 U13362 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n11847) );
  AOI22_X1 U13363 ( .A1(n12127), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12269), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11833) );
  AOI22_X1 U13364 ( .A1(n11979), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12197), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11832) );
  AOI22_X1 U13365 ( .A1(n12271), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12218), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11831) );
  AOI22_X1 U13366 ( .A1(n10956), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11585), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11830) );
  NAND4_X1 U13367 ( .A1(n11833), .A2(n11832), .A3(n11831), .A4(n11830), .ZN(
        n11840) );
  AOI22_X1 U13368 ( .A1(n12223), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12247), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11838) );
  AOI22_X1 U13369 ( .A1(n10953), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12270), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11837) );
  AOI22_X1 U13370 ( .A1(n12264), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n12101), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11836) );
  AOI22_X1 U13371 ( .A1(n12263), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n11968), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11835) );
  NAND4_X1 U13372 ( .A1(n11838), .A2(n11837), .A3(n11836), .A4(n11835), .ZN(
        n11839) );
  NAND2_X1 U13373 ( .A1(n12343), .A2(n12443), .ZN(n11842) );
  NAND2_X1 U13374 ( .A1(n12302), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n11841) );
  NAND2_X1 U13375 ( .A1(n11848), .A2(n11849), .ZN(n12434) );
  NAND2_X1 U13376 ( .A1(n12434), .A2(n11991), .ZN(n11846) );
  NOR2_X1 U13377 ( .A1(n11843), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11844) );
  OR2_X1 U13378 ( .A1(n11855), .A2(n11844), .ZN(n21460) );
  AOI22_X1 U13379 ( .A1(n21460), .A2(n12291), .B1(n12294), .B2(
        P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n11845) );
  INV_X1 U13380 ( .A(n11848), .ZN(n11851) );
  NAND2_X1 U13381 ( .A1(n11851), .A2(n11850), .ZN(n12433) );
  INV_X1 U13382 ( .A(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11853) );
  NAND2_X1 U13383 ( .A1(n12343), .A2(n12453), .ZN(n11852) );
  OAI21_X1 U13384 ( .B1(n11853), .B2(n12333), .A(n11852), .ZN(n11854) );
  INV_X1 U13385 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n11859) );
  NOR2_X1 U13386 ( .A1(n11855), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11856) );
  OR2_X1 U13387 ( .A1(n11877), .A2(n11856), .ZN(n21477) );
  INV_X1 U13388 ( .A(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n21467) );
  NOR2_X1 U13389 ( .A1(n12023), .A2(n21467), .ZN(n11857) );
  AOI21_X1 U13390 ( .B1(n21477), .B2(n12291), .A(n11857), .ZN(n11858) );
  OAI21_X1 U13391 ( .B1(n11822), .B2(n11859), .A(n11858), .ZN(n11860) );
  AOI21_X1 U13392 ( .B1(n12441), .B2(n11991), .A(n11860), .ZN(n14461) );
  NOR2_X2 U13393 ( .A1(n14306), .A2(n14461), .ZN(n11861) );
  AOI22_X1 U13394 ( .A1(n12263), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n12218), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11865) );
  AOI22_X1 U13395 ( .A1(n12271), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12270), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11864) );
  AOI22_X1 U13396 ( .A1(n12127), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n11968), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11863) );
  NAND4_X1 U13397 ( .A1(n11865), .A2(n11864), .A3(n11863), .A4(n11862), .ZN(
        n11871) );
  AOI22_X1 U13398 ( .A1(n10951), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11979), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11869) );
  AOI22_X1 U13399 ( .A1(n10955), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12269), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11868) );
  AOI22_X1 U13400 ( .A1(n12247), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12197), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11867) );
  AOI22_X1 U13401 ( .A1(n12223), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12101), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11866) );
  NAND4_X1 U13402 ( .A1(n11869), .A2(n11868), .A3(n11867), .A4(n11866), .ZN(
        n11870) );
  OAI21_X1 U13403 ( .B1(n11871), .B2(n11870), .A(n11991), .ZN(n11875) );
  NAND2_X1 U13404 ( .A1(n12285), .A2(P1_EAX_REG_8__SCAN_IN), .ZN(n11874) );
  XNOR2_X1 U13405 ( .A(n11877), .B(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n14917) );
  NAND2_X1 U13406 ( .A1(n14917), .A2(n12291), .ZN(n11873) );
  NAND2_X1 U13407 ( .A1(n12294), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11872) );
  NAND4_X1 U13408 ( .A1(n11875), .A2(n11874), .A3(n11873), .A4(n11872), .ZN(
        n14497) );
  INV_X1 U13409 ( .A(n14497), .ZN(n11876) );
  XNOR2_X1 U13410 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .B(n11902), .ZN(
        n21478) );
  AOI22_X1 U13411 ( .A1(n12127), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n11878), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11882) );
  AOI22_X1 U13412 ( .A1(n11979), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n11545), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11881) );
  AOI22_X1 U13413 ( .A1(n12218), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n11585), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11880) );
  AOI22_X1 U13414 ( .A1(n12264), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n12270), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11879) );
  NAND4_X1 U13415 ( .A1(n11882), .A2(n11881), .A3(n11880), .A4(n11879), .ZN(
        n11888) );
  AOI22_X1 U13416 ( .A1(n12096), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12197), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11886) );
  AOI22_X1 U13417 ( .A1(n10955), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12263), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11885) );
  AOI22_X1 U13418 ( .A1(n10954), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n11968), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11884) );
  AOI22_X1 U13419 ( .A1(n12247), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12101), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11883) );
  NAND4_X1 U13420 ( .A1(n11886), .A2(n11885), .A3(n11884), .A4(n11883), .ZN(
        n11887) );
  OR2_X1 U13421 ( .A1(n11888), .A2(n11887), .ZN(n11889) );
  AOI22_X1 U13422 ( .A1(n11991), .A2(n11889), .B1(n12294), .B2(
        P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n11891) );
  NAND2_X1 U13423 ( .A1(n11772), .A2(P1_EAX_REG_9__SCAN_IN), .ZN(n11890) );
  OAI211_X1 U13424 ( .C1(n21478), .C2(n11799), .A(n11891), .B(n11890), .ZN(
        n14870) );
  AOI22_X1 U13425 ( .A1(n10954), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n10956), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11895) );
  AOI22_X1 U13426 ( .A1(n12127), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12269), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11894) );
  AOI22_X1 U13427 ( .A1(n12271), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12218), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11893) );
  AOI22_X1 U13428 ( .A1(n12264), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n12270), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11892) );
  NAND4_X1 U13429 ( .A1(n11895), .A2(n11894), .A3(n11893), .A4(n11892), .ZN(
        n11901) );
  AOI22_X1 U13430 ( .A1(n11979), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n12247), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11899) );
  AOI22_X1 U13431 ( .A1(n12263), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n11968), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11898) );
  AOI22_X1 U13432 ( .A1(n12223), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12101), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11897) );
  NAND4_X1 U13433 ( .A1(n11899), .A2(n11898), .A3(n11897), .A4(n11896), .ZN(
        n11900) );
  NOR2_X1 U13434 ( .A1(n11901), .A2(n11900), .ZN(n11905) );
  XNOR2_X1 U13435 ( .A(n11906), .B(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n19988) );
  NAND2_X1 U13436 ( .A1(n19988), .A2(n12291), .ZN(n11904) );
  AOI22_X1 U13437 ( .A1(n11772), .A2(P1_EAX_REG_10__SCAN_IN), .B1(n12294), 
        .B2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n11903) );
  OAI211_X1 U13438 ( .C1(n11905), .C2(n11958), .A(n11904), .B(n11903), .ZN(
        n14951) );
  INV_X1 U13439 ( .A(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n11909) );
  OAI21_X1 U13440 ( .B1(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n11907), .A(
        n11953), .ZN(n21503) );
  NAND2_X1 U13441 ( .A1(n21503), .A2(n12291), .ZN(n11908) );
  OAI21_X1 U13442 ( .B1(n11909), .B2(n12023), .A(n11908), .ZN(n11910) );
  AOI21_X1 U13443 ( .B1(n12285), .B2(P1_EAX_REG_11__SCAN_IN), .A(n11910), .ZN(
        n15076) );
  INV_X1 U13444 ( .A(n15076), .ZN(n11911) );
  AOI22_X1 U13445 ( .A1(n12127), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12269), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11915) );
  AOI22_X1 U13446 ( .A1(n12197), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n12264), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11914) );
  AOI22_X1 U13447 ( .A1(n12271), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12218), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11913) );
  AOI22_X1 U13448 ( .A1(n10956), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11585), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11912) );
  NAND4_X1 U13449 ( .A1(n11915), .A2(n11914), .A3(n11913), .A4(n11912), .ZN(
        n11921) );
  AOI22_X1 U13450 ( .A1(n11979), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12247), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11919) );
  AOI22_X1 U13451 ( .A1(n10953), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12270), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11918) );
  AOI22_X1 U13452 ( .A1(n12223), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12101), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11917) );
  AOI22_X1 U13453 ( .A1(n12263), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n11968), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11916) );
  NAND4_X1 U13454 ( .A1(n11919), .A2(n11918), .A3(n11917), .A4(n11916), .ZN(
        n11920) );
  OR2_X1 U13455 ( .A1(n11921), .A2(n11920), .ZN(n11922) );
  NAND2_X1 U13456 ( .A1(n11991), .A2(n11922), .ZN(n15083) );
  INV_X1 U13457 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n11925) );
  XNOR2_X1 U13458 ( .A(n11961), .B(n11925), .ZN(n21530) );
  OR2_X1 U13459 ( .A1(n21530), .A2(n11799), .ZN(n11942) );
  AOI22_X1 U13460 ( .A1(n12096), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12264), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11929) );
  AOI22_X1 U13461 ( .A1(n12223), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12197), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11928) );
  AOI22_X1 U13462 ( .A1(n12247), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12263), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11927) );
  AOI22_X1 U13463 ( .A1(n12271), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12101), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11926) );
  NAND4_X1 U13464 ( .A1(n11929), .A2(n11928), .A3(n11927), .A4(n11926), .ZN(
        n11936) );
  AOI22_X1 U13465 ( .A1(n10951), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11979), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11934) );
  AOI22_X1 U13466 ( .A1(n12218), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11968), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11933) );
  AOI22_X1 U13467 ( .A1(n12127), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12270), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11932) );
  NAND4_X1 U13468 ( .A1(n11934), .A2(n11933), .A3(n11932), .A4(n11931), .ZN(
        n11935) );
  NOR2_X1 U13469 ( .A1(n11936), .A2(n11935), .ZN(n11939) );
  NAND2_X1 U13470 ( .A1(n11772), .A2(P1_EAX_REG_13__SCAN_IN), .ZN(n11938) );
  NAND2_X1 U13471 ( .A1(n12294), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n11937) );
  OAI211_X1 U13472 ( .C1(n11958), .C2(n11939), .A(n11938), .B(n11937), .ZN(
        n11940) );
  INV_X1 U13473 ( .A(n11940), .ZN(n11941) );
  NAND2_X1 U13474 ( .A1(n11942), .A2(n11941), .ZN(n15087) );
  AOI22_X1 U13475 ( .A1(n10952), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n10956), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11946) );
  AOI22_X1 U13476 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n11979), .B1(
        n11545), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11945) );
  AOI22_X1 U13477 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n12197), .B1(
        n12263), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11944) );
  AOI22_X1 U13478 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n12223), .B1(
        n12218), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11943) );
  NAND4_X1 U13479 ( .A1(n11946), .A2(n11945), .A3(n11944), .A4(n11943), .ZN(
        n11952) );
  AOI22_X1 U13480 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n12127), .B1(
        n12247), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11950) );
  AOI22_X1 U13481 ( .A1(n12096), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12264), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11949) );
  AOI22_X1 U13482 ( .A1(n11585), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n11968), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11948) );
  AOI22_X1 U13483 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n12101), .B1(
        n12270), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11947) );
  NAND4_X1 U13484 ( .A1(n11950), .A2(n11949), .A3(n11948), .A4(n11947), .ZN(
        n11951) );
  NOR2_X1 U13485 ( .A1(n11952), .A2(n11951), .ZN(n11957) );
  XNOR2_X1 U13486 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B(n11953), .ZN(
        n21516) );
  OAI22_X1 U13487 ( .A1(n21516), .A2(n11799), .B1(n12023), .B2(n11924), .ZN(
        n11954) );
  INV_X1 U13488 ( .A(n11954), .ZN(n11956) );
  NAND2_X1 U13489 ( .A1(n11772), .A2(P1_EAX_REG_12__SCAN_IN), .ZN(n11955) );
  OAI211_X1 U13490 ( .C1(n11958), .C2(n11957), .A(n11956), .B(n11955), .ZN(
        n15095) );
  NAND2_X1 U13491 ( .A1(n15087), .A2(n15095), .ZN(n11959) );
  XOR2_X1 U13492 ( .A(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B(n11978), .Z(
        n21534) );
  AOI22_X1 U13493 ( .A1(n12127), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12223), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11967) );
  AOI22_X1 U13494 ( .A1(n10956), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12247), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11966) );
  AOI22_X1 U13495 ( .A1(n11962), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n12270), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11965) );
  AOI22_X1 U13496 ( .A1(n12271), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12101), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11964) );
  NAND4_X1 U13497 ( .A1(n11967), .A2(n11966), .A3(n11965), .A4(n11964), .ZN(
        n11974) );
  AOI22_X1 U13498 ( .A1(n10953), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12264), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11972) );
  AOI22_X1 U13499 ( .A1(n11979), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n12263), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11971) );
  AOI22_X1 U13500 ( .A1(n12096), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12218), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11969) );
  NAND4_X1 U13501 ( .A1(n11972), .A2(n11971), .A3(n11970), .A4(n11969), .ZN(
        n11973) );
  OR2_X1 U13502 ( .A1(n11974), .A2(n11973), .ZN(n11975) );
  AOI22_X1 U13503 ( .A1(n11991), .A2(n11975), .B1(n12294), .B2(
        P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n11977) );
  NAND2_X1 U13504 ( .A1(n11772), .A2(P1_EAX_REG_14__SCAN_IN), .ZN(n11976) );
  OAI211_X1 U13505 ( .C1(n21534), .C2(n11799), .A(n11977), .B(n11976), .ZN(
        n15704) );
  XNOR2_X1 U13506 ( .A(n11994), .B(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n21545) );
  AOI22_X1 U13507 ( .A1(n10952), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11537), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11983) );
  AOI22_X1 U13508 ( .A1(n12127), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12247), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11982) );
  AOI22_X1 U13509 ( .A1(n11979), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n12223), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11981) );
  AOI22_X1 U13510 ( .A1(n12271), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11963), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11980) );
  NAND4_X1 U13511 ( .A1(n11983), .A2(n11982), .A3(n11981), .A4(n11980), .ZN(
        n11989) );
  AOI22_X1 U13512 ( .A1(n10956), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12096), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11987) );
  AOI22_X1 U13513 ( .A1(n12263), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n12264), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11986) );
  AOI22_X1 U13514 ( .A1(n12218), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n11997), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11985) );
  AOI22_X1 U13515 ( .A1(n12270), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11585), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11984) );
  NAND4_X1 U13516 ( .A1(n11987), .A2(n11986), .A3(n11985), .A4(n11984), .ZN(
        n11988) );
  OR2_X1 U13517 ( .A1(n11989), .A2(n11988), .ZN(n11990) );
  AOI22_X1 U13518 ( .A1(n11991), .A2(n11990), .B1(n12294), .B2(
        P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n11993) );
  NAND2_X1 U13519 ( .A1(n11772), .A2(P1_EAX_REG_15__SCAN_IN), .ZN(n11992) );
  OAI211_X1 U13520 ( .C1(n21545), .C2(n11799), .A(n11993), .B(n11992), .ZN(
        n15698) );
  NAND2_X1 U13521 ( .A1(n15697), .A2(n15698), .ZN(n15620) );
  OR2_X1 U13522 ( .A1(n11995), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n11996) );
  NAND2_X1 U13523 ( .A1(n11996), .A2(n12027), .ZN(n21552) );
  AOI22_X1 U13524 ( .A1(n10955), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11537), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12001) );
  AOI22_X1 U13525 ( .A1(n10951), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11979), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12000) );
  AOI22_X1 U13526 ( .A1(n12127), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11968), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11999) );
  AOI22_X1 U13527 ( .A1(n12223), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12101), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11998) );
  NAND4_X1 U13528 ( .A1(n12001), .A2(n12000), .A3(n11999), .A4(n11998), .ZN(
        n12007) );
  AOI22_X1 U13529 ( .A1(n12247), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n12263), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12005) );
  AOI22_X1 U13530 ( .A1(n12096), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12218), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12004) );
  AOI22_X1 U13531 ( .A1(n12264), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12270), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12003) );
  NAND4_X1 U13532 ( .A1(n12005), .A2(n12004), .A3(n12003), .A4(n12002), .ZN(
        n12006) );
  NOR2_X1 U13533 ( .A1(n12007), .A2(n12006), .ZN(n12008) );
  NOR2_X1 U13534 ( .A1(n12287), .A2(n12008), .ZN(n12011) );
  INV_X1 U13535 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n15688) );
  NAND2_X1 U13536 ( .A1(n21910), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12009) );
  OAI211_X1 U13537 ( .C1(n11822), .C2(n15688), .A(n11799), .B(n12009), .ZN(
        n12010) );
  OAI22_X1 U13538 ( .A1(n21552), .A2(n11799), .B1(n12011), .B2(n12010), .ZN(
        n15619) );
  AOI22_X1 U13539 ( .A1(n10955), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12247), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12015) );
  AOI22_X1 U13540 ( .A1(n10952), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11537), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12014) );
  AOI22_X1 U13541 ( .A1(n12127), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n11997), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12013) );
  AOI22_X1 U13542 ( .A1(n12101), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n12270), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12012) );
  NAND4_X1 U13543 ( .A1(n12015), .A2(n12014), .A3(n12013), .A4(n12012), .ZN(
        n12021) );
  AOI22_X1 U13544 ( .A1(n11979), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n11545), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12019) );
  AOI22_X1 U13545 ( .A1(n12223), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12263), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12018) );
  AOI22_X1 U13546 ( .A1(n11641), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12218), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12016) );
  NAND4_X1 U13547 ( .A1(n12019), .A2(n12018), .A3(n12017), .A4(n12016), .ZN(
        n12020) );
  OAI21_X1 U13548 ( .B1(n12021), .B2(n12020), .A(n12256), .ZN(n12026) );
  XNOR2_X1 U13549 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B(n12027), .ZN(
        n15788) );
  INV_X1 U13550 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n12022) );
  OAI22_X1 U13551 ( .A1(n15788), .A2(n11799), .B1(n12023), .B2(n12022), .ZN(
        n12024) );
  AOI21_X1 U13552 ( .B1(n12285), .B2(P1_EAX_REG_17__SCAN_IN), .A(n12024), .ZN(
        n12025) );
  OR2_X1 U13553 ( .A1(n12028), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n12029) );
  NAND2_X1 U13554 ( .A1(n12029), .A2(n12059), .ZN(n21565) );
  AOI22_X1 U13555 ( .A1(n12127), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11979), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12033) );
  AOI22_X1 U13556 ( .A1(n12096), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12247), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12032) );
  AOI22_X1 U13557 ( .A1(n12197), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n11545), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12031) );
  AOI22_X1 U13558 ( .A1(n10954), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12218), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12030) );
  NAND4_X1 U13559 ( .A1(n12033), .A2(n12032), .A3(n12031), .A4(n12030), .ZN(
        n12039) );
  AOI22_X1 U13560 ( .A1(n12223), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12263), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12037) );
  AOI22_X1 U13561 ( .A1(n12264), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12101), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12036) );
  AOI22_X1 U13562 ( .A1(n10956), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12270), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12035) );
  AOI22_X1 U13563 ( .A1(n11585), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n11997), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12034) );
  NAND4_X1 U13564 ( .A1(n12037), .A2(n12036), .A3(n12035), .A4(n12034), .ZN(
        n12038) );
  NOR2_X1 U13565 ( .A1(n12039), .A2(n12038), .ZN(n12040) );
  NOR2_X1 U13566 ( .A1(n12287), .A2(n12040), .ZN(n12043) );
  INV_X1 U13567 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n15675) );
  NAND2_X1 U13568 ( .A1(n21910), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n12041) );
  OAI211_X1 U13569 ( .C1(n11822), .C2(n15675), .A(n11799), .B(n12041), .ZN(
        n12042) );
  OAI22_X1 U13570 ( .A1(n21565), .A2(n11799), .B1(n12043), .B2(n12042), .ZN(
        n15609) );
  AOI22_X1 U13571 ( .A1(n10952), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11979), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12047) );
  AOI22_X1 U13572 ( .A1(n11537), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n12264), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12046) );
  AOI22_X1 U13573 ( .A1(n10955), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12270), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12045) );
  AOI22_X1 U13574 ( .A1(n11878), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11963), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12044) );
  NAND4_X1 U13575 ( .A1(n12047), .A2(n12046), .A3(n12045), .A4(n12044), .ZN(
        n12053) );
  AOI22_X1 U13576 ( .A1(n12271), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12263), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12051) );
  AOI22_X1 U13577 ( .A1(n12127), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11997), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12050) );
  AOI22_X1 U13578 ( .A1(n12096), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12218), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12049) );
  NAND4_X1 U13579 ( .A1(n12051), .A2(n12050), .A3(n12049), .A4(n12048), .ZN(
        n12052) );
  NOR2_X1 U13580 ( .A1(n12053), .A2(n12052), .ZN(n12056) );
  AOI21_X1 U13581 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n21573), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n12054) );
  AOI21_X1 U13582 ( .B1(n12285), .B2(P1_EAX_REG_19__SCAN_IN), .A(n12054), .ZN(
        n12055) );
  OAI21_X1 U13583 ( .B1(n12287), .B2(n12056), .A(n12055), .ZN(n12058) );
  XNOR2_X1 U13584 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B(n12059), .ZN(
        n21578) );
  NAND2_X1 U13585 ( .A1(n21578), .A2(n12291), .ZN(n12057) );
  OR2_X1 U13586 ( .A1(n12060), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12061) );
  NAND2_X1 U13587 ( .A1(n12061), .A2(n12093), .ZN(n21590) );
  INV_X1 U13588 ( .A(n21590), .ZN(n12076) );
  AOI22_X1 U13589 ( .A1(n11979), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n11537), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12065) );
  AOI22_X1 U13590 ( .A1(n12096), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12264), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12064) );
  AOI22_X1 U13591 ( .A1(n12127), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n11968), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12063) );
  AOI22_X1 U13592 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n12270), .B1(
        n12218), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12062) );
  NAND4_X1 U13593 ( .A1(n12065), .A2(n12064), .A3(n12063), .A4(n12062), .ZN(
        n12071) );
  AOI22_X1 U13594 ( .A1(n10952), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n10955), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12069) );
  AOI22_X1 U13595 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n12247), .B1(
        n12263), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12068) );
  AOI22_X1 U13596 ( .A1(n12223), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n11585), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12067) );
  AOI22_X1 U13597 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n12271), .B1(
        n12101), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12066) );
  NAND4_X1 U13598 ( .A1(n12069), .A2(n12068), .A3(n12067), .A4(n12066), .ZN(
        n12070) );
  OR2_X1 U13599 ( .A1(n12071), .A2(n12070), .ZN(n12074) );
  INV_X1 U13600 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n15667) );
  NAND2_X1 U13601 ( .A1(n21910), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12072) );
  OAI211_X1 U13602 ( .C1(n11822), .C2(n15667), .A(n11799), .B(n12072), .ZN(
        n12073) );
  AOI21_X1 U13603 ( .B1(n12256), .B2(n12074), .A(n12073), .ZN(n12075) );
  AOI21_X1 U13604 ( .B1(n12076), .B2(n12291), .A(n12075), .ZN(n15595) );
  AOI22_X1 U13605 ( .A1(n10955), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11979), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12080) );
  AOI22_X1 U13606 ( .A1(n12096), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12263), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12079) );
  AOI22_X1 U13607 ( .A1(n12247), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12264), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12078) );
  AOI22_X1 U13608 ( .A1(n12223), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11963), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12077) );
  NAND4_X1 U13609 ( .A1(n12080), .A2(n12079), .A3(n12078), .A4(n12077), .ZN(
        n12086) );
  AOI22_X1 U13610 ( .A1(n10953), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12218), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12084) );
  AOI22_X1 U13611 ( .A1(n12271), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12270), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12083) );
  AOI22_X1 U13612 ( .A1(n12127), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11968), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12082) );
  AOI22_X1 U13613 ( .A1(n11537), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11585), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12081) );
  NAND4_X1 U13614 ( .A1(n12084), .A2(n12083), .A3(n12082), .A4(n12081), .ZN(
        n12085) );
  NOR2_X1 U13615 ( .A1(n12086), .A2(n12085), .ZN(n12090) );
  NAND2_X1 U13616 ( .A1(n21910), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12087) );
  NAND2_X1 U13617 ( .A1(n11799), .A2(n12087), .ZN(n12088) );
  AOI21_X1 U13618 ( .B1(n12285), .B2(P1_EAX_REG_21__SCAN_IN), .A(n12088), .ZN(
        n12089) );
  OAI21_X1 U13619 ( .B1(n12287), .B2(n12090), .A(n12089), .ZN(n12092) );
  XNOR2_X1 U13620 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B(n12093), .ZN(
        n21597) );
  NAND2_X1 U13621 ( .A1(n21597), .A2(n12291), .ZN(n12091) );
  NAND2_X1 U13622 ( .A1(n12092), .A2(n12091), .ZN(n15590) );
  INV_X1 U13623 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n21593) );
  OR2_X1 U13624 ( .A1(n12094), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n12095) );
  NAND2_X1 U13625 ( .A1(n12095), .A2(n12139), .ZN(n21605) );
  AOI22_X1 U13626 ( .A1(n10956), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12247), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12100) );
  AOI22_X1 U13627 ( .A1(n12096), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12197), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12099) );
  AOI22_X1 U13628 ( .A1(n12218), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11968), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12098) );
  AOI22_X1 U13629 ( .A1(n12271), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12270), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12097) );
  NAND4_X1 U13630 ( .A1(n12100), .A2(n12099), .A3(n12098), .A4(n12097), .ZN(
        n12107) );
  AOI22_X1 U13631 ( .A1(n10954), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12127), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12105) );
  AOI22_X1 U13632 ( .A1(n12263), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n12264), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12104) );
  AOI22_X1 U13633 ( .A1(n11979), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n11585), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12103) );
  AOI22_X1 U13634 ( .A1(n12223), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12101), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12102) );
  NAND4_X1 U13635 ( .A1(n12105), .A2(n12104), .A3(n12103), .A4(n12102), .ZN(
        n12106) );
  NOR2_X1 U13636 ( .A1(n12107), .A2(n12106), .ZN(n12108) );
  NOR2_X1 U13637 ( .A1(n12287), .A2(n12108), .ZN(n12111) );
  INV_X1 U13638 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n15659) );
  NAND2_X1 U13639 ( .A1(n21910), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n12109) );
  OAI211_X1 U13640 ( .C1(n11822), .C2(n15659), .A(n11799), .B(n12109), .ZN(
        n12110) );
  OAI22_X1 U13641 ( .A1(n21605), .A2(n11799), .B1(n12111), .B2(n12110), .ZN(
        n15582) );
  INV_X1 U13642 ( .A(n15582), .ZN(n12112) );
  AOI22_X1 U13643 ( .A1(n12223), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11962), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12116) );
  AOI22_X1 U13644 ( .A1(n11979), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n12271), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12115) );
  AOI22_X1 U13645 ( .A1(n12269), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12270), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12113) );
  NAND4_X1 U13646 ( .A1(n12116), .A2(n12115), .A3(n12114), .A4(n12113), .ZN(
        n12122) );
  AOI22_X1 U13647 ( .A1(n10954), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12127), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12120) );
  AOI22_X1 U13648 ( .A1(n12247), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12263), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12119) );
  AOI22_X1 U13649 ( .A1(n10955), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12218), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12118) );
  AOI22_X1 U13650 ( .A1(n12264), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12101), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12117) );
  NAND4_X1 U13651 ( .A1(n12120), .A2(n12119), .A3(n12118), .A4(n12117), .ZN(
        n12121) );
  NOR2_X1 U13652 ( .A1(n12122), .A2(n12121), .ZN(n12143) );
  AOI22_X1 U13653 ( .A1(n12223), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12264), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12126) );
  AOI22_X1 U13654 ( .A1(n11979), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n12101), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12125) );
  AOI22_X1 U13655 ( .A1(n12096), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12270), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12124) );
  AOI22_X1 U13656 ( .A1(n12218), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n11968), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12123) );
  NAND4_X1 U13657 ( .A1(n12126), .A2(n12125), .A3(n12124), .A4(n12123), .ZN(
        n12133) );
  AOI22_X1 U13658 ( .A1(n12127), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n10955), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12131) );
  AOI22_X1 U13659 ( .A1(n12197), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n12271), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12130) );
  AOI22_X1 U13660 ( .A1(n12247), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12263), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12129) );
  AOI22_X1 U13661 ( .A1(n10952), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11585), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12128) );
  NAND4_X1 U13662 ( .A1(n12131), .A2(n12130), .A3(n12129), .A4(n12128), .ZN(
        n12132) );
  NOR2_X1 U13663 ( .A1(n12133), .A2(n12132), .ZN(n12142) );
  XOR2_X1 U13664 ( .A(n12143), .B(n12142), .Z(n12134) );
  NAND2_X1 U13665 ( .A1(n12134), .A2(n12256), .ZN(n12138) );
  INV_X1 U13666 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n15757) );
  AOI21_X1 U13667 ( .B1(n15757), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n12135) );
  AOI21_X1 U13668 ( .B1(n12285), .B2(P1_EAX_REG_23__SCAN_IN), .A(n12135), .ZN(
        n12137) );
  XNOR2_X1 U13669 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .B(n12139), .ZN(
        n15761) );
  AOI21_X1 U13670 ( .B1(n12138), .B2(n12137), .A(n12136), .ZN(n15552) );
  OR2_X1 U13671 ( .A1(n12140), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n12141) );
  NAND2_X1 U13672 ( .A1(n12141), .A2(n12177), .ZN(n21619) );
  NOR2_X1 U13673 ( .A1(n12143), .A2(n12142), .ZN(n12170) );
  AOI22_X1 U13674 ( .A1(n10954), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12127), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12147) );
  AOI22_X1 U13675 ( .A1(n12096), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12263), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12146) );
  AOI22_X1 U13676 ( .A1(n12218), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n11968), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12145) );
  AOI22_X1 U13677 ( .A1(n10955), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11585), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12144) );
  NAND4_X1 U13678 ( .A1(n12147), .A2(n12146), .A3(n12145), .A4(n12144), .ZN(
        n12153) );
  AOI22_X1 U13679 ( .A1(n11979), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n12223), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12151) );
  AOI22_X1 U13680 ( .A1(n12197), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n12264), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12150) );
  AOI22_X1 U13681 ( .A1(n12247), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12270), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12149) );
  AOI22_X1 U13682 ( .A1(n12271), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n12101), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12148) );
  NAND4_X1 U13683 ( .A1(n12151), .A2(n12150), .A3(n12149), .A4(n12148), .ZN(
        n12152) );
  OR2_X1 U13684 ( .A1(n12153), .A2(n12152), .ZN(n12169) );
  XNOR2_X1 U13685 ( .A(n12170), .B(n12169), .ZN(n12157) );
  INV_X1 U13686 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n12154) );
  AOI21_X1 U13687 ( .B1(n12154), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n12155) );
  AOI21_X1 U13688 ( .B1(n12285), .B2(P1_EAX_REG_24__SCAN_IN), .A(n12155), .ZN(
        n12156) );
  OAI21_X1 U13689 ( .B1(n12157), .B2(n12287), .A(n12156), .ZN(n12158) );
  OAI21_X1 U13690 ( .B1(n21619), .B2(n11799), .A(n12158), .ZN(n15576) );
  AOI22_X1 U13691 ( .A1(n12096), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12218), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12162) );
  AOI22_X1 U13692 ( .A1(n11979), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n12101), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12161) );
  AOI22_X1 U13693 ( .A1(n12264), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12270), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12160) );
  NAND4_X1 U13694 ( .A1(n12162), .A2(n12161), .A3(n12160), .A4(n12159), .ZN(
        n12168) );
  AOI22_X1 U13695 ( .A1(n12127), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n10955), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12166) );
  AOI22_X1 U13696 ( .A1(n12247), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12197), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12165) );
  AOI22_X1 U13697 ( .A1(n12223), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12271), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12164) );
  AOI22_X1 U13698 ( .A1(n10953), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12263), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12163) );
  NAND4_X1 U13699 ( .A1(n12166), .A2(n12165), .A3(n12164), .A4(n12163), .ZN(
        n12167) );
  NOR2_X1 U13700 ( .A1(n12168), .A2(n12167), .ZN(n12181) );
  NAND2_X1 U13701 ( .A1(n12170), .A2(n12169), .ZN(n12180) );
  XOR2_X1 U13702 ( .A(n12181), .B(n12180), .Z(n12173) );
  INV_X1 U13703 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n15646) );
  NAND2_X1 U13704 ( .A1(n21910), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n12171) );
  OAI211_X1 U13705 ( .C1(n11822), .C2(n15646), .A(n11799), .B(n12171), .ZN(
        n12172) );
  AOI21_X1 U13706 ( .B1(n12173), .B2(n12256), .A(n12172), .ZN(n12174) );
  INV_X1 U13707 ( .A(n12174), .ZN(n12176) );
  XNOR2_X1 U13708 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .B(n12177), .ZN(
        n21628) );
  NAND2_X1 U13709 ( .A1(n21628), .A2(n12291), .ZN(n12175) );
  INV_X1 U13710 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n21637) );
  OR2_X1 U13711 ( .A1(n12178), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12179) );
  NAND2_X1 U13712 ( .A1(n12179), .A2(n12234), .ZN(n21643) );
  NOR2_X1 U13713 ( .A1(n12181), .A2(n12180), .ZN(n12209) );
  AOI22_X1 U13714 ( .A1(n10951), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12127), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12185) );
  AOI22_X1 U13715 ( .A1(n12096), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12263), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12184) );
  AOI22_X1 U13716 ( .A1(n12218), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n11997), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12183) );
  NAND4_X1 U13717 ( .A1(n12185), .A2(n12184), .A3(n12183), .A4(n12182), .ZN(
        n12191) );
  AOI22_X1 U13718 ( .A1(n11979), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n12223), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12189) );
  AOI22_X1 U13719 ( .A1(n12197), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12264), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12188) );
  AOI22_X1 U13720 ( .A1(n12247), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12270), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12187) );
  AOI22_X1 U13721 ( .A1(n12271), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12101), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12186) );
  NAND4_X1 U13722 ( .A1(n12189), .A2(n12188), .A3(n12187), .A4(n12186), .ZN(
        n12190) );
  OR2_X1 U13723 ( .A1(n12191), .A2(n12190), .ZN(n12208) );
  XNOR2_X1 U13724 ( .A(n12209), .B(n12208), .ZN(n12195) );
  NAND2_X1 U13725 ( .A1(n21910), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12192) );
  NAND2_X1 U13726 ( .A1(n11799), .A2(n12192), .ZN(n12193) );
  AOI21_X1 U13727 ( .B1(n12285), .B2(P1_EAX_REG_26__SCAN_IN), .A(n12193), .ZN(
        n12194) );
  OAI21_X1 U13728 ( .B1(n12195), .B2(n12287), .A(n12194), .ZN(n12196) );
  OAI21_X1 U13729 ( .B1(n21643), .B2(n11799), .A(n12196), .ZN(n15640) );
  AOI22_X1 U13730 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n12247), .B1(
        n12197), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12201) );
  AOI22_X1 U13731 ( .A1(n11878), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12264), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12200) );
  AOI22_X1 U13732 ( .A1(n11585), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n11997), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12199) );
  AOI22_X1 U13733 ( .A1(n12263), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n12218), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12198) );
  NAND4_X1 U13734 ( .A1(n12201), .A2(n12200), .A3(n12199), .A4(n12198), .ZN(
        n12207) );
  AOI22_X1 U13735 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n12127), .B1(
        n10956), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12205) );
  AOI22_X1 U13736 ( .A1(n10953), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12269), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12204) );
  AOI22_X1 U13737 ( .A1(n11979), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n12270), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12203) );
  AOI22_X1 U13738 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n12271), .B1(
        n12101), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12202) );
  NAND4_X1 U13739 ( .A1(n12205), .A2(n12204), .A3(n12203), .A4(n12202), .ZN(
        n12206) );
  NOR2_X1 U13740 ( .A1(n12207), .A2(n12206), .ZN(n12217) );
  NAND2_X1 U13741 ( .A1(n12209), .A2(n12208), .ZN(n12216) );
  XOR2_X1 U13742 ( .A(n12217), .B(n12216), .Z(n12210) );
  NAND2_X1 U13743 ( .A1(n12210), .A2(n12256), .ZN(n12215) );
  NAND2_X1 U13744 ( .A1(n21910), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n12211) );
  NAND2_X1 U13745 ( .A1(n11799), .A2(n12211), .ZN(n12212) );
  AOI21_X1 U13746 ( .B1(n12285), .B2(P1_EAX_REG_27__SCAN_IN), .A(n12212), .ZN(
        n12214) );
  XNOR2_X1 U13747 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .B(n12234), .ZN(
        n15739) );
  AOI21_X1 U13748 ( .B1(n12215), .B2(n12214), .A(n12213), .ZN(n15540) );
  NOR2_X1 U13749 ( .A1(n12217), .A2(n12216), .ZN(n12255) );
  AOI22_X1 U13750 ( .A1(n10951), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12127), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12222) );
  AOI22_X1 U13751 ( .A1(n11641), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12263), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12221) );
  AOI22_X1 U13752 ( .A1(n12218), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11997), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12220) );
  NAND4_X1 U13753 ( .A1(n12222), .A2(n12221), .A3(n12220), .A4(n12219), .ZN(
        n12229) );
  AOI22_X1 U13754 ( .A1(n11979), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n12223), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12227) );
  AOI22_X1 U13755 ( .A1(n11537), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12264), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12226) );
  AOI22_X1 U13756 ( .A1(n12247), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12270), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12225) );
  AOI22_X1 U13757 ( .A1(n12271), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12101), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12224) );
  NAND4_X1 U13758 ( .A1(n12227), .A2(n12226), .A3(n12225), .A4(n12224), .ZN(
        n12228) );
  OR2_X1 U13759 ( .A1(n12229), .A2(n12228), .ZN(n12254) );
  INV_X1 U13760 ( .A(n12254), .ZN(n12230) );
  XNOR2_X1 U13761 ( .A(n12255), .B(n12230), .ZN(n12231) );
  NAND2_X1 U13762 ( .A1(n12231), .A2(n12256), .ZN(n12242) );
  NAND2_X1 U13763 ( .A1(n21910), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12232) );
  NAND2_X1 U13764 ( .A1(n11799), .A2(n12232), .ZN(n12233) );
  AOI21_X1 U13765 ( .B1(n12285), .B2(P1_EAX_REG_28__SCAN_IN), .A(n12233), .ZN(
        n12241) );
  INV_X1 U13766 ( .A(n12234), .ZN(n12235) );
  INV_X1 U13767 ( .A(n12236), .ZN(n12238) );
  INV_X1 U13768 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n12237) );
  NAND2_X1 U13769 ( .A1(n12238), .A2(n12237), .ZN(n12239) );
  NAND2_X1 U13770 ( .A1(n12289), .A2(n12239), .ZN(n15729) );
  NOR2_X1 U13771 ( .A1(n15729), .A2(n11799), .ZN(n12240) );
  AOI21_X1 U13772 ( .B1(n12242), .B2(n12241), .A(n12240), .ZN(n15527) );
  AOI22_X1 U13773 ( .A1(n10953), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n10956), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12246) );
  AOI22_X1 U13774 ( .A1(n11878), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12264), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12245) );
  AOI22_X1 U13775 ( .A1(n12218), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n11997), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12244) );
  NAND4_X1 U13776 ( .A1(n12246), .A2(n12245), .A3(n12244), .A4(n12243), .ZN(
        n12253) );
  AOI22_X1 U13777 ( .A1(n12127), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12269), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12251) );
  AOI22_X1 U13778 ( .A1(n11979), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n11537), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12250) );
  AOI22_X1 U13779 ( .A1(n12247), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12270), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12249) );
  AOI22_X1 U13780 ( .A1(n12271), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n12101), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12248) );
  NAND4_X1 U13781 ( .A1(n12251), .A2(n12250), .A3(n12249), .A4(n12248), .ZN(
        n12252) );
  NOR2_X1 U13782 ( .A1(n12253), .A2(n12252), .ZN(n12280) );
  NAND2_X1 U13783 ( .A1(n12255), .A2(n12254), .ZN(n12279) );
  XOR2_X1 U13784 ( .A(n12280), .B(n12279), .Z(n12257) );
  NAND2_X1 U13785 ( .A1(n12257), .A2(n12256), .ZN(n12262) );
  NAND2_X1 U13786 ( .A1(n21910), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12258) );
  NAND2_X1 U13787 ( .A1(n11799), .A2(n12258), .ZN(n12259) );
  AOI21_X1 U13788 ( .B1(n12285), .B2(P1_EAX_REG_29__SCAN_IN), .A(n12259), .ZN(
        n12261) );
  XNOR2_X1 U13789 ( .A(n12289), .B(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15496) );
  AND2_X1 U13790 ( .A1(n15496), .A2(n12291), .ZN(n12260) );
  AOI22_X1 U13791 ( .A1(n10955), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12263), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12268) );
  AOI22_X1 U13792 ( .A1(n12247), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11537), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12267) );
  AOI22_X1 U13793 ( .A1(n11979), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n12264), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12266) );
  AOI22_X1 U13794 ( .A1(n12218), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n11997), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12265) );
  NAND4_X1 U13795 ( .A1(n12268), .A2(n12267), .A3(n12266), .A4(n12265), .ZN(
        n12278) );
  AOI22_X1 U13796 ( .A1(n10954), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12269), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12276) );
  AOI22_X1 U13797 ( .A1(n11878), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12270), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12275) );
  AOI22_X1 U13798 ( .A1(n12271), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n12101), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12274) );
  AOI22_X1 U13799 ( .A1(n12127), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11585), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12273) );
  NAND4_X1 U13800 ( .A1(n12276), .A2(n12275), .A3(n12274), .A4(n12273), .ZN(
        n12277) );
  NOR2_X1 U13801 ( .A1(n12278), .A2(n12277), .ZN(n12282) );
  NOR2_X1 U13802 ( .A1(n12280), .A2(n12279), .ZN(n12281) );
  XOR2_X1 U13803 ( .A(n12282), .B(n12281), .Z(n12288) );
  NAND2_X1 U13804 ( .A1(n21910), .A2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12283) );
  NAND2_X1 U13805 ( .A1(n11799), .A2(n12283), .ZN(n12284) );
  AOI21_X1 U13806 ( .B1(n12285), .B2(P1_EAX_REG_30__SCAN_IN), .A(n12284), .ZN(
        n12286) );
  OAI21_X1 U13807 ( .B1(n12288), .B2(n12287), .A(n12286), .ZN(n12293) );
  INV_X1 U13808 ( .A(n12289), .ZN(n12290) );
  NAND2_X1 U13809 ( .A1(n12290), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12493) );
  XNOR2_X1 U13810 ( .A(n12493), .B(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15717) );
  NAND2_X1 U13811 ( .A1(n15717), .A2(n12291), .ZN(n12292) );
  NAND2_X1 U13812 ( .A1(n12293), .A2(n12292), .ZN(n15513) );
  AOI22_X1 U13813 ( .A1(n11772), .A2(P1_EAX_REG_31__SCAN_IN), .B1(n12294), 
        .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n12295) );
  MUX2_X1 U13814 ( .A(n11700), .B(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .S(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n12317) );
  NOR2_X1 U13815 ( .A1(n21864), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12297) );
  NAND2_X1 U13816 ( .A1(n21864), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12296) );
  NAND2_X1 U13817 ( .A1(n12317), .A2(n12318), .ZN(n12299) );
  NAND2_X1 U13818 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n11700), .ZN(
        n12298) );
  INV_X1 U13819 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n12300) );
  MUX2_X1 U13820 ( .A(n12300), .B(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .S(
        n11492), .Z(n12301) );
  XNOR2_X1 U13821 ( .A(n12330), .B(n12301), .ZN(n12327) );
  XNOR2_X1 U13822 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n12307), .ZN(
        n12303) );
  XNOR2_X1 U13823 ( .A(n12303), .B(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n12350) );
  INV_X1 U13824 ( .A(n12350), .ZN(n12304) );
  AOI211_X1 U13825 ( .C1(n12343), .C2(n13732), .A(n12304), .B(n12305), .ZN(
        n12316) );
  AOI21_X1 U13826 ( .B1(n12320), .B2(n12440), .A(n12350), .ZN(n12315) );
  INV_X1 U13827 ( .A(n12305), .ZN(n12306) );
  NAND2_X1 U13828 ( .A1(n12306), .A2(n14298), .ZN(n12313) );
  OAI21_X1 U13829 ( .B1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n21877), .A(
        n12307), .ZN(n12309) );
  OAI21_X1 U13830 ( .B1(n12320), .B2(n12309), .A(n12341), .ZN(n12312) );
  INV_X1 U13831 ( .A(n12309), .ZN(n12310) );
  OAI211_X1 U13832 ( .C1(n13905), .C2(n13570), .A(n12322), .B(n12310), .ZN(
        n12311) );
  OAI211_X1 U13833 ( .C1(n12350), .C2(n12313), .A(n12312), .B(n12311), .ZN(
        n12314) );
  OAI21_X1 U13834 ( .B1(n12316), .B2(n12315), .A(n12314), .ZN(n12326) );
  XOR2_X1 U13835 ( .A(n12318), .B(n12317), .Z(n12351) );
  INV_X1 U13836 ( .A(n12351), .ZN(n12319) );
  INV_X1 U13837 ( .A(n12324), .ZN(n12321) );
  OAI211_X1 U13838 ( .C1(n12333), .C2(n12351), .A(n12322), .B(n12321), .ZN(
        n12325) );
  INV_X1 U13839 ( .A(n12322), .ZN(n12323) );
  INV_X1 U13840 ( .A(n12327), .ZN(n12332) );
  NOR2_X1 U13841 ( .A1(n11492), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n12328) );
  NOR2_X1 U13842 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n16773), .ZN(
        n12331) );
  NAND2_X1 U13843 ( .A1(n12333), .A2(n12349), .ZN(n12336) );
  INV_X1 U13844 ( .A(n12341), .ZN(n12335) );
  NAND2_X1 U13845 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n16773), .ZN(
        n12337) );
  NAND2_X1 U13846 ( .A1(n12338), .A2(n12337), .ZN(n12340) );
  NAND2_X1 U13847 ( .A1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n11775), .ZN(
        n12339) );
  AND2_X4 U13848 ( .A1(n12345), .A2(n12344), .ZN(n13735) );
  INV_X1 U13849 ( .A(n13725), .ZN(n13597) );
  AND2_X4 U13850 ( .A1(n13732), .A2(n13747), .ZN(n13663) );
  NAND2_X1 U13851 ( .A1(n13597), .A2(n13663), .ZN(n13741) );
  NAND2_X1 U13852 ( .A1(READY1), .A2(READY11_REG_SCAN_IN), .ZN(n21675) );
  AND2_X1 U13853 ( .A1(n13460), .A2(n11615), .ZN(n12346) );
  NAND2_X1 U13854 ( .A1(n16006), .A2(n12346), .ZN(n13466) );
  OAI21_X1 U13855 ( .B1(n13741), .B2(n21712), .A(n13466), .ZN(n12347) );
  NAND2_X1 U13856 ( .A1(n13735), .A2(n12347), .ZN(n12356) );
  INV_X1 U13857 ( .A(n12348), .ZN(n16702) );
  INV_X1 U13858 ( .A(n12349), .ZN(n12354) );
  AND2_X1 U13859 ( .A1(n12351), .A2(n12350), .ZN(n12353) );
  NAND3_X1 U13860 ( .A1(n16702), .A2(n13729), .A3(n21675), .ZN(n12355) );
  NAND2_X1 U13861 ( .A1(n12356), .A2(n12355), .ZN(n13606) );
  AND4_X1 U13862 ( .A1(n15506), .A2(n14173), .A3(n20029), .A4(n12357), .ZN(
        n13658) );
  NAND2_X1 U13863 ( .A1(n13584), .A2(n13658), .ZN(n12358) );
  AND2_X1 U13864 ( .A1(n15703), .A2(n15506), .ZN(n12360) );
  NOR4_X1 U13865 ( .A1(P1_ADDRESS_REG_15__SCAN_IN), .A2(
        P1_ADDRESS_REG_13__SCAN_IN), .A3(P1_ADDRESS_REG_12__SCAN_IN), .A4(
        P1_ADDRESS_REG_11__SCAN_IN), .ZN(n12364) );
  NOR4_X1 U13866 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(
        P1_ADDRESS_REG_17__SCAN_IN), .A3(P1_ADDRESS_REG_14__SCAN_IN), .A4(
        P1_ADDRESS_REG_16__SCAN_IN), .ZN(n12363) );
  NOR4_X1 U13867 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(
        P1_ADDRESS_REG_5__SCAN_IN), .A3(P1_ADDRESS_REG_4__SCAN_IN), .A4(
        P1_ADDRESS_REG_3__SCAN_IN), .ZN(n12362) );
  NOR4_X1 U13868 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(
        P1_ADDRESS_REG_7__SCAN_IN), .A3(P1_ADDRESS_REG_9__SCAN_IN), .A4(
        P1_ADDRESS_REG_8__SCAN_IN), .ZN(n12361) );
  AND4_X1 U13869 ( .A1(n12364), .A2(n12363), .A3(n12362), .A4(n12361), .ZN(
        n12369) );
  NOR4_X1 U13870 ( .A1(P1_ADDRESS_REG_2__SCAN_IN), .A2(
        P1_ADDRESS_REG_1__SCAN_IN), .A3(P1_ADDRESS_REG_26__SCAN_IN), .A4(
        P1_ADDRESS_REG_28__SCAN_IN), .ZN(n12367) );
  NOR4_X1 U13871 ( .A1(P1_ADDRESS_REG_22__SCAN_IN), .A2(
        P1_ADDRESS_REG_21__SCAN_IN), .A3(P1_ADDRESS_REG_20__SCAN_IN), .A4(
        P1_ADDRESS_REG_19__SCAN_IN), .ZN(n12366) );
  NOR4_X1 U13872 ( .A1(P1_ADDRESS_REG_27__SCAN_IN), .A2(
        P1_ADDRESS_REG_25__SCAN_IN), .A3(P1_ADDRESS_REG_24__SCAN_IN), .A4(
        P1_ADDRESS_REG_23__SCAN_IN), .ZN(n12365) );
  INV_X1 U13873 ( .A(P1_ADDRESS_REG_0__SCAN_IN), .ZN(n19886) );
  AND4_X1 U13874 ( .A1(n12367), .A2(n12366), .A3(n12365), .A4(n19886), .ZN(
        n12368) );
  NAND2_X1 U13875 ( .A1(n12369), .A2(n12368), .ZN(n12370) );
  NOR3_X1 U13876 ( .A1(n15707), .A2(n11614), .A3(n14376), .ZN(n12371) );
  AOI22_X1 U13877 ( .A1(n15694), .A2(BUF1_REG_31__SCAN_IN), .B1(
        P1_EAX_REG_31__SCAN_IN), .B2(n15707), .ZN(n12372) );
  INV_X1 U13878 ( .A(n12372), .ZN(n12375) );
  NOR2_X1 U13879 ( .A1(n11614), .A2(n14301), .ZN(n12373) );
  NAND2_X1 U13880 ( .A1(n15703), .A2(n12373), .ZN(n15689) );
  INV_X1 U13881 ( .A(DATAI_31_), .ZN(n13935) );
  NOR2_X1 U13882 ( .A1(n15689), .A2(n13935), .ZN(n12374) );
  NOR2_X1 U13883 ( .A1(n12375), .A2(n12374), .ZN(n12376) );
  NAND2_X1 U13884 ( .A1(n12377), .A2(n12376), .ZN(P1_U2873) );
  NAND3_X1 U13885 ( .A1(n21321), .A2(P1_STATEBS16_REG_SCAN_IN), .A3(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n21676) );
  INV_X1 U13886 ( .A(n21676), .ZN(n12382) );
  NAND2_X1 U13887 ( .A1(n12396), .A2(n12395), .ZN(n12409) );
  INV_X1 U13888 ( .A(n12383), .ZN(n12408) );
  XNOR2_X1 U13889 ( .A(n12409), .B(n12408), .ZN(n12385) );
  AND2_X1 U13890 ( .A1(n13905), .A2(n12384), .ZN(n12389) );
  AOI21_X1 U13891 ( .B1(n12385), .B2(n21319), .A(n12389), .ZN(n12386) );
  NAND2_X1 U13892 ( .A1(n12387), .A2(n12386), .ZN(n13761) );
  INV_X1 U13893 ( .A(n12389), .ZN(n12390) );
  OAI21_X1 U13894 ( .B1(n14295), .B2(n12395), .A(n12390), .ZN(n12391) );
  INV_X1 U13895 ( .A(n12391), .ZN(n12392) );
  OR2_X1 U13896 ( .A1(n12394), .A2(n11443), .ZN(n12400) );
  XNOR2_X1 U13897 ( .A(n12396), .B(n12395), .ZN(n12397) );
  INV_X1 U13898 ( .A(n12398), .ZN(n12399) );
  NAND2_X1 U13899 ( .A1(n12400), .A2(n12399), .ZN(n12401) );
  INV_X1 U13900 ( .A(n12401), .ZN(n12402) );
  OR2_X1 U13901 ( .A1(n19971), .A2(n12402), .ZN(n12403) );
  NAND2_X1 U13902 ( .A1(n13762), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12405) );
  INV_X1 U13903 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n12406) );
  OR2_X1 U13904 ( .A1(n12407), .A2(n11443), .ZN(n12413) );
  NAND2_X1 U13905 ( .A1(n12409), .A2(n12408), .ZN(n12410) );
  NAND2_X1 U13906 ( .A1(n12410), .A2(n12411), .ZN(n12426) );
  OAI211_X1 U13907 ( .C1(n12411), .C2(n12410), .A(n12426), .B(n21319), .ZN(
        n12412) );
  NAND2_X1 U13908 ( .A1(n12413), .A2(n12412), .ZN(n13872) );
  NAND2_X1 U13909 ( .A1(n12414), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12415) );
  NAND2_X1 U13910 ( .A1(n12416), .A2(n12440), .ZN(n12419) );
  XNOR2_X1 U13911 ( .A(n12426), .B(n12424), .ZN(n12417) );
  NAND2_X1 U13912 ( .A1(n12417), .A2(n21319), .ZN(n12418) );
  NAND2_X1 U13913 ( .A1(n12419), .A2(n12418), .ZN(n12420) );
  INV_X1 U13914 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n12543) );
  XNOR2_X1 U13915 ( .A(n12420), .B(n12543), .ZN(n14097) );
  NAND2_X1 U13916 ( .A1(n14098), .A2(n14097), .ZN(n12422) );
  NAND2_X1 U13917 ( .A1(n12420), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12421) );
  NAND2_X1 U13918 ( .A1(n12423), .A2(n12440), .ZN(n12430) );
  INV_X1 U13919 ( .A(n12424), .ZN(n12425) );
  NOR2_X1 U13920 ( .A1(n12426), .A2(n12425), .ZN(n12428) );
  NAND2_X1 U13921 ( .A1(n12428), .A2(n12427), .ZN(n12442) );
  OAI211_X1 U13922 ( .C1(n12428), .C2(n12427), .A(n12442), .B(n21319), .ZN(
        n12429) );
  NAND2_X1 U13923 ( .A1(n12430), .A2(n12429), .ZN(n12431) );
  OR2_X1 U13924 ( .A1(n12431), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12432) );
  NAND3_X1 U13925 ( .A1(n12433), .A2(n12440), .A3(n12434), .ZN(n12437) );
  XNOR2_X1 U13926 ( .A(n12442), .B(n12443), .ZN(n12435) );
  NAND2_X1 U13927 ( .A1(n12435), .A2(n21319), .ZN(n12436) );
  NAND2_X1 U13928 ( .A1(n12437), .A2(n12436), .ZN(n12438) );
  INV_X1 U13929 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n14476) );
  XNOR2_X1 U13930 ( .A(n12438), .B(n14476), .ZN(n14468) );
  NAND2_X1 U13931 ( .A1(n12438), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12439) );
  NAND2_X1 U13932 ( .A1(n12441), .A2(n12440), .ZN(n12447) );
  INV_X1 U13933 ( .A(n12442), .ZN(n12444) );
  NAND2_X1 U13934 ( .A1(n12444), .A2(n12443), .ZN(n12455) );
  XNOR2_X1 U13935 ( .A(n12455), .B(n12453), .ZN(n12445) );
  NAND2_X1 U13936 ( .A1(n12445), .A2(n21319), .ZN(n12446) );
  NAND2_X1 U13937 ( .A1(n12447), .A2(n12446), .ZN(n12448) );
  INV_X1 U13938 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n14883) );
  XNOR2_X1 U13939 ( .A(n12448), .B(n14883), .ZN(n14877) );
  AND2_X1 U13940 ( .A1(n12448), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12449) );
  AOI21_X2 U13941 ( .B1(n14876), .B2(n14877), .A(n12449), .ZN(n14906) );
  INV_X1 U13942 ( .A(n12450), .ZN(n12451) );
  NOR2_X1 U13943 ( .A1(n12451), .A2(n11443), .ZN(n12452) );
  NAND2_X1 U13944 ( .A1(n21319), .A2(n12453), .ZN(n12454) );
  OR2_X1 U13945 ( .A1(n12455), .A2(n12454), .ZN(n12456) );
  NAND2_X1 U13946 ( .A1(n12469), .A2(n12456), .ZN(n12457) );
  INV_X1 U13947 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n12560) );
  XNOR2_X1 U13948 ( .A(n12457), .B(n12560), .ZN(n14907) );
  NOR2_X1 U13949 ( .A1(n12457), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12458) );
  XNOR2_X1 U13950 ( .A(n15881), .B(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n14922) );
  INV_X1 U13951 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n14934) );
  XNOR2_X1 U13952 ( .A(n12469), .B(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n15800) );
  INV_X1 U13953 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n15988) );
  NAND2_X1 U13954 ( .A1(n15881), .A2(n15988), .ZN(n15798) );
  INV_X1 U13955 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n12581) );
  NAND2_X1 U13956 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15794) );
  OAI21_X1 U13957 ( .B1(n12581), .B2(n15794), .A(n15881), .ZN(n12460) );
  NAND2_X1 U13958 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15899) );
  INV_X1 U13959 ( .A(n15899), .ZN(n15781) );
  NAND2_X1 U13960 ( .A1(n15781), .A2(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n12461) );
  NOR2_X1 U13961 ( .A1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n12465) );
  NOR2_X1 U13962 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n12462) );
  OR2_X1 U13963 ( .A1(n15881), .A2(n12462), .ZN(n15795) );
  OR2_X1 U13964 ( .A1(n15881), .A2(n15988), .ZN(n15797) );
  NOR2_X1 U13965 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n12463) );
  OR2_X1 U13966 ( .A1(n15881), .A2(n12463), .ZN(n15929) );
  INV_X1 U13967 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15932) );
  OR2_X1 U13968 ( .A1(n15881), .A2(n15932), .ZN(n12464) );
  OAI211_X1 U13969 ( .C1(n12465), .C2(n15881), .A(n15930), .B(n15782), .ZN(
        n12466) );
  INV_X1 U13970 ( .A(n12466), .ZN(n12467) );
  INV_X1 U13971 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n12468) );
  NAND2_X1 U13972 ( .A1(n12470), .A2(n15994), .ZN(n15763) );
  INV_X1 U13973 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15901) );
  INV_X1 U13974 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15917) );
  INV_X1 U13975 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n15900) );
  AND3_X1 U13976 ( .A1(n15901), .A2(n15917), .A3(n15900), .ZN(n12471) );
  OR2_X1 U13977 ( .A1(n15881), .A2(n12471), .ZN(n12472) );
  AND2_X2 U13978 ( .A1(n15763), .A2(n12472), .ZN(n15897) );
  AND4_X1 U13979 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A4(
        P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n15909) );
  INV_X1 U13980 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15885) );
  INV_X1 U13981 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15889) );
  INV_X1 U13982 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n21398) );
  NAND2_X1 U13983 ( .A1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15872) );
  INV_X1 U13984 ( .A(n15872), .ZN(n12474) );
  NAND2_X1 U13985 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n12474), .ZN(
        n15826) );
  NAND2_X1 U13986 ( .A1(n15881), .A2(n15826), .ZN(n15723) );
  INV_X1 U13987 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15741) );
  NOR2_X1 U13988 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15858) );
  AND2_X1 U13989 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15860) );
  INV_X1 U13990 ( .A(n15860), .ZN(n15836) );
  NAND2_X1 U13991 ( .A1(n15881), .A2(n15836), .ZN(n12477) );
  INV_X1 U13992 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15850) );
  AND2_X1 U13993 ( .A1(n15881), .A2(n15850), .ZN(n12480) );
  INV_X1 U13994 ( .A(n12480), .ZN(n12478) );
  OR2_X1 U13995 ( .A1(n15881), .A2(n15850), .ZN(n12503) );
  OAI21_X1 U13996 ( .B1(n15714), .B2(n12480), .A(n12479), .ZN(n12481) );
  OAI21_X1 U13997 ( .B1(n12508), .B2(n15714), .A(n12481), .ZN(n15857) );
  INV_X1 U13998 ( .A(n15857), .ZN(n12485) );
  OR2_X1 U13999 ( .A1(n13634), .A2(n11640), .ZN(n12483) );
  AND2_X1 U14000 ( .A1(n12483), .A2(n12482), .ZN(n13577) );
  NAND2_X1 U14001 ( .A1(n16740), .A2(n13905), .ZN(n12484) );
  NAND3_X1 U14002 ( .A1(n13577), .A2(n11615), .A3(n12484), .ZN(n13598) );
  NOR2_X1 U14003 ( .A1(n13598), .A2(n13570), .ZN(n13468) );
  NAND2_X1 U14004 ( .A1(n21915), .A2(n12489), .ZN(n21323) );
  NAND2_X1 U14005 ( .A1(n21323), .A2(n21321), .ZN(n12486) );
  NAND2_X1 U14006 ( .A1(n14152), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n12488) );
  NOR2_X1 U14007 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n21910), .ZN(n16765) );
  INV_X1 U14008 ( .A(n16765), .ZN(n12487) );
  NAND2_X1 U14009 ( .A1(n12488), .A2(n12487), .ZN(n19974) );
  INV_X1 U14010 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n15499) );
  NAND2_X1 U14011 ( .A1(n10970), .A2(P1_REIP_REG_29__SCAN_IN), .ZN(n15852) );
  OAI21_X1 U14012 ( .B1(n19987), .B2(n15499), .A(n15852), .ZN(n12490) );
  AOI21_X1 U14013 ( .B1(n15496), .B2(n20005), .A(n12490), .ZN(n12491) );
  INV_X2 U14014 ( .A(n20018), .ZN(n20009) );
  INV_X1 U14015 ( .A(n12493), .ZN(n12494) );
  NAND2_X1 U14016 ( .A1(n12494), .A2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12496) );
  INV_X1 U14017 ( .A(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n12495) );
  INV_X2 U14018 ( .A(n19987), .ZN(n20022) );
  INV_X1 U14019 ( .A(P1_REIP_REG_31__SCAN_IN), .ZN(n19929) );
  NOR2_X1 U14020 ( .A1(n21386), .A2(n19929), .ZN(n15829) );
  AOI21_X1 U14021 ( .B1(n20022), .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n15829), .ZN(n12497) );
  OAI21_X1 U14022 ( .B1(n20028), .B2(n13952), .A(n12497), .ZN(n12498) );
  AOI21_X1 U14023 ( .B1(n12519), .B2(n20009), .A(n12498), .ZN(n12509) );
  INV_X1 U14024 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n15821) );
  XNOR2_X1 U14025 ( .A(n12469), .B(n15821), .ZN(n12500) );
  INV_X1 U14026 ( .A(n12500), .ZN(n12499) );
  INV_X1 U14027 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15838) );
  NAND2_X1 U14028 ( .A1(n15881), .A2(n15838), .ZN(n12502) );
  NAND2_X1 U14029 ( .A1(n12499), .A2(n12502), .ZN(n12507) );
  NOR2_X1 U14030 ( .A1(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n12501) );
  OAI211_X1 U14031 ( .C1(n12501), .C2(n15881), .A(n12508), .B(n12500), .ZN(
        n12506) );
  OAI211_X1 U14032 ( .C1(n15881), .C2(n15838), .A(n12503), .B(n12502), .ZN(
        n12504) );
  NAND2_X1 U14033 ( .A1(n12504), .A2(n15821), .ZN(n12505) );
  NAND2_X1 U14034 ( .A1(n13735), .A2(n12510), .ZN(n12514) );
  INV_X1 U14035 ( .A(n13729), .ZN(n12512) );
  NOR2_X1 U14036 ( .A1(n12511), .A2(n12512), .ZN(n13463) );
  INV_X1 U14037 ( .A(n13463), .ZN(n12513) );
  AOI21_X2 U14038 ( .B1(n12514), .B2(n12513), .A(n21689), .ZN(n21324) );
  NOR2_X1 U14039 ( .A1(P1_STATEBS16_REG_SCAN_IN), .A2(n16772), .ZN(n12515) );
  NAND2_X1 U14040 ( .A1(n16772), .A2(n21910), .ZN(n21320) );
  OAI21_X1 U14041 ( .B1(n21868), .B2(n21320), .A(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n16737) );
  OAI21_X1 U14042 ( .B1(P1_STATE2_REG_0__SCAN_IN), .B2(n12515), .A(n16737), 
        .ZN(n12516) );
  NOR2_X1 U14043 ( .A1(n12516), .A2(n16765), .ZN(n12517) );
  NOR2_X1 U14044 ( .A1(n13952), .A2(n16772), .ZN(n12518) );
  AND4_X1 U14045 ( .A1(P1_REIP_REG_9__SCAN_IN), .A2(P1_REIP_REG_8__SCAN_IN), 
        .A3(P1_REIP_REG_7__SCAN_IN), .A4(P1_REIP_REG_10__SCAN_IN), .ZN(n21490)
         );
  NAND4_X1 U14046 ( .A1(P1_REIP_REG_2__SCAN_IN), .A2(P1_REIP_REG_1__SCAN_IN), 
        .A3(P1_REIP_REG_3__SCAN_IN), .A4(P1_REIP_REG_4__SCAN_IN), .ZN(n21458)
         );
  INV_X1 U14047 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n20034) );
  AND2_X1 U14048 ( .A1(n12520), .A2(n20034), .ZN(n21718) );
  OAI21_X1 U14049 ( .B1(n13732), .B2(n21718), .A(n21675), .ZN(n13724) );
  INV_X1 U14050 ( .A(n12637), .ZN(n12522) );
  AND2_X2 U14051 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n12521), .ZN(n12633) );
  INV_X1 U14052 ( .A(P1_REIP_REG_6__SCAN_IN), .ZN(n21463) );
  INV_X1 U14053 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n21509) );
  NAND2_X1 U14054 ( .A1(n21515), .A2(P1_REIP_REG_12__SCAN_IN), .ZN(n21532) );
  INV_X1 U14055 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n21522) );
  INV_X1 U14056 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n19904) );
  INV_X1 U14057 ( .A(P1_REIP_REG_17__SCAN_IN), .ZN(n21366) );
  NOR2_X2 U14058 ( .A1(n11009), .A2(n21366), .ZN(n21563) );
  INV_X1 U14059 ( .A(P1_REIP_REG_19__SCAN_IN), .ZN(n21582) );
  INV_X1 U14060 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n21601) );
  INV_X1 U14061 ( .A(P1_REIP_REG_23__SCAN_IN), .ZN(n19913) );
  INV_X1 U14062 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n19919) );
  NOR2_X2 U14063 ( .A1(n21616), .A2(n19919), .ZN(n21638) );
  INV_X1 U14064 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n19925) );
  INV_X1 U14065 ( .A(P1_REIP_REG_30__SCAN_IN), .ZN(n19931) );
  OR2_X1 U14066 ( .A1(n13680), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12526) );
  INV_X1 U14067 ( .A(P1_EBX_REG_30__SCAN_IN), .ZN(n12524) );
  NAND2_X1 U14068 ( .A1(n13663), .A2(n12524), .ZN(n12525) );
  NAND2_X1 U14069 ( .A1(n12526), .A2(n12525), .ZN(n15518) );
  AND2_X2 U14070 ( .A1(n15514), .A2(n13663), .ZN(n12617) );
  INV_X1 U14071 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n21425) );
  NAND2_X1 U14072 ( .A1(n12617), .A2(n21425), .ZN(n12531) );
  INV_X1 U14073 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n12527) );
  NAND2_X1 U14074 ( .A1(n12592), .A2(n12527), .ZN(n12529) );
  NAND2_X1 U14075 ( .A1(n13663), .A2(n21425), .ZN(n12528) );
  NAND3_X1 U14076 ( .A1(n12529), .A2(n12613), .A3(n12528), .ZN(n12530) );
  NAND2_X1 U14077 ( .A1(n12531), .A2(n12530), .ZN(n12535) );
  NAND2_X1 U14078 ( .A1(n12592), .A2(P1_EBX_REG_0__SCAN_IN), .ZN(n12534) );
  INV_X1 U14079 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n14081) );
  NAND2_X1 U14080 ( .A1(n12613), .A2(n14081), .ZN(n12533) );
  NAND2_X1 U14081 ( .A1(n12534), .A2(n12533), .ZN(n13679) );
  XNOR2_X1 U14082 ( .A(n12535), .B(n13679), .ZN(n21424) );
  INV_X1 U14083 ( .A(n12535), .ZN(n12536) );
  AOI21_X1 U14084 ( .B1(n21424), .B2(n13663), .A(n12536), .ZN(n13768) );
  INV_X1 U14085 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n13760) );
  NAND2_X1 U14086 ( .A1(n12592), .A2(n13760), .ZN(n12538) );
  INV_X1 U14087 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n13947) );
  NAND2_X1 U14088 ( .A1(n13663), .A2(n13947), .ZN(n12537) );
  NAND3_X1 U14089 ( .A1(n12538), .A2(n12613), .A3(n12537), .ZN(n12539) );
  OAI21_X1 U14090 ( .B1(n12627), .B2(P1_EBX_REG_2__SCAN_IN), .A(n12539), .ZN(
        n13767) );
  MUX2_X1 U14091 ( .A(n12614), .B(n12613), .S(P1_EBX_REG_3__SCAN_IN), .Z(
        n12540) );
  INV_X1 U14092 ( .A(n12540), .ZN(n12542) );
  NOR2_X1 U14093 ( .A1(n13680), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12541) );
  NOR2_X1 U14094 ( .A1(n12542), .A2(n12541), .ZN(n13874) );
  NAND2_X1 U14095 ( .A1(n13875), .A2(n13874), .ZN(n14100) );
  INV_X1 U14096 ( .A(P1_EBX_REG_4__SCAN_IN), .ZN(n21434) );
  NAND2_X1 U14097 ( .A1(n12617), .A2(n21434), .ZN(n12547) );
  NAND2_X1 U14098 ( .A1(n12592), .A2(n12543), .ZN(n12545) );
  NAND2_X1 U14099 ( .A1(n13663), .A2(n21434), .ZN(n12544) );
  NAND3_X1 U14100 ( .A1(n12545), .A2(n12613), .A3(n12544), .ZN(n12546) );
  AND2_X1 U14101 ( .A1(n12547), .A2(n12546), .ZN(n14099) );
  INV_X1 U14102 ( .A(P1_EBX_REG_5__SCAN_IN), .ZN(n12550) );
  NAND2_X1 U14103 ( .A1(n13663), .A2(n12550), .ZN(n12552) );
  NAND2_X1 U14104 ( .A1(n12613), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12551) );
  NAND3_X1 U14105 ( .A1(n12552), .A2(n12592), .A3(n12551), .ZN(n12553) );
  OAI21_X1 U14106 ( .B1(n12614), .B2(P1_EBX_REG_5__SCAN_IN), .A(n12553), .ZN(
        n14257) );
  NAND2_X1 U14107 ( .A1(n12592), .A2(n14476), .ZN(n12555) );
  INV_X1 U14108 ( .A(P1_EBX_REG_6__SCAN_IN), .ZN(n21455) );
  NAND2_X1 U14109 ( .A1(n13663), .A2(n21455), .ZN(n12554) );
  NAND3_X1 U14110 ( .A1(n12555), .A2(n12613), .A3(n12554), .ZN(n12556) );
  OAI21_X1 U14111 ( .B1(n12627), .B2(P1_EBX_REG_6__SCAN_IN), .A(n12556), .ZN(
        n14309) );
  INV_X1 U14112 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n21469) );
  NAND2_X1 U14113 ( .A1(n13663), .A2(n21469), .ZN(n12558) );
  NAND2_X1 U14114 ( .A1(n12613), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12557) );
  NAND3_X1 U14115 ( .A1(n12558), .A2(n12592), .A3(n12557), .ZN(n12559) );
  OAI21_X1 U14116 ( .B1(n12614), .B2(P1_EBX_REG_7__SCAN_IN), .A(n12559), .ZN(
        n14463) );
  INV_X1 U14117 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n14505) );
  NAND2_X1 U14118 ( .A1(n12617), .A2(n14505), .ZN(n12564) );
  NAND2_X1 U14119 ( .A1(n12592), .A2(n12560), .ZN(n12562) );
  NAND2_X1 U14120 ( .A1(n13663), .A2(n14505), .ZN(n12561) );
  NAND3_X1 U14121 ( .A1(n12562), .A2(n12613), .A3(n12561), .ZN(n12563) );
  MUX2_X1 U14122 ( .A(n12614), .B(n12613), .S(P1_EBX_REG_9__SCAN_IN), .Z(
        n12565) );
  NAND2_X1 U14123 ( .A1(n11482), .A2(n12565), .ZN(n14873) );
  INV_X1 U14124 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15997) );
  NAND2_X1 U14125 ( .A1(n12592), .A2(n15997), .ZN(n12567) );
  INV_X1 U14126 ( .A(P1_EBX_REG_10__SCAN_IN), .ZN(n14955) );
  NAND2_X1 U14127 ( .A1(n13663), .A2(n14955), .ZN(n12566) );
  NAND3_X1 U14128 ( .A1(n12567), .A2(n12613), .A3(n12566), .ZN(n12568) );
  OAI21_X1 U14129 ( .B1(n12627), .B2(P1_EBX_REG_10__SCAN_IN), .A(n12568), .ZN(
        n14952) );
  MUX2_X1 U14130 ( .A(n12614), .B(n12613), .S(P1_EBX_REG_11__SCAN_IN), .Z(
        n12569) );
  INV_X1 U14131 ( .A(n12569), .ZN(n12571) );
  NOR2_X1 U14132 ( .A1(n13680), .A2(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n12570) );
  NOR2_X1 U14133 ( .A1(n12571), .A2(n12570), .ZN(n15080) );
  INV_X1 U14134 ( .A(P1_EBX_REG_12__SCAN_IN), .ZN(n15105) );
  NAND2_X1 U14135 ( .A1(n12613), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n12572) );
  NAND2_X1 U14136 ( .A1(n12592), .A2(n12572), .ZN(n12574) );
  NAND2_X1 U14137 ( .A1(n13663), .A2(n15105), .ZN(n12573) );
  AOI22_X1 U14138 ( .A1(n12617), .A2(n15105), .B1(n12574), .B2(n12573), .ZN(
        n15101) );
  MUX2_X1 U14139 ( .A(n12614), .B(n12613), .S(P1_EBX_REG_13__SCAN_IN), .Z(
        n12575) );
  OAI21_X1 U14140 ( .B1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n13680), .A(
        n12575), .ZN(n15091) );
  OR2_X2 U14141 ( .A1(n15104), .A2(n15091), .ZN(n15974) );
  INV_X1 U14142 ( .A(n12614), .ZN(n12576) );
  INV_X1 U14143 ( .A(P1_EBX_REG_15__SCAN_IN), .ZN(n21542) );
  NAND2_X1 U14144 ( .A1(n12576), .A2(n21542), .ZN(n12580) );
  NAND2_X1 U14145 ( .A1(n13663), .A2(n21542), .ZN(n12578) );
  NAND2_X1 U14146 ( .A1(n12613), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n12577) );
  NAND3_X1 U14147 ( .A1(n12578), .A2(n12592), .A3(n12577), .ZN(n12579) );
  AND2_X1 U14148 ( .A1(n12580), .A2(n12579), .ZN(n15952) );
  INV_X1 U14149 ( .A(P1_EBX_REG_14__SCAN_IN), .ZN(n19964) );
  NAND2_X1 U14150 ( .A1(n12617), .A2(n19964), .ZN(n12585) );
  NAND2_X1 U14151 ( .A1(n12592), .A2(n12581), .ZN(n12583) );
  NAND2_X1 U14152 ( .A1(n13663), .A2(n19964), .ZN(n12582) );
  NAND3_X1 U14153 ( .A1(n12583), .A2(n12613), .A3(n12582), .ZN(n12584) );
  NAND2_X1 U14154 ( .A1(n12585), .A2(n12584), .ZN(n15973) );
  NAND2_X1 U14155 ( .A1(n15952), .A2(n15973), .ZN(n12586) );
  NOR2_X2 U14156 ( .A1(n15974), .A2(n12586), .ZN(n15949) );
  INV_X1 U14157 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n12587) );
  NAND2_X1 U14158 ( .A1(n12592), .A2(n12587), .ZN(n12589) );
  INV_X1 U14159 ( .A(P1_EBX_REG_16__SCAN_IN), .ZN(n15625) );
  NAND2_X1 U14160 ( .A1(n13663), .A2(n15625), .ZN(n12588) );
  NAND3_X1 U14161 ( .A1(n12589), .A2(n12532), .A3(n12588), .ZN(n12590) );
  OAI21_X1 U14162 ( .B1(n12627), .B2(P1_EBX_REG_16__SCAN_IN), .A(n12590), .ZN(
        n15622) );
  NAND2_X1 U14163 ( .A1(n15949), .A2(n15622), .ZN(n15624) );
  MUX2_X1 U14164 ( .A(n12614), .B(n12532), .S(P1_EBX_REG_17__SCAN_IN), .Z(
        n12591) );
  OAI21_X1 U14165 ( .B1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n13680), .A(
        n12591), .ZN(n15563) );
  OR2_X2 U14166 ( .A1(n15624), .A2(n15563), .ZN(n15612) );
  INV_X1 U14167 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n21560) );
  NAND2_X1 U14168 ( .A1(n12617), .A2(n21560), .ZN(n12596) );
  NAND2_X1 U14169 ( .A1(n12592), .A2(n12468), .ZN(n12594) );
  NAND2_X1 U14170 ( .A1(n13663), .A2(n21560), .ZN(n12593) );
  NAND3_X1 U14171 ( .A1(n12594), .A2(n12613), .A3(n12593), .ZN(n12595) );
  MUX2_X1 U14172 ( .A(n12614), .B(n12532), .S(P1_EBX_REG_19__SCAN_IN), .Z(
        n12597) );
  INV_X1 U14173 ( .A(n12597), .ZN(n12599) );
  NOR2_X1 U14174 ( .A1(n13680), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n12598) );
  NOR2_X1 U14175 ( .A1(n12599), .A2(n12598), .ZN(n15605) );
  NAND2_X1 U14176 ( .A1(n12592), .A2(n15917), .ZN(n12601) );
  INV_X1 U14177 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n15599) );
  NAND2_X1 U14178 ( .A1(n13663), .A2(n15599), .ZN(n12600) );
  NAND3_X1 U14179 ( .A1(n12601), .A2(n12532), .A3(n12600), .ZN(n12602) );
  OAI21_X1 U14180 ( .B1(n12627), .B2(P1_EBX_REG_20__SCAN_IN), .A(n12602), .ZN(
        n15597) );
  MUX2_X1 U14181 ( .A(n12614), .B(n12532), .S(P1_EBX_REG_21__SCAN_IN), .Z(
        n12603) );
  NAND2_X1 U14182 ( .A1(n11480), .A2(n12603), .ZN(n15593) );
  INV_X1 U14183 ( .A(P1_EBX_REG_22__SCAN_IN), .ZN(n15587) );
  NAND2_X1 U14184 ( .A1(n12617), .A2(n15587), .ZN(n12607) );
  INV_X1 U14185 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15908) );
  NAND2_X1 U14186 ( .A1(n12592), .A2(n15908), .ZN(n12605) );
  NAND2_X1 U14187 ( .A1(n13663), .A2(n15587), .ZN(n12604) );
  NAND3_X1 U14188 ( .A1(n12605), .A2(n12532), .A3(n12604), .ZN(n12606) );
  AND2_X1 U14189 ( .A1(n12607), .A2(n12606), .ZN(n15584) );
  MUX2_X1 U14190 ( .A(n12614), .B(n12532), .S(P1_EBX_REG_23__SCAN_IN), .Z(
        n12608) );
  OAI21_X1 U14191 ( .B1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n13680), .A(
        n12608), .ZN(n15553) );
  NOR2_X2 U14192 ( .A1(n15586), .A2(n15553), .ZN(n15579) );
  NAND2_X1 U14193 ( .A1(n12592), .A2(n15885), .ZN(n12610) );
  INV_X1 U14194 ( .A(P1_EBX_REG_24__SCAN_IN), .ZN(n21618) );
  NAND2_X1 U14195 ( .A1(n13663), .A2(n21618), .ZN(n12609) );
  NAND3_X1 U14196 ( .A1(n12610), .A2(n12613), .A3(n12609), .ZN(n12611) );
  OAI21_X1 U14197 ( .B1(n12627), .B2(P1_EBX_REG_24__SCAN_IN), .A(n12611), .ZN(
        n15578) );
  MUX2_X1 U14198 ( .A(n12614), .B(n12532), .S(P1_EBX_REG_25__SCAN_IN), .Z(
        n12612) );
  NAND2_X1 U14199 ( .A1(n11481), .A2(n12612), .ZN(n15574) );
  MUX2_X1 U14200 ( .A(n12614), .B(n12613), .S(P1_EBX_REG_27__SCAN_IN), .Z(
        n12615) );
  OAI21_X1 U14201 ( .B1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n13680), .A(
        n12615), .ZN(n12616) );
  INV_X1 U14202 ( .A(n12616), .ZN(n15543) );
  INV_X1 U14203 ( .A(P1_EBX_REG_26__SCAN_IN), .ZN(n21641) );
  NAND2_X1 U14204 ( .A1(n12617), .A2(n21641), .ZN(n12621) );
  NAND2_X1 U14205 ( .A1(n12592), .A2(n15741), .ZN(n12619) );
  NAND2_X1 U14206 ( .A1(n13663), .A2(n21641), .ZN(n12618) );
  NAND3_X1 U14207 ( .A1(n12619), .A2(n12613), .A3(n12618), .ZN(n12620) );
  NAND2_X1 U14208 ( .A1(n12621), .A2(n12620), .ZN(n15869) );
  INV_X1 U14209 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n12622) );
  NAND2_X1 U14210 ( .A1(n12592), .A2(n12622), .ZN(n12625) );
  INV_X1 U14211 ( .A(P1_EBX_REG_28__SCAN_IN), .ZN(n12623) );
  NAND2_X1 U14212 ( .A1(n13663), .A2(n12623), .ZN(n12624) );
  NAND3_X1 U14213 ( .A1(n12625), .A2(n12532), .A3(n12624), .ZN(n12626) );
  OAI21_X1 U14214 ( .B1(n12627), .B2(P1_EBX_REG_28__SCAN_IN), .A(n12626), .ZN(
        n15529) );
  OR2_X1 U14215 ( .A1(n13680), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12628) );
  INV_X1 U14216 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n15510) );
  NAND2_X1 U14217 ( .A1(n13663), .A2(n15510), .ZN(n12629) );
  NAND2_X1 U14218 ( .A1(n12628), .A2(n12629), .ZN(n15515) );
  MUX2_X1 U14219 ( .A(n15515), .B(n12629), .S(n15514), .Z(n15494) );
  MUX2_X1 U14220 ( .A(n15518), .B(n12532), .S(n11011), .Z(n12632) );
  INV_X1 U14221 ( .A(n13663), .ZN(n12630) );
  OAI22_X1 U14222 ( .A1(n13680), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        n12630), .B2(P1_EBX_REG_31__SCAN_IN), .ZN(n12631) );
  XNOR2_X2 U14223 ( .A(n12632), .B(n12631), .ZN(n15806) );
  AND2_X1 U14224 ( .A1(n13732), .A2(P1_EBX_REG_31__SCAN_IN), .ZN(n12636) );
  INV_X1 U14225 ( .A(n12633), .ZN(n13944) );
  AOI21_X1 U14226 ( .B1(n21675), .B2(n14152), .A(n13944), .ZN(n12634) );
  AND2_X1 U14227 ( .A1(n13747), .A2(n12634), .ZN(n12635) );
  NAND2_X1 U14228 ( .A1(n21645), .A2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n12640) );
  NOR2_X1 U14229 ( .A1(n11049), .A2(n12636), .ZN(n12638) );
  NAND2_X1 U14230 ( .A1(n21626), .A2(P1_EBX_REG_31__SCAN_IN), .ZN(n12639) );
  NAND2_X1 U14231 ( .A1(n12642), .A2(n21639), .ZN(n15525) );
  INV_X1 U14232 ( .A(n13142), .ZN(n12665) );
  AOI22_X1 U14233 ( .A1(n12665), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n10957), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12644) );
  AND2_X1 U14234 ( .A1(n12644), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12652) );
  AOI22_X1 U14235 ( .A1(n12866), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12738), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12651) );
  AND2_X4 U14236 ( .A1(n12873), .A2(n14027), .ZN(n13107) );
  AOI22_X1 U14237 ( .A1(n16064), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n13107), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12650) );
  AND3_X4 U14238 ( .A1(n12647), .A2(n12646), .A3(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n16063) );
  AND3_X4 U14239 ( .A1(n12648), .A2(n12646), .A3(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n16068) );
  AOI22_X1 U14240 ( .A1(n16063), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n16068), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12649) );
  NAND4_X1 U14241 ( .A1(n12652), .A2(n12651), .A3(n12650), .A4(n12649), .ZN(
        n12659) );
  AOI22_X1 U14242 ( .A1(n12665), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12738), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12653) );
  AOI22_X1 U14243 ( .A1(n16063), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n16068), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12656) );
  AOI22_X1 U14244 ( .A1(n16064), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n13107), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12655) );
  INV_X2 U14245 ( .A(n16061), .ZN(n13049) );
  AOI22_X1 U14246 ( .A1(n10957), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n12866), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12654) );
  NAND4_X1 U14247 ( .A1(n12657), .A2(n12656), .A3(n12655), .A4(n12654), .ZN(
        n12658) );
  AND2_X2 U14248 ( .A1(n12659), .A2(n12658), .ZN(n12763) );
  AOI22_X1 U14249 ( .A1(n12665), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n12738), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12660) );
  AND2_X1 U14250 ( .A1(n12660), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12664) );
  AOI22_X1 U14251 ( .A1(n13107), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n13049), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12663) );
  AOI22_X1 U14252 ( .A1(n16063), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n16068), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12662) );
  AOI22_X1 U14253 ( .A1(n16064), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12866), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12661) );
  NAND4_X1 U14254 ( .A1(n12664), .A2(n12663), .A3(n12662), .A4(n12661), .ZN(
        n12672) );
  AOI22_X1 U14255 ( .A1(n12665), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12738), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12666) );
  AND2_X1 U14256 ( .A1(n12666), .A2(n12681), .ZN(n12670) );
  AOI22_X1 U14257 ( .A1(n16064), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12866), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12669) );
  AOI22_X1 U14258 ( .A1(n13049), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n13107), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12668) );
  AOI22_X1 U14259 ( .A1(n16063), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n16068), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12667) );
  NAND4_X1 U14260 ( .A1(n12670), .A2(n12669), .A3(n12668), .A4(n12667), .ZN(
        n12671) );
  NAND2_X2 U14261 ( .A1(n12672), .A2(n12671), .ZN(n12753) );
  OR2_X2 U14262 ( .A1(n12754), .A2(n12753), .ZN(n12748) );
  INV_X1 U14263 ( .A(n12763), .ZN(n12754) );
  NAND2_X1 U14264 ( .A1(n12754), .A2(n12753), .ZN(n12768) );
  AOI22_X1 U14265 ( .A1(n16064), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12866), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12676) );
  AOI22_X1 U14266 ( .A1(n16063), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n16068), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12675) );
  AOI22_X1 U14267 ( .A1(n16067), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n12738), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12674) );
  AOI22_X1 U14268 ( .A1(n13049), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n13107), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12673) );
  AOI22_X1 U14269 ( .A1(n16064), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n12866), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12680) );
  AOI22_X1 U14270 ( .A1(n16063), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n16068), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12679) );
  AOI22_X1 U14271 ( .A1(n16067), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n12738), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12678) );
  AOI22_X1 U14272 ( .A1(n13049), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n13107), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12677) );
  AOI22_X1 U14273 ( .A1(n13107), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n13049), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12685) );
  AOI22_X1 U14274 ( .A1(n16064), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12866), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12684) );
  AOI22_X1 U14275 ( .A1(n16067), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n12738), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12683) );
  AOI22_X1 U14276 ( .A1(n16063), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n16068), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12682) );
  AOI22_X1 U14277 ( .A1(n13107), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n13049), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12689) );
  AOI22_X1 U14278 ( .A1(n16063), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n16068), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12688) );
  AOI22_X1 U14279 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n12866), .B1(
        n16064), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12687) );
  AOI22_X1 U14280 ( .A1(n16067), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12738), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12686) );
  AOI22_X1 U14281 ( .A1(n16067), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12738), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12693) );
  AOI22_X1 U14282 ( .A1(n13107), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n10957), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12692) );
  AOI22_X1 U14283 ( .A1(n16063), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n16068), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12691) );
  AOI22_X1 U14284 ( .A1(n16064), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12866), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12690) );
  NAND4_X1 U14285 ( .A1(n12693), .A2(n12692), .A3(n12691), .A4(n12690), .ZN(
        n12694) );
  AOI22_X1 U14286 ( .A1(n16064), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12866), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12698) );
  AOI22_X1 U14287 ( .A1(n16063), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n16068), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12697) );
  AOI22_X1 U14288 ( .A1(n13107), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n16067), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12696) );
  AOI22_X1 U14289 ( .A1(n13049), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n12738), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12695) );
  NAND4_X1 U14290 ( .A1(n12698), .A2(n12697), .A3(n12696), .A4(n12695), .ZN(
        n12699) );
  NAND2_X1 U14291 ( .A1(n13998), .A2(n14008), .ZN(n12706) );
  NAND2_X2 U14292 ( .A1(n12763), .A2(n12753), .ZN(n12769) );
  INV_X1 U14293 ( .A(n12732), .ZN(n12703) );
  AOI22_X1 U14294 ( .A1(n16064), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12866), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12710) );
  AOI22_X1 U14295 ( .A1(n16063), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n16068), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12709) );
  AOI22_X1 U14296 ( .A1(n13107), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n13049), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12708) );
  AOI22_X1 U14297 ( .A1(n16058), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n12738), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12707) );
  NAND4_X1 U14298 ( .A1(n12710), .A2(n12709), .A3(n12708), .A4(n12707), .ZN(
        n12711) );
  NAND2_X1 U14299 ( .A1(n12711), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12718) );
  AOI22_X1 U14300 ( .A1(n13107), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n10957), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12715) );
  AOI22_X1 U14301 ( .A1(n16063), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n16068), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12714) );
  AOI22_X1 U14302 ( .A1(n16064), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n12866), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12713) );
  AOI22_X1 U14303 ( .A1(n16058), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n12738), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12712) );
  NAND4_X1 U14304 ( .A1(n12715), .A2(n12714), .A3(n12713), .A4(n12712), .ZN(
        n12716) );
  NAND2_X1 U14305 ( .A1(n12716), .A2(n12681), .ZN(n12717) );
  NAND2_X2 U14306 ( .A1(n12718), .A2(n12717), .ZN(n13265) );
  AOI22_X1 U14307 ( .A1(n16064), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12866), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12722) );
  AOI22_X1 U14308 ( .A1(n16063), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n16068), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12721) );
  AOI22_X1 U14309 ( .A1(n13107), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n10957), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12720) );
  AOI22_X1 U14310 ( .A1(n16058), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n12738), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12719) );
  NAND4_X1 U14311 ( .A1(n12722), .A2(n12721), .A3(n12720), .A4(n12719), .ZN(
        n12723) );
  NAND2_X1 U14312 ( .A1(n12723), .A2(n12681), .ZN(n12730) );
  AOI22_X1 U14313 ( .A1(n16064), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12866), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12727) );
  AOI22_X1 U14314 ( .A1(n16063), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n16068), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12726) );
  AOI22_X1 U14315 ( .A1(n13107), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n13049), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12725) );
  AOI22_X1 U14316 ( .A1(n16058), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n12738), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12724) );
  NAND4_X1 U14317 ( .A1(n12727), .A2(n12726), .A3(n12725), .A4(n12724), .ZN(
        n12728) );
  NAND2_X2 U14318 ( .A1(n13265), .A2(n14994), .ZN(n13184) );
  OAI21_X1 U14319 ( .B1(n12751), .B2(n12753), .A(n12771), .ZN(n12731) );
  AOI22_X1 U14320 ( .A1(n16063), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n16068), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12735) );
  AOI22_X1 U14321 ( .A1(n13107), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n13049), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12734) );
  AOI22_X1 U14322 ( .A1(n16067), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n12738), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12733) );
  NAND4_X1 U14323 ( .A1(n12736), .A2(n12735), .A3(n12734), .A4(n12733), .ZN(
        n12737) );
  AOI22_X1 U14324 ( .A1(n16064), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12866), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12742) );
  AOI22_X1 U14325 ( .A1(n16063), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n16068), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12741) );
  AOI22_X1 U14326 ( .A1(n13107), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n13049), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12740) );
  AOI22_X1 U14327 ( .A1(n16067), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12738), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12739) );
  NAND4_X1 U14328 ( .A1(n12742), .A2(n12741), .A3(n12740), .A4(n12739), .ZN(
        n12743) );
  NAND2_X1 U14329 ( .A1(n12743), .A2(n12681), .ZN(n12744) );
  AND2_X1 U14330 ( .A1(n12763), .A2(n12746), .ZN(n12750) );
  NAND2_X1 U14331 ( .A1(n12749), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12762) );
  AND2_X1 U14332 ( .A1(n14008), .A2(n12862), .ZN(n12752) );
  NAND3_X1 U14333 ( .A1(n12750), .A2(n12755), .A3(n12752), .ZN(n14998) );
  NAND3_X1 U14334 ( .A1(n14998), .A2(n19559), .A3(n13265), .ZN(n12759) );
  NAND2_X1 U14335 ( .A1(n12759), .A2(n12758), .ZN(n13551) );
  INV_X1 U14336 ( .A(n13551), .ZN(n12761) );
  NAND2_X1 U14337 ( .A1(n14994), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n13228) );
  NAND2_X1 U14338 ( .A1(n12761), .A2(n12760), .ZN(n12794) );
  NAND2_X1 U14339 ( .A1(n12762), .A2(n12794), .ZN(n12808) );
  NAND2_X1 U14340 ( .A1(n12808), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12767) );
  NOR2_X1 U14341 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n12823) );
  INV_X1 U14342 ( .A(n12823), .ZN(n18627) );
  NAND2_X1 U14343 ( .A1(n12767), .A2(n12766), .ZN(n12783) );
  INV_X1 U14344 ( .A(n12783), .ZN(n12781) );
  NOR2_X1 U14345 ( .A1(n12768), .A2(n13265), .ZN(n12770) );
  INV_X1 U14346 ( .A(n12769), .ZN(n13250) );
  INV_X1 U14347 ( .A(n12771), .ZN(n12774) );
  INV_X1 U14348 ( .A(n12772), .ZN(n12773) );
  AND2_X2 U14349 ( .A1(n12776), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12810) );
  INV_X1 U14350 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n12779) );
  INV_X1 U14351 ( .A(P2_EBX_REG_1__SCAN_IN), .ZN(n12777) );
  NAND2_X1 U14352 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n12778) );
  AOI21_X2 U14353 ( .B1(n12810), .B2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n12780), .ZN(n12782) );
  NAND2_X1 U14354 ( .A1(n12781), .A2(n12782), .ZN(n12807) );
  INV_X1 U14355 ( .A(n12782), .ZN(n12784) );
  NAND2_X1 U14356 ( .A1(n12784), .A2(n12783), .ZN(n12785) );
  NAND2_X1 U14357 ( .A1(n13498), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12786) );
  NOR2_X1 U14358 ( .A1(n12786), .A2(n14000), .ZN(n12789) );
  INV_X1 U14359 ( .A(n12790), .ZN(n12791) );
  AOI22_X1 U14360 ( .A1(n12791), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(n12823), 
        .B2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n12792) );
  NAND2_X1 U14361 ( .A1(n12793), .A2(n12792), .ZN(n12848) );
  NAND2_X1 U14362 ( .A1(n12810), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12806) );
  INV_X1 U14363 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n18102) );
  OAI21_X1 U14364 ( .B1(n15436), .B2(n18102), .A(n12794), .ZN(n12797) );
  INV_X1 U14365 ( .A(P2_EBX_REG_0__SCAN_IN), .ZN(n18103) );
  NAND2_X1 U14366 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n12795) );
  OAI211_X1 U14367 ( .C1(n12787), .C2(n18103), .A(n18627), .B(n12795), .ZN(
        n12796) );
  NOR2_X1 U14368 ( .A1(n12797), .A2(n12796), .ZN(n12805) );
  INV_X1 U14369 ( .A(n12798), .ZN(n12799) );
  NAND2_X1 U14370 ( .A1(n12800), .A2(n12799), .ZN(n12802) );
  NAND2_X1 U14371 ( .A1(n12802), .A2(n12801), .ZN(n12803) );
  NAND2_X1 U14372 ( .A1(n12803), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12804) );
  NAND3_X1 U14373 ( .A1(n12806), .A2(n12805), .A3(n12804), .ZN(n12847) );
  OAI21_X1 U14374 ( .B1(n19231), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n16719), 
        .ZN(n12809) );
  NAND2_X1 U14375 ( .A1(n12811), .A2(P2_EBX_REG_2__SCAN_IN), .ZN(n12816) );
  INV_X1 U14376 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n12813) );
  NAND2_X1 U14377 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n12812) );
  OAI21_X1 U14378 ( .B1(n10963), .B2(n12813), .A(n12812), .ZN(n12814) );
  NAND2_X1 U14379 ( .A1(n12816), .A2(n12815), .ZN(n12817) );
  NAND2_X1 U14380 ( .A1(n12818), .A2(n12819), .ZN(n12821) );
  INV_X1 U14381 ( .A(n12818), .ZN(n12820) );
  NAND2_X1 U14382 ( .A1(n12808), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12825) );
  NAND2_X1 U14383 ( .A1(n12823), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n12824) );
  INV_X1 U14384 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n18602) );
  AOI22_X1 U14385 ( .A1(n15227), .A2(P2_EBX_REG_3__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12827) );
  NAND2_X1 U14386 ( .A1(n15440), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n12826) );
  BUF_X1 U14387 ( .A(n14816), .Z(n13704) );
  NAND2_X1 U14388 ( .A1(n13554), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n14078) );
  OR2_X2 U14389 ( .A1(n13704), .A2(n14078), .ZN(n12832) );
  NAND2_X1 U14390 ( .A1(n19232), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n12842) );
  INV_X1 U14391 ( .A(n12842), .ZN(n12829) );
  NAND2_X1 U14392 ( .A1(n12829), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n16666) );
  NOR2_X2 U14393 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19316) );
  NAND2_X1 U14394 ( .A1(n12842), .A2(n19200), .ZN(n12830) );
  AND3_X1 U14395 ( .A1(n16666), .A2(n19316), .A3(n12830), .ZN(n19175) );
  AOI21_X1 U14396 ( .B1(n12853), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n19175), .ZN(n12831) );
  NAND2_X1 U14397 ( .A1(n12832), .A2(n12831), .ZN(n12836) );
  INV_X1 U14398 ( .A(n12836), .ZN(n12833) );
  NAND2_X1 U14399 ( .A1(n11477), .A2(n12828), .ZN(n13063) );
  INV_X1 U14400 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n16683) );
  OR2_X1 U14401 ( .A1(n13063), .A2(n16683), .ZN(n12834) );
  NAND2_X1 U14402 ( .A1(n12833), .A2(n12834), .ZN(n12837) );
  INV_X1 U14403 ( .A(n12834), .ZN(n12835) );
  NAND2_X1 U14404 ( .A1(n12836), .A2(n12835), .ZN(n12864) );
  INV_X1 U14405 ( .A(n12839), .ZN(n12840) );
  XNOR2_X2 U14406 ( .A(n12838), .B(n12840), .ZN(n14807) );
  INV_X1 U14407 ( .A(n19316), .ZN(n19326) );
  INV_X1 U14408 ( .A(n19232), .ZN(n19294) );
  NAND2_X1 U14409 ( .A1(n19294), .A2(n19231), .ZN(n12841) );
  NAND2_X1 U14410 ( .A1(n12842), .A2(n12841), .ZN(n19176) );
  NOR2_X1 U14411 ( .A1(n19326), .A2(n19176), .ZN(n12843) );
  AOI21_X1 U14412 ( .B1(n12853), .B2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n12843), .ZN(n12844) );
  INV_X1 U14413 ( .A(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n19601) );
  NOR2_X1 U14414 ( .A1(n13063), .A2(n19601), .ZN(n12845) );
  AOI22_X1 U14415 ( .A1(n12853), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n19332), .B2(n19323), .ZN(n12850) );
  INV_X1 U14416 ( .A(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n19651) );
  INV_X1 U14417 ( .A(n14078), .ZN(n12856) );
  NAND2_X1 U14418 ( .A1(n12853), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12854) );
  NAND2_X1 U14419 ( .A1(n19323), .A2(n19296), .ZN(n19280) );
  AND2_X1 U14420 ( .A1(n19294), .A2(n19280), .ZN(n19248) );
  NAND2_X1 U14421 ( .A1(n19332), .A2(n19248), .ZN(n19308) );
  NAND2_X1 U14422 ( .A1(n12854), .A2(n19308), .ZN(n12855) );
  NAND2_X1 U14423 ( .A1(n13646), .A2(n13645), .ZN(n12860) );
  INV_X1 U14424 ( .A(n12857), .ZN(n12858) );
  NAND2_X1 U14425 ( .A1(n12862), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n12863) );
  AND2_X2 U14426 ( .A1(n16064), .A2(n12681), .ZN(n12884) );
  AND2_X2 U14427 ( .A1(n16062), .A2(n12681), .ZN(n13360) );
  AOI22_X1 U14428 ( .A1(n12884), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n13360), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12871) );
  AND2_X2 U14429 ( .A1(n16064), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13484) );
  NOR2_X1 U14430 ( .A1(n12867), .A2(n12681), .ZN(n13482) );
  AOI22_X1 U14431 ( .A1(n13484), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n13354), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12870) );
  AND2_X2 U14432 ( .A1(n16062), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13280) );
  AOI22_X1 U14433 ( .A1(n13280), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12898), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12869) );
  AND2_X2 U14434 ( .A1(n16058), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12954) );
  AOI22_X1 U14435 ( .A1(n12954), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n13366), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12868) );
  NAND4_X1 U14436 ( .A1(n12871), .A2(n12870), .A3(n12869), .A4(n12868), .ZN(
        n12881) );
  AND2_X2 U14437 ( .A1(n16057), .A2(n12681), .ZN(n13361) );
  AOI22_X1 U14438 ( .A1(n12885), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n13361), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12879) );
  AOI22_X1 U14439 ( .A1(n13343), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n13368), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12878) );
  AND2_X1 U14440 ( .A1(n12645), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12872) );
  AND2_X2 U14441 ( .A1(n13041), .A2(n12872), .ZN(n13373) );
  AOI22_X1 U14442 ( .A1(n13373), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n12903), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12877) );
  AND2_X1 U14443 ( .A1(n13211), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12874) );
  AND2_X1 U14444 ( .A1(n13041), .A2(n12875), .ZN(n12891) );
  AOI22_X1 U14445 ( .A1(n12890), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n12891), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12876) );
  NAND4_X1 U14446 ( .A1(n12879), .A2(n12878), .A3(n12877), .A4(n12876), .ZN(
        n12880) );
  INV_X1 U14447 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n19348) );
  NAND2_X1 U14448 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n13883) );
  NOR2_X1 U14449 ( .A1(n19348), .A2(n13883), .ZN(n13840) );
  AND2_X1 U14450 ( .A1(n13842), .A2(n13840), .ZN(n12882) );
  INV_X1 U14451 ( .A(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n19506) );
  NOR2_X1 U14452 ( .A1(n13063), .A2(n19506), .ZN(n13891) );
  AOI22_X1 U14453 ( .A1(n12884), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n13360), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12889) );
  INV_X1 U14454 ( .A(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n19609) );
  AOI22_X1 U14455 ( .A1(n13484), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n13354), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12888) );
  AOI22_X1 U14456 ( .A1(n13280), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12898), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12887) );
  AOI22_X1 U14457 ( .A1(n12885), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n13361), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12886) );
  NAND4_X1 U14458 ( .A1(n12889), .A2(n12888), .A3(n12887), .A4(n12886), .ZN(
        n12897) );
  AOI22_X1 U14459 ( .A1(n12954), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n13366), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12895) );
  AOI22_X1 U14460 ( .A1(n13343), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n13368), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12894) );
  AOI22_X1 U14461 ( .A1(n13373), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n12903), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12893) );
  AOI22_X1 U14462 ( .A1(n12890), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n12891), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12892) );
  NAND4_X1 U14463 ( .A1(n12895), .A2(n12894), .A3(n12893), .A4(n12892), .ZN(
        n12896) );
  AOI22_X1 U14464 ( .A1(n13360), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n13280), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12902) );
  AOI22_X1 U14465 ( .A1(n13484), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n13354), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12901) );
  AOI22_X1 U14466 ( .A1(n12884), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12898), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12900) );
  AOI22_X1 U14467 ( .A1(n12954), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n13361), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12899) );
  NAND4_X1 U14468 ( .A1(n12902), .A2(n12901), .A3(n12900), .A4(n12899), .ZN(
        n12909) );
  AOI22_X1 U14469 ( .A1(n13366), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12885), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12907) );
  AOI22_X1 U14470 ( .A1(n13343), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n13368), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12906) );
  AOI22_X1 U14471 ( .A1(n13373), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n12903), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12905) );
  AOI22_X1 U14472 ( .A1(n12890), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n12891), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12904) );
  NAND4_X1 U14473 ( .A1(n12907), .A2(n12906), .A3(n12905), .A4(n12904), .ZN(
        n12908) );
  AOI22_X1 U14474 ( .A1(n12884), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n13360), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12913) );
  AOI22_X1 U14475 ( .A1(n13484), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n13354), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12912) );
  AOI22_X1 U14476 ( .A1(n13280), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12898), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12911) );
  AOI22_X1 U14477 ( .A1(n12885), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n13361), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12910) );
  NAND4_X1 U14478 ( .A1(n12913), .A2(n12912), .A3(n12911), .A4(n12910), .ZN(
        n12919) );
  AOI22_X1 U14479 ( .A1(n12954), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n13366), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12917) );
  AOI22_X1 U14480 ( .A1(n13343), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n13368), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12916) );
  AOI22_X1 U14481 ( .A1(n13373), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n12903), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12915) );
  AOI22_X1 U14482 ( .A1(n12890), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n12891), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12914) );
  NAND4_X1 U14483 ( .A1(n12917), .A2(n12916), .A3(n12915), .A4(n12914), .ZN(
        n12918) );
  AOI22_X1 U14484 ( .A1(n12884), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n13360), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12923) );
  AOI22_X1 U14485 ( .A1(n13484), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n13354), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12922) );
  AOI22_X1 U14486 ( .A1(n13280), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n12898), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12921) );
  AOI22_X1 U14487 ( .A1(n12885), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n13361), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12920) );
  NAND4_X1 U14488 ( .A1(n12923), .A2(n12922), .A3(n12921), .A4(n12920), .ZN(
        n12929) );
  AOI22_X1 U14489 ( .A1(n12954), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n13366), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12927) );
  AOI22_X1 U14490 ( .A1(n13343), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n13368), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12926) );
  AOI22_X1 U14491 ( .A1(n13373), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n12903), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12925) );
  AOI22_X1 U14492 ( .A1(n12890), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n12891), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12924) );
  NAND4_X1 U14493 ( .A1(n12927), .A2(n12926), .A3(n12925), .A4(n12924), .ZN(
        n12928) );
  AOI22_X1 U14494 ( .A1(n12884), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n13360), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12933) );
  AOI22_X1 U14495 ( .A1(n13484), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n13354), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12932) );
  AOI22_X1 U14496 ( .A1(n13280), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12898), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12931) );
  AOI22_X1 U14497 ( .A1(n12885), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n13361), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12930) );
  NAND4_X1 U14498 ( .A1(n12933), .A2(n12932), .A3(n12931), .A4(n12930), .ZN(
        n12939) );
  AOI22_X1 U14499 ( .A1(n12954), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n13366), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12937) );
  AOI22_X1 U14500 ( .A1(n13343), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n13368), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12936) );
  AOI22_X1 U14501 ( .A1(n13373), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n12903), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12935) );
  AOI22_X1 U14502 ( .A1(n12890), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n12891), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12934) );
  NAND4_X1 U14503 ( .A1(n12937), .A2(n12936), .A3(n12935), .A4(n12934), .ZN(
        n12938) );
  AOI22_X1 U14504 ( .A1(n13484), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n13280), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12943) );
  AOI22_X1 U14505 ( .A1(n12884), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n13360), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12942) );
  AOI22_X1 U14506 ( .A1(n12898), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n13354), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12941) );
  AOI22_X1 U14507 ( .A1(n13366), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n13361), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12940) );
  NAND4_X1 U14508 ( .A1(n12943), .A2(n12942), .A3(n12941), .A4(n12940), .ZN(
        n12949) );
  AOI22_X1 U14509 ( .A1(n12954), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n12885), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12947) );
  AOI22_X1 U14510 ( .A1(n13343), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n13368), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12946) );
  AOI22_X1 U14511 ( .A1(n12890), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n13373), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12945) );
  AOI22_X1 U14512 ( .A1(n12891), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12903), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12944) );
  NAND4_X1 U14513 ( .A1(n12947), .A2(n12946), .A3(n12945), .A4(n12944), .ZN(
        n12948) );
  AOI22_X1 U14514 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n13360), .B1(
        n12884), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12953) );
  AOI22_X1 U14515 ( .A1(n13484), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__7__SCAN_IN), .B2(n13354), .ZN(n12952) );
  AOI22_X1 U14516 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n13280), .B1(
        n12898), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12951) );
  AOI22_X1 U14517 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n13361), .B1(
        n12885), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12950) );
  NAND4_X1 U14518 ( .A1(n12953), .A2(n12952), .A3(n12951), .A4(n12950), .ZN(
        n12960) );
  AOI22_X1 U14519 ( .A1(n12954), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n13366), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12958) );
  AOI22_X1 U14520 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n13368), .B1(
        n13343), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12957) );
  AOI22_X1 U14521 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n13373), .B1(
        n12903), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12956) );
  AOI22_X1 U14522 ( .A1(n12890), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n12891), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12955) );
  NAND4_X1 U14523 ( .A1(n12958), .A2(n12957), .A3(n12956), .A4(n12955), .ZN(
        n12959) );
  NOR2_X1 U14524 ( .A1(n12960), .A2(n12959), .ZN(n14795) );
  OR2_X2 U14525 ( .A1(n14794), .A2(n14795), .ZN(n14940) );
  AOI22_X1 U14526 ( .A1(n12884), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n13360), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12964) );
  AOI22_X1 U14527 ( .A1(n13484), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n13354), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12963) );
  AOI22_X1 U14528 ( .A1(n13280), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n12898), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12962) );
  AOI22_X1 U14529 ( .A1(n12885), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n13361), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12961) );
  NAND4_X1 U14530 ( .A1(n12964), .A2(n12963), .A3(n12962), .A4(n12961), .ZN(
        n12970) );
  AOI22_X1 U14531 ( .A1(n12954), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n13366), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12968) );
  AOI22_X1 U14532 ( .A1(n13343), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n13368), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12967) );
  AOI22_X1 U14533 ( .A1(n13373), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n12903), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12966) );
  AOI22_X1 U14534 ( .A1(n12890), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12891), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12965) );
  NAND4_X1 U14535 ( .A1(n12968), .A2(n12967), .A3(n12966), .A4(n12965), .ZN(
        n12969) );
  NOR2_X1 U14536 ( .A1(n12970), .A2(n12969), .ZN(n14939) );
  AOI22_X1 U14537 ( .A1(n12884), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n13360), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12974) );
  AOI22_X1 U14538 ( .A1(n13484), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n13354), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12973) );
  AOI22_X1 U14539 ( .A1(n13280), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n12898), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12972) );
  AOI22_X1 U14540 ( .A1(n12885), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n13361), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12971) );
  NAND4_X1 U14541 ( .A1(n12974), .A2(n12973), .A3(n12972), .A4(n12971), .ZN(
        n12980) );
  AOI22_X1 U14542 ( .A1(n12954), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n13366), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12978) );
  AOI22_X1 U14543 ( .A1(n13343), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n13368), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12977) );
  AOI22_X1 U14544 ( .A1(n13373), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n12903), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12976) );
  AOI22_X1 U14545 ( .A1(n12890), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n12891), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12975) );
  NAND4_X1 U14546 ( .A1(n12978), .A2(n12977), .A3(n12976), .A4(n12975), .ZN(
        n12979) );
  NOR2_X1 U14547 ( .A1(n12980), .A2(n12979), .ZN(n15056) );
  AOI22_X1 U14548 ( .A1(n12884), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n13360), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12984) );
  AOI22_X1 U14549 ( .A1(n13484), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n13354), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12983) );
  AOI22_X1 U14550 ( .A1(n13280), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n12898), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12982) );
  AOI22_X1 U14551 ( .A1(n12885), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n13361), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12981) );
  NAND4_X1 U14552 ( .A1(n12984), .A2(n12983), .A3(n12982), .A4(n12981), .ZN(
        n12990) );
  AOI22_X1 U14553 ( .A1(n12954), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n13366), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12988) );
  AOI22_X1 U14554 ( .A1(n13343), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n13368), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12987) );
  AOI22_X1 U14555 ( .A1(n13373), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n12903), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12986) );
  AOI22_X1 U14556 ( .A1(n12890), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12891), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12985) );
  NAND4_X1 U14557 ( .A1(n12988), .A2(n12987), .A3(n12986), .A4(n12985), .ZN(
        n12989) );
  OR2_X1 U14558 ( .A1(n12990), .A2(n12989), .ZN(n16159) );
  AOI22_X1 U14559 ( .A1(n12884), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n13360), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12994) );
  AOI22_X1 U14560 ( .A1(n13484), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n13354), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12993) );
  AOI22_X1 U14561 ( .A1(n13280), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12898), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12992) );
  AOI22_X1 U14562 ( .A1(n12885), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n13361), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12991) );
  NAND4_X1 U14563 ( .A1(n12994), .A2(n12993), .A3(n12992), .A4(n12991), .ZN(
        n13000) );
  AOI22_X1 U14564 ( .A1(n12954), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n13366), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12998) );
  AOI22_X1 U14565 ( .A1(n13343), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n13368), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12997) );
  AOI22_X1 U14566 ( .A1(n13373), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n12903), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12996) );
  AOI22_X1 U14567 ( .A1(n12890), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12891), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12995) );
  NAND4_X1 U14568 ( .A1(n12998), .A2(n12997), .A3(n12996), .A4(n12995), .ZN(
        n12999) );
  NOR2_X1 U14569 ( .A1(n13000), .A2(n12999), .ZN(n16152) );
  AOI22_X1 U14570 ( .A1(n12884), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n13360), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n13004) );
  AOI22_X1 U14571 ( .A1(n13484), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n13354), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n13003) );
  AOI22_X1 U14572 ( .A1(n13280), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n12898), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n13002) );
  AOI22_X1 U14573 ( .A1(n12885), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n13361), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n13001) );
  NAND4_X1 U14574 ( .A1(n13004), .A2(n13003), .A3(n13002), .A4(n13001), .ZN(
        n13010) );
  AOI22_X1 U14575 ( .A1(n12954), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n13366), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n13008) );
  AOI22_X1 U14576 ( .A1(n13343), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n13368), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n13007) );
  AOI22_X1 U14577 ( .A1(n13373), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n12903), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n13006) );
  AOI22_X1 U14578 ( .A1(n12890), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n12891), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n13005) );
  NAND4_X1 U14579 ( .A1(n13008), .A2(n13007), .A3(n13006), .A4(n13005), .ZN(
        n13009) );
  OR2_X1 U14580 ( .A1(n13010), .A2(n13009), .ZN(n16145) );
  AOI22_X1 U14581 ( .A1(n12884), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n13360), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n13014) );
  AOI22_X1 U14582 ( .A1(n13484), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n13354), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n13013) );
  AOI22_X1 U14583 ( .A1(n12885), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n13361), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n13012) );
  AOI22_X1 U14584 ( .A1(n13280), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12898), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n13011) );
  NAND4_X1 U14585 ( .A1(n13014), .A2(n13013), .A3(n13012), .A4(n13011), .ZN(
        n13020) );
  AOI22_X1 U14586 ( .A1(n12954), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n13366), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n13018) );
  AOI22_X1 U14587 ( .A1(n13343), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n13368), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n13017) );
  AOI22_X1 U14588 ( .A1(n13373), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n12903), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n13016) );
  AOI22_X1 U14589 ( .A1(n12891), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12890), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n13015) );
  NAND4_X1 U14590 ( .A1(n13018), .A2(n13017), .A3(n13016), .A4(n13015), .ZN(
        n13019) );
  NOR2_X1 U14591 ( .A1(n13020), .A2(n13019), .ZN(n16140) );
  AOI22_X1 U14592 ( .A1(n12884), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n13360), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n13024) );
  AOI22_X1 U14593 ( .A1(n13484), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n13354), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n13023) );
  AOI22_X1 U14594 ( .A1(n13280), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n12898), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n13022) );
  AOI22_X1 U14595 ( .A1(n12885), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n13361), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n13021) );
  NAND4_X1 U14596 ( .A1(n13024), .A2(n13023), .A3(n13022), .A4(n13021), .ZN(
        n13030) );
  AOI22_X1 U14597 ( .A1(n12954), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n13366), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n13028) );
  AOI22_X1 U14598 ( .A1(n13343), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n13368), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n13027) );
  AOI22_X1 U14599 ( .A1(n13373), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n12903), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n13026) );
  AOI22_X1 U14600 ( .A1(n12890), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12891), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n13025) );
  NAND4_X1 U14601 ( .A1(n13028), .A2(n13027), .A3(n13026), .A4(n13025), .ZN(
        n13029) );
  OR2_X1 U14602 ( .A1(n13030), .A2(n13029), .ZN(n16132) );
  AOI22_X1 U14603 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n12884), .B1(
        n13360), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n13034) );
  AOI22_X1 U14604 ( .A1(n13484), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__7__SCAN_IN), .B2(n13354), .ZN(n13033) );
  AOI22_X1 U14605 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n13280), .B1(
        n12898), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n13032) );
  AOI22_X1 U14606 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n13361), .B1(
        n12885), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n13031) );
  NAND4_X1 U14607 ( .A1(n13034), .A2(n13033), .A3(n13032), .A4(n13031), .ZN(
        n13040) );
  AOI22_X1 U14608 ( .A1(n12954), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n13366), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n13038) );
  AOI22_X1 U14609 ( .A1(n13343), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n13368), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n13037) );
  AOI22_X1 U14610 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n12903), .B1(
        n13373), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n13036) );
  AOI22_X1 U14611 ( .A1(n12890), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n12891), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n13035) );
  NAND4_X1 U14612 ( .A1(n13038), .A2(n13037), .A3(n13036), .A4(n13035), .ZN(
        n13039) );
  NOR2_X1 U14613 ( .A1(n13040), .A2(n13039), .ZN(n13059) );
  AOI22_X1 U14614 ( .A1(n16062), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n13107), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n13048) );
  AND2_X1 U14615 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13042) );
  OR2_X1 U14616 ( .A1(n13042), .A2(n13041), .ZN(n16070) );
  INV_X1 U14617 ( .A(n16070), .ZN(n13123) );
  NAND2_X1 U14618 ( .A1(n16057), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n13044) );
  NAND2_X1 U14619 ( .A1(n16063), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n13043) );
  AND3_X1 U14620 ( .A1(n13123), .A2(n13044), .A3(n13043), .ZN(n13047) );
  AOI22_X1 U14621 ( .A1(n16064), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n16068), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n13046) );
  AOI22_X1 U14622 ( .A1(n16058), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n10957), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n13045) );
  NAND4_X1 U14623 ( .A1(n13048), .A2(n13047), .A3(n13046), .A4(n13045), .ZN(
        n13057) );
  AOI22_X1 U14624 ( .A1(n16062), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n13107), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n13055) );
  AOI22_X1 U14625 ( .A1(n16064), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n16068), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n13054) );
  AOI22_X1 U14626 ( .A1(n16058), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n13049), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n13053) );
  NAND2_X1 U14627 ( .A1(n16057), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n13051) );
  NAND2_X1 U14628 ( .A1(n16063), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n13050) );
  AND3_X1 U14629 ( .A1(n13051), .A2(n13050), .A3(n16070), .ZN(n13052) );
  NAND4_X1 U14630 ( .A1(n13055), .A2(n13054), .A3(n13053), .A4(n13052), .ZN(
        n13056) );
  NAND2_X1 U14631 ( .A1(n13057), .A2(n13056), .ZN(n13060) );
  XNOR2_X1 U14632 ( .A(n13059), .B(n13060), .ZN(n16127) );
  INV_X1 U14633 ( .A(n13059), .ZN(n13062) );
  INV_X1 U14634 ( .A(n13060), .ZN(n13061) );
  NAND2_X1 U14635 ( .A1(n13062), .A2(n13061), .ZN(n13079) );
  OAI22_X2 U14636 ( .A1(n16126), .A2(n16127), .B1(n18090), .B2(n13079), .ZN(
        n16122) );
  INV_X1 U14637 ( .A(n13063), .ZN(n13136) );
  INV_X1 U14638 ( .A(n13079), .ZN(n13064) );
  NAND2_X1 U14639 ( .A1(n13136), .A2(n13064), .ZN(n13081) );
  AOI22_X1 U14640 ( .A1(n16064), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n16062), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n13070) );
  AOI22_X1 U14641 ( .A1(n13107), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n16068), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n13069) );
  AOI22_X1 U14642 ( .A1(n13049), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n16057), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n13068) );
  NAND2_X1 U14643 ( .A1(n16058), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n13066) );
  NAND2_X1 U14644 ( .A1(n16063), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n13065) );
  AND3_X1 U14645 ( .A1(n13123), .A2(n13066), .A3(n13065), .ZN(n13067) );
  NAND4_X1 U14646 ( .A1(n13070), .A2(n13069), .A3(n13068), .A4(n13067), .ZN(
        n13078) );
  AOI22_X1 U14647 ( .A1(n16062), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n13107), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n13076) );
  INV_X1 U14648 ( .A(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n19630) );
  AOI22_X1 U14649 ( .A1(n16064), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n16063), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n13075) );
  AOI22_X1 U14650 ( .A1(n16058), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n10957), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n13074) );
  NAND2_X1 U14651 ( .A1(n16057), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n13072) );
  NAND2_X1 U14652 ( .A1(n16068), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n13071) );
  AND3_X1 U14653 ( .A1(n13072), .A2(n13071), .A3(n16070), .ZN(n13073) );
  NAND4_X1 U14654 ( .A1(n13076), .A2(n13075), .A3(n13074), .A4(n13073), .ZN(
        n13077) );
  NAND2_X1 U14655 ( .A1(n13078), .A2(n13077), .ZN(n13080) );
  NOR2_X1 U14656 ( .A1(n13079), .A2(n13080), .ZN(n13096) );
  AOI22_X1 U14657 ( .A1(n13081), .A2(n13080), .B1(n13096), .B2(n18090), .ZN(
        n16121) );
  AOI22_X1 U14658 ( .A1(n16062), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n13107), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n13087) );
  NAND2_X1 U14659 ( .A1(n16057), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n13083) );
  NAND2_X1 U14660 ( .A1(n16063), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n13082) );
  AND3_X1 U14661 ( .A1(n13123), .A2(n13083), .A3(n13082), .ZN(n13086) );
  AOI22_X1 U14662 ( .A1(n16064), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n16068), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n13085) );
  AOI22_X1 U14663 ( .A1(n16058), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n10957), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n13084) );
  NAND4_X1 U14664 ( .A1(n13087), .A2(n13086), .A3(n13085), .A4(n13084), .ZN(
        n13095) );
  AOI22_X1 U14665 ( .A1(n16062), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n13107), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n13093) );
  AOI22_X1 U14666 ( .A1(n16064), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n16068), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n13092) );
  AOI22_X1 U14667 ( .A1(n16058), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n13049), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n13091) );
  NAND2_X1 U14668 ( .A1(n16057), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n13089) );
  NAND2_X1 U14669 ( .A1(n16063), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(
        n13088) );
  AND3_X1 U14670 ( .A1(n13089), .A2(n13088), .A3(n16070), .ZN(n13090) );
  NAND4_X1 U14671 ( .A1(n13093), .A2(n13092), .A3(n13091), .A4(n13090), .ZN(
        n13094) );
  AND2_X1 U14672 ( .A1(n13095), .A2(n13094), .ZN(n13098) );
  NAND2_X1 U14673 ( .A1(n13096), .A2(n13098), .ZN(n13120) );
  OAI211_X1 U14674 ( .C1(n13096), .C2(n13098), .A(n13120), .B(n13136), .ZN(
        n13100) );
  INV_X1 U14675 ( .A(n13098), .ZN(n13099) );
  NOR2_X1 U14676 ( .A1(n18090), .A2(n13099), .ZN(n16115) );
  NAND2_X1 U14677 ( .A1(n16116), .A2(n16115), .ZN(n16114) );
  AOI22_X1 U14678 ( .A1(n16062), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n13107), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n13106) );
  NAND2_X1 U14679 ( .A1(n16057), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n13102) );
  NAND2_X1 U14680 ( .A1(n16063), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n13101) );
  AND3_X1 U14681 ( .A1(n13123), .A2(n13102), .A3(n13101), .ZN(n13105) );
  AOI22_X1 U14682 ( .A1(n16064), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n16068), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n13104) );
  AOI22_X1 U14683 ( .A1(n16058), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n13049), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n13103) );
  NAND4_X1 U14684 ( .A1(n13106), .A2(n13105), .A3(n13104), .A4(n13103), .ZN(
        n13115) );
  AOI22_X1 U14685 ( .A1(n16062), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n13107), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n13113) );
  AOI22_X1 U14686 ( .A1(n16064), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n16068), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n13112) );
  AOI22_X1 U14687 ( .A1(n16058), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n13049), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n13111) );
  NAND2_X1 U14688 ( .A1(n16057), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n13109) );
  NAND2_X1 U14689 ( .A1(n16063), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n13108) );
  AND3_X1 U14690 ( .A1(n13109), .A2(n13108), .A3(n16070), .ZN(n13110) );
  NAND4_X1 U14691 ( .A1(n13113), .A2(n13112), .A3(n13111), .A4(n13110), .ZN(
        n13114) );
  AND2_X1 U14692 ( .A1(n13115), .A2(n13114), .ZN(n13118) );
  XNOR2_X1 U14693 ( .A(n13120), .B(n13118), .ZN(n13116) );
  NAND2_X1 U14694 ( .A1(n19605), .A2(n13118), .ZN(n16109) );
  NOR2_X2 U14695 ( .A1(n16108), .A2(n11486), .ZN(n13156) );
  INV_X1 U14696 ( .A(n13118), .ZN(n13119) );
  NOR2_X1 U14697 ( .A1(n13120), .A2(n13119), .ZN(n13137) );
  AOI22_X1 U14698 ( .A1(n16062), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n13107), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n13127) );
  NAND2_X1 U14699 ( .A1(n16057), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n13122) );
  NAND2_X1 U14700 ( .A1(n16063), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n13121) );
  AND3_X1 U14701 ( .A1(n13123), .A2(n13122), .A3(n13121), .ZN(n13126) );
  AOI22_X1 U14702 ( .A1(n16064), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n16068), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n13125) );
  AOI22_X1 U14703 ( .A1(n16058), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n13049), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n13124) );
  NAND4_X1 U14704 ( .A1(n13127), .A2(n13126), .A3(n13125), .A4(n13124), .ZN(
        n13135) );
  AOI22_X1 U14705 ( .A1(n16062), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n13107), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n13133) );
  AOI22_X1 U14706 ( .A1(n16064), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n16068), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n13132) );
  AOI22_X1 U14707 ( .A1(n16058), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n10957), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n13131) );
  NAND2_X1 U14708 ( .A1(n16057), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n13129) );
  NAND2_X1 U14709 ( .A1(n16063), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n13128) );
  AND3_X1 U14710 ( .A1(n13129), .A2(n13128), .A3(n16070), .ZN(n13130) );
  NAND4_X1 U14711 ( .A1(n13133), .A2(n13132), .A3(n13131), .A4(n13130), .ZN(
        n13134) );
  AND2_X1 U14712 ( .A1(n13135), .A2(n13134), .ZN(n13138) );
  NAND2_X1 U14713 ( .A1(n13137), .A2(n13138), .ZN(n16087) );
  OAI211_X1 U14714 ( .C1(n13137), .C2(n13138), .A(n13136), .B(n16087), .ZN(
        n13155) );
  INV_X1 U14715 ( .A(n13138), .ZN(n13139) );
  NOR2_X1 U14716 ( .A1(n18090), .A2(n13139), .ZN(n16098) );
  AOI22_X1 U14717 ( .A1(n16062), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n13107), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n13141) );
  AOI22_X1 U14718 ( .A1(n16064), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n16068), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n13140) );
  NAND2_X1 U14719 ( .A1(n13141), .A2(n13140), .ZN(n13154) );
  INV_X1 U14720 ( .A(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n13145) );
  AOI21_X1 U14721 ( .B1(n16063), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A(
        n16070), .ZN(n13144) );
  AOI22_X1 U14722 ( .A1(n13049), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n16057), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n13143) );
  OAI211_X1 U14723 ( .C1(n13142), .C2(n13145), .A(n13144), .B(n13143), .ZN(
        n13153) );
  AOI22_X1 U14724 ( .A1(n16062), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n13107), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13147) );
  AOI22_X1 U14725 ( .A1(n16064), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n16063), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n13146) );
  NAND2_X1 U14726 ( .A1(n13147), .A2(n13146), .ZN(n13152) );
  AOI22_X1 U14727 ( .A1(n16058), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n10957), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n13150) );
  NAND2_X1 U14728 ( .A1(n16057), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n13149) );
  NAND2_X1 U14729 ( .A1(n16068), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n13148) );
  NAND4_X1 U14730 ( .A1(n13150), .A2(n16070), .A3(n13149), .A4(n13148), .ZN(
        n13151) );
  OAI22_X1 U14731 ( .A1(n13154), .A2(n13153), .B1(n13152), .B2(n13151), .ZN(
        n13174) );
  INV_X1 U14732 ( .A(n13174), .ZN(n16088) );
  NAND2_X1 U14733 ( .A1(n13156), .A2(n13155), .ZN(n16095) );
  AOI22_X1 U14734 ( .A1(n16064), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n13107), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n13158) );
  AOI22_X1 U14735 ( .A1(n16062), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n16068), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n13157) );
  NAND2_X1 U14736 ( .A1(n13158), .A2(n13157), .ZN(n13170) );
  INV_X1 U14737 ( .A(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n13161) );
  AOI21_X1 U14738 ( .B1(n16063), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A(
        n16070), .ZN(n13160) );
  AOI22_X1 U14739 ( .A1(n10957), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n16057), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n13159) );
  OAI211_X1 U14740 ( .C1(n13142), .C2(n13161), .A(n13160), .B(n13159), .ZN(
        n13169) );
  AOI22_X1 U14741 ( .A1(n16062), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n13107), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n13163) );
  AOI22_X1 U14742 ( .A1(n16064), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n16068), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n13162) );
  NAND2_X1 U14743 ( .A1(n13163), .A2(n13162), .ZN(n13168) );
  AOI22_X1 U14744 ( .A1(n16058), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n13049), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n13166) );
  NAND2_X1 U14745 ( .A1(n16057), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n13165) );
  NAND2_X1 U14746 ( .A1(n16063), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n13164) );
  NAND4_X1 U14747 ( .A1(n13166), .A2(n13165), .A3(n13164), .A4(n16070), .ZN(
        n13167) );
  OAI22_X1 U14748 ( .A1(n13170), .A2(n13169), .B1(n13168), .B2(n13167), .ZN(
        n13171) );
  NOR2_X1 U14749 ( .A1(n13172), .A2(n13171), .ZN(n16052) );
  NAND2_X1 U14750 ( .A1(n13172), .A2(n13171), .ZN(n16053) );
  INV_X1 U14751 ( .A(n16053), .ZN(n13173) );
  NOR2_X1 U14752 ( .A1(n16052), .A2(n13173), .ZN(n13175) );
  NOR3_X1 U14753 ( .A1(n16087), .A2(n19605), .A3(n13174), .ZN(n16054) );
  XNOR2_X1 U14754 ( .A(n13175), .B(n16054), .ZN(n16086) );
  XNOR2_X1 U14755 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n13218) );
  NAND2_X1 U14756 ( .A1(n13218), .A2(n13213), .ZN(n13177) );
  NAND2_X1 U14757 ( .A1(n19296), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13176) );
  NAND2_X1 U14758 ( .A1(n13177), .A2(n13176), .ZN(n13210) );
  XNOR2_X1 U14759 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n13208) );
  NAND2_X1 U14760 ( .A1(n13210), .A2(n13208), .ZN(n13179) );
  NAND2_X1 U14761 ( .A1(n19231), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13178) );
  INV_X1 U14762 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n16722) );
  NOR2_X1 U14763 ( .A1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n16722), .ZN(
        n13182) );
  NAND3_X1 U14764 ( .A1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n13183), .A3(
        n14054), .ZN(n13480) );
  NOR2_X1 U14765 ( .A1(n13480), .A2(n13184), .ZN(n13185) );
  OR2_X1 U14766 ( .A1(n13489), .A2(n13185), .ZN(n13226) );
  AOI22_X1 U14767 ( .A1(n12884), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n13360), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n13189) );
  AOI22_X1 U14768 ( .A1(n13484), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n13354), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n13188) );
  AOI22_X1 U14769 ( .A1(n13280), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12898), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n13187) );
  AOI22_X1 U14770 ( .A1(n12885), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n13361), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n13186) );
  NAND4_X1 U14771 ( .A1(n13189), .A2(n13188), .A3(n13187), .A4(n13186), .ZN(
        n13195) );
  AOI22_X1 U14772 ( .A1(n12954), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n13366), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n13193) );
  AOI22_X1 U14773 ( .A1(n13343), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n13368), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n13192) );
  AOI22_X1 U14774 ( .A1(n13373), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n12903), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n13191) );
  AOI22_X1 U14775 ( .A1(n12890), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n12891), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n13190) );
  NAND4_X1 U14776 ( .A1(n13193), .A2(n13192), .A3(n13191), .A4(n13190), .ZN(
        n13194) );
  MUX2_X1 U14777 ( .A(n13480), .B(n13335), .S(n13498), .Z(n14889) );
  AOI22_X1 U14778 ( .A1(n12884), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n13360), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n13199) );
  AOI22_X1 U14779 ( .A1(n13484), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n13354), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n13198) );
  AOI22_X1 U14780 ( .A1(n13280), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12898), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n13197) );
  AOI22_X1 U14781 ( .A1(n12885), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n13361), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n13196) );
  NAND4_X1 U14782 ( .A1(n13199), .A2(n13198), .A3(n13197), .A4(n13196), .ZN(
        n13205) );
  AOI22_X1 U14783 ( .A1(n12954), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n13366), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n13203) );
  AOI22_X1 U14784 ( .A1(n13343), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n13368), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n13202) );
  AOI22_X1 U14785 ( .A1(n13373), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n12903), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n13201) );
  AOI22_X1 U14786 ( .A1(n12890), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n12891), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n13200) );
  NAND4_X1 U14787 ( .A1(n13203), .A2(n13202), .A3(n13201), .A4(n13200), .ZN(
        n13204) );
  XNOR2_X1 U14788 ( .A(n13207), .B(n13206), .ZN(n13479) );
  MUX2_X1 U14789 ( .A(n14831), .B(n13479), .S(n13184), .Z(n14857) );
  NAND2_X1 U14790 ( .A1(n14889), .A2(n14857), .ZN(n13488) );
  INV_X1 U14791 ( .A(n13208), .ZN(n13209) );
  XNOR2_X1 U14792 ( .A(n13210), .B(n13209), .ZN(n13478) );
  NAND2_X1 U14793 ( .A1(n13184), .A2(n13478), .ZN(n13522) );
  INV_X1 U14794 ( .A(n13522), .ZN(n13223) );
  AOI21_X1 U14795 ( .B1(n13228), .B2(n18090), .A(n13478), .ZN(n13222) );
  INV_X1 U14796 ( .A(n13478), .ZN(n13216) );
  AND2_X1 U14797 ( .A1(n13211), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n13212) );
  NOR2_X1 U14798 ( .A1(n13213), .A2(n13212), .ZN(n13500) );
  INV_X1 U14799 ( .A(n13213), .ZN(n13214) );
  XNOR2_X1 U14800 ( .A(n13214), .B(n13218), .ZN(n13244) );
  OAI21_X1 U14801 ( .B1(n18090), .B2(n13500), .A(n13244), .ZN(n13215) );
  OAI21_X1 U14802 ( .B1(n13216), .B2(n18090), .A(n13215), .ZN(n13217) );
  NAND2_X1 U14803 ( .A1(n13217), .A2(n19676), .ZN(n13220) );
  NAND2_X1 U14804 ( .A1(n13500), .A2(n13218), .ZN(n13486) );
  NAND2_X1 U14805 ( .A1(n13498), .A2(n13486), .ZN(n13219) );
  NAND2_X1 U14806 ( .A1(n13220), .A2(n13219), .ZN(n13221) );
  OAI21_X1 U14807 ( .B1(n13223), .B2(n13222), .A(n13221), .ZN(n13224) );
  AOI22_X1 U14808 ( .A1(n13488), .A2(n13184), .B1(n13479), .B2(n13224), .ZN(
        n13225) );
  NOR2_X1 U14809 ( .A1(n13226), .A2(n13225), .ZN(n13227) );
  MUX2_X1 U14810 ( .A(n14054), .B(n13227), .S(P2_STATE2_REG_0__SCAN_IN), .Z(
        n14995) );
  AND2_X1 U14811 ( .A1(n13489), .A2(n12760), .ZN(n13229) );
  NAND2_X1 U14812 ( .A1(n12769), .A2(n14993), .ZN(n13996) );
  NAND2_X1 U14813 ( .A1(n13996), .A2(n19559), .ZN(n13238) );
  AND2_X1 U14814 ( .A1(n19605), .A2(n14994), .ZN(n13491) );
  NAND2_X1 U14815 ( .A1(n13232), .A2(n13491), .ZN(n13999) );
  NAND2_X1 U14816 ( .A1(n19605), .A2(n14993), .ZN(n13239) );
  AOI21_X1 U14817 ( .B1(n13239), .B2(n19676), .A(n13233), .ZN(n13234) );
  OR2_X1 U14818 ( .A1(n13234), .A2(n14999), .ZN(n13235) );
  NAND4_X1 U14819 ( .A1(n13999), .A2(n14000), .A3(n13236), .A4(n13235), .ZN(
        n13237) );
  AOI21_X1 U14820 ( .B1(n13230), .B2(n13238), .A(n13237), .ZN(n13545) );
  INV_X1 U14821 ( .A(n13239), .ZN(n13240) );
  NAND2_X1 U14822 ( .A1(n16640), .A2(n15030), .ZN(n13547) );
  NAND2_X1 U14823 ( .A1(n13242), .A2(n13241), .ZN(n14005) );
  NAND2_X1 U14824 ( .A1(n13547), .A2(n14005), .ZN(n13243) );
  NAND2_X1 U14825 ( .A1(n13243), .A2(n18099), .ZN(n13249) );
  AND4_X1 U14826 ( .A1(n13480), .A2(n13478), .A3(n13479), .A4(n13244), .ZN(
        n13245) );
  OR2_X1 U14827 ( .A1(n13489), .A2(n13245), .ZN(n15004) );
  NAND2_X1 U14828 ( .A1(n13230), .A2(n11133), .ZN(n15043) );
  INV_X1 U14829 ( .A(n15043), .ZN(n13246) );
  OR2_X1 U14830 ( .A1(n15004), .A2(n13246), .ZN(n14040) );
  INV_X1 U14831 ( .A(n18099), .ZN(n18649) );
  NAND2_X1 U14832 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n21729) );
  NAND2_X1 U14833 ( .A1(n18095), .A2(n14039), .ZN(n13248) );
  NOR2_X2 U14834 ( .A1(n19652), .A2(n13251), .ZN(n19653) );
  NOR4_X1 U14835 ( .A1(P2_ADDRESS_REG_15__SCAN_IN), .A2(
        P2_ADDRESS_REG_13__SCAN_IN), .A3(P2_ADDRESS_REG_12__SCAN_IN), .A4(
        P2_ADDRESS_REG_11__SCAN_IN), .ZN(n13255) );
  NOR4_X1 U14836 ( .A1(P2_ADDRESS_REG_18__SCAN_IN), .A2(
        P2_ADDRESS_REG_17__SCAN_IN), .A3(P2_ADDRESS_REG_14__SCAN_IN), .A4(
        P2_ADDRESS_REG_16__SCAN_IN), .ZN(n13254) );
  NOR4_X1 U14837 ( .A1(P2_ADDRESS_REG_6__SCAN_IN), .A2(
        P2_ADDRESS_REG_5__SCAN_IN), .A3(P2_ADDRESS_REG_4__SCAN_IN), .A4(
        P2_ADDRESS_REG_3__SCAN_IN), .ZN(n13253) );
  NOR4_X1 U14838 ( .A1(P2_ADDRESS_REG_10__SCAN_IN), .A2(
        P2_ADDRESS_REG_7__SCAN_IN), .A3(P2_ADDRESS_REG_9__SCAN_IN), .A4(
        P2_ADDRESS_REG_8__SCAN_IN), .ZN(n13252) );
  NAND4_X1 U14839 ( .A1(n13255), .A2(n13254), .A3(n13253), .A4(n13252), .ZN(
        n13260) );
  NOR4_X1 U14840 ( .A1(P2_ADDRESS_REG_2__SCAN_IN), .A2(
        P2_ADDRESS_REG_1__SCAN_IN), .A3(P2_ADDRESS_REG_26__SCAN_IN), .A4(
        P2_ADDRESS_REG_28__SCAN_IN), .ZN(n13258) );
  NOR4_X1 U14841 ( .A1(P2_ADDRESS_REG_22__SCAN_IN), .A2(
        P2_ADDRESS_REG_21__SCAN_IN), .A3(P2_ADDRESS_REG_20__SCAN_IN), .A4(
        P2_ADDRESS_REG_19__SCAN_IN), .ZN(n13257) );
  NOR4_X1 U14842 ( .A1(P2_ADDRESS_REG_27__SCAN_IN), .A2(
        P2_ADDRESS_REG_25__SCAN_IN), .A3(P2_ADDRESS_REG_24__SCAN_IN), .A4(
        P2_ADDRESS_REG_23__SCAN_IN), .ZN(n13256) );
  INV_X1 U14843 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n19791) );
  NAND4_X1 U14844 ( .A1(n13258), .A2(n13257), .A3(n13256), .A4(n19791), .ZN(
        n13259) );
  AOI22_X1 U14845 ( .A1(n16679), .A2(BUF1_REG_13__SCAN_IN), .B1(
        BUF2_REG_13__SCAN_IN), .B2(n16678), .ZN(n19122) );
  INV_X1 U14846 ( .A(n19122), .ZN(n13433) );
  NAND2_X1 U14847 ( .A1(n15456), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n13262) );
  NAND2_X1 U14848 ( .A1(n13265), .A2(n19203), .ZN(n13409) );
  INV_X2 U14849 ( .A(n13409), .ZN(n13405) );
  AOI22_X1 U14850 ( .A1(n15461), .A2(P2_EAX_REG_17__SCAN_IN), .B1(n13405), 
        .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n13261) );
  NAND2_X1 U14851 ( .A1(n13262), .A2(n13261), .ZN(n15058) );
  NAND2_X1 U14852 ( .A1(n15456), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n13264) );
  AOI22_X1 U14853 ( .A1(n15461), .A2(P2_EAX_REG_16__SCAN_IN), .B1(n13405), 
        .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n13263) );
  NOR2_X1 U14854 ( .A1(n13265), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n13266) );
  AOI22_X1 U14855 ( .A1(n13484), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n13280), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n13270) );
  AOI22_X1 U14856 ( .A1(n12884), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n13354), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13269) );
  AOI22_X1 U14857 ( .A1(n13360), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12898), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n13268) );
  AOI22_X1 U14858 ( .A1(n13366), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n13361), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n13267) );
  NAND4_X1 U14859 ( .A1(n13270), .A2(n13269), .A3(n13268), .A4(n13267), .ZN(
        n13276) );
  AOI22_X1 U14860 ( .A1(n12954), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n12885), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n13274) );
  AOI22_X1 U14861 ( .A1(n13343), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n13368), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n13273) );
  AOI22_X1 U14862 ( .A1(n12890), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n13373), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n13272) );
  AOI22_X1 U14863 ( .A1(n12891), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n12903), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n13271) );
  NAND4_X1 U14864 ( .A1(n13274), .A2(n13273), .A3(n13272), .A4(n13271), .ZN(
        n13275) );
  NOR2_X1 U14865 ( .A1(n13276), .A2(n13275), .ZN(n15132) );
  INV_X1 U14866 ( .A(n15132), .ZN(n13353) );
  NAND2_X1 U14867 ( .A1(n13323), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n13279) );
  AOI22_X1 U14868 ( .A1(n13277), .A2(P2_EAX_REG_1__SCAN_IN), .B1(n13405), .B2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n13278) );
  NAND2_X1 U14869 ( .A1(n13279), .A2(n13278), .ZN(n13308) );
  INV_X1 U14870 ( .A(n13308), .ZN(n13294) );
  AOI22_X1 U14871 ( .A1(n12884), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n13484), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n13284) );
  AOI22_X1 U14872 ( .A1(n13360), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n13280), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n13283) );
  AOI22_X1 U14873 ( .A1(n12898), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n13354), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n13282) );
  AOI22_X1 U14874 ( .A1(n12885), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n13361), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n13281) );
  NAND4_X1 U14875 ( .A1(n13284), .A2(n13283), .A3(n13282), .A4(n13281), .ZN(
        n13290) );
  INV_X1 U14876 ( .A(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n19787) );
  AOI22_X1 U14877 ( .A1(n12954), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n13366), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n13288) );
  AOI22_X1 U14878 ( .A1(n13343), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n13368), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n13287) );
  AOI22_X1 U14879 ( .A1(n13373), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n12891), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n13286) );
  AOI22_X1 U14880 ( .A1(n12890), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n12903), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n13285) );
  NAND4_X1 U14881 ( .A1(n13288), .A2(n13287), .A3(n13286), .A4(n13285), .ZN(
        n13289) );
  INV_X1 U14882 ( .A(n13499), .ZN(n13507) );
  OR2_X1 U14883 ( .A1(n13409), .A2(n12769), .ZN(n13321) );
  OAI21_X1 U14884 ( .B1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n19203), .A(
        n11125), .ZN(n13291) );
  NAND2_X1 U14885 ( .A1(n13323), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n13293) );
  INV_X1 U14886 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n13675) );
  NAND2_X1 U14887 ( .A1(n18090), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13292) );
  NAND2_X1 U14888 ( .A1(n13293), .A2(n11025), .ZN(n13670) );
  XNOR2_X1 U14889 ( .A(n13294), .B(n13668), .ZN(n13689) );
  AOI22_X1 U14890 ( .A1(n12884), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n13360), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n13298) );
  AOI22_X1 U14891 ( .A1(n13484), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n13354), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n13297) );
  AOI22_X1 U14892 ( .A1(n13280), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12898), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n13296) );
  AOI22_X1 U14893 ( .A1(n12885), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n13361), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n13295) );
  NAND4_X1 U14894 ( .A1(n13298), .A2(n13297), .A3(n13296), .A4(n13295), .ZN(
        n13304) );
  AOI22_X1 U14895 ( .A1(n12954), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n13366), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n13302) );
  AOI22_X1 U14896 ( .A1(n13343), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n13368), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n13301) );
  AOI22_X1 U14897 ( .A1(n13373), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n12903), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n13300) );
  AOI22_X1 U14898 ( .A1(n12890), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n12891), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n13299) );
  NAND4_X1 U14899 ( .A1(n13302), .A2(n13301), .A3(n13300), .A4(n13299), .ZN(
        n13303) );
  INV_X1 U14900 ( .A(n13518), .ZN(n13511) );
  OR2_X1 U14901 ( .A1(n13408), .A2(n13511), .ZN(n13307) );
  NAND2_X1 U14902 ( .A1(n12769), .A2(n13305), .ZN(n13306) );
  OAI211_X1 U14903 ( .C1(n19203), .C2(n19296), .A(n13307), .B(n13306), .ZN(
        n13688) );
  INV_X1 U14904 ( .A(n13688), .ZN(n13310) );
  NOR2_X1 U14905 ( .A1(n13668), .A2(n13308), .ZN(n13309) );
  AOI22_X1 U14906 ( .A1(n12884), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n13360), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n13314) );
  AOI22_X1 U14907 ( .A1(n13484), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n13354), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n13313) );
  AOI22_X1 U14908 ( .A1(n13280), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12898), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n13312) );
  AOI22_X1 U14909 ( .A1(n12885), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n13361), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n13311) );
  NAND4_X1 U14910 ( .A1(n13314), .A2(n13313), .A3(n13312), .A4(n13311), .ZN(
        n13320) );
  AOI22_X1 U14911 ( .A1(n12954), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n13366), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n13318) );
  AOI22_X1 U14912 ( .A1(n13343), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n13368), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n13317) );
  AOI22_X1 U14913 ( .A1(n13373), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n12903), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n13316) );
  AOI22_X1 U14914 ( .A1(n12890), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n12891), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n13315) );
  NAND4_X1 U14915 ( .A1(n13318), .A2(n13317), .A3(n13316), .A4(n13315), .ZN(
        n13319) );
  INV_X1 U14916 ( .A(n13513), .ZN(n14849) );
  NAND2_X1 U14917 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n13322) );
  OAI211_X1 U14918 ( .C1(n13408), .C2(n14849), .A(n13322), .B(n13321), .ZN(
        n13326) );
  XNOR2_X1 U14919 ( .A(n13327), .B(n13326), .ZN(n13865) );
  NAND2_X1 U14920 ( .A1(n13323), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n13325) );
  AOI22_X1 U14921 ( .A1(n13277), .A2(P2_EAX_REG_2__SCAN_IN), .B1(n13405), .B2(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n13324) );
  NAND2_X1 U14922 ( .A1(n13325), .A2(n13324), .ZN(n13864) );
  NOR2_X1 U14923 ( .A1(n13865), .A2(n13864), .ZN(n13329) );
  NOR2_X1 U14924 ( .A1(n13327), .A2(n13326), .ZN(n13328) );
  NAND2_X1 U14925 ( .A1(n15456), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n13334) );
  INV_X1 U14926 ( .A(n14831), .ZN(n13330) );
  OR2_X1 U14927 ( .A1(n13408), .A2(n13330), .ZN(n13333) );
  AOI22_X1 U14928 ( .A1(n13277), .A2(P2_EAX_REG_3__SCAN_IN), .B1(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n13332) );
  NAND2_X1 U14929 ( .A1(n13405), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13331) );
  NAND4_X1 U14930 ( .A1(n13334), .A2(n13333), .A3(n13332), .A4(n13331), .ZN(
        n14137) );
  NAND2_X1 U14931 ( .A1(n15456), .A2(P2_REIP_REG_4__SCAN_IN), .ZN(n13338) );
  AOI22_X1 U14932 ( .A1(n13277), .A2(P2_EAX_REG_4__SCAN_IN), .B1(n13405), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n13337) );
  INV_X1 U14933 ( .A(n13335), .ZN(n14958) );
  OR2_X1 U14934 ( .A1(n13408), .A2(n14958), .ZN(n13336) );
  AOI22_X1 U14935 ( .A1(n13323), .A2(P2_REIP_REG_5__SCAN_IN), .B1(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n13405), .ZN(n13351) );
  AOI22_X1 U14936 ( .A1(n12884), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n13360), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n13342) );
  AOI22_X1 U14937 ( .A1(n13484), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n13354), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n13341) );
  AOI22_X1 U14938 ( .A1(n13280), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12898), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n13340) );
  AOI22_X1 U14939 ( .A1(n12885), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n13361), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n13339) );
  NAND4_X1 U14940 ( .A1(n13342), .A2(n13341), .A3(n13340), .A4(n13339), .ZN(
        n13349) );
  AOI22_X1 U14941 ( .A1(n12954), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n13366), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n13347) );
  AOI22_X1 U14942 ( .A1(n13343), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n13368), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n13346) );
  AOI22_X1 U14943 ( .A1(n13373), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n12903), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n13345) );
  AOI22_X1 U14944 ( .A1(n12890), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n12891), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13344) );
  NAND4_X1 U14945 ( .A1(n13347), .A2(n13346), .A3(n13345), .A4(n13344), .ZN(
        n13348) );
  AOI22_X1 U14946 ( .A1(n13394), .A2(n15017), .B1(P2_EAX_REG_5__SCAN_IN), .B2(
        n15461), .ZN(n13350) );
  NAND2_X1 U14947 ( .A1(n13351), .A2(n13350), .ZN(n15042) );
  INV_X1 U14948 ( .A(n15041), .ZN(n13352) );
  AOI21_X1 U14949 ( .B1(n13394), .B2(n13353), .A(n13352), .ZN(n13682) );
  AOI222_X1 U14950 ( .A1(P2_REIP_REG_6__SCAN_IN), .A2(n15456), .B1(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n13405), .C1(
        P2_EAX_REG_6__SCAN_IN), .C2(n15461), .ZN(n13681) );
  NAND2_X1 U14951 ( .A1(n12884), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n13359) );
  NAND2_X1 U14952 ( .A1(n13484), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n13358) );
  NAND2_X1 U14953 ( .A1(n12898), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n13357) );
  INV_X1 U14954 ( .A(n13354), .ZN(n13355) );
  INV_X1 U14955 ( .A(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n19150) );
  OR2_X1 U14956 ( .A1(n13355), .A2(n19150), .ZN(n13356) );
  NAND2_X1 U14957 ( .A1(n13360), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n13365) );
  NAND2_X1 U14958 ( .A1(n13280), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n13364) );
  NAND2_X1 U14959 ( .A1(n12885), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n13363) );
  NAND2_X1 U14960 ( .A1(n13361), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n13362) );
  AOI22_X1 U14961 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n12954), .B1(
        n13366), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n13381) );
  INV_X1 U14962 ( .A(n13367), .ZN(n13372) );
  INV_X1 U14963 ( .A(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n19196) );
  INV_X1 U14964 ( .A(n13368), .ZN(n13370) );
  INV_X1 U14965 ( .A(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n13369) );
  OR2_X1 U14966 ( .A1(n13370), .A2(n13369), .ZN(n13371) );
  OAI21_X1 U14967 ( .B1(n13372), .B2(n19196), .A(n13371), .ZN(n13379) );
  NAND2_X1 U14968 ( .A1(n12890), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n13377) );
  NAND2_X1 U14969 ( .A1(n13373), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n13376) );
  NAND2_X1 U14970 ( .A1(n12891), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n13375) );
  NAND2_X1 U14971 ( .A1(n12903), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n13374) );
  NAND4_X1 U14972 ( .A1(n13377), .A2(n13376), .A3(n13375), .A4(n13374), .ZN(
        n13378) );
  NOR2_X1 U14973 ( .A1(n13379), .A2(n13378), .ZN(n13380) );
  AND4_X2 U14974 ( .A1(n13383), .A2(n13382), .A3(n13381), .A4(n13380), .ZN(
        n15139) );
  INV_X1 U14975 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16623) );
  INV_X1 U14976 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n17109) );
  INV_X1 U14977 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n17133) );
  OAI222_X1 U14978 ( .A1(n13409), .A2(n16623), .B1(n13384), .B2(n17109), .C1(
        n15463), .C2(n17133), .ZN(n13684) );
  NAND2_X1 U14979 ( .A1(n15456), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n13388) );
  AOI22_X1 U14980 ( .A1(n13277), .A2(P2_EAX_REG_8__SCAN_IN), .B1(n13405), .B2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n13387) );
  INV_X1 U14981 ( .A(n13842), .ZN(n13385) );
  OR2_X1 U14982 ( .A1(n13408), .A2(n13385), .ZN(n13386) );
  AOI22_X1 U14983 ( .A1(n15456), .A2(P2_REIP_REG_9__SCAN_IN), .B1(n13277), 
        .B2(P2_EAX_REG_9__SCAN_IN), .ZN(n13390) );
  AOI22_X1 U14984 ( .A1(n13394), .A2(n13928), .B1(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n13405), .ZN(n13389) );
  NAND2_X1 U14985 ( .A1(n13390), .A2(n13389), .ZN(n13722) );
  INV_X1 U14986 ( .A(n13391), .ZN(n13929) );
  AOI22_X1 U14987 ( .A1(n13277), .A2(P2_EAX_REG_10__SCAN_IN), .B1(n13405), 
        .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n13392) );
  OAI21_X1 U14988 ( .B1(n13929), .B2(n13408), .A(n13392), .ZN(n13393) );
  AOI21_X1 U14989 ( .B1(P2_REIP_REG_10__SCAN_IN), .B2(n15456), .A(n13393), 
        .ZN(n16590) );
  AOI22_X1 U14990 ( .A1(n15456), .A2(P2_REIP_REG_11__SCAN_IN), .B1(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n13405), .ZN(n13396) );
  AOI22_X1 U14991 ( .A1(n13394), .A2(n14222), .B1(n13277), .B2(
        P2_EAX_REG_11__SCAN_IN), .ZN(n13395) );
  NAND2_X1 U14992 ( .A1(n13396), .A2(n13395), .ZN(n13862) );
  NAND2_X1 U14993 ( .A1(n13863), .A2(n13862), .ZN(n13861) );
  INV_X1 U14994 ( .A(n13397), .ZN(n14223) );
  AOI22_X1 U14995 ( .A1(n13277), .A2(P2_EAX_REG_12__SCAN_IN), .B1(n13405), 
        .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n13398) );
  OAI21_X1 U14996 ( .B1(n14223), .B2(n13408), .A(n13398), .ZN(n13399) );
  AOI21_X1 U14997 ( .B1(P2_REIP_REG_12__SCAN_IN), .B2(n13323), .A(n13399), 
        .ZN(n14087) );
  NAND2_X1 U14998 ( .A1(n15456), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n13401) );
  AOI22_X1 U14999 ( .A1(n13277), .A2(P2_EAX_REG_13__SCAN_IN), .B1(n13405), 
        .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n13400) );
  OAI211_X1 U15000 ( .C1(n11426), .C2(n13408), .A(n13401), .B(n13400), .ZN(
        n14293) );
  INV_X1 U15001 ( .A(n14494), .ZN(n13404) );
  NAND2_X1 U15002 ( .A1(n13323), .A2(P2_REIP_REG_14__SCAN_IN), .ZN(n13403) );
  AOI22_X1 U15003 ( .A1(n13277), .A2(P2_EAX_REG_14__SCAN_IN), .B1(n13405), 
        .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n13402) );
  OAI211_X1 U15004 ( .C1(n13404), .C2(n13408), .A(n13403), .B(n13402), .ZN(
        n14449) );
  NAND2_X1 U15005 ( .A1(n13323), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n13407) );
  AOI22_X1 U15006 ( .A1(n15461), .A2(P2_EAX_REG_15__SCAN_IN), .B1(n13405), 
        .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n13406) );
  OAI211_X1 U15007 ( .C1(n14795), .C2(n13408), .A(n13407), .B(n13406), .ZN(
        n14789) );
  NAND2_X1 U15008 ( .A1(n15456), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n13411) );
  AOI22_X1 U15009 ( .A1(n15461), .A2(P2_EAX_REG_18__SCAN_IN), .B1(n13405), 
        .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n13410) );
  NAND2_X1 U15010 ( .A1(n15456), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n13413) );
  AOI22_X1 U15011 ( .A1(n15461), .A2(P2_EAX_REG_19__SCAN_IN), .B1(n13405), 
        .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n13412) );
  NAND2_X1 U15012 ( .A1(n15456), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n13415) );
  AOI22_X1 U15013 ( .A1(n15461), .A2(P2_EAX_REG_20__SCAN_IN), .B1(n13405), 
        .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n13414) );
  NAND2_X1 U15014 ( .A1(n13415), .A2(n13414), .ZN(n16476) );
  NAND2_X1 U15015 ( .A1(n15456), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n13417) );
  AOI22_X1 U15016 ( .A1(n15461), .A2(P2_EAX_REG_21__SCAN_IN), .B1(n13405), 
        .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n13416) );
  NAND2_X1 U15017 ( .A1(n13417), .A2(n13416), .ZN(n16227) );
  NAND2_X1 U15018 ( .A1(n15456), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n13419) );
  AOI22_X1 U15019 ( .A1(n15461), .A2(P2_EAX_REG_22__SCAN_IN), .B1(n13405), 
        .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n13418) );
  NAND2_X1 U15020 ( .A1(n15456), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n13421) );
  AOI22_X1 U15021 ( .A1(n15461), .A2(P2_EAX_REG_23__SCAN_IN), .B1(n13405), 
        .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n13420) );
  AND2_X1 U15022 ( .A1(n13421), .A2(n13420), .ZN(n15351) );
  NAND2_X1 U15023 ( .A1(n13323), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n13423) );
  AOI22_X1 U15024 ( .A1(n15461), .A2(P2_EAX_REG_24__SCAN_IN), .B1(n13405), 
        .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n13422) );
  AND2_X1 U15025 ( .A1(n13423), .A2(n13422), .ZN(n15380) );
  NOR2_X2 U15026 ( .A1(n15381), .A2(n15380), .ZN(n15383) );
  INV_X1 U15027 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n18410) );
  AOI22_X1 U15028 ( .A1(n15461), .A2(P2_EAX_REG_25__SCAN_IN), .B1(n13405), 
        .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n13424) );
  OAI21_X1 U15029 ( .B1(n15463), .B2(n18410), .A(n13424), .ZN(n15323) );
  NAND2_X1 U15030 ( .A1(n13323), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n13426) );
  AOI22_X1 U15031 ( .A1(n15461), .A2(P2_EAX_REG_26__SCAN_IN), .B1(n13405), 
        .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n13425) );
  AND2_X1 U15032 ( .A1(n13426), .A2(n13425), .ZN(n16199) );
  NAND2_X1 U15033 ( .A1(n15456), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n13428) );
  AOI22_X1 U15034 ( .A1(n15461), .A2(P2_EAX_REG_27__SCAN_IN), .B1(n13405), 
        .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n13427) );
  AND2_X1 U15035 ( .A1(n13428), .A2(n13427), .ZN(n16186) );
  INV_X1 U15036 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n18454) );
  AOI22_X1 U15037 ( .A1(n15461), .A2(P2_EAX_REG_28__SCAN_IN), .B1(n13405), 
        .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n13429) );
  OAI21_X1 U15038 ( .B1(n15463), .B2(n18454), .A(n13429), .ZN(n16175) );
  AOI22_X1 U15039 ( .A1(n15461), .A2(P2_EAX_REG_29__SCAN_IN), .B1(n13405), 
        .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n13430) );
  OAI21_X1 U15040 ( .B1(n15463), .B2(n18468), .A(n13430), .ZN(n13431) );
  NAND2_X1 U15041 ( .A1(n16176), .A2(n13431), .ZN(n15455) );
  OAI21_X1 U15042 ( .B1(n16176), .B2(n13431), .A(n15455), .ZN(n16412) );
  INV_X1 U15043 ( .A(P2_EAX_REG_29__SCAN_IN), .ZN(n13799) );
  OAI22_X1 U15044 ( .A1(n19658), .A2(n16412), .B1(n13799), .B2(n19401), .ZN(
        n13432) );
  AOI21_X1 U15045 ( .B1(n19653), .B2(n13433), .A(n13432), .ZN(n13436) );
  NAND2_X1 U15046 ( .A1(n19401), .A2(n11021), .ZN(n13434) );
  NOR2_X2 U15047 ( .A1(n13434), .A2(n16678), .ZN(n19654) );
  NOR2_X2 U15048 ( .A1(n13434), .A2(n16679), .ZN(n19655) );
  AOI22_X1 U15049 ( .A1(n19654), .A2(BUF1_REG_29__SCAN_IN), .B1(n19655), .B2(
        BUF2_REG_29__SCAN_IN), .ZN(n13435) );
  AND2_X1 U15050 ( .A1(n13436), .A2(n13435), .ZN(n13437) );
  OAI21_X1 U15051 ( .B1(n16086), .B2(n19659), .A(n13437), .ZN(P2_U2890) );
  NOR2_X1 U15052 ( .A1(P2_BE_N_REG_3__SCAN_IN), .A2(P2_BE_N_REG_2__SCAN_IN), 
        .ZN(n13439) );
  NOR4_X1 U15053 ( .A1(P2_BE_N_REG_1__SCAN_IN), .A2(P2_BE_N_REG_0__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n13438) );
  NAND4_X1 U15054 ( .A1(n13439), .A2(P2_M_IO_N_REG_SCAN_IN), .A3(
        P2_W_R_N_REG_SCAN_IN), .A4(n13438), .ZN(n13442) );
  INV_X1 U15055 ( .A(P1_M_IO_N_REG_SCAN_IN), .ZN(n22220) );
  INV_X1 U15056 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n20102) );
  NOR4_X1 U15057 ( .A1(P1_BE_N_REG_2__SCAN_IN), .A2(P1_BE_N_REG_0__SCAN_IN), 
        .A3(n22220), .A4(n20102), .ZN(n13441) );
  NOR4_X1 U15058 ( .A1(P1_ADS_N_REG_SCAN_IN), .A2(P1_D_C_N_REG_SCAN_IN), .A3(
        P1_BE_N_REG_1__SCAN_IN), .A4(P1_BE_N_REG_3__SCAN_IN), .ZN(n13440) );
  NAND3_X1 U15059 ( .A1(n14301), .A2(n13441), .A3(n13440), .ZN(U214) );
  OR2_X1 U15060 ( .A1(n16226), .A2(n13442), .ZN(n20037) );
  OR2_X1 U15061 ( .A1(n13230), .A2(n18649), .ZN(n13640) );
  NOR2_X1 U15062 ( .A1(n15004), .A2(n13640), .ZN(n18119) );
  INV_X1 U15063 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .ZN(n17091) );
  AND2_X1 U15064 ( .A1(n19316), .A2(n16719), .ZN(n13497) );
  INV_X1 U15065 ( .A(n13497), .ZN(n13446) );
  NAND2_X1 U15066 ( .A1(n13443), .A2(n18099), .ZN(n13444) );
  OAI211_X1 U15067 ( .C1(n18119), .C2(n17091), .A(n13446), .B(n16029), .ZN(
        P2_U2814) );
  NOR2_X1 U15068 ( .A1(n18095), .A2(P2_READREQUEST_REG_SCAN_IN), .ZN(n13447)
         );
  INV_X1 U15069 ( .A(n13247), .ZN(n13445) );
  AOI22_X1 U15070 ( .A1(n13447), .A2(n13446), .B1(n13445), .B2(n18095), .ZN(
        P2_U3612) );
  AOI22_X1 U15071 ( .A1(n16679), .A2(BUF1_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n16678), .ZN(n14793) );
  INV_X1 U15072 ( .A(n19670), .ZN(n13456) );
  OR2_X1 U15073 ( .A1(n13456), .A2(n19667), .ZN(n19116) );
  INV_X1 U15074 ( .A(P2_LWORD_REG_15__SCAN_IN), .ZN(n13450) );
  INV_X1 U15075 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n17129) );
  OAI222_X1 U15076 ( .A1(n19670), .A2(n14793), .B1(n19116), .B2(n13450), .C1(
        n16026), .C2(n17129), .ZN(P2_U2982) );
  AND2_X1 U15077 ( .A1(n12510), .A2(n20029), .ZN(n13451) );
  INV_X1 U15078 ( .A(n21915), .ZN(n21857) );
  AND2_X1 U15079 ( .A1(n21857), .A2(n16772), .ZN(n14504) );
  INV_X1 U15080 ( .A(P1_MEMORYFETCH_REG_SCAN_IN), .ZN(n13452) );
  AOI21_X1 U15081 ( .B1(n13463), .B2(n20029), .A(n13452), .ZN(n13453) );
  OR3_X1 U15082 ( .A1(n14297), .A2(n14504), .A3(n13453), .ZN(P1_U2801) );
  INV_X1 U15083 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n13793) );
  NAND2_X1 U15084 ( .A1(n19668), .A2(P2_UWORD_REG_10__SCAN_IN), .ZN(n13457) );
  INV_X1 U15085 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n20055) );
  OR2_X1 U15086 ( .A1(n16678), .A2(n20055), .ZN(n13455) );
  NAND2_X1 U15087 ( .A1(n16678), .A2(BUF2_REG_10__SCAN_IN), .ZN(n13454) );
  NAND2_X1 U15088 ( .A1(n13455), .A2(n13454), .ZN(n19129) );
  NAND2_X1 U15089 ( .A1(n13456), .A2(n19129), .ZN(n13458) );
  OAI211_X1 U15090 ( .C1(n13793), .C2(n16026), .A(n13457), .B(n13458), .ZN(
        P2_U2962) );
  INV_X1 U15091 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n17117) );
  NAND2_X1 U15092 ( .A1(n19668), .A2(P2_LWORD_REG_10__SCAN_IN), .ZN(n13459) );
  OAI211_X1 U15093 ( .C1(n17117), .C2(n16026), .A(n13459), .B(n13458), .ZN(
        P2_U2977) );
  NOR2_X1 U15094 ( .A1(n14504), .A2(P1_READREQUEST_REG_SCAN_IN), .ZN(n13462)
         );
  OAI21_X1 U15095 ( .B1(n13460), .B2(n15514), .A(n21324), .ZN(n13461) );
  OAI21_X1 U15096 ( .B1(n21324), .B2(n13462), .A(n13461), .ZN(P1_U3487) );
  INV_X1 U15097 ( .A(n12510), .ZN(n13464) );
  INV_X1 U15098 ( .A(n13945), .ZN(n13573) );
  INV_X1 U15099 ( .A(n21718), .ZN(n13727) );
  OAI21_X1 U15100 ( .B1(n13573), .B2(n21319), .A(n13727), .ZN(n13465) );
  NAND2_X1 U15101 ( .A1(n13465), .A2(n21675), .ZN(n21318) );
  NAND2_X1 U15102 ( .A1(n20030), .A2(n21318), .ZN(n16755) );
  AND2_X1 U15103 ( .A1(n16755), .A2(n20029), .ZN(n21657) );
  INV_X1 U15104 ( .A(P1_MORE_REG_SCAN_IN), .ZN(n16948) );
  INV_X1 U15105 ( .A(n13466), .ZN(n13467) );
  NOR2_X1 U15106 ( .A1(n13468), .A2(n13467), .ZN(n13742) );
  OR2_X1 U15107 ( .A1(n13469), .A2(n13905), .ZN(n13470) );
  AND2_X1 U15108 ( .A1(n13742), .A2(n13470), .ZN(n13475) );
  NAND2_X1 U15109 ( .A1(n16006), .A2(n13471), .ZN(n13745) );
  INV_X1 U15110 ( .A(n13745), .ZN(n13472) );
  NAND2_X1 U15111 ( .A1(n13735), .A2(n13472), .ZN(n13474) );
  OR2_X1 U15112 ( .A1(n12511), .A2(n13729), .ZN(n13473) );
  OAI211_X1 U15113 ( .C1(n13735), .C2(n13475), .A(n13474), .B(n13473), .ZN(
        n13476) );
  AND2_X1 U15114 ( .A1(n13476), .A2(n13662), .ZN(n16756) );
  NAND2_X1 U15115 ( .A1(n21657), .A2(n16756), .ZN(n13477) );
  OAI21_X1 U15116 ( .B1(n21657), .B2(n16948), .A(n13477), .ZN(P1_U3484) );
  AND4_X1 U15117 ( .A1(n13480), .A2(n13479), .A3(n13478), .A4(n13500), .ZN(
        n13481) );
  OAI21_X1 U15118 ( .B1(n15004), .B2(n13481), .A(n16719), .ZN(n13485) );
  OR2_X1 U15119 ( .A1(n13482), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n14044) );
  NOR2_X1 U15120 ( .A1(n16719), .A2(P2_FLUSH_REG_SCAN_IN), .ZN(n13483) );
  OAI21_X1 U15121 ( .B1(n13484), .B2(n14044), .A(n13483), .ZN(n17063) );
  NAND2_X1 U15122 ( .A1(n13485), .A2(n17063), .ZN(n18638) );
  NOR2_X1 U15123 ( .A1(n14998), .A2(n13184), .ZN(n15029) );
  INV_X1 U15124 ( .A(n15029), .ZN(n14050) );
  OR2_X1 U15125 ( .A1(n18638), .A2(n14050), .ZN(n13494) );
  AND2_X1 U15126 ( .A1(n13522), .A2(n13486), .ZN(n13487) );
  NOR2_X1 U15127 ( .A1(n13488), .A2(n13487), .ZN(n13490) );
  OR2_X1 U15128 ( .A1(n13490), .A2(n13489), .ZN(n14047) );
  INV_X1 U15129 ( .A(n14047), .ZN(n13493) );
  INV_X1 U15130 ( .A(n13491), .ZN(n13492) );
  NOR2_X1 U15131 ( .A1(n14998), .A2(n13492), .ZN(n15013) );
  NAND2_X1 U15132 ( .A1(n13493), .A2(n15013), .ZN(n15001) );
  NAND2_X1 U15133 ( .A1(n13494), .A2(n15001), .ZN(n14043) );
  NAND2_X1 U15134 ( .A1(n19203), .A2(n17064), .ZN(n18098) );
  NOR2_X1 U15135 ( .A1(n18098), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n13495) );
  NOR2_X1 U15136 ( .A1(n16719), .A2(n21695), .ZN(n16718) );
  INV_X1 U15137 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n18528) );
  NAND2_X1 U15138 ( .A1(n19605), .A2(n13499), .ZN(n13512) );
  INV_X1 U15139 ( .A(n13512), .ZN(n13496) );
  NOR2_X1 U15140 ( .A1(n13496), .A2(n18528), .ZN(n13508) );
  AOI21_X1 U15141 ( .B1(n18528), .B2(n13496), .A(n13508), .ZN(n18515) );
  AND2_X2 U15142 ( .A1(n13497), .A2(n13554), .ZN(n18572) );
  AND2_X1 U15143 ( .A1(n18572), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n18520) );
  MUX2_X1 U15144 ( .A(n13500), .B(n13499), .S(n13498), .Z(n13501) );
  MUX2_X1 U15145 ( .A(n13501), .B(P2_EBX_REG_0__SCAN_IN), .S(n16684), .Z(
        n18106) );
  XNOR2_X1 U15146 ( .A(n18106), .B(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n18517) );
  NOR2_X1 U15147 ( .A1(n17058), .A2(n18517), .ZN(n13502) );
  AOI211_X1 U15148 ( .C1(n17047), .C2(n18515), .A(n18520), .B(n13502), .ZN(
        n13505) );
  NAND2_X1 U15149 ( .A1(n21695), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n13503) );
  NAND2_X1 U15150 ( .A1(n14078), .A2(n13503), .ZN(n13506) );
  OAI21_X1 U15151 ( .B1(n17052), .B2(n13506), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13504) );
  OAI211_X1 U15152 ( .C1(n17062), .C2(n18108), .A(n13505), .B(n13504), .ZN(
        P2_U3014) );
  AOI21_X1 U15153 ( .B1(n18120), .B2(n16041), .A(n14865), .ZN(n16039) );
  XNOR2_X1 U15154 ( .A(n13518), .B(n13507), .ZN(n13509) );
  NAND2_X1 U15155 ( .A1(n13509), .A2(n13508), .ZN(n13510) );
  XOR2_X1 U15156 ( .A(n13509), .B(n13508), .Z(n13538) );
  NAND2_X1 U15157 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n13538), .ZN(
        n13537) );
  NAND2_X1 U15158 ( .A1(n13510), .A2(n13537), .ZN(n14854) );
  XOR2_X1 U15159 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n14854), .Z(
        n13515) );
  OR2_X1 U15160 ( .A1(n13512), .A2(n13511), .ZN(n14850) );
  XOR2_X1 U15161 ( .A(n13513), .B(n14850), .Z(n13514) );
  NAND2_X1 U15162 ( .A1(n13515), .A2(n13514), .ZN(n14856) );
  OAI21_X1 U15163 ( .B1(n13515), .B2(n13514), .A(n14856), .ZN(n18618) );
  AND2_X1 U15164 ( .A1(n18572), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n18611) );
  INV_X1 U15165 ( .A(n18611), .ZN(n13517) );
  OR2_X1 U15166 ( .A1(n17022), .A2(n16041), .ZN(n13516) );
  OAI211_X1 U15167 ( .C1(n17042), .C2(n18618), .A(n13517), .B(n13516), .ZN(
        n13531) );
  NAND2_X1 U15168 ( .A1(n18106), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13521) );
  NOR2_X1 U15169 ( .A1(P2_EBX_REG_0__SCAN_IN), .A2(P2_EBX_REG_1__SCAN_IN), 
        .ZN(n13519) );
  MUX2_X1 U15170 ( .A(n13519), .B(n13518), .S(n15131), .Z(n13525) );
  INV_X1 U15171 ( .A(n13525), .ZN(n13527) );
  NAND3_X1 U15172 ( .A1(n16684), .A2(P2_EBX_REG_1__SCAN_IN), .A3(
        P2_EBX_REG_0__SCAN_IN), .ZN(n13520) );
  NAND2_X1 U15173 ( .A1(n13527), .A2(n13520), .ZN(n18113) );
  NAND2_X1 U15174 ( .A1(n13521), .A2(n18113), .ZN(n13533) );
  INV_X1 U15175 ( .A(n13533), .ZN(n13536) );
  NOR2_X1 U15176 ( .A1(n13521), .A2(n18113), .ZN(n13535) );
  NOR2_X1 U15177 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n13535), .ZN(
        n13534) );
  NOR2_X1 U15178 ( .A1(n13536), .A2(n13534), .ZN(n14863) );
  OAI21_X1 U15179 ( .B1(n14849), .B2(n13184), .A(n13522), .ZN(n13524) );
  INV_X1 U15180 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n13523) );
  MUX2_X1 U15181 ( .A(n13524), .B(n13523), .S(n16684), .Z(n13526) );
  INV_X1 U15182 ( .A(n13526), .ZN(n13528) );
  NAND2_X1 U15183 ( .A1(n13528), .A2(n13527), .ZN(n13529) );
  NAND2_X1 U15184 ( .A1(n11279), .A2(n13529), .ZN(n16040) );
  XNOR2_X1 U15185 ( .A(n16040), .B(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n14862) );
  XNOR2_X1 U15186 ( .A(n14863), .B(n14862), .ZN(n18607) );
  NOR2_X1 U15187 ( .A1(n18607), .A2(n17058), .ZN(n13530) );
  AOI211_X1 U15188 ( .C1(n17055), .C2(n16039), .A(n13531), .B(n13530), .ZN(
        n13532) );
  OAI21_X1 U15189 ( .B1(n14807), .B2(n17062), .A(n13532), .ZN(P2_U3012) );
  AOI222_X1 U15190 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n13536), .B1(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n13535), .C1(n13534), .C2(
        n13533), .ZN(n18525) );
  OAI21_X1 U15191 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n13538), .A(
        n13537), .ZN(n13539) );
  INV_X1 U15192 ( .A(n13539), .ZN(n18530) );
  NAND2_X1 U15193 ( .A1(n17047), .A2(n18530), .ZN(n13540) );
  NAND2_X1 U15194 ( .A1(n18572), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n18535) );
  OAI211_X1 U15195 ( .C1(n17022), .C2(n18120), .A(n13540), .B(n18535), .ZN(
        n13542) );
  NOR2_X1 U15196 ( .A1(n17046), .A2(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13541) );
  AOI211_X1 U15197 ( .C1(n17019), .C2(n18526), .A(n13542), .B(n13541), .ZN(
        n13543) );
  OAI21_X1 U15198 ( .B1(n18525), .B2(n17058), .A(n13543), .ZN(P2_U3013) );
  INV_X1 U15199 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n21745) );
  NAND2_X2 U15200 ( .A1(n21734), .A2(n21745), .ZN(n17138) );
  NOR2_X1 U15201 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(P2_STATE_REG_0__SCAN_IN), 
        .ZN(n21731) );
  NAND2_X1 U15202 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(n21731), .ZN(n17130) );
  NAND2_X1 U15203 ( .A1(n17138), .A2(n17130), .ZN(n21735) );
  NAND2_X1 U15204 ( .A1(n21729), .A2(n21735), .ZN(n14076) );
  OR2_X1 U15205 ( .A1(n13230), .A2(n14076), .ZN(n13553) );
  INV_X1 U15206 ( .A(n14039), .ZN(n13548) );
  INV_X1 U15207 ( .A(n14076), .ZN(n14992) );
  OR2_X1 U15208 ( .A1(n15004), .A2(n13544), .ZN(n13546) );
  AND2_X1 U15209 ( .A1(n13546), .A2(n13545), .ZN(n15002) );
  OAI211_X1 U15210 ( .C1(n13548), .C2(n14040), .A(n13547), .B(n15002), .ZN(
        n13549) );
  INV_X1 U15211 ( .A(n13549), .ZN(n13552) );
  INV_X1 U15212 ( .A(n16640), .ZN(n14052) );
  NAND2_X1 U15213 ( .A1(n13550), .A2(n13551), .ZN(n15044) );
  INV_X1 U15214 ( .A(n15044), .ZN(n14046) );
  NAND2_X1 U15215 ( .A1(n14052), .A2(n14046), .ZN(n13648) );
  OAI211_X1 U15216 ( .C1(n15011), .C2(n13553), .A(n13552), .B(n13648), .ZN(
        n14058) );
  NAND2_X1 U15217 ( .A1(n14058), .A2(n18099), .ZN(n13556) );
  NOR2_X1 U15218 ( .A1(n13554), .A2(n17064), .ZN(n16721) );
  AOI22_X1 U15219 ( .A1(n13554), .A2(P2_STATE2_REG_3__SCAN_IN), .B1(n16721), 
        .B2(P2_FLUSH_REG_SCAN_IN), .ZN(n13555) );
  NAND2_X1 U15220 ( .A1(n13556), .A2(n13555), .ZN(n16652) );
  NOR2_X1 U15221 ( .A1(n13230), .A2(n18090), .ZN(n14045) );
  NAND2_X1 U15222 ( .A1(n16719), .A2(n19203), .ZN(n18628) );
  INV_X1 U15223 ( .A(n18628), .ZN(n16656) );
  NAND2_X1 U15224 ( .A1(n14045), .A2(n16656), .ZN(n13557) );
  NAND2_X1 U15225 ( .A1(n16652), .A2(n13557), .ZN(n13558) );
  OAI211_X1 U15226 ( .C1(n16652), .C2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(
        n13558), .B(n14044), .ZN(n13559) );
  INV_X1 U15227 ( .A(n13559), .ZN(P2_U3595) );
  INV_X1 U15228 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n14347) );
  INV_X1 U15229 ( .A(n16744), .ZN(n13560) );
  NAND2_X1 U15230 ( .A1(n12510), .A2(n14298), .ZN(n16764) );
  NAND2_X1 U15231 ( .A1(n13560), .A2(n16764), .ZN(n13562) );
  NAND2_X1 U15232 ( .A1(n13735), .A2(n21718), .ZN(n16763) );
  NOR2_X1 U15233 ( .A1(n21689), .A2(n16763), .ZN(n13561) );
  NAND2_X1 U15234 ( .A1(n19854), .A2(n13747), .ZN(n13714) );
  NAND2_X1 U15235 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n21667) );
  NOR2_X1 U15236 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n21667), .ZN(n19869) );
  CLKBUF_X2 U15237 ( .A(n19869), .Z(n21325) );
  NOR2_X4 U15238 ( .A1(n19854), .A2(n21325), .ZN(n19866) );
  AOI22_X1 U15239 ( .A1(n19869), .A2(P1_UWORD_REG_7__SCAN_IN), .B1(n19866), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n13563) );
  OAI21_X1 U15240 ( .B1(n14347), .B2(n13714), .A(n13563), .ZN(P1_U2913) );
  INV_X1 U15241 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n15651) );
  AOI22_X1 U15242 ( .A1(n21325), .A2(P1_UWORD_REG_8__SCAN_IN), .B1(n19866), 
        .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n13564) );
  OAI21_X1 U15243 ( .B1(n15651), .B2(n13714), .A(n13564), .ZN(P1_U2912) );
  INV_X1 U15244 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n14394) );
  AOI22_X1 U15245 ( .A1(n21325), .A2(P1_UWORD_REG_5__SCAN_IN), .B1(n19866), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n13565) );
  OAI21_X1 U15246 ( .B1(n14394), .B2(n13714), .A(n13565), .ZN(P1_U2915) );
  AOI22_X1 U15247 ( .A1(n21325), .A2(P1_UWORD_REG_9__SCAN_IN), .B1(n19866), 
        .B2(P1_DATAO_REG_25__SCAN_IN), .ZN(n13566) );
  OAI21_X1 U15248 ( .B1(n15646), .B2(n13714), .A(n13566), .ZN(P1_U2911) );
  AOI22_X1 U15249 ( .A1(n21325), .A2(P1_UWORD_REG_6__SCAN_IN), .B1(n19866), 
        .B2(P1_DATAO_REG_22__SCAN_IN), .ZN(n13567) );
  OAI21_X1 U15250 ( .B1(n15659), .B2(n13714), .A(n13567), .ZN(P1_U2914) );
  OAI22_X1 U15251 ( .A1(n11615), .A2(n13905), .B1(n13568), .B2(n14182), .ZN(
        n13569) );
  INV_X1 U15252 ( .A(n13569), .ZN(n13576) );
  INV_X1 U15253 ( .A(n13570), .ZN(n13572) );
  NAND2_X1 U15254 ( .A1(n13572), .A2(n13571), .ZN(n13574) );
  NAND2_X1 U15255 ( .A1(n13574), .A2(n13573), .ZN(n13575) );
  OAI211_X1 U15256 ( .C1(n13577), .C2(n12613), .A(n13576), .B(n13575), .ZN(
        n13578) );
  INV_X1 U15257 ( .A(n13578), .ZN(n13582) );
  AOI21_X1 U15258 ( .B1(n13579), .B2(n13732), .A(n13905), .ZN(n13580) );
  NAND2_X1 U15259 ( .A1(n13581), .A2(n13580), .ZN(n13599) );
  INV_X1 U15260 ( .A(n13748), .ZN(n13583) );
  NOR2_X1 U15261 ( .A1(n13584), .A2(n13583), .ZN(n13585) );
  NAND3_X1 U15262 ( .A1(n12348), .A2(n13585), .A3(n13725), .ZN(n13586) );
  NOR2_X1 U15263 ( .A1(n13750), .A2(n13586), .ZN(n16739) );
  XNOR2_X1 U15264 ( .A(n13622), .B(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13590) );
  NAND4_X1 U15265 ( .A1(n16006), .A2(n11615), .A3(n14295), .A4(n13945), .ZN(
        n13617) );
  INV_X1 U15266 ( .A(n13617), .ZN(n13589) );
  XNOR2_X1 U15267 ( .A(n13587), .B(n13622), .ZN(n13594) );
  INV_X1 U15268 ( .A(n13594), .ZN(n13588) );
  AOI22_X1 U15269 ( .A1(n16744), .A2(n13590), .B1(n13589), .B2(n13588), .ZN(
        n13592) );
  NAND3_X1 U15270 ( .A1(n16739), .A2(n11613), .A3(n13594), .ZN(n13591) );
  OAI211_X1 U15271 ( .C1(n21860), .C2(n16739), .A(n13592), .B(n13591), .ZN(
        n13981) );
  INV_X1 U15272 ( .A(n21666), .ZN(n16703) );
  INV_X1 U15273 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n21658) );
  NOR2_X1 U15274 ( .A1(n16772), .A2(n21658), .ZN(n16013) );
  AOI22_X1 U15275 ( .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n15821), .B1(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n12527), .ZN(n16014) );
  INV_X1 U15276 ( .A(n16014), .ZN(n13595) );
  AOI222_X1 U15277 ( .A1(n13981), .A2(n16703), .B1(n16013), .B2(n13595), .C1(
        n21683), .C2(n13594), .ZN(n13612) );
  INV_X1 U15278 ( .A(n16763), .ZN(n13596) );
  OAI211_X1 U15279 ( .C1(n16744), .C2(n13597), .A(n13596), .B(n21675), .ZN(
        n13602) );
  INV_X1 U15280 ( .A(n13598), .ZN(n13600) );
  NAND2_X1 U15281 ( .A1(n13600), .A2(n13599), .ZN(n13601) );
  NAND2_X1 U15282 ( .A1(n13601), .A2(n12511), .ZN(n13733) );
  OAI211_X1 U15283 ( .C1(n13945), .C2(n11617), .A(n13602), .B(n13733), .ZN(
        n13603) );
  INV_X1 U15284 ( .A(n13603), .ZN(n13604) );
  OAI21_X1 U15285 ( .B1(n13735), .B2(n13745), .A(n13604), .ZN(n13605) );
  OR2_X1 U15286 ( .A1(n13606), .A2(n13605), .ZN(n13983) );
  NAND2_X1 U15287 ( .A1(n13983), .A2(n20029), .ZN(n13610) );
  INV_X1 U15288 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n21656) );
  INV_X1 U15289 ( .A(n21667), .ZN(n13902) );
  NAND2_X1 U15290 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n13902), .ZN(n21680) );
  NOR2_X1 U15291 ( .A1(n21656), .A2(n21680), .ZN(n13608) );
  NOR2_X1 U15292 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n21868), .ZN(n13607) );
  NOR2_X1 U15293 ( .A1(n13608), .A2(n13607), .ZN(n13609) );
  NAND2_X1 U15294 ( .A1(n13610), .A2(n13609), .ZN(n21661) );
  NAND2_X1 U15295 ( .A1(n21663), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13611) );
  OAI21_X1 U15296 ( .B1(n13612), .B2(n21663), .A(n13611), .ZN(P1_U3472) );
  INV_X1 U15297 ( .A(n21769), .ZN(n13628) );
  XNOR2_X1 U15298 ( .A(n13613), .B(n11492), .ZN(n13621) );
  INV_X1 U15299 ( .A(n13614), .ZN(n13619) );
  INV_X1 U15300 ( .A(n13615), .ZN(n13616) );
  MUX2_X1 U15301 ( .A(n13616), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n13587), .Z(n13618) );
  AOI21_X1 U15302 ( .B1(n13619), .B2(n13618), .A(n13617), .ZN(n13620) );
  AOI21_X1 U15303 ( .B1(n16744), .B2(n13621), .A(n13620), .ZN(n13627) );
  INV_X1 U15304 ( .A(n13587), .ZN(n13623) );
  OAI21_X1 U15305 ( .B1(n13623), .B2(n13622), .A(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13624) );
  NAND2_X1 U15306 ( .A1(n13625), .A2(n13624), .ZN(n13629) );
  NAND3_X1 U15307 ( .A1(n16739), .A2(n11613), .A3(n13629), .ZN(n13626) );
  OAI211_X1 U15308 ( .C1(n13628), .C2(n16739), .A(n13627), .B(n13626), .ZN(
        n13982) );
  AOI22_X1 U15309 ( .A1(n13982), .A2(n16703), .B1(n21683), .B2(n13629), .ZN(
        n13631) );
  NAND2_X1 U15310 ( .A1(n21663), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13630) );
  OAI21_X1 U15311 ( .B1(n13631), .B2(n21663), .A(n13630), .ZN(P1_U3469) );
  OR2_X1 U15312 ( .A1(n14376), .A2(BUF1_REG_0__SCAN_IN), .ZN(n13633) );
  INV_X1 U15313 ( .A(DATAI_0_), .ZN(n16927) );
  NAND2_X1 U15314 ( .A1(n14376), .A2(n16927), .ZN(n13632) );
  NAND2_X1 U15315 ( .A1(n13633), .A2(n13632), .ZN(n15690) );
  NAND2_X1 U15316 ( .A1(n13634), .A2(n13662), .ZN(n13635) );
  INV_X1 U15317 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n19856) );
  NAND2_X2 U15318 ( .A1(n15703), .A2(n13635), .ZN(n15711) );
  NAND2_X1 U15319 ( .A1(n13637), .A2(n13636), .ZN(n13638) );
  NAND2_X1 U15320 ( .A1(n13639), .A2(n13638), .ZN(n19977) );
  OAI222_X1 U15321 ( .A1(n15690), .A2(n15701), .B1(n15703), .B2(n19856), .C1(
        n15711), .C2(n19977), .ZN(P1_U2904) );
  INV_X1 U15322 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n13643) );
  OAI21_X1 U15323 ( .B1(n15011), .B2(n13640), .A(n16026), .ZN(n13641) );
  NOR2_X1 U15324 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n17064), .ZN(n17115) );
  NOR2_X4 U15325 ( .A1(n17095), .A2(n17126), .ZN(n17114) );
  AOI22_X1 U15326 ( .A1(n17115), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n17114), 
        .B2(P2_DATAO_REG_18__SCAN_IN), .ZN(n13642) );
  OAI21_X1 U15327 ( .B1(n13643), .B2(n13808), .A(n13642), .ZN(P2_U2933) );
  INV_X1 U15328 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n15059) );
  AOI22_X1 U15329 ( .A1(n17115), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n17114), 
        .B2(P2_DATAO_REG_17__SCAN_IN), .ZN(n13644) );
  OAI21_X1 U15330 ( .B1(n15059), .B2(n13808), .A(n13644), .ZN(P2_U2934) );
  INV_X1 U15331 ( .A(n13647), .ZN(n15031) );
  NAND2_X1 U15332 ( .A1(n13648), .A2(n15031), .ZN(n13649) );
  INV_X2 U15333 ( .A(n16102), .ZN(n16111) );
  MUX2_X1 U15334 ( .A(n14808), .B(n12777), .S(n16111), .Z(n13650) );
  OAI21_X1 U15335 ( .B1(n19152), .B2(n16167), .A(n13650), .ZN(P2_U2886) );
  NAND2_X1 U15336 ( .A1(n18090), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n13651) );
  AND4_X1 U15337 ( .A1(n13651), .A2(n12828), .A3(P2_STATE2_REG_0__SCAN_IN), 
        .A4(n19203), .ZN(n13652) );
  MUX2_X1 U15338 ( .A(n18108), .B(n18103), .S(n16111), .Z(n13653) );
  OAI21_X1 U15339 ( .B1(n19147), .B2(n16167), .A(n13653), .ZN(P2_U2887) );
  INV_X1 U15340 ( .A(n13654), .ZN(n13655) );
  XNOR2_X1 U15341 ( .A(n13656), .B(n13655), .ZN(n21428) );
  INV_X1 U15342 ( .A(n21428), .ZN(n13717) );
  OR2_X1 U15343 ( .A1(n13745), .A2(n21689), .ZN(n13661) );
  INV_X1 U15344 ( .A(n13657), .ZN(n13659) );
  NAND3_X1 U15345 ( .A1(n13659), .A2(n13663), .A3(n13658), .ZN(n13660) );
  XNOR2_X1 U15346 ( .A(n21424), .B(n13663), .ZN(n13754) );
  AOI22_X1 U15347 ( .A1(n19961), .A2(n13754), .B1(n15617), .B2(
        P1_EBX_REG_1__SCAN_IN), .ZN(n13664) );
  OAI21_X1 U15348 ( .B1(n13717), .B2(n19966), .A(n13664), .ZN(P1_U2871) );
  MUX2_X1 U15349 ( .A(n14807), .B(n13523), .S(n16111), .Z(n13667) );
  OAI21_X1 U15350 ( .B1(n19219), .B2(n16167), .A(n13667), .ZN(P2_U2885) );
  INV_X1 U15351 ( .A(n19403), .ZN(n19130) );
  INV_X1 U15352 ( .A(BUF1_REG_0__SCAN_IN), .ZN(n20039) );
  INV_X1 U15353 ( .A(BUF2_REG_0__SCAN_IN), .ZN(n20135) );
  AOI22_X1 U15354 ( .A1(n16679), .A2(n20039), .B1(n20135), .B2(n16226), .ZN(
        n19665) );
  INV_X1 U15355 ( .A(n13668), .ZN(n13674) );
  INV_X1 U15356 ( .A(n13669), .ZN(n13672) );
  INV_X1 U15357 ( .A(n13670), .ZN(n13671) );
  NAND2_X1 U15358 ( .A1(n13672), .A2(n13671), .ZN(n13673) );
  NAND2_X1 U15359 ( .A1(n13674), .A2(n13673), .ZN(n18518) );
  OAI22_X1 U15360 ( .A1(n19658), .A2(n18518), .B1(n19401), .B2(n13675), .ZN(
        n13677) );
  NOR2_X1 U15361 ( .A1(n19147), .A2(n18518), .ZN(n13691) );
  AOI211_X1 U15362 ( .C1(n19147), .C2(n18518), .A(n19659), .B(n13691), .ZN(
        n13676) );
  AOI211_X1 U15363 ( .C1(n19130), .C2(n19665), .A(n13677), .B(n13676), .ZN(
        n13678) );
  INV_X1 U15364 ( .A(n13678), .ZN(P2_U2919) );
  OAI21_X1 U15365 ( .B1(n13680), .B2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n13679), .ZN(n21407) );
  OAI222_X1 U15366 ( .A1(n21407), .A2(n19965), .B1(n19969), .B2(n14081), .C1(
        n19977), .C2(n19966), .ZN(P1_U2872) );
  INV_X1 U15367 ( .A(BUF1_REG_6__SCAN_IN), .ZN(n20048) );
  INV_X1 U15368 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n20145) );
  AOI22_X1 U15369 ( .A1(n16679), .A2(n20048), .B1(n20145), .B2(n16226), .ZN(
        n19349) );
  INV_X1 U15370 ( .A(n19349), .ZN(n19358) );
  XNOR2_X1 U15371 ( .A(n13682), .B(n13681), .ZN(n18162) );
  INV_X1 U15372 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n17107) );
  OAI222_X1 U15373 ( .A1(n19403), .A2(n19358), .B1(n18162), .B2(n19410), .C1(
        n19401), .C2(n17107), .ZN(P2_U2913) );
  AOI22_X1 U15374 ( .A1(n16679), .A2(BUF1_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n16678), .ZN(n19146) );
  OAI21_X1 U15375 ( .B1(n13685), .B2(n13684), .A(n13683), .ZN(n18176) );
  OAI222_X1 U15376 ( .A1(n19403), .A2(n19146), .B1(n18176), .B2(n19410), .C1(
        n19401), .C2(n17109), .ZN(P2_U2912) );
  AOI22_X1 U15377 ( .A1(n16679), .A2(BUF1_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n16226), .ZN(n19138) );
  AOI21_X1 U15378 ( .B1(n13686), .B2(n13683), .A(n13723), .ZN(n18566) );
  INV_X1 U15379 ( .A(n18566), .ZN(n13687) );
  INV_X1 U15380 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n17111) );
  OAI222_X1 U15381 ( .A1(n19403), .A2(n19138), .B1(n13687), .B2(n19410), .C1(
        n19401), .C2(n17111), .ZN(P2_U2911) );
  XNOR2_X1 U15382 ( .A(n13689), .B(n13688), .ZN(n18116) );
  NAND2_X1 U15383 ( .A1(n19152), .A2(n18116), .ZN(n13866) );
  OAI21_X1 U15384 ( .B1(n19152), .B2(n18116), .A(n13866), .ZN(n13690) );
  NOR2_X1 U15385 ( .A1(n13690), .A2(n13691), .ZN(n13868) );
  AOI21_X1 U15386 ( .B1(n13691), .B2(n13690), .A(n13868), .ZN(n13694) );
  INV_X1 U15387 ( .A(n18116), .ZN(n18527) );
  AOI22_X1 U15388 ( .A1(n19548), .A2(n18527), .B1(n19652), .B2(
        P2_EAX_REG_1__SCAN_IN), .ZN(n13693) );
  AOI22_X1 U15389 ( .A1(n16679), .A2(BUF1_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n16226), .ZN(n19604) );
  INV_X1 U15390 ( .A(n19604), .ZN(n15062) );
  NAND2_X1 U15391 ( .A1(n19130), .A2(n15062), .ZN(n13692) );
  OAI211_X1 U15392 ( .C1(n13694), .C2(n19659), .A(n13693), .B(n13692), .ZN(
        P2_U2918) );
  XNOR2_X1 U15393 ( .A(n13695), .B(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13759) );
  AOI22_X1 U15394 ( .A1(n20022), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B1(
        n10970), .B2(P1_REIP_REG_1__SCAN_IN), .ZN(n13696) );
  OAI21_X1 U15395 ( .B1(n20028), .B2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n13696), .ZN(n13697) );
  AOI21_X1 U15396 ( .B1(n21428), .B2(n20009), .A(n13697), .ZN(n13698) );
  OAI21_X1 U15397 ( .B1(n13759), .B2(n21655), .A(n13698), .ZN(P1_U2998) );
  AOI22_X1 U15398 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n19866), .B1(n19869), 
        .B2(P1_UWORD_REG_0__SCAN_IN), .ZN(n13699) );
  OAI21_X1 U15399 ( .B1(n15688), .B2(n13714), .A(n13699), .ZN(P1_U2920) );
  INV_X1 U15400 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n14360) );
  AOI22_X1 U15401 ( .A1(n19869), .A2(P1_UWORD_REG_1__SCAN_IN), .B1(n19866), 
        .B2(P1_DATAO_REG_17__SCAN_IN), .ZN(n13700) );
  OAI21_X1 U15402 ( .B1(n14360), .B2(n13714), .A(n13700), .ZN(P1_U2919) );
  INV_X1 U15403 ( .A(P2_EBX_REG_3__SCAN_IN), .ZN(n16034) );
  MUX2_X1 U15404 ( .A(n14816), .B(n16034), .S(n16111), .Z(n13705) );
  OAI21_X1 U15405 ( .B1(n19328), .B2(n16167), .A(n13705), .ZN(P2_U2884) );
  INV_X1 U15406 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n14375) );
  AOI22_X1 U15407 ( .A1(n21325), .A2(P1_UWORD_REG_13__SCAN_IN), .B1(n19866), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n13706) );
  OAI21_X1 U15408 ( .B1(n14375), .B2(n13714), .A(n13706), .ZN(P1_U2907) );
  INV_X1 U15409 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n14339) );
  AOI22_X1 U15410 ( .A1(n21325), .A2(P1_UWORD_REG_10__SCAN_IN), .B1(n19866), 
        .B2(P1_DATAO_REG_26__SCAN_IN), .ZN(n13707) );
  OAI21_X1 U15411 ( .B1(n14339), .B2(n13714), .A(n13707), .ZN(P1_U2910) );
  INV_X1 U15412 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n14331) );
  AOI22_X1 U15413 ( .A1(n21325), .A2(P1_UWORD_REG_12__SCAN_IN), .B1(n19866), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n13708) );
  OAI21_X1 U15414 ( .B1(n14331), .B2(n13714), .A(n13708), .ZN(P1_U2908) );
  INV_X1 U15415 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n14386) );
  AOI22_X1 U15416 ( .A1(n21325), .A2(P1_UWORD_REG_14__SCAN_IN), .B1(n19866), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .ZN(n13709) );
  OAI21_X1 U15417 ( .B1(n14386), .B2(n13714), .A(n13709), .ZN(P1_U2906) );
  INV_X1 U15418 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n14355) );
  AOI22_X1 U15419 ( .A1(n21325), .A2(P1_UWORD_REG_3__SCAN_IN), .B1(n19866), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n13710) );
  OAI21_X1 U15420 ( .B1(n14355), .B2(n13714), .A(n13710), .ZN(P1_U2917) );
  AOI22_X1 U15421 ( .A1(n21325), .A2(P1_UWORD_REG_2__SCAN_IN), .B1(n19866), 
        .B2(P1_DATAO_REG_18__SCAN_IN), .ZN(n13711) );
  OAI21_X1 U15422 ( .B1(n15675), .B2(n13714), .A(n13711), .ZN(P1_U2918) );
  INV_X1 U15423 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n14383) );
  AOI22_X1 U15424 ( .A1(n21325), .A2(P1_UWORD_REG_11__SCAN_IN), .B1(n19866), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n13712) );
  OAI21_X1 U15425 ( .B1(n14383), .B2(n13714), .A(n13712), .ZN(P1_U2909) );
  AOI22_X1 U15426 ( .A1(n21325), .A2(P1_UWORD_REG_4__SCAN_IN), .B1(n19866), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n13713) );
  OAI21_X1 U15427 ( .B1(n15667), .B2(n13714), .A(n13713), .ZN(P1_U2916) );
  OR2_X1 U15428 ( .A1(n14376), .A2(BUF1_REG_1__SCAN_IN), .ZN(n13716) );
  INV_X1 U15429 ( .A(DATAI_1_), .ZN(n16926) );
  NAND2_X1 U15430 ( .A1(n14376), .A2(n16926), .ZN(n13715) );
  NAND2_X1 U15431 ( .A1(n13716), .A2(n13715), .ZN(n14344) );
  INV_X1 U15432 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n19858) );
  OAI222_X1 U15433 ( .A1(n14344), .A2(n15701), .B1(n15703), .B2(n19858), .C1(
        n15711), .C2(n13717), .ZN(P1_U2903) );
  INV_X1 U15434 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n13718) );
  OR2_X1 U15435 ( .A1(n16678), .A2(n13718), .ZN(n13720) );
  NAND2_X1 U15436 ( .A1(n16678), .A2(BUF2_REG_9__SCAN_IN), .ZN(n13719) );
  AND2_X1 U15437 ( .A1(n13720), .A2(n13719), .ZN(n19135) );
  INV_X1 U15438 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n17113) );
  OAI21_X1 U15439 ( .B1(n13723), .B2(n13722), .A(n13721), .ZN(n18201) );
  OAI222_X1 U15440 ( .A1(n19403), .A2(n19135), .B1(n19401), .B2(n17113), .C1(
        n19410), .C2(n18201), .ZN(P2_U2910) );
  OAI211_X1 U15441 ( .C1(n13725), .C2(n13724), .A(n13747), .B(n11614), .ZN(
        n13726) );
  NAND2_X1 U15442 ( .A1(n13735), .A2(n13726), .ZN(n13731) );
  AOI21_X1 U15443 ( .B1(n13732), .B2(n13727), .A(n21712), .ZN(n13728) );
  NAND2_X1 U15444 ( .A1(n13729), .A2(n13728), .ZN(n13730) );
  MUX2_X1 U15445 ( .A(n13731), .B(n13730), .S(n11617), .Z(n13738) );
  NAND2_X1 U15446 ( .A1(n16006), .A2(n13732), .ZN(n13734) );
  OAI21_X1 U15447 ( .B1(n13735), .B2(n13734), .A(n13733), .ZN(n13736) );
  INV_X1 U15448 ( .A(n13736), .ZN(n13737) );
  OR2_X1 U15449 ( .A1(n13739), .A2(n14173), .ZN(n13740) );
  NAND4_X1 U15450 ( .A1(n13742), .A2(n12348), .A3(n13741), .A4(n13740), .ZN(
        n13743) );
  INV_X1 U15451 ( .A(n13753), .ZN(n13744) );
  INV_X1 U15452 ( .A(n15987), .ZN(n21413) );
  OAI21_X1 U15453 ( .B1(n13748), .B2(n13747), .A(n13746), .ZN(n13749) );
  OR2_X1 U15454 ( .A1(n13750), .A2(n13749), .ZN(n13751) );
  OAI22_X1 U15455 ( .A1(n10970), .A2(n13753), .B1(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n21412), .ZN(n15903) );
  OAI21_X1 U15456 ( .B1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n21413), .A(
        n15982), .ZN(n21415) );
  INV_X1 U15457 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n19947) );
  NOR2_X1 U15458 ( .A1(n15987), .A2(n15938), .ZN(n21351) );
  INV_X1 U15459 ( .A(n21351), .ZN(n15820) );
  NAND2_X1 U15460 ( .A1(n21658), .A2(n15967), .ZN(n13764) );
  NAND3_X1 U15461 ( .A1(n12527), .A2(n15820), .A3(n13764), .ZN(n13756) );
  OAI21_X1 U15462 ( .B1(n13739), .B2(n11640), .A(n16764), .ZN(n13752) );
  NAND2_X1 U15463 ( .A1(n21409), .A2(n13754), .ZN(n13755) );
  OAI211_X1 U15464 ( .C1(n19947), .C2(n21386), .A(n13756), .B(n13755), .ZN(
        n13757) );
  AOI21_X1 U15465 ( .B1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n21415), .A(
        n13757), .ZN(n13758) );
  OAI21_X1 U15466 ( .B1(n13759), .B2(n21353), .A(n13758), .ZN(P1_U3030) );
  XNOR2_X1 U15467 ( .A(n13761), .B(n13760), .ZN(n13763) );
  XNOR2_X1 U15468 ( .A(n13763), .B(n13762), .ZN(n13783) );
  NAND2_X1 U15469 ( .A1(n15938), .A2(n13764), .ZN(n15823) );
  OR3_X1 U15470 ( .A1(n12527), .A2(n15823), .A3(
        P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n13774) );
  INV_X1 U15471 ( .A(n15938), .ZN(n15984) );
  NAND2_X1 U15472 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n13765) );
  OAI22_X1 U15473 ( .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n15984), .B1(
        n13765), .B2(n21413), .ZN(n13766) );
  OR2_X1 U15474 ( .A1(n13766), .A2(n15903), .ZN(n13772) );
  NOR2_X1 U15475 ( .A1(n13768), .A2(n13767), .ZN(n13769) );
  OR2_X1 U15476 ( .A1(n13875), .A2(n13769), .ZN(n13946) );
  AOI21_X1 U15477 ( .B1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n14879) );
  NAND2_X1 U15478 ( .A1(n15987), .A2(n14879), .ZN(n13770) );
  NAND2_X1 U15479 ( .A1(n10970), .A2(P1_REIP_REG_2__SCAN_IN), .ZN(n13780) );
  OAI211_X1 U15480 ( .C1(n21352), .C2(n13946), .A(n13770), .B(n13780), .ZN(
        n13771) );
  AOI21_X1 U15481 ( .B1(n13772), .B2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A(
        n13771), .ZN(n13773) );
  OAI211_X1 U15482 ( .C1(n13783), .C2(n21353), .A(n13774), .B(n13773), .ZN(
        P1_U3029) );
  INV_X1 U15483 ( .A(n13775), .ZN(n13776) );
  AOI21_X1 U15484 ( .B1(n13778), .B2(n13777), .A(n13776), .ZN(n13784) );
  NAND2_X1 U15485 ( .A1(n20022), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13779) );
  OAI211_X1 U15486 ( .C1(n20028), .C2(n13954), .A(n13780), .B(n13779), .ZN(
        n13781) );
  AOI21_X1 U15487 ( .B1(n13784), .B2(n20009), .A(n13781), .ZN(n13782) );
  OAI21_X1 U15488 ( .B1(n21655), .B2(n13783), .A(n13782), .ZN(P1_U2997) );
  INV_X1 U15489 ( .A(n13784), .ZN(n13958) );
  INV_X1 U15490 ( .A(n13946), .ZN(n13785) );
  AOI22_X1 U15491 ( .A1(n19961), .A2(n13785), .B1(n15617), .B2(
        P1_EBX_REG_2__SCAN_IN), .ZN(n13786) );
  OAI21_X1 U15492 ( .B1(n13958), .B2(n19966), .A(n13786), .ZN(P1_U2870) );
  INV_X1 U15493 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n13788) );
  AOI22_X1 U15494 ( .A1(P2_DATAO_REG_16__SCAN_IN), .A2(n17114), .B1(n17126), 
        .B2(P2_UWORD_REG_0__SCAN_IN), .ZN(n13787) );
  OAI21_X1 U15495 ( .B1(n13788), .B2(n13808), .A(n13787), .ZN(P2_U2935) );
  INV_X1 U15496 ( .A(BUF1_REG_2__SCAN_IN), .ZN(n13789) );
  OR2_X1 U15497 ( .A1(n14376), .A2(n13789), .ZN(n13791) );
  NAND2_X1 U15498 ( .A1(n14376), .A2(DATAI_2_), .ZN(n13790) );
  AND2_X1 U15499 ( .A1(n13791), .A2(n13790), .ZN(n15677) );
  INV_X1 U15500 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n19860) );
  OAI222_X1 U15501 ( .A1(n13958), .A2(n15711), .B1(n15701), .B2(n15677), .C1(
        n15703), .C2(n19860), .ZN(P1_U2902) );
  AOI22_X1 U15502 ( .A1(n17126), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(n17114), 
        .B2(P2_DATAO_REG_26__SCAN_IN), .ZN(n13792) );
  OAI21_X1 U15503 ( .B1(n13793), .B2(n13808), .A(n13792), .ZN(P2_U2925) );
  INV_X1 U15504 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n13795) );
  AOI22_X1 U15505 ( .A1(n17126), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n17114), 
        .B2(P2_DATAO_REG_20__SCAN_IN), .ZN(n13794) );
  OAI21_X1 U15506 ( .B1(n13795), .B2(n13808), .A(n13794), .ZN(P2_U2931) );
  INV_X1 U15507 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n16179) );
  AOI22_X1 U15508 ( .A1(n17126), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(n17114), 
        .B2(P2_DATAO_REG_28__SCAN_IN), .ZN(n13796) );
  OAI21_X1 U15509 ( .B1(n16179), .B2(n13808), .A(n13796), .ZN(P2_U2923) );
  INV_X1 U15510 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n16210) );
  AOI22_X1 U15511 ( .A1(n17126), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(n17114), 
        .B2(P2_DATAO_REG_24__SCAN_IN), .ZN(n13797) );
  OAI21_X1 U15512 ( .B1(n16210), .B2(n13808), .A(n13797), .ZN(P2_U2927) );
  AOI22_X1 U15513 ( .A1(n17126), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(n17114), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n13798) );
  OAI21_X1 U15514 ( .B1(n13799), .B2(n13808), .A(n13798), .ZN(P2_U2922) );
  INV_X1 U15515 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n16204) );
  AOI22_X1 U15516 ( .A1(n17126), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(n17114), 
        .B2(P2_DATAO_REG_25__SCAN_IN), .ZN(n13800) );
  OAI21_X1 U15517 ( .B1(n16204), .B2(n13808), .A(n13800), .ZN(P2_U2926) );
  INV_X1 U15518 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n16230) );
  AOI22_X1 U15519 ( .A1(n17126), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n17114), 
        .B2(P2_DATAO_REG_21__SCAN_IN), .ZN(n13801) );
  OAI21_X1 U15520 ( .B1(n16230), .B2(n13808), .A(n13801), .ZN(P2_U2930) );
  INV_X1 U15521 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n16218) );
  AOI22_X1 U15522 ( .A1(n17126), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n17114), 
        .B2(P2_DATAO_REG_23__SCAN_IN), .ZN(n13802) );
  OAI21_X1 U15523 ( .B1(n16218), .B2(n13808), .A(n13802), .ZN(P2_U2928) );
  INV_X1 U15524 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n13804) );
  AOI22_X1 U15525 ( .A1(n17126), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(n17114), 
        .B2(P2_DATAO_REG_22__SCAN_IN), .ZN(n13803) );
  OAI21_X1 U15526 ( .B1(n13804), .B2(n13808), .A(n13803), .ZN(P2_U2929) );
  INV_X1 U15527 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n16189) );
  AOI22_X1 U15528 ( .A1(n17126), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(n17114), 
        .B2(P2_DATAO_REG_27__SCAN_IN), .ZN(n13805) );
  OAI21_X1 U15529 ( .B1(n16189), .B2(n13808), .A(n13805), .ZN(P2_U2924) );
  INV_X1 U15530 ( .A(P2_EAX_REG_30__SCAN_IN), .ZN(n16168) );
  AOI22_X1 U15531 ( .A1(n17115), .A2(P2_UWORD_REG_14__SCAN_IN), .B1(n17114), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .ZN(n13806) );
  OAI21_X1 U15532 ( .B1(n16168), .B2(n13808), .A(n13806), .ZN(P2_U2921) );
  INV_X1 U15533 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n16240) );
  AOI22_X1 U15534 ( .A1(n17115), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n17114), 
        .B2(P2_DATAO_REG_19__SCAN_IN), .ZN(n13807) );
  OAI21_X1 U15535 ( .B1(n16240), .B2(n13808), .A(n13807), .ZN(P2_U2932) );
  INV_X1 U15536 ( .A(n13822), .ZN(n13924) );
  NAND2_X1 U15537 ( .A1(n13924), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13814) );
  INV_X1 U15538 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n13811) );
  NAND2_X1 U15539 ( .A1(n15227), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n13810) );
  NAND2_X1 U15540 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n13809) );
  OAI211_X1 U15541 ( .C1(n15436), .C2(n13811), .A(n13810), .B(n13809), .ZN(
        n13812) );
  INV_X1 U15542 ( .A(n13812), .ZN(n13813) );
  NAND2_X1 U15543 ( .A1(n13814), .A2(n13813), .ZN(n13838) );
  INV_X1 U15544 ( .A(n13816), .ZN(n13817) );
  NAND2_X1 U15545 ( .A1(n13815), .A2(n13817), .ZN(n13821) );
  OR2_X1 U15546 ( .A1(n13819), .A2(n13818), .ZN(n13820) );
  NAND2_X1 U15547 ( .A1(n13821), .A2(n13820), .ZN(n13888) );
  INV_X1 U15548 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n13825) );
  NAND2_X1 U15549 ( .A1(n15227), .A2(P2_EBX_REG_4__SCAN_IN), .ZN(n13824) );
  NAND2_X1 U15550 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n13823) );
  OAI211_X1 U15551 ( .C1(n15436), .C2(n13825), .A(n13824), .B(n13823), .ZN(
        n13826) );
  AOI21_X1 U15552 ( .B1(n13924), .B2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A(
        n13826), .ZN(n13887) );
  INV_X1 U15553 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n13830) );
  NAND2_X1 U15554 ( .A1(n15227), .A2(P2_EBX_REG_5__SCAN_IN), .ZN(n13829) );
  NAND2_X1 U15555 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n13828) );
  OAI211_X1 U15556 ( .C1(n15436), .C2(n13830), .A(n13829), .B(n13828), .ZN(
        n13831) );
  AOI21_X1 U15557 ( .B1(n13924), .B2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A(
        n13831), .ZN(n13846) );
  INV_X1 U15558 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n13834) );
  NAND2_X1 U15559 ( .A1(n13924), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13833) );
  AOI22_X1 U15560 ( .A1(n15227), .A2(P2_EBX_REG_6__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13832) );
  OAI211_X1 U15561 ( .C1(n15436), .C2(n13834), .A(n13833), .B(n13832), .ZN(
        n13879) );
  NAND2_X1 U15562 ( .A1(n15227), .A2(P2_EBX_REG_7__SCAN_IN), .ZN(n13836) );
  NAND2_X1 U15563 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n13835) );
  OAI211_X1 U15564 ( .C1(n10963), .C2(n17133), .A(n13836), .B(n13835), .ZN(
        n13837) );
  AOI21_X1 U15565 ( .B1(n13924), .B2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n13837), .ZN(n13960) );
  OAI21_X1 U15566 ( .B1(n13838), .B2(n13961), .A(n13857), .ZN(n18192) );
  AND2_X1 U15567 ( .A1(n13839), .A2(n13891), .ZN(n13841) );
  AND2_X1 U15568 ( .A1(n13841), .A2(n13840), .ZN(n13843) );
  OAI211_X1 U15569 ( .C1(n13843), .C2(n13842), .A(n13931), .B(n16141), .ZN(
        n13845) );
  NAND2_X1 U15570 ( .A1(n16111), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n13844) );
  OAI211_X1 U15571 ( .C1(n18192), .C2(n16157), .A(n13845), .B(n13844), .ZN(
        P2_U2879) );
  NAND2_X1 U15572 ( .A1(n13839), .A2(n13891), .ZN(n13893) );
  XOR2_X1 U15573 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B(n13893), .Z(n13850)
         );
  AND2_X1 U15574 ( .A1(n13890), .A2(n13846), .ZN(n13847) );
  OR2_X1 U15575 ( .A1(n13847), .A2(n13880), .ZN(n18149) );
  INV_X1 U15576 ( .A(P2_EBX_REG_5__SCAN_IN), .ZN(n13848) );
  MUX2_X1 U15577 ( .A(n18149), .B(n13848), .S(n16111), .Z(n13849) );
  OAI21_X1 U15578 ( .B1(n13850), .B2(n16167), .A(n13849), .ZN(P2_U2882) );
  XOR2_X1 U15579 ( .A(n13928), .B(n13931), .Z(n13860) );
  INV_X1 U15580 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n13853) );
  NAND2_X1 U15581 ( .A1(n15227), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n13852) );
  NAND2_X1 U15582 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n13851) );
  OAI211_X1 U15583 ( .C1(n15436), .C2(n13853), .A(n13852), .B(n13851), .ZN(
        n13854) );
  AOI21_X1 U15584 ( .B1(n13924), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n13854), .ZN(n13856) );
  NAND2_X1 U15585 ( .A1(n13857), .A2(n13856), .ZN(n13858) );
  AND2_X1 U15586 ( .A1(n13926), .A2(n13858), .ZN(n17004) );
  INV_X1 U15587 ( .A(n17004), .ZN(n18202) );
  INV_X1 U15588 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n18197) );
  MUX2_X1 U15589 ( .A(n18202), .B(n18197), .S(n16111), .Z(n13859) );
  OAI21_X1 U15590 ( .B1(n13860), .B2(n16167), .A(n13859), .ZN(P2_U2878) );
  AOI22_X1 U15591 ( .A1(n16679), .A2(BUF1_REG_11__SCAN_IN), .B1(
        BUF2_REG_11__SCAN_IN), .B2(n16678), .ZN(n19128) );
  INV_X1 U15592 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n17119) );
  OAI21_X1 U15593 ( .B1(n13863), .B2(n13862), .A(n13861), .ZN(n18229) );
  OAI222_X1 U15594 ( .A1(n19403), .A2(n19128), .B1(n19401), .B2(n17119), .C1(
        n18229), .C2(n19410), .ZN(P2_U2908) );
  XNOR2_X1 U15595 ( .A(n13865), .B(n13864), .ZN(n18621) );
  INV_X1 U15596 ( .A(n13866), .ZN(n13867) );
  NOR2_X1 U15597 ( .A1(n13868), .A2(n13867), .ZN(n14143) );
  XOR2_X1 U15598 ( .A(n18621), .B(n14143), .Z(n14141) );
  XNOR2_X1 U15599 ( .A(n14141), .B(n17077), .ZN(n13871) );
  INV_X1 U15600 ( .A(BUF2_REG_2__SCAN_IN), .ZN(n20139) );
  AOI22_X1 U15601 ( .A1(n16679), .A2(n13789), .B1(n20139), .B2(n16678), .ZN(
        n19554) );
  AOI22_X1 U15602 ( .A1(n19130), .A2(n19554), .B1(n19652), .B2(
        P2_EAX_REG_2__SCAN_IN), .ZN(n13870) );
  NAND2_X1 U15603 ( .A1(n18621), .A2(n19548), .ZN(n13869) );
  OAI211_X1 U15604 ( .C1(n13871), .C2(n19659), .A(n13870), .B(n13869), .ZN(
        P2_U2917) );
  XNOR2_X1 U15605 ( .A(n13873), .B(n13872), .ZN(n14096) );
  AND2_X1 U15606 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n14930) );
  OAI21_X1 U15607 ( .B1(n15984), .B2(n14930), .A(n15982), .ZN(n14880) );
  AOI21_X1 U15608 ( .B1(n15987), .B2(n14879), .A(n14880), .ZN(n14320) );
  INV_X1 U15609 ( .A(n14320), .ZN(n14105) );
  AOI21_X1 U15610 ( .B1(n14930), .B2(n15981), .A(n15987), .ZN(n14933) );
  NOR2_X1 U15611 ( .A1(n14879), .A2(n14933), .ZN(n14477) );
  AOI22_X1 U15612 ( .A1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n14105), .B1(
        n14477), .B2(n12406), .ZN(n13878) );
  OAI21_X1 U15613 ( .B1(n13875), .B2(n13874), .A(n14100), .ZN(n13918) );
  INV_X1 U15614 ( .A(n13918), .ZN(n13971) );
  INV_X1 U15615 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n13876) );
  NOR2_X1 U15616 ( .A1(n21386), .A2(n13876), .ZN(n14090) );
  AOI21_X1 U15617 ( .B1(n21409), .B2(n13971), .A(n14090), .ZN(n13877) );
  OAI211_X1 U15618 ( .C1(n14096), .C2(n21353), .A(n13878), .B(n13877), .ZN(
        P1_U3028) );
  OR2_X1 U15619 ( .A1(n13880), .A2(n13879), .ZN(n13882) );
  NAND2_X1 U15620 ( .A1(n13882), .A2(n13881), .ZN(n18161) );
  INV_X1 U15621 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n16688) );
  NOR2_X1 U15622 ( .A1(n13893), .A2(n16688), .ZN(n13884) );
  OR2_X1 U15623 ( .A1(n13893), .A2(n13883), .ZN(n13959) );
  OAI211_X1 U15624 ( .C1(n13884), .C2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A(
        n16141), .B(n13959), .ZN(n13886) );
  NAND2_X1 U15625 ( .A1(n16157), .A2(P2_EBX_REG_6__SCAN_IN), .ZN(n13885) );
  OAI211_X1 U15626 ( .C1(n18161), .C2(n16111), .A(n13886), .B(n13885), .ZN(
        P2_U2881) );
  NAND2_X1 U15627 ( .A1(n13888), .A2(n13887), .ZN(n13889) );
  NAND2_X1 U15628 ( .A1(n13890), .A2(n13889), .ZN(n18581) );
  OR2_X1 U15629 ( .A1(n13839), .A2(n13891), .ZN(n13892) );
  NAND2_X1 U15630 ( .A1(n13893), .A2(n13892), .ZN(n19405) );
  INV_X1 U15631 ( .A(n19405), .ZN(n13894) );
  NAND2_X1 U15632 ( .A1(n13894), .A2(n16141), .ZN(n13896) );
  NAND2_X1 U15633 ( .A1(n16157), .A2(P2_EBX_REG_4__SCAN_IN), .ZN(n13895) );
  OAI211_X1 U15634 ( .C1(n18581), .C2(n16111), .A(n13896), .B(n13895), .ZN(
        P2_U2883) );
  INV_X1 U15635 ( .A(n22169), .ZN(n13912) );
  INV_X1 U15636 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n20067) );
  INV_X1 U15637 ( .A(DATAI_16_), .ZN(n13899) );
  OAI22_X1 U15638 ( .A1(n20067), .A2(n14243), .B1(n13899), .B2(n13898), .ZN(
        n21921) );
  INV_X1 U15639 ( .A(n21921), .ZN(n21903) );
  AND2_X1 U15640 ( .A1(n21909), .A2(n12300), .ZN(n13907) );
  NAND2_X1 U15641 ( .A1(n14157), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n21796) );
  OR2_X1 U15642 ( .A1(n21860), .A2(n13978), .ZN(n21811) );
  INV_X1 U15643 ( .A(n21811), .ZN(n14410) );
  AND2_X1 U15644 ( .A1(n13900), .A2(n16743), .ZN(n21904) );
  AOI21_X1 U15645 ( .B1(n14410), .B2(n21904), .A(n13901), .ZN(n13906) );
  OAI211_X1 U15646 ( .C1(n14158), .C2(n21796), .A(n21857), .B(n13906), .ZN(
        n13903) );
  INV_X1 U15647 ( .A(n21320), .ZN(n21684) );
  OAI211_X1 U15648 ( .C1(n21857), .C2(n13907), .A(n13903), .B(n21918), .ZN(
        n14277) );
  NAND2_X1 U15649 ( .A1(n14277), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n13911) );
  INV_X1 U15650 ( .A(DATAI_24_), .ZN(n16793) );
  INV_X1 U15651 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n20084) );
  OAI22_X2 U15652 ( .A1(n16793), .A2(n13898), .B1(n20084), .B2(n14243), .ZN(
        n21900) );
  INV_X1 U15653 ( .A(n21913), .ZN(n21865) );
  INV_X1 U15654 ( .A(n13906), .ZN(n13908) );
  AOI22_X1 U15655 ( .A1(n13908), .A2(n21857), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n13907), .ZN(n14278) );
  INV_X1 U15656 ( .A(n21914), .ZN(n21876) );
  OAI22_X1 U15657 ( .A1(n21865), .A2(n14279), .B1(n14278), .B2(n21876), .ZN(
        n13909) );
  AOI21_X1 U15658 ( .B1(n22162), .B2(n21900), .A(n13909), .ZN(n13910) );
  OAI211_X1 U15659 ( .C1(n13912), .C2(n21903), .A(n13911), .B(n13910), .ZN(
        P1_U3089) );
  OAI21_X1 U15660 ( .B1(n13914), .B2(n13913), .A(n14204), .ZN(n14089) );
  INV_X1 U15661 ( .A(BUF1_REG_3__SCAN_IN), .ZN(n13915) );
  OR2_X1 U15662 ( .A1(n14376), .A2(n13915), .ZN(n13917) );
  NAND2_X1 U15663 ( .A1(n14376), .A2(DATAI_3_), .ZN(n13916) );
  AND2_X1 U15664 ( .A1(n13917), .A2(n13916), .ZN(n14334) );
  INV_X1 U15665 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n19862) );
  OAI222_X1 U15666 ( .A1(n14089), .A2(n15711), .B1(n15701), .B2(n14334), .C1(
        n15703), .C2(n19862), .ZN(P1_U2901) );
  INV_X1 U15667 ( .A(P1_EBX_REG_3__SCAN_IN), .ZN(n13919) );
  OAI222_X1 U15668 ( .A1(n14089), .A2(n19966), .B1(n19969), .B2(n13919), .C1(
        n13918), .C2(n19965), .ZN(P1_U2869) );
  INV_X1 U15669 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n13922) );
  NAND2_X1 U15670 ( .A1(n15227), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n13921) );
  NAND2_X1 U15671 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n13920) );
  OAI211_X1 U15672 ( .C1(n10963), .C2(n13922), .A(n13921), .B(n13920), .ZN(
        n13923) );
  AOI21_X1 U15673 ( .B1(n13924), .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n13923), .ZN(n13925) );
  AND2_X1 U15674 ( .A1(n13926), .A2(n13925), .ZN(n13927) );
  OR2_X1 U15675 ( .A1(n13927), .A2(n14287), .ZN(n18215) );
  INV_X1 U15676 ( .A(n13928), .ZN(n13930) );
  OAI21_X1 U15677 ( .B1(n13931), .B2(n13930), .A(n13929), .ZN(n13932) );
  NAND3_X1 U15678 ( .A1(n13932), .A2(n16141), .A3(n14285), .ZN(n13934) );
  NAND2_X1 U15679 ( .A1(n16157), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n13933) );
  OAI211_X1 U15680 ( .C1(n18215), .C2(n16111), .A(n13934), .B(n13933), .ZN(
        P2_U2877) );
  INV_X1 U15681 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n20099) );
  OAI22_X1 U15682 ( .A1(n13935), .A2(n13898), .B1(n20099), .B2(n14243), .ZN(
        n22203) );
  NAND2_X1 U15683 ( .A1(n14277), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n13940) );
  INV_X1 U15684 ( .A(DATAI_23_), .ZN(n16886) );
  INV_X1 U15685 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n20082) );
  OAI22_X1 U15686 ( .A1(n16886), .A2(n13898), .B1(n20082), .B2(n14243), .ZN(
        n22214) );
  NOR2_X2 U15687 ( .A1(n14244), .A2(n15506), .ZN(n22210) );
  INV_X1 U15688 ( .A(n22210), .ZN(n22187) );
  OR2_X1 U15689 ( .A1(n14376), .A2(BUF1_REG_7__SCAN_IN), .ZN(n13937) );
  INV_X1 U15690 ( .A(DATAI_7_), .ZN(n16912) );
  NAND2_X1 U15691 ( .A1(n14376), .A2(n16912), .ZN(n13936) );
  NAND2_X1 U15692 ( .A1(n13937), .A2(n13936), .ZN(n14787) );
  INV_X1 U15693 ( .A(n22211), .ZN(n22193) );
  OAI22_X1 U15694 ( .A1(n22187), .A2(n14279), .B1(n14278), .B2(n22193), .ZN(
        n13938) );
  AOI21_X1 U15695 ( .B1(n22169), .B2(n22214), .A(n13938), .ZN(n13939) );
  OAI211_X1 U15696 ( .C1(n14283), .C2(n11083), .A(n13940), .B(n13939), .ZN(
        P1_U3096) );
  INV_X1 U15697 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n20091) );
  INV_X1 U15698 ( .A(DATAI_27_), .ZN(n16882) );
  INV_X1 U15699 ( .A(n22018), .ZN(n22027) );
  NAND2_X1 U15700 ( .A1(n14277), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n13943) );
  INV_X1 U15701 ( .A(DATAI_19_), .ZN(n16889) );
  INV_X1 U15702 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n20073) );
  OAI22_X1 U15703 ( .A1(n16889), .A2(n13898), .B1(n20073), .B2(n14243), .ZN(
        n22024) );
  NOR2_X2 U15704 ( .A1(n14244), .A2(n12523), .ZN(n22022) );
  INV_X1 U15705 ( .A(n22022), .ZN(n22011) );
  INV_X1 U15706 ( .A(n22023), .ZN(n22015) );
  OAI22_X1 U15707 ( .A1(n22011), .A2(n14279), .B1(n14278), .B2(n22015), .ZN(
        n13941) );
  AOI21_X1 U15708 ( .B1(n22169), .B2(n22024), .A(n13941), .ZN(n13942) );
  OAI211_X1 U15709 ( .C1(n14283), .C2(n22027), .A(n13943), .B(n13942), .ZN(
        P1_U3092) );
  INV_X1 U15710 ( .A(n21449), .ZN(n14086) );
  NOR2_X1 U15711 ( .A1(n13945), .A2(n13944), .ZN(n13968) );
  INV_X1 U15712 ( .A(n13968), .ZN(n21431) );
  NOR2_X1 U15713 ( .A1(P1_REIP_REG_2__SCAN_IN), .A2(n21439), .ZN(n13967) );
  OAI22_X1 U15714 ( .A1(n13947), .A2(n21640), .B1(n21646), .B2(n13946), .ZN(
        n13948) );
  AOI21_X1 U15715 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n13967), .A(n13948), .ZN(
        n13951) );
  INV_X1 U15716 ( .A(n21439), .ZN(n21602) );
  INV_X1 U15717 ( .A(n21422), .ZN(n21459) );
  AOI21_X1 U15718 ( .B1(n19947), .B2(n21602), .A(n21459), .ZN(n13949) );
  INV_X1 U15719 ( .A(n13949), .ZN(n13966) );
  NAND2_X1 U15720 ( .A1(P1_REIP_REG_2__SCAN_IN), .A2(n13966), .ZN(n13950) );
  OAI211_X1 U15721 ( .C1(n21860), .C2(n21431), .A(n13951), .B(n13950), .ZN(
        n13956) );
  NOR2_X1 U15722 ( .A1(n21642), .A2(n13954), .ZN(n13955) );
  AOI211_X1 U15723 ( .C1(n21645), .C2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .A(
        n13956), .B(n13955), .ZN(n13957) );
  OAI21_X1 U15724 ( .B1(n13958), .B2(n14086), .A(n13957), .ZN(P1_U2838) );
  XOR2_X1 U15725 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B(n13959), .Z(n13965)
         );
  NAND2_X1 U15726 ( .A1(n13960), .A2(n13881), .ZN(n13963) );
  INV_X1 U15727 ( .A(n13961), .ZN(n13962) );
  NAND2_X1 U15728 ( .A1(n13963), .A2(n13962), .ZN(n18175) );
  INV_X1 U15729 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n18171) );
  MUX2_X1 U15730 ( .A(n18175), .B(n18171), .S(n16111), .Z(n13964) );
  OAI21_X1 U15731 ( .B1(n13965), .B2(n16167), .A(n13964), .ZN(P2_U2880) );
  OAI21_X1 U15732 ( .B1(n13967), .B2(n13966), .A(P1_REIP_REG_3__SCAN_IN), .ZN(
        n13970) );
  NAND2_X1 U15733 ( .A1(n21769), .A2(n13968), .ZN(n13969) );
  OAI211_X1 U15734 ( .C1(n21642), .C2(n14092), .A(n13970), .B(n13969), .ZN(
        n13975) );
  NAND3_X1 U15735 ( .A1(P1_REIP_REG_2__SCAN_IN), .A2(P1_REIP_REG_1__SCAN_IN), 
        .A3(n21602), .ZN(n13973) );
  AOI22_X1 U15736 ( .A1(P1_EBX_REG_3__SCAN_IN), .A2(n21626), .B1(n21633), .B2(
        n13971), .ZN(n13972) );
  OAI21_X1 U15737 ( .B1(P1_REIP_REG_3__SCAN_IN), .B2(n13973), .A(n13972), .ZN(
        n13974) );
  AOI211_X1 U15738 ( .C1(n21645), .C2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A(
        n13975), .B(n13974), .ZN(n13976) );
  OAI21_X1 U15739 ( .B1(n14086), .B2(n14089), .A(n13976), .ZN(P1_U2837) );
  NAND2_X1 U15740 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n21656), .ZN(n13988) );
  INV_X1 U15741 ( .A(n13977), .ZN(n13987) );
  INV_X1 U15742 ( .A(n13978), .ZN(n21859) );
  NOR2_X1 U15743 ( .A1(n13979), .A2(n21859), .ZN(n13980) );
  XOR2_X1 U15744 ( .A(n11775), .B(n13980), .Z(n21432) );
  NOR2_X1 U15745 ( .A1(n21432), .A2(n12348), .ZN(n13985) );
  INV_X1 U15746 ( .A(n13983), .ZN(n16748) );
  AOI22_X1 U15747 ( .A1(n16748), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n13981), .B2(n13983), .ZN(n16752) );
  AOI22_X1 U15748 ( .A1(n16748), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n13982), .B2(n13983), .ZN(n16738) );
  OAI22_X1 U15749 ( .A1(n13983), .A2(n11775), .B1(n16752), .B2(n16738), .ZN(
        n13984) );
  OAI21_X1 U15750 ( .B1(n13985), .B2(n13984), .A(n16772), .ZN(n13986) );
  OAI21_X1 U15751 ( .B1(n13988), .B2(n13987), .A(n13986), .ZN(n16759) );
  INV_X1 U15752 ( .A(n16011), .ZN(n13990) );
  INV_X1 U15753 ( .A(n13988), .ZN(n13989) );
  AOI22_X1 U15754 ( .A1(n16759), .A2(n13990), .B1(n13989), .B2(
        P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n13991) );
  INV_X1 U15755 ( .A(n13991), .ZN(n21668) );
  NOR2_X1 U15756 ( .A1(n21668), .A2(P1_FLUSH_REG_SCAN_IN), .ZN(n13992) );
  OAI21_X1 U15757 ( .B1(n13992), .B2(n21680), .A(n21771), .ZN(n21674) );
  INV_X1 U15758 ( .A(n21674), .ZN(n14119) );
  AOI21_X1 U15759 ( .B1(n14401), .B2(n21796), .A(n21915), .ZN(n14121) );
  INV_X1 U15760 ( .A(n21796), .ZN(n14113) );
  NAND2_X1 U15761 ( .A1(n11056), .A2(n14113), .ZN(n14108) );
  INV_X1 U15762 ( .A(n21860), .ZN(n21768) );
  NOR2_X1 U15763 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n16772), .ZN(n21670) );
  INV_X1 U15764 ( .A(n21670), .ZN(n14116) );
  AOI22_X1 U15765 ( .A1(n14121), .A2(n14108), .B1(n21768), .B2(n14116), .ZN(
        n13994) );
  OR2_X1 U15766 ( .A1(n21674), .A2(n11700), .ZN(n13993) );
  OAI21_X1 U15767 ( .B1(n14119), .B2(n13994), .A(n13993), .ZN(P1_U3476) );
  MUX2_X1 U15768 ( .A(n19559), .B(n13995), .S(n19676), .Z(n14011) );
  INV_X1 U15769 ( .A(n13996), .ZN(n13997) );
  OAI21_X1 U15770 ( .B1(n13998), .B2(n13997), .A(n18090), .ZN(n14056) );
  NAND2_X1 U15771 ( .A1(n14056), .A2(n13999), .ZN(n14009) );
  AND2_X1 U15772 ( .A1(n19464), .A2(n14000), .ZN(n14006) );
  NAND3_X1 U15773 ( .A1(n14003), .A2(n14002), .A3(n14001), .ZN(n14004) );
  OAI211_X1 U15774 ( .C1(n14006), .C2(n13247), .A(n14005), .B(n14004), .ZN(
        n14007) );
  AOI21_X1 U15775 ( .B1(n14009), .B2(n14008), .A(n14007), .ZN(n14010) );
  OR2_X1 U15776 ( .A1(n14816), .A2(n15032), .ZN(n14022) );
  OR2_X1 U15777 ( .A1(n15030), .A2(n14046), .ZN(n14024) );
  NOR2_X1 U15778 ( .A1(n12875), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n14025) );
  INV_X1 U15779 ( .A(n14025), .ZN(n14030) );
  NAND2_X1 U15780 ( .A1(n14012), .A2(n14013), .ZN(n14014) );
  NAND2_X1 U15781 ( .A1(n14014), .A2(n13142), .ZN(n14015) );
  AOI21_X1 U15782 ( .B1(n14024), .B2(n14030), .A(n14015), .ZN(n14020) );
  AOI21_X1 U15783 ( .B1(n12790), .B2(n15031), .A(n16058), .ZN(n14031) );
  INV_X1 U15784 ( .A(n14031), .ZN(n14017) );
  NAND2_X1 U15785 ( .A1(n14012), .A2(n12867), .ZN(n14016) );
  NAND2_X1 U15786 ( .A1(n14017), .A2(n14016), .ZN(n14018) );
  NOR2_X1 U15787 ( .A1(n14025), .A2(n14018), .ZN(n14019) );
  MUX2_X1 U15788 ( .A(n14020), .B(n14019), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n14021) );
  AND2_X1 U15789 ( .A1(n14022), .A2(n14021), .ZN(n16660) );
  NOR2_X1 U15790 ( .A1(n14058), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n14023) );
  AOI21_X1 U15791 ( .B1(n16660), .B2(n14058), .A(n14023), .ZN(n14075) );
  OR2_X1 U15792 ( .A1(n14807), .A2(n15032), .ZN(n14036) );
  OAI21_X1 U15793 ( .B1(n16058), .B2(n14025), .A(n14024), .ZN(n14034) );
  INV_X1 U15794 ( .A(n14026), .ZN(n14029) );
  NAND2_X1 U15795 ( .A1(n14027), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n14028) );
  NAND2_X1 U15796 ( .A1(n14029), .A2(n14028), .ZN(n14032) );
  AOI22_X1 U15797 ( .A1(n14012), .A2(n14032), .B1(n14031), .B2(n14030), .ZN(
        n14033) );
  AND2_X1 U15798 ( .A1(n14034), .A2(n14033), .ZN(n14035) );
  NAND2_X1 U15799 ( .A1(n14036), .A2(n14035), .ZN(n16657) );
  INV_X1 U15800 ( .A(n16657), .ZN(n14038) );
  NOR2_X1 U15801 ( .A1(n14058), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n14037) );
  AOI21_X1 U15802 ( .B1(n14038), .B2(n14058), .A(n14037), .ZN(n14074) );
  NOR3_X1 U15803 ( .A1(n14040), .A2(n14992), .A3(n14039), .ZN(n18650) );
  OAI21_X1 U15804 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(P2_MORE_REG_SCAN_IN), .A(
        n18650), .ZN(n14041) );
  INV_X1 U15805 ( .A(n14041), .ZN(n14042) );
  AOI211_X1 U15806 ( .C1(n14045), .C2(n14044), .A(n14043), .B(n14042), .ZN(
        n14053) );
  INV_X1 U15807 ( .A(n18638), .ZN(n15007) );
  NAND2_X1 U15808 ( .A1(n16640), .A2(n14046), .ZN(n14049) );
  AOI22_X1 U15809 ( .A1(n15013), .A2(n14047), .B1(n15004), .B2(n15043), .ZN(
        n14048) );
  OAI211_X1 U15810 ( .C1(n15007), .C2(n14050), .A(n14049), .B(n14048), .ZN(
        n14051) );
  AOI21_X1 U15811 ( .B1(n14052), .B2(n15030), .A(n14051), .ZN(n18652) );
  OAI211_X1 U15812 ( .C1(n14054), .C2(n14058), .A(n14053), .B(n18652), .ZN(
        n14073) );
  INV_X1 U15813 ( .A(n14074), .ZN(n14068) );
  INV_X1 U15814 ( .A(n15032), .ZN(n14060) );
  INV_X1 U15815 ( .A(n13550), .ZN(n14055) );
  NAND2_X1 U15816 ( .A1(n14056), .A2(n14055), .ZN(n14061) );
  MUX2_X1 U15817 ( .A(n14061), .B(n14012), .S(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Z(n14057) );
  AOI21_X1 U15818 ( .B1(n18521), .B2(n14060), .A(n14057), .ZN(n16644) );
  INV_X1 U15819 ( .A(n14058), .ZN(n14059) );
  AOI21_X1 U15820 ( .B1(n16644), .B2(n19232), .A(n14059), .ZN(n14066) );
  NAND2_X1 U15821 ( .A1(n18526), .A2(n14060), .ZN(n14064) );
  NOR2_X1 U15822 ( .A1(n12873), .A2(n12875), .ZN(n14062) );
  AOI22_X1 U15823 ( .A1(n14012), .A2(n12648), .B1(n14062), .B2(n14061), .ZN(
        n14063) );
  AND2_X1 U15824 ( .A1(n14064), .A2(n14063), .ZN(n16650) );
  OAI211_X1 U15825 ( .C1(n16644), .C2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(
        n16650), .B(n19280), .ZN(n14065) );
  OAI211_X1 U15826 ( .C1(n14074), .C2(n19231), .A(n14066), .B(n14065), .ZN(
        n14067) );
  OAI21_X1 U15827 ( .B1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n14068), .A(
        n14067), .ZN(n14069) );
  OAI21_X1 U15828 ( .B1(n14075), .B2(n19200), .A(n14069), .ZN(n14071) );
  NAND2_X1 U15829 ( .A1(n14075), .A2(n19200), .ZN(n14070) );
  AOI21_X1 U15830 ( .B1(n14071), .B2(n14070), .A(
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n14072) );
  AOI211_X1 U15831 ( .C1(n14075), .C2(n14074), .A(n14073), .B(n14072), .ZN(
        n18648) );
  NAND3_X1 U15832 ( .A1(n18648), .A2(P2_STATE2_REG_2__SCAN_IN), .A3(n16719), 
        .ZN(n14079) );
  OR2_X1 U15833 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n14076), .ZN(n16025) );
  NOR3_X1 U15834 ( .A1(n11133), .A2(n18090), .A3(n16025), .ZN(n14077) );
  AOI21_X1 U15835 ( .B1(n14079), .B2(n14078), .A(n14077), .ZN(n18641) );
  OAI21_X1 U15836 ( .B1(n18641), .B2(n13554), .A(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n14080) );
  INV_X1 U15837 ( .A(n16721), .ZN(n18637) );
  NAND2_X1 U15838 ( .A1(n14080), .A2(n18637), .ZN(P2_U3593) );
  OAI21_X1 U15839 ( .B1(n21645), .B2(n21627), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n14085) );
  INV_X1 U15840 ( .A(n16743), .ZN(n21669) );
  NOR2_X1 U15841 ( .A1(n21669), .A2(n21431), .ZN(n14083) );
  OAI22_X1 U15842 ( .A1(n21640), .A2(n14081), .B1(n21407), .B2(n21646), .ZN(
        n14082) );
  AOI211_X1 U15843 ( .C1(n21639), .C2(P1_REIP_REG_0__SCAN_IN), .A(n14083), .B(
        n14082), .ZN(n14084) );
  OAI211_X1 U15844 ( .C1(n14086), .C2(n19977), .A(n14085), .B(n14084), .ZN(
        P1_U2840) );
  AOI22_X1 U15845 ( .A1(n16679), .A2(BUF1_REG_12__SCAN_IN), .B1(
        BUF2_REG_12__SCAN_IN), .B2(n16226), .ZN(n19125) );
  AOI21_X1 U15846 ( .B1(n13861), .B2(n14087), .A(n14292), .ZN(n18246) );
  INV_X1 U15847 ( .A(n18246), .ZN(n14088) );
  INV_X1 U15848 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n17121) );
  OAI222_X1 U15849 ( .A1(n19403), .A2(n19125), .B1(n14088), .B2(n19410), .C1(
        n19401), .C2(n17121), .ZN(P2_U2907) );
  INV_X1 U15850 ( .A(n14089), .ZN(n14094) );
  AOI21_X1 U15851 ( .B1(n20022), .B2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A(
        n14090), .ZN(n14091) );
  OAI21_X1 U15852 ( .B1(n20028), .B2(n14092), .A(n14091), .ZN(n14093) );
  AOI21_X1 U15853 ( .B1(n14094), .B2(n20009), .A(n14093), .ZN(n14095) );
  OAI21_X1 U15854 ( .B1(n14096), .B2(n21655), .A(n14095), .ZN(P1_U2996) );
  XNOR2_X1 U15855 ( .A(n14098), .B(n14097), .ZN(n14212) );
  NAND2_X1 U15856 ( .A1(n14100), .A2(n14099), .ZN(n14101) );
  NAND2_X1 U15857 ( .A1(n14258), .A2(n14101), .ZN(n21433) );
  NAND2_X1 U15858 ( .A1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n14318) );
  OAI211_X1 U15859 ( .C1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A(n14477), .B(n14318), .ZN(n14103) );
  INV_X1 U15860 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n21437) );
  NOR2_X1 U15861 ( .A1(n21386), .A2(n21437), .ZN(n14208) );
  INV_X1 U15862 ( .A(n14208), .ZN(n14102) );
  OAI211_X1 U15863 ( .C1(n21352), .C2(n21433), .A(n14103), .B(n14102), .ZN(
        n14104) );
  AOI21_X1 U15864 ( .B1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n14105), .A(
        n14104), .ZN(n14106) );
  OAI21_X1 U15865 ( .B1(n21353), .B2(n14212), .A(n14106), .ZN(P1_U3027) );
  OAI21_X1 U15866 ( .B1(n21885), .B2(n21796), .A(n21857), .ZN(n21920) );
  AOI21_X1 U15867 ( .B1(n12407), .B2(n14108), .A(n21920), .ZN(n14109) );
  AOI21_X1 U15868 ( .B1(n14116), .B2(n21769), .A(n14109), .ZN(n14111) );
  NAND2_X1 U15869 ( .A1(n14119), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n14110) );
  OAI21_X1 U15870 ( .B1(n14119), .B2(n14111), .A(n14110), .ZN(P1_U3475) );
  INV_X1 U15871 ( .A(n10973), .ZN(n21890) );
  INV_X1 U15872 ( .A(n14157), .ZN(n14114) );
  AOI211_X1 U15873 ( .C1(n14114), .C2(n14152), .A(n21915), .B(n14113), .ZN(
        n14115) );
  AOI21_X1 U15874 ( .B1(n21890), .B2(n14116), .A(n14115), .ZN(n14118) );
  NAND2_X1 U15875 ( .A1(n14119), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n14117) );
  OAI21_X1 U15876 ( .B1(n14119), .B2(n14118), .A(n14117), .ZN(P1_U3477) );
  NAND3_X1 U15877 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n11700), .ZN(n21846) );
  INV_X1 U15878 ( .A(n21846), .ZN(n14120) );
  AOI21_X1 U15879 ( .B1(n21822), .B2(n14121), .A(n14120), .ZN(n14123) );
  INV_X1 U15880 ( .A(n21918), .ZN(n14122) );
  INV_X1 U15881 ( .A(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n14128) );
  AND2_X1 U15882 ( .A1(n21769), .A2(n21860), .ZN(n21842) );
  NOR2_X1 U15883 ( .A1(n21877), .A2(n21846), .ZN(n14266) );
  AOI21_X1 U15884 ( .B1(n21842), .B2(n21904), .A(n14266), .ZN(n14124) );
  OAI22_X1 U15885 ( .A1(n14124), .A2(n21915), .B1(n21846), .B2(n21910), .ZN(
        n14267) );
  AOI22_X1 U15886 ( .A1(n14267), .A2(n21914), .B1(n21913), .B2(n14266), .ZN(
        n14125) );
  OAI21_X1 U15887 ( .B1(n14269), .B2(n21903), .A(n14125), .ZN(n14126) );
  AOI21_X1 U15888 ( .B1(n21900), .B2(n22180), .A(n14126), .ZN(n14127) );
  OAI21_X1 U15889 ( .B1(n14273), .B2(n14128), .A(n14127), .ZN(P1_U3121) );
  INV_X1 U15890 ( .A(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n14132) );
  INV_X1 U15891 ( .A(n22214), .ZN(n22208) );
  AOI22_X1 U15892 ( .A1(n14267), .A2(n22211), .B1(n22210), .B2(n14266), .ZN(
        n14129) );
  OAI21_X1 U15893 ( .B1(n14269), .B2(n22208), .A(n14129), .ZN(n14130) );
  AOI21_X1 U15894 ( .B1(n11084), .B2(n22180), .A(n14130), .ZN(n14131) );
  OAI21_X1 U15895 ( .B1(n14273), .B2(n14132), .A(n14131), .ZN(P1_U3128) );
  INV_X1 U15896 ( .A(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n14136) );
  INV_X1 U15897 ( .A(n22024), .ZN(n22021) );
  AOI22_X1 U15898 ( .A1(n14267), .A2(n22023), .B1(n22022), .B2(n14266), .ZN(
        n14133) );
  OAI21_X1 U15899 ( .B1(n14269), .B2(n22021), .A(n14133), .ZN(n14134) );
  AOI21_X1 U15900 ( .B1(n22018), .B2(n22180), .A(n14134), .ZN(n14135) );
  OAI21_X1 U15901 ( .B1(n14273), .B2(n14136), .A(n14135), .ZN(P1_U3124) );
  OR2_X1 U15902 ( .A1(n14138), .A2(n14137), .ZN(n14140) );
  NAND2_X1 U15903 ( .A1(n14140), .A2(n14139), .ZN(n18595) );
  NAND2_X1 U15904 ( .A1(n14141), .A2(n17077), .ZN(n14146) );
  INV_X1 U15905 ( .A(n18595), .ZN(n14142) );
  XNOR2_X1 U15906 ( .A(n19328), .B(n14142), .ZN(n14144) );
  NAND2_X1 U15907 ( .A1(n14143), .A2(n18621), .ZN(n14145) );
  NAND3_X1 U15908 ( .A1(n14146), .A2(n14144), .A3(n14145), .ZN(n14456) );
  INV_X1 U15909 ( .A(n14456), .ZN(n14148) );
  AOI21_X1 U15910 ( .B1(n14146), .B2(n14145), .A(n14144), .ZN(n14147) );
  INV_X1 U15911 ( .A(n19659), .ZN(n19549) );
  OAI21_X1 U15912 ( .B1(n14148), .B2(n14147), .A(n19549), .ZN(n14150) );
  AOI22_X1 U15913 ( .A1(n16679), .A2(BUF1_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n16226), .ZN(n19509) );
  INV_X1 U15914 ( .A(n19509), .ZN(n16246) );
  AOI22_X1 U15915 ( .A1(n19130), .A2(n16246), .B1(n19652), .B2(
        P2_EAX_REG_3__SCAN_IN), .ZN(n14149) );
  OAI211_X1 U15916 ( .C1(n18595), .C2(n19658), .A(n14150), .B(n14149), .ZN(
        P2_U2916) );
  NAND3_X1 U15917 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n12300), .A3(
        n21864), .ZN(n14404) );
  INV_X1 U15918 ( .A(n14404), .ZN(n14154) );
  INV_X1 U15919 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n14152) );
  INV_X1 U15920 ( .A(n14151), .ZN(n21878) );
  NOR2_X1 U15921 ( .A1(n21877), .A2(n14404), .ZN(n14245) );
  AOI21_X1 U15922 ( .B1(n14410), .B2(n21878), .A(n14245), .ZN(n14159) );
  OAI211_X1 U15923 ( .C1(n14158), .C2(n14152), .A(n21881), .B(n14159), .ZN(
        n14153) );
  OAI211_X1 U15924 ( .C1(n21881), .C2(n14154), .A(n14153), .B(n21918), .ZN(
        n14155) );
  INV_X1 U15925 ( .A(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n14163) );
  INV_X1 U15926 ( .A(n21855), .ZN(n14156) );
  OAI22_X1 U15927 ( .A1(n14159), .A2(n21915), .B1(n14404), .B2(n21910), .ZN(
        n14246) );
  AOI22_X1 U15928 ( .A1(n14246), .A2(n22211), .B1(n22210), .B2(n14245), .ZN(
        n14160) );
  OAI21_X1 U15929 ( .B1(n14248), .B2(n22208), .A(n14160), .ZN(n14161) );
  AOI21_X1 U15930 ( .B1(n14407), .B2(n11084), .A(n14161), .ZN(n14162) );
  OAI21_X1 U15931 ( .B1(n14252), .B2(n14163), .A(n14162), .ZN(P1_U3080) );
  INV_X1 U15932 ( .A(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n14170) );
  INV_X1 U15933 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n20095) );
  INV_X1 U15934 ( .A(DATAI_29_), .ZN(n16787) );
  INV_X1 U15935 ( .A(DATAI_21_), .ZN(n16894) );
  INV_X1 U15936 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n20077) );
  OAI22_X1 U15937 ( .A1(n16894), .A2(n13898), .B1(n20077), .B2(n14243), .ZN(
        n22095) );
  INV_X1 U15938 ( .A(n22095), .ZN(n22092) );
  INV_X1 U15939 ( .A(BUF1_REG_5__SCAN_IN), .ZN(n14164) );
  OR2_X1 U15940 ( .A1(n14376), .A2(n14164), .ZN(n14166) );
  NAND2_X1 U15941 ( .A1(n14376), .A2(DATAI_5_), .ZN(n14165) );
  AND2_X1 U15942 ( .A1(n14166), .A2(n14165), .ZN(n14367) );
  NOR2_X2 U15943 ( .A1(n14244), .A2(n11148), .ZN(n22093) );
  AOI22_X1 U15944 ( .A1(n14246), .A2(n22094), .B1(n22093), .B2(n14245), .ZN(
        n14167) );
  OAI21_X1 U15945 ( .B1(n14248), .B2(n22092), .A(n14167), .ZN(n14168) );
  AOI21_X1 U15946 ( .B1(n14407), .B2(n22089), .A(n14168), .ZN(n14169) );
  OAI21_X1 U15947 ( .B1(n14252), .B2(n14170), .A(n14169), .ZN(P1_U3078) );
  INV_X1 U15948 ( .A(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n14177) );
  INV_X1 U15949 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n20093) );
  INV_X1 U15950 ( .A(DATAI_28_), .ZN(n16783) );
  OAI22_X1 U15951 ( .A1(n20093), .A2(n14243), .B1(n16783), .B2(n13898), .ZN(
        n22053) );
  INV_X1 U15952 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n20075) );
  INV_X1 U15953 ( .A(DATAI_20_), .ZN(n16780) );
  OAI22_X1 U15954 ( .A1(n20075), .A2(n14243), .B1(n16780), .B2(n13898), .ZN(
        n22059) );
  INV_X1 U15955 ( .A(n22059), .ZN(n22056) );
  OR2_X1 U15956 ( .A1(n14376), .A2(BUF1_REG_4__SCAN_IN), .ZN(n14172) );
  INV_X1 U15957 ( .A(DATAI_4_), .ZN(n16923) );
  NAND2_X1 U15958 ( .A1(n14376), .A2(n16923), .ZN(n14171) );
  NAND2_X1 U15959 ( .A1(n14172), .A2(n14171), .ZN(n15668) );
  AOI22_X1 U15960 ( .A1(n14246), .A2(n22058), .B1(n22057), .B2(n14245), .ZN(
        n14174) );
  OAI21_X1 U15961 ( .B1(n14248), .B2(n22056), .A(n14174), .ZN(n14175) );
  AOI21_X1 U15962 ( .B1(n14407), .B2(n22053), .A(n14175), .ZN(n14176) );
  OAI21_X1 U15963 ( .B1(n14252), .B2(n14177), .A(n14176), .ZN(P1_U3077) );
  INV_X1 U15964 ( .A(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n14181) );
  AOI22_X1 U15965 ( .A1(n14246), .A2(n22023), .B1(n22022), .B2(n14245), .ZN(
        n14178) );
  OAI21_X1 U15966 ( .B1(n14248), .B2(n22021), .A(n14178), .ZN(n14179) );
  AOI21_X1 U15967 ( .B1(n14407), .B2(n22018), .A(n14179), .ZN(n14180) );
  OAI21_X1 U15968 ( .B1(n14252), .B2(n14181), .A(n14180), .ZN(P1_U3076) );
  INV_X1 U15969 ( .A(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n14186) );
  INV_X1 U15970 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n20088) );
  INV_X1 U15971 ( .A(DATAI_26_), .ZN(n16873) );
  OAI22_X1 U15972 ( .A1(n20088), .A2(n14243), .B1(n16873), .B2(n13898), .ZN(
        n21984) );
  INV_X1 U15973 ( .A(DATAI_18_), .ZN(n16899) );
  INV_X1 U15974 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n20071) );
  OAI22_X1 U15975 ( .A1(n16899), .A2(n13898), .B1(n20071), .B2(n14243), .ZN(
        n21990) );
  INV_X1 U15976 ( .A(n21990), .ZN(n21987) );
  NOR2_X2 U15977 ( .A1(n14244), .A2(n14182), .ZN(n21988) );
  AOI22_X1 U15978 ( .A1(n14246), .A2(n21989), .B1(n21988), .B2(n14245), .ZN(
        n14183) );
  OAI21_X1 U15979 ( .B1(n14248), .B2(n21987), .A(n14183), .ZN(n14184) );
  AOI21_X1 U15980 ( .B1(n14407), .B2(n21984), .A(n14184), .ZN(n14185) );
  OAI21_X1 U15981 ( .B1(n14252), .B2(n14186), .A(n14185), .ZN(P1_U3075) );
  INV_X1 U15982 ( .A(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n14190) );
  AOI22_X1 U15983 ( .A1(n14246), .A2(n21914), .B1(n21913), .B2(n14245), .ZN(
        n14187) );
  OAI21_X1 U15984 ( .B1(n14248), .B2(n21903), .A(n14187), .ZN(n14188) );
  AOI21_X1 U15985 ( .B1(n14407), .B2(n21900), .A(n14188), .ZN(n14189) );
  OAI21_X1 U15986 ( .B1(n14252), .B2(n14190), .A(n14189), .ZN(P1_U3073) );
  INV_X1 U15987 ( .A(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n14194) );
  AOI22_X1 U15988 ( .A1(n14267), .A2(n22094), .B1(n22093), .B2(n14266), .ZN(
        n14191) );
  OAI21_X1 U15989 ( .B1(n14269), .B2(n22092), .A(n14191), .ZN(n14192) );
  AOI21_X1 U15990 ( .B1(n22089), .B2(n22180), .A(n14192), .ZN(n14193) );
  OAI21_X1 U15991 ( .B1(n14273), .B2(n14194), .A(n14193), .ZN(P1_U3126) );
  INV_X1 U15992 ( .A(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n14198) );
  AOI22_X1 U15993 ( .A1(n14267), .A2(n22058), .B1(n22057), .B2(n14266), .ZN(
        n14195) );
  OAI21_X1 U15994 ( .B1(n14269), .B2(n22056), .A(n14195), .ZN(n14196) );
  AOI21_X1 U15995 ( .B1(n22053), .B2(n22180), .A(n14196), .ZN(n14197) );
  OAI21_X1 U15996 ( .B1(n14273), .B2(n14198), .A(n14197), .ZN(P1_U3125) );
  INV_X1 U15997 ( .A(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n14202) );
  AOI22_X1 U15998 ( .A1(n14267), .A2(n21989), .B1(n21988), .B2(n14266), .ZN(
        n14199) );
  OAI21_X1 U15999 ( .B1(n14269), .B2(n21987), .A(n14199), .ZN(n14200) );
  AOI21_X1 U16000 ( .B1(n21984), .B2(n22180), .A(n14200), .ZN(n14201) );
  OAI21_X1 U16001 ( .B1(n14273), .B2(n14202), .A(n14201), .ZN(P1_U3123) );
  OR2_X1 U16002 ( .A1(n14204), .A2(n14205), .ZN(n14253) );
  INV_X1 U16003 ( .A(n14253), .ZN(n14203) );
  AOI21_X1 U16004 ( .B1(n14205), .B2(n14204), .A(n14203), .ZN(n21441) );
  INV_X1 U16005 ( .A(n21441), .ZN(n14305) );
  INV_X1 U16006 ( .A(n21433), .ZN(n14206) );
  AOI22_X1 U16007 ( .A1(n19961), .A2(n14206), .B1(n15617), .B2(
        P1_EBX_REG_4__SCAN_IN), .ZN(n14207) );
  OAI21_X1 U16008 ( .B1(n14305), .B2(n19966), .A(n14207), .ZN(P1_U2868) );
  AOI21_X1 U16009 ( .B1(n20022), .B2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n14208), .ZN(n14209) );
  OAI21_X1 U16010 ( .B1(n20028), .B2(n21444), .A(n14209), .ZN(n14210) );
  AOI21_X1 U16011 ( .B1(n21441), .B2(n20009), .A(n14210), .ZN(n14211) );
  OAI21_X1 U16012 ( .B1(n21655), .B2(n14212), .A(n14211), .ZN(P1_U2995) );
  INV_X1 U16013 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15249) );
  AOI22_X1 U16014 ( .A1(n15227), .A2(P2_EBX_REG_11__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), 
        .ZN(n14214) );
  NAND2_X1 U16015 ( .A1(n15440), .A2(P2_REIP_REG_11__SCAN_IN), .ZN(n14213) );
  OAI211_X1 U16016 ( .C1(n15443), .C2(n15249), .A(n14214), .B(n14213), .ZN(
        n14286) );
  INV_X1 U16017 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n14217) );
  NAND2_X1 U16018 ( .A1(n15227), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n14216) );
  NAND2_X1 U16019 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n14215) );
  OAI211_X1 U16020 ( .C1(n10963), .C2(n14217), .A(n14216), .B(n14215), .ZN(
        n14218) );
  AOI21_X1 U16021 ( .B1(n13924), .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n14218), .ZN(n14219) );
  INV_X1 U16022 ( .A(n14219), .ZN(n14221) );
  OAI21_X1 U16023 ( .B1(n14220), .B2(n14221), .A(n14489), .ZN(n18249) );
  INV_X1 U16024 ( .A(n14222), .ZN(n14284) );
  OAI21_X1 U16025 ( .B1(n14285), .B2(n14284), .A(n14223), .ZN(n14224) );
  NAND3_X1 U16026 ( .A1(n11427), .A2(n16141), .A3(n14224), .ZN(n14226) );
  NAND2_X1 U16027 ( .A1(n16111), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n14225) );
  OAI211_X1 U16028 ( .C1(n18249), .C2(n16111), .A(n14226), .B(n14225), .ZN(
        P2_U2875) );
  INV_X1 U16029 ( .A(n22089), .ZN(n22098) );
  NAND2_X1 U16030 ( .A1(n14277), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n14229) );
  INV_X1 U16031 ( .A(n22093), .ZN(n22082) );
  INV_X1 U16032 ( .A(n22094), .ZN(n22086) );
  OAI22_X1 U16033 ( .A1(n22082), .A2(n14279), .B1(n14278), .B2(n22086), .ZN(
        n14227) );
  AOI21_X1 U16034 ( .B1(n22169), .B2(n22095), .A(n14227), .ZN(n14228) );
  OAI211_X1 U16035 ( .C1(n14283), .C2(n22098), .A(n14229), .B(n14228), .ZN(
        P1_U3094) );
  INV_X1 U16036 ( .A(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n14235) );
  INV_X1 U16037 ( .A(BUF1_REG_30__SCAN_IN), .ZN(n20097) );
  INV_X1 U16038 ( .A(DATAI_30_), .ZN(n16879) );
  INV_X1 U16039 ( .A(DATAI_22_), .ZN(n16895) );
  INV_X1 U16040 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n20079) );
  OAI22_X1 U16041 ( .A1(n16895), .A2(n13898), .B1(n20079), .B2(n14243), .ZN(
        n22129) );
  INV_X1 U16042 ( .A(n22129), .ZN(n22126) );
  OR2_X1 U16043 ( .A1(n14376), .A2(BUF1_REG_6__SCAN_IN), .ZN(n14231) );
  INV_X1 U16044 ( .A(DATAI_6_), .ZN(n16914) );
  NAND2_X1 U16045 ( .A1(n14376), .A2(n16914), .ZN(n14230) );
  NAND2_X1 U16046 ( .A1(n14231), .A2(n14230), .ZN(n15660) );
  NOR2_X2 U16047 ( .A1(n14244), .A2(n11631), .ZN(n22127) );
  AOI22_X1 U16048 ( .A1(n14246), .A2(n22128), .B1(n22127), .B2(n14245), .ZN(
        n14232) );
  OAI21_X1 U16049 ( .B1(n14248), .B2(n22126), .A(n14232), .ZN(n14233) );
  AOI21_X1 U16050 ( .B1(n14407), .B2(n22123), .A(n14233), .ZN(n14234) );
  OAI21_X1 U16051 ( .B1(n14252), .B2(n14235), .A(n14234), .ZN(P1_U3079) );
  INV_X1 U16052 ( .A(n22053), .ZN(n22062) );
  NAND2_X1 U16053 ( .A1(n14277), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n14238) );
  INV_X1 U16054 ( .A(n22057), .ZN(n22046) );
  OAI22_X1 U16055 ( .A1(n22046), .A2(n14279), .B1(n14278), .B2(n22050), .ZN(
        n14236) );
  AOI21_X1 U16056 ( .B1(n22169), .B2(n22059), .A(n14236), .ZN(n14237) );
  OAI211_X1 U16057 ( .C1(n14283), .C2(n22062), .A(n14238), .B(n14237), .ZN(
        P1_U3093) );
  INV_X1 U16058 ( .A(n21984), .ZN(n21993) );
  NAND2_X1 U16059 ( .A1(n14277), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n14241) );
  INV_X1 U16060 ( .A(n21988), .ZN(n21977) );
  INV_X1 U16061 ( .A(n21989), .ZN(n21981) );
  OAI22_X1 U16062 ( .A1(n21977), .A2(n14279), .B1(n14278), .B2(n21981), .ZN(
        n14239) );
  AOI21_X1 U16063 ( .B1(n22169), .B2(n21990), .A(n14239), .ZN(n14240) );
  OAI211_X1 U16064 ( .C1(n14283), .C2(n21993), .A(n14241), .B(n14240), .ZN(
        P1_U3091) );
  INV_X1 U16065 ( .A(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n14251) );
  INV_X1 U16066 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n20086) );
  INV_X1 U16067 ( .A(DATAI_25_), .ZN(n14242) );
  INV_X1 U16068 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n20069) );
  INV_X1 U16069 ( .A(DATAI_17_), .ZN(n16803) );
  OAI22_X1 U16070 ( .A1(n20069), .A2(n14243), .B1(n16803), .B2(n13898), .ZN(
        n21955) );
  INV_X1 U16071 ( .A(n21955), .ZN(n21952) );
  NOR2_X2 U16072 ( .A1(n14244), .A2(n14298), .ZN(n21953) );
  AOI22_X1 U16073 ( .A1(n14246), .A2(n21954), .B1(n21953), .B2(n14245), .ZN(
        n14247) );
  OAI21_X1 U16074 ( .B1(n14248), .B2(n21952), .A(n14247), .ZN(n14249) );
  AOI21_X1 U16075 ( .B1(n14407), .B2(n21949), .A(n14249), .ZN(n14250) );
  OAI21_X1 U16076 ( .B1(n14252), .B2(n14251), .A(n14250), .ZN(P1_U3074) );
  AND2_X1 U16077 ( .A1(n14254), .A2(n14253), .ZN(n14256) );
  OR2_X1 U16078 ( .A1(n14256), .A2(n14255), .ZN(n21445) );
  AND2_X1 U16079 ( .A1(n14258), .A2(n14257), .ZN(n14259) );
  OR2_X1 U16080 ( .A1(n14310), .A2(n14259), .ZN(n21453) );
  INV_X1 U16081 ( .A(n21453), .ZN(n14260) );
  AOI22_X1 U16082 ( .A1(n19961), .A2(n14260), .B1(n15617), .B2(
        P1_EBX_REG_5__SCAN_IN), .ZN(n14261) );
  OAI21_X1 U16083 ( .B1(n21445), .B2(n19966), .A(n14261), .ZN(P1_U2867) );
  INV_X1 U16084 ( .A(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n14265) );
  AOI22_X1 U16085 ( .A1(n14267), .A2(n22128), .B1(n22127), .B2(n14266), .ZN(
        n14262) );
  OAI21_X1 U16086 ( .B1(n14269), .B2(n22126), .A(n14262), .ZN(n14263) );
  AOI21_X1 U16087 ( .B1(n22123), .B2(n22180), .A(n14263), .ZN(n14264) );
  OAI21_X1 U16088 ( .B1(n14273), .B2(n14265), .A(n14264), .ZN(P1_U3127) );
  INV_X1 U16089 ( .A(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n14272) );
  AOI22_X1 U16090 ( .A1(n14267), .A2(n21954), .B1(n21953), .B2(n14266), .ZN(
        n14268) );
  OAI21_X1 U16091 ( .B1(n14269), .B2(n21952), .A(n14268), .ZN(n14270) );
  AOI21_X1 U16092 ( .B1(n21949), .B2(n22180), .A(n14270), .ZN(n14271) );
  OAI21_X1 U16093 ( .B1(n14273), .B2(n14272), .A(n14271), .ZN(P1_U3122) );
  INV_X1 U16094 ( .A(n22123), .ZN(n22132) );
  NAND2_X1 U16095 ( .A1(n14277), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n14276) );
  INV_X1 U16096 ( .A(n22127), .ZN(n22116) );
  INV_X1 U16097 ( .A(n22128), .ZN(n22120) );
  OAI22_X1 U16098 ( .A1(n22116), .A2(n14279), .B1(n14278), .B2(n22120), .ZN(
        n14274) );
  AOI21_X1 U16099 ( .B1(n22169), .B2(n22129), .A(n14274), .ZN(n14275) );
  OAI211_X1 U16100 ( .C1(n14283), .C2(n22132), .A(n14276), .B(n14275), .ZN(
        P1_U3095) );
  INV_X1 U16101 ( .A(n21949), .ZN(n21958) );
  NAND2_X1 U16102 ( .A1(n14277), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n14282) );
  INV_X1 U16103 ( .A(n21953), .ZN(n21942) );
  INV_X1 U16104 ( .A(n21954), .ZN(n21946) );
  OAI22_X1 U16105 ( .A1(n21942), .A2(n14279), .B1(n14278), .B2(n21946), .ZN(
        n14280) );
  AOI21_X1 U16106 ( .B1(n22169), .B2(n21955), .A(n14280), .ZN(n14281) );
  OAI211_X1 U16107 ( .C1(n14283), .C2(n21958), .A(n14282), .B(n14281), .ZN(
        P1_U3090) );
  OAI222_X1 U16108 ( .A1(n21445), .A2(n15711), .B1(n15701), .B2(n14367), .C1(
        n15703), .C2(n11769), .ZN(P1_U2899) );
  XNOR2_X1 U16109 ( .A(n14285), .B(n14284), .ZN(n14291) );
  OR2_X1 U16110 ( .A1(n14287), .A2(n14286), .ZN(n14288) );
  AND2_X1 U16111 ( .A1(n14289), .A2(n14288), .ZN(n17018) );
  INV_X1 U16112 ( .A(n17018), .ZN(n18230) );
  INV_X1 U16113 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n18225) );
  MUX2_X1 U16114 ( .A(n18230), .B(n18225), .S(n16111), .Z(n14290) );
  OAI21_X1 U16115 ( .B1(n14291), .B2(n16167), .A(n14290), .ZN(P2_U2876) );
  NOR2_X1 U16116 ( .A1(n14293), .A2(n14292), .ZN(n14294) );
  OR2_X1 U16117 ( .A1(n14450), .A2(n14294), .ZN(n18258) );
  INV_X1 U16118 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n17123) );
  OAI222_X1 U16119 ( .A1(n19403), .A2(n19122), .B1(n18258), .B2(n19410), .C1(
        n19401), .C2(n17123), .ZN(P2_U2906) );
  NAND2_X2 U16120 ( .A1(n14297), .A2(n14298), .ZN(n14393) );
  INV_X1 U16121 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n15702) );
  NAND2_X1 U16122 ( .A1(n14295), .A2(n21712), .ZN(n14296) );
  NOR2_X2 U16123 ( .A1(n14395), .A2(n14298), .ZN(n14379) );
  INV_X1 U16124 ( .A(n14379), .ZN(n14304) );
  INV_X1 U16125 ( .A(DATAI_15_), .ZN(n14299) );
  NOR2_X1 U16126 ( .A1(n14301), .A2(n14299), .ZN(n14300) );
  AOI21_X1 U16127 ( .B1(n14301), .B2(BUF1_REG_15__SCAN_IN), .A(n14300), .ZN(
        n15700) );
  INV_X1 U16128 ( .A(P1_LWORD_REG_15__SCAN_IN), .ZN(n14303) );
  OAI222_X1 U16129 ( .A1(n14393), .A2(n15702), .B1(n14304), .B2(n15700), .C1(
        n14303), .C2(n14302), .ZN(P1_U2967) );
  INV_X1 U16130 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n19864) );
  OAI222_X1 U16131 ( .A1(n15701), .A2(n15668), .B1(n15703), .B2(n19864), .C1(
        n15711), .C2(n14305), .ZN(P1_U2900) );
  OR2_X1 U16132 ( .A1(n14255), .A2(n14307), .ZN(n14308) );
  AND2_X1 U16133 ( .A1(n14306), .A2(n14308), .ZN(n14474) );
  INV_X1 U16134 ( .A(n14474), .ZN(n21461) );
  OR2_X1 U16135 ( .A1(n14310), .A2(n14309), .ZN(n14311) );
  NAND2_X1 U16136 ( .A1(n14464), .A2(n14311), .ZN(n21454) );
  INV_X1 U16137 ( .A(n21454), .ZN(n14479) );
  AOI22_X1 U16138 ( .A1(n19961), .A2(n14479), .B1(n15617), .B2(
        P1_EBX_REG_6__SCAN_IN), .ZN(n14312) );
  OAI21_X1 U16139 ( .B1(n21461), .B2(n19966), .A(n14312), .ZN(P1_U2866) );
  XNOR2_X1 U16140 ( .A(n14314), .B(n14313), .ZN(n19979) );
  INV_X1 U16141 ( .A(n19979), .ZN(n14323) );
  INV_X1 U16142 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n14319) );
  AND2_X1 U16143 ( .A1(n14477), .A2(n14319), .ZN(n14317) );
  INV_X1 U16144 ( .A(n14318), .ZN(n14316) );
  NAND2_X1 U16145 ( .A1(n10970), .A2(P1_REIP_REG_5__SCAN_IN), .ZN(n19980) );
  OAI21_X1 U16146 ( .B1(n21352), .B2(n21453), .A(n19980), .ZN(n14315) );
  AOI21_X1 U16147 ( .B1(n14317), .B2(n14316), .A(n14315), .ZN(n14322) );
  NOR2_X1 U16148 ( .A1(n14319), .A2(n14318), .ZN(n14878) );
  OAI21_X1 U16149 ( .B1(n21351), .B2(n14878), .A(n14320), .ZN(n14482) );
  NAND2_X1 U16150 ( .A1(n14482), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n14321) );
  OAI211_X1 U16151 ( .C1(n14323), .C2(n21353), .A(n14322), .B(n14321), .ZN(
        P1_U3026) );
  INV_X1 U16152 ( .A(n15677), .ZN(n14324) );
  NAND2_X1 U16153 ( .A1(n14379), .A2(n14324), .ZN(n14357) );
  NAND2_X1 U16154 ( .A1(n14398), .A2(P1_LWORD_REG_2__SCAN_IN), .ZN(n14325) );
  OAI211_X1 U16155 ( .C1(n19860), .C2(n14393), .A(n14357), .B(n14325), .ZN(
        P1_U2954) );
  INV_X1 U16156 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n19875) );
  OR2_X1 U16157 ( .A1(n14376), .A2(BUF1_REG_10__SCAN_IN), .ZN(n14327) );
  INV_X1 U16158 ( .A(DATAI_10_), .ZN(n16872) );
  NAND2_X1 U16159 ( .A1(n14376), .A2(n16872), .ZN(n14326) );
  NAND2_X1 U16160 ( .A1(n14327), .A2(n14326), .ZN(n15642) );
  INV_X1 U16161 ( .A(n15642), .ZN(n14328) );
  NAND2_X1 U16162 ( .A1(n14379), .A2(n14328), .ZN(n14338) );
  NAND2_X1 U16163 ( .A1(n14398), .A2(P1_LWORD_REG_10__SCAN_IN), .ZN(n14329) );
  OAI211_X1 U16164 ( .C1(n19875), .C2(n14393), .A(n14338), .B(n14329), .ZN(
        P1_U2962) );
  MUX2_X1 U16165 ( .A(BUF1_REG_12__SCAN_IN), .B(DATAI_12_), .S(n14376), .Z(
        n15633) );
  NAND2_X1 U16166 ( .A1(n14379), .A2(n15633), .ZN(n14333) );
  NAND2_X1 U16167 ( .A1(n14398), .A2(P1_UWORD_REG_12__SCAN_IN), .ZN(n14330) );
  OAI211_X1 U16168 ( .C1(n14331), .C2(n14393), .A(n14333), .B(n14330), .ZN(
        P1_U2949) );
  INV_X1 U16169 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n19879) );
  NAND2_X1 U16170 ( .A1(n14398), .A2(P1_LWORD_REG_12__SCAN_IN), .ZN(n14332) );
  OAI211_X1 U16171 ( .C1(n19879), .C2(n14393), .A(n14333), .B(n14332), .ZN(
        P1_U2964) );
  INV_X1 U16172 ( .A(n14334), .ZN(n15672) );
  NAND2_X1 U16173 ( .A1(n14379), .A2(n15672), .ZN(n14354) );
  NAND2_X1 U16174 ( .A1(n14398), .A2(P1_LWORD_REG_3__SCAN_IN), .ZN(n14335) );
  OAI211_X1 U16175 ( .C1(n19862), .C2(n14393), .A(n14354), .B(n14335), .ZN(
        P1_U2955) );
  INV_X1 U16176 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n19883) );
  MUX2_X1 U16177 ( .A(BUF1_REG_14__SCAN_IN), .B(DATAI_14_), .S(n14376), .Z(
        n15708) );
  NAND2_X1 U16178 ( .A1(n14379), .A2(n15708), .ZN(n14385) );
  NAND2_X1 U16179 ( .A1(n14398), .A2(P1_LWORD_REG_14__SCAN_IN), .ZN(n14336) );
  OAI211_X1 U16180 ( .C1(n19883), .C2(n14393), .A(n14385), .B(n14336), .ZN(
        P1_U2966) );
  NAND2_X1 U16181 ( .A1(n14395), .A2(P1_UWORD_REG_10__SCAN_IN), .ZN(n14337) );
  OAI211_X1 U16182 ( .C1(n14339), .C2(n14393), .A(n14338), .B(n14337), .ZN(
        P1_U2947) );
  OR2_X1 U16183 ( .A1(n14376), .A2(BUF1_REG_9__SCAN_IN), .ZN(n14341) );
  INV_X1 U16184 ( .A(DATAI_9_), .ZN(n16915) );
  NAND2_X1 U16185 ( .A1(n14376), .A2(n16915), .ZN(n14340) );
  NAND2_X1 U16186 ( .A1(n14341), .A2(n14340), .ZN(n15647) );
  INV_X1 U16187 ( .A(n15647), .ZN(n14342) );
  NAND2_X1 U16188 ( .A1(n14379), .A2(n14342), .ZN(n14400) );
  NAND2_X1 U16189 ( .A1(n14395), .A2(P1_UWORD_REG_9__SCAN_IN), .ZN(n14343) );
  OAI211_X1 U16190 ( .C1(n15646), .C2(n14393), .A(n14400), .B(n14343), .ZN(
        P1_U2946) );
  INV_X1 U16191 ( .A(n14344), .ZN(n15683) );
  NAND2_X1 U16192 ( .A1(n14379), .A2(n15683), .ZN(n14359) );
  NAND2_X1 U16193 ( .A1(n14398), .A2(P1_LWORD_REG_1__SCAN_IN), .ZN(n14345) );
  OAI211_X1 U16194 ( .C1(n19858), .C2(n14393), .A(n14359), .B(n14345), .ZN(
        P1_U2953) );
  INV_X1 U16195 ( .A(n14787), .ZN(n15656) );
  NAND2_X1 U16196 ( .A1(n14379), .A2(n15656), .ZN(n14390) );
  NAND2_X1 U16197 ( .A1(n14395), .A2(P1_UWORD_REG_7__SCAN_IN), .ZN(n14346) );
  OAI211_X1 U16198 ( .C1(n14347), .C2(n14393), .A(n14390), .B(n14346), .ZN(
        P1_U2944) );
  INV_X1 U16199 ( .A(n15660), .ZN(n14348) );
  NAND2_X1 U16200 ( .A1(n14379), .A2(n14348), .ZN(n14351) );
  NAND2_X1 U16201 ( .A1(n14395), .A2(P1_UWORD_REG_6__SCAN_IN), .ZN(n14349) );
  OAI211_X1 U16202 ( .C1(n15659), .C2(n14393), .A(n14351), .B(n14349), .ZN(
        P1_U2943) );
  NAND2_X1 U16203 ( .A1(n14395), .A2(P1_LWORD_REG_6__SCAN_IN), .ZN(n14350) );
  OAI211_X1 U16204 ( .C1(n11847), .C2(n14393), .A(n14351), .B(n14350), .ZN(
        P1_U2958) );
  INV_X1 U16205 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n19881) );
  MUX2_X1 U16206 ( .A(BUF1_REG_13__SCAN_IN), .B(DATAI_13_), .S(n14376), .Z(
        n15507) );
  NAND2_X1 U16207 ( .A1(n14379), .A2(n15507), .ZN(n14374) );
  NAND2_X1 U16208 ( .A1(n14398), .A2(P1_LWORD_REG_13__SCAN_IN), .ZN(n14352) );
  OAI211_X1 U16209 ( .C1(n19881), .C2(n14393), .A(n14374), .B(n14352), .ZN(
        P1_U2965) );
  NAND2_X1 U16210 ( .A1(n14395), .A2(P1_UWORD_REG_3__SCAN_IN), .ZN(n14353) );
  OAI211_X1 U16211 ( .C1(n14355), .C2(n14393), .A(n14354), .B(n14353), .ZN(
        P1_U2940) );
  NAND2_X1 U16212 ( .A1(n14395), .A2(P1_UWORD_REG_2__SCAN_IN), .ZN(n14356) );
  OAI211_X1 U16213 ( .C1(n15675), .C2(n14393), .A(n14357), .B(n14356), .ZN(
        P1_U2939) );
  NAND2_X1 U16214 ( .A1(n14395), .A2(P1_UWORD_REG_1__SCAN_IN), .ZN(n14358) );
  OAI211_X1 U16215 ( .C1(n14360), .C2(n14393), .A(n14359), .B(n14358), .ZN(
        P1_U2938) );
  INV_X1 U16216 ( .A(n15690), .ZN(n14361) );
  NAND2_X1 U16217 ( .A1(n14379), .A2(n14361), .ZN(n14388) );
  NAND2_X1 U16218 ( .A1(n14395), .A2(P1_UWORD_REG_0__SCAN_IN), .ZN(n14362) );
  OAI211_X1 U16219 ( .C1(n15688), .C2(n14393), .A(n14388), .B(n14362), .ZN(
        P1_U2937) );
  INV_X1 U16220 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n19871) );
  OR2_X1 U16221 ( .A1(n14376), .A2(BUF1_REG_8__SCAN_IN), .ZN(n14364) );
  INV_X1 U16222 ( .A(DATAI_8_), .ZN(n16911) );
  NAND2_X1 U16223 ( .A1(n14376), .A2(n16911), .ZN(n14363) );
  NAND2_X1 U16224 ( .A1(n14364), .A2(n14363), .ZN(n15652) );
  INV_X1 U16225 ( .A(n15652), .ZN(n14365) );
  NAND2_X1 U16226 ( .A1(n14379), .A2(n14365), .ZN(n14397) );
  NAND2_X1 U16227 ( .A1(n14398), .A2(P1_LWORD_REG_8__SCAN_IN), .ZN(n14366) );
  OAI211_X1 U16228 ( .C1(n19871), .C2(n14393), .A(n14397), .B(n14366), .ZN(
        P1_U2960) );
  INV_X1 U16229 ( .A(n14367), .ZN(n15664) );
  NAND2_X1 U16230 ( .A1(n14379), .A2(n15664), .ZN(n14392) );
  NAND2_X1 U16231 ( .A1(n14398), .A2(P1_LWORD_REG_5__SCAN_IN), .ZN(n14368) );
  OAI211_X1 U16232 ( .C1(n11769), .C2(n14393), .A(n14392), .B(n14368), .ZN(
        P1_U2957) );
  INV_X1 U16233 ( .A(n15668), .ZN(n14369) );
  NAND2_X1 U16234 ( .A1(n14379), .A2(n14369), .ZN(n14372) );
  NAND2_X1 U16235 ( .A1(n14398), .A2(P1_LWORD_REG_4__SCAN_IN), .ZN(n14370) );
  OAI211_X1 U16236 ( .C1(n19864), .C2(n14393), .A(n14372), .B(n14370), .ZN(
        P1_U2956) );
  NAND2_X1 U16237 ( .A1(n14395), .A2(P1_UWORD_REG_4__SCAN_IN), .ZN(n14371) );
  OAI211_X1 U16238 ( .C1(n15667), .C2(n14393), .A(n14372), .B(n14371), .ZN(
        P1_U2941) );
  NAND2_X1 U16239 ( .A1(n14398), .A2(P1_UWORD_REG_13__SCAN_IN), .ZN(n14373) );
  OAI211_X1 U16240 ( .C1(n14375), .C2(n14393), .A(n14374), .B(n14373), .ZN(
        P1_U2950) );
  INV_X1 U16241 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n19877) );
  OR2_X1 U16242 ( .A1(n14376), .A2(BUF1_REG_11__SCAN_IN), .ZN(n14378) );
  INV_X1 U16243 ( .A(DATAI_11_), .ZN(n16811) );
  NAND2_X1 U16244 ( .A1(n14376), .A2(n16811), .ZN(n14377) );
  NAND2_X1 U16245 ( .A1(n14378), .A2(n14377), .ZN(n15079) );
  INV_X1 U16246 ( .A(n15079), .ZN(n15637) );
  NAND2_X1 U16247 ( .A1(n14379), .A2(n15637), .ZN(n14382) );
  NAND2_X1 U16248 ( .A1(n14398), .A2(P1_LWORD_REG_11__SCAN_IN), .ZN(n14380) );
  OAI211_X1 U16249 ( .C1(n19877), .C2(n14393), .A(n14382), .B(n14380), .ZN(
        P1_U2963) );
  NAND2_X1 U16250 ( .A1(n14398), .A2(P1_UWORD_REG_11__SCAN_IN), .ZN(n14381) );
  OAI211_X1 U16251 ( .C1(n14383), .C2(n14393), .A(n14382), .B(n14381), .ZN(
        P1_U2948) );
  NAND2_X1 U16252 ( .A1(n14398), .A2(P1_UWORD_REG_14__SCAN_IN), .ZN(n14384) );
  OAI211_X1 U16253 ( .C1(n14386), .C2(n14393), .A(n14385), .B(n14384), .ZN(
        P1_U2951) );
  NAND2_X1 U16254 ( .A1(n14398), .A2(P1_LWORD_REG_0__SCAN_IN), .ZN(n14387) );
  OAI211_X1 U16255 ( .C1(n19856), .C2(n14393), .A(n14388), .B(n14387), .ZN(
        P1_U2952) );
  NAND2_X1 U16256 ( .A1(n14395), .A2(P1_LWORD_REG_7__SCAN_IN), .ZN(n14389) );
  OAI211_X1 U16257 ( .C1(n11859), .C2(n14393), .A(n14390), .B(n14389), .ZN(
        P1_U2959) );
  NAND2_X1 U16258 ( .A1(n14395), .A2(P1_UWORD_REG_5__SCAN_IN), .ZN(n14391) );
  OAI211_X1 U16259 ( .C1(n14394), .C2(n14393), .A(n14392), .B(n14391), .ZN(
        P1_U2942) );
  NAND2_X1 U16260 ( .A1(n14395), .A2(P1_UWORD_REG_8__SCAN_IN), .ZN(n14396) );
  OAI211_X1 U16261 ( .C1(n14393), .C2(n15651), .A(n14397), .B(n14396), .ZN(
        P1_U2945) );
  INV_X1 U16262 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n19873) );
  NAND2_X1 U16263 ( .A1(n14398), .A2(P1_LWORD_REG_9__SCAN_IN), .ZN(n14399) );
  OAI211_X1 U16264 ( .C1(n19873), .C2(n14393), .A(n14400), .B(n14399), .ZN(
        P1_U2961) );
  OAI222_X1 U16265 ( .A1(n15701), .A2(n15660), .B1(n15703), .B2(n11847), .C1(
        n15711), .C2(n21461), .ZN(P1_U2898) );
  INV_X1 U16266 ( .A(n14402), .ZN(n21766) );
  OAI21_X1 U16267 ( .B1(n22155), .B2(n14407), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n14403) );
  OAI21_X1 U16268 ( .B1(n21890), .B2(n21811), .A(n14403), .ZN(n14405) );
  NOR2_X1 U16269 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n14404), .ZN(
        n14442) );
  AOI21_X1 U16270 ( .B1(n14405), .B2(n21868), .A(n14442), .ZN(n14406) );
  NOR2_X1 U16271 ( .A1(n14408), .A2(n21910), .ZN(n21845) );
  INV_X1 U16272 ( .A(n21898), .ZN(n21814) );
  INV_X1 U16273 ( .A(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n14416) );
  INV_X1 U16274 ( .A(n21823), .ZN(n21843) );
  NOR2_X1 U16275 ( .A1(n21824), .A2(n21843), .ZN(n21776) );
  INV_X1 U16276 ( .A(n21776), .ZN(n14412) );
  INV_X1 U16277 ( .A(n14408), .ZN(n14409) );
  NOR2_X1 U16278 ( .A1(n14409), .A2(n21910), .ZN(n21862) );
  INV_X1 U16279 ( .A(n21862), .ZN(n21893) );
  NAND3_X1 U16280 ( .A1(n14410), .A2(n21857), .A3(n10973), .ZN(n14411) );
  OAI21_X1 U16281 ( .B1(n14412), .B2(n21893), .A(n14411), .ZN(n14441) );
  AOI22_X1 U16282 ( .A1(n21988), .A2(n14442), .B1(n21989), .B2(n14441), .ZN(
        n14413) );
  OAI21_X1 U16283 ( .B1(n14444), .B2(n21987), .A(n14413), .ZN(n14414) );
  AOI21_X1 U16284 ( .B1(n22155), .B2(n21984), .A(n14414), .ZN(n14415) );
  OAI21_X1 U16285 ( .B1(n14448), .B2(n14416), .A(n14415), .ZN(P1_U3067) );
  INV_X1 U16286 ( .A(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n14420) );
  AOI22_X1 U16287 ( .A1(n21953), .A2(n14442), .B1(n21954), .B2(n14441), .ZN(
        n14417) );
  OAI21_X1 U16288 ( .B1(n14444), .B2(n21952), .A(n14417), .ZN(n14418) );
  AOI21_X1 U16289 ( .B1(n22155), .B2(n21949), .A(n14418), .ZN(n14419) );
  OAI21_X1 U16290 ( .B1(n14448), .B2(n14420), .A(n14419), .ZN(P1_U3066) );
  INV_X1 U16291 ( .A(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n14424) );
  AOI22_X1 U16292 ( .A1(n22210), .A2(n14442), .B1(n22211), .B2(n14441), .ZN(
        n14421) );
  OAI21_X1 U16293 ( .B1(n14444), .B2(n22208), .A(n14421), .ZN(n14422) );
  AOI21_X1 U16294 ( .B1(n22155), .B2(n11084), .A(n14422), .ZN(n14423) );
  OAI21_X1 U16295 ( .B1(n14448), .B2(n14424), .A(n14423), .ZN(P1_U3072) );
  INV_X1 U16296 ( .A(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n14428) );
  AOI22_X1 U16297 ( .A1(n22057), .A2(n14442), .B1(n22058), .B2(n14441), .ZN(
        n14425) );
  OAI21_X1 U16298 ( .B1(n14444), .B2(n22056), .A(n14425), .ZN(n14426) );
  AOI21_X1 U16299 ( .B1(n22155), .B2(n22053), .A(n14426), .ZN(n14427) );
  OAI21_X1 U16300 ( .B1(n14448), .B2(n14428), .A(n14427), .ZN(P1_U3069) );
  INV_X1 U16301 ( .A(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n14432) );
  AOI22_X1 U16302 ( .A1(n22093), .A2(n14442), .B1(n22094), .B2(n14441), .ZN(
        n14429) );
  OAI21_X1 U16303 ( .B1(n14444), .B2(n22092), .A(n14429), .ZN(n14430) );
  AOI21_X1 U16304 ( .B1(n22155), .B2(n22089), .A(n14430), .ZN(n14431) );
  OAI21_X1 U16305 ( .B1(n14448), .B2(n14432), .A(n14431), .ZN(P1_U3070) );
  INV_X1 U16306 ( .A(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n14436) );
  AOI22_X1 U16307 ( .A1(n21913), .A2(n14442), .B1(n21914), .B2(n14441), .ZN(
        n14433) );
  OAI21_X1 U16308 ( .B1(n14444), .B2(n21903), .A(n14433), .ZN(n14434) );
  AOI21_X1 U16309 ( .B1(n22155), .B2(n21900), .A(n14434), .ZN(n14435) );
  OAI21_X1 U16310 ( .B1(n14448), .B2(n14436), .A(n14435), .ZN(P1_U3065) );
  INV_X1 U16311 ( .A(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n14440) );
  AOI22_X1 U16312 ( .A1(n22127), .A2(n14442), .B1(n22128), .B2(n14441), .ZN(
        n14437) );
  OAI21_X1 U16313 ( .B1(n14444), .B2(n22126), .A(n14437), .ZN(n14438) );
  AOI21_X1 U16314 ( .B1(n22155), .B2(n22123), .A(n14438), .ZN(n14439) );
  OAI21_X1 U16315 ( .B1(n14448), .B2(n14440), .A(n14439), .ZN(P1_U3071) );
  INV_X1 U16316 ( .A(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n14447) );
  AOI22_X1 U16317 ( .A1(n22022), .A2(n14442), .B1(n22023), .B2(n14441), .ZN(
        n14443) );
  OAI21_X1 U16318 ( .B1(n14444), .B2(n22021), .A(n14443), .ZN(n14445) );
  AOI21_X1 U16319 ( .B1(n22155), .B2(n22018), .A(n14445), .ZN(n14446) );
  OAI21_X1 U16320 ( .B1(n14448), .B2(n14447), .A(n14446), .ZN(P1_U3068) );
  AOI22_X1 U16321 ( .A1(n16679), .A2(BUF1_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n16678), .ZN(n19119) );
  NOR2_X1 U16322 ( .A1(n14450), .A2(n14449), .ZN(n14451) );
  NOR2_X1 U16323 ( .A1(n14791), .A2(n14451), .ZN(n18538) );
  INV_X1 U16324 ( .A(n18538), .ZN(n14452) );
  INV_X1 U16325 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n17125) );
  OAI222_X1 U16326 ( .A1(n19403), .A2(n19119), .B1(n14452), .B2(n19410), .C1(
        n19401), .C2(n17125), .ZN(P2_U2905) );
  INV_X1 U16327 ( .A(BUF1_REG_4__SCAN_IN), .ZN(n20045) );
  INV_X1 U16328 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n20657) );
  AOI22_X1 U16329 ( .A1(n16679), .A2(n20045), .B1(n20657), .B2(n16226), .ZN(
        n19453) );
  INV_X1 U16330 ( .A(n19453), .ZN(n19462) );
  NAND2_X1 U16331 ( .A1(n19328), .A2(n18595), .ZN(n14455) );
  AOI21_X1 U16332 ( .B1(n14454), .B2(n14139), .A(n14453), .ZN(n18579) );
  AOI21_X1 U16333 ( .B1(n14456), .B2(n14455), .A(n18579), .ZN(n19406) );
  XOR2_X1 U16334 ( .A(n19405), .B(n19406), .Z(n14457) );
  NAND2_X1 U16335 ( .A1(n14457), .A2(n19549), .ZN(n14459) );
  AOI22_X1 U16336 ( .A1(n19548), .A2(n18579), .B1(n19652), .B2(
        P2_EAX_REG_4__SCAN_IN), .ZN(n14458) );
  OAI211_X1 U16337 ( .C1(n19462), .C2(n19403), .A(n14459), .B(n14458), .ZN(
        P2_U2915) );
  NAND2_X1 U16338 ( .A1(n14306), .A2(n14461), .ZN(n14462) );
  AND2_X1 U16339 ( .A1(n14460), .A2(n14462), .ZN(n21474) );
  INV_X1 U16340 ( .A(n21474), .ZN(n14786) );
  XNOR2_X1 U16341 ( .A(n14464), .B(n14463), .ZN(n21468) );
  INV_X1 U16342 ( .A(n21468), .ZN(n14465) );
  AOI22_X1 U16343 ( .A1(n19961), .A2(n14465), .B1(n15617), .B2(
        P1_EBX_REG_7__SCAN_IN), .ZN(n14466) );
  OAI21_X1 U16344 ( .B1(n14786), .B2(n19966), .A(n14466), .ZN(P1_U2865) );
  OAI21_X1 U16345 ( .B1(n14469), .B2(n14468), .A(n14467), .ZN(n14485) );
  NOR2_X1 U16346 ( .A1(n21386), .A2(n21463), .ZN(n14478) );
  AOI21_X1 U16347 ( .B1(n20022), .B2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n14478), .ZN(n14472) );
  INV_X1 U16348 ( .A(n21460), .ZN(n14470) );
  NAND2_X1 U16349 ( .A1(n20005), .A2(n14470), .ZN(n14471) );
  NAND2_X1 U16350 ( .A1(n14472), .A2(n14471), .ZN(n14473) );
  AOI21_X1 U16351 ( .B1(n14474), .B2(n20009), .A(n14473), .ZN(n14475) );
  OAI21_X1 U16352 ( .B1(n14485), .B2(n21655), .A(n14475), .ZN(P1_U2993) );
  NAND3_X1 U16353 ( .A1(n14878), .A2(n14477), .A3(n14476), .ZN(n14481) );
  AOI21_X1 U16354 ( .B1(n21409), .B2(n14479), .A(n14478), .ZN(n14480) );
  AND2_X1 U16355 ( .A1(n14481), .A2(n14480), .ZN(n14484) );
  NAND2_X1 U16356 ( .A1(n14482), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n14483) );
  OAI211_X1 U16357 ( .C1(n14485), .C2(n21353), .A(n14484), .B(n14483), .ZN(
        P1_U3025) );
  INV_X1 U16358 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n16391) );
  NAND2_X1 U16359 ( .A1(n15227), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n14487) );
  NAND2_X1 U16360 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n14486) );
  OAI211_X1 U16361 ( .C1(n15436), .C2(n16391), .A(n14487), .B(n14486), .ZN(
        n14488) );
  AOI21_X1 U16362 ( .B1(n13924), .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n14488), .ZN(n14516) );
  INV_X1 U16363 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n15191) );
  AOI22_X1 U16364 ( .A1(n15227), .A2(P2_EBX_REG_14__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), 
        .ZN(n14491) );
  NAND2_X1 U16365 ( .A1(n15440), .A2(P2_REIP_REG_14__SCAN_IN), .ZN(n14490) );
  OAI211_X1 U16366 ( .C1(n15443), .C2(n15191), .A(n14491), .B(n14490), .ZN(
        n14492) );
  NOR2_X1 U16367 ( .A1(n11043), .A2(n14492), .ZN(n14493) );
  OR2_X1 U16368 ( .A1(n14801), .A2(n14493), .ZN(n18540) );
  OAI211_X1 U16369 ( .C1(n14512), .C2(n14494), .A(n14794), .B(n16141), .ZN(
        n14496) );
  NAND2_X1 U16370 ( .A1(n16157), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n14495) );
  OAI211_X1 U16371 ( .C1(n18540), .C2(n16111), .A(n14496), .B(n14495), .ZN(
        P2_U2873) );
  XNOR2_X1 U16372 ( .A(n14460), .B(n14497), .ZN(n14919) );
  INV_X1 U16373 ( .A(n14919), .ZN(n14788) );
  NAND2_X1 U16374 ( .A1(n14499), .A2(n14498), .ZN(n14500) );
  NAND2_X1 U16375 ( .A1(n14872), .A2(n14500), .ZN(n14908) );
  INV_X1 U16376 ( .A(n14908), .ZN(n14501) );
  AOI22_X1 U16377 ( .A1(n19961), .A2(n14501), .B1(n15617), .B2(
        P1_EBX_REG_8__SCAN_IN), .ZN(n14502) );
  OAI21_X1 U16378 ( .B1(n14788), .B2(n19966), .A(n14502), .ZN(P1_U2864) );
  INV_X1 U16379 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n14503) );
  OAI22_X1 U16380 ( .A1(n14917), .A2(n21642), .B1(n21636), .B2(n14503), .ZN(
        n14507) );
  NAND2_X1 U16381 ( .A1(n21422), .A2(n14504), .ZN(n21571) );
  OAI22_X1 U16382 ( .A1(n14505), .A2(n21640), .B1(n21646), .B2(n14908), .ZN(
        n14506) );
  NOR3_X1 U16383 ( .A1(n14507), .A2(n21562), .A3(n14506), .ZN(n14511) );
  INV_X1 U16384 ( .A(P1_REIP_REG_8__SCAN_IN), .ZN(n19895) );
  NAND2_X1 U16385 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(n21488), .ZN(n14508) );
  NAND2_X1 U16386 ( .A1(n19895), .A2(n14508), .ZN(n14509) );
  NAND3_X1 U16387 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(P1_REIP_REG_7__SCAN_IN), 
        .A3(n21488), .ZN(n21487) );
  NAND3_X1 U16388 ( .A1(n14509), .A2(n21487), .A3(n21639), .ZN(n14510) );
  OAI211_X1 U16389 ( .C1(n14788), .C2(n21648), .A(n14511), .B(n14510), .ZN(
        P1_U2832) );
  INV_X1 U16390 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n14520) );
  INV_X1 U16391 ( .A(n14512), .ZN(n14513) );
  OAI211_X1 U16392 ( .C1(n14515), .C2(n14514), .A(n14513), .B(n16141), .ZN(
        n14519) );
  AND2_X1 U16393 ( .A1(n14489), .A2(n14516), .ZN(n14517) );
  OR2_X1 U16394 ( .A1(n14517), .A2(n11043), .ZN(n18259) );
  INV_X1 U16395 ( .A(n18259), .ZN(n16550) );
  NAND2_X1 U16396 ( .A1(n16550), .A2(n16102), .ZN(n14518) );
  OAI211_X1 U16397 ( .C1(n16102), .C2(n14520), .A(n14519), .B(n14518), .ZN(
        P2_U2874) );
  INV_X1 U16398 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n20882) );
  INV_X1 U16399 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n20881) );
  INV_X1 U16400 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n20894) );
  OAI21_X1 U16401 ( .B1(n20882), .B2(n20881), .A(n20894), .ZN(n20846) );
  INV_X1 U16402 ( .A(n20846), .ZN(n20885) );
  INV_X4 U16403 ( .A(n17391), .ZN(n17546) );
  AOI22_X1 U16404 ( .A1(n10967), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n10966), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n14521) );
  OAI21_X1 U16405 ( .B1(n17208), .B2(n17523), .A(n14521), .ZN(n14530) );
  AOI22_X1 U16406 ( .A1(n17539), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n17286), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n14528) );
  AOI22_X1 U16407 ( .A1(n14603), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n10965), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n14527) );
  NOR2_X2 U16408 ( .A1(n20829), .A2(n20192), .ZN(n20181) );
  NAND2_X1 U16409 ( .A1(n21260), .A2(n20181), .ZN(n20193) );
  AOI22_X1 U16410 ( .A1(n14589), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n20216), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n14526) );
  AOI22_X1 U16411 ( .A1(n10968), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n17540), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n14525) );
  NAND4_X1 U16412 ( .A1(n14528), .A2(n14527), .A3(n14526), .A4(n14525), .ZN(
        n14529) );
  AOI22_X1 U16413 ( .A1(n17539), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n17286), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n14543) );
  AOI22_X1 U16414 ( .A1(n10961), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n14603), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n14542) );
  INV_X1 U16415 ( .A(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n17347) );
  AOI22_X1 U16416 ( .A1(n10958), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n10967), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n14534) );
  OAI21_X1 U16417 ( .B1(n17208), .B2(n17347), .A(n14534), .ZN(n14540) );
  AOI22_X1 U16418 ( .A1(n10960), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n10971), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n14538) );
  AOI22_X1 U16419 ( .A1(n17546), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10965), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n14537) );
  AOI22_X1 U16420 ( .A1(n14589), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n20216), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n14536) );
  AOI22_X1 U16421 ( .A1(n10968), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n14682), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n14535) );
  NAND4_X1 U16422 ( .A1(n14538), .A2(n14537), .A3(n14536), .A4(n14535), .ZN(
        n14539) );
  INV_X2 U16423 ( .A(n20166), .ZN(n19013) );
  NOR2_X1 U16424 ( .A1(n14680), .A2(n19013), .ZN(n17149) );
  AOI22_X1 U16425 ( .A1(n17546), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n10976), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n14548) );
  CLKBUF_X3 U16426 ( .A(n14561), .Z(n17537) );
  AOI22_X1 U16427 ( .A1(n17205), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n17537), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n14547) );
  AOI22_X1 U16428 ( .A1(n17540), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n14589), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n14546) );
  AOI22_X1 U16429 ( .A1(n10968), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n20216), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n14545) );
  NAND4_X1 U16430 ( .A1(n14548), .A2(n14547), .A3(n14546), .A4(n14545), .ZN(
        n14555) );
  AOI22_X1 U16431 ( .A1(n10958), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n10967), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n14553) );
  AOI22_X1 U16432 ( .A1(n10977), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n10971), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n14552) );
  AOI22_X1 U16433 ( .A1(n17505), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17538), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n14551) );
  AOI22_X1 U16434 ( .A1(n14603), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n17539), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n14550) );
  NAND4_X1 U16435 ( .A1(n14553), .A2(n14552), .A3(n14551), .A4(n14550), .ZN(
        n14554) );
  AOI22_X1 U16436 ( .A1(n17545), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17548), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n14560) );
  AOI22_X1 U16437 ( .A1(n17505), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n10976), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n14559) );
  AOI22_X1 U16438 ( .A1(n17540), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n14589), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n14558) );
  AOI22_X1 U16439 ( .A1(n10968), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n20216), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n14557) );
  NAND4_X1 U16440 ( .A1(n14560), .A2(n14559), .A3(n14558), .A4(n14557), .ZN(
        n14567) );
  AOI22_X1 U16441 ( .A1(n17205), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17546), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n14565) );
  AOI22_X1 U16442 ( .A1(n17538), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n17539), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n14564) );
  AOI22_X1 U16443 ( .A1(n10958), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n10967), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n14563) );
  AOI22_X1 U16444 ( .A1(n10971), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17286), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n14562) );
  NAND4_X1 U16445 ( .A1(n14565), .A2(n14564), .A3(n14563), .A4(n14562), .ZN(
        n14566) );
  AOI22_X1 U16446 ( .A1(n10958), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n14603), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n14571) );
  AOI22_X1 U16447 ( .A1(n17538), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n10966), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n14570) );
  AOI22_X1 U16448 ( .A1(n10968), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n20216), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n14569) );
  AOI22_X1 U16449 ( .A1(n17540), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n14589), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n14568) );
  NAND4_X1 U16450 ( .A1(n14571), .A2(n14570), .A3(n14569), .A4(n14568), .ZN(
        n14578) );
  AOI22_X1 U16451 ( .A1(n10975), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17539), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n14576) );
  AOI22_X1 U16452 ( .A1(n10961), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17286), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n14575) );
  AOI22_X1 U16453 ( .A1(n17205), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17546), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n14574) );
  AOI22_X1 U16454 ( .A1(n10960), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10967), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n14573) );
  NAND4_X1 U16455 ( .A1(n14576), .A2(n14575), .A3(n14574), .A4(n14573), .ZN(
        n14577) );
  AOI22_X1 U16456 ( .A1(n10977), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17538), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n14582) );
  AOI22_X1 U16457 ( .A1(n17205), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n10966), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n14581) );
  AOI22_X1 U16458 ( .A1(n10968), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n14589), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n14580) );
  AOI22_X1 U16459 ( .A1(n17540), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n20216), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n14579) );
  NAND4_X1 U16460 ( .A1(n14582), .A2(n14581), .A3(n14580), .A4(n14579), .ZN(
        n14588) );
  AOI22_X1 U16461 ( .A1(n14603), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n17539), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n14586) );
  AOI22_X1 U16462 ( .A1(n10958), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n10967), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n14585) );
  AOI22_X1 U16463 ( .A1(n10961), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n10976), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n14584) );
  AOI22_X1 U16464 ( .A1(n17546), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17286), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n14583) );
  NAND4_X1 U16465 ( .A1(n14586), .A2(n14585), .A3(n14584), .A4(n14583), .ZN(
        n14587) );
  AOI22_X1 U16466 ( .A1(n17546), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n14603), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n14593) );
  AOI22_X1 U16467 ( .A1(n10967), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n10966), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n14592) );
  AOI22_X1 U16468 ( .A1(n10968), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n14589), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n14591) );
  AOI22_X1 U16469 ( .A1(n17540), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n20216), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n14590) );
  NAND4_X1 U16470 ( .A1(n14593), .A2(n14592), .A3(n14591), .A4(n14590), .ZN(
        n14600) );
  AOI22_X1 U16471 ( .A1(n10961), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n10965), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n14598) );
  AOI22_X1 U16472 ( .A1(n17538), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n17286), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n14597) );
  AOI22_X1 U16473 ( .A1(n10959), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n10977), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n14596) );
  AOI22_X1 U16474 ( .A1(n17205), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17539), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n14595) );
  NAND4_X1 U16475 ( .A1(n14598), .A2(n14597), .A3(n14596), .A4(n14595), .ZN(
        n14599) );
  AOI22_X1 U16476 ( .A1(n17205), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n10961), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n14611) );
  AOI22_X1 U16477 ( .A1(n17545), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17539), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n14610) );
  AOI22_X1 U16478 ( .A1(n10966), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n10965), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n14602) );
  OAI21_X1 U16479 ( .B1(n17208), .B2(n17453), .A(n14602), .ZN(n14609) );
  AOI22_X1 U16480 ( .A1(n17546), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17286), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n14608) );
  AOI22_X1 U16481 ( .A1(n14604), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n14603), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n14607) );
  AOI22_X1 U16482 ( .A1(n10968), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17540), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n14606) );
  AOI22_X1 U16483 ( .A1(n14589), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n20216), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n14605) );
  NAND3_X1 U16484 ( .A1(n14666), .A2(n14661), .A3(n20809), .ZN(n17148) );
  NAND3_X1 U16485 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n20844) );
  NAND2_X1 U16486 ( .A1(n19013), .A2(n20171), .ZN(n14629) );
  INV_X1 U16487 ( .A(n14666), .ZN(n14621) );
  NAND3_X1 U16488 ( .A1(n14614), .A2(n14662), .A3(n14613), .ZN(n14620) );
  NAND2_X1 U16489 ( .A1(n14616), .A2(n14615), .ZN(n14618) );
  NAND2_X1 U16490 ( .A1(n18925), .A2(n18844), .ZN(n14672) );
  NOR2_X1 U16491 ( .A1(n14622), .A2(n14672), .ZN(n14617) );
  INV_X1 U16492 ( .A(n18844), .ZN(n14623) );
  NAND2_X1 U16493 ( .A1(n20711), .A2(n19013), .ZN(n14632) );
  NAND2_X1 U16494 ( .A1(n20673), .A2(n14622), .ZN(n14658) );
  NAND2_X1 U16495 ( .A1(n14624), .A2(n14678), .ZN(n14667) );
  AND2_X1 U16496 ( .A1(n20711), .A2(n20609), .ZN(n14626) );
  INV_X1 U16497 ( .A(n14679), .ZN(n14635) );
  NOR2_X1 U16498 ( .A1(n14680), .A2(n14666), .ZN(n20806) );
  NAND2_X1 U16499 ( .A1(n18925), .A2(n14629), .ZN(n14664) );
  AOI21_X1 U16500 ( .B1(n20711), .B2(n14658), .A(n18844), .ZN(n14630) );
  AOI21_X1 U16501 ( .B1(n14658), .B2(n14664), .A(n14630), .ZN(n14634) );
  NOR2_X1 U16502 ( .A1(n20687), .A2(n20795), .ZN(n20616) );
  NOR3_X1 U16503 ( .A1(n19013), .A2(n20616), .A3(n20171), .ZN(n14663) );
  AOI211_X1 U16504 ( .C1(n18885), .C2(n14632), .A(n14663), .B(n14631), .ZN(
        n14633) );
  NAND2_X1 U16505 ( .A1(n14634), .A2(n14633), .ZN(n20828) );
  NOR2_X1 U16506 ( .A1(n21006), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n21173) );
  AOI221_X1 U16507 ( .B1(n20885), .B2(n21256), .C1(n20844), .C2(n21256), .A(
        n21173), .ZN(n20925) );
  NOR2_X1 U16508 ( .A1(n20894), .A2(n20882), .ZN(n20897) );
  INV_X1 U16509 ( .A(n20897), .ZN(n14781) );
  NOR2_X2 U16510 ( .A1(n14679), .A2(n20828), .ZN(n20807) );
  INV_X1 U16511 ( .A(n14678), .ZN(n14636) );
  NAND2_X1 U16512 ( .A1(n20807), .A2(n14636), .ZN(n20836) );
  NAND2_X1 U16513 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n21262), .ZN(
        n14646) );
  AOI22_X1 U16514 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B1(n18692), .B2(n20822), .ZN(
        n14643) );
  OAI21_X1 U16515 ( .B1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n20822), .A(
        n14639), .ZN(n14640) );
  OAI22_X1 U16516 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n16711), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n14640), .ZN(n14647) );
  NOR2_X1 U16517 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n16711), .ZN(
        n14641) );
  NAND2_X1 U16518 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n14640), .ZN(
        n14648) );
  AOI22_X1 U16519 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n14647), .B1(
        n14641), .B2(n14648), .ZN(n14652) );
  OAI21_X1 U16520 ( .B1(n14644), .B2(n14643), .A(n14652), .ZN(n14642) );
  AOI21_X1 U16521 ( .B1(n14644), .B2(n14643), .A(n14642), .ZN(n14645) );
  OAI21_X1 U16522 ( .B1(n21262), .B2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n14646), .ZN(n14657) );
  XNOR2_X1 U16523 ( .A(n14646), .B(n14651), .ZN(n14650) );
  AOI21_X1 U16524 ( .B1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n14648), .A(
        n14647), .ZN(n14649) );
  OAI21_X1 U16525 ( .B1(n14654), .B2(n14657), .A(n21250), .ZN(n17566) );
  INV_X1 U16526 ( .A(n17566), .ZN(n21252) );
  NAND2_X1 U16527 ( .A1(n21252), .A2(n20171), .ZN(n14659) );
  INV_X1 U16528 ( .A(n14651), .ZN(n14653) );
  NAND2_X1 U16529 ( .A1(n14653), .A2(n14652), .ZN(n14656) );
  OAI22_X1 U16530 ( .A1(n20674), .A2(n14659), .B1(n21255), .B2(n14658), .ZN(
        n14675) );
  INV_X2 U16531 ( .A(n21710), .ZN(n21756) );
  NAND2_X1 U16532 ( .A1(P3_STATE_REG_2__SCAN_IN), .A2(n21706), .ZN(n21753) );
  AOI21_X1 U16533 ( .B1(n21756), .B2(n21753), .A(n18071), .ZN(n20164) );
  XOR2_X1 U16534 ( .A(n18925), .B(n14680), .Z(n14660) );
  NAND2_X1 U16535 ( .A1(READY2), .A2(READY22_REG_SCAN_IN), .ZN(n21755) );
  OAI21_X1 U16536 ( .B1(n20164), .B2(n14660), .A(n21755), .ZN(n21279) );
  NOR3_X1 U16537 ( .A1(n14661), .A2(n21280), .A3(n21279), .ZN(n14674) );
  INV_X1 U16538 ( .A(n14662), .ZN(n14673) );
  INV_X1 U16539 ( .A(n14663), .ZN(n14671) );
  INV_X1 U16540 ( .A(n14664), .ZN(n14665) );
  OAI211_X1 U16541 ( .C1(n20795), .C2(n18844), .A(n14666), .B(n14665), .ZN(
        n14668) );
  OAI21_X1 U16542 ( .B1(n14669), .B2(n14668), .A(n14667), .ZN(n14670) );
  OAI211_X1 U16543 ( .C1(n14673), .C2(n14672), .A(n14671), .B(n14670), .ZN(
        n16694) );
  AOI211_X1 U16544 ( .C1(n18925), .C2(n14675), .A(n14674), .B(n16694), .ZN(
        n14676) );
  AOI221_X4 U16545 ( .B1(n18844), .B2(n14676), .C1(n21255), .C2(n14676), .A(
        n21310), .ZN(n21117) );
  AOI221_X1 U16546 ( .B1(n14781), .B2(n21229), .C1(n20844), .C2(n21229), .A(
        n21234), .ZN(n14677) );
  NOR2_X1 U16547 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n21301) );
  NAND2_X1 U16548 ( .A1(n21301), .A2(n21296), .ZN(n17530) );
  OR2_X2 U16549 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n17530), .ZN(n21223) );
  INV_X2 U16550 ( .A(n21223), .ZN(n21238) );
  AOI21_X1 U16551 ( .B1(n20925), .B2(n14677), .A(n21238), .ZN(n20920) );
  NOR2_X1 U16552 ( .A1(n21223), .A2(n20250), .ZN(n14780) );
  INV_X1 U16553 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n20845) );
  AOI22_X1 U16554 ( .A1(n10958), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17546), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n14693) );
  AOI22_X1 U16555 ( .A1(n17505), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n10971), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n14692) );
  AOI22_X1 U16556 ( .A1(n17540), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n14589), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n14683) );
  OAI21_X1 U16557 ( .B1(n14730), .B2(n17453), .A(n14683), .ZN(n14690) );
  AOI22_X1 U16558 ( .A1(n17547), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n10977), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n14688) );
  AOI22_X1 U16559 ( .A1(n10967), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17548), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n14687) );
  AOI22_X1 U16560 ( .A1(n17539), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17537), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n14686) );
  AOI22_X1 U16561 ( .A1(n17538), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n10975), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n14685) );
  NAND4_X1 U16562 ( .A1(n14688), .A2(n14687), .A3(n14686), .A4(n14685), .ZN(
        n14689) );
  AOI211_X1 U16563 ( .C1(n10968), .C2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A(
        n14690), .B(n14689), .ZN(n14691) );
  NAND3_X1 U16564 ( .A1(n14693), .A2(n14692), .A3(n14691), .ZN(n20642) );
  AOI22_X1 U16565 ( .A1(n17546), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n10976), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n14697) );
  AOI22_X1 U16566 ( .A1(n10959), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n10966), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n14696) );
  AOI22_X1 U16567 ( .A1(n10968), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17540), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n14695) );
  AOI22_X1 U16568 ( .A1(n14589), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n20216), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n14694) );
  NAND4_X1 U16569 ( .A1(n14697), .A2(n14696), .A3(n14695), .A4(n14694), .ZN(
        n14703) );
  AOI22_X1 U16570 ( .A1(n10972), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n17537), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n14701) );
  AOI22_X1 U16571 ( .A1(n10961), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17548), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n14700) );
  AOI22_X1 U16572 ( .A1(n10967), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n17539), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n14699) );
  INV_X2 U16573 ( .A(n11012), .ZN(n17547) );
  AOI22_X1 U16574 ( .A1(n17547), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17545), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n14698) );
  NAND4_X1 U16575 ( .A1(n14701), .A2(n14700), .A3(n14699), .A4(n14698), .ZN(
        n14702) );
  AOI22_X1 U16576 ( .A1(n17538), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n10971), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n14707) );
  AOI22_X1 U16577 ( .A1(n17547), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n10967), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n14706) );
  AOI22_X1 U16578 ( .A1(n17540), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n14589), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n14705) );
  AOI22_X1 U16579 ( .A1(n10968), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n20216), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n14704) );
  NAND4_X1 U16580 ( .A1(n14707), .A2(n14706), .A3(n14705), .A4(n14704), .ZN(
        n14713) );
  AOI22_X1 U16581 ( .A1(n17546), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n10975), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n14711) );
  AOI22_X1 U16582 ( .A1(n17505), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17548), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n14710) );
  AOI22_X1 U16583 ( .A1(n10958), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17545), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n14709) );
  AOI22_X1 U16584 ( .A1(n17539), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17537), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n14708) );
  NAND4_X1 U16585 ( .A1(n14711), .A2(n14710), .A3(n14709), .A4(n14708), .ZN(
        n14712) );
  AOI22_X1 U16586 ( .A1(n17546), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17539), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n14720) );
  AOI22_X1 U16587 ( .A1(n10959), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n10966), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n14719) );
  INV_X1 U16588 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17369) );
  AOI22_X1 U16589 ( .A1(n14682), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n14589), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n14714) );
  OAI21_X1 U16590 ( .B1(n14730), .B2(n17369), .A(n14714), .ZN(n14718) );
  AOI22_X1 U16591 ( .A1(n17547), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n10972), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n14717) );
  AOI22_X1 U16592 ( .A1(n17545), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n17548), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n14716) );
  AOI22_X1 U16593 ( .A1(n10975), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n17537), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n14715) );
  AOI22_X1 U16594 ( .A1(n10972), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n10965), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n14728) );
  AOI22_X1 U16595 ( .A1(n10967), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n17539), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n14727) );
  AOI22_X1 U16596 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n14682), .B1(
        P3_INSTQUEUE_REG_4__1__SCAN_IN), .B2(n14681), .ZN(n14721) );
  OAI21_X1 U16597 ( .B1(n17523), .B2(n14730), .A(n14721), .ZN(n14726) );
  AOI22_X1 U16598 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n17537), .B1(
        n10977), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n14725) );
  AOI22_X1 U16599 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n17546), .B1(
        P3_INSTQUEUE_REG_5__1__SCAN_IN), .B2(n14603), .ZN(n14724) );
  AOI22_X1 U16600 ( .A1(n10961), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n10966), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n14723) );
  AOI22_X1 U16601 ( .A1(n17547), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n10959), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n14722) );
  NAND2_X1 U16602 ( .A1(n14761), .A2(n20783), .ZN(n14766) );
  AOI22_X1 U16603 ( .A1(n10959), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17548), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n14739) );
  AOI22_X1 U16604 ( .A1(n17545), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17546), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n14738) );
  INV_X1 U16605 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17380) );
  AOI22_X1 U16606 ( .A1(n17540), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n14589), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n14729) );
  OAI21_X1 U16607 ( .B1(n14730), .B2(n17380), .A(n14729), .ZN(n14736) );
  AOI22_X1 U16608 ( .A1(n17538), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n10967), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n14734) );
  AOI22_X1 U16609 ( .A1(n10971), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17537), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n14733) );
  AOI22_X1 U16610 ( .A1(n17505), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17539), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n14732) );
  AOI22_X1 U16611 ( .A1(n17547), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n10976), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n14731) );
  NAND4_X1 U16612 ( .A1(n14734), .A2(n14733), .A3(n14732), .A4(n14731), .ZN(
        n14735) );
  AOI211_X1 U16613 ( .C1(n10968), .C2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A(
        n14736), .B(n14735), .ZN(n14737) );
  NAND3_X1 U16614 ( .A1(n14739), .A2(n14738), .A3(n14737), .ZN(n20652) );
  NAND2_X1 U16615 ( .A1(n14741), .A2(n20652), .ZN(n14740) );
  XOR2_X1 U16616 ( .A(n20642), .B(n17567), .Z(n17569) );
  XNOR2_X1 U16617 ( .A(n20845), .B(n17569), .ZN(n14760) );
  XOR2_X1 U16618 ( .A(n20646), .B(n14740), .Z(n14756) );
  XOR2_X1 U16619 ( .A(n20652), .B(n14741), .Z(n14742) );
  NAND2_X1 U16620 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n14742), .ZN(
        n14755) );
  INV_X1 U16621 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n20914) );
  XNOR2_X1 U16622 ( .A(n20914), .B(n14742), .ZN(n17927) );
  XOR2_X1 U16623 ( .A(n20661), .B(n14766), .Z(n17938) );
  INV_X1 U16624 ( .A(n14761), .ZN(n20666) );
  XOR2_X1 U16625 ( .A(n20666), .B(n20783), .Z(n14743) );
  OR2_X1 U16626 ( .A1(n20894), .A2(n14743), .ZN(n14754) );
  XNOR2_X1 U16627 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n14743), .ZN(
        n17951) );
  AOI22_X1 U16628 ( .A1(n14603), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17537), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n14747) );
  AOI22_X1 U16629 ( .A1(n17546), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10976), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n14746) );
  AOI22_X1 U16630 ( .A1(n10968), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n14589), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n14745) );
  AOI22_X1 U16631 ( .A1(n17540), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n20216), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n14744) );
  NAND4_X1 U16632 ( .A1(n14747), .A2(n14746), .A3(n14745), .A4(n14744), .ZN(
        n14753) );
  AOI22_X1 U16633 ( .A1(n17547), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n17539), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n14751) );
  AOI22_X1 U16634 ( .A1(n17505), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n10972), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n14750) );
  AOI22_X1 U16635 ( .A1(n17545), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10971), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n14749) );
  AOI22_X1 U16636 ( .A1(n10959), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n10967), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n14748) );
  NAND4_X1 U16637 ( .A1(n14751), .A2(n14750), .A3(n14749), .A4(n14748), .ZN(
        n14752) );
  NOR2_X1 U16638 ( .A1(n14753), .A2(n14752), .ZN(n14767) );
  NOR2_X1 U16639 ( .A1(n14767), .A2(n20881), .ZN(n17965) );
  OAI21_X1 U16640 ( .B1(n20882), .B2(n20783), .A(n17956), .ZN(n17950) );
  NAND2_X1 U16641 ( .A1(n17951), .A2(n17950), .ZN(n17949) );
  INV_X1 U16642 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n20915) );
  NAND2_X1 U16643 ( .A1(n14755), .A2(n17925), .ZN(n14757) );
  NAND2_X1 U16644 ( .A1(n14756), .A2(n14757), .ZN(n14758) );
  XOR2_X1 U16645 ( .A(n14757), .B(n14756), .Z(n17915) );
  NAND2_X1 U16646 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n17915), .ZN(
        n17914) );
  OAI21_X1 U16647 ( .B1(n14760), .B2(n14759), .A(n17570), .ZN(n17904) );
  INV_X1 U16648 ( .A(n14767), .ZN(n20788) );
  NOR2_X1 U16649 ( .A1(n20661), .A2(n14764), .ZN(n14774) );
  NAND2_X1 U16650 ( .A1(n14774), .A2(n20652), .ZN(n14777) );
  XOR2_X1 U16651 ( .A(n20646), .B(n14777), .Z(n14762) );
  NAND2_X1 U16652 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n14762), .ZN(
        n14776) );
  XOR2_X1 U16653 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B(n14762), .Z(
        n17911) );
  XOR2_X1 U16654 ( .A(n20661), .B(n14764), .Z(n14763) );
  NAND2_X1 U16655 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n14763), .ZN(
        n14772) );
  XNOR2_X1 U16656 ( .A(n20915), .B(n14763), .ZN(n17935) );
  OAI21_X1 U16657 ( .B1(n14767), .B2(n14766), .A(n14765), .ZN(n14768) );
  NAND2_X1 U16658 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n14768), .ZN(
        n14771) );
  XOR2_X1 U16659 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n14768), .Z(
        n17947) );
  NOR2_X1 U16660 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n20783), .ZN(
        n14770) );
  NOR2_X1 U16661 ( .A1(n20788), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n17964) );
  INV_X1 U16662 ( .A(n17964), .ZN(n17958) );
  NOR2_X1 U16663 ( .A1(n17959), .A2(n17958), .ZN(n17957) );
  NOR3_X1 U16664 ( .A1(n14770), .A2(n14769), .A3(n17957), .ZN(n17946) );
  NAND2_X1 U16665 ( .A1(n17947), .A2(n17946), .ZN(n17945) );
  NAND2_X1 U16666 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n14773), .ZN(
        n14775) );
  XOR2_X1 U16667 ( .A(n20652), .B(n14774), .Z(n17921) );
  NAND2_X1 U16668 ( .A1(n17922), .A2(n17921), .ZN(n17920) );
  NOR2_X1 U16669 ( .A1(n20646), .A2(n14777), .ZN(n17555) );
  XOR2_X1 U16670 ( .A(n20642), .B(n17555), .Z(n17558) );
  NAND2_X1 U16671 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n14778), .ZN(
        n17559) );
  OAI21_X1 U16672 ( .B1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n14778), .A(
        n17559), .ZN(n17902) );
  OAI22_X1 U16673 ( .A1(n20929), .A2(n17904), .B1(n21048), .B2(n17902), .ZN(
        n14779) );
  AOI211_X1 U16674 ( .C1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .C2(n20920), .A(
        n14780), .B(n14779), .ZN(n14785) );
  INV_X1 U16675 ( .A(n20844), .ZN(n14783) );
  OAI21_X1 U16676 ( .B1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n21237), .A(
        n21229), .ZN(n20880) );
  OAI22_X1 U16677 ( .A1(n20885), .A2(n11276), .B1(n14781), .B2(n20880), .ZN(
        n20923) );
  NAND2_X1 U16678 ( .A1(n21117), .A2(n20923), .ZN(n20913) );
  INV_X1 U16679 ( .A(n20913), .ZN(n14782) );
  NAND3_X1 U16680 ( .A1(n14783), .A2(n20845), .A3(n14782), .ZN(n14784) );
  NAND2_X1 U16681 ( .A1(n14785), .A2(n14784), .ZN(P3_U2856) );
  OAI222_X1 U16682 ( .A1(n15701), .A2(n14787), .B1(n15703), .B2(n11859), .C1(
        n15711), .C2(n14786), .ZN(P1_U2897) );
  OAI222_X1 U16683 ( .A1(n15701), .A2(n15652), .B1(n15711), .B2(n14788), .C1(
        n19871), .C2(n15703), .ZN(P1_U2896) );
  INV_X1 U16684 ( .A(n14789), .ZN(n14790) );
  XNOR2_X1 U16685 ( .A(n14791), .B(n14790), .ZN(n18285) );
  INV_X1 U16686 ( .A(n18285), .ZN(n14792) );
  OAI222_X1 U16687 ( .A1(n19403), .A2(n14793), .B1(n19401), .B2(n17129), .C1(
        n19410), .C2(n14792), .ZN(P2_U2904) );
  INV_X1 U16688 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n18280) );
  INV_X1 U16689 ( .A(n14794), .ZN(n14797) );
  INV_X1 U16690 ( .A(n14795), .ZN(n14796) );
  OAI211_X1 U16691 ( .C1(n14797), .C2(n14796), .A(n16141), .B(n14940), .ZN(
        n14804) );
  INV_X1 U16692 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n16531) );
  AOI22_X1 U16693 ( .A1(n15227), .A2(P2_EBX_REG_15__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), 
        .ZN(n14799) );
  NAND2_X1 U16694 ( .A1(n15440), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n14798) );
  OAI211_X1 U16695 ( .C1(n15443), .C2(n16531), .A(n14799), .B(n14798), .ZN(
        n14800) );
  OR2_X1 U16696 ( .A1(n14801), .A2(n14800), .ZN(n14802) );
  AND2_X1 U16697 ( .A1(n14946), .A2(n14802), .ZN(n18286) );
  NAND2_X1 U16698 ( .A1(n18286), .A2(n16102), .ZN(n14803) );
  OAI211_X1 U16699 ( .C1(n16102), .C2(n18280), .A(n14804), .B(n14803), .ZN(
        P2_U2872) );
  NOR2_X2 U16700 ( .A1(n14821), .A2(n14806), .ZN(n15111) );
  AOI22_X1 U16701 ( .A1(n15112), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n15111), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n14815) );
  AOI22_X1 U16702 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19204), .B1(
        n14960), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n14814) );
  AOI22_X1 U16703 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19235), .B1(
        n14967), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n14813) );
  INV_X1 U16704 ( .A(n14819), .ZN(n14809) );
  NOR2_X2 U16705 ( .A1(n14821), .A2(n14809), .ZN(n14966) );
  AOI22_X1 U16706 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n14966), .B1(
        n19214), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n14812) );
  AOI22_X1 U16707 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19310), .B1(
        n19301), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n14827) );
  AOI22_X1 U16708 ( .A1(n14968), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n16673), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n14826) );
  AOI22_X1 U16709 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19324), .B1(
        n14970), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n14825) );
  INV_X1 U16710 ( .A(n14822), .ZN(n14820) );
  NOR2_X2 U16711 ( .A1(n14821), .A2(n14820), .ZN(n14969) );
  AOI22_X1 U16712 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n14969), .B1(
        n14961), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n14824) );
  NAND2_X1 U16713 ( .A1(n14829), .A2(n14828), .ZN(n14830) );
  NAND2_X1 U16714 ( .A1(n14830), .A2(n18090), .ZN(n14833) );
  NAND2_X1 U16715 ( .A1(n14831), .A2(n19605), .ZN(n14832) );
  AOI22_X1 U16716 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19214), .B1(
        n14968), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n14837) );
  AOI22_X1 U16717 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19301), .B1(
        n14970), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n14836) );
  AOI22_X1 U16718 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19310), .B1(
        n15111), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n14835) );
  AOI22_X1 U16719 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19204), .B1(
        n14961), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n14834) );
  INV_X1 U16720 ( .A(n14960), .ZN(n14839) );
  INV_X1 U16721 ( .A(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n14838) );
  INV_X1 U16722 ( .A(n19324), .ZN(n19335) );
  INV_X1 U16723 ( .A(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n14840) );
  NOR2_X1 U16724 ( .A1(n14842), .A2(n14841), .ZN(n14847) );
  AOI22_X1 U16725 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n14969), .B1(
        n14966), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n14844) );
  AOI22_X1 U16726 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n15112), .B1(
        n14967), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n14843) );
  AND2_X1 U16727 ( .A1(n14844), .A2(n14843), .ZN(n14846) );
  NAND4_X1 U16728 ( .A1(n14848), .A2(n14847), .A3(n14846), .A4(n14845), .ZN(
        n14852) );
  NAND2_X1 U16729 ( .A1(n14850), .A2(n14849), .ZN(n14851) );
  NAND2_X1 U16730 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n14854), .ZN(
        n14855) );
  NAND2_X1 U16731 ( .A1(n14856), .A2(n14855), .ZN(n14894) );
  XNOR2_X1 U16732 ( .A(n14894), .B(n18602), .ZN(n14892) );
  XNOR2_X1 U16733 ( .A(n14893), .B(n14892), .ZN(n18590) );
  NAND2_X1 U16734 ( .A1(n14893), .A2(n15139), .ZN(n14860) );
  MUX2_X1 U16735 ( .A(n14857), .B(n16034), .S(n16684), .Z(n14858) );
  OAI21_X1 U16736 ( .B1(n14859), .B2(n14858), .A(n15015), .ZN(n16030) );
  NAND2_X1 U16737 ( .A1(n14860), .A2(n16030), .ZN(n15023) );
  XNOR2_X1 U16738 ( .A(n15023), .B(n18602), .ZN(n14888) );
  INV_X1 U16739 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18626) );
  NOR2_X1 U16740 ( .A1(n16040), .A2(n18626), .ZN(n14861) );
  AOI21_X1 U16741 ( .B1(n14863), .B2(n14862), .A(n14861), .ZN(n15021) );
  XNOR2_X1 U16742 ( .A(n14888), .B(n15021), .ZN(n18599) );
  NAND2_X1 U16743 ( .A1(n18599), .A2(n17039), .ZN(n14869) );
  INV_X1 U16744 ( .A(n13704), .ZN(n14864) );
  INV_X1 U16745 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n16027) );
  NAND2_X1 U16746 ( .A1(n18572), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n18593) );
  OAI21_X1 U16747 ( .B1(n17022), .B2(n16027), .A(n18593), .ZN(n14867) );
  OAI21_X1 U16748 ( .B1(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n14865), .A(
        n14900), .ZN(n18135) );
  NOR2_X1 U16749 ( .A1(n17046), .A2(n18135), .ZN(n14866) );
  AOI211_X1 U16750 ( .C1(n14864), .C2(n17019), .A(n14867), .B(n14866), .ZN(
        n14868) );
  OAI211_X1 U16751 ( .C1(n18590), .C2(n17042), .A(n14869), .B(n14868), .ZN(
        P2_U3011) );
  NOR2_X1 U16752 ( .A1(n11048), .A2(n14870), .ZN(n14871) );
  NOR2_X1 U16753 ( .A1(n14871), .A2(n10984), .ZN(n21484) );
  INV_X1 U16754 ( .A(n21484), .ZN(n14875) );
  AOI21_X1 U16755 ( .B1(n14873), .B2(n14872), .A(n14953), .ZN(n21482) );
  AOI22_X1 U16756 ( .A1(n21482), .A2(n19961), .B1(P1_EBX_REG_9__SCAN_IN), .B2(
        n15617), .ZN(n14874) );
  OAI21_X1 U16757 ( .B1(n14875), .B2(n15628), .A(n14874), .ZN(P1_U2863) );
  OAI222_X1 U16758 ( .A1(n14875), .A2(n15711), .B1(n15703), .B2(n19873), .C1(
        n15647), .C2(n15701), .ZN(P1_U2895) );
  XOR2_X1 U16759 ( .A(n14877), .B(n14876), .Z(n19984) );
  INV_X1 U16760 ( .A(n19984), .ZN(n14887) );
  NAND2_X1 U16761 ( .A1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n14878), .ZN(
        n14929) );
  NOR2_X1 U16762 ( .A1(n14879), .A2(n14929), .ZN(n14928) );
  INV_X1 U16763 ( .A(n14880), .ZN(n14881) );
  AOI22_X1 U16764 ( .A1(n21351), .A2(n15982), .B1(n14928), .B2(n14881), .ZN(
        n14914) );
  INV_X1 U16765 ( .A(n14928), .ZN(n14882) );
  NOR2_X1 U16766 ( .A1(n14933), .A2(n14882), .ZN(n14910) );
  NAND2_X1 U16767 ( .A1(n14910), .A2(n14883), .ZN(n14884) );
  NAND2_X1 U16768 ( .A1(n10970), .A2(P1_REIP_REG_7__SCAN_IN), .ZN(n19985) );
  OAI211_X1 U16769 ( .C1(n21352), .C2(n21468), .A(n14884), .B(n19985), .ZN(
        n14885) );
  AOI21_X1 U16770 ( .B1(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n14914), .A(
        n14885), .ZN(n14886) );
  OAI21_X1 U16771 ( .B1(n14887), .B2(n21353), .A(n14886), .ZN(P1_U3024) );
  INV_X1 U16772 ( .A(n15021), .ZN(n15026) );
  AOI22_X1 U16773 ( .A1(n14888), .A2(n15026), .B1(
        P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n15023), .ZN(n14891) );
  INV_X1 U16774 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n18125) );
  MUX2_X1 U16775 ( .A(n14889), .B(n18125), .S(n16684), .Z(n15014) );
  XNOR2_X1 U16776 ( .A(n15014), .B(n15015), .ZN(n18126) );
  XNOR2_X1 U16777 ( .A(n18126), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n14890) );
  XNOR2_X1 U16778 ( .A(n14891), .B(n14890), .ZN(n18584) );
  NAND2_X1 U16779 ( .A1(n14893), .A2(n14892), .ZN(n14896) );
  NAND2_X1 U16780 ( .A1(n14894), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n14895) );
  NAND2_X1 U16781 ( .A1(n14896), .A2(n14895), .ZN(n14987) );
  XNOR2_X1 U16782 ( .A(n14959), .B(n14958), .ZN(n14988) );
  XNOR2_X1 U16783 ( .A(n14987), .B(n14988), .ZN(n14898) );
  INV_X1 U16784 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n15038) );
  OR2_X1 U16785 ( .A1(n14898), .A2(n15038), .ZN(n14899) );
  NAND2_X1 U16786 ( .A1(n14898), .A2(n15038), .ZN(n14991) );
  AND2_X1 U16787 ( .A1(n14899), .A2(n14991), .ZN(n18583) );
  NOR2_X1 U16788 ( .A1(n18583), .A2(n17042), .ZN(n14904) );
  NOR2_X1 U16789 ( .A1(n18581), .A2(n17062), .ZN(n14903) );
  INV_X2 U16790 ( .A(n18572), .ZN(n18589) );
  OAI22_X1 U16791 ( .A1(n18124), .A2(n17022), .B1(n13825), .B2(n18589), .ZN(
        n14902) );
  AOI21_X1 U16792 ( .B1(n18124), .B2(n14900), .A(n16979), .ZN(n18147) );
  AND2_X1 U16793 ( .A1(n17055), .A2(n18147), .ZN(n14901) );
  NOR4_X1 U16794 ( .A1(n14904), .A2(n14903), .A3(n14902), .A4(n14901), .ZN(
        n14905) );
  OAI21_X1 U16795 ( .B1(n18584), .B2(n17058), .A(n14905), .ZN(P2_U3010) );
  XOR2_X1 U16796 ( .A(n14907), .B(n14906), .Z(n14921) );
  OAI22_X1 U16797 ( .A1(n21352), .A2(n14908), .B1(n19895), .B2(n21386), .ZN(
        n14913) );
  NAND2_X1 U16798 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n14909) );
  OAI211_X1 U16799 ( .C1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A(n14910), .B(n14909), .ZN(n14911) );
  INV_X1 U16800 ( .A(n14911), .ZN(n14912) );
  AOI211_X1 U16801 ( .C1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .C2(n14914), .A(
        n14913), .B(n14912), .ZN(n14915) );
  OAI21_X1 U16802 ( .B1(n14921), .B2(n21353), .A(n14915), .ZN(P1_U3023) );
  AOI22_X1 U16803 ( .A1(n20022), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B1(
        n10970), .B2(P1_REIP_REG_8__SCAN_IN), .ZN(n14916) );
  OAI21_X1 U16804 ( .B1(n20028), .B2(n14917), .A(n14916), .ZN(n14918) );
  AOI21_X1 U16805 ( .B1(n14919), .B2(n20009), .A(n14918), .ZN(n14920) );
  OAI21_X1 U16806 ( .B1(n14921), .B2(n21655), .A(n14920), .ZN(P1_U2991) );
  OAI21_X1 U16807 ( .B1(n14923), .B2(n14922), .A(n15996), .ZN(n14938) );
  INV_X1 U16808 ( .A(n21478), .ZN(n14925) );
  AND2_X1 U16809 ( .A1(n10970), .A2(P1_REIP_REG_9__SCAN_IN), .ZN(n14935) );
  AOI21_X1 U16810 ( .B1(n20022), .B2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .A(
        n14935), .ZN(n14924) );
  OAI21_X1 U16811 ( .B1(n20028), .B2(n14925), .A(n14924), .ZN(n14926) );
  AOI21_X1 U16812 ( .B1(n21484), .B2(n20009), .A(n14926), .ZN(n14927) );
  OAI21_X1 U16813 ( .B1(n14938), .B2(n21655), .A(n14927), .ZN(P1_U2990) );
  NAND3_X1 U16814 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(n14928), .ZN(n15811) );
  INV_X1 U16815 ( .A(n14929), .ZN(n14931) );
  NAND4_X1 U16816 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(n14931), .A4(n14930), .ZN(
        n15807) );
  AOI22_X1 U16817 ( .A1(n15987), .A2(n15811), .B1(n15938), .B2(n15807), .ZN(
        n14932) );
  NAND2_X1 U16818 ( .A1(n15982), .A2(n14932), .ZN(n16003) );
  NOR2_X1 U16819 ( .A1(n14933), .A2(n15811), .ZN(n16001) );
  AOI22_X1 U16820 ( .A1(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n16003), .B1(
        n16001), .B2(n14934), .ZN(n14937) );
  AOI21_X1 U16821 ( .B1(n21409), .B2(n21482), .A(n14935), .ZN(n14936) );
  OAI211_X1 U16822 ( .C1(n14938), .C2(n21353), .A(n14937), .B(n14936), .ZN(
        P1_U3022) );
  NAND2_X1 U16823 ( .A1(n14940), .A2(n14939), .ZN(n14941) );
  NAND2_X1 U16824 ( .A1(n15055), .A2(n14941), .ZN(n19660) );
  INV_X1 U16825 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n14944) );
  NAND2_X1 U16826 ( .A1(n15227), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n14943) );
  NAND2_X1 U16827 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n14942) );
  OAI211_X1 U16828 ( .C1(n10963), .C2(n14944), .A(n14943), .B(n14942), .ZN(
        n14945) );
  AOI21_X1 U16829 ( .B1(n13924), .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n14945), .ZN(n14947) );
  NAND2_X1 U16830 ( .A1(n14946), .A2(n14947), .ZN(n14948) );
  NAND2_X1 U16831 ( .A1(n15070), .A2(n14948), .ZN(n18301) );
  NOR2_X1 U16832 ( .A1(n18301), .A2(n16157), .ZN(n14949) );
  AOI21_X1 U16833 ( .B1(P2_EBX_REG_16__SCAN_IN), .B2(n16157), .A(n14949), .ZN(
        n14950) );
  OAI21_X1 U16834 ( .B1(n19660), .B2(n16167), .A(n14950), .ZN(P2_U2871) );
  XOR2_X1 U16835 ( .A(n14951), .B(n10984), .Z(n21495) );
  NOR2_X1 U16836 ( .A1(n14953), .A2(n14952), .ZN(n14954) );
  OR2_X1 U16837 ( .A1(n15081), .A2(n14954), .ZN(n21492) );
  OAI22_X1 U16838 ( .A1(n19965), .A2(n21492), .B1(n14955), .B2(n19969), .ZN(
        n14956) );
  AOI21_X1 U16839 ( .B1(n21495), .B2(n19962), .A(n14956), .ZN(n14957) );
  INV_X1 U16840 ( .A(n14957), .ZN(P1_U2862) );
  INV_X1 U16841 ( .A(n14985), .ZN(n14983) );
  AOI22_X1 U16842 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19204), .B1(
        n14960), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n14965) );
  AOI22_X1 U16843 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19310), .B1(
        n19235), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n14964) );
  AOI22_X1 U16844 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n16673), .B1(
        n19301), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n14963) );
  AOI22_X1 U16845 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19324), .B1(
        n14961), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n14962) );
  AOI22_X1 U16846 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n14966), .B1(
        n14967), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n14978) );
  AOI22_X1 U16847 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19214), .B1(
        n14968), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n14977) );
  AOI22_X1 U16848 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n14969), .B1(
        n14970), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n14976) );
  INV_X1 U16849 ( .A(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n19436) );
  INV_X1 U16850 ( .A(n15111), .ZN(n14973) );
  INV_X1 U16851 ( .A(n15112), .ZN(n14972) );
  INV_X1 U16852 ( .A(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n14971) );
  OAI22_X1 U16853 ( .A1(n19436), .A2(n14973), .B1(n14972), .B2(n14971), .ZN(
        n14974) );
  INV_X1 U16854 ( .A(n14974), .ZN(n14975) );
  INV_X1 U16855 ( .A(n15017), .ZN(n14979) );
  NAND2_X1 U16856 ( .A1(n14979), .A2(n19605), .ZN(n14980) );
  INV_X1 U16857 ( .A(n14984), .ZN(n14982) );
  NAND2_X1 U16858 ( .A1(n14983), .A2(n14982), .ZN(n14986) );
  INV_X1 U16859 ( .A(n14987), .ZN(n14989) );
  NAND2_X1 U16860 ( .A1(n14989), .A2(n14988), .ZN(n14990) );
  INV_X1 U16861 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n15265) );
  XNOR2_X1 U16862 ( .A(n15267), .B(n15265), .ZN(n16981) );
  NAND2_X1 U16863 ( .A1(n14999), .A2(n14992), .ZN(n15010) );
  OAI21_X1 U16864 ( .B1(n14995), .B2(n14994), .A(n14993), .ZN(n14996) );
  INV_X1 U16865 ( .A(n14996), .ZN(n14997) );
  NAND2_X1 U16866 ( .A1(n14997), .A2(n15011), .ZN(n15009) );
  NOR2_X1 U16867 ( .A1(n14998), .A2(n19605), .ZN(n15006) );
  NAND2_X1 U16868 ( .A1(n15000), .A2(n21729), .ZN(n15003) );
  OAI211_X1 U16869 ( .C1(n15004), .C2(n15003), .A(n15002), .B(n15001), .ZN(
        n15005) );
  AOI21_X1 U16870 ( .B1(n15007), .B2(n15006), .A(n15005), .ZN(n15008) );
  OAI211_X1 U16871 ( .C1(n15011), .C2(n15010), .A(n15009), .B(n15008), .ZN(
        n15012) );
  INV_X1 U16872 ( .A(n15014), .ZN(n15016) );
  MUX2_X1 U16873 ( .A(n13848), .B(n15017), .S(n15131), .Z(n15018) );
  OAI21_X1 U16874 ( .B1(n15019), .B2(n15018), .A(n15134), .ZN(n18141) );
  XNOR2_X1 U16875 ( .A(n15108), .B(n15265), .ZN(n15107) );
  NOR2_X1 U16876 ( .A1(n18126), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n15024) );
  AOI21_X1 U16877 ( .B1(n15021), .B2(n18602), .A(n15024), .ZN(n15022) );
  NAND2_X1 U16878 ( .A1(n15023), .A2(n15022), .ZN(n15028) );
  NOR2_X1 U16879 ( .A1(n15024), .A2(n18602), .ZN(n15025) );
  AOI22_X1 U16880 ( .A1(n15026), .A2(n15025), .B1(n18126), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n15027) );
  NAND2_X1 U16881 ( .A1(n15028), .A2(n15027), .ZN(n15106) );
  XNOR2_X1 U16882 ( .A(n15107), .B(n15106), .ZN(n16980) );
  NAND2_X1 U16883 ( .A1(n15032), .A2(n15031), .ZN(n15033) );
  NAND2_X1 U16884 ( .A1(n15049), .A2(n15033), .ZN(n16616) );
  NAND2_X1 U16885 ( .A1(n18608), .A2(n16616), .ZN(n18555) );
  INV_X1 U16886 ( .A(n18555), .ZN(n18524) );
  NAND2_X1 U16887 ( .A1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18604) );
  INV_X1 U16888 ( .A(n18604), .ZN(n18613) );
  AOI21_X1 U16889 ( .B1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n18613), .A(
        n16616), .ZN(n15034) );
  NAND2_X1 U16890 ( .A1(n18626), .A2(n18604), .ZN(n18610) );
  NOR2_X1 U16891 ( .A1(n18572), .A2(n15049), .ZN(n18516) );
  INV_X1 U16892 ( .A(n18516), .ZN(n18625) );
  OAI21_X1 U16893 ( .B1(n18608), .B2(n18610), .A(n18625), .ZN(n16618) );
  NOR2_X1 U16894 ( .A1(n15034), .A2(n16618), .ZN(n18601) );
  OAI21_X1 U16895 ( .B1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n18524), .A(
        n18601), .ZN(n18580) );
  INV_X1 U16896 ( .A(n18608), .ZN(n15036) );
  NAND2_X1 U16897 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n18613), .ZN(
        n18609) );
  INV_X1 U16898 ( .A(n18609), .ZN(n15035) );
  OAI211_X1 U16899 ( .C1(n15036), .C2(n15035), .A(n18610), .B(n18555), .ZN(
        n18603) );
  INV_X1 U16900 ( .A(n18603), .ZN(n15037) );
  NAND2_X1 U16901 ( .A1(n15037), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n18582) );
  AOI221_X1 U16902 ( .B1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .C1(n15038), .C2(n15265), .A(
        n18582), .ZN(n15040) );
  NOR2_X1 U16903 ( .A1(n13830), .A2(n18589), .ZN(n15039) );
  AOI211_X1 U16904 ( .C1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .C2(n18580), .A(
        n15040), .B(n15039), .ZN(n15052) );
  OAI21_X1 U16905 ( .B1(n14453), .B2(n15042), .A(n15041), .ZN(n19409) );
  NAND2_X1 U16906 ( .A1(n15043), .A2(n18090), .ZN(n15045) );
  NAND2_X1 U16907 ( .A1(n15045), .A2(n15044), .ZN(n15046) );
  NAND2_X1 U16908 ( .A1(n14012), .A2(n19605), .ZN(n15047) );
  NAND2_X1 U16909 ( .A1(n15047), .A2(n12790), .ZN(n15048) );
  OAI22_X1 U16910 ( .A1(n19409), .A2(n18594), .B1(n18605), .B2(n18149), .ZN(
        n15050) );
  INV_X1 U16911 ( .A(n15050), .ZN(n15051) );
  OAI211_X1 U16912 ( .C1(n16980), .C2(n18606), .A(n15052), .B(n15051), .ZN(
        n15053) );
  INV_X1 U16913 ( .A(n15053), .ZN(n15054) );
  OAI21_X1 U16914 ( .B1(n16981), .B2(n18617), .A(n15054), .ZN(P2_U3041) );
  AOI21_X1 U16915 ( .B1(n15056), .B2(n15055), .A(n16160), .ZN(n15057) );
  INV_X1 U16916 ( .A(n15057), .ZN(n15074) );
  XOR2_X1 U16917 ( .A(n16523), .B(n15058), .Z(n18553) );
  INV_X1 U16918 ( .A(n18553), .ZN(n15060) );
  OAI22_X1 U16919 ( .A1(n19658), .A2(n15060), .B1(n15059), .B2(n19401), .ZN(
        n15061) );
  AOI21_X1 U16920 ( .B1(n19653), .B2(n15062), .A(n15061), .ZN(n15064) );
  AOI22_X1 U16921 ( .A1(n19654), .A2(BUF1_REG_17__SCAN_IN), .B1(n19655), .B2(
        BUF2_REG_17__SCAN_IN), .ZN(n15063) );
  OAI211_X1 U16922 ( .C1(n15074), .C2(n19659), .A(n15064), .B(n15063), .ZN(
        P2_U2902) );
  NAND2_X1 U16923 ( .A1(n16111), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n15073) );
  INV_X1 U16924 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n15067) );
  NAND2_X1 U16925 ( .A1(n15227), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n15066) );
  NAND2_X1 U16926 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n15065) );
  OAI211_X1 U16927 ( .C1(n15436), .C2(n15067), .A(n15066), .B(n15065), .ZN(
        n15068) );
  AOI21_X1 U16928 ( .B1(n13924), .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n15068), .ZN(n15071) );
  INV_X1 U16929 ( .A(n16162), .ZN(n15069) );
  AOI21_X1 U16930 ( .B1(n15071), .B2(n15070), .A(n15069), .ZN(n18554) );
  NAND2_X1 U16931 ( .A1(n18554), .A2(n16102), .ZN(n15072) );
  OAI211_X1 U16932 ( .C1(n15074), .C2(n16167), .A(n15073), .B(n15072), .ZN(
        P2_U2870) );
  INV_X1 U16933 ( .A(n21495), .ZN(n15075) );
  OAI222_X1 U16934 ( .A1(n15701), .A2(n15642), .B1(n15711), .B2(n15075), .C1(
        n19875), .C2(n15703), .ZN(P1_U2894) );
  NAND2_X1 U16935 ( .A1(n15077), .A2(n15076), .ZN(n15078) );
  NAND2_X1 U16936 ( .A1(n15085), .A2(n15078), .ZN(n15084) );
  XNOR2_X1 U16937 ( .A(n15084), .B(n15083), .ZN(n21502) );
  OAI222_X1 U16938 ( .A1(n21502), .A2(n15711), .B1(n15703), .B2(n19877), .C1(
        n15701), .C2(n15079), .ZN(P1_U2893) );
  OAI21_X1 U16939 ( .B1(n15081), .B2(n15080), .A(n15102), .ZN(n21340) );
  INV_X1 U16940 ( .A(P1_EBX_REG_11__SCAN_IN), .ZN(n15082) );
  OAI222_X1 U16941 ( .A1(n19965), .A2(n21340), .B1(n19969), .B2(n15082), .C1(
        n19966), .C2(n21502), .ZN(P1_U2861) );
  OR2_X1 U16942 ( .A1(n15084), .A2(n15083), .ZN(n15086) );
  NAND2_X1 U16943 ( .A1(n15086), .A2(n15085), .ZN(n15094) );
  NAND2_X1 U16944 ( .A1(n15094), .A2(n15095), .ZN(n15098) );
  INV_X1 U16945 ( .A(n15087), .ZN(n15089) );
  AOI21_X1 U16946 ( .B1(n15098), .B2(n15089), .A(n15088), .ZN(n15804) );
  INV_X1 U16947 ( .A(n15804), .ZN(n21528) );
  AOI22_X1 U16948 ( .A1(n15709), .A2(n15507), .B1(P1_EAX_REG_13__SCAN_IN), 
        .B2(n15707), .ZN(n15090) );
  OAI21_X1 U16949 ( .B1(n21528), .B2(n15711), .A(n15090), .ZN(P1_U2891) );
  NAND2_X1 U16950 ( .A1(n15104), .A2(n15091), .ZN(n15092) );
  AND2_X1 U16951 ( .A1(n15974), .A2(n15092), .ZN(n21520) );
  AOI22_X1 U16952 ( .A1(n21520), .A2(n19961), .B1(n15617), .B2(
        P1_EBX_REG_13__SCAN_IN), .ZN(n15093) );
  OAI21_X1 U16953 ( .B1(n21528), .B2(n15628), .A(n15093), .ZN(P1_U2859) );
  INV_X1 U16954 ( .A(n15094), .ZN(n15097) );
  INV_X1 U16955 ( .A(n15095), .ZN(n15096) );
  NAND2_X1 U16956 ( .A1(n15097), .A2(n15096), .ZN(n15099) );
  AOI22_X1 U16957 ( .A1(n15709), .A2(n15633), .B1(P1_EAX_REG_12__SCAN_IN), 
        .B2(n15707), .ZN(n15100) );
  OAI21_X1 U16958 ( .B1(n21519), .B2(n15711), .A(n15100), .ZN(P1_U2892) );
  NAND2_X1 U16959 ( .A1(n15102), .A2(n15101), .ZN(n15103) );
  NAND2_X1 U16960 ( .A1(n15104), .A2(n15103), .ZN(n21512) );
  OAI222_X1 U16961 ( .A1(n21519), .A2(n19966), .B1(n19969), .B2(n15105), .C1(
        n21512), .C2(n19965), .ZN(P1_U2860) );
  NAND2_X1 U16962 ( .A1(n15107), .A2(n15106), .ZN(n15110) );
  NAND2_X1 U16963 ( .A1(n15108), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n15109) );
  AOI22_X1 U16964 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n15111), .B1(
        n15112), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n15116) );
  AOI22_X1 U16965 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19204), .B1(
        n14960), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n15115) );
  AOI22_X1 U16966 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n14967), .B1(
        n19235), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n15114) );
  AOI22_X1 U16967 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n14966), .B1(
        n19214), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n15113) );
  NAND4_X1 U16968 ( .A1(n15116), .A2(n15115), .A3(n15114), .A4(n15113), .ZN(
        n15126) );
  AOI22_X1 U16969 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19301), .B1(
        n19310), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n15124) );
  AOI22_X1 U16970 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n14961), .B1(
        n14969), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n15123) );
  AOI22_X1 U16971 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n14970), .B1(
        n19324), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n15122) );
  INV_X1 U16972 ( .A(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n19400) );
  INV_X1 U16973 ( .A(n16673), .ZN(n15117) );
  INV_X1 U16974 ( .A(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n15118) );
  OAI22_X1 U16975 ( .A1(n19400), .A2(n15117), .B1(n15119), .B2(n15118), .ZN(
        n15120) );
  INV_X1 U16976 ( .A(n15120), .ZN(n15121) );
  NAND4_X1 U16977 ( .A1(n15124), .A2(n15123), .A3(n15122), .A4(n15121), .ZN(
        n15125) );
  NAND2_X1 U16978 ( .A1(n15132), .A2(n19605), .ZN(n15127) );
  MUX2_X1 U16979 ( .A(P2_EBX_REG_6__SCAN_IN), .B(n15132), .S(n15131), .Z(
        n15133) );
  INV_X1 U16980 ( .A(n15143), .ZN(n15136) );
  NAND2_X1 U16981 ( .A1(n15134), .A2(n15133), .ZN(n15135) );
  NAND2_X1 U16982 ( .A1(n15136), .A2(n15135), .ZN(n18155) );
  INV_X1 U16983 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n15243) );
  NAND2_X1 U16984 ( .A1(n15137), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n15138) );
  MUX2_X1 U16985 ( .A(n18171), .B(n15420), .S(n15131), .Z(n15142) );
  INV_X1 U16986 ( .A(P2_EBX_REG_8__SCAN_IN), .ZN(n18183) );
  NOR2_X1 U16987 ( .A1(n15131), .A2(n18183), .ZN(n15140) );
  NAND2_X1 U16988 ( .A1(n15419), .A2(n15140), .ZN(n15141) );
  NAND2_X1 U16989 ( .A1(n15151), .A2(n15141), .ZN(n18181) );
  NOR2_X1 U16990 ( .A1(n18181), .A2(n15139), .ZN(n15146) );
  NAND2_X1 U16991 ( .A1(n15146), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n16989) );
  OR2_X1 U16992 ( .A1(n15143), .A2(n15142), .ZN(n15144) );
  NAND2_X1 U16993 ( .A1(n15419), .A2(n15144), .ZN(n18174) );
  INV_X1 U16994 ( .A(n18174), .ZN(n15145) );
  NAND2_X1 U16995 ( .A1(n15145), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16990) );
  NAND2_X1 U16996 ( .A1(n16989), .A2(n16990), .ZN(n15150) );
  INV_X1 U16997 ( .A(n15146), .ZN(n15148) );
  INV_X1 U16998 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n15147) );
  NAND2_X1 U16999 ( .A1(n15148), .A2(n15147), .ZN(n16988) );
  NAND2_X1 U17000 ( .A1(n18174), .A2(n16623), .ZN(n16992) );
  AND2_X1 U17001 ( .A1(n16988), .A2(n16992), .ZN(n15149) );
  XNOR2_X1 U17002 ( .A(n15151), .B(n11067), .ZN(n18196) );
  AOI21_X1 U17003 ( .B1(n18196), .B2(n15420), .A(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n16609) );
  NAND2_X1 U17004 ( .A1(n16684), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n15152) );
  OR2_X1 U17005 ( .A1(n15153), .A2(n15152), .ZN(n15154) );
  AND2_X1 U17006 ( .A1(n15154), .A2(n15161), .ZN(n18209) );
  NAND2_X1 U17007 ( .A1(n18209), .A2(n15420), .ZN(n15155) );
  INV_X1 U17008 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16583) );
  NAND2_X1 U17009 ( .A1(n15155), .A2(n16583), .ZN(n16586) );
  INV_X1 U17010 ( .A(n15155), .ZN(n15156) );
  NAND2_X1 U17011 ( .A1(n15156), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n16587) );
  AND2_X1 U17012 ( .A1(n15420), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n15157) );
  NAND2_X1 U17013 ( .A1(n18196), .A2(n15157), .ZN(n16584) );
  AND2_X1 U17014 ( .A1(n16587), .A2(n16584), .ZN(n15158) );
  NOR2_X1 U17015 ( .A1(n15131), .A2(n18225), .ZN(n15160) );
  INV_X1 U17016 ( .A(n15160), .ZN(n15159) );
  XNOR2_X1 U17017 ( .A(n15161), .B(n15159), .ZN(n18224) );
  NAND2_X1 U17018 ( .A1(n18224), .A2(n15420), .ZN(n16569) );
  INV_X1 U17019 ( .A(P2_EBX_REG_12__SCAN_IN), .ZN(n18237) );
  NOR2_X1 U17020 ( .A1(n15131), .A2(n18237), .ZN(n15162) );
  AND2_X1 U17021 ( .A1(n15163), .A2(n15162), .ZN(n15164) );
  OR2_X1 U17022 ( .A1(n15164), .A2(n15182), .ZN(n18235) );
  NOR2_X1 U17023 ( .A1(n18235), .A2(n15139), .ZN(n15185) );
  NAND2_X1 U17024 ( .A1(n15185), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n16558) );
  OAI21_X1 U17025 ( .B1(n15249), .B2(n16569), .A(n16558), .ZN(n15165) );
  NAND2_X1 U17026 ( .A1(n16684), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n15181) );
  NAND2_X1 U17027 ( .A1(n16684), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n15187) );
  NOR2_X1 U17028 ( .A1(n15131), .A2(n18280), .ZN(n15177) );
  INV_X1 U17029 ( .A(P2_EBX_REG_16__SCAN_IN), .ZN(n18291) );
  NOR2_X1 U17030 ( .A1(n15131), .A2(n18291), .ZN(n15171) );
  NAND2_X1 U17031 ( .A1(n16684), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n15198) );
  NAND2_X1 U17032 ( .A1(n16684), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n15195) );
  INV_X1 U17033 ( .A(P2_EBX_REG_19__SCAN_IN), .ZN(n18333) );
  NOR2_X1 U17034 ( .A1(n15131), .A2(n18333), .ZN(n15168) );
  INV_X1 U17035 ( .A(P2_EBX_REG_20__SCAN_IN), .ZN(n18351) );
  NOR2_X1 U17036 ( .A1(n15131), .A2(n18351), .ZN(n15218) );
  INV_X1 U17037 ( .A(P2_EBX_REG_21__SCAN_IN), .ZN(n18359) );
  NOR2_X1 U17038 ( .A1(n15131), .A2(n18359), .ZN(n15224) );
  INV_X1 U17039 ( .A(n15224), .ZN(n15166) );
  XNOR2_X1 U17040 ( .A(n15225), .B(n15166), .ZN(n18361) );
  NAND2_X1 U17041 ( .A1(n18361), .A2(n15420), .ZN(n15167) );
  INV_X1 U17042 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n16461) );
  NAND2_X1 U17043 ( .A1(n15167), .A2(n16461), .ZN(n16303) );
  NAND2_X1 U17044 ( .A1(n11030), .A2(n15168), .ZN(n15169) );
  NAND2_X1 U17045 ( .A1(n11010), .A2(n15169), .ZN(n18330) );
  OR2_X1 U17046 ( .A1(n18330), .A2(n15139), .ZN(n15170) );
  INV_X1 U17047 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n16492) );
  NAND2_X1 U17048 ( .A1(n15170), .A2(n16492), .ZN(n16342) );
  AND2_X1 U17049 ( .A1(n15179), .A2(n15171), .ZN(n15172) );
  OR2_X1 U17050 ( .A1(n15172), .A2(n15199), .ZN(n15175) );
  INV_X1 U17051 ( .A(n15175), .ZN(n18293) );
  AND2_X1 U17052 ( .A1(n15420), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15173) );
  NAND2_X1 U17053 ( .A1(n18293), .A2(n15173), .ZN(n16313) );
  INV_X1 U17054 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15174) );
  OAI21_X1 U17055 ( .B1(n15175), .B2(n15139), .A(n15174), .ZN(n15176) );
  NAND2_X1 U17056 ( .A1(n16313), .A2(n15176), .ZN(n16312) );
  NAND2_X1 U17057 ( .A1(n15190), .A2(n15177), .ZN(n15178) );
  NAND2_X1 U17058 ( .A1(n15179), .A2(n15178), .ZN(n18281) );
  OR2_X1 U17059 ( .A1(n18281), .A2(n15139), .ZN(n15180) );
  NAND2_X1 U17060 ( .A1(n15180), .A2(n16531), .ZN(n16380) );
  NOR2_X1 U17061 ( .A1(n15182), .A2(n15181), .ZN(n15183) );
  OR2_X1 U17062 ( .A1(n15188), .A2(n15183), .ZN(n15211) );
  INV_X1 U17063 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15184) );
  OAI21_X1 U17064 ( .B1(n15211), .B2(n15139), .A(n15184), .ZN(n16388) );
  INV_X1 U17065 ( .A(n15185), .ZN(n15186) );
  INV_X1 U17066 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n16563) );
  NAND2_X1 U17067 ( .A1(n15186), .A2(n16563), .ZN(n16557) );
  AND2_X1 U17068 ( .A1(n16388), .A2(n16557), .ZN(n15193) );
  OR2_X1 U17069 ( .A1(n15188), .A2(n15187), .ZN(n15189) );
  AND2_X1 U17070 ( .A1(n15190), .A2(n15189), .ZN(n18269) );
  NAND2_X1 U17071 ( .A1(n18269), .A2(n15420), .ZN(n15192) );
  NAND2_X1 U17072 ( .A1(n15192), .A2(n15191), .ZN(n16378) );
  AND3_X1 U17073 ( .A1(n16380), .A2(n15193), .A3(n16378), .ZN(n16308) );
  NAND2_X1 U17074 ( .A1(n16308), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n15194) );
  NOR2_X1 U17075 ( .A1(n16312), .A2(n15194), .ZN(n15203) );
  OR2_X1 U17076 ( .A1(n15201), .A2(n15195), .ZN(n15196) );
  AND2_X1 U17077 ( .A1(n11030), .A2(n15196), .ZN(n18320) );
  NAND2_X1 U17078 ( .A1(n18320), .A2(n15420), .ZN(n15197) );
  INV_X1 U17079 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n16326) );
  NAND2_X1 U17080 ( .A1(n15197), .A2(n16326), .ZN(n16353) );
  NOR2_X1 U17081 ( .A1(n15199), .A2(n15198), .ZN(n15200) );
  OR2_X1 U17082 ( .A1(n15201), .A2(n15200), .ZN(n18306) );
  INV_X1 U17083 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15202) );
  OAI21_X1 U17084 ( .B1(n18306), .B2(n15139), .A(n15202), .ZN(n16363) );
  AND4_X1 U17085 ( .A1(n16342), .A2(n15203), .A3(n16353), .A4(n16363), .ZN(
        n15204) );
  AND2_X1 U17086 ( .A1(n16303), .A2(n15204), .ZN(n15205) );
  AND2_X1 U17087 ( .A1(n15420), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15206) );
  NAND2_X1 U17088 ( .A1(n18361), .A2(n15206), .ZN(n16302) );
  INV_X1 U17089 ( .A(n18320), .ZN(n15208) );
  NAND2_X1 U17090 ( .A1(n15420), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15207) );
  NAND2_X1 U17091 ( .A1(n15420), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15209) );
  OR2_X1 U17092 ( .A1(n18281), .A2(n15209), .ZN(n16379) );
  AND2_X1 U17093 ( .A1(n15420), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n15210) );
  NAND2_X1 U17094 ( .A1(n18269), .A2(n15210), .ZN(n16377) );
  INV_X1 U17095 ( .A(n15211), .ZN(n18253) );
  AND2_X1 U17096 ( .A1(n15420), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n15212) );
  NAND2_X1 U17097 ( .A1(n18253), .A2(n15212), .ZN(n16387) );
  AND3_X1 U17098 ( .A1(n16379), .A2(n16377), .A3(n16387), .ZN(n16309) );
  NAND2_X1 U17099 ( .A1(n15420), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n15213) );
  OR2_X1 U17100 ( .A1(n18306), .A2(n15213), .ZN(n16362) );
  AND4_X1 U17101 ( .A1(n16352), .A2(n16309), .A3(n16313), .A4(n16362), .ZN(
        n15215) );
  NAND2_X1 U17102 ( .A1(n15420), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15214) );
  NAND3_X1 U17103 ( .A1(n16302), .A2(n15215), .A3(n16341), .ZN(n15216) );
  AOI21_X1 U17104 ( .B1(n15221), .B2(n15217), .A(n15216), .ZN(n15223) );
  INV_X1 U17105 ( .A(n15218), .ZN(n15219) );
  XNOR2_X1 U17106 ( .A(n11010), .B(n15219), .ZN(n18349) );
  INV_X1 U17107 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n16475) );
  NAND2_X1 U17108 ( .A1(n16684), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n15300) );
  NOR2_X2 U17109 ( .A1(n15225), .A2(n15224), .ZN(n15301) );
  XOR2_X1 U17110 ( .A(n15300), .B(n15301), .Z(n18374) );
  NAND2_X1 U17111 ( .A1(n18374), .A2(n15420), .ZN(n15297) );
  INV_X1 U17112 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15298) );
  XNOR2_X1 U17113 ( .A(n15297), .B(n15298), .ZN(n15226) );
  XNOR2_X1 U17114 ( .A(n15299), .B(n15226), .ZN(n15296) );
  INV_X1 U17115 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n16356) );
  NAND2_X1 U17116 ( .A1(n15227), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n15229) );
  NAND2_X1 U17117 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n15228) );
  OAI211_X1 U17118 ( .C1(n15436), .C2(n16356), .A(n15229), .B(n15228), .ZN(
        n15230) );
  AOI21_X1 U17119 ( .B1(n13924), .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n15230), .ZN(n16161) );
  AOI22_X1 U17120 ( .A1(n15227), .A2(P2_EBX_REG_19__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), 
        .ZN(n15232) );
  NAND2_X1 U17121 ( .A1(n15440), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n15231) );
  OAI211_X1 U17122 ( .C1(n15443), .C2(n16492), .A(n15232), .B(n15231), .ZN(
        n16155) );
  INV_X1 U17123 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n18350) );
  NAND2_X1 U17124 ( .A1(n15227), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n15234) );
  NAND2_X1 U17125 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n15233) );
  OAI211_X1 U17126 ( .C1(n15436), .C2(n18350), .A(n15234), .B(n15233), .ZN(
        n15235) );
  AOI21_X1 U17127 ( .B1(n13924), .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n15235), .ZN(n16146) );
  INV_X1 U17128 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n18358) );
  NAND2_X1 U17129 ( .A1(n15227), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n15237) );
  NAND2_X1 U17130 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n15236) );
  OAI211_X1 U17131 ( .C1(n10963), .C2(n18358), .A(n15237), .B(n15236), .ZN(
        n15238) );
  AOI21_X1 U17132 ( .B1(n13924), .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n15238), .ZN(n16136) );
  AOI22_X1 U17133 ( .A1(n15227), .A2(P2_EBX_REG_22__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), 
        .ZN(n15240) );
  NAND2_X1 U17134 ( .A1(n15440), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n15239) );
  OAI211_X1 U17135 ( .C1(n15443), .C2(n15298), .A(n15240), .B(n15239), .ZN(
        n15241) );
  NOR2_X1 U17136 ( .A1(n16137), .A2(n15241), .ZN(n15242) );
  OR2_X1 U17137 ( .A1(n15349), .A2(n15242), .ZN(n16133) );
  INV_X1 U17138 ( .A(n16133), .ZN(n18375) );
  NAND3_X1 U17139 ( .A1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n16630) );
  NOR2_X1 U17140 ( .A1(n15243), .A2(n16630), .ZN(n15245) );
  NAND4_X1 U17141 ( .A1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A3(n15245), .A4(n18610), .ZN(
        n15254) );
  INV_X1 U17142 ( .A(n15254), .ZN(n15244) );
  OAI21_X1 U17143 ( .B1(n18608), .B2(n15244), .A(n18625), .ZN(n16469) );
  INV_X1 U17144 ( .A(n15245), .ZN(n16622) );
  NOR2_X1 U17145 ( .A1(n18609), .A2(n16622), .ZN(n16617) );
  NAND3_X1 U17146 ( .A1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(n16617), .ZN(n15253) );
  INV_X1 U17147 ( .A(n15253), .ZN(n16516) );
  NOR2_X1 U17148 ( .A1(n16616), .A2(n16516), .ZN(n15246) );
  OR2_X1 U17149 ( .A1(n16469), .A2(n15246), .ZN(n16601) );
  AND4_X1 U17150 ( .A1(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A4(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15248) );
  NAND2_X1 U17151 ( .A1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n15259) );
  INV_X1 U17152 ( .A(n15259), .ZN(n15247) );
  INV_X1 U17153 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n16603) );
  NOR3_X1 U17154 ( .A1(n15249), .A2(n16583), .A3(n16603), .ZN(n16547) );
  AND3_X1 U17155 ( .A1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A3(n16547), .ZN(n18548) );
  NAND2_X1 U17156 ( .A1(n11081), .A2(n16532), .ZN(n15250) );
  AND2_X1 U17157 ( .A1(n18555), .A2(n15250), .ZN(n15251) );
  NOR2_X1 U17158 ( .A1(n16601), .A2(n15251), .ZN(n16462) );
  INV_X1 U17159 ( .A(n15352), .ZN(n15252) );
  AOI21_X1 U17160 ( .B1(n11079), .B2(n16228), .A(n15252), .ZN(n19351) );
  NOR2_X1 U17161 ( .A1(n16616), .A2(n15253), .ZN(n15256) );
  NOR2_X1 U17162 ( .A1(n18608), .A2(n15254), .ZN(n15255) );
  AND2_X1 U17163 ( .A1(n16532), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15257) );
  NAND3_X1 U17164 ( .A1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A3(n16514), .ZN(n16473) );
  INV_X1 U17165 ( .A(n16473), .ZN(n15258) );
  NAND2_X1 U17166 ( .A1(n16474), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n16484) );
  NOR2_X1 U17167 ( .A1(n16484), .A2(n15259), .ZN(n15327) );
  INV_X1 U17168 ( .A(n15327), .ZN(n15357) );
  NAND2_X1 U17169 ( .A1(P2_REIP_REG_22__SCAN_IN), .A2(n18572), .ZN(n15260) );
  OAI21_X1 U17170 ( .B1(n15357), .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n15260), .ZN(n15261) );
  AOI21_X1 U17171 ( .B1(n18622), .B2(n19351), .A(n15261), .ZN(n15262) );
  OAI21_X1 U17172 ( .B1(n16462), .B2(n15298), .A(n15262), .ZN(n15263) );
  AOI21_X1 U17173 ( .B1(n18375), .B2(n18591), .A(n15263), .ZN(n15286) );
  AND2_X1 U17174 ( .A1(n15020), .A2(n15265), .ZN(n15264) );
  OR2_X1 U17175 ( .A1(n15266), .A2(n15264), .ZN(n15268) );
  INV_X1 U17176 ( .A(n15020), .ZN(n15270) );
  NAND3_X1 U17177 ( .A1(n15270), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A3(
        n15269), .ZN(n15271) );
  NAND2_X1 U17178 ( .A1(n15273), .A2(n15272), .ZN(n15274) );
  XNOR2_X1 U17179 ( .A(n15280), .B(n15139), .ZN(n15276) );
  XNOR2_X1 U17180 ( .A(n15276), .B(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16396) );
  NAND2_X1 U17181 ( .A1(n16397), .A2(n16396), .ZN(n15279) );
  INV_X1 U17182 ( .A(n15276), .ZN(n15277) );
  NAND2_X1 U17183 ( .A1(n15277), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15278) );
  NAND2_X1 U17184 ( .A1(n15282), .A2(n15420), .ZN(n15281) );
  XNOR2_X1 U17185 ( .A(n15281), .B(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n16996) );
  NAND3_X1 U17186 ( .A1(n15282), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A3(
        n15420), .ZN(n15283) );
  INV_X1 U17187 ( .A(n16327), .ZN(n15284) );
  NAND2_X1 U17188 ( .A1(n15284), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15360) );
  NAND2_X1 U17189 ( .A1(n16327), .A2(n15298), .ZN(n15293) );
  NAND3_X1 U17190 ( .A1(n15360), .A2(n18568), .A3(n15293), .ZN(n15285) );
  OAI211_X1 U17191 ( .C1(n15296), .C2(n18606), .A(n15286), .B(n15285), .ZN(
        P2_U3024) );
  INV_X1 U17192 ( .A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n16367) );
  INV_X1 U17193 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n16325) );
  INV_X1 U17194 ( .A(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n15288) );
  AND2_X1 U17195 ( .A1(n16322), .A2(n15288), .ZN(n15287) );
  OR2_X1 U17196 ( .A1(n15287), .A2(n15364), .ZN(n18377) );
  INV_X1 U17197 ( .A(n18377), .ZN(n15290) );
  INV_X1 U17198 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n18371) );
  OAI22_X1 U17199 ( .A1(n17022), .A2(n15288), .B1(n18371), .B2(n18589), .ZN(
        n15289) );
  AOI21_X1 U17200 ( .B1(n15290), .B2(n17055), .A(n15289), .ZN(n15291) );
  OAI21_X1 U17201 ( .B1(n16133), .B2(n17062), .A(n15291), .ZN(n15292) );
  INV_X1 U17202 ( .A(n15292), .ZN(n15295) );
  NAND3_X1 U17203 ( .A1(n15360), .A2(n17047), .A3(n15293), .ZN(n15294) );
  OAI211_X1 U17204 ( .C1(n15296), .C2(n17058), .A(n15295), .B(n15294), .ZN(
        P2_U2992) );
  NAND2_X1 U17205 ( .A1(n16684), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n15302) );
  NOR2_X1 U17206 ( .A1(n15303), .A2(n15302), .ZN(n15304) );
  OR2_X1 U17207 ( .A1(n15306), .A2(n15304), .ZN(n18385) );
  INV_X1 U17208 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15361) );
  OAI21_X1 U17209 ( .B1(n18385), .B2(n15139), .A(n15361), .ZN(n15343) );
  NOR3_X1 U17210 ( .A1(n18385), .A2(n15139), .A3(n15361), .ZN(n15345) );
  INV_X1 U17211 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15325) );
  NAND2_X1 U17212 ( .A1(n16684), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n15305) );
  XOR2_X1 U17213 ( .A(n15305), .B(n15306), .Z(n18399) );
  NAND2_X1 U17214 ( .A1(n18399), .A2(n15420), .ZN(n15374) );
  INV_X1 U17215 ( .A(P2_EBX_REG_25__SCAN_IN), .ZN(n18411) );
  XNOR2_X1 U17216 ( .A(n15399), .B(n11078), .ZN(n18413) );
  NOR2_X1 U17217 ( .A1(n15307), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n16289) );
  INV_X1 U17218 ( .A(n16289), .ZN(n15309) );
  INV_X1 U17219 ( .A(n15307), .ZN(n15308) );
  INV_X1 U17220 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n16448) );
  NAND2_X1 U17221 ( .A1(n15309), .A2(n16290), .ZN(n15310) );
  XNOR2_X1 U17222 ( .A(n16291), .B(n15310), .ZN(n15341) );
  AOI22_X1 U17223 ( .A1(n15227), .A2(P2_EBX_REG_23__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), 
        .ZN(n15312) );
  NAND2_X1 U17224 ( .A1(n15440), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n15311) );
  OAI211_X1 U17225 ( .C1(n15443), .C2(n15361), .A(n15312), .B(n15311), .ZN(
        n15348) );
  NAND2_X1 U17226 ( .A1(n15349), .A2(n15348), .ZN(n15347) );
  INV_X1 U17227 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n18396) );
  NAND2_X1 U17228 ( .A1(n15227), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n15314) );
  NAND2_X1 U17229 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n15313) );
  OAI211_X1 U17230 ( .C1(n15436), .C2(n18396), .A(n15314), .B(n15313), .ZN(
        n15315) );
  AOI21_X1 U17231 ( .B1(n13924), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n15315), .ZN(n15379) );
  NAND2_X1 U17232 ( .A1(n15227), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n15317) );
  NAND2_X1 U17233 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n15316) );
  OAI211_X1 U17234 ( .C1(n15436), .C2(n18410), .A(n15317), .B(n15316), .ZN(
        n15318) );
  AOI21_X1 U17235 ( .B1(n13924), .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n15318), .ZN(n15319) );
  AND2_X1 U17236 ( .A1(n15377), .A2(n15319), .ZN(n15320) );
  OR2_X1 U17237 ( .A1(n15320), .A2(n16107), .ZN(n16117) );
  NAND2_X1 U17238 ( .A1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15350) );
  INV_X1 U17239 ( .A(n15350), .ZN(n15321) );
  OAI21_X1 U17240 ( .B1(n15321), .B2(n18524), .A(n16462), .ZN(n15385) );
  NOR2_X1 U17241 ( .A1(n15350), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15322) );
  AND2_X1 U17242 ( .A1(n15327), .A2(n15322), .ZN(n15384) );
  NOR2_X1 U17243 ( .A1(n15385), .A2(n15384), .ZN(n16453) );
  NOR2_X1 U17244 ( .A1(n16453), .A2(n16448), .ZN(n15330) );
  OR2_X1 U17245 ( .A1(n15383), .A2(n15323), .ZN(n15324) );
  NAND2_X1 U17246 ( .A1(n16198), .A2(n15324), .ZN(n18414) );
  NAND2_X1 U17247 ( .A1(n18572), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n15333) );
  NOR2_X1 U17248 ( .A1(n15350), .A2(n15325), .ZN(n15326) );
  AND2_X1 U17249 ( .A1(n15327), .A2(n15326), .ZN(n16445) );
  NAND2_X1 U17250 ( .A1(n16445), .A2(n16448), .ZN(n15328) );
  OAI211_X1 U17251 ( .C1(n18594), .C2(n18414), .A(n15333), .B(n15328), .ZN(
        n15329) );
  AOI211_X1 U17252 ( .C1(n18416), .C2(n18591), .A(n15330), .B(n15329), .ZN(
        n15332) );
  NOR2_X1 U17253 ( .A1(n15425), .A2(n16448), .ZN(n16298) );
  INV_X1 U17254 ( .A(n16298), .ZN(n15338) );
  NAND2_X1 U17255 ( .A1(n15425), .A2(n16448), .ZN(n15337) );
  NAND3_X1 U17256 ( .A1(n15338), .A2(n18568), .A3(n15337), .ZN(n15331) );
  OAI211_X1 U17257 ( .C1(n15341), .C2(n18606), .A(n15332), .B(n15331), .ZN(
        P2_U3021) );
  INV_X1 U17258 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n15335) );
  INV_X1 U17259 ( .A(n15447), .ZN(n16295) );
  AOI21_X1 U17260 ( .B1(n15335), .B2(n15390), .A(n16295), .ZN(n18418) );
  NAND2_X1 U17261 ( .A1(n18418), .A2(n17055), .ZN(n15334) );
  OAI211_X1 U17262 ( .C1(n17022), .C2(n15335), .A(n15334), .B(n15333), .ZN(
        n15336) );
  AOI21_X1 U17263 ( .B1(n18416), .B2(n17019), .A(n15336), .ZN(n15340) );
  NAND3_X1 U17264 ( .A1(n15338), .A2(n17047), .A3(n15337), .ZN(n15339) );
  OAI211_X1 U17265 ( .C1(n15341), .C2(n17058), .A(n15340), .B(n15339), .ZN(
        P2_U2989) );
  INV_X1 U17266 ( .A(n15343), .ZN(n15344) );
  NOR2_X1 U17267 ( .A1(n15345), .A2(n15344), .ZN(n15346) );
  XNOR2_X1 U17268 ( .A(n15342), .B(n15346), .ZN(n15372) );
  OAI21_X1 U17269 ( .B1(n15349), .B2(n15348), .A(n15347), .ZN(n16128) );
  INV_X1 U17270 ( .A(n16128), .ZN(n18389) );
  NOR2_X1 U17271 ( .A1(n16462), .A2(n15361), .ZN(n15359) );
  OAI21_X1 U17272 ( .B1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(n15350), .ZN(n15356) );
  NAND2_X1 U17273 ( .A1(n15352), .A2(n15351), .ZN(n15353) );
  NAND2_X1 U17274 ( .A1(n15381), .A2(n15353), .ZN(n18395) );
  INV_X1 U17275 ( .A(n18395), .ZN(n15354) );
  NAND2_X1 U17276 ( .A1(n18622), .A2(n15354), .ZN(n15355) );
  NAND2_X1 U17277 ( .A1(n18572), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n15367) );
  OAI211_X1 U17278 ( .C1(n15357), .C2(n15356), .A(n15355), .B(n15367), .ZN(
        n15358) );
  AOI211_X1 U17279 ( .C1(n18389), .C2(n18591), .A(n15359), .B(n15358), .ZN(
        n15363) );
  AOI21_X1 U17280 ( .B1(n15361), .B2(n15360), .A(n15373), .ZN(n15369) );
  NAND2_X1 U17281 ( .A1(n15369), .A2(n18568), .ZN(n15362) );
  OAI211_X1 U17282 ( .C1(n15372), .C2(n18606), .A(n15363), .B(n15362), .ZN(
        P2_U3023) );
  NOR2_X1 U17283 ( .A1(n15364), .A2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15365) );
  OR2_X1 U17284 ( .A1(n15391), .A2(n15365), .ZN(n18391) );
  NAND2_X1 U17285 ( .A1(n17052), .A2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15366) );
  OAI211_X1 U17286 ( .C1(n18391), .C2(n17046), .A(n15367), .B(n15366), .ZN(
        n15368) );
  AOI21_X1 U17287 ( .B1(n18389), .B2(n17019), .A(n15368), .ZN(n15371) );
  NAND2_X1 U17288 ( .A1(n15369), .A2(n17047), .ZN(n15370) );
  OAI211_X1 U17289 ( .C1(n15372), .C2(n17058), .A(n15371), .B(n15370), .ZN(
        P2_U2991) );
  OAI21_X1 U17290 ( .B1(n15373), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n15425), .ZN(n15398) );
  XNOR2_X1 U17291 ( .A(n15374), .B(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15375) );
  XNOR2_X1 U17292 ( .A(n15376), .B(n15375), .ZN(n15396) );
  INV_X1 U17293 ( .A(n15377), .ZN(n15378) );
  AOI21_X1 U17294 ( .B1(n15379), .B2(n15347), .A(n15378), .ZN(n18401) );
  INV_X1 U17295 ( .A(n18401), .ZN(n16123) );
  AND2_X1 U17296 ( .A1(n15381), .A2(n15380), .ZN(n15382) );
  NOR2_X1 U17297 ( .A1(n15383), .A2(n15382), .ZN(n18400) );
  NOR2_X1 U17298 ( .A1(n18589), .A2(n18396), .ZN(n15392) );
  AOI211_X1 U17299 ( .C1(n18622), .C2(n18400), .A(n15384), .B(n15392), .ZN(
        n15387) );
  NAND2_X1 U17300 ( .A1(n15385), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15386) );
  OAI211_X1 U17301 ( .C1(n16123), .C2(n18605), .A(n15387), .B(n15386), .ZN(
        n15388) );
  AOI21_X1 U17302 ( .B1(n15396), .B2(n18598), .A(n15388), .ZN(n15389) );
  OAI21_X1 U17303 ( .B1(n18617), .B2(n15398), .A(n15389), .ZN(P2_U3022) );
  OAI21_X1 U17304 ( .B1(n15391), .B2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n15390), .ZN(n18404) );
  NAND2_X1 U17305 ( .A1(n18401), .A2(n17019), .ZN(n15394) );
  AOI21_X1 U17306 ( .B1(n17052), .B2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n15392), .ZN(n15393) );
  OAI211_X1 U17307 ( .C1(n17046), .C2(n18404), .A(n15394), .B(n15393), .ZN(
        n15395) );
  AOI21_X1 U17308 ( .B1(n15396), .B2(n17039), .A(n15395), .ZN(n15397) );
  OAI21_X1 U17309 ( .B1(n17042), .B2(n15398), .A(n15397), .ZN(P2_U2990) );
  INV_X1 U17310 ( .A(P2_EBX_REG_26__SCAN_IN), .ZN(n18426) );
  NOR2_X1 U17311 ( .A1(n15131), .A2(n18426), .ZN(n15402) );
  XOR2_X1 U17312 ( .A(n15402), .B(n15403), .Z(n18428) );
  INV_X1 U17313 ( .A(n18428), .ZN(n15400) );
  NOR2_X1 U17314 ( .A1(n15400), .A2(n15139), .ZN(n15401) );
  NAND3_X1 U17315 ( .A1(n18428), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        n15420), .ZN(n15409) );
  OAI21_X1 U17316 ( .B1(n15401), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n15409), .ZN(n16293) );
  NAND2_X1 U17317 ( .A1(n16684), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n15404) );
  NOR2_X1 U17318 ( .A1(n11022), .A2(n15404), .ZN(n15405) );
  INV_X1 U17319 ( .A(n18441), .ZN(n15406) );
  NAND2_X1 U17320 ( .A1(n15406), .A2(n15420), .ZN(n16280) );
  INV_X1 U17321 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n16413) );
  NAND2_X1 U17322 ( .A1(n16280), .A2(n16413), .ZN(n16271) );
  NAND2_X1 U17323 ( .A1(n16684), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n15410) );
  XOR2_X1 U17324 ( .A(n15410), .B(n15411), .Z(n18458) );
  OAI21_X1 U17325 ( .B1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(n16273), .ZN(n15408) );
  INV_X1 U17326 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n16427) );
  INV_X1 U17327 ( .A(n16273), .ZN(n15407) );
  NAND2_X1 U17328 ( .A1(n15409), .A2(n16290), .ZN(n16269) );
  INV_X1 U17329 ( .A(P2_EBX_REG_29__SCAN_IN), .ZN(n18469) );
  NOR2_X1 U17330 ( .A1(n15131), .A2(n18469), .ZN(n15412) );
  XOR2_X1 U17331 ( .A(n15412), .B(n15413), .Z(n18472) );
  AOI21_X1 U17332 ( .B1(n18472), .B2(n15420), .A(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16257) );
  INV_X1 U17333 ( .A(P2_EBX_REG_30__SCAN_IN), .ZN(n15414) );
  NOR2_X1 U17334 ( .A1(n15131), .A2(n15414), .ZN(n15416) );
  XNOR2_X1 U17335 ( .A(n15417), .B(n15416), .ZN(n18488) );
  INV_X1 U17336 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15487) );
  OAI21_X1 U17337 ( .B1(n18488), .B2(n15139), .A(n15487), .ZN(n15476) );
  NOR2_X1 U17338 ( .A1(n15417), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n15418) );
  MUX2_X1 U17339 ( .A(n15419), .B(n15418), .S(n16684), .Z(n18500) );
  NAND2_X1 U17340 ( .A1(n18500), .A2(n15420), .ZN(n15421) );
  XOR2_X1 U17341 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n15421), .Z(
        n15422) );
  XNOR2_X1 U17342 ( .A(n15423), .B(n15422), .ZN(n15474) );
  AND2_X1 U17343 ( .A1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n16447) );
  INV_X1 U17344 ( .A(n16447), .ZN(n15424) );
  NAND4_X1 U17345 ( .A1(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A4(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15465) );
  NOR2_X1 U17346 ( .A1(n16297), .A2(n15465), .ZN(n15480) );
  XOR2_X1 U17347 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n15480), .Z(
        n15472) );
  INV_X1 U17348 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n16452) );
  AOI22_X1 U17349 ( .A1(n15227), .A2(P2_EBX_REG_26__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), 
        .ZN(n15427) );
  NAND2_X1 U17350 ( .A1(n15440), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n15426) );
  OAI211_X1 U17351 ( .C1(n15443), .C2(n16452), .A(n15427), .B(n15426), .ZN(
        n16106) );
  INV_X1 U17352 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n18438) );
  NAND2_X1 U17353 ( .A1(n15227), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n15429) );
  NAND2_X1 U17354 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n15428) );
  OAI211_X1 U17355 ( .C1(n10963), .C2(n18438), .A(n15429), .B(n15428), .ZN(
        n15430) );
  AOI21_X1 U17356 ( .B1(n13924), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n15430), .ZN(n16101) );
  NAND2_X1 U17357 ( .A1(n15227), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n15432) );
  NAND2_X1 U17358 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n15431) );
  OAI211_X1 U17359 ( .C1(n10963), .C2(n18454), .A(n15432), .B(n15431), .ZN(
        n15433) );
  AOI21_X1 U17360 ( .B1(n13924), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n15433), .ZN(n16092) );
  INV_X1 U17361 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n18468) );
  NAND2_X1 U17362 ( .A1(n15227), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n15435) );
  NAND2_X1 U17363 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n15434) );
  OAI211_X1 U17364 ( .C1(n10963), .C2(n18468), .A(n15435), .B(n15434), .ZN(
        n15437) );
  AOI21_X1 U17365 ( .B1(n13924), .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n15437), .ZN(n16081) );
  AOI22_X1 U17366 ( .A1(n15227), .A2(P2_EBX_REG_30__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), 
        .ZN(n15439) );
  NAND2_X1 U17367 ( .A1(n15440), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n15438) );
  OAI211_X1 U17368 ( .C1(n15443), .C2(n15487), .A(n15439), .B(n15438), .ZN(
        n15481) );
  NAND2_X1 U17369 ( .A1(n16082), .A2(n15481), .ZN(n15445) );
  INV_X1 U17370 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n16018) );
  AOI22_X1 U17371 ( .A1(n15227), .A2(P2_EBX_REG_31__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n15442) );
  NAND2_X1 U17372 ( .A1(n15440), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n15441) );
  OAI211_X1 U17373 ( .C1(n15443), .C2(n16018), .A(n15442), .B(n15441), .ZN(
        n15444) );
  INV_X1 U17374 ( .A(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n15446) );
  INV_X1 U17375 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n18442) );
  INV_X1 U17376 ( .A(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n16264) );
  INV_X1 U17377 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n18501) );
  NOR2_X1 U17378 ( .A1(n18589), .A2(n18501), .ZN(n15466) );
  AOI21_X1 U17379 ( .B1(n17052), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n15466), .ZN(n15449) );
  INV_X1 U17380 ( .A(n15450), .ZN(n15451) );
  AOI21_X1 U17381 ( .B1(n15472), .B2(n17047), .A(n15453), .ZN(n15454) );
  OAI21_X1 U17382 ( .B1(n15474), .B2(n17058), .A(n15454), .ZN(P2_U2983) );
  NAND2_X1 U17383 ( .A1(n18508), .A2(n18591), .ZN(n15470) );
  INV_X1 U17384 ( .A(n15455), .ZN(n15460) );
  NAND2_X1 U17385 ( .A1(n15456), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n15458) );
  AOI22_X1 U17386 ( .A1(n15461), .A2(P2_EAX_REG_30__SCAN_IN), .B1(n13405), 
        .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15457) );
  AND2_X1 U17387 ( .A1(n15458), .A2(n15457), .ZN(n15482) );
  INV_X1 U17388 ( .A(n15482), .ZN(n15459) );
  NAND2_X1 U17389 ( .A1(n15460), .A2(n15459), .ZN(n15484) );
  AOI22_X1 U17390 ( .A1(n15461), .A2(P2_EAX_REG_31__SCAN_IN), .B1(n13405), 
        .B2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n15462) );
  OAI21_X1 U17391 ( .B1(n18501), .B2(n15463), .A(n15462), .ZN(n15464) );
  XNOR2_X1 U17392 ( .A(n15484), .B(n15464), .ZN(n19113) );
  OAI21_X1 U17393 ( .B1(n16447), .B2(n18524), .A(n16453), .ZN(n16434) );
  AOI21_X1 U17394 ( .B1(n15465), .B2(n18555), .A(n16434), .ZN(n15488) );
  NAND2_X1 U17395 ( .A1(n16445), .A2(n16447), .ZN(n16416) );
  AOI21_X1 U17396 ( .B1(n15472), .B2(n18568), .A(n15471), .ZN(n15473) );
  OAI21_X1 U17397 ( .B1(n15474), .B2(n18606), .A(n15473), .ZN(P2_U3015) );
  NOR2_X1 U17398 ( .A1(n15475), .A2(n16256), .ZN(n15478) );
  NAND2_X1 U17399 ( .A1(n10985), .A2(n15476), .ZN(n15477) );
  XNOR2_X1 U17400 ( .A(n15478), .B(n15477), .ZN(n16255) );
  AND2_X1 U17401 ( .A1(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15479) );
  AOI21_X1 U17402 ( .B1(n16260), .B2(n15487), .A(n15480), .ZN(n16253) );
  NAND2_X1 U17403 ( .A1(n15455), .A2(n15482), .ZN(n15483) );
  NAND3_X1 U17404 ( .A1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15485) );
  INV_X1 U17405 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n18485) );
  NOR2_X1 U17406 ( .A1(n18589), .A2(n18485), .ZN(n16250) );
  INV_X1 U17407 ( .A(n16250), .ZN(n15486) );
  OAI211_X1 U17408 ( .C1(n15488), .C2(n15487), .A(n11478), .B(n15486), .ZN(
        n15489) );
  NAND3_X1 U17409 ( .A1(n15533), .A2(P1_REIP_REG_29__SCAN_IN), .A3(n21639), 
        .ZN(n15503) );
  NAND2_X1 U17410 ( .A1(n15531), .A2(n15494), .ZN(n15495) );
  NAND2_X1 U17411 ( .A1(n11011), .A2(n15495), .ZN(n15853) );
  INV_X1 U17412 ( .A(n15853), .ZN(n15501) );
  NAND2_X1 U17413 ( .A1(n21627), .A2(n15496), .ZN(n15498) );
  NAND2_X1 U17414 ( .A1(n21626), .A2(P1_EBX_REG_29__SCAN_IN), .ZN(n15497) );
  OAI211_X1 U17415 ( .C1(n21636), .C2(n15499), .A(n15498), .B(n15497), .ZN(
        n15500) );
  AOI21_X1 U17416 ( .B1(n15501), .B2(n21633), .A(n15500), .ZN(n15502) );
  OAI211_X1 U17417 ( .C1(n15533), .C2(P1_REIP_REG_29__SCAN_IN), .A(n15503), 
        .B(n15502), .ZN(n15504) );
  INV_X1 U17418 ( .A(n15504), .ZN(n15505) );
  OAI21_X1 U17419 ( .B1(n15493), .B2(n21648), .A(n15505), .ZN(P1_U2811) );
  AOI22_X1 U17420 ( .A1(n15682), .A2(DATAI_29_), .B1(P1_EAX_REG_29__SCAN_IN), 
        .B2(n15707), .ZN(n15509) );
  AOI22_X1 U17421 ( .A1(n15684), .A2(n15507), .B1(n15694), .B2(
        BUF1_REG_29__SCAN_IN), .ZN(n15508) );
  OAI211_X1 U17422 ( .C1(n15493), .C2(n15711), .A(n15509), .B(n15508), .ZN(
        P1_U2875) );
  OAI222_X1 U17423 ( .A1(n15510), .A2(n19969), .B1(n19965), .B2(n15853), .C1(
        n15493), .C2(n19966), .ZN(P1_U2843) );
  AND2_X1 U17424 ( .A1(n15511), .A2(n19931), .ZN(n15526) );
  NAND2_X1 U17425 ( .A1(n15721), .A2(n21611), .ZN(n15524) );
  NAND2_X1 U17426 ( .A1(n11011), .A2(n15514), .ZN(n15517) );
  OR2_X1 U17427 ( .A1(n15531), .A2(n15515), .ZN(n15516) );
  NAND2_X1 U17428 ( .A1(n15517), .A2(n15516), .ZN(n15519) );
  XNOR2_X1 U17429 ( .A(n15519), .B(n15518), .ZN(n15846) );
  INV_X1 U17430 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n15719) );
  NAND2_X1 U17431 ( .A1(n21627), .A2(n15717), .ZN(n15521) );
  NAND2_X1 U17432 ( .A1(n21626), .A2(P1_EBX_REG_30__SCAN_IN), .ZN(n15520) );
  OAI211_X1 U17433 ( .C1(n21636), .C2(n15719), .A(n15521), .B(n15520), .ZN(
        n15522) );
  AOI21_X1 U17434 ( .B1(n15846), .B2(n21633), .A(n15522), .ZN(n15523) );
  OAI211_X1 U17435 ( .C1(n15526), .C2(n15525), .A(n15524), .B(n15523), .ZN(
        P1_U2810) );
  INV_X1 U17436 ( .A(n15527), .ZN(n15528) );
  AOI21_X1 U17437 ( .B1(n15528), .B2(n10983), .A(n12379), .ZN(n15731) );
  INV_X1 U17438 ( .A(n15731), .ZN(n15636) );
  OR2_X1 U17439 ( .A1(n11019), .A2(n15529), .ZN(n15530) );
  AND2_X1 U17440 ( .A1(n15531), .A2(n15530), .ZN(n15866) );
  AOI22_X1 U17441 ( .A1(n21645), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .B1(
        n21626), .B2(P1_EBX_REG_28__SCAN_IN), .ZN(n15532) );
  OAI21_X1 U17442 ( .B1(n15729), .B2(n21642), .A(n15532), .ZN(n15537) );
  AOI21_X1 U17443 ( .B1(P1_REIP_REG_28__SCAN_IN), .B2(n21639), .A(n15550), 
        .ZN(n15535) );
  INV_X1 U17444 ( .A(n15533), .ZN(n15534) );
  NOR2_X1 U17445 ( .A1(n15535), .A2(n15534), .ZN(n15536) );
  AOI211_X1 U17446 ( .C1(n21633), .C2(n15866), .A(n15537), .B(n15536), .ZN(
        n15538) );
  OAI21_X1 U17447 ( .B1(n15636), .B2(n21648), .A(n15538), .ZN(P1_U2812) );
  AOI21_X1 U17448 ( .B1(P1_REIP_REG_27__SCAN_IN), .B2(n21639), .A(n21654), 
        .ZN(n15549) );
  INV_X1 U17449 ( .A(n15736), .ZN(n15542) );
  NAND2_X1 U17450 ( .A1(n15542), .A2(n21611), .ZN(n15548) );
  INV_X1 U17451 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n15735) );
  INV_X1 U17452 ( .A(P1_EBX_REG_27__SCAN_IN), .ZN(n15571) );
  OAI22_X1 U17453 ( .A1(n21636), .A2(n15735), .B1(n21640), .B2(n15571), .ZN(
        n15546) );
  INV_X1 U17454 ( .A(n15871), .ZN(n15573) );
  AOI21_X1 U17455 ( .B1(n15573), .B2(n15869), .A(n15543), .ZN(n15544) );
  OR2_X1 U17456 ( .A1(n15544), .A2(n11019), .ZN(n21382) );
  NOR2_X1 U17457 ( .A1(n21382), .A2(n21646), .ZN(n15545) );
  AOI211_X1 U17458 ( .C1(n21627), .C2(n15739), .A(n15546), .B(n15545), .ZN(
        n15547) );
  OAI211_X1 U17459 ( .C1(n15550), .C2(n15549), .A(n15548), .B(n15547), .ZN(
        P1_U2813) );
  OAI21_X1 U17460 ( .B1(n11028), .B2(n15552), .A(n15551), .ZN(n15758) );
  AND2_X1 U17461 ( .A1(n15586), .A2(n15553), .ZN(n15554) );
  NOR2_X1 U17462 ( .A1(n15579), .A2(n15554), .ZN(n21402) );
  AOI22_X1 U17463 ( .A1(n15761), .A2(n21627), .B1(P1_EBX_REG_23__SCAN_IN), 
        .B2(n21626), .ZN(n15555) );
  OAI21_X1 U17464 ( .B1(n15757), .B2(n21636), .A(n15555), .ZN(n15557) );
  AOI211_X1 U17465 ( .C1(n11060), .C2(n19913), .A(n21523), .B(n21617), .ZN(
        n15556) );
  AOI211_X1 U17466 ( .C1(n21402), .C2(n21633), .A(n15557), .B(n15556), .ZN(
        n15558) );
  OAI21_X1 U17467 ( .B1(n15758), .B2(n21648), .A(n15558), .ZN(P1_U2817) );
  AOI21_X1 U17468 ( .B1(n15561), .B2(n15559), .A(n15560), .ZN(n15792) );
  INV_X1 U17469 ( .A(n15792), .ZN(n15687) );
  INV_X1 U17470 ( .A(n15612), .ZN(n15562) );
  AOI21_X1 U17471 ( .B1(n15563), .B2(n15624), .A(n15562), .ZN(n21360) );
  AOI22_X1 U17472 ( .A1(n15788), .A2(n21627), .B1(P1_EBX_REG_17__SCAN_IN), 
        .B2(n21626), .ZN(n15564) );
  OAI211_X1 U17473 ( .C1(n21636), .C2(n12022), .A(n15564), .B(n21571), .ZN(
        n15566) );
  OR2_X1 U17474 ( .A1(n21563), .A2(n21523), .ZN(n21581) );
  AOI21_X1 U17475 ( .B1(n11009), .B2(n21366), .A(n21581), .ZN(n15565) );
  AOI211_X1 U17476 ( .C1(n21360), .C2(n21633), .A(n15566), .B(n15565), .ZN(
        n15567) );
  OAI21_X1 U17477 ( .B1(n15687), .B2(n21648), .A(n15567), .ZN(P1_U2823) );
  INV_X1 U17478 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n15568) );
  OAI22_X1 U17479 ( .A1(n15806), .A2(n19965), .B1(n15568), .B2(n19969), .ZN(
        P1_U2841) );
  INV_X1 U17480 ( .A(n15721), .ZN(n15632) );
  AOI22_X1 U17481 ( .A1(n15846), .A2(n19961), .B1(n15617), .B2(
        P1_EBX_REG_30__SCAN_IN), .ZN(n15569) );
  OAI21_X1 U17482 ( .B1(n15632), .B2(n19966), .A(n15569), .ZN(P1_U2842) );
  AOI22_X1 U17483 ( .A1(n15866), .A2(n19961), .B1(n15617), .B2(
        P1_EBX_REG_28__SCAN_IN), .ZN(n15570) );
  OAI21_X1 U17484 ( .B1(n15636), .B2(n15628), .A(n15570), .ZN(P1_U2844) );
  OAI222_X1 U17485 ( .A1(n15571), .A2(n19969), .B1(n19965), .B2(n21382), .C1(
        n15736), .C2(n19966), .ZN(P1_U2845) );
  AOI21_X1 U17486 ( .B1(n15574), .B2(n15577), .A(n15573), .ZN(n21632) );
  AOI22_X1 U17487 ( .A1(n21632), .A2(n19961), .B1(P1_EBX_REG_25__SCAN_IN), 
        .B2(n15617), .ZN(n15575) );
  OAI21_X1 U17488 ( .B1(n21630), .B2(n15628), .A(n15575), .ZN(P1_U2847) );
  AOI21_X1 U17489 ( .B1(n15576), .B2(n15551), .A(n15572), .ZN(n20025) );
  INV_X1 U17490 ( .A(n20025), .ZN(n21621) );
  OAI21_X1 U17491 ( .B1(n15579), .B2(n15578), .A(n15577), .ZN(n21620) );
  INV_X1 U17492 ( .A(n21620), .ZN(n15892) );
  AOI22_X1 U17493 ( .A1(n15892), .A2(n19961), .B1(n15617), .B2(
        P1_EBX_REG_24__SCAN_IN), .ZN(n15580) );
  OAI21_X1 U17494 ( .B1(n21621), .B2(n15628), .A(n15580), .ZN(P1_U2848) );
  AOI22_X1 U17495 ( .A1(n21402), .A2(n19961), .B1(P1_EBX_REG_23__SCAN_IN), 
        .B2(n15617), .ZN(n15581) );
  OAI21_X1 U17496 ( .B1(n15758), .B2(n15628), .A(n15581), .ZN(P1_U2849) );
  AND2_X1 U17497 ( .A1(n11018), .A2(n15582), .ZN(n15583) );
  NAND2_X1 U17498 ( .A1(n15592), .A2(n15584), .ZN(n15585) );
  NAND2_X1 U17499 ( .A1(n15586), .A2(n15585), .ZN(n21604) );
  OAI22_X1 U17500 ( .A1(n21604), .A2(n19965), .B1(n15587), .B2(n19969), .ZN(
        n15588) );
  INV_X1 U17501 ( .A(n15588), .ZN(n15589) );
  OAI21_X1 U17502 ( .B1(n21603), .B2(n15628), .A(n15589), .ZN(P1_U2850) );
  INV_X1 U17503 ( .A(n15590), .ZN(n15591) );
  OAI21_X1 U17504 ( .B1(n10987), .B2(n15591), .A(n11018), .ZN(n21594) );
  AOI21_X1 U17505 ( .B1(n15593), .B2(n10999), .A(n11300), .ZN(n21591) );
  AOI22_X1 U17506 ( .A1(n21591), .A2(n19961), .B1(P1_EBX_REG_21__SCAN_IN), 
        .B2(n15617), .ZN(n15594) );
  OAI21_X1 U17507 ( .B1(n21594), .B2(n15628), .A(n15594), .ZN(P1_U2851) );
  INV_X1 U17508 ( .A(n15596), .ZN(n15603) );
  AOI21_X1 U17509 ( .B1(n11468), .B2(n15603), .A(n10987), .ZN(n20014) );
  INV_X1 U17510 ( .A(n20014), .ZN(n21584) );
  OR2_X1 U17511 ( .A1(n15607), .A2(n15597), .ZN(n15598) );
  NAND2_X1 U17512 ( .A1(n10999), .A2(n15598), .ZN(n21583) );
  OAI22_X1 U17513 ( .A1(n21583), .A2(n19965), .B1(n15599), .B2(n19969), .ZN(
        n15600) );
  INV_X1 U17514 ( .A(n15600), .ZN(n15601) );
  OAI21_X1 U17515 ( .B1(n21584), .B2(n15628), .A(n15601), .ZN(P1_U2852) );
  OAI21_X1 U17516 ( .B1(n15604), .B2(n15602), .A(n15603), .ZN(n21575) );
  INV_X1 U17517 ( .A(P1_EBX_REG_19__SCAN_IN), .ZN(n15608) );
  NOR2_X1 U17518 ( .A1(n15613), .A2(n15605), .ZN(n15606) );
  OR2_X1 U17519 ( .A1(n15607), .A2(n15606), .ZN(n21368) );
  OAI222_X1 U17520 ( .A1(n21575), .A2(n15628), .B1(n19969), .B2(n15608), .C1(
        n21368), .C2(n19965), .ZN(P1_U2853) );
  AND2_X1 U17521 ( .A1(n11471), .A2(n15609), .ZN(n15610) );
  NOR2_X1 U17522 ( .A1(n15602), .A2(n15610), .ZN(n21567) );
  INV_X1 U17523 ( .A(n21567), .ZN(n15681) );
  AND2_X1 U17524 ( .A1(n15612), .A2(n15611), .ZN(n15614) );
  OR2_X1 U17525 ( .A1(n15614), .A2(n15613), .ZN(n21559) );
  OAI22_X1 U17526 ( .A1(n21559), .A2(n19965), .B1(n21560), .B2(n19969), .ZN(
        n15615) );
  INV_X1 U17527 ( .A(n15615), .ZN(n15616) );
  OAI21_X1 U17528 ( .B1(n15681), .B2(n15628), .A(n15616), .ZN(P1_U2854) );
  AOI22_X1 U17529 ( .A1(n21360), .A2(n19961), .B1(P1_EBX_REG_17__SCAN_IN), 
        .B2(n15617), .ZN(n15618) );
  OAI21_X1 U17530 ( .B1(n15687), .B2(n15628), .A(n15618), .ZN(P1_U2855) );
  NAND2_X1 U17531 ( .A1(n15620), .A2(n15619), .ZN(n15621) );
  AND2_X1 U17532 ( .A1(n15559), .A2(n15621), .ZN(n21554) );
  INV_X1 U17533 ( .A(n21554), .ZN(n15696) );
  OR2_X1 U17534 ( .A1(n15949), .A2(n15622), .ZN(n15623) );
  NAND2_X1 U17535 ( .A1(n15624), .A2(n15623), .ZN(n21558) );
  OAI22_X1 U17536 ( .A1(n21558), .A2(n19965), .B1(n15625), .B2(n19969), .ZN(
        n15626) );
  INV_X1 U17537 ( .A(n15626), .ZN(n15627) );
  OAI21_X1 U17538 ( .B1(n15696), .B2(n15628), .A(n15627), .ZN(P1_U2856) );
  OAI22_X1 U17539 ( .A1(n15689), .A2(n16879), .B1(n14386), .B2(n15703), .ZN(
        n15629) );
  INV_X1 U17540 ( .A(n15629), .ZN(n15631) );
  AOI22_X1 U17541 ( .A1(n15684), .A2(n15708), .B1(n15694), .B2(
        BUF1_REG_30__SCAN_IN), .ZN(n15630) );
  OAI211_X1 U17542 ( .C1(n15632), .C2(n15711), .A(n15631), .B(n15630), .ZN(
        P1_U2874) );
  AOI22_X1 U17543 ( .A1(n15682), .A2(DATAI_28_), .B1(P1_EAX_REG_28__SCAN_IN), 
        .B2(n15707), .ZN(n15635) );
  AOI22_X1 U17544 ( .A1(n15684), .A2(n15633), .B1(n15694), .B2(
        BUF1_REG_28__SCAN_IN), .ZN(n15634) );
  OAI211_X1 U17545 ( .C1(n15636), .C2(n15711), .A(n15635), .B(n15634), .ZN(
        P1_U2876) );
  AOI22_X1 U17546 ( .A1(n15682), .A2(DATAI_27_), .B1(P1_EAX_REG_27__SCAN_IN), 
        .B2(n15707), .ZN(n15639) );
  AOI22_X1 U17547 ( .A1(n15684), .A2(n15637), .B1(n15694), .B2(
        BUF1_REG_27__SCAN_IN), .ZN(n15638) );
  OAI211_X1 U17548 ( .C1(n15736), .C2(n15711), .A(n15639), .B(n15638), .ZN(
        P1_U2877) );
  AND2_X1 U17549 ( .A1(n10982), .A2(n15640), .ZN(n15641) );
  OAI22_X1 U17550 ( .A1(n15689), .A2(n16873), .B1(n14339), .B2(n15703), .ZN(
        n15644) );
  INV_X1 U17551 ( .A(n15684), .ZN(n15691) );
  NOR2_X1 U17552 ( .A1(n15691), .A2(n15642), .ZN(n15643) );
  AOI211_X1 U17553 ( .C1(n15694), .C2(BUF1_REG_26__SCAN_IN), .A(n15644), .B(
        n15643), .ZN(n15645) );
  OAI21_X1 U17554 ( .B1(n21649), .B2(n15711), .A(n15645), .ZN(P1_U2878) );
  OAI22_X1 U17555 ( .A1(n15689), .A2(n14242), .B1(n15646), .B2(n15703), .ZN(
        n15649) );
  NOR2_X1 U17556 ( .A1(n15691), .A2(n15647), .ZN(n15648) );
  AOI211_X1 U17557 ( .C1(BUF1_REG_25__SCAN_IN), .C2(n15694), .A(n15649), .B(
        n15648), .ZN(n15650) );
  OAI21_X1 U17558 ( .B1(n21630), .B2(n15711), .A(n15650), .ZN(P1_U2879) );
  OAI22_X1 U17559 ( .A1(n15689), .A2(n16793), .B1(n15651), .B2(n15703), .ZN(
        n15654) );
  NOR2_X1 U17560 ( .A1(n15691), .A2(n15652), .ZN(n15653) );
  AOI211_X1 U17561 ( .C1(n15694), .C2(BUF1_REG_24__SCAN_IN), .A(n15654), .B(
        n15653), .ZN(n15655) );
  OAI21_X1 U17562 ( .B1(n21621), .B2(n15711), .A(n15655), .ZN(P1_U2880) );
  AOI22_X1 U17563 ( .A1(n15682), .A2(DATAI_23_), .B1(P1_EAX_REG_23__SCAN_IN), 
        .B2(n15707), .ZN(n15658) );
  AOI22_X1 U17564 ( .A1(n15684), .A2(n15656), .B1(n15694), .B2(
        BUF1_REG_23__SCAN_IN), .ZN(n15657) );
  OAI211_X1 U17565 ( .C1(n15758), .C2(n15711), .A(n15658), .B(n15657), .ZN(
        P1_U2881) );
  OAI22_X1 U17566 ( .A1(n15689), .A2(n16895), .B1(n15659), .B2(n15703), .ZN(
        n15662) );
  NOR2_X1 U17567 ( .A1(n15691), .A2(n15660), .ZN(n15661) );
  AOI211_X1 U17568 ( .C1(n15694), .C2(BUF1_REG_22__SCAN_IN), .A(n15662), .B(
        n15661), .ZN(n15663) );
  OAI21_X1 U17569 ( .B1(n21603), .B2(n15711), .A(n15663), .ZN(P1_U2882) );
  AOI22_X1 U17570 ( .A1(n15682), .A2(DATAI_21_), .B1(P1_EAX_REG_21__SCAN_IN), 
        .B2(n15707), .ZN(n15666) );
  AOI22_X1 U17571 ( .A1(n15684), .A2(n15664), .B1(n15694), .B2(
        BUF1_REG_21__SCAN_IN), .ZN(n15665) );
  OAI211_X1 U17572 ( .C1(n21594), .C2(n15711), .A(n15666), .B(n15665), .ZN(
        P1_U2883) );
  OAI22_X1 U17573 ( .A1(n15689), .A2(n16780), .B1(n15667), .B2(n15703), .ZN(
        n15670) );
  NOR2_X1 U17574 ( .A1(n15691), .A2(n15668), .ZN(n15669) );
  AOI211_X1 U17575 ( .C1(n15694), .C2(BUF1_REG_20__SCAN_IN), .A(n15670), .B(
        n15669), .ZN(n15671) );
  OAI21_X1 U17576 ( .B1(n21584), .B2(n15711), .A(n15671), .ZN(P1_U2884) );
  AOI22_X1 U17577 ( .A1(n15682), .A2(DATAI_19_), .B1(P1_EAX_REG_19__SCAN_IN), 
        .B2(n15707), .ZN(n15674) );
  AOI22_X1 U17578 ( .A1(n15684), .A2(n15672), .B1(n15694), .B2(
        BUF1_REG_19__SCAN_IN), .ZN(n15673) );
  OAI211_X1 U17579 ( .C1(n21575), .C2(n15711), .A(n15674), .B(n15673), .ZN(
        P1_U2885) );
  NOR2_X1 U17580 ( .A1(n15703), .A2(n15675), .ZN(n15679) );
  INV_X1 U17581 ( .A(n15694), .ZN(n15676) );
  OAI22_X1 U17582 ( .A1(n15691), .A2(n15677), .B1(n15676), .B2(n20071), .ZN(
        n15678) );
  AOI211_X1 U17583 ( .C1(DATAI_18_), .C2(n15682), .A(n15679), .B(n15678), .ZN(
        n15680) );
  OAI21_X1 U17584 ( .B1(n15681), .B2(n15711), .A(n15680), .ZN(P1_U2886) );
  AOI22_X1 U17585 ( .A1(n15682), .A2(DATAI_17_), .B1(P1_EAX_REG_17__SCAN_IN), 
        .B2(n15707), .ZN(n15686) );
  AOI22_X1 U17586 ( .A1(n15684), .A2(n15683), .B1(n15694), .B2(
        BUF1_REG_17__SCAN_IN), .ZN(n15685) );
  OAI211_X1 U17587 ( .C1(n15687), .C2(n15711), .A(n15686), .B(n15685), .ZN(
        P1_U2887) );
  OAI22_X1 U17588 ( .A1(n15689), .A2(n13899), .B1(n15688), .B2(n15703), .ZN(
        n15693) );
  NOR2_X1 U17589 ( .A1(n15691), .A2(n15690), .ZN(n15692) );
  AOI211_X1 U17590 ( .C1(n15694), .C2(BUF1_REG_16__SCAN_IN), .A(n15693), .B(
        n15692), .ZN(n15695) );
  OAI21_X1 U17591 ( .B1(n15696), .B2(n15711), .A(n15695), .ZN(P1_U2888) );
  XOR2_X1 U17592 ( .A(n15698), .B(n15697), .Z(n21547) );
  INV_X1 U17593 ( .A(n21547), .ZN(n15699) );
  OAI222_X1 U17594 ( .A1(n15703), .A2(n15702), .B1(n15701), .B2(n15700), .C1(
        n15711), .C2(n15699), .ZN(P1_U2889) );
  INV_X1 U17595 ( .A(n15704), .ZN(n15706) );
  INV_X1 U17596 ( .A(n15088), .ZN(n15705) );
  AOI21_X1 U17597 ( .B1(n15706), .B2(n15705), .A(n15697), .ZN(n21535) );
  INV_X1 U17598 ( .A(n21535), .ZN(n15712) );
  AOI22_X1 U17599 ( .A1(n15709), .A2(n15708), .B1(P1_EAX_REG_14__SCAN_IN), 
        .B2(n15707), .ZN(n15710) );
  OAI21_X1 U17600 ( .B1(n15712), .B2(n15711), .A(n15710), .ZN(P1_U2890) );
  NAND2_X1 U17601 ( .A1(n15994), .A2(n15858), .ZN(n15713) );
  NAND2_X1 U17602 ( .A1(n15860), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15827) );
  MUX2_X1 U17603 ( .A(n15713), .B(n15827), .S(n15734), .Z(n15715) );
  XNOR2_X1 U17604 ( .A(n15716), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15848) );
  NAND2_X1 U17605 ( .A1(n20005), .A2(n15717), .ZN(n15718) );
  NAND2_X1 U17606 ( .A1(n10970), .A2(P1_REIP_REG_30__SCAN_IN), .ZN(n15841) );
  OAI211_X1 U17607 ( .C1(n15719), .C2(n19987), .A(n15718), .B(n15841), .ZN(
        n15720) );
  AOI21_X1 U17608 ( .B1(n15721), .B2(n20009), .A(n15720), .ZN(n15722) );
  OAI21_X1 U17609 ( .B1(n15848), .B2(n21655), .A(n15722), .ZN(P1_U2969) );
  INV_X1 U17610 ( .A(n15882), .ZN(n15880) );
  NAND3_X1 U17611 ( .A1(n15880), .A2(n15741), .A3(n11082), .ZN(n15726) );
  NAND3_X1 U17612 ( .A1(n15882), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A3(
        n15723), .ZN(n15725) );
  MUX2_X1 U17613 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .B(n15741), .S(
        n15881), .Z(n15724) );
  AOI21_X1 U17614 ( .B1(n15726), .B2(n15725), .A(n15724), .ZN(n15727) );
  XNOR2_X1 U17615 ( .A(n15727), .B(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n15868) );
  NAND2_X1 U17616 ( .A1(n10970), .A2(P1_REIP_REG_28__SCAN_IN), .ZN(n15864) );
  NAND2_X1 U17617 ( .A1(n20022), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n15728) );
  OAI211_X1 U17618 ( .C1(n20028), .C2(n15729), .A(n15864), .B(n15728), .ZN(
        n15730) );
  AOI21_X1 U17619 ( .B1(n15731), .B2(n20009), .A(n15730), .ZN(n15732) );
  OAI21_X1 U17620 ( .B1(n21655), .B2(n15868), .A(n15732), .ZN(P1_U2971) );
  XNOR2_X1 U17621 ( .A(n12469), .B(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15733) );
  XNOR2_X1 U17622 ( .A(n15734), .B(n15733), .ZN(n21381) );
  INV_X1 U17623 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n21385) );
  OAI22_X1 U17624 ( .A1(n19987), .A2(n15735), .B1(n21386), .B2(n21385), .ZN(
        n15738) );
  NOR2_X1 U17625 ( .A1(n15736), .A2(n20018), .ZN(n15737) );
  OAI21_X1 U17626 ( .B1(n21381), .B2(n21655), .A(n15740), .ZN(P1_U2972) );
  XNOR2_X1 U17627 ( .A(n15742), .B(n15741), .ZN(n15879) );
  INV_X1 U17628 ( .A(n21649), .ZN(n15745) );
  NAND2_X1 U17629 ( .A1(n10970), .A2(P1_REIP_REG_26__SCAN_IN), .ZN(n15875) );
  NAND2_X1 U17630 ( .A1(n20022), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15743) );
  OAI211_X1 U17631 ( .C1(n21643), .C2(n20028), .A(n15875), .B(n15743), .ZN(
        n15744) );
  AOI21_X1 U17632 ( .B1(n15745), .B2(n20009), .A(n15744), .ZN(n15746) );
  OAI21_X1 U17633 ( .B1(n21655), .B2(n15879), .A(n15746), .ZN(P1_U2973) );
  OAI21_X1 U17634 ( .B1(n15882), .B2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n15872), .ZN(n15748) );
  NAND2_X1 U17635 ( .A1(n15994), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15755) );
  NAND3_X1 U17636 ( .A1(n15748), .A2(n15747), .A3(n15755), .ZN(n15749) );
  XNOR2_X1 U17637 ( .A(n15749), .B(n21398), .ZN(n21394) );
  INV_X1 U17638 ( .A(n21630), .ZN(n15753) );
  INV_X1 U17639 ( .A(n21628), .ZN(n15751) );
  AOI22_X1 U17640 ( .A1(n20022), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .B1(
        n10970), .B2(P1_REIP_REG_25__SCAN_IN), .ZN(n15750) );
  OAI21_X1 U17641 ( .B1(n20028), .B2(n15751), .A(n15750), .ZN(n15752) );
  AOI21_X1 U17642 ( .B1(n15753), .B2(n20009), .A(n15752), .ZN(n15754) );
  OAI21_X1 U17643 ( .B1(n21655), .B2(n21394), .A(n15754), .ZN(P1_U2974) );
  OAI21_X1 U17644 ( .B1(n15994), .B2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n15755), .ZN(n15756) );
  XNOR2_X1 U17645 ( .A(n15880), .B(n15756), .ZN(n21401) );
  OAI22_X1 U17646 ( .A1(n19987), .A2(n15757), .B1(n21386), .B2(n19913), .ZN(
        n15760) );
  NOR2_X1 U17647 ( .A1(n15758), .A2(n20018), .ZN(n15759) );
  AOI211_X1 U17648 ( .C1(n20005), .C2(n15761), .A(n15760), .B(n15759), .ZN(
        n15762) );
  OAI21_X1 U17649 ( .B1(n21401), .B2(n21655), .A(n15762), .ZN(P1_U2976) );
  XNOR2_X1 U17650 ( .A(n15881), .B(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15776) );
  AOI22_X1 U17651 ( .A1(n15777), .A2(n15776), .B1(n15994), .B2(
        P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n15916) );
  NOR2_X1 U17652 ( .A1(n15901), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15919) );
  OAI21_X1 U17653 ( .B1(n15994), .B2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n15763), .ZN(n15915) );
  AOI211_X1 U17654 ( .C1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .C2(n15916), .A(
        n15919), .B(n15915), .ZN(n15764) );
  XNOR2_X1 U17655 ( .A(n15764), .B(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n21376) );
  INV_X1 U17656 ( .A(n21594), .ZN(n15768) );
  INV_X1 U17657 ( .A(n21597), .ZN(n15766) );
  AOI22_X1 U17658 ( .A1(n20022), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B1(
        n10970), .B2(P1_REIP_REG_21__SCAN_IN), .ZN(n15765) );
  OAI21_X1 U17659 ( .B1(n20028), .B2(n15766), .A(n15765), .ZN(n15767) );
  AOI21_X1 U17660 ( .B1(n15768), .B2(n20009), .A(n15767), .ZN(n15769) );
  OAI21_X1 U17661 ( .B1(n21655), .B2(n21376), .A(n15769), .ZN(P1_U2978) );
  XNOR2_X1 U17662 ( .A(n12469), .B(n15901), .ZN(n15770) );
  XNOR2_X1 U17663 ( .A(n15916), .B(n15770), .ZN(n21367) );
  INV_X1 U17664 ( .A(n21575), .ZN(n15774) );
  INV_X1 U17665 ( .A(n21578), .ZN(n15772) );
  AOI22_X1 U17666 ( .A1(n20022), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B1(
        n10970), .B2(P1_REIP_REG_19__SCAN_IN), .ZN(n15771) );
  OAI21_X1 U17667 ( .B1(n20028), .B2(n15772), .A(n15771), .ZN(n15773) );
  AOI21_X1 U17668 ( .B1(n15774), .B2(n20009), .A(n15773), .ZN(n15775) );
  OAI21_X1 U17669 ( .B1(n21367), .B2(n21655), .A(n15775), .ZN(P1_U2980) );
  XNOR2_X1 U17670 ( .A(n15777), .B(n15776), .ZN(n21354) );
  AOI22_X1 U17671 ( .A1(n20022), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B1(
        n10970), .B2(P1_REIP_REG_18__SCAN_IN), .ZN(n15778) );
  OAI21_X1 U17672 ( .B1(n20028), .B2(n21565), .A(n15778), .ZN(n15779) );
  AOI21_X1 U17673 ( .B1(n21567), .B2(n20009), .A(n15779), .ZN(n15780) );
  OAI21_X1 U17674 ( .B1(n21354), .B2(n21655), .A(n15780), .ZN(P1_U2981) );
  NAND2_X1 U17675 ( .A1(n15881), .A2(n15781), .ZN(n15786) );
  INV_X1 U17676 ( .A(n15995), .ZN(n19992) );
  NAND2_X1 U17677 ( .A1(n19992), .A2(n15930), .ZN(n15961) );
  INV_X1 U17678 ( .A(n15782), .ZN(n15783) );
  AOI21_X1 U17679 ( .B1(n15961), .B2(n15784), .A(n15783), .ZN(n15785) );
  MUX2_X1 U17680 ( .A(n15786), .B(n15933), .S(n15785), .Z(n15787) );
  INV_X1 U17681 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15808) );
  XNOR2_X1 U17682 ( .A(n15787), .B(n15808), .ZN(n21359) );
  INV_X1 U17683 ( .A(n15788), .ZN(n15790) );
  AOI22_X1 U17684 ( .A1(n20022), .A2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B1(
        n10970), .B2(P1_REIP_REG_17__SCAN_IN), .ZN(n15789) );
  OAI21_X1 U17685 ( .B1(n20028), .B2(n15790), .A(n15789), .ZN(n15791) );
  AOI21_X1 U17686 ( .B1(n15792), .B2(n20009), .A(n15791), .ZN(n15793) );
  OAI21_X1 U17687 ( .B1(n21359), .B2(n21655), .A(n15793), .ZN(P1_U2982) );
  NAND2_X1 U17688 ( .A1(n15881), .A2(n15794), .ZN(n15959) );
  INV_X1 U17689 ( .A(n15795), .ZN(n15796) );
  AOI21_X1 U17690 ( .B1(n15995), .B2(n15959), .A(n15796), .ZN(n15979) );
  AND2_X1 U17691 ( .A1(n15797), .A2(n15798), .ZN(n15978) );
  NAND2_X1 U17692 ( .A1(n15979), .A2(n15978), .ZN(n15977) );
  NAND2_X1 U17693 ( .A1(n15977), .A2(n15798), .ZN(n15799) );
  XOR2_X1 U17694 ( .A(n15800), .B(n15799), .Z(n21333) );
  INV_X1 U17695 ( .A(n21530), .ZN(n15802) );
  AOI22_X1 U17696 ( .A1(n20022), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .B1(
        n10970), .B2(P1_REIP_REG_13__SCAN_IN), .ZN(n15801) );
  OAI21_X1 U17697 ( .B1(n20028), .B2(n15802), .A(n15801), .ZN(n15803) );
  AOI21_X1 U17698 ( .B1(n15804), .B2(n20009), .A(n15803), .ZN(n15805) );
  OAI21_X1 U17699 ( .B1(n21333), .B2(n21655), .A(n15805), .ZN(P1_U2986) );
  NOR2_X1 U17700 ( .A1(n15806), .A2(n21352), .ZN(n15831) );
  INV_X1 U17701 ( .A(n15826), .ZN(n15816) );
  NAND2_X1 U17702 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n16000) );
  NOR2_X1 U17703 ( .A1(n15807), .A2(n16000), .ZN(n15983) );
  NAND3_X1 U17704 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A3(n15983), .ZN(n21328) );
  INV_X1 U17705 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n21337) );
  NOR4_X1 U17706 ( .A1(n15808), .A2(n21337), .A3(n12581), .A4(n15899), .ZN(
        n21350) );
  NAND2_X1 U17707 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n21350), .ZN(
        n15810) );
  NOR2_X1 U17708 ( .A1(n21328), .A2(n15810), .ZN(n15902) );
  NAND4_X1 U17709 ( .A1(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A4(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15813) );
  INV_X1 U17710 ( .A(n15813), .ZN(n15809) );
  NAND2_X1 U17711 ( .A1(n15902), .A2(n15809), .ZN(n15824) );
  INV_X1 U17712 ( .A(n15810), .ZN(n15812) );
  NOR2_X1 U17713 ( .A1(n16000), .A2(n15811), .ZN(n15920) );
  NAND2_X1 U17714 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n15920), .ZN(
        n15986) );
  NOR2_X1 U17715 ( .A1(n15988), .A2(n15986), .ZN(n15937) );
  NAND2_X1 U17716 ( .A1(n15812), .A2(n15937), .ZN(n15905) );
  NOR2_X1 U17717 ( .A1(n15813), .A2(n15905), .ZN(n15825) );
  AOI21_X1 U17718 ( .B1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n15825), .A(
        n21413), .ZN(n15814) );
  AOI211_X1 U17719 ( .C1(n15938), .C2(n15824), .A(n15814), .B(n15903), .ZN(
        n15887) );
  AOI22_X1 U17720 ( .A1(n15970), .A2(n15872), .B1(n15987), .B2(n15885), .ZN(
        n15815) );
  OAI211_X1 U17721 ( .C1(n15816), .C2(n15967), .A(n15887), .B(n15815), .ZN(
        n15817) );
  NOR2_X1 U17722 ( .A1(n15820), .A2(n15817), .ZN(n15819) );
  INV_X1 U17723 ( .A(n15817), .ZN(n21399) );
  NAND2_X1 U17724 ( .A1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n21399), .ZN(
        n15873) );
  NOR2_X1 U17725 ( .A1(n21398), .A2(n15873), .ZN(n15834) );
  NOR2_X1 U17726 ( .A1(n15819), .A2(n15834), .ZN(n21390) );
  INV_X1 U17727 ( .A(n21390), .ZN(n15818) );
  NAND2_X1 U17728 ( .A1(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n15818), .ZN(
        n15840) );
  INV_X1 U17729 ( .A(n15819), .ZN(n15835) );
  OAI21_X1 U17730 ( .B1(n15836), .B2(n15840), .A(n15835), .ZN(n15822) );
  NAND2_X1 U17731 ( .A1(n15820), .A2(n15850), .ZN(n15839) );
  AOI21_X1 U17732 ( .B1(n15822), .B2(n15839), .A(n15821), .ZN(n15830) );
  NOR2_X1 U17733 ( .A1(n15824), .A2(n15823), .ZN(n15888) );
  AOI21_X1 U17734 ( .B1(n15825), .B2(n15987), .A(n15888), .ZN(n21406) );
  NOR2_X1 U17735 ( .A1(n21406), .A2(n15826), .ZN(n15874) );
  NAND2_X1 U17736 ( .A1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n15874), .ZN(
        n15859) );
  OR2_X1 U17737 ( .A1(n15859), .A2(n15827), .ZN(n15843) );
  NOR3_X1 U17738 ( .A1(n15843), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n15838), .ZN(n15828) );
  NOR4_X1 U17739 ( .A1(n15831), .A2(n15830), .A3(n15829), .A4(n15828), .ZN(
        n15832) );
  OAI21_X1 U17740 ( .B1(n15833), .B2(n21353), .A(n15832), .ZN(P1_U3000) );
  INV_X1 U17741 ( .A(n15834), .ZN(n15837) );
  OAI21_X1 U17742 ( .B1(n15837), .B2(n15836), .A(n15835), .ZN(n15849) );
  AOI21_X1 U17743 ( .B1(n15849), .B2(n15839), .A(n15838), .ZN(n15845) );
  INV_X1 U17744 ( .A(n15840), .ZN(n15842) );
  OAI21_X1 U17745 ( .B1(n15843), .B2(n15842), .A(n15841), .ZN(n15844) );
  AOI211_X1 U17746 ( .C1(n15846), .C2(n21409), .A(n15845), .B(n15844), .ZN(
        n15847) );
  OAI21_X1 U17747 ( .B1(n15848), .B2(n21353), .A(n15847), .ZN(P1_U3001) );
  INV_X1 U17748 ( .A(n15849), .ZN(n15855) );
  INV_X1 U17749 ( .A(n15859), .ZN(n21389) );
  NAND3_X1 U17750 ( .A1(n21389), .A2(n15860), .A3(n15850), .ZN(n15851) );
  OAI211_X1 U17751 ( .C1(n15853), .C2(n21352), .A(n15852), .B(n15851), .ZN(
        n15854) );
  AOI21_X1 U17752 ( .B1(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n15855), .A(
        n15854), .ZN(n15856) );
  OAI21_X1 U17753 ( .B1(n15857), .B2(n21353), .A(n15856), .ZN(P1_U3002) );
  INV_X1 U17754 ( .A(n15858), .ZN(n15862) );
  NOR2_X1 U17755 ( .A1(n15860), .A2(n15859), .ZN(n15861) );
  AOI22_X1 U17756 ( .A1(n15862), .A2(n15861), .B1(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n21390), .ZN(n15863) );
  NAND2_X1 U17757 ( .A1(n15864), .A2(n15863), .ZN(n15865) );
  AOI21_X1 U17758 ( .B1(n15866), .B2(n21409), .A(n15865), .ZN(n15867) );
  OAI21_X1 U17759 ( .B1(n15868), .B2(n21353), .A(n15867), .ZN(P1_U3003) );
  INV_X1 U17760 ( .A(n15869), .ZN(n15870) );
  XNOR2_X1 U17761 ( .A(n15871), .B(n15870), .ZN(n21647) );
  NOR3_X1 U17762 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n21406), .A3(
        n15872), .ZN(n21393) );
  OAI22_X1 U17763 ( .A1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n15874), .B1(
        n21393), .B2(n15873), .ZN(n15876) );
  OAI211_X1 U17764 ( .C1(n21647), .C2(n21352), .A(n15876), .B(n15875), .ZN(
        n15877) );
  INV_X1 U17765 ( .A(n15877), .ZN(n15878) );
  OAI21_X1 U17766 ( .B1(n15879), .B2(n21353), .A(n15878), .ZN(P1_U3005) );
  NAND3_X1 U17767 ( .A1(n15880), .A2(n15994), .A3(n15889), .ZN(n15884) );
  NAND3_X1 U17768 ( .A1(n15882), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        n15881), .ZN(n15883) );
  NAND2_X1 U17769 ( .A1(n15884), .A2(n15883), .ZN(n15886) );
  XNOR2_X1 U17770 ( .A(n15886), .B(n15885), .ZN(n20023) );
  INV_X1 U17771 ( .A(n20023), .ZN(n15895) );
  INV_X1 U17772 ( .A(n15887), .ZN(n21400) );
  OAI221_X1 U17773 ( .B1(n21400), .B2(n15888), .C1(n21400), .C2(n15889), .A(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15894) );
  NOR3_X1 U17774 ( .A1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n21406), .A3(
        n15889), .ZN(n15891) );
  INV_X1 U17775 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n19915) );
  NOR2_X1 U17776 ( .A1(n21386), .A2(n19915), .ZN(n15890) );
  AOI211_X1 U17777 ( .C1(n15892), .C2(n21409), .A(n15891), .B(n15890), .ZN(
        n15893) );
  OAI211_X1 U17778 ( .C1(n15895), .C2(n21353), .A(n15894), .B(n15893), .ZN(
        P1_U3007) );
  NAND2_X1 U17779 ( .A1(n15897), .A2(n15896), .ZN(n15898) );
  XNOR2_X1 U17780 ( .A(n15898), .B(n15908), .ZN(n20017) );
  AOI22_X1 U17781 ( .A1(n15987), .A2(n15920), .B1(n15983), .B2(n15981), .ZN(
        n21343) );
  NAND3_X1 U17782 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15966) );
  NOR2_X1 U17783 ( .A1(n21343), .A2(n15966), .ZN(n15971) );
  NAND2_X1 U17784 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n15971), .ZN(
        n15955) );
  NOR2_X1 U17785 ( .A1(n15899), .A2(n15955), .ZN(n21363) );
  NAND2_X1 U17786 ( .A1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n21363), .ZN(
        n21358) );
  NOR2_X1 U17787 ( .A1(n12468), .A2(n21358), .ZN(n21372) );
  NAND4_X1 U17788 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(n21372), .A4(n15900), .ZN(
        n21378) );
  INV_X1 U17789 ( .A(n21378), .ZN(n15907) );
  NOR2_X1 U17790 ( .A1(n15917), .A2(n15901), .ZN(n15906) );
  NOR2_X1 U17791 ( .A1(n15984), .A2(n15902), .ZN(n15904) );
  AOI211_X1 U17792 ( .C1(n15987), .C2(n15905), .A(n15904), .B(n15903), .ZN(
        n21370) );
  AOI22_X1 U17793 ( .A1(n15906), .A2(n21370), .B1(n21351), .B2(n15982), .ZN(
        n21375) );
  OAI21_X1 U17794 ( .B1(n15907), .B2(n21375), .A(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15914) );
  INV_X1 U17795 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n21615) );
  OAI22_X1 U17796 ( .A1(n21604), .A2(n21352), .B1(n21615), .B2(n21386), .ZN(
        n15912) );
  NAND2_X1 U17797 ( .A1(n15909), .A2(n15908), .ZN(n15910) );
  NOR2_X1 U17798 ( .A1(n21358), .A2(n15910), .ZN(n15911) );
  NOR2_X1 U17799 ( .A1(n15912), .A2(n15911), .ZN(n15913) );
  OAI211_X1 U17800 ( .C1(n20017), .C2(n21353), .A(n15914), .B(n15913), .ZN(
        P1_U3009) );
  AOI21_X1 U17801 ( .B1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n15916), .A(
        n15915), .ZN(n15918) );
  XNOR2_X1 U17802 ( .A(n15918), .B(n15917), .ZN(n20013) );
  AOI22_X1 U17803 ( .A1(n10970), .A2(P1_REIP_REG_20__SCAN_IN), .B1(n21372), 
        .B2(n15919), .ZN(n15926) );
  AND2_X1 U17804 ( .A1(n15987), .A2(n15920), .ZN(n15923) );
  INV_X1 U17805 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n21347) );
  NOR2_X1 U17806 ( .A1(n15988), .A2(n21347), .ZN(n15922) );
  NOR3_X1 U17807 ( .A1(n21658), .A2(n21412), .A3(n21328), .ZN(n15921) );
  AOI21_X1 U17808 ( .B1(n15923), .B2(n15922), .A(n15921), .ZN(n15965) );
  OAI221_X1 U17809 ( .B1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n15965), 
        .C1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n15967), .A(n21370), .ZN(
        n15924) );
  NAND2_X1 U17810 ( .A1(n15924), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15925) );
  OAI211_X1 U17811 ( .C1(n21583), .C2(n21352), .A(n15926), .B(n15925), .ZN(
        n15927) );
  AOI21_X1 U17812 ( .B1(n20013), .B2(n21410), .A(n15927), .ZN(n15928) );
  INV_X1 U17813 ( .A(n15928), .ZN(P1_U3011) );
  XNOR2_X1 U17814 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .B(
        P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15944) );
  NAND3_X1 U17815 ( .A1(n15931), .A2(n15930), .A3(n15929), .ZN(n15946) );
  MUX2_X1 U17816 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B(n15932), .S(
        n15881), .Z(n15947) );
  NOR2_X1 U17817 ( .A1(n15946), .A2(n15947), .ZN(n15945) );
  AOI21_X1 U17818 ( .B1(n15932), .B2(n15881), .A(n15945), .ZN(n15936) );
  INV_X1 U17819 ( .A(n15933), .ZN(n15934) );
  AOI21_X1 U17820 ( .B1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n15881), .A(
        n15934), .ZN(n15935) );
  XNOR2_X1 U17821 ( .A(n15936), .B(n15935), .ZN(n20010) );
  NAND2_X1 U17822 ( .A1(n20010), .A2(n21410), .ZN(n15943) );
  NOR2_X1 U17823 ( .A1(n21337), .A2(n12581), .ZN(n15939) );
  OAI21_X1 U17824 ( .B1(n15937), .B2(n21413), .A(n15982), .ZN(n15969) );
  AOI21_X1 U17825 ( .B1(n15938), .B2(n21328), .A(n15969), .ZN(n21349) );
  OAI21_X1 U17826 ( .B1(n21351), .B2(n15939), .A(n21349), .ZN(n15954) );
  INV_X1 U17827 ( .A(P1_REIP_REG_16__SCAN_IN), .ZN(n15940) );
  OAI22_X1 U17828 ( .A1(n21558), .A2(n21352), .B1(n21386), .B2(n15940), .ZN(
        n15941) );
  AOI21_X1 U17829 ( .B1(n15954), .B2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n15941), .ZN(n15942) );
  OAI211_X1 U17830 ( .C1(n15944), .C2(n15955), .A(n15943), .B(n15942), .ZN(
        P1_U3015) );
  AOI21_X1 U17831 ( .B1(n15947), .B2(n15946), .A(n15945), .ZN(n20008) );
  INV_X1 U17832 ( .A(n15973), .ZN(n15948) );
  NOR2_X1 U17833 ( .A1(n15974), .A2(n15948), .ZN(n15951) );
  INV_X1 U17834 ( .A(n15949), .ZN(n15950) );
  OAI21_X1 U17835 ( .B1(n15952), .B2(n15951), .A(n15950), .ZN(n19959) );
  OAI22_X1 U17836 ( .A1(n19959), .A2(n21352), .B1(n21386), .B2(n19904), .ZN(
        n15953) );
  AOI21_X1 U17837 ( .B1(n15954), .B2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n15953), .ZN(n15958) );
  INV_X1 U17838 ( .A(n15955), .ZN(n15956) );
  NAND2_X1 U17839 ( .A1(n15956), .A2(n15932), .ZN(n15957) );
  OAI211_X1 U17840 ( .C1(n20008), .C2(n21353), .A(n15958), .B(n15957), .ZN(
        P1_U3016) );
  MUX2_X1 U17841 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B(n12581), .S(
        n15881), .Z(n15964) );
  NAND3_X1 U17842 ( .A1(n15961), .A2(n15960), .A3(n15959), .ZN(n15962) );
  OAI21_X1 U17843 ( .B1(n21337), .B2(n12469), .A(n15962), .ZN(n15963) );
  XOR2_X1 U17844 ( .A(n15964), .B(n15963), .Z(n20004) );
  NOR2_X1 U17845 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n15965), .ZN(
        n21329) );
  INV_X1 U17846 ( .A(n15966), .ZN(n15968) );
  AOI21_X1 U17847 ( .B1(n15983), .B2(n15968), .A(n15967), .ZN(n21331) );
  AOI211_X1 U17848 ( .C1(n15970), .C2(n21328), .A(n21331), .B(n15969), .ZN(
        n21338) );
  NAND2_X1 U17849 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n21338), .ZN(
        n15972) );
  OAI22_X1 U17850 ( .A1(n21329), .A2(n15972), .B1(n15971), .B2(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n15976) );
  XNOR2_X1 U17851 ( .A(n15974), .B(n15973), .ZN(n21533) );
  AOI22_X1 U17852 ( .A1(n21533), .A2(n21409), .B1(n10970), .B2(
        P1_REIP_REG_14__SCAN_IN), .ZN(n15975) );
  OAI211_X1 U17853 ( .C1(n20004), .C2(n21353), .A(n15976), .B(n15975), .ZN(
        P1_U3017) );
  OAI21_X1 U17854 ( .B1(n15979), .B2(n15978), .A(n15977), .ZN(n15980) );
  INV_X1 U17855 ( .A(n15980), .ZN(n20001) );
  OAI21_X1 U17856 ( .B1(n15984), .B2(n15983), .A(n15982), .ZN(n15985) );
  AOI21_X1 U17857 ( .B1(n15987), .B2(n15986), .A(n15985), .ZN(n21348) );
  OAI21_X1 U17858 ( .B1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n15823), .A(
        n21348), .ZN(n15992) );
  NOR2_X1 U17859 ( .A1(n21343), .A2(n21347), .ZN(n15989) );
  AOI22_X1 U17860 ( .A1(n10970), .A2(P1_REIP_REG_12__SCAN_IN), .B1(n15989), 
        .B2(n15988), .ZN(n15990) );
  OAI21_X1 U17861 ( .B1(n21512), .B2(n21352), .A(n15990), .ZN(n15991) );
  AOI21_X1 U17862 ( .B1(n15992), .B2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n15991), .ZN(n15993) );
  OAI21_X1 U17863 ( .B1(n20001), .B2(n21353), .A(n15993), .ZN(P1_U3019) );
  MUX2_X1 U17864 ( .A(n15996), .B(n15995), .S(n15994), .Z(n15998) );
  INV_X1 U17865 ( .A(n15998), .ZN(n15999) );
  OR2_X2 U17866 ( .A1(n15998), .A2(n15997), .ZN(n19994) );
  OAI21_X1 U17867 ( .B1(n15999), .B2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n19994), .ZN(n19991) );
  OAI211_X1 U17868 ( .C1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A(n16001), .B(n16000), .ZN(n16005) );
  INV_X1 U17869 ( .A(P1_REIP_REG_10__SCAN_IN), .ZN(n19897) );
  OAI22_X1 U17870 ( .A1(n21352), .A2(n21492), .B1(n19897), .B2(n21386), .ZN(
        n16002) );
  AOI21_X1 U17871 ( .B1(n16003), .B2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n16002), .ZN(n16004) );
  OAI211_X1 U17872 ( .C1(n19991), .C2(n21353), .A(n16005), .B(n16004), .ZN(
        P1_U3021) );
  NOR2_X1 U17873 ( .A1(n16011), .A2(n13587), .ZN(n16007) );
  AOI22_X1 U17874 ( .A1(n16744), .A2(n11493), .B1(n16007), .B2(n16006), .ZN(
        n16008) );
  OAI21_X1 U17875 ( .B1(n10973), .B2(n16739), .A(n16008), .ZN(n16009) );
  INV_X1 U17876 ( .A(n16009), .ZN(n16747) );
  NOR3_X1 U17877 ( .A1(n16011), .A2(n13587), .A3(n16010), .ZN(n16012) );
  AOI21_X1 U17878 ( .B1(n16014), .B2(n16013), .A(n16012), .ZN(n16015) );
  OAI21_X1 U17879 ( .B1(n16747), .B2(n21666), .A(n16015), .ZN(n16016) );
  MUX2_X1 U17880 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n16016), .S(
        n21661), .Z(P1_U3473) );
  INV_X1 U17881 ( .A(n18119), .ZN(n18133) );
  AOI22_X1 U17882 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n13554), .ZN(n18112) );
  AOI22_X1 U17883 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n18120), .B2(n13554), .ZN(
        n16648) );
  NAND2_X1 U17884 ( .A1(n18112), .A2(n16648), .ZN(n16647) );
  NOR2_X1 U17885 ( .A1(n16039), .A2(n16647), .ZN(n18136) );
  NOR2_X1 U17886 ( .A1(n16641), .A2(n18136), .ZN(n16019) );
  XNOR2_X1 U17887 ( .A(n16019), .B(n18135), .ZN(n16020) );
  NOR4_X1 U17888 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(P2_STATE2_REG_2__SCAN_IN), .A3(P2_STATEBS16_REG_SCAN_IN), .A4(n16719), .ZN(n18261) );
  NAND2_X1 U17889 ( .A1(n16020), .A2(n18493), .ZN(n16037) );
  INV_X1 U17890 ( .A(n21729), .ZN(n18630) );
  INV_X1 U17891 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n18505) );
  OAI21_X1 U17892 ( .B1(P2_STATEBS16_REG_SCAN_IN), .B2(n18630), .A(n18505), 
        .ZN(n16021) );
  OAI21_X1 U17893 ( .B1(n16021), .B2(n16029), .A(n16026), .ZN(n16022) );
  OR2_X1 U17894 ( .A1(n18572), .A2(n18493), .ZN(n16023) );
  INV_X1 U17895 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n19264) );
  NAND2_X1 U17896 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19264), .ZN(n18636) );
  NOR3_X1 U17897 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(n19203), .A3(n18636), 
        .ZN(n18640) );
  OR2_X1 U17898 ( .A1(n16023), .A2(n18640), .ZN(n16024) );
  OAI22_X1 U17899 ( .A1(n16027), .A2(n18486), .B1(n18453), .B2(n18595), .ZN(
        n16032) );
  OAI211_X1 U17900 ( .C1(P2_STATEBS16_REG_SCAN_IN), .C2(n18630), .A(n18090), 
        .B(P2_EBX_REG_31__SCAN_IN), .ZN(n16028) );
  INV_X1 U17901 ( .A(n18457), .ZN(n18504) );
  NOR2_X1 U17902 ( .A1(n18504), .A2(n16030), .ZN(n16031) );
  AOI211_X1 U17903 ( .C1(n18331), .C2(P2_REIP_REG_3__SCAN_IN), .A(n16032), .B(
        n16031), .ZN(n16033) );
  OAI21_X1 U17904 ( .B1(n16034), .B2(n18440), .A(n16033), .ZN(n16035) );
  AOI21_X1 U17905 ( .B1(n14864), .B2(n18509), .A(n16035), .ZN(n16036) );
  OAI211_X1 U17906 ( .C1(n19328), .C2(n18133), .A(n16037), .B(n16036), .ZN(
        P2_U2852) );
  NAND2_X1 U17907 ( .A1(n10964), .A2(n16647), .ZN(n16038) );
  XNOR2_X1 U17908 ( .A(n16039), .B(n16038), .ZN(n16050) );
  INV_X2 U17909 ( .A(n18250), .ZN(n18440) );
  INV_X1 U17910 ( .A(n16040), .ZN(n16043) );
  OAI22_X1 U17911 ( .A1(n16041), .A2(n18486), .B1(n12813), .B2(n18502), .ZN(
        n16042) );
  AOI21_X1 U17912 ( .B1(n18471), .B2(n16043), .A(n16042), .ZN(n16044) );
  OAI21_X1 U17913 ( .B1(n18440), .B2(n13523), .A(n16044), .ZN(n16045) );
  AOI21_X1 U17914 ( .B1(n16046), .B2(n18509), .A(n16045), .ZN(n16048) );
  NAND2_X1 U17915 ( .A1(n18621), .A2(n18510), .ZN(n16047) );
  OAI211_X1 U17916 ( .C1(n19219), .C2(n18133), .A(n16048), .B(n16047), .ZN(
        n16049) );
  AOI21_X1 U17917 ( .B1(n16050), .B2(n18493), .A(n16049), .ZN(n16051) );
  INV_X1 U17918 ( .A(n16051), .ZN(P2_U2853) );
  MUX2_X1 U17919 ( .A(n18508), .B(P2_EBX_REG_31__SCAN_IN), .S(n16111), .Z(
        P2_U2856) );
  AOI22_X1 U17920 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n16062), .B1(
        n13107), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n16056) );
  AOI22_X1 U17921 ( .A1(n16064), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n16068), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n16055) );
  NAND2_X1 U17922 ( .A1(n16056), .A2(n16055), .ZN(n16076) );
  AOI21_X1 U17923 ( .B1(n16063), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A(
        n16070), .ZN(n16060) );
  AOI22_X1 U17924 ( .A1(n16058), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n16057), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n16059) );
  OAI211_X1 U17925 ( .C1(n19150), .C2(n16061), .A(n16060), .B(n16059), .ZN(
        n16075) );
  AOI22_X1 U17926 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n16062), .B1(
        n13107), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n16066) );
  AOI22_X1 U17927 ( .A1(n16064), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n16063), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n16065) );
  NAND2_X1 U17928 ( .A1(n16066), .A2(n16065), .ZN(n16074) );
  AOI22_X1 U17929 ( .A1(n16067), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n10957), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n16072) );
  NAND2_X1 U17930 ( .A1(n16057), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n16071) );
  NAND2_X1 U17931 ( .A1(n16068), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n16069) );
  NAND4_X1 U17932 ( .A1(n16072), .A2(n16071), .A3(n16070), .A4(n16069), .ZN(
        n16073) );
  OAI22_X1 U17933 ( .A1(n16076), .A2(n16075), .B1(n16074), .B2(n16073), .ZN(
        n16077) );
  XNOR2_X1 U17934 ( .A(n16078), .B(n16077), .ZN(n16174) );
  NOR2_X1 U17935 ( .A1(n18498), .A2(n16111), .ZN(n16079) );
  AOI21_X1 U17936 ( .B1(P2_EBX_REG_30__SCAN_IN), .B2(n16157), .A(n16079), .ZN(
        n16080) );
  OAI21_X1 U17937 ( .B1(n16174), .B2(n16167), .A(n16080), .ZN(P2_U2857) );
  AND2_X1 U17938 ( .A1(n16090), .A2(n16081), .ZN(n16083) );
  NOR2_X1 U17939 ( .A1(n18474), .A2(n16111), .ZN(n16084) );
  AOI21_X1 U17940 ( .B1(P2_EBX_REG_29__SCAN_IN), .B2(n16157), .A(n16084), .ZN(
        n16085) );
  OAI21_X1 U17941 ( .B1(n16086), .B2(n16167), .A(n16085), .ZN(P2_U2858) );
  NAND2_X1 U17942 ( .A1(n16096), .A2(n16087), .ZN(n16089) );
  XNOR2_X1 U17943 ( .A(n16089), .B(n16088), .ZN(n16185) );
  NAND2_X1 U17944 ( .A1(n16111), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n16094) );
  INV_X1 U17945 ( .A(n16090), .ZN(n16091) );
  AOI21_X1 U17946 ( .B1(n16092), .B2(n16099), .A(n16091), .ZN(n18460) );
  NAND2_X1 U17947 ( .A1(n18460), .A2(n16102), .ZN(n16093) );
  OAI211_X1 U17948 ( .C1(n16185), .C2(n16167), .A(n16094), .B(n16093), .ZN(
        P2_U2859) );
  NAND2_X1 U17949 ( .A1(n16096), .A2(n16095), .ZN(n16097) );
  XOR2_X1 U17950 ( .A(n16098), .B(n16097), .Z(n16194) );
  NAND2_X1 U17951 ( .A1(n16157), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n16104) );
  INV_X1 U17952 ( .A(n16099), .ZN(n16100) );
  AOI21_X1 U17953 ( .B1(n16101), .B2(n16105), .A(n16100), .ZN(n18445) );
  NAND2_X1 U17954 ( .A1(n18445), .A2(n16102), .ZN(n16103) );
  OAI211_X1 U17955 ( .C1(n16194), .C2(n16167), .A(n16104), .B(n16103), .ZN(
        P2_U2860) );
  OAI21_X1 U17956 ( .B1(n16107), .B2(n16106), .A(n16105), .ZN(n16294) );
  AOI21_X1 U17957 ( .B1(n16110), .B2(n16109), .A(n16108), .ZN(n16195) );
  NAND2_X1 U17958 ( .A1(n16195), .A2(n16141), .ZN(n16113) );
  NAND2_X1 U17959 ( .A1(n16111), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n16112) );
  OAI211_X1 U17960 ( .C1(n16294), .C2(n16157), .A(n16113), .B(n16112), .ZN(
        P2_U2861) );
  OAI21_X1 U17961 ( .B1(n16116), .B2(n16115), .A(n16114), .ZN(n16209) );
  NOR2_X1 U17962 ( .A1(n16117), .A2(n16111), .ZN(n16118) );
  AOI21_X1 U17963 ( .B1(P2_EBX_REG_25__SCAN_IN), .B2(n16157), .A(n16118), .ZN(
        n16119) );
  OAI21_X1 U17964 ( .B1(n16209), .B2(n16167), .A(n16119), .ZN(P2_U2862) );
  OAI21_X1 U17965 ( .B1(n16122), .B2(n16121), .A(n16120), .ZN(n16217) );
  NOR2_X1 U17966 ( .A1(n16123), .A2(n16111), .ZN(n16124) );
  AOI21_X1 U17967 ( .B1(P2_EBX_REG_24__SCAN_IN), .B2(n16157), .A(n16124), .ZN(
        n16125) );
  OAI21_X1 U17968 ( .B1(n16217), .B2(n16167), .A(n16125), .ZN(P2_U2863) );
  XNOR2_X1 U17969 ( .A(n16126), .B(n16127), .ZN(n16224) );
  NOR2_X1 U17970 ( .A1(n16128), .A2(n16111), .ZN(n16129) );
  AOI21_X1 U17971 ( .B1(P2_EBX_REG_23__SCAN_IN), .B2(n16157), .A(n16129), .ZN(
        n16130) );
  OAI21_X1 U17972 ( .B1(n16224), .B2(n16167), .A(n16130), .ZN(P2_U2864) );
  OAI21_X1 U17973 ( .B1(n16139), .B2(n16132), .A(n16126), .ZN(n19350) );
  NOR2_X1 U17974 ( .A1(n16133), .A2(n16111), .ZN(n16134) );
  AOI21_X1 U17975 ( .B1(P2_EBX_REG_22__SCAN_IN), .B2(n16157), .A(n16134), .ZN(
        n16135) );
  OAI21_X1 U17976 ( .B1(n19350), .B2(n16167), .A(n16135), .ZN(P2_U2865) );
  AND2_X1 U17977 ( .A1(n16148), .A2(n16136), .ZN(n16138) );
  OR2_X1 U17978 ( .A1(n16138), .A2(n16137), .ZN(n16321) );
  AOI21_X1 U17979 ( .B1(n16140), .B2(n16144), .A(n16139), .ZN(n16225) );
  NAND2_X1 U17980 ( .A1(n16225), .A2(n16141), .ZN(n16143) );
  NAND2_X1 U17981 ( .A1(n16111), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n16142) );
  OAI211_X1 U17982 ( .C1(n16321), .C2(n16157), .A(n16143), .B(n16142), .ZN(
        P2_U2866) );
  OAI21_X1 U17983 ( .B1(n11040), .B2(n16145), .A(n16144), .ZN(n19454) );
  NAND2_X1 U17984 ( .A1(n16154), .A2(n16146), .ZN(n16147) );
  NAND2_X1 U17985 ( .A1(n16148), .A2(n16147), .ZN(n16333) );
  NOR2_X1 U17986 ( .A1(n16333), .A2(n16157), .ZN(n16149) );
  AOI21_X1 U17987 ( .B1(P2_EBX_REG_20__SCAN_IN), .B2(n16157), .A(n16149), .ZN(
        n16150) );
  OAI21_X1 U17988 ( .B1(n19454), .B2(n16167), .A(n16150), .ZN(P2_U2867) );
  AOI21_X1 U17989 ( .B1(n16152), .B2(n16151), .A(n11040), .ZN(n16153) );
  INV_X1 U17990 ( .A(n16153), .ZN(n16248) );
  OAI21_X1 U17991 ( .B1(n16163), .B2(n16155), .A(n16154), .ZN(n16491) );
  NOR2_X1 U17992 ( .A1(n16491), .A2(n16111), .ZN(n16156) );
  AOI21_X1 U17993 ( .B1(P2_EBX_REG_19__SCAN_IN), .B2(n16157), .A(n16156), .ZN(
        n16158) );
  OAI21_X1 U17994 ( .B1(n16248), .B2(n16167), .A(n16158), .ZN(P2_U2868) );
  OAI21_X1 U17995 ( .B1(n16160), .B2(n16159), .A(n16151), .ZN(n19546) );
  AND2_X1 U17996 ( .A1(n16162), .A2(n16161), .ZN(n16164) );
  OR2_X1 U17997 ( .A1(n16164), .A2(n16163), .ZN(n18321) );
  NOR2_X1 U17998 ( .A1(n18321), .A2(n16111), .ZN(n16165) );
  AOI21_X1 U17999 ( .B1(P2_EBX_REG_18__SCAN_IN), .B2(n16157), .A(n16165), .ZN(
        n16166) );
  OAI21_X1 U18000 ( .B1(n19546), .B2(n16167), .A(n16166), .ZN(P2_U2869) );
  INV_X1 U18001 ( .A(n19119), .ZN(n16171) );
  INV_X1 U18002 ( .A(n18491), .ZN(n16169) );
  OAI22_X1 U18003 ( .A1(n19658), .A2(n16169), .B1(n16168), .B2(n19401), .ZN(
        n16170) );
  AOI21_X1 U18004 ( .B1(n19653), .B2(n16171), .A(n16170), .ZN(n16173) );
  AOI22_X1 U18005 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n19654), .B1(n19655), .B2(
        BUF2_REG_30__SCAN_IN), .ZN(n16172) );
  OAI211_X1 U18006 ( .C1(n16174), .C2(n19659), .A(n16173), .B(n16172), .ZN(
        P2_U2889) );
  INV_X1 U18007 ( .A(n19125), .ZN(n16182) );
  INV_X1 U18008 ( .A(n16175), .ZN(n16178) );
  INV_X1 U18009 ( .A(n16187), .ZN(n16177) );
  AOI21_X1 U18010 ( .B1(n16178), .B2(n16177), .A(n16176), .ZN(n18459) );
  INV_X1 U18011 ( .A(n18459), .ZN(n16180) );
  OAI22_X1 U18012 ( .A1(n19658), .A2(n16180), .B1(n16179), .B2(n19401), .ZN(
        n16181) );
  AOI21_X1 U18013 ( .B1(n19653), .B2(n16182), .A(n16181), .ZN(n16184) );
  AOI22_X1 U18014 ( .A1(n19654), .A2(BUF1_REG_28__SCAN_IN), .B1(n19655), .B2(
        BUF2_REG_28__SCAN_IN), .ZN(n16183) );
  OAI211_X1 U18015 ( .C1(n16185), .C2(n19659), .A(n16184), .B(n16183), .ZN(
        P2_U2891) );
  INV_X1 U18016 ( .A(n19128), .ZN(n16191) );
  AND2_X1 U18017 ( .A1(n16196), .A2(n16186), .ZN(n16188) );
  OR2_X1 U18018 ( .A1(n16188), .A2(n16187), .ZN(n18452) );
  OAI22_X1 U18019 ( .A1(n19658), .A2(n18452), .B1(n16189), .B2(n19401), .ZN(
        n16190) );
  AOI21_X1 U18020 ( .B1(n19653), .B2(n16191), .A(n16190), .ZN(n16193) );
  AOI22_X1 U18021 ( .A1(n19654), .A2(BUF1_REG_27__SCAN_IN), .B1(n19655), .B2(
        BUF2_REG_27__SCAN_IN), .ZN(n16192) );
  OAI211_X1 U18022 ( .C1(n16194), .C2(n19659), .A(n16193), .B(n16192), .ZN(
        P2_U2892) );
  NAND2_X1 U18023 ( .A1(n16195), .A2(n19549), .ZN(n16203) );
  INV_X1 U18024 ( .A(n16196), .ZN(n16197) );
  AOI21_X1 U18025 ( .B1(n16199), .B2(n16198), .A(n16197), .ZN(n18429) );
  AOI22_X1 U18026 ( .A1(n19548), .A2(n18429), .B1(P2_EAX_REG_26__SCAN_IN), 
        .B2(n19652), .ZN(n16202) );
  AOI22_X1 U18027 ( .A1(n19654), .A2(BUF1_REG_26__SCAN_IN), .B1(n19655), .B2(
        BUF2_REG_26__SCAN_IN), .ZN(n16201) );
  NAND2_X1 U18028 ( .A1(n19653), .A2(n19129), .ZN(n16200) );
  NAND4_X1 U18029 ( .A1(n16203), .A2(n16202), .A3(n16201), .A4(n16200), .ZN(
        P2_U2893) );
  INV_X1 U18030 ( .A(n19135), .ZN(n16206) );
  OAI22_X1 U18031 ( .A1(n19658), .A2(n18414), .B1(n16204), .B2(n19401), .ZN(
        n16205) );
  AOI21_X1 U18032 ( .B1(n19653), .B2(n16206), .A(n16205), .ZN(n16208) );
  AOI22_X1 U18033 ( .A1(n19654), .A2(BUF1_REG_25__SCAN_IN), .B1(n19655), .B2(
        BUF2_REG_25__SCAN_IN), .ZN(n16207) );
  OAI211_X1 U18034 ( .C1(n16209), .C2(n19659), .A(n16208), .B(n16207), .ZN(
        P2_U2894) );
  INV_X1 U18035 ( .A(n19138), .ZN(n16215) );
  INV_X1 U18036 ( .A(n18400), .ZN(n16211) );
  OAI22_X1 U18037 ( .A1(n19658), .A2(n16211), .B1(n16210), .B2(n19401), .ZN(
        n16214) );
  INV_X1 U18038 ( .A(n19654), .ZN(n16243) );
  INV_X1 U18039 ( .A(n19655), .ZN(n16242) );
  INV_X1 U18040 ( .A(BUF2_REG_24__SCAN_IN), .ZN(n16212) );
  OAI22_X1 U18041 ( .A1(n16243), .A2(n20084), .B1(n16242), .B2(n16212), .ZN(
        n16213) );
  AOI211_X1 U18042 ( .C1(n19653), .C2(n16215), .A(n16214), .B(n16213), .ZN(
        n16216) );
  OAI21_X1 U18043 ( .B1(n16217), .B2(n19659), .A(n16216), .ZN(P2_U2895) );
  INV_X1 U18044 ( .A(n19146), .ZN(n16222) );
  OAI22_X1 U18045 ( .A1(n19658), .A2(n18395), .B1(n16218), .B2(n19401), .ZN(
        n16221) );
  INV_X1 U18046 ( .A(BUF2_REG_23__SCAN_IN), .ZN(n16219) );
  OAI22_X1 U18047 ( .A1(n16243), .A2(n20082), .B1(n16242), .B2(n16219), .ZN(
        n16220) );
  AOI211_X1 U18048 ( .C1(n19653), .C2(n16222), .A(n16221), .B(n16220), .ZN(
        n16223) );
  OAI21_X1 U18049 ( .B1(n16224), .B2(n19659), .A(n16223), .ZN(P2_U2896) );
  INV_X1 U18050 ( .A(n16225), .ZN(n16237) );
  AOI22_X1 U18051 ( .A1(n16679), .A2(BUF1_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n16226), .ZN(n19413) );
  INV_X1 U18052 ( .A(n19413), .ZN(n16235) );
  OR2_X1 U18053 ( .A1(n16478), .A2(n16227), .ZN(n16229) );
  AND2_X1 U18054 ( .A1(n16229), .A2(n16228), .ZN(n18362) );
  INV_X1 U18055 ( .A(n18362), .ZN(n16231) );
  OAI22_X1 U18056 ( .A1(n19658), .A2(n16231), .B1(n16230), .B2(n19401), .ZN(
        n16234) );
  INV_X1 U18057 ( .A(BUF2_REG_21__SCAN_IN), .ZN(n16232) );
  OAI22_X1 U18058 ( .A1(n16243), .A2(n20077), .B1(n16242), .B2(n16232), .ZN(
        n16233) );
  AOI211_X1 U18059 ( .C1(n19653), .C2(n16235), .A(n16234), .B(n16233), .ZN(
        n16236) );
  OAI21_X1 U18060 ( .B1(n16237), .B2(n19659), .A(n16236), .ZN(P2_U2898) );
  AND2_X1 U18061 ( .A1(n11008), .A2(n16238), .ZN(n16239) );
  NOR2_X1 U18062 ( .A1(n16477), .A2(n16239), .ZN(n18336) );
  INV_X1 U18063 ( .A(n18336), .ZN(n16496) );
  OAI22_X1 U18064 ( .A1(n19658), .A2(n16496), .B1(n16240), .B2(n19401), .ZN(
        n16245) );
  INV_X1 U18065 ( .A(BUF2_REG_19__SCAN_IN), .ZN(n16241) );
  OAI22_X1 U18066 ( .A1(n16243), .A2(n20073), .B1(n16242), .B2(n16241), .ZN(
        n16244) );
  AOI211_X1 U18067 ( .C1(n19653), .C2(n16246), .A(n16245), .B(n16244), .ZN(
        n16247) );
  OAI21_X1 U18068 ( .B1(n16248), .B2(n19659), .A(n16247), .ZN(P2_U2900) );
  XNOR2_X1 U18069 ( .A(n16263), .B(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n18494) );
  NOR2_X1 U18070 ( .A1(n18494), .A2(n17046), .ZN(n16249) );
  AOI211_X1 U18071 ( .C1(n17052), .C2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n16250), .B(n16249), .ZN(n16251) );
  OAI21_X1 U18072 ( .B1(n18498), .B2(n17062), .A(n16251), .ZN(n16252) );
  AOI21_X1 U18073 ( .B1(n16253), .B2(n17047), .A(n16252), .ZN(n16254) );
  OAI21_X1 U18074 ( .B1(n16255), .B2(n17058), .A(n16254), .ZN(P2_U2984) );
  NOR2_X1 U18075 ( .A1(n16257), .A2(n16256), .ZN(n16259) );
  XOR2_X1 U18076 ( .A(n16259), .B(n16258), .Z(n16422) );
  INV_X1 U18077 ( .A(n16260), .ZN(n16262) );
  AOI21_X1 U18078 ( .B1(n16286), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16261) );
  NOR2_X1 U18079 ( .A1(n16262), .A2(n16261), .ZN(n16420) );
  AOI21_X1 U18080 ( .B1(n16264), .B2(n11068), .A(n16263), .ZN(n18478) );
  NAND2_X1 U18081 ( .A1(n18572), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n16414) );
  OAI21_X1 U18082 ( .B1(n17022), .B2(n16264), .A(n16414), .ZN(n16265) );
  AOI21_X1 U18083 ( .B1(n18478), .B2(n17055), .A(n16265), .ZN(n16266) );
  OAI21_X1 U18084 ( .B1(n18474), .B2(n17062), .A(n16266), .ZN(n16267) );
  AOI21_X1 U18085 ( .B1(n16420), .B2(n17047), .A(n16267), .ZN(n16268) );
  OAI21_X1 U18086 ( .B1(n16422), .B2(n17058), .A(n16268), .ZN(P2_U2985) );
  NOR2_X1 U18087 ( .A1(n16270), .A2(n16269), .ZN(n16282) );
  INV_X1 U18088 ( .A(n16271), .ZN(n16272) );
  OAI22_X1 U18089 ( .A1(n16282), .A2(n16272), .B1(n16280), .B2(n16413), .ZN(
        n16275) );
  XNOR2_X1 U18090 ( .A(n16273), .B(n16427), .ZN(n16274) );
  XNOR2_X1 U18091 ( .A(n16275), .B(n16274), .ZN(n16433) );
  OAI21_X1 U18092 ( .B1(n16283), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n11068), .ZN(n18462) );
  NOR2_X1 U18093 ( .A1(n18589), .A2(n18454), .ZN(n16425) );
  AOI21_X1 U18094 ( .B1(n17052), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n16425), .ZN(n16276) );
  OAI21_X1 U18095 ( .B1(n18462), .B2(n17046), .A(n16276), .ZN(n16277) );
  AOI21_X1 U18096 ( .B1(n18460), .B2(n17019), .A(n16277), .ZN(n16279) );
  XNOR2_X1 U18097 ( .A(n16286), .B(n16427), .ZN(n16430) );
  NAND2_X1 U18098 ( .A1(n16430), .A2(n17047), .ZN(n16278) );
  OAI211_X1 U18099 ( .C1(n16433), .C2(n17058), .A(n16279), .B(n16278), .ZN(
        P2_U2986) );
  XNOR2_X1 U18100 ( .A(n16280), .B(n16413), .ZN(n16281) );
  XNOR2_X1 U18101 ( .A(n16282), .B(n16281), .ZN(n16444) );
  AOI21_X1 U18102 ( .B1(n18442), .B2(n11064), .A(n16283), .ZN(n18447) );
  NAND2_X1 U18103 ( .A1(n18447), .A2(n17055), .ZN(n16284) );
  NAND2_X1 U18104 ( .A1(n18572), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n16435) );
  OAI211_X1 U18105 ( .C1(n17022), .C2(n18442), .A(n16284), .B(n16435), .ZN(
        n16285) );
  AOI21_X1 U18106 ( .B1(n18445), .B2(n17019), .A(n16285), .ZN(n16288) );
  AOI21_X1 U18107 ( .B1(n16413), .B2(n16297), .A(n16286), .ZN(n16441) );
  NAND2_X1 U18108 ( .A1(n16441), .A2(n17047), .ZN(n16287) );
  OAI211_X1 U18109 ( .C1(n16444), .C2(n17058), .A(n16288), .B(n16287), .ZN(
        P2_U2987) );
  AOI21_X1 U18110 ( .B1(n16291), .B2(n16290), .A(n16289), .ZN(n16292) );
  XOR2_X1 U18111 ( .A(n16293), .B(n16292), .Z(n16456) );
  INV_X1 U18112 ( .A(n16294), .ZN(n18430) );
  OAI21_X1 U18113 ( .B1(n16295), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n11064), .ZN(n18432) );
  INV_X1 U18114 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n18425) );
  NOR2_X1 U18115 ( .A1(n18589), .A2(n18425), .ZN(n16450) );
  AOI21_X1 U18116 ( .B1(n17052), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n16450), .ZN(n16296) );
  OAI21_X1 U18117 ( .B1(n18432), .B2(n17046), .A(n16296), .ZN(n16300) );
  NOR2_X1 U18118 ( .A1(n16454), .A2(n17042), .ZN(n16299) );
  AOI211_X1 U18119 ( .C1(n17019), .C2(n18430), .A(n16300), .B(n16299), .ZN(
        n16301) );
  OAI21_X1 U18120 ( .B1(n16456), .B2(n17058), .A(n16301), .ZN(P2_U2988) );
  NAND2_X1 U18121 ( .A1(n16305), .A2(n16569), .ZN(n16307) );
  AND2_X1 U18122 ( .A1(n16309), .A2(n16558), .ZN(n16310) );
  NAND2_X1 U18123 ( .A1(n16311), .A2(n16310), .ZN(n16522) );
  INV_X1 U18124 ( .A(n16312), .ZN(n16521) );
  INV_X1 U18125 ( .A(n16362), .ZN(n16314) );
  AND2_X1 U18126 ( .A1(n16342), .A2(n16353), .ZN(n16315) );
  NAND2_X1 U18127 ( .A1(n16316), .A2(n16315), .ZN(n16317) );
  NOR2_X1 U18128 ( .A1(n16317), .A2(n16318), .ZN(n16319) );
  INV_X1 U18129 ( .A(n16319), .ZN(n16320) );
  INV_X1 U18130 ( .A(n16322), .ZN(n16323) );
  AOI21_X1 U18131 ( .B1(n16325), .B2(n16334), .A(n16323), .ZN(n18364) );
  NAND2_X1 U18132 ( .A1(n18364), .A2(n17055), .ZN(n16324) );
  NAND2_X1 U18133 ( .A1(n18572), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n16457) );
  OAI211_X1 U18134 ( .C1(n17022), .C2(n16325), .A(n16324), .B(n16457), .ZN(
        n16330) );
  OAI21_X1 U18135 ( .B1(n16339), .B2(n16475), .A(n16461), .ZN(n16328) );
  NOR2_X1 U18136 ( .A1(n16463), .A2(n17042), .ZN(n16329) );
  AOI211_X1 U18137 ( .C1(n17019), .C2(n18363), .A(n16330), .B(n16329), .ZN(
        n16331) );
  OAI21_X1 U18138 ( .B1(n16465), .B2(n17058), .A(n16331), .ZN(P2_U2993) );
  XNOR2_X1 U18139 ( .A(n16339), .B(n16475), .ZN(n16489) );
  OR2_X1 U18140 ( .A1(n16332), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n16467) );
  NAND3_X1 U18141 ( .A1(n16467), .A2(n16466), .A3(n17039), .ZN(n16338) );
  INV_X1 U18142 ( .A(n16333), .ZN(n18353) );
  OAI21_X1 U18143 ( .B1(n11041), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n16334), .ZN(n18341) );
  NOR2_X1 U18144 ( .A1(n18589), .A2(n18350), .ZN(n16481) );
  AOI21_X1 U18145 ( .B1(n17052), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n16481), .ZN(n16335) );
  OAI21_X1 U18146 ( .B1(n18341), .B2(n17046), .A(n16335), .ZN(n16336) );
  AOI21_X1 U18147 ( .B1(n18353), .B2(n17019), .A(n16336), .ZN(n16337) );
  OAI211_X1 U18148 ( .C1(n16489), .C2(n17042), .A(n16338), .B(n16337), .ZN(
        P2_U2994) );
  OAI21_X1 U18149 ( .B1(n16350), .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n16339), .ZN(n16501) );
  INV_X1 U18150 ( .A(n16353), .ZN(n16340) );
  OAI21_X1 U18151 ( .B1(n16354), .B2(n16340), .A(n16352), .ZN(n16344) );
  NAND2_X1 U18152 ( .A1(n16342), .A2(n16341), .ZN(n16343) );
  XNOR2_X1 U18153 ( .A(n16344), .B(n16343), .ZN(n16490) );
  AOI21_X1 U18154 ( .B1(n16357), .B2(n16345), .A(n11041), .ZN(n18342) );
  NAND2_X1 U18155 ( .A1(n18572), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n16495) );
  OAI21_X1 U18156 ( .B1(n17022), .B2(n16345), .A(n16495), .ZN(n16346) );
  AOI21_X1 U18157 ( .B1(n18342), .B2(n17055), .A(n16346), .ZN(n16347) );
  OAI21_X1 U18158 ( .B1(n16491), .B2(n17062), .A(n16347), .ZN(n16348) );
  AOI21_X1 U18159 ( .B1(n16490), .B2(n17039), .A(n16348), .ZN(n16349) );
  OAI21_X1 U18160 ( .B1(n17042), .B2(n16501), .A(n16349), .ZN(P2_U2995) );
  INV_X1 U18161 ( .A(n16370), .ZN(n16351) );
  OAI21_X1 U18162 ( .B1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n16351), .A(
        n11240), .ZN(n16513) );
  NAND2_X1 U18163 ( .A1(n16353), .A2(n16352), .ZN(n16355) );
  XOR2_X1 U18164 ( .A(n16355), .B(n16354), .Z(n16511) );
  NOR2_X1 U18165 ( .A1(n18589), .A2(n16356), .ZN(n16505) );
  OAI21_X1 U18166 ( .B1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n16366), .A(
        n16357), .ZN(n18326) );
  NOR2_X1 U18167 ( .A1(n18326), .A2(n17046), .ZN(n16358) );
  AOI211_X1 U18168 ( .C1(n17052), .C2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n16505), .B(n16358), .ZN(n16359) );
  OAI21_X1 U18169 ( .B1(n18321), .B2(n17062), .A(n16359), .ZN(n16360) );
  AOI21_X1 U18170 ( .B1(n16511), .B2(n17039), .A(n16360), .ZN(n16361) );
  OAI21_X1 U18171 ( .B1(n17042), .B2(n16513), .A(n16361), .ZN(P2_U2996) );
  NAND2_X1 U18172 ( .A1(n16363), .A2(n16362), .ZN(n16364) );
  XNOR2_X1 U18173 ( .A(n16365), .B(n16364), .ZN(n18559) );
  INV_X1 U18174 ( .A(n18559), .ZN(n16374) );
  AOI21_X1 U18175 ( .B1(n16367), .B2(n17049), .A(n16366), .ZN(n18305) );
  INV_X1 U18176 ( .A(n18305), .ZN(n18314) );
  NAND2_X1 U18177 ( .A1(n18572), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n18563) );
  NAND2_X1 U18178 ( .A1(n17052), .A2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n16368) );
  OAI211_X1 U18179 ( .C1(n18314), .C2(n17046), .A(n18563), .B(n16368), .ZN(
        n16369) );
  AOI21_X1 U18180 ( .B1(n18554), .B2(n17019), .A(n16369), .ZN(n16373) );
  NAND2_X1 U18181 ( .A1(n11013), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n17048) );
  INV_X1 U18182 ( .A(n17048), .ZN(n16371) );
  OAI211_X1 U18183 ( .C1(n16371), .C2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n17047), .B(n16370), .ZN(n16372) );
  OAI211_X1 U18184 ( .C1(n16374), .C2(n17058), .A(n16373), .B(n16372), .ZN(
        P2_U2997) );
  NAND2_X1 U18185 ( .A1(n16375), .A2(n16557), .ZN(n16389) );
  NAND2_X1 U18186 ( .A1(n16389), .A2(n16387), .ZN(n16376) );
  NAND2_X1 U18187 ( .A1(n16376), .A2(n16388), .ZN(n17036) );
  AND2_X1 U18188 ( .A1(n16378), .A2(n16377), .ZN(n17035) );
  NAND2_X1 U18189 ( .A1(n17036), .A2(n17035), .ZN(n17038) );
  NAND2_X1 U18190 ( .A1(n17038), .A2(n16378), .ZN(n16382) );
  NAND2_X1 U18191 ( .A1(n16380), .A2(n16379), .ZN(n16381) );
  XNOR2_X1 U18192 ( .A(n16382), .B(n16381), .ZN(n16537) );
  AOI21_X1 U18193 ( .B1(n18282), .B2(n17031), .A(n17050), .ZN(n18294) );
  NAND2_X1 U18194 ( .A1(n17055), .A2(n18294), .ZN(n16383) );
  NAND2_X1 U18195 ( .A1(n18572), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n16535) );
  OAI211_X1 U18196 ( .C1(n17022), .C2(n18282), .A(n16383), .B(n16535), .ZN(
        n16384) );
  AOI21_X1 U18197 ( .B1(n18286), .B2(n17019), .A(n16384), .ZN(n16386) );
  AOI21_X1 U18198 ( .B1(n16531), .B2(n17033), .A(n11013), .ZN(n16530) );
  NAND2_X1 U18199 ( .A1(n16530), .A2(n17047), .ZN(n16385) );
  OAI211_X1 U18200 ( .C1(n16537), .C2(n17058), .A(n16386), .B(n16385), .ZN(
        P2_U2999) );
  NAND2_X1 U18201 ( .A1(n16600), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n16599) );
  NAND2_X1 U18202 ( .A1(n16582), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n16568) );
  NOR2_X1 U18203 ( .A1(n16568), .A2(n16563), .ZN(n16560) );
  NAND2_X1 U18204 ( .A1(n16600), .A2(n18548), .ZN(n17032) );
  OAI21_X1 U18205 ( .B1(n16560), .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n17032), .ZN(n16556) );
  NAND2_X1 U18206 ( .A1(n16388), .A2(n16387), .ZN(n16390) );
  XOR2_X1 U18207 ( .A(n16390), .B(n16389), .Z(n16554) );
  AOI21_X1 U18208 ( .B1(n17024), .B2(n18265), .A(n11042), .ZN(n18254) );
  OAI22_X1 U18209 ( .A1(n17022), .A2(n18265), .B1(n16391), .B2(n18589), .ZN(
        n16392) );
  AOI21_X1 U18210 ( .B1(n17055), .B2(n18254), .A(n16392), .ZN(n16393) );
  OAI21_X1 U18211 ( .B1(n18259), .B2(n17062), .A(n16393), .ZN(n16394) );
  AOI21_X1 U18212 ( .B1(n16554), .B2(n17039), .A(n16394), .ZN(n16395) );
  OAI21_X1 U18213 ( .B1(n16556), .B2(n17042), .A(n16395), .ZN(P2_U3001) );
  XNOR2_X1 U18214 ( .A(n16397), .B(n16396), .ZN(n16629) );
  NAND2_X1 U18215 ( .A1(n16990), .A2(n16992), .ZN(n16399) );
  XNOR2_X1 U18216 ( .A(n16398), .B(n16399), .ZN(n16627) );
  INV_X1 U18217 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n16400) );
  OAI21_X1 U18218 ( .B1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n16407), .A(
        n16987), .ZN(n18186) );
  OAI22_X1 U18219 ( .A1(n16400), .A2(n17022), .B1(n17046), .B2(n18186), .ZN(
        n16402) );
  OAI22_X1 U18220 ( .A1(n17062), .A2(n18175), .B1(n18589), .B2(n17133), .ZN(
        n16401) );
  AOI211_X1 U18221 ( .C1(n16627), .C2(n17039), .A(n16402), .B(n16401), .ZN(
        n16403) );
  OAI21_X1 U18222 ( .B1(n16629), .B2(n17042), .A(n16403), .ZN(P2_U3007) );
  XNOR2_X1 U18223 ( .A(n16404), .B(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n16639) );
  XOR2_X1 U18224 ( .A(n16406), .B(n16405), .Z(n16637) );
  AOI21_X1 U18225 ( .B1(n18167), .B2(n16978), .A(n16407), .ZN(n18169) );
  OAI22_X1 U18226 ( .A1(n18167), .A2(n17022), .B1(n13834), .B2(n18589), .ZN(
        n16408) );
  AOI21_X1 U18227 ( .B1(n17055), .B2(n18169), .A(n16408), .ZN(n16409) );
  OAI21_X1 U18228 ( .B1(n18161), .B2(n17062), .A(n16409), .ZN(n16410) );
  AOI21_X1 U18229 ( .B1(n16637), .B2(n17039), .A(n16410), .ZN(n16411) );
  OAI21_X1 U18230 ( .B1(n16639), .B2(n17042), .A(n16411), .ZN(P2_U3008) );
  OR2_X1 U18231 ( .A1(n16413), .A2(n16416), .ZN(n16423) );
  XNOR2_X1 U18232 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .B(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16415) );
  OAI21_X1 U18233 ( .B1(n16423), .B2(n16415), .A(n16414), .ZN(n16419) );
  NOR2_X1 U18234 ( .A1(n16416), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n16437) );
  NOR2_X1 U18235 ( .A1(n16434), .A2(n16437), .ZN(n16428) );
  INV_X1 U18236 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16417) );
  NOR2_X1 U18237 ( .A1(n16428), .A2(n16417), .ZN(n16418) );
  OAI21_X1 U18238 ( .B1(n16422), .B2(n18606), .A(n16421), .ZN(P2_U3017) );
  NOR2_X1 U18239 ( .A1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n16423), .ZN(
        n16424) );
  AOI211_X1 U18240 ( .C1(n18622), .C2(n18459), .A(n16425), .B(n16424), .ZN(
        n16426) );
  OAI21_X1 U18241 ( .B1(n16428), .B2(n16427), .A(n16426), .ZN(n16429) );
  AOI21_X1 U18242 ( .B1(n18460), .B2(n18591), .A(n16429), .ZN(n16432) );
  NAND2_X1 U18243 ( .A1(n16430), .A2(n18568), .ZN(n16431) );
  OAI211_X1 U18244 ( .C1(n16433), .C2(n18606), .A(n16432), .B(n16431), .ZN(
        P2_U3018) );
  NAND2_X1 U18245 ( .A1(n16434), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n16439) );
  INV_X1 U18246 ( .A(n16435), .ZN(n16436) );
  NOR2_X1 U18247 ( .A1(n16437), .A2(n16436), .ZN(n16438) );
  OAI211_X1 U18248 ( .C1(n18594), .C2(n18452), .A(n16439), .B(n16438), .ZN(
        n16440) );
  AOI21_X1 U18249 ( .B1(n18445), .B2(n18591), .A(n16440), .ZN(n16443) );
  NAND2_X1 U18250 ( .A1(n16441), .A2(n18568), .ZN(n16442) );
  OAI211_X1 U18251 ( .C1(n16444), .C2(n18606), .A(n16443), .B(n16442), .ZN(
        P2_U3019) );
  INV_X1 U18252 ( .A(n16445), .ZN(n16446) );
  AOI211_X1 U18253 ( .C1(n16448), .C2(n16452), .A(n16447), .B(n16446), .ZN(
        n16449) );
  AOI211_X1 U18254 ( .C1(n18622), .C2(n18429), .A(n16450), .B(n16449), .ZN(
        n16451) );
  OAI21_X1 U18255 ( .B1(n16453), .B2(n16452), .A(n16451), .ZN(n16455) );
  INV_X1 U18256 ( .A(n16457), .ZN(n16459) );
  NOR3_X1 U18257 ( .A1(n16484), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(
        n16475), .ZN(n16458) );
  AOI211_X1 U18258 ( .C1(n18622), .C2(n18362), .A(n16459), .B(n16458), .ZN(
        n16460) );
  OAI21_X1 U18259 ( .B1(n16462), .B2(n16461), .A(n16460), .ZN(n16464) );
  NAND3_X1 U18260 ( .A1(n16467), .A2(n16466), .A3(n18598), .ZN(n16488) );
  NOR2_X1 U18261 ( .A1(n18608), .A2(n16532), .ZN(n16468) );
  NOR2_X1 U18262 ( .A1(n16469), .A2(n16468), .ZN(n16519) );
  NAND3_X1 U18263 ( .A1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n16471) );
  INV_X1 U18264 ( .A(n16616), .ZN(n18614) );
  NAND2_X1 U18265 ( .A1(n16532), .A2(n16516), .ZN(n16470) );
  AOI22_X1 U18266 ( .A1(n18555), .A2(n16471), .B1(n18614), .B2(n16470), .ZN(
        n16472) );
  NAND2_X1 U18267 ( .A1(n16519), .A2(n16472), .ZN(n16507) );
  NOR2_X1 U18268 ( .A1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n16473), .ZN(
        n16506) );
  NOR2_X1 U18269 ( .A1(n16507), .A2(n16506), .ZN(n16493) );
  NAND2_X1 U18270 ( .A1(n16474), .A2(n16492), .ZN(n16494) );
  AOI21_X1 U18271 ( .B1(n16493), .B2(n16494), .A(n16475), .ZN(n16486) );
  INV_X1 U18272 ( .A(n16476), .ZN(n16480) );
  INV_X1 U18273 ( .A(n16477), .ZN(n16479) );
  AOI21_X1 U18274 ( .B1(n16480), .B2(n16479), .A(n16478), .ZN(n19455) );
  NAND2_X1 U18275 ( .A1(n18622), .A2(n19455), .ZN(n16483) );
  INV_X1 U18276 ( .A(n16481), .ZN(n16482) );
  OAI211_X1 U18277 ( .C1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .C2(n16484), .A(
        n16483), .B(n16482), .ZN(n16485) );
  AOI211_X1 U18278 ( .C1(n18353), .C2(n18591), .A(n16486), .B(n16485), .ZN(
        n16487) );
  OAI211_X1 U18279 ( .C1(n16489), .C2(n18617), .A(n16488), .B(n16487), .ZN(
        P2_U3026) );
  NAND2_X1 U18280 ( .A1(n16490), .A2(n18598), .ZN(n16500) );
  INV_X1 U18281 ( .A(n16491), .ZN(n18337) );
  NOR2_X1 U18282 ( .A1(n16493), .A2(n16492), .ZN(n16498) );
  OAI211_X1 U18283 ( .C1(n18594), .C2(n16496), .A(n16495), .B(n16494), .ZN(
        n16497) );
  AOI211_X1 U18284 ( .C1(n18337), .C2(n18591), .A(n16498), .B(n16497), .ZN(
        n16499) );
  OAI211_X1 U18285 ( .C1(n16501), .C2(n18617), .A(n16500), .B(n16499), .ZN(
        P2_U3027) );
  NAND2_X1 U18286 ( .A1(n16503), .A2(n16502), .ZN(n16504) );
  AND2_X1 U18287 ( .A1(n11008), .A2(n16504), .ZN(n19547) );
  AOI211_X1 U18288 ( .C1(n18622), .C2(n19547), .A(n16506), .B(n16505), .ZN(
        n16509) );
  NAND2_X1 U18289 ( .A1(n16507), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n16508) );
  OAI211_X1 U18290 ( .C1(n18321), .C2(n18605), .A(n16509), .B(n16508), .ZN(
        n16510) );
  AOI21_X1 U18291 ( .B1(n16511), .B2(n18598), .A(n16510), .ZN(n16512) );
  OAI21_X1 U18292 ( .B1(n18617), .B2(n16513), .A(n16512), .ZN(P2_U3028) );
  AOI21_X1 U18293 ( .B1(n11013), .B2(n18568), .A(n16514), .ZN(n18561) );
  NAND3_X1 U18294 ( .A1(n18617), .A2(n18608), .A3(
        P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n16515) );
  NAND2_X1 U18295 ( .A1(n17048), .A2(n16515), .ZN(n18558) );
  NAND3_X1 U18296 ( .A1(n16532), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A3(
        n16516), .ZN(n16517) );
  NAND2_X1 U18297 ( .A1(n18614), .A2(n16517), .ZN(n16518) );
  NAND2_X1 U18298 ( .A1(n16519), .A2(n16518), .ZN(n16540) );
  INV_X1 U18299 ( .A(n16540), .ZN(n18556) );
  AOI22_X1 U18300 ( .A1(n15174), .A2(n18561), .B1(n18558), .B2(n18556), .ZN(
        n16529) );
  OAI21_X1 U18301 ( .B1(n16522), .B2(n16521), .A(n16520), .ZN(n17059) );
  NOR2_X1 U18302 ( .A1(n17059), .A2(n18606), .ZN(n16528) );
  AOI21_X1 U18303 ( .B1(n16525), .B2(n16524), .A(n16523), .ZN(n19656) );
  AOI22_X1 U18304 ( .A1(n18622), .A2(n19656), .B1(P2_REIP_REG_16__SCAN_IN), 
        .B2(n18572), .ZN(n16526) );
  OAI21_X1 U18305 ( .B1(n18301), .B2(n18605), .A(n16526), .ZN(n16527) );
  OR3_X1 U18306 ( .A1(n16529), .A2(n16528), .A3(n16527), .ZN(P2_U3030) );
  INV_X1 U18307 ( .A(n16530), .ZN(n16542) );
  NAND2_X1 U18308 ( .A1(n18286), .A2(n18591), .ZN(n16536) );
  NAND3_X1 U18309 ( .A1(n18547), .A2(n16532), .A3(n16531), .ZN(n16534) );
  NAND2_X1 U18310 ( .A1(n18622), .A2(n18285), .ZN(n16533) );
  NAND4_X1 U18311 ( .A1(n16536), .A2(n16535), .A3(n16534), .A4(n16533), .ZN(
        n16539) );
  NOR2_X1 U18312 ( .A1(n16537), .A2(n18606), .ZN(n16538) );
  AOI211_X1 U18313 ( .C1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n16540), .A(
        n16539), .B(n16538), .ZN(n16541) );
  OAI21_X1 U18314 ( .B1(n18617), .B2(n16542), .A(n16541), .ZN(P2_U3031) );
  INV_X1 U18315 ( .A(n16547), .ZN(n16544) );
  NOR2_X1 U18316 ( .A1(n18516), .A2(n18555), .ZN(n16571) );
  INV_X1 U18317 ( .A(n16571), .ZN(n16543) );
  OAI21_X1 U18318 ( .B1(n16601), .B2(n16544), .A(n16543), .ZN(n16546) );
  NAND2_X1 U18319 ( .A1(n18547), .A2(n16563), .ZN(n16545) );
  NAND2_X1 U18320 ( .A1(n16546), .A2(n16545), .ZN(n18545) );
  INV_X1 U18321 ( .A(n18545), .ZN(n16561) );
  NAND2_X1 U18322 ( .A1(n16547), .A2(n18547), .ZN(n16562) );
  NOR2_X1 U18323 ( .A1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n16562), .ZN(
        n18546) );
  NAND2_X1 U18324 ( .A1(n18546), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n16552) );
  NOR2_X1 U18325 ( .A1(n16391), .A2(n18589), .ZN(n16549) );
  NOR2_X1 U18326 ( .A1(n18594), .A2(n18258), .ZN(n16548) );
  AOI211_X1 U18327 ( .C1(n16550), .C2(n18591), .A(n16549), .B(n16548), .ZN(
        n16551) );
  OAI211_X1 U18328 ( .C1(n15184), .C2(n16561), .A(n16552), .B(n16551), .ZN(
        n16553) );
  AOI21_X1 U18329 ( .B1(n16554), .B2(n18598), .A(n16553), .ZN(n16555) );
  OAI21_X1 U18330 ( .B1(n16556), .B2(n18617), .A(n16555), .ZN(P2_U3033) );
  NAND2_X1 U18331 ( .A1(n16558), .A2(n16557), .ZN(n16559) );
  AOI21_X1 U18332 ( .B1(n16563), .B2(n16568), .A(n16560), .ZN(n17028) );
  NAND2_X1 U18333 ( .A1(n17028), .A2(n18568), .ZN(n16567) );
  AOI21_X1 U18334 ( .B1(n16563), .B2(n16562), .A(n16561), .ZN(n16565) );
  OAI22_X1 U18335 ( .A1(n18249), .A2(n18605), .B1(n14217), .B2(n18589), .ZN(
        n16564) );
  AOI211_X1 U18336 ( .C1(n18246), .C2(n18622), .A(n16565), .B(n16564), .ZN(
        n16566) );
  OAI211_X1 U18337 ( .C1(n17026), .C2(n18606), .A(n16567), .B(n16566), .ZN(
        P2_U3034) );
  OAI21_X1 U18338 ( .B1(n16582), .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n16568), .ZN(n17016) );
  XNOR2_X1 U18339 ( .A(n16569), .B(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n16570) );
  INV_X1 U18340 ( .A(n17015), .ZN(n16580) );
  INV_X1 U18341 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n16574) );
  INV_X1 U18342 ( .A(n16601), .ZN(n16572) );
  AOI21_X1 U18343 ( .B1(n16572), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n16571), .ZN(n16593) );
  AND3_X1 U18344 ( .A1(n16583), .A2(n18547), .A3(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n16592) );
  OAI21_X1 U18345 ( .B1(n16593), .B2(n16592), .A(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16573) );
  OAI21_X1 U18346 ( .B1(n18589), .B2(n16574), .A(n16573), .ZN(n16577) );
  INV_X1 U18347 ( .A(n18547), .ZN(n16575) );
  NOR4_X1 U18348 ( .A1(n16575), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A3(
        n16583), .A4(n16603), .ZN(n16576) );
  AOI211_X1 U18349 ( .C1(n18591), .C2(n17018), .A(n16577), .B(n16576), .ZN(
        n16578) );
  OAI21_X1 U18350 ( .B1(n18229), .B2(n18594), .A(n16578), .ZN(n16579) );
  AOI21_X1 U18351 ( .B1(n16580), .B2(n18598), .A(n16579), .ZN(n16581) );
  OAI21_X1 U18352 ( .B1(n17016), .B2(n18617), .A(n16581), .ZN(P2_U3035) );
  AOI21_X1 U18353 ( .B1(n16583), .B2(n16599), .A(n16582), .ZN(n17009) );
  INV_X1 U18354 ( .A(n17009), .ZN(n16598) );
  INV_X1 U18355 ( .A(n16584), .ZN(n16610) );
  OR2_X1 U18356 ( .A1(n16585), .A2(n16610), .ZN(n16589) );
  NAND2_X1 U18357 ( .A1(n16587), .A2(n16586), .ZN(n16588) );
  XNOR2_X1 U18358 ( .A(n16589), .B(n16588), .ZN(n17011) );
  XNOR2_X1 U18359 ( .A(n13721), .B(n16590), .ZN(n19132) );
  NOR2_X1 U18360 ( .A1(n13922), .A2(n18589), .ZN(n16591) );
  AOI211_X1 U18361 ( .C1(n16593), .C2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n16592), .B(n16591), .ZN(n16595) );
  INV_X1 U18362 ( .A(n18215), .ZN(n17010) );
  NAND2_X1 U18363 ( .A1(n18591), .A2(n17010), .ZN(n16594) );
  OAI211_X1 U18364 ( .C1(n19132), .C2(n18594), .A(n16595), .B(n16594), .ZN(
        n16596) );
  AOI21_X1 U18365 ( .B1(n17011), .B2(n18598), .A(n16596), .ZN(n16597) );
  OAI21_X1 U18366 ( .B1(n16598), .B2(n18617), .A(n16597), .ZN(P2_U3036) );
  OAI21_X1 U18367 ( .B1(n16600), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n16599), .ZN(n17002) );
  INV_X1 U18368 ( .A(n18201), .ZN(n16608) );
  NAND2_X1 U18369 ( .A1(n16601), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n16606) );
  NOR2_X1 U18370 ( .A1(n13853), .A2(n18589), .ZN(n16602) );
  AOI21_X1 U18371 ( .B1(n18591), .B2(n17004), .A(n16602), .ZN(n16605) );
  NAND2_X1 U18372 ( .A1(n18547), .A2(n16603), .ZN(n16604) );
  NAND3_X1 U18373 ( .A1(n16606), .A2(n16605), .A3(n16604), .ZN(n16607) );
  AOI21_X1 U18374 ( .B1(n16608), .B2(n18622), .A(n16607), .ZN(n16614) );
  OR2_X1 U18375 ( .A1(n16610), .A2(n16609), .ZN(n16611) );
  XNOR2_X1 U18376 ( .A(n16612), .B(n16611), .ZN(n17001) );
  OR2_X1 U18377 ( .A1(n17001), .A2(n18606), .ZN(n16613) );
  OAI211_X1 U18378 ( .C1(n17002), .C2(n18617), .A(n16614), .B(n16613), .ZN(
        P2_U3037) );
  INV_X1 U18379 ( .A(n16630), .ZN(n16615) );
  OAI22_X1 U18380 ( .A1(n16617), .A2(n16616), .B1(n18608), .B2(n16615), .ZN(
        n16619) );
  OR2_X1 U18381 ( .A1(n16619), .A2(n16618), .ZN(n16633) );
  INV_X1 U18382 ( .A(n16633), .ZN(n16620) );
  OAI21_X1 U18383 ( .B1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n18608), .A(
        n16620), .ZN(n18567) );
  OAI22_X1 U18384 ( .A1(n18605), .A2(n18175), .B1(n17133), .B2(n18589), .ZN(
        n16621) );
  AOI21_X1 U18385 ( .B1(n18567), .B2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n16621), .ZN(n16625) );
  NOR2_X1 U18386 ( .A1(n16622), .A2(n18603), .ZN(n18574) );
  NAND2_X1 U18387 ( .A1(n18574), .A2(n16623), .ZN(n16624) );
  OAI211_X1 U18388 ( .C1(n18176), .C2(n18594), .A(n16625), .B(n16624), .ZN(
        n16626) );
  AOI21_X1 U18389 ( .B1(n16627), .B2(n18598), .A(n16626), .ZN(n16628) );
  OAI21_X1 U18390 ( .B1(n16629), .B2(n18617), .A(n16628), .ZN(P2_U3039) );
  NOR2_X1 U18391 ( .A1(n18162), .A2(n18594), .ZN(n16636) );
  NOR2_X1 U18392 ( .A1(n13834), .A2(n18589), .ZN(n16632) );
  NOR3_X1 U18393 ( .A1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n16630), .A3(
        n18603), .ZN(n16631) );
  AOI211_X1 U18394 ( .C1(n16633), .C2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n16632), .B(n16631), .ZN(n16634) );
  OAI21_X1 U18395 ( .B1(n18161), .B2(n18605), .A(n16634), .ZN(n16635) );
  AOI211_X1 U18396 ( .C1(n16637), .C2(n18598), .A(n16636), .B(n16635), .ZN(
        n16638) );
  OAI21_X1 U18397 ( .B1(n16639), .B2(n18617), .A(n16638), .ZN(P2_U3040) );
  INV_X1 U18398 ( .A(n18112), .ZN(n16642) );
  OAI22_X1 U18399 ( .A1(n10964), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        n16642), .B2(n16641), .ZN(n16649) );
  INV_X1 U18400 ( .A(n16649), .ZN(n16643) );
  OAI222_X1 U18401 ( .A1(n16669), .A2(n16645), .B1(n18628), .B2(n16644), .C1(
        n16719), .C2(n16643), .ZN(n16646) );
  MUX2_X1 U18402 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B(n16646), .S(
        n16652), .Z(P2_U3601) );
  INV_X1 U18403 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18537) );
  OAI211_X1 U18404 ( .C1(n18112), .C2(n16648), .A(n10964), .B(n16647), .ZN(
        n18123) );
  OAI21_X1 U18405 ( .B1(n10964), .B2(n18537), .A(n18123), .ZN(n16655) );
  NOR2_X1 U18406 ( .A1(n16719), .A2(n16649), .ZN(n16654) );
  INV_X1 U18407 ( .A(n16654), .ZN(n16651) );
  OAI222_X1 U18408 ( .A1(n19152), .A2(n16669), .B1(n16655), .B2(n16651), .C1(
        n16650), .C2(n18628), .ZN(n16653) );
  INV_X1 U18409 ( .A(n16652), .ZN(n16661) );
  MUX2_X1 U18410 ( .A(n16653), .B(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .S(
        n16661), .Z(P2_U3600) );
  INV_X1 U18411 ( .A(n16669), .ZN(n18642) );
  AOI222_X1 U18412 ( .A1(n16657), .A2(n16656), .B1(n16655), .B2(n16654), .C1(
        n18642), .C2(n17077), .ZN(n16659) );
  NAND2_X1 U18413 ( .A1(n16661), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n16658) );
  OAI21_X1 U18414 ( .B1(n16659), .B2(n16661), .A(n16658), .ZN(P2_U3599) );
  OAI22_X1 U18415 ( .A1(n19328), .A2(n16669), .B1(n16660), .B2(n18628), .ZN(
        n16662) );
  MUX2_X1 U18416 ( .A(n16662), .B(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n16661), .Z(P2_U3596) );
  INV_X1 U18417 ( .A(n19169), .ZN(n16664) );
  INV_X1 U18418 ( .A(n19278), .ZN(n16663) );
  NOR2_X1 U18419 ( .A1(n19784), .A2(n19779), .ZN(n16665) );
  OAI21_X1 U18420 ( .B1(n16665), .B2(n21695), .A(n19332), .ZN(n16676) );
  INV_X1 U18421 ( .A(n16666), .ZN(n19677) );
  AOI21_X1 U18422 ( .B1(n16719), .B2(n19264), .A(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n18644) );
  NAND2_X1 U18423 ( .A1(n16667), .A2(n19203), .ZN(n19334) );
  OAI21_X1 U18424 ( .B1(n15117), .B2(n19334), .A(n19252), .ZN(n16670) );
  OAI21_X1 U18425 ( .B1(n16676), .B2(n19677), .A(n16670), .ZN(n16672) );
  NAND2_X1 U18426 ( .A1(n19231), .A2(n19200), .ZN(n19322) );
  NOR2_X1 U18427 ( .A1(n19280), .A2(n19322), .ZN(n19778) );
  INV_X1 U18428 ( .A(n19778), .ZN(n16671) );
  NOR2_X1 U18429 ( .A1(n19677), .A2(n19778), .ZN(n16675) );
  OAI21_X1 U18430 ( .B1(n16673), .B2(n19778), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n16674) );
  INV_X1 U18431 ( .A(BUF2_REG_27__SCAN_IN), .ZN(n18660) );
  INV_X1 U18432 ( .A(n19537), .ZN(n19545) );
  AOI22_X1 U18433 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n19672), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n19671), .ZN(n19540) );
  NOR2_X2 U18434 ( .A1(n12702), .A2(n19675), .ZN(n19541) );
  AOI22_X1 U18435 ( .A1(n19542), .A2(n19779), .B1(n19778), .B2(n19541), .ZN(
        n16680) );
  OAI21_X1 U18436 ( .B1(n19545), .B2(n19562), .A(n16680), .ZN(n16681) );
  AOI21_X1 U18437 ( .B1(n19781), .B2(n16677), .A(n16681), .ZN(n16682) );
  OAI21_X1 U18438 ( .B1(n19788), .B2(n16683), .A(n16682), .ZN(P2_U3051) );
  NOR2_X2 U18439 ( .A1(n19413), .A2(n19673), .ZN(n19448) );
  INV_X1 U18440 ( .A(BUF2_REG_29__SCAN_IN), .ZN(n18657) );
  AOI22_X1 U18441 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n19672), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n19671), .ZN(n19431) );
  NOR2_X2 U18442 ( .A1(n16684), .A2(n19675), .ZN(n19447) );
  AOI22_X1 U18443 ( .A1(n19449), .A2(n19779), .B1(n19778), .B2(n19447), .ZN(
        n16685) );
  OAI21_X1 U18444 ( .B1(n19452), .B2(n19562), .A(n16685), .ZN(n16686) );
  AOI21_X1 U18445 ( .B1(n19781), .B2(n19448), .A(n16686), .ZN(n16687) );
  OAI21_X1 U18446 ( .B1(n19788), .B2(n16688), .A(n16687), .ZN(P2_U3053) );
  NAND2_X1 U18447 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18707) );
  NAND2_X1 U18448 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n17879) );
  INV_X1 U18449 ( .A(n17879), .ZN(n17924) );
  INV_X1 U18450 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n21288) );
  NOR2_X1 U18451 ( .A1(n20798), .A2(n21288), .ZN(n17531) );
  NOR2_X1 U18452 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n17531), .ZN(n17533) );
  INV_X1 U18453 ( .A(n17533), .ZN(n20108) );
  NOR2_X1 U18454 ( .A1(n17924), .A2(n20108), .ZN(n16691) );
  NAND2_X1 U18455 ( .A1(n21262), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n18704) );
  NAND2_X1 U18456 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n17531), .ZN(n21295) );
  INV_X1 U18457 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n16701) );
  OAI21_X1 U18458 ( .B1(n16689), .B2(n20825), .A(n16701), .ZN(n16699) );
  NOR2_X1 U18459 ( .A1(n17205), .A2(n16699), .ZN(n17532) );
  INV_X1 U18460 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n21316) );
  INV_X1 U18461 ( .A(n21300), .ZN(n16690) );
  OAI221_X1 U18462 ( .B1(n21295), .B2(n17532), .C1(n21295), .C2(n21316), .A(
        n19010), .ZN(n17976) );
  NAND2_X1 U18463 ( .A1(n18704), .A2(n17976), .ZN(n17977) );
  AOI221_X1 U18464 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n18707), .C1(n16691), 
        .C2(n18707), .A(n17977), .ZN(n17974) );
  AOI21_X1 U18465 ( .B1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(
        P3_STATE2_REG_3__SCAN_IN), .A(n16691), .ZN(n16692) );
  INV_X1 U18466 ( .A(n16692), .ZN(n17975) );
  OAI221_X1 U18467 ( .B1(n18703), .B2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .C1(n18703), .C2(n17975), .A(n17976), .ZN(n17972) );
  AOI22_X1 U18468 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n17974), .B1(
        n17972), .B2(n18692), .ZN(P3_U2865) );
  NOR2_X1 U18469 ( .A1(n21255), .A2(n17148), .ZN(n16696) );
  OR2_X2 U18470 ( .A1(n16698), .A2(n20111), .ZN(n20613) );
  INV_X1 U18471 ( .A(n20613), .ZN(n16693) );
  NAND2_X1 U18472 ( .A1(n20164), .A2(n16713), .ZN(n16712) );
  AOI211_X1 U18473 ( .C1(n16693), .C2(n16712), .A(n21707), .B(n21280), .ZN(
        n16695) );
  NOR2_X1 U18474 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n21296), .ZN(n18685) );
  NOR2_X1 U18475 ( .A1(n21316), .A2(n21295), .ZN(n16697) );
  AND2_X1 U18476 ( .A1(n16699), .A2(n16698), .ZN(n21258) );
  NAND2_X1 U18477 ( .A1(n20798), .A2(n21296), .ZN(n20802) );
  INV_X1 U18478 ( .A(n20802), .ZN(n20839) );
  NAND3_X1 U18479 ( .A1(n20841), .A2(n21258), .A3(n20839), .ZN(n16700) );
  OAI21_X1 U18480 ( .B1(n20841), .B2(n16701), .A(n16700), .ZN(P3_U3284) );
  INV_X1 U18481 ( .A(n21432), .ZN(n16704) );
  NAND4_X1 U18482 ( .A1(n16704), .A2(n16703), .A3(n16702), .A4(n21661), .ZN(
        n16705) );
  OAI21_X1 U18483 ( .B1(n21661), .B2(n11775), .A(n16705), .ZN(P1_U3468) );
  INV_X1 U18484 ( .A(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(n16706) );
  INV_X1 U18485 ( .A(P3_STATE_REG_1__SCAN_IN), .ZN(n21747) );
  OAI21_X1 U18486 ( .B1(P3_STATE_REG_2__SCAN_IN), .B2(n21747), .A(
        P3_STATE_REG_0__SCAN_IN), .ZN(n18041) );
  NAND2_X1 U18487 ( .A1(n21756), .A2(n18041), .ZN(n16708) );
  INV_X1 U18488 ( .A(n16708), .ZN(n21703) );
  INV_X1 U18489 ( .A(BS16), .ZN(n16734) );
  NAND2_X1 U18490 ( .A1(n21758), .A2(n21747), .ZN(n21705) );
  AOI21_X1 U18491 ( .B1(n16734), .B2(n21705), .A(n16707), .ZN(n21699) );
  AOI21_X1 U18492 ( .B1(n16706), .B2(n16707), .A(n21699), .ZN(P3_U3280) );
  AND2_X1 U18493 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n16707), .ZN(P3_U3028) );
  AND2_X1 U18494 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n16707), .ZN(P3_U3027) );
  AND2_X1 U18495 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n16707), .ZN(P3_U3026) );
  AND2_X1 U18496 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n16707), .ZN(P3_U3025) );
  AND2_X1 U18497 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n16707), .ZN(P3_U3024) );
  AND2_X1 U18498 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n16707), .ZN(P3_U3023) );
  AND2_X1 U18499 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n16707), .ZN(P3_U3022) );
  AND2_X1 U18500 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n16707), .ZN(P3_U3021) );
  AND2_X1 U18501 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n16707), .ZN(
        P3_U3020) );
  AND2_X1 U18502 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n16707), .ZN(
        P3_U3019) );
  AND2_X1 U18503 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n16707), .ZN(
        P3_U3018) );
  AND2_X1 U18504 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n16707), .ZN(
        P3_U3017) );
  AND2_X1 U18505 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n16707), .ZN(
        P3_U3016) );
  AND2_X1 U18506 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n16708), .ZN(
        P3_U3015) );
  AND2_X1 U18507 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n16708), .ZN(
        P3_U3014) );
  AND2_X1 U18508 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n16708), .ZN(
        P3_U3013) );
  AND2_X1 U18509 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n16708), .ZN(
        P3_U3012) );
  AND2_X1 U18510 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n16708), .ZN(
        P3_U3011) );
  AND2_X1 U18511 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n16708), .ZN(
        P3_U3010) );
  AND2_X1 U18512 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n16708), .ZN(
        P3_U3009) );
  AND2_X1 U18513 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n16708), .ZN(
        P3_U3008) );
  AND2_X1 U18514 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n16708), .ZN(
        P3_U3007) );
  AND2_X1 U18515 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n16708), .ZN(
        P3_U3006) );
  AND2_X1 U18516 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n16708), .ZN(
        P3_U3005) );
  AND2_X1 U18517 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n16708), .ZN(
        P3_U3004) );
  AND2_X1 U18518 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n16707), .ZN(
        P3_U3003) );
  AND2_X1 U18519 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n16707), .ZN(
        P3_U3002) );
  AND2_X1 U18520 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n16707), .ZN(
        P3_U3001) );
  AND2_X1 U18521 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n16707), .ZN(
        P3_U3000) );
  AND2_X1 U18522 ( .A1(P3_DATAWIDTH_REG_31__SCAN_IN), .A2(n16708), .ZN(
        P3_U2999) );
  OAI21_X1 U18523 ( .B1(n21309), .B2(n20798), .A(n21288), .ZN(n16709) );
  NAND4_X1 U18524 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_0__SCAN_IN), .A3(n21707), .A4(n21288), .ZN(n21292) );
  OAI211_X1 U18525 ( .C1(n17924), .C2(n16709), .A(n21295), .B(n21292), .ZN(
        n16710) );
  INV_X1 U18526 ( .A(n16710), .ZN(P3_U2998) );
  NOR2_X1 U18527 ( .A1(n16711), .A2(n17976), .ZN(P3_U2867) );
  NAND2_X1 U18528 ( .A1(n21309), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n17967) );
  NOR2_X4 U18529 ( .A1(n21248), .A2(n18019), .ZN(n18032) );
  AND2_X1 U18530 ( .A1(n18032), .A2(P3_DATAO_REG_31__SCAN_IN), .ZN(P3_U2736)
         );
  INV_X1 U18531 ( .A(n20165), .ZN(n16715) );
  AND2_X1 U18532 ( .A1(n17530), .A2(n16715), .ZN(n16716) );
  INV_X1 U18533 ( .A(P3_READREQUEST_REG_SCAN_IN), .ZN(n16714) );
  AOI22_X1 U18534 ( .A1(n20104), .A2(n20165), .B1(n16716), .B2(n16714), .ZN(
        P3_U3298) );
  INV_X1 U18535 ( .A(P3_MEMORYFETCH_REG_SCAN_IN), .ZN(n17998) );
  NOR2_X1 U18536 ( .A1(n20166), .A2(n16715), .ZN(n20601) );
  AOI21_X1 U18537 ( .B1(n16716), .B2(n17998), .A(n20601), .ZN(P3_U3299) );
  NOR2_X1 U18538 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(n21728), .ZN(n21736) );
  AOI21_X1 U18539 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(n21736), .A(n21731), 
        .ZN(n16717) );
  INV_X1 U18540 ( .A(n16717), .ZN(n21698) );
  INV_X1 U18541 ( .A(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n16733) );
  NAND2_X1 U18542 ( .A1(n21745), .A2(n21728), .ZN(n21727) );
  AOI21_X1 U18543 ( .B1(n16734), .B2(n21727), .A(n17093), .ZN(n21694) );
  AOI21_X1 U18544 ( .B1(n17093), .B2(n16733), .A(n21694), .ZN(P2_U3591) );
  AND2_X1 U18545 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n17093), .ZN(P2_U3208) );
  AND2_X1 U18546 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n16717), .ZN(P2_U3207) );
  AND2_X1 U18547 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n17093), .ZN(P2_U3206) );
  AND2_X1 U18548 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n17093), .ZN(P2_U3205) );
  AND2_X1 U18549 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n17093), .ZN(P2_U3204) );
  AND2_X1 U18550 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n17093), .ZN(P2_U3203) );
  AND2_X1 U18551 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n16717), .ZN(P2_U3202) );
  AND2_X1 U18552 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n16717), .ZN(P2_U3201) );
  AND2_X1 U18553 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n16717), .ZN(
        P2_U3200) );
  AND2_X1 U18554 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n16717), .ZN(
        P2_U3199) );
  AND2_X1 U18555 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n16717), .ZN(
        P2_U3198) );
  AND2_X1 U18556 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n16717), .ZN(
        P2_U3197) );
  AND2_X1 U18557 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n16717), .ZN(
        P2_U3196) );
  AND2_X1 U18558 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n16717), .ZN(
        P2_U3195) );
  AND2_X1 U18559 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n16717), .ZN(
        P2_U3194) );
  AND2_X1 U18560 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n16717), .ZN(
        P2_U3193) );
  AND2_X1 U18561 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n16717), .ZN(
        P2_U3192) );
  AND2_X1 U18562 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n16717), .ZN(
        P2_U3191) );
  AND2_X1 U18563 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n17093), .ZN(
        P2_U3190) );
  AND2_X1 U18564 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n17093), .ZN(
        P2_U3189) );
  AND2_X1 U18565 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n17093), .ZN(
        P2_U3188) );
  AND2_X1 U18566 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n17093), .ZN(
        P2_U3187) );
  AND2_X1 U18567 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n16717), .ZN(
        P2_U3186) );
  AND2_X1 U18568 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n17093), .ZN(
        P2_U3185) );
  AND2_X1 U18569 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n17093), .ZN(
        P2_U3184) );
  AND2_X1 U18570 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n17093), .ZN(
        P2_U3183) );
  AND2_X1 U18571 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n17093), .ZN(
        P2_U3182) );
  AND2_X1 U18572 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n17093), .ZN(
        P2_U3181) );
  AND2_X1 U18573 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n17093), .ZN(
        P2_U3180) );
  AND2_X1 U18574 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n17093), .ZN(
        P2_U3179) );
  NAND2_X1 U18575 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n21729), .ZN(n18629) );
  AOI21_X1 U18576 ( .B1(n16718), .B2(n13554), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n16720) );
  AOI221_X1 U18577 ( .B1(n18629), .B2(n16720), .C1(n16719), .C2(n16720), .A(
        n16721), .ZN(P2_U3178) );
  AOI221_X1 U18578 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(n16721), .C1(n18638), .C2(
        n16721), .A(n19331), .ZN(n17082) );
  INV_X1 U18579 ( .A(n17082), .ZN(n17080) );
  NOR2_X1 U18580 ( .A1(n16722), .A2(n17080), .ZN(P2_U3047) );
  AND2_X1 U18581 ( .A1(n17114), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(P2_U2920)
         );
  NOR4_X1 U18582 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_12__SCAN_IN), .A3(P2_DATAWIDTH_REG_11__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_10__SCAN_IN), .ZN(n16726) );
  NOR4_X1 U18583 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_16__SCAN_IN), .A3(P2_DATAWIDTH_REG_15__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_14__SCAN_IN), .ZN(n16725) );
  NOR4_X1 U18584 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_4__SCAN_IN), .A3(P2_DATAWIDTH_REG_3__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_2__SCAN_IN), .ZN(n16724) );
  NOR4_X1 U18585 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_8__SCAN_IN), .A3(P2_DATAWIDTH_REG_7__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_6__SCAN_IN), .ZN(n16723) );
  NAND4_X1 U18586 ( .A1(n16726), .A2(n16725), .A3(n16724), .A4(n16723), .ZN(
        n16732) );
  NOR4_X1 U18587 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_28__SCAN_IN), .A3(P2_DATAWIDTH_REG_27__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_26__SCAN_IN), .ZN(n16730) );
  AOI211_X1 U18588 ( .C1(P2_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_1__SCAN_IN), .A(P2_DATAWIDTH_REG_31__SCAN_IN), .B(
        P2_DATAWIDTH_REG_30__SCAN_IN), .ZN(n16729) );
  NOR4_X1 U18589 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_20__SCAN_IN), .A3(P2_DATAWIDTH_REG_19__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_18__SCAN_IN), .ZN(n16728) );
  NOR4_X1 U18590 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_24__SCAN_IN), .A3(P2_DATAWIDTH_REG_23__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_22__SCAN_IN), .ZN(n16727) );
  NAND4_X1 U18591 ( .A1(n16730), .A2(n16729), .A3(n16728), .A4(n16727), .ZN(
        n16731) );
  NOR2_X1 U18592 ( .A1(n16732), .A2(n16731), .ZN(n17089) );
  INV_X1 U18593 ( .A(n17089), .ZN(n17088) );
  NOR2_X1 U18594 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n17088), .ZN(n17083) );
  INV_X1 U18595 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n21697) );
  NAND3_X1 U18596 ( .A1(n18102), .A2(n21697), .A3(n16733), .ZN(n17087) );
  INV_X1 U18597 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n17142) );
  AOI22_X1 U18598 ( .A1(n17083), .A2(n17087), .B1(n17088), .B2(n17142), .ZN(
        P2_U2821) );
  INV_X1 U18599 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n17140) );
  AOI22_X1 U18600 ( .A1(n17083), .A2(n18102), .B1(n17088), .B2(n17140), .ZN(
        P2_U2820) );
  NAND2_X1 U18601 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(n20034), .ZN(n22219) );
  NAND2_X1 U18602 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n21711), .ZN(n16774) );
  INV_X1 U18603 ( .A(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(n16735) );
  AOI221_X1 U18604 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n16734), .C1(
        P1_STATE_REG_2__SCAN_IN), .C2(n16734), .A(n16736), .ZN(n21692) );
  AOI21_X1 U18605 ( .B1(n16736), .B2(n16735), .A(n21692), .ZN(P1_U3464) );
  AND2_X1 U18606 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n16736), .ZN(P1_U3193) );
  AND2_X1 U18607 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n16736), .ZN(P1_U3192) );
  AND2_X1 U18608 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n16736), .ZN(P1_U3191) );
  AND2_X1 U18609 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n16736), .ZN(P1_U3190) );
  AND2_X1 U18610 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n16736), .ZN(P1_U3189) );
  AND2_X1 U18611 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n16736), .ZN(P1_U3188) );
  AND2_X1 U18612 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n16736), .ZN(P1_U3187) );
  AND2_X1 U18613 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n16736), .ZN(P1_U3186) );
  AND2_X1 U18614 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n16736), .ZN(
        P1_U3185) );
  AND2_X1 U18615 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(n16736), .ZN(
        P1_U3184) );
  AND2_X1 U18616 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n16736), .ZN(
        P1_U3183) );
  AND2_X1 U18617 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(n16736), .ZN(
        P1_U3182) );
  AND2_X1 U18618 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n16736), .ZN(
        P1_U3181) );
  AND2_X1 U18619 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n16736), .ZN(
        P1_U3179) );
  AND2_X1 U18620 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n16736), .ZN(
        P1_U3178) );
  AND2_X1 U18621 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n16736), .ZN(
        P1_U3177) );
  AND2_X1 U18622 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n16736), .ZN(
        P1_U3176) );
  AND2_X1 U18623 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n16736), .ZN(
        P1_U3175) );
  AND2_X1 U18624 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n16736), .ZN(
        P1_U3174) );
  AND2_X1 U18625 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n16736), .ZN(
        P1_U3173) );
  AND2_X1 U18626 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n16736), .ZN(
        P1_U3172) );
  AND2_X1 U18627 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n16736), .ZN(
        P1_U3171) );
  AND2_X1 U18628 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n16736), .ZN(
        P1_U3170) );
  AND2_X1 U18629 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n16736), .ZN(
        P1_U3169) );
  AND2_X1 U18630 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n16736), .ZN(
        P1_U3168) );
  AND2_X1 U18631 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n16736), .ZN(
        P1_U3167) );
  AND2_X1 U18632 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n16736), .ZN(
        P1_U3166) );
  AND2_X1 U18633 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n16736), .ZN(
        P1_U3165) );
  AND2_X1 U18634 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n16736), .ZN(
        P1_U3164) );
  INV_X1 U18635 ( .A(n16737), .ZN(n16768) );
  INV_X1 U18636 ( .A(n16738), .ZN(n16754) );
  INV_X1 U18637 ( .A(n16739), .ZN(n16742) );
  NOR2_X1 U18638 ( .A1(n16740), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n16741) );
  AOI21_X1 U18639 ( .B1(n16743), .B2(n16742), .A(n16741), .ZN(n21660) );
  NAND2_X1 U18640 ( .A1(n16744), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n21665) );
  AND2_X1 U18641 ( .A1(n21665), .A2(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n16745) );
  AND2_X1 U18642 ( .A1(n21660), .A2(n16745), .ZN(n16746) );
  INV_X1 U18643 ( .A(n16746), .ZN(n16750) );
  OAI22_X1 U18644 ( .A1(n16748), .A2(n16747), .B1(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n16746), .ZN(n16749) );
  OAI21_X1 U18645 ( .B1(n16750), .B2(n21864), .A(n16749), .ZN(n16751) );
  AOI222_X1 U18646 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n16752), 
        .B1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n16751), .C1(n16752), 
        .C2(n16751), .ZN(n16753) );
  AOI222_X1 U18647 ( .A1(n16754), .A2(n16753), .B1(n16754), .B2(n12300), .C1(
        n16753), .C2(n12300), .ZN(n16761) );
  AOI21_X1 U18648 ( .B1(n16948), .B2(n21656), .A(n16755), .ZN(n16757) );
  NOR4_X1 U18649 ( .A1(n16759), .A2(n16758), .A3(n16757), .A4(n16756), .ZN(
        n16760) );
  OAI21_X1 U18650 ( .B1(n16761), .B2(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A(
        n16760), .ZN(n16762) );
  INV_X1 U18651 ( .A(n16762), .ZN(n21690) );
  NOR4_X1 U18652 ( .A1(n16764), .A2(n21712), .A3(P1_STATEBS16_REG_SCAN_IN), 
        .A4(n16763), .ZN(n16767) );
  NOR2_X1 U18653 ( .A1(n16766), .A2(n16765), .ZN(n21677) );
  AOI211_X1 U18654 ( .C1(P1_STATE2_REG_1__SCAN_IN), .C2(n21675), .A(n16767), 
        .B(n21677), .ZN(n16769) );
  OAI221_X1 U18655 ( .B1(P1_STATE2_REG_1__SCAN_IN), .B2(
        P1_STATE2_REG_0__SCAN_IN), .C1(P1_STATE2_REG_1__SCAN_IN), .C2(n21690), 
        .A(n16769), .ZN(n21681) );
  OAI211_X1 U18656 ( .C1(P1_STATE2_REG_2__SCAN_IN), .C2(n21675), .A(n16768), 
        .B(n21681), .ZN(n21686) );
  OAI221_X1 U18657 ( .B1(P1_STATE2_REG_0__SCAN_IN), .B2(n14152), .C1(n21321), 
        .C2(n21712), .A(n21910), .ZN(n16771) );
  NOR2_X1 U18658 ( .A1(n16772), .A2(n16769), .ZN(n16770) );
  AOI22_X1 U18659 ( .A1(n21686), .A2(n16772), .B1(n16771), .B2(n16770), .ZN(
        P1_U3162) );
  NOR2_X1 U18660 ( .A1(n16773), .A2(n21674), .ZN(P1_U3032) );
  AND2_X1 U18661 ( .A1(n19866), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(P1_U2905)
         );
  OAI21_X1 U18662 ( .B1(n16774), .B2(P1_ADS_N_REG_SCAN_IN), .A(n22219), .ZN(
        n16775) );
  INV_X1 U18663 ( .A(n16775), .ZN(P1_U2802) );
  NAND2_X1 U18664 ( .A1(n16736), .A2(P1_DATAWIDTH_REG_15__SCAN_IN), .ZN(n16976) );
  OAI22_X1 U18665 ( .A1(P1_REIP_REG_20__SCAN_IN), .A2(keyinput_63), .B1(
        keyinput_61), .B2(P1_REIP_REG_22__SCAN_IN), .ZN(n16776) );
  AOI221_X1 U18666 ( .B1(P1_REIP_REG_20__SCAN_IN), .B2(keyinput_63), .C1(
        P1_REIP_REG_22__SCAN_IN), .C2(keyinput_61), .A(n16776), .ZN(n16866) );
  INV_X1 U18667 ( .A(keyinput_60), .ZN(n16864) );
  INV_X1 U18668 ( .A(keyinput_59), .ZN(n16862) );
  OAI22_X1 U18669 ( .A1(P1_REIP_REG_31__SCAN_IN), .A2(keyinput_52), .B1(
        keyinput_53), .B2(P1_REIP_REG_30__SCAN_IN), .ZN(n16777) );
  AOI221_X1 U18670 ( .B1(P1_REIP_REG_31__SCAN_IN), .B2(keyinput_52), .C1(
        P1_REIP_REG_30__SCAN_IN), .C2(keyinput_53), .A(n16777), .ZN(n16856) );
  INV_X1 U18671 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n19934) );
  INV_X1 U18672 ( .A(keyinput_51), .ZN(n16852) );
  INV_X1 U18673 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n19950) );
  INV_X1 U18674 ( .A(keyinput_50), .ZN(n16850) );
  INV_X1 U18675 ( .A(keyinput_49), .ZN(n16848) );
  INV_X1 U18676 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n19954) );
  AOI22_X1 U18677 ( .A1(P1_REQUESTPENDING_REG_SCAN_IN), .A2(keyinput_43), .B1(
        P1_STATEBS16_REG_SCAN_IN), .B2(keyinput_44), .ZN(n16778) );
  OAI221_X1 U18678 ( .B1(P1_REQUESTPENDING_REG_SCAN_IN), .B2(keyinput_43), 
        .C1(P1_STATEBS16_REG_SCAN_IN), .C2(keyinput_44), .A(n16778), .ZN(
        n16841) );
  XOR2_X1 U18679 ( .A(keyinput_29), .B(DATAI_3_), .Z(n16827) );
  INV_X1 U18680 ( .A(keyinput_28), .ZN(n16821) );
  AOI22_X1 U18681 ( .A1(n16780), .A2(keyinput_12), .B1(keyinput_13), .B2(
        n16889), .ZN(n16779) );
  OAI221_X1 U18682 ( .B1(n16780), .B2(keyinput_12), .C1(n16889), .C2(
        keyinput_13), .A(n16779), .ZN(n16800) );
  XNOR2_X1 U18683 ( .A(DATAI_26_), .B(keyinput_6), .ZN(n16791) );
  INV_X1 U18684 ( .A(keyinput_5), .ZN(n16789) );
  OAI22_X1 U18685 ( .A1(DATAI_31_), .A2(keyinput_1), .B1(keyinput_0), .B2(
        P1_MEMORYFETCH_REG_SCAN_IN), .ZN(n16781) );
  AOI221_X1 U18686 ( .B1(DATAI_31_), .B2(keyinput_1), .C1(
        P1_MEMORYFETCH_REG_SCAN_IN), .C2(keyinput_0), .A(n16781), .ZN(n16785)
         );
  AOI22_X1 U18687 ( .A1(DATAI_30_), .A2(keyinput_2), .B1(n16783), .B2(
        keyinput_4), .ZN(n16782) );
  OAI221_X1 U18688 ( .B1(DATAI_30_), .B2(keyinput_2), .C1(n16783), .C2(
        keyinput_4), .A(n16782), .ZN(n16784) );
  AOI211_X1 U18689 ( .C1(n16787), .C2(keyinput_3), .A(n16785), .B(n16784), 
        .ZN(n16786) );
  OAI21_X1 U18690 ( .B1(n16787), .B2(keyinput_3), .A(n16786), .ZN(n16788) );
  OAI221_X1 U18691 ( .B1(DATAI_27_), .B2(n16789), .C1(n16882), .C2(keyinput_5), 
        .A(n16788), .ZN(n16790) );
  AOI22_X1 U18692 ( .A1(n16791), .A2(n16790), .B1(keyinput_8), .B2(n16793), 
        .ZN(n16792) );
  OAI21_X1 U18693 ( .B1(keyinput_8), .B2(n16793), .A(n16792), .ZN(n16798) );
  AOI22_X1 U18694 ( .A1(DATAI_23_), .A2(keyinput_9), .B1(DATAI_25_), .B2(
        keyinput_7), .ZN(n16794) );
  OAI221_X1 U18695 ( .B1(DATAI_23_), .B2(keyinput_9), .C1(DATAI_25_), .C2(
        keyinput_7), .A(n16794), .ZN(n16797) );
  OAI22_X1 U18696 ( .A1(DATAI_22_), .A2(keyinput_10), .B1(DATAI_21_), .B2(
        keyinput_11), .ZN(n16795) );
  AOI221_X1 U18697 ( .B1(DATAI_22_), .B2(keyinput_10), .C1(keyinput_11), .C2(
        DATAI_21_), .A(n16795), .ZN(n16796) );
  OAI21_X1 U18698 ( .B1(n16798), .B2(n16797), .A(n16796), .ZN(n16799) );
  OAI22_X1 U18699 ( .A1(n16800), .A2(n16799), .B1(n16899), .B2(keyinput_14), 
        .ZN(n16801) );
  AOI21_X1 U18700 ( .B1(n16899), .B2(keyinput_14), .A(n16801), .ZN(n16809) );
  OAI22_X1 U18701 ( .A1(n16803), .A2(keyinput_15), .B1(DATAI_16_), .B2(
        keyinput_16), .ZN(n16802) );
  AOI221_X1 U18702 ( .B1(n16803), .B2(keyinput_15), .C1(keyinput_16), .C2(
        DATAI_16_), .A(n16802), .ZN(n16808) );
  INV_X1 U18703 ( .A(DATAI_14_), .ZN(n16905) );
  INV_X1 U18704 ( .A(DATAI_12_), .ZN(n16902) );
  AOI22_X1 U18705 ( .A1(n16905), .A2(keyinput_18), .B1(keyinput_20), .B2(
        n16902), .ZN(n16804) );
  OAI221_X1 U18706 ( .B1(n16905), .B2(keyinput_18), .C1(n16902), .C2(
        keyinput_20), .A(n16804), .ZN(n16807) );
  INV_X1 U18707 ( .A(DATAI_13_), .ZN(n16903) );
  AOI22_X1 U18708 ( .A1(DATAI_15_), .A2(keyinput_17), .B1(n16903), .B2(
        keyinput_19), .ZN(n16805) );
  OAI221_X1 U18709 ( .B1(DATAI_15_), .B2(keyinput_17), .C1(n16903), .C2(
        keyinput_19), .A(n16805), .ZN(n16806) );
  AOI211_X1 U18710 ( .C1(n16809), .C2(n16808), .A(n16807), .B(n16806), .ZN(
        n16817) );
  AOI22_X1 U18711 ( .A1(n16872), .A2(keyinput_22), .B1(n16811), .B2(
        keyinput_21), .ZN(n16810) );
  OAI221_X1 U18712 ( .B1(n16872), .B2(keyinput_22), .C1(n16811), .C2(
        keyinput_21), .A(n16810), .ZN(n16816) );
  OAI22_X1 U18713 ( .A1(n16914), .A2(keyinput_26), .B1(keyinput_23), .B2(
        DATAI_9_), .ZN(n16812) );
  AOI221_X1 U18714 ( .B1(n16914), .B2(keyinput_26), .C1(DATAI_9_), .C2(
        keyinput_23), .A(n16812), .ZN(n16815) );
  OAI22_X1 U18715 ( .A1(n16911), .A2(keyinput_24), .B1(DATAI_7_), .B2(
        keyinput_25), .ZN(n16813) );
  AOI221_X1 U18716 ( .B1(n16911), .B2(keyinput_24), .C1(keyinput_25), .C2(
        DATAI_7_), .A(n16813), .ZN(n16814) );
  OAI211_X1 U18717 ( .C1(n16817), .C2(n16816), .A(n16815), .B(n16814), .ZN(
        n16818) );
  AOI21_X1 U18718 ( .B1(DATAI_5_), .B2(keyinput_27), .A(n16818), .ZN(n16819)
         );
  OAI21_X1 U18719 ( .B1(DATAI_5_), .B2(keyinput_27), .A(n16819), .ZN(n16820)
         );
  OAI221_X1 U18720 ( .B1(DATAI_4_), .B2(n16821), .C1(n16923), .C2(keyinput_28), 
        .A(n16820), .ZN(n16826) );
  INV_X1 U18721 ( .A(HOLD), .ZN(n21757) );
  AOI22_X1 U18722 ( .A1(keyinput_30), .A2(DATAI_2_), .B1(n21757), .B2(
        keyinput_33), .ZN(n16822) );
  OAI221_X1 U18723 ( .B1(keyinput_30), .B2(DATAI_2_), .C1(n21757), .C2(
        keyinput_33), .A(n16822), .ZN(n16825) );
  AOI22_X1 U18724 ( .A1(DATAI_0_), .A2(keyinput_32), .B1(DATAI_1_), .B2(
        keyinput_31), .ZN(n16823) );
  OAI221_X1 U18725 ( .B1(DATAI_0_), .B2(keyinput_32), .C1(DATAI_1_), .C2(
        keyinput_31), .A(n16823), .ZN(n16824) );
  AOI211_X1 U18726 ( .C1(n16827), .C2(n16826), .A(n16825), .B(n16824), .ZN(
        n16835) );
  OAI22_X1 U18727 ( .A1(READY1), .A2(keyinput_36), .B1(READY2), .B2(
        keyinput_37), .ZN(n16828) );
  AOI221_X1 U18728 ( .B1(READY1), .B2(keyinput_36), .C1(keyinput_37), .C2(
        READY2), .A(n16828), .ZN(n16834) );
  INV_X1 U18729 ( .A(NA), .ZN(n21759) );
  AOI22_X1 U18730 ( .A1(BS16), .A2(keyinput_35), .B1(n21759), .B2(keyinput_34), 
        .ZN(n16829) );
  OAI221_X1 U18731 ( .B1(BS16), .B2(keyinput_35), .C1(n21759), .C2(keyinput_34), .A(n16829), .ZN(n16833) );
  INV_X1 U18732 ( .A(P1_READREQUEST_REG_SCAN_IN), .ZN(n16831) );
  AOI22_X1 U18733 ( .A1(P1_CODEFETCH_REG_SCAN_IN), .A2(keyinput_40), .B1(
        n16831), .B2(keyinput_38), .ZN(n16830) );
  OAI221_X1 U18734 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(keyinput_40), .C1(
        n16831), .C2(keyinput_38), .A(n16830), .ZN(n16832) );
  AOI221_X1 U18735 ( .B1(n16835), .B2(n16834), .C1(n16833), .C2(n16834), .A(
        n16832), .ZN(n16838) );
  OAI22_X1 U18736 ( .A1(n22220), .A2(keyinput_41), .B1(P1_D_C_N_REG_SCAN_IN), 
        .B2(keyinput_42), .ZN(n16836) );
  AOI221_X1 U18737 ( .B1(n22220), .B2(keyinput_41), .C1(keyinput_42), .C2(
        P1_D_C_N_REG_SCAN_IN), .A(n16836), .ZN(n16837) );
  OAI211_X1 U18738 ( .C1(P1_ADS_N_REG_SCAN_IN), .C2(keyinput_39), .A(n16838), 
        .B(n16837), .ZN(n16839) );
  AOI21_X1 U18739 ( .B1(P1_ADS_N_REG_SCAN_IN), .B2(keyinput_39), .A(n16839), 
        .ZN(n16840) );
  OAI22_X1 U18740 ( .A1(keyinput_45), .A2(n16948), .B1(n16841), .B2(n16840), 
        .ZN(n16842) );
  AOI21_X1 U18741 ( .B1(keyinput_45), .B2(n16948), .A(n16842), .ZN(n16845) );
  AOI22_X1 U18742 ( .A1(P1_BYTEENABLE_REG_0__SCAN_IN), .A2(keyinput_48), .B1(
        P1_W_R_N_REG_SCAN_IN), .B2(keyinput_47), .ZN(n16843) );
  OAI221_X1 U18743 ( .B1(P1_BYTEENABLE_REG_0__SCAN_IN), .B2(keyinput_48), .C1(
        P1_W_R_N_REG_SCAN_IN), .C2(keyinput_47), .A(n16843), .ZN(n16844) );
  AOI211_X1 U18744 ( .C1(P1_FLUSH_REG_SCAN_IN), .C2(keyinput_46), .A(n16845), 
        .B(n16844), .ZN(n16846) );
  OAI21_X1 U18745 ( .B1(P1_FLUSH_REG_SCAN_IN), .B2(keyinput_46), .A(n16846), 
        .ZN(n16847) );
  OAI221_X1 U18746 ( .B1(P1_BYTEENABLE_REG_1__SCAN_IN), .B2(n16848), .C1(
        n19954), .C2(keyinput_49), .A(n16847), .ZN(n16849) );
  OAI221_X1 U18747 ( .B1(P1_BYTEENABLE_REG_2__SCAN_IN), .B2(keyinput_50), .C1(
        n19950), .C2(n16850), .A(n16849), .ZN(n16851) );
  OAI221_X1 U18748 ( .B1(P1_BYTEENABLE_REG_3__SCAN_IN), .B2(keyinput_51), .C1(
        n19934), .C2(n16852), .A(n16851), .ZN(n16855) );
  INV_X1 U18749 ( .A(P1_REIP_REG_28__SCAN_IN), .ZN(n19924) );
  AOI22_X1 U18750 ( .A1(P1_REIP_REG_29__SCAN_IN), .A2(keyinput_54), .B1(n19924), .B2(keyinput_55), .ZN(n16853) );
  OAI221_X1 U18751 ( .B1(P1_REIP_REG_29__SCAN_IN), .B2(keyinput_54), .C1(
        n19924), .C2(keyinput_55), .A(n16853), .ZN(n16854) );
  AOI21_X1 U18752 ( .B1(n16856), .B2(n16855), .A(n16854), .ZN(n16859) );
  AOI22_X1 U18753 ( .A1(n21385), .A2(keyinput_56), .B1(keyinput_58), .B2(
        n19919), .ZN(n16857) );
  OAI221_X1 U18754 ( .B1(n21385), .B2(keyinput_56), .C1(n19919), .C2(
        keyinput_58), .A(n16857), .ZN(n16858) );
  AOI211_X1 U18755 ( .C1(P1_REIP_REG_26__SCAN_IN), .C2(keyinput_57), .A(n16859), .B(n16858), .ZN(n16860) );
  OAI21_X1 U18756 ( .B1(P1_REIP_REG_26__SCAN_IN), .B2(keyinput_57), .A(n16860), 
        .ZN(n16861) );
  OAI221_X1 U18757 ( .B1(P1_REIP_REG_24__SCAN_IN), .B2(keyinput_59), .C1(
        n19915), .C2(n16862), .A(n16861), .ZN(n16863) );
  OAI221_X1 U18758 ( .B1(P1_REIP_REG_23__SCAN_IN), .B2(n16864), .C1(n19913), 
        .C2(keyinput_60), .A(n16863), .ZN(n16865) );
  OAI211_X1 U18759 ( .C1(P1_REIP_REG_21__SCAN_IN), .C2(keyinput_62), .A(n16866), .B(n16865), .ZN(n16867) );
  AOI21_X1 U18760 ( .B1(P1_REIP_REG_21__SCAN_IN), .B2(keyinput_62), .A(n16867), 
        .ZN(n16974) );
  INV_X1 U18761 ( .A(keyinput_124), .ZN(n16969) );
  INV_X1 U18762 ( .A(keyinput_123), .ZN(n16967) );
  OAI22_X1 U18763 ( .A1(n21385), .A2(keyinput_120), .B1(keyinput_122), .B2(
        P1_REIP_REG_25__SCAN_IN), .ZN(n16868) );
  AOI221_X1 U18764 ( .B1(n21385), .B2(keyinput_120), .C1(
        P1_REIP_REG_25__SCAN_IN), .C2(keyinput_122), .A(n16868), .ZN(n16964)
         );
  INV_X1 U18765 ( .A(keyinput_115), .ZN(n16957) );
  INV_X1 U18766 ( .A(keyinput_114), .ZN(n16955) );
  INV_X1 U18767 ( .A(keyinput_113), .ZN(n16953) );
  INV_X1 U18768 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n19957) );
  OAI22_X1 U18769 ( .A1(n20102), .A2(keyinput_111), .B1(n19957), .B2(
        keyinput_112), .ZN(n16869) );
  AOI221_X1 U18770 ( .B1(n20102), .B2(keyinput_111), .C1(keyinput_112), .C2(
        n19957), .A(n16869), .ZN(n16950) );
  INV_X1 U18771 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n21714) );
  OAI22_X1 U18772 ( .A1(n21714), .A2(keyinput_107), .B1(keyinput_108), .B2(
        P1_STATEBS16_REG_SCAN_IN), .ZN(n16870) );
  AOI221_X1 U18773 ( .B1(n21714), .B2(keyinput_107), .C1(
        P1_STATEBS16_REG_SCAN_IN), .C2(keyinput_108), .A(n16870), .ZN(n16946)
         );
  XNOR2_X1 U18774 ( .A(DATAI_3_), .B(keyinput_93), .ZN(n16932) );
  INV_X1 U18775 ( .A(keyinput_92), .ZN(n16924) );
  OAI22_X1 U18776 ( .A1(n16872), .A2(keyinput_86), .B1(keyinput_85), .B2(
        DATAI_11_), .ZN(n16871) );
  AOI221_X1 U18777 ( .B1(n16872), .B2(keyinput_86), .C1(DATAI_11_), .C2(
        keyinput_85), .A(n16871), .ZN(n16919) );
  XNOR2_X1 U18778 ( .A(keyinput_70), .B(n16873), .ZN(n16884) );
  INV_X1 U18779 ( .A(keyinput_69), .ZN(n16881) );
  OAI22_X1 U18780 ( .A1(DATAI_31_), .A2(keyinput_65), .B1(keyinput_64), .B2(
        P1_MEMORYFETCH_REG_SCAN_IN), .ZN(n16874) );
  AOI221_X1 U18781 ( .B1(DATAI_31_), .B2(keyinput_65), .C1(
        P1_MEMORYFETCH_REG_SCAN_IN), .C2(keyinput_64), .A(n16874), .ZN(n16878)
         );
  OAI22_X1 U18782 ( .A1(DATAI_29_), .A2(keyinput_67), .B1(DATAI_28_), .B2(
        keyinput_68), .ZN(n16875) );
  AOI221_X1 U18783 ( .B1(DATAI_29_), .B2(keyinput_67), .C1(keyinput_68), .C2(
        DATAI_28_), .A(n16875), .ZN(n16876) );
  OAI21_X1 U18784 ( .B1(n16879), .B2(keyinput_66), .A(n16876), .ZN(n16877) );
  AOI211_X1 U18785 ( .C1(n16879), .C2(keyinput_66), .A(n16878), .B(n16877), 
        .ZN(n16880) );
  AOI221_X1 U18786 ( .B1(DATAI_27_), .B2(keyinput_69), .C1(n16882), .C2(n16881), .A(n16880), .ZN(n16883) );
  OAI22_X1 U18787 ( .A1(n16884), .A2(n16883), .B1(n16886), .B2(keyinput_73), 
        .ZN(n16885) );
  AOI21_X1 U18788 ( .B1(n16886), .B2(keyinput_73), .A(n16885), .ZN(n16892) );
  OAI22_X1 U18789 ( .A1(DATAI_25_), .A2(keyinput_71), .B1(keyinput_72), .B2(
        DATAI_24_), .ZN(n16887) );
  AOI221_X1 U18790 ( .B1(DATAI_25_), .B2(keyinput_71), .C1(DATAI_24_), .C2(
        keyinput_72), .A(n16887), .ZN(n16891) );
  AOI22_X1 U18791 ( .A1(DATAI_20_), .A2(keyinput_76), .B1(n16889), .B2(
        keyinput_77), .ZN(n16888) );
  OAI221_X1 U18792 ( .B1(DATAI_20_), .B2(keyinput_76), .C1(n16889), .C2(
        keyinput_77), .A(n16888), .ZN(n16890) );
  AOI21_X1 U18793 ( .B1(n16892), .B2(n16891), .A(n16890), .ZN(n16897) );
  OAI22_X1 U18794 ( .A1(n16895), .A2(keyinput_74), .B1(n16894), .B2(
        keyinput_75), .ZN(n16893) );
  AOI221_X1 U18795 ( .B1(n16895), .B2(keyinput_74), .C1(keyinput_75), .C2(
        n16894), .A(n16893), .ZN(n16896) );
  AOI22_X1 U18796 ( .A1(n16897), .A2(n16896), .B1(keyinput_78), .B2(n16899), 
        .ZN(n16898) );
  OAI21_X1 U18797 ( .B1(keyinput_78), .B2(n16899), .A(n16898), .ZN(n16909) );
  AOI22_X1 U18798 ( .A1(DATAI_16_), .A2(keyinput_80), .B1(DATAI_17_), .B2(
        keyinput_79), .ZN(n16900) );
  OAI221_X1 U18799 ( .B1(DATAI_16_), .B2(keyinput_80), .C1(DATAI_17_), .C2(
        keyinput_79), .A(n16900), .ZN(n16908) );
  OAI22_X1 U18800 ( .A1(n16903), .A2(keyinput_83), .B1(n16902), .B2(
        keyinput_84), .ZN(n16901) );
  AOI221_X1 U18801 ( .B1(n16903), .B2(keyinput_83), .C1(keyinput_84), .C2(
        n16902), .A(n16901), .ZN(n16907) );
  OAI22_X1 U18802 ( .A1(n16905), .A2(keyinput_82), .B1(DATAI_15_), .B2(
        keyinput_81), .ZN(n16904) );
  AOI221_X1 U18803 ( .B1(n16905), .B2(keyinput_82), .C1(keyinput_81), .C2(
        DATAI_15_), .A(n16904), .ZN(n16906) );
  OAI211_X1 U18804 ( .C1(n16909), .C2(n16908), .A(n16907), .B(n16906), .ZN(
        n16918) );
  AOI22_X1 U18805 ( .A1(n16912), .A2(keyinput_89), .B1(n16911), .B2(
        keyinput_88), .ZN(n16910) );
  OAI221_X1 U18806 ( .B1(n16912), .B2(keyinput_89), .C1(n16911), .C2(
        keyinput_88), .A(n16910), .ZN(n16917) );
  AOI22_X1 U18807 ( .A1(n16915), .A2(keyinput_87), .B1(keyinput_90), .B2(
        n16914), .ZN(n16913) );
  OAI221_X1 U18808 ( .B1(n16915), .B2(keyinput_87), .C1(n16914), .C2(
        keyinput_90), .A(n16913), .ZN(n16916) );
  AOI211_X1 U18809 ( .C1(n16919), .C2(n16918), .A(n16917), .B(n16916), .ZN(
        n16921) );
  NAND2_X1 U18810 ( .A1(DATAI_5_), .A2(keyinput_91), .ZN(n16920) );
  OAI211_X1 U18811 ( .C1(DATAI_5_), .C2(keyinput_91), .A(n16921), .B(n16920), 
        .ZN(n16922) );
  OAI221_X1 U18812 ( .B1(DATAI_4_), .B2(n16924), .C1(n16923), .C2(keyinput_92), 
        .A(n16922), .ZN(n16931) );
  AOI22_X1 U18813 ( .A1(n16927), .A2(keyinput_96), .B1(n16926), .B2(
        keyinput_95), .ZN(n16925) );
  OAI221_X1 U18814 ( .B1(n16927), .B2(keyinput_96), .C1(n16926), .C2(
        keyinput_95), .A(n16925), .ZN(n16930) );
  AOI22_X1 U18815 ( .A1(HOLD), .A2(keyinput_97), .B1(DATAI_2_), .B2(
        keyinput_94), .ZN(n16928) );
  OAI221_X1 U18816 ( .B1(HOLD), .B2(keyinput_97), .C1(DATAI_2_), .C2(
        keyinput_94), .A(n16928), .ZN(n16929) );
  AOI211_X1 U18817 ( .C1(n16932), .C2(n16931), .A(n16930), .B(n16929), .ZN(
        n16940) );
  INV_X1 U18818 ( .A(READY2), .ZN(n16934) );
  OAI22_X1 U18819 ( .A1(n16934), .A2(keyinput_101), .B1(keyinput_100), .B2(
        READY1), .ZN(n16933) );
  AOI221_X1 U18820 ( .B1(n16934), .B2(keyinput_101), .C1(READY1), .C2(
        keyinput_100), .A(n16933), .ZN(n16939) );
  AOI22_X1 U18821 ( .A1(BS16), .A2(keyinput_99), .B1(NA), .B2(keyinput_98), 
        .ZN(n16935) );
  OAI221_X1 U18822 ( .B1(BS16), .B2(keyinput_99), .C1(NA), .C2(keyinput_98), 
        .A(n16935), .ZN(n16938) );
  AOI22_X1 U18823 ( .A1(P1_D_C_N_REG_SCAN_IN), .A2(keyinput_106), .B1(n22220), 
        .B2(keyinput_105), .ZN(n16936) );
  OAI221_X1 U18824 ( .B1(P1_D_C_N_REG_SCAN_IN), .B2(keyinput_106), .C1(n22220), 
        .C2(keyinput_105), .A(n16936), .ZN(n16937) );
  AOI221_X1 U18825 ( .B1(n16940), .B2(n16939), .C1(n16938), .C2(n16939), .A(
        n16937), .ZN(n16944) );
  INV_X1 U18826 ( .A(P1_CODEFETCH_REG_SCAN_IN), .ZN(n20031) );
  AOI22_X1 U18827 ( .A1(P1_ADS_N_REG_SCAN_IN), .A2(keyinput_103), .B1(n20031), 
        .B2(keyinput_104), .ZN(n16941) );
  OAI221_X1 U18828 ( .B1(P1_ADS_N_REG_SCAN_IN), .B2(keyinput_103), .C1(n20031), 
        .C2(keyinput_104), .A(n16941), .ZN(n16942) );
  AOI21_X1 U18829 ( .B1(P1_READREQUEST_REG_SCAN_IN), .B2(keyinput_102), .A(
        n16942), .ZN(n16943) );
  OAI211_X1 U18830 ( .C1(P1_READREQUEST_REG_SCAN_IN), .C2(keyinput_102), .A(
        n16944), .B(n16943), .ZN(n16945) );
  AOI22_X1 U18831 ( .A1(keyinput_109), .A2(n16948), .B1(n16946), .B2(n16945), 
        .ZN(n16947) );
  OAI21_X1 U18832 ( .B1(n16948), .B2(keyinput_109), .A(n16947), .ZN(n16949) );
  OAI211_X1 U18833 ( .C1(P1_FLUSH_REG_SCAN_IN), .C2(keyinput_110), .A(n16950), 
        .B(n16949), .ZN(n16951) );
  AOI21_X1 U18834 ( .B1(P1_FLUSH_REG_SCAN_IN), .B2(keyinput_110), .A(n16951), 
        .ZN(n16952) );
  AOI221_X1 U18835 ( .B1(P1_BYTEENABLE_REG_1__SCAN_IN), .B2(keyinput_113), 
        .C1(n19954), .C2(n16953), .A(n16952), .ZN(n16954) );
  AOI221_X1 U18836 ( .B1(P1_BYTEENABLE_REG_2__SCAN_IN), .B2(keyinput_114), 
        .C1(n19950), .C2(n16955), .A(n16954), .ZN(n16956) );
  AOI221_X1 U18837 ( .B1(P1_BYTEENABLE_REG_3__SCAN_IN), .B2(n16957), .C1(
        n19934), .C2(keyinput_115), .A(n16956), .ZN(n16962) );
  AOI22_X1 U18838 ( .A1(P1_REIP_REG_30__SCAN_IN), .A2(keyinput_117), .B1(
        n19929), .B2(keyinput_116), .ZN(n16958) );
  OAI221_X1 U18839 ( .B1(P1_REIP_REG_30__SCAN_IN), .B2(keyinput_117), .C1(
        n19929), .C2(keyinput_116), .A(n16958), .ZN(n16961) );
  OAI22_X1 U18840 ( .A1(n19925), .A2(keyinput_118), .B1(keyinput_119), .B2(
        P1_REIP_REG_28__SCAN_IN), .ZN(n16959) );
  AOI221_X1 U18841 ( .B1(n19925), .B2(keyinput_118), .C1(
        P1_REIP_REG_28__SCAN_IN), .C2(keyinput_119), .A(n16959), .ZN(n16960)
         );
  OAI21_X1 U18842 ( .B1(n16962), .B2(n16961), .A(n16960), .ZN(n16963) );
  OAI211_X1 U18843 ( .C1(P1_REIP_REG_26__SCAN_IN), .C2(keyinput_121), .A(
        n16964), .B(n16963), .ZN(n16965) );
  AOI21_X1 U18844 ( .B1(P1_REIP_REG_26__SCAN_IN), .B2(keyinput_121), .A(n16965), .ZN(n16966) );
  AOI221_X1 U18845 ( .B1(P1_REIP_REG_24__SCAN_IN), .B2(keyinput_123), .C1(
        n19915), .C2(n16967), .A(n16966), .ZN(n16968) );
  AOI221_X1 U18846 ( .B1(P1_REIP_REG_23__SCAN_IN), .B2(keyinput_124), .C1(
        n19913), .C2(n16969), .A(n16968), .ZN(n16973) );
  XNOR2_X1 U18847 ( .A(P1_REIP_REG_21__SCAN_IN), .B(keyinput_126), .ZN(n16972)
         );
  INV_X1 U18848 ( .A(P1_REIP_REG_20__SCAN_IN), .ZN(n19909) );
  AOI22_X1 U18849 ( .A1(n21615), .A2(keyinput_125), .B1(n19909), .B2(
        keyinput_127), .ZN(n16970) );
  OAI221_X1 U18850 ( .B1(n21615), .B2(keyinput_125), .C1(n19909), .C2(
        keyinput_127), .A(n16970), .ZN(n16971) );
  NOR4_X1 U18851 ( .A1(n16974), .A2(n16973), .A3(n16972), .A4(n16971), .ZN(
        n16975) );
  XNOR2_X1 U18852 ( .A(n16976), .B(n16975), .ZN(P1_U3180) );
  INV_X1 U18853 ( .A(P2_CODEFETCH_REG_SCAN_IN), .ZN(n16977) );
  OAI22_X1 U18854 ( .A1(n18095), .A2(n16977), .B1(n18636), .B2(n18628), .ZN(
        P2_U2816) );
  OAI21_X1 U18855 ( .B1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n16979), .A(
        n16978), .ZN(n18158) );
  AOI22_X1 U18856 ( .A1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n17052), .B1(
        P2_REIP_REG_5__SCAN_IN), .B2(n18572), .ZN(n16985) );
  INV_X1 U18857 ( .A(n18149), .ZN(n16983) );
  OAI22_X1 U18858 ( .A1(n16981), .A2(n17042), .B1(n17058), .B2(n16980), .ZN(
        n16982) );
  AOI21_X1 U18859 ( .B1(n17019), .B2(n16983), .A(n16982), .ZN(n16984) );
  OAI211_X1 U18860 ( .C1(n17046), .C2(n18158), .A(n16985), .B(n16984), .ZN(
        P2_U3009) );
  AOI21_X1 U18861 ( .B1(n16999), .B2(n16987), .A(n16986), .ZN(n18194) );
  AOI22_X1 U18862 ( .A1(P2_REIP_REG_8__SCAN_IN), .A2(n18572), .B1(n17055), 
        .B2(n18194), .ZN(n16998) );
  NAND2_X1 U18863 ( .A1(n16989), .A2(n16988), .ZN(n16994) );
  INV_X1 U18864 ( .A(n16990), .ZN(n16991) );
  AOI21_X1 U18865 ( .B1(n16398), .B2(n16992), .A(n16991), .ZN(n16993) );
  XOR2_X1 U18866 ( .A(n16994), .B(n16993), .Z(n18571) );
  INV_X1 U18867 ( .A(n18192), .ZN(n18570) );
  XOR2_X1 U18868 ( .A(n16996), .B(n16995), .Z(n18569) );
  AOI222_X1 U18869 ( .A1(n18571), .A2(n17039), .B1(n17019), .B2(n18570), .C1(
        n18569), .C2(n17047), .ZN(n16997) );
  OAI211_X1 U18870 ( .C1(n16999), .C2(n17022), .A(n16998), .B(n16997), .ZN(
        P2_U3006) );
  AOI21_X1 U18871 ( .B1(n17007), .B2(n17000), .A(n17008), .ZN(n18211) );
  AOI22_X1 U18872 ( .A1(P2_REIP_REG_9__SCAN_IN), .A2(n18572), .B1(n17055), 
        .B2(n18211), .ZN(n17006) );
  OAI22_X1 U18873 ( .A1(n17002), .A2(n17042), .B1(n17058), .B2(n17001), .ZN(
        n17003) );
  AOI21_X1 U18874 ( .B1(n17019), .B2(n17004), .A(n17003), .ZN(n17005) );
  OAI211_X1 U18875 ( .C1(n17007), .C2(n17022), .A(n17006), .B(n17005), .ZN(
        P2_U3005) );
  OAI21_X1 U18876 ( .B1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n17008), .A(
        n17014), .ZN(n18210) );
  AOI22_X1 U18877 ( .A1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n17052), .B1(
        P2_REIP_REG_10__SCAN_IN), .B2(n18572), .ZN(n17013) );
  AOI222_X1 U18878 ( .A1(n17011), .A2(n17039), .B1(n17019), .B2(n17010), .C1(
        n17047), .C2(n17009), .ZN(n17012) );
  OAI211_X1 U18879 ( .C1(n17046), .C2(n18210), .A(n17013), .B(n17012), .ZN(
        P2_U3004) );
  AOI21_X1 U18880 ( .B1(n17023), .B2(n17014), .A(n17025), .ZN(n18241) );
  AOI22_X1 U18881 ( .A1(P2_REIP_REG_11__SCAN_IN), .A2(n18572), .B1(n17055), 
        .B2(n18241), .ZN(n17021) );
  OAI22_X1 U18882 ( .A1(n17016), .A2(n17042), .B1(n17015), .B2(n17058), .ZN(
        n17017) );
  AOI21_X1 U18883 ( .B1(n17019), .B2(n17018), .A(n17017), .ZN(n17020) );
  OAI211_X1 U18884 ( .C1(n17023), .C2(n17022), .A(n17021), .B(n17020), .ZN(
        P2_U3003) );
  OAI21_X1 U18885 ( .B1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n17025), .A(
        n17024), .ZN(n18240) );
  AOI22_X1 U18886 ( .A1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n17052), .B1(
        P2_REIP_REG_12__SCAN_IN), .B2(n18572), .ZN(n17030) );
  OAI22_X1 U18887 ( .A1(n17026), .A2(n17058), .B1(n17062), .B2(n18249), .ZN(
        n17027) );
  AOI21_X1 U18888 ( .B1(n17028), .B2(n17047), .A(n17027), .ZN(n17029) );
  OAI211_X1 U18889 ( .C1(n17046), .C2(n18240), .A(n17030), .B(n17029), .ZN(
        P2_U3002) );
  OAI21_X1 U18890 ( .B1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n11042), .A(
        n17031), .ZN(n18270) );
  AOI22_X1 U18891 ( .A1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n17052), .B1(
        P2_REIP_REG_14__SCAN_IN), .B2(n18572), .ZN(n17045) );
  NAND2_X1 U18892 ( .A1(n17032), .A2(n15191), .ZN(n17034) );
  NAND2_X1 U18893 ( .A1(n17034), .A2(n17033), .ZN(n18543) );
  OR2_X1 U18894 ( .A1(n17036), .A2(n17035), .ZN(n17037) );
  NAND2_X1 U18895 ( .A1(n17038), .A2(n17037), .ZN(n18539) );
  NAND2_X1 U18896 ( .A1(n18539), .A2(n17039), .ZN(n17041) );
  OR2_X1 U18897 ( .A1(n18540), .A2(n17062), .ZN(n17040) );
  OAI211_X1 U18898 ( .C1(n18543), .C2(n17042), .A(n17041), .B(n17040), .ZN(
        n17043) );
  INV_X1 U18899 ( .A(n17043), .ZN(n17044) );
  OAI211_X1 U18900 ( .C1(n17046), .C2(n18270), .A(n17045), .B(n17044), .ZN(
        P2_U3000) );
  OAI211_X1 U18901 ( .C1(n11013), .C2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n17048), .B(n17047), .ZN(n17057) );
  OAI21_X1 U18902 ( .B1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n17050), .A(
        n17049), .ZN(n17051) );
  INV_X1 U18903 ( .A(n17051), .ZN(n18303) );
  AOI22_X1 U18904 ( .A1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n17052), .B1(
        P2_REIP_REG_16__SCAN_IN), .B2(n18572), .ZN(n17053) );
  INV_X1 U18905 ( .A(n17053), .ZN(n17054) );
  AOI21_X1 U18906 ( .B1(n18303), .B2(n17055), .A(n17054), .ZN(n17056) );
  OAI211_X1 U18907 ( .C1(n17059), .C2(n17058), .A(n17057), .B(n17056), .ZN(
        n17060) );
  INV_X1 U18908 ( .A(n17060), .ZN(n17061) );
  OAI21_X1 U18909 ( .B1(n17062), .B2(n18301), .A(n17061), .ZN(P2_U2998) );
  INV_X1 U18910 ( .A(n17063), .ZN(n17065) );
  OAI22_X1 U18911 ( .A1(n19147), .A2(n18098), .B1(n17065), .B2(n17064), .ZN(
        n17066) );
  AOI21_X1 U18912 ( .B1(n19323), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n17066), 
        .ZN(n17067) );
  OAI22_X1 U18913 ( .A1(n19323), .A2(n17080), .B1(n17082), .B2(n17067), .ZN(
        P2_U3605) );
  NAND2_X1 U18914 ( .A1(n19168), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19295) );
  NAND2_X1 U18915 ( .A1(n19295), .A2(n19316), .ZN(n17073) );
  AND2_X1 U18916 ( .A1(n17073), .A2(n18628), .ZN(n17078) );
  NAND2_X1 U18917 ( .A1(n18621), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n17070) );
  INV_X1 U18918 ( .A(n19295), .ZN(n17068) );
  NAND3_X1 U18919 ( .A1(n19219), .A2(n19332), .A3(n17068), .ZN(n17069) );
  OAI211_X1 U18920 ( .C1(n17078), .C2(n19219), .A(n17070), .B(n17069), .ZN(
        n17071) );
  INV_X1 U18921 ( .A(n17071), .ZN(n17072) );
  AOI22_X1 U18922 ( .A1(n17082), .A2(n19231), .B1(n17072), .B2(n17080), .ZN(
        P2_U3603) );
  AOI21_X1 U18923 ( .B1(n21695), .B2(n19152), .A(n17073), .ZN(n17075) );
  OAI22_X1 U18924 ( .A1(n19152), .A2(n18628), .B1(n19203), .B2(n18116), .ZN(
        n17074) );
  NOR2_X1 U18925 ( .A1(n17075), .A2(n17074), .ZN(n17076) );
  AOI22_X1 U18926 ( .A1(n17082), .A2(n19296), .B1(n17076), .B2(n17080), .ZN(
        P2_U3604) );
  NOR2_X1 U18927 ( .A1(n21695), .A2(n19217), .ZN(n19197) );
  NOR2_X1 U18928 ( .A1(n19267), .A2(n19295), .ZN(n19245) );
  OAI22_X1 U18929 ( .A1(n19328), .A2(n17078), .B1(n19203), .B2(n18595), .ZN(
        n17079) );
  AOI221_X1 U18930 ( .B1(n19197), .B2(n19316), .C1(n19245), .C2(n19332), .A(
        n17079), .ZN(n17081) );
  AOI22_X1 U18931 ( .A1(n17082), .A2(n19200), .B1(n17081), .B2(n17080), .ZN(
        P2_U3602) );
  NAND2_X1 U18932 ( .A1(n17083), .A2(n21697), .ZN(n17086) );
  OAI21_X1 U18933 ( .B1(n12779), .B2(n18102), .A(n17089), .ZN(n17084) );
  OAI21_X1 U18934 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n17089), .A(n17084), 
        .ZN(n17085) );
  OAI221_X1 U18935 ( .B1(n17086), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n17086), .C2(P2_REIP_REG_0__SCAN_IN), .A(n17085), .ZN(P2_U2822) );
  INV_X1 U18936 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n17145) );
  OAI221_X1 U18937 ( .B1(n17089), .B2(n17145), .C1(n17088), .C2(n17087), .A(
        n17086), .ZN(P2_U2823) );
  INV_X1 U18938 ( .A(P2_M_IO_N_REG_SCAN_IN), .ZN(n17090) );
  AOI22_X1 U18939 ( .A1(n21734), .A2(n17091), .B1(n17090), .B2(n17143), .ZN(
        P2_U3611) );
  INV_X1 U18940 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n17092) );
  AOI22_X1 U18941 ( .A1(n21734), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n17092), 
        .B2(n17143), .ZN(P2_U3608) );
  INV_X1 U18942 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n21739) );
  INV_X1 U18943 ( .A(P2_ADS_N_REG_SCAN_IN), .ZN(n17094) );
  OAI21_X1 U18944 ( .B1(n21739), .B2(n17094), .A(n17093), .ZN(P2_U2815) );
  AOI22_X1 U18945 ( .A1(n17126), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n17114), 
        .B2(P2_DATAO_REG_0__SCAN_IN), .ZN(n17096) );
  OAI21_X1 U18946 ( .B1(n13675), .B2(n17128), .A(n17096), .ZN(P2_U2951) );
  INV_X1 U18947 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n17098) );
  AOI22_X1 U18948 ( .A1(n17126), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n17114), 
        .B2(P2_DATAO_REG_1__SCAN_IN), .ZN(n17097) );
  OAI21_X1 U18949 ( .B1(n17098), .B2(n17128), .A(n17097), .ZN(P2_U2950) );
  INV_X1 U18950 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n17100) );
  AOI22_X1 U18951 ( .A1(n17126), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n17114), 
        .B2(P2_DATAO_REG_2__SCAN_IN), .ZN(n17099) );
  OAI21_X1 U18952 ( .B1(n17100), .B2(n17128), .A(n17099), .ZN(P2_U2949) );
  INV_X1 U18953 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n17102) );
  AOI22_X1 U18954 ( .A1(n17115), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n17114), 
        .B2(P2_DATAO_REG_3__SCAN_IN), .ZN(n17101) );
  OAI21_X1 U18955 ( .B1(n17102), .B2(n17128), .A(n17101), .ZN(P2_U2948) );
  INV_X1 U18956 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n17104) );
  AOI22_X1 U18957 ( .A1(n17126), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n17114), 
        .B2(P2_DATAO_REG_4__SCAN_IN), .ZN(n17103) );
  OAI21_X1 U18958 ( .B1(n17104), .B2(n17128), .A(n17103), .ZN(P2_U2947) );
  INV_X1 U18959 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n19402) );
  AOI22_X1 U18960 ( .A1(n17115), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n17114), 
        .B2(P2_DATAO_REG_5__SCAN_IN), .ZN(n17105) );
  OAI21_X1 U18961 ( .B1(n19402), .B2(n17128), .A(n17105), .ZN(P2_U2946) );
  AOI22_X1 U18962 ( .A1(n17115), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n17114), 
        .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n17106) );
  OAI21_X1 U18963 ( .B1(n17107), .B2(n17128), .A(n17106), .ZN(P2_U2945) );
  AOI22_X1 U18964 ( .A1(n17115), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n17114), 
        .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n17108) );
  OAI21_X1 U18965 ( .B1(n17109), .B2(n17128), .A(n17108), .ZN(P2_U2944) );
  AOI22_X1 U18966 ( .A1(n17115), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n17114), 
        .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n17110) );
  OAI21_X1 U18967 ( .B1(n17111), .B2(n17128), .A(n17110), .ZN(P2_U2943) );
  AOI22_X1 U18968 ( .A1(n17126), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n17114), 
        .B2(P2_DATAO_REG_9__SCAN_IN), .ZN(n17112) );
  OAI21_X1 U18969 ( .B1(n17113), .B2(n17128), .A(n17112), .ZN(P2_U2942) );
  AOI22_X1 U18970 ( .A1(n17115), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(n17114), 
        .B2(P2_DATAO_REG_10__SCAN_IN), .ZN(n17116) );
  OAI21_X1 U18971 ( .B1(n17117), .B2(n17128), .A(n17116), .ZN(P2_U2941) );
  AOI22_X1 U18972 ( .A1(n17126), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n17114), 
        .B2(P2_DATAO_REG_11__SCAN_IN), .ZN(n17118) );
  OAI21_X1 U18973 ( .B1(n17119), .B2(n17128), .A(n17118), .ZN(P2_U2940) );
  AOI22_X1 U18974 ( .A1(n17126), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(n17114), 
        .B2(P2_DATAO_REG_12__SCAN_IN), .ZN(n17120) );
  OAI21_X1 U18975 ( .B1(n17121), .B2(n17128), .A(n17120), .ZN(P2_U2939) );
  AOI22_X1 U18976 ( .A1(n17126), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n17114), 
        .B2(P2_DATAO_REG_13__SCAN_IN), .ZN(n17122) );
  OAI21_X1 U18977 ( .B1(n17123), .B2(n17128), .A(n17122), .ZN(P2_U2938) );
  AOI22_X1 U18978 ( .A1(n17126), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n17114), 
        .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n17124) );
  OAI21_X1 U18979 ( .B1(n17125), .B2(n17128), .A(n17124), .ZN(P2_U2937) );
  AOI22_X1 U18980 ( .A1(n17126), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n17114), 
        .B2(P2_DATAO_REG_15__SCAN_IN), .ZN(n17127) );
  OAI21_X1 U18981 ( .B1(n17129), .B2(n17128), .A(n17127), .ZN(P2_U2936) );
  AOI21_X1 U18982 ( .B1(n21739), .B2(n17130), .A(P2_D_C_N_REG_SCAN_IN), .ZN(
        n17131) );
  AOI21_X1 U18983 ( .B1(P2_CODEFETCH_REG_SCAN_IN), .B2(n21734), .A(n17131), 
        .ZN(P2_U2817) );
  OAI222_X1 U18984 ( .A1(n17138), .A2(n12813), .B1(n19791), .B2(n21734), .C1(
        n12779), .C2(n17137), .ZN(P2_U3212) );
  INV_X1 U18985 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n17132) );
  INV_X1 U18986 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n19793) );
  OAI222_X1 U18987 ( .A1(n17138), .A2(n17132), .B1(n19793), .B2(n21734), .C1(
        n12813), .C2(n17137), .ZN(P2_U3213) );
  INV_X1 U18988 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n19795) );
  OAI222_X1 U18989 ( .A1(n17138), .A2(n13825), .B1(n19795), .B2(n21734), .C1(
        n17132), .C2(n17137), .ZN(P2_U3214) );
  INV_X1 U18990 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n19797) );
  OAI222_X1 U18991 ( .A1(n17138), .A2(n13830), .B1(n19797), .B2(n21734), .C1(
        n13825), .C2(n17137), .ZN(P2_U3215) );
  INV_X1 U18992 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n19799) );
  OAI222_X1 U18993 ( .A1(n17138), .A2(n13834), .B1(n19799), .B2(n21734), .C1(
        n13830), .C2(n17137), .ZN(P2_U3216) );
  INV_X1 U18994 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n19801) );
  OAI222_X1 U18995 ( .A1(n17138), .A2(n17133), .B1(n19801), .B2(n21734), .C1(
        n13834), .C2(n17137), .ZN(P2_U3217) );
  INV_X1 U18996 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n19803) );
  OAI222_X1 U18997 ( .A1(n17138), .A2(n13811), .B1(n19803), .B2(n21734), .C1(
        n17133), .C2(n17137), .ZN(P2_U3218) );
  INV_X1 U18998 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n19805) );
  OAI222_X1 U18999 ( .A1(n17138), .A2(n13853), .B1(n19805), .B2(n21734), .C1(
        n13811), .C2(n17137), .ZN(P2_U3219) );
  INV_X1 U19000 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n19807) );
  OAI222_X1 U19001 ( .A1(n17137), .A2(n13853), .B1(n19807), .B2(n21734), .C1(
        n13922), .C2(n17138), .ZN(P2_U3220) );
  INV_X1 U19002 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n19809) );
  OAI222_X1 U19003 ( .A1(n17137), .A2(n13922), .B1(n19809), .B2(n21734), .C1(
        n16574), .C2(n17138), .ZN(P2_U3221) );
  INV_X1 U19004 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n19811) );
  OAI222_X1 U19005 ( .A1(n17137), .A2(n16574), .B1(n19811), .B2(n21734), .C1(
        n14217), .C2(n17138), .ZN(P2_U3222) );
  INV_X1 U19006 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n19813) );
  OAI222_X1 U19007 ( .A1(n17137), .A2(n14217), .B1(n19813), .B2(n21734), .C1(
        n16391), .C2(n17138), .ZN(P2_U3223) );
  INV_X1 U19008 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n19815) );
  INV_X1 U19009 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n17134) );
  OAI222_X1 U19010 ( .A1(n17137), .A2(n16391), .B1(n19815), .B2(n21734), .C1(
        n17134), .C2(n17138), .ZN(P2_U3224) );
  INV_X1 U19011 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n19817) );
  INV_X1 U19012 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n17135) );
  OAI222_X1 U19013 ( .A1(n17137), .A2(n17134), .B1(n19817), .B2(n21734), .C1(
        n17135), .C2(n17138), .ZN(P2_U3225) );
  INV_X1 U19014 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n19819) );
  OAI222_X1 U19015 ( .A1(n17137), .A2(n17135), .B1(n19819), .B2(n21734), .C1(
        n14944), .C2(n17138), .ZN(P2_U3226) );
  INV_X1 U19016 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n19821) );
  OAI222_X1 U19017 ( .A1(n17137), .A2(n14944), .B1(n19821), .B2(n21734), .C1(
        n15067), .C2(n17138), .ZN(P2_U3227) );
  INV_X1 U19018 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n19823) );
  OAI222_X1 U19019 ( .A1(n17137), .A2(n15067), .B1(n19823), .B2(n21734), .C1(
        n16356), .C2(n17138), .ZN(P2_U3228) );
  INV_X1 U19020 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n17136) );
  INV_X1 U19021 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n19825) );
  OAI222_X1 U19022 ( .A1(n17138), .A2(n17136), .B1(n19825), .B2(n21734), .C1(
        n16356), .C2(n17137), .ZN(P2_U3229) );
  INV_X1 U19023 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n19827) );
  OAI222_X1 U19024 ( .A1(n17137), .A2(n17136), .B1(n19827), .B2(n21734), .C1(
        n18350), .C2(n17138), .ZN(P2_U3230) );
  INV_X1 U19025 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n19829) );
  OAI222_X1 U19026 ( .A1(n17138), .A2(n18358), .B1(n19829), .B2(n21734), .C1(
        n18350), .C2(n17137), .ZN(P2_U3231) );
  INV_X1 U19027 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n19831) );
  OAI222_X1 U19028 ( .A1(n17138), .A2(n18371), .B1(n19831), .B2(n21734), .C1(
        n18358), .C2(n17137), .ZN(P2_U3232) );
  INV_X1 U19029 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n18383) );
  INV_X1 U19030 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n19833) );
  OAI222_X1 U19031 ( .A1(n17138), .A2(n18383), .B1(n19833), .B2(n21734), .C1(
        n18371), .C2(n17137), .ZN(P2_U3233) );
  INV_X1 U19032 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n19835) );
  OAI222_X1 U19033 ( .A1(n17138), .A2(n18396), .B1(n19835), .B2(n21734), .C1(
        n18383), .C2(n17137), .ZN(P2_U3234) );
  INV_X1 U19034 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n19837) );
  OAI222_X1 U19035 ( .A1(n17138), .A2(n18410), .B1(n19837), .B2(n21734), .C1(
        n18396), .C2(n17137), .ZN(P2_U3235) );
  INV_X1 U19036 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n19840) );
  OAI222_X1 U19037 ( .A1(n17137), .A2(n18410), .B1(n19840), .B2(n21734), .C1(
        n18425), .C2(n17138), .ZN(P2_U3236) );
  INV_X1 U19038 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n19842) );
  OAI222_X1 U19039 ( .A1(n17138), .A2(n18438), .B1(n19842), .B2(n21734), .C1(
        n18425), .C2(n17137), .ZN(P2_U3237) );
  INV_X1 U19040 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n19844) );
  OAI222_X1 U19041 ( .A1(n17137), .A2(n18438), .B1(n19844), .B2(n21734), .C1(
        n18454), .C2(n17138), .ZN(P2_U3238) );
  INV_X1 U19042 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n19846) );
  OAI222_X1 U19043 ( .A1(n17137), .A2(n18454), .B1(n19846), .B2(n21734), .C1(
        n18468), .C2(n17138), .ZN(P2_U3239) );
  INV_X1 U19044 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n19848) );
  OAI222_X1 U19045 ( .A1(n17137), .A2(n18468), .B1(n19848), .B2(n21734), .C1(
        n18485), .C2(n17138), .ZN(P2_U3240) );
  INV_X1 U19046 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n19851) );
  OAI222_X1 U19047 ( .A1(n17138), .A2(n18501), .B1(n19851), .B2(n21734), .C1(
        n18485), .C2(n17137), .ZN(P2_U3241) );
  INV_X1 U19048 ( .A(P2_BE_N_REG_0__SCAN_IN), .ZN(n17139) );
  AOI22_X1 U19049 ( .A1(n21734), .A2(n17140), .B1(n17139), .B2(n17143), .ZN(
        P2_U3588) );
  INV_X1 U19050 ( .A(P2_BE_N_REG_1__SCAN_IN), .ZN(n17141) );
  AOI22_X1 U19051 ( .A1(n21734), .A2(n17142), .B1(n17141), .B2(n17143), .ZN(
        P2_U3587) );
  MUX2_X1 U19052 ( .A(P2_BE_N_REG_2__SCAN_IN), .B(P2_BYTEENABLE_REG_2__SCAN_IN), .S(n21734), .Z(P2_U3586) );
  INV_X1 U19053 ( .A(P2_BE_N_REG_3__SCAN_IN), .ZN(n17144) );
  AOI22_X1 U19054 ( .A1(n21734), .A2(n17145), .B1(n17144), .B2(n17143), .ZN(
        P2_U3585) );
  NAND3_X1 U19055 ( .A1(n20687), .A2(n18844), .A3(n17146), .ZN(n17147) );
  NAND2_X1 U19056 ( .A1(n17149), .A2(n20610), .ZN(n17525) );
  NAND2_X1 U19057 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n17521) );
  INV_X1 U19058 ( .A(n17521), .ZN(n17154) );
  AND2_X1 U19059 ( .A1(P3_EBX_REG_2__SCAN_IN), .A2(n17154), .ZN(n17150) );
  NAND3_X1 U19060 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(P3_EBX_REG_3__SCAN_IN), 
        .A3(n17150), .ZN(n17218) );
  NOR2_X1 U19061 ( .A1(n17525), .A2(n17218), .ZN(n17174) );
  INV_X1 U19062 ( .A(n17174), .ZN(n17188) );
  NOR2_X1 U19063 ( .A1(n20711), .A2(n17188), .ZN(n17239) );
  INV_X2 U19064 ( .A(n17526), .ZN(n17522) );
  NOR2_X1 U19065 ( .A1(n20711), .A2(n17525), .ZN(n17225) );
  AND2_X1 U19066 ( .A1(n17150), .A2(n17225), .ZN(n17155) );
  AND2_X1 U19067 ( .A1(P3_EBX_REG_3__SCAN_IN), .A2(n17155), .ZN(n17153) );
  AOI21_X1 U19068 ( .B1(P3_EBX_REG_4__SCAN_IN), .B2(n17522), .A(n17153), .ZN(
        n17151) );
  OAI22_X1 U19069 ( .A1(n17239), .A2(n17151), .B1(n17380), .B2(n17522), .ZN(
        P3_U2699) );
  AOI21_X1 U19070 ( .B1(P3_EBX_REG_3__SCAN_IN), .B2(n17522), .A(n17155), .ZN(
        n17152) );
  INV_X1 U19071 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17254) );
  OAI22_X1 U19072 ( .A1(n17153), .A2(n17152), .B1(n17254), .B2(n17522), .ZN(
        P3_U2700) );
  AOI21_X1 U19073 ( .B1(n17154), .B2(n17524), .A(P3_EBX_REG_2__SCAN_IN), .ZN(
        n17156) );
  AOI221_X1 U19074 ( .B1(n17156), .B2(n17522), .C1(n17369), .C2(n17526), .A(
        n17155), .ZN(P3_U2701) );
  AOI22_X1 U19075 ( .A1(n17546), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n17548), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n17160) );
  AOI22_X1 U19076 ( .A1(n17205), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n10966), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n17159) );
  AOI22_X1 U19077 ( .A1(n10968), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n14589), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n17158) );
  AOI22_X1 U19078 ( .A1(n17540), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n20216), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n17157) );
  NAND4_X1 U19079 ( .A1(n17160), .A2(n17159), .A3(n17158), .A4(n17157), .ZN(
        n17166) );
  AOI22_X1 U19080 ( .A1(n10958), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17286), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n17164) );
  AOI22_X1 U19081 ( .A1(n10972), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n10965), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n17163) );
  AOI22_X1 U19082 ( .A1(n10960), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n17505), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n17162) );
  AOI22_X1 U19083 ( .A1(n10967), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n17539), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n17161) );
  NAND4_X1 U19084 ( .A1(n17164), .A2(n17163), .A3(n17162), .A4(n17161), .ZN(
        n17165) );
  NOR2_X1 U19085 ( .A1(n17166), .A2(n17165), .ZN(n20782) );
  INV_X1 U19086 ( .A(P3_EBX_REG_8__SCAN_IN), .ZN(n20275) );
  NAND2_X1 U19087 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(P3_EBX_REG_5__SCAN_IN), 
        .ZN(n17187) );
  NOR2_X1 U19088 ( .A1(n17187), .A2(n17188), .ZN(n17168) );
  NAND2_X1 U19089 ( .A1(P3_EBX_REG_7__SCAN_IN), .A2(n17168), .ZN(n17293) );
  XNOR2_X1 U19090 ( .A(n20275), .B(n17293), .ZN(n17167) );
  AOI22_X1 U19091 ( .A1(n17526), .A2(n20782), .B1(n17167), .B2(n17522), .ZN(
        P3_U2695) );
  INV_X1 U19092 ( .A(n17168), .ZN(n17278) );
  INV_X1 U19093 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n17169) );
  OAI33_X1 U19094 ( .A1(P3_EBX_REG_7__SCAN_IN), .A2(n20711), .A3(n17278), .B1(
        n17169), .B2(n17526), .B3(n17168), .ZN(n17170) );
  AOI21_X1 U19095 ( .B1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B2(n17526), .A(
        n17170), .ZN(n17171) );
  INV_X1 U19096 ( .A(n17171), .ZN(P3_U2696) );
  NAND2_X1 U19097 ( .A1(P3_EBX_REG_5__SCAN_IN), .A2(n17239), .ZN(n17173) );
  NAND3_X1 U19098 ( .A1(n17173), .A2(P3_EBX_REG_6__SCAN_IN), .A3(n17522), .ZN(
        n17172) );
  OAI221_X1 U19099 ( .B1(n17173), .B2(P3_EBX_REG_6__SCAN_IN), .C1(n17522), 
        .C2(n17453), .A(n17172), .ZN(P3_U2697) );
  INV_X1 U19100 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n17176) );
  OAI211_X1 U19101 ( .C1(P3_EBX_REG_5__SCAN_IN), .C2(n17174), .A(n17173), .B(
        n17522), .ZN(n17175) );
  OAI21_X1 U19102 ( .B1(n17522), .B2(n17176), .A(n17175), .ZN(P3_U2698) );
  AOI22_X1 U19103 ( .A1(n17546), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n10967), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n17180) );
  AOI22_X1 U19104 ( .A1(n17205), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n17505), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n17179) );
  AOI22_X1 U19105 ( .A1(n17540), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n14589), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n17178) );
  AOI22_X1 U19106 ( .A1(n10968), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n20216), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n17177) );
  NAND4_X1 U19107 ( .A1(n17180), .A2(n17179), .A3(n17178), .A4(n17177), .ZN(
        n17186) );
  AOI22_X1 U19108 ( .A1(n17538), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17286), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n17184) );
  AOI22_X1 U19109 ( .A1(n10959), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17539), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n17183) );
  AOI22_X1 U19110 ( .A1(n10971), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17548), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n17182) );
  AOI22_X1 U19111 ( .A1(n17545), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n10965), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n17181) );
  NAND4_X1 U19112 ( .A1(n17184), .A2(n17183), .A3(n17182), .A4(n17181), .ZN(
        n17185) );
  NOR2_X1 U19113 ( .A1(n17186), .A2(n17185), .ZN(n20763) );
  INV_X1 U19114 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n20371) );
  INV_X1 U19115 ( .A(P3_EBX_REG_14__SCAN_IN), .ZN(n20362) );
  INV_X1 U19116 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n17224) );
  NOR2_X1 U19117 ( .A1(n20362), .A2(n17224), .ZN(n17297) );
  INV_X1 U19118 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n20316) );
  INV_X1 U19119 ( .A(P3_EBX_REG_10__SCAN_IN), .ZN(n20295) );
  NAND3_X1 U19120 ( .A1(P3_EBX_REG_9__SCAN_IN), .A2(P3_EBX_REG_8__SCAN_IN), 
        .A3(P3_EBX_REG_7__SCAN_IN), .ZN(n17279) );
  NOR4_X1 U19121 ( .A1(n20316), .A2(n20295), .A3(n17279), .A4(n17187), .ZN(
        n17240) );
  NAND2_X1 U19122 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n17240), .ZN(n17219) );
  NOR2_X1 U19123 ( .A1(n17219), .A2(n17188), .ZN(n17220) );
  NAND2_X1 U19124 ( .A1(n17297), .A2(n17220), .ZN(n17191) );
  NOR2_X1 U19125 ( .A1(n20371), .A2(n17191), .ZN(n17204) );
  NAND2_X1 U19126 ( .A1(n17204), .A2(P3_EBX_REG_16__SCAN_IN), .ZN(n17189) );
  OAI211_X1 U19127 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n17204), .A(n17522), .B(
        n17189), .ZN(n17190) );
  OAI21_X1 U19128 ( .B1(n20763), .B2(n17522), .A(n17190), .ZN(P3_U2687) );
  NAND2_X1 U19129 ( .A1(n20371), .A2(n17191), .ZN(n17192) );
  NAND2_X1 U19130 ( .A1(n17192), .A2(n17522), .ZN(n17203) );
  AOI22_X1 U19131 ( .A1(n10959), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n17505), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n17196) );
  AOI22_X1 U19132 ( .A1(n10967), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n17548), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n17195) );
  AOI22_X1 U19133 ( .A1(n10968), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n20216), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n17194) );
  AOI22_X1 U19134 ( .A1(n17540), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n14589), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n17193) );
  NAND4_X1 U19135 ( .A1(n17196), .A2(n17195), .A3(n17194), .A4(n17193), .ZN(
        n17202) );
  AOI22_X1 U19136 ( .A1(n10960), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n17286), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n17200) );
  AOI22_X1 U19137 ( .A1(n10972), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n10965), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n17199) );
  AOI22_X1 U19138 ( .A1(n17205), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n17539), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n17198) );
  AOI22_X1 U19139 ( .A1(n17546), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n10966), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n17197) );
  NAND4_X1 U19140 ( .A1(n17200), .A2(n17199), .A3(n17198), .A4(n17197), .ZN(
        n17201) );
  NOR2_X1 U19141 ( .A1(n17202), .A2(n17201), .ZN(n20774) );
  OAI22_X1 U19142 ( .A1(n17204), .A2(n17203), .B1(n20774), .B2(n17522), .ZN(
        P3_U2688) );
  AOI22_X1 U19143 ( .A1(n17205), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17546), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n17217) );
  AOI22_X1 U19144 ( .A1(n17505), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n10971), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n17216) );
  INV_X1 U19145 ( .A(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n17207) );
  AOI22_X1 U19146 ( .A1(n10967), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17539), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n17206) );
  OAI21_X1 U19147 ( .B1(n17208), .B2(n17207), .A(n17206), .ZN(n17214) );
  AOI22_X1 U19148 ( .A1(n10959), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17286), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n17212) );
  AOI22_X1 U19149 ( .A1(n14603), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10965), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n17211) );
  AOI22_X1 U19150 ( .A1(n17540), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n20216), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n17210) );
  AOI22_X1 U19151 ( .A1(n10968), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n14589), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n17209) );
  NAND4_X1 U19152 ( .A1(n17212), .A2(n17211), .A3(n17210), .A4(n17209), .ZN(
        n17213) );
  AOI211_X1 U19153 ( .C1(n10977), .C2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A(
        n17214), .B(n17213), .ZN(n17215) );
  NAND3_X1 U19154 ( .A1(n17217), .A2(n17216), .A3(n17215), .ZN(n20617) );
  NOR2_X1 U19155 ( .A1(n17219), .A2(n17218), .ZN(n17298) );
  INV_X1 U19156 ( .A(n17225), .ZN(n17528) );
  NOR2_X1 U19157 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(n17528), .ZN(n17221) );
  NOR2_X1 U19158 ( .A1(n17526), .A2(n17220), .ZN(n17223) );
  AOI222_X1 U19159 ( .A1(n20617), .A2(n17526), .B1(n17298), .B2(n17221), .C1(
        P3_EBX_REG_13__SCAN_IN), .C2(n17223), .ZN(n17222) );
  INV_X1 U19160 ( .A(n17222), .ZN(P3_U2690) );
  AOI21_X1 U19161 ( .B1(n17225), .B2(n17224), .A(n17223), .ZN(n17238) );
  NAND2_X1 U19162 ( .A1(n20362), .A2(n17238), .ZN(n17237) );
  AOI22_X1 U19163 ( .A1(n17539), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17286), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n17235) );
  AOI22_X1 U19164 ( .A1(n10958), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n10967), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n17234) );
  AOI22_X1 U19165 ( .A1(n17505), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17546), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n17226) );
  OAI21_X1 U19166 ( .B1(n14684), .B2(n17453), .A(n17226), .ZN(n17232) );
  AOI22_X1 U19167 ( .A1(n10971), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17548), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n17230) );
  AOI22_X1 U19168 ( .A1(n10960), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17538), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n17229) );
  AOI22_X1 U19169 ( .A1(n10968), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n20216), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n17228) );
  AOI22_X1 U19170 ( .A1(n17540), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n14589), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n17227) );
  NAND4_X1 U19171 ( .A1(n17230), .A2(n17229), .A3(n17228), .A4(n17227), .ZN(
        n17231) );
  AOI211_X1 U19172 ( .C1(n17205), .C2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A(
        n17232), .B(n17231), .ZN(n17233) );
  NAND3_X1 U19173 ( .A1(n17235), .A2(n17234), .A3(n17233), .ZN(n20765) );
  NAND2_X1 U19174 ( .A1(n17526), .A2(n20765), .ZN(n17236) );
  OAI221_X1 U19175 ( .B1(n20362), .B2(n17238), .C1(n17237), .C2(n20711), .A(
        n17236), .ZN(P3_U2689) );
  NAND2_X1 U19176 ( .A1(n17240), .A2(n17239), .ZN(n17252) );
  AOI22_X1 U19177 ( .A1(n10960), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n17546), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n17244) );
  AOI22_X1 U19178 ( .A1(n17547), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n10972), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n17243) );
  AOI22_X1 U19179 ( .A1(n10968), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17540), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n17242) );
  AOI22_X1 U19180 ( .A1(n14589), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n20216), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n17241) );
  NAND4_X1 U19181 ( .A1(n17244), .A2(n17243), .A3(n17242), .A4(n17241), .ZN(
        n17250) );
  AOI22_X1 U19182 ( .A1(n10971), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17548), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n17248) );
  AOI22_X1 U19183 ( .A1(n10967), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n10965), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17247) );
  AOI22_X1 U19184 ( .A1(n10959), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17539), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n17246) );
  AOI22_X1 U19185 ( .A1(n17505), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17286), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n17245) );
  NAND4_X1 U19186 ( .A1(n17248), .A2(n17247), .A3(n17246), .A4(n17245), .ZN(
        n17249) );
  NOR2_X1 U19187 ( .A1(n17250), .A2(n17249), .ZN(n20622) );
  NAND3_X1 U19188 ( .A1(n17252), .A2(P3_EBX_REG_12__SCAN_IN), .A3(n17522), 
        .ZN(n17251) );
  OAI221_X1 U19189 ( .B1(n17252), .B2(P3_EBX_REG_12__SCAN_IN), .C1(n17522), 
        .C2(n20622), .A(n17251), .ZN(P3_U2691) );
  NOR2_X1 U19190 ( .A1(n17279), .A2(n17278), .ZN(n17277) );
  AOI21_X1 U19191 ( .B1(P3_EBX_REG_10__SCAN_IN), .B2(n17277), .A(
        P3_EBX_REG_11__SCAN_IN), .ZN(n17266) );
  NAND2_X1 U19192 ( .A1(n17522), .A2(n17252), .ZN(n17265) );
  AOI22_X1 U19193 ( .A1(n17546), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n17548), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n17263) );
  AOI22_X1 U19194 ( .A1(n10959), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17539), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n17262) );
  AOI22_X1 U19195 ( .A1(n10966), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17286), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n17253) );
  OAI21_X1 U19196 ( .B1(n14684), .B2(n17254), .A(n17253), .ZN(n17260) );
  AOI22_X1 U19197 ( .A1(n17545), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n10967), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n17258) );
  AOI22_X1 U19198 ( .A1(n17205), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17505), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n17257) );
  AOI22_X1 U19199 ( .A1(n10968), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n20216), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n17256) );
  AOI22_X1 U19200 ( .A1(n17540), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n14589), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n17255) );
  NAND4_X1 U19201 ( .A1(n17258), .A2(n17257), .A3(n17256), .A4(n17255), .ZN(
        n17259) );
  AOI211_X1 U19202 ( .C1(n10972), .C2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A(
        n17260), .B(n17259), .ZN(n17261) );
  NAND3_X1 U19203 ( .A1(n17263), .A2(n17262), .A3(n17261), .ZN(n20625) );
  INV_X1 U19204 ( .A(n20625), .ZN(n17264) );
  OAI22_X1 U19205 ( .A1(n17266), .A2(n17265), .B1(n17264), .B2(n17522), .ZN(
        P3_U2692) );
  AOI22_X1 U19206 ( .A1(n10960), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n17538), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n17270) );
  AOI22_X1 U19207 ( .A1(n17205), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n17505), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n17269) );
  AOI22_X1 U19208 ( .A1(n17540), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n20216), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n17268) );
  AOI22_X1 U19209 ( .A1(n10968), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n14589), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n17267) );
  NAND4_X1 U19210 ( .A1(n17270), .A2(n17269), .A3(n17268), .A4(n17267), .ZN(
        n17276) );
  AOI22_X1 U19211 ( .A1(n17546), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n10967), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n17274) );
  AOI22_X1 U19212 ( .A1(n14603), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n10965), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17273) );
  AOI22_X1 U19213 ( .A1(n17539), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17286), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n17272) );
  AOI22_X1 U19214 ( .A1(n10958), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n10966), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n17271) );
  NAND4_X1 U19215 ( .A1(n17274), .A2(n17273), .A3(n17272), .A4(n17271), .ZN(
        n17275) );
  NOR2_X1 U19216 ( .A1(n17276), .A2(n17275), .ZN(n20629) );
  NOR2_X1 U19217 ( .A1(n17526), .A2(n17277), .ZN(n17294) );
  NOR3_X1 U19218 ( .A1(n20711), .A2(n17279), .A3(n17278), .ZN(n17280) );
  AOI22_X1 U19219 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n17294), .B1(n17280), 
        .B2(n20295), .ZN(n17281) );
  OAI21_X1 U19220 ( .B1(n20629), .B2(n17522), .A(n17281), .ZN(P3_U2693) );
  AOI22_X1 U19221 ( .A1(n10958), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_6__1__SCAN_IN), .B2(n14603), .ZN(n17285) );
  AOI22_X1 U19222 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n17539), .B1(
        n10967), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n17284) );
  AOI22_X1 U19223 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n17540), .B1(
        P3_INSTQUEUE_REG_5__1__SCAN_IN), .B2(n10968), .ZN(n17283) );
  AOI22_X1 U19224 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n14589), .B1(
        P3_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n20216), .ZN(n17282) );
  NAND4_X1 U19225 ( .A1(n17285), .A2(n17284), .A3(n17283), .A4(n17282), .ZN(
        n17292) );
  AOI22_X1 U19226 ( .A1(n10960), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_0__1__SCAN_IN), .B2(n10976), .ZN(n17290) );
  AOI22_X1 U19227 ( .A1(n17505), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n17286), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n17289) );
  AOI22_X1 U19228 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n10971), .B1(
        n17546), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n17288) );
  AOI22_X1 U19229 ( .A1(n17205), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_2__1__SCAN_IN), .B2(n17538), .ZN(n17287) );
  NAND4_X1 U19230 ( .A1(n17290), .A2(n17289), .A3(n17288), .A4(n17287), .ZN(
        n17291) );
  NOR2_X1 U19231 ( .A1(n17292), .A2(n17291), .ZN(n20634) );
  NOR2_X1 U19232 ( .A1(n20275), .A2(n17293), .ZN(n17295) );
  OAI21_X1 U19233 ( .B1(P3_EBX_REG_9__SCAN_IN), .B2(n17295), .A(n17294), .ZN(
        n17296) );
  OAI21_X1 U19234 ( .B1(n20634), .B2(n17522), .A(n17296), .ZN(P3_U2694) );
  INV_X1 U19235 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n20589) );
  AND3_X1 U19236 ( .A1(P3_EBX_REG_23__SCAN_IN), .A2(P3_EBX_REG_22__SCAN_IN), 
        .A3(P3_EBX_REG_21__SCAN_IN), .ZN(n17301) );
  INV_X1 U19237 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n20560) );
  INV_X1 U19238 ( .A(P3_EBX_REG_26__SCAN_IN), .ZN(n20515) );
  INV_X1 U19239 ( .A(P3_EBX_REG_20__SCAN_IN), .ZN(n20440) );
  INV_X1 U19240 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n17501) );
  INV_X1 U19241 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n17518) );
  NAND4_X1 U19242 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(P3_EBX_REG_15__SCAN_IN), 
        .A3(n17298), .A4(n17297), .ZN(n17517) );
  NOR2_X1 U19243 ( .A1(n17518), .A2(n17517), .ZN(n17516) );
  NAND2_X1 U19244 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n17489), .ZN(n17488) );
  NOR3_X1 U19245 ( .A1(n20440), .A2(n17501), .A3(n17488), .ZN(n17414) );
  INV_X1 U19246 ( .A(n17414), .ZN(n17415) );
  NAND2_X1 U19247 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(P3_EBX_REG_27__SCAN_IN), 
        .ZN(n17299) );
  NOR4_X1 U19248 ( .A1(n20560), .A2(n20515), .A3(n17415), .A4(n17299), .ZN(
        n17300) );
  NAND4_X1 U19249 ( .A1(P3_EBX_REG_25__SCAN_IN), .A2(P3_EBX_REG_24__SCAN_IN), 
        .A3(n17301), .A4(n17300), .ZN(n17304) );
  NOR2_X1 U19250 ( .A1(n20589), .A2(n17304), .ZN(n17403) );
  NAND2_X1 U19251 ( .A1(n17522), .A2(P3_EBX_REG_31__SCAN_IN), .ZN(n17303) );
  NAND2_X1 U19252 ( .A1(n17403), .A2(n20687), .ZN(n17302) );
  OAI22_X1 U19253 ( .A1(n17403), .A2(n17303), .B1(P3_EBX_REG_31__SCAN_IN), 
        .B2(n17302), .ZN(P3_U2672) );
  NAND2_X1 U19254 ( .A1(n20589), .A2(n17304), .ZN(n17305) );
  NAND2_X1 U19255 ( .A1(n17305), .A2(n17522), .ZN(n17402) );
  AOI22_X1 U19256 ( .A1(n17546), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n10965), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n17309) );
  AOI22_X1 U19257 ( .A1(n10966), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n17539), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n17308) );
  AOI22_X1 U19258 ( .A1(n10958), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n17505), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n17307) );
  AOI22_X1 U19259 ( .A1(n10960), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n10967), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n17306) );
  NAND4_X1 U19260 ( .A1(n17309), .A2(n17308), .A3(n17307), .A4(n17306), .ZN(
        n17315) );
  AOI22_X1 U19261 ( .A1(n10972), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n17537), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n17313) );
  AOI22_X1 U19262 ( .A1(n17205), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n17548), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n17312) );
  AOI22_X1 U19263 ( .A1(n10968), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n20216), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n17311) );
  AOI22_X1 U19264 ( .A1(n17540), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n14589), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n17310) );
  NAND4_X1 U19265 ( .A1(n17313), .A2(n17312), .A3(n17311), .A4(n17310), .ZN(
        n17314) );
  NOR2_X1 U19266 ( .A1(n17315), .A2(n17314), .ZN(n17401) );
  AOI22_X1 U19267 ( .A1(n10960), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17548), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n17319) );
  AOI22_X1 U19268 ( .A1(n17547), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n10958), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n17318) );
  AOI22_X1 U19269 ( .A1(n10968), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n20216), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n17317) );
  AOI22_X1 U19270 ( .A1(n17540), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n14589), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n17316) );
  NAND4_X1 U19271 ( .A1(n17319), .A2(n17318), .A3(n17317), .A4(n17316), .ZN(
        n17325) );
  AOI22_X1 U19272 ( .A1(n17505), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10967), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n17323) );
  AOI22_X1 U19273 ( .A1(n17546), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n17537), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n17322) );
  AOI22_X1 U19274 ( .A1(n17538), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17539), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n17321) );
  AOI22_X1 U19275 ( .A1(n10971), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n10965), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n17320) );
  NAND4_X1 U19276 ( .A1(n17323), .A2(n17322), .A3(n17321), .A4(n17320), .ZN(
        n17324) );
  NOR2_X1 U19277 ( .A1(n17325), .A2(n17324), .ZN(n17425) );
  AOI22_X1 U19278 ( .A1(n17546), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n10976), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n17329) );
  AOI22_X1 U19279 ( .A1(n17547), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n17539), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n17328) );
  AOI22_X1 U19280 ( .A1(n10968), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n14589), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n17327) );
  AOI22_X1 U19281 ( .A1(n17540), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n20216), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n17326) );
  NAND4_X1 U19282 ( .A1(n17329), .A2(n17328), .A3(n17327), .A4(n17326), .ZN(
        n17335) );
  AOI22_X1 U19283 ( .A1(n10967), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17548), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n17333) );
  AOI22_X1 U19284 ( .A1(n10959), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n10972), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n17332) );
  AOI22_X1 U19285 ( .A1(n17505), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17537), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n17331) );
  AOI22_X1 U19286 ( .A1(n10977), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n10966), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n17330) );
  NAND4_X1 U19287 ( .A1(n17333), .A2(n17332), .A3(n17331), .A4(n17330), .ZN(
        n17334) );
  NOR2_X1 U19288 ( .A1(n17335), .A2(n17334), .ZN(n17431) );
  AOI22_X1 U19289 ( .A1(n17538), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n10971), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n17339) );
  AOI22_X1 U19290 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n10975), .B1(
        n17546), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n17338) );
  AOI22_X1 U19291 ( .A1(n10968), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n17540), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n17337) );
  AOI22_X1 U19292 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n20216), .B1(
        P3_INSTQUEUE_REG_11__1__SCAN_IN), .B2(n14589), .ZN(n17336) );
  NAND4_X1 U19293 ( .A1(n17339), .A2(n17338), .A3(n17337), .A4(n17336), .ZN(
        n17345) );
  AOI22_X1 U19294 ( .A1(n17505), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_14__1__SCAN_IN), .B2(n17539), .ZN(n17343) );
  AOI22_X1 U19295 ( .A1(n10959), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_5__1__SCAN_IN), .B2(n17537), .ZN(n17342) );
  AOI22_X1 U19296 ( .A1(n10977), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_8__1__SCAN_IN), .B2(n14603), .ZN(n17341) );
  AOI22_X1 U19297 ( .A1(n17547), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_13__1__SCAN_IN), .B2(n10967), .ZN(n17340) );
  NAND4_X1 U19298 ( .A1(n17343), .A2(n17342), .A3(n17341), .A4(n17340), .ZN(
        n17344) );
  NOR2_X1 U19299 ( .A1(n17345), .A2(n17344), .ZN(n17441) );
  AOI22_X1 U19300 ( .A1(n17505), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10966), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n17356) );
  AOI22_X1 U19301 ( .A1(n10972), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17539), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n17355) );
  AOI22_X1 U19302 ( .A1(n10967), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10975), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n17346) );
  OAI21_X1 U19303 ( .B1(n17391), .B2(n17347), .A(n17346), .ZN(n17353) );
  AOI22_X1 U19304 ( .A1(n17545), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17537), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n17351) );
  AOI22_X1 U19305 ( .A1(n17547), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n17548), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n17350) );
  AOI22_X1 U19306 ( .A1(n17540), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n20216), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n17349) );
  AOI22_X1 U19307 ( .A1(n10968), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n14589), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n17348) );
  NAND4_X1 U19308 ( .A1(n17351), .A2(n17350), .A3(n17349), .A4(n17348), .ZN(
        n17352) );
  AOI211_X1 U19309 ( .C1(n10959), .C2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A(
        n17353), .B(n17352), .ZN(n17354) );
  NAND3_X1 U19310 ( .A1(n17356), .A2(n17355), .A3(n17354), .ZN(n17448) );
  AOI22_X1 U19311 ( .A1(n17538), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n17537), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n17367) );
  AOI22_X1 U19312 ( .A1(n14603), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n17539), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n17366) );
  INV_X1 U19313 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n17358) );
  AOI22_X1 U19314 ( .A1(n17546), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n10967), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n17357) );
  OAI21_X1 U19315 ( .B1(n11012), .B2(n17358), .A(n17357), .ZN(n17364) );
  AOI22_X1 U19316 ( .A1(n10958), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17505), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n17362) );
  AOI22_X1 U19317 ( .A1(n10966), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n10976), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n17361) );
  AOI22_X1 U19318 ( .A1(n17540), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n14589), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n17360) );
  AOI22_X1 U19319 ( .A1(n10968), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n20216), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n17359) );
  NAND4_X1 U19320 ( .A1(n17362), .A2(n17361), .A3(n17360), .A4(n17359), .ZN(
        n17363) );
  AOI211_X1 U19321 ( .C1(n10977), .C2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A(
        n17364), .B(n17363), .ZN(n17365) );
  NAND3_X1 U19322 ( .A1(n17367), .A2(n17366), .A3(n17365), .ZN(n17449) );
  NAND2_X1 U19323 ( .A1(n17448), .A2(n17449), .ZN(n17447) );
  NOR2_X1 U19324 ( .A1(n17441), .A2(n17447), .ZN(n17440) );
  AOI22_X1 U19325 ( .A1(n17547), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n10977), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n17378) );
  AOI22_X1 U19326 ( .A1(n10958), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17537), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n17377) );
  AOI22_X1 U19327 ( .A1(n10972), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n17548), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n17368) );
  OAI21_X1 U19328 ( .B1(n17391), .B2(n17369), .A(n17368), .ZN(n17375) );
  AOI22_X1 U19329 ( .A1(n10967), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n10971), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n17373) );
  AOI22_X1 U19330 ( .A1(n10976), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n17539), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n17372) );
  AOI22_X1 U19331 ( .A1(n17540), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n20216), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n17371) );
  AOI22_X1 U19332 ( .A1(n10968), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n14589), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n17370) );
  NAND4_X1 U19333 ( .A1(n17373), .A2(n17372), .A3(n17371), .A4(n17370), .ZN(
        n17374) );
  AOI211_X1 U19334 ( .C1(n17505), .C2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A(
        n17375), .B(n17374), .ZN(n17376) );
  NAND3_X1 U19335 ( .A1(n17378), .A2(n17377), .A3(n17376), .ZN(n17436) );
  NAND2_X1 U19336 ( .A1(n17440), .A2(n17436), .ZN(n17435) );
  NOR2_X1 U19337 ( .A1(n17431), .A2(n17435), .ZN(n17430) );
  AOI22_X1 U19338 ( .A1(n17505), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n10966), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n17389) );
  AOI22_X1 U19339 ( .A1(n10958), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n10967), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n17388) );
  AOI22_X1 U19340 ( .A1(n10975), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17537), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n17379) );
  OAI21_X1 U19341 ( .B1(n17391), .B2(n17380), .A(n17379), .ZN(n17386) );
  AOI22_X1 U19342 ( .A1(n17545), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17538), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n17384) );
  AOI22_X1 U19343 ( .A1(n14603), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17539), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n17383) );
  AOI22_X1 U19344 ( .A1(n10968), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n20216), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n17382) );
  AOI22_X1 U19345 ( .A1(n17540), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n14589), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n17381) );
  NAND4_X1 U19346 ( .A1(n17384), .A2(n17383), .A3(n17382), .A4(n17381), .ZN(
        n17385) );
  AOI211_X1 U19347 ( .C1(n17547), .C2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A(
        n17386), .B(n17385), .ZN(n17387) );
  NAND3_X1 U19348 ( .A1(n17389), .A2(n17388), .A3(n17387), .ZN(n17417) );
  NAND2_X1 U19349 ( .A1(n17430), .A2(n17417), .ZN(n17424) );
  NOR2_X1 U19350 ( .A1(n17425), .A2(n17424), .ZN(n17423) );
  AOI22_X1 U19351 ( .A1(n17547), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n10967), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n17400) );
  AOI22_X1 U19352 ( .A1(n17505), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17537), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n17399) );
  AOI22_X1 U19353 ( .A1(n10971), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n10975), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n17390) );
  OAI21_X1 U19354 ( .B1(n17391), .B2(n17453), .A(n17390), .ZN(n17397) );
  AOI22_X1 U19355 ( .A1(n17545), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17548), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n17395) );
  AOI22_X1 U19356 ( .A1(n10972), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17539), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n17394) );
  AOI22_X1 U19357 ( .A1(n14589), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n20216), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n17393) );
  AOI22_X1 U19358 ( .A1(n10968), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17540), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n17392) );
  NAND4_X1 U19359 ( .A1(n17395), .A2(n17394), .A3(n17393), .A4(n17392), .ZN(
        n17396) );
  AOI211_X1 U19360 ( .C1(n10959), .C2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A(
        n17397), .B(n17396), .ZN(n17398) );
  NAND3_X1 U19361 ( .A1(n17400), .A2(n17399), .A3(n17398), .ZN(n17420) );
  NAND2_X1 U19362 ( .A1(n17423), .A2(n17420), .ZN(n17419) );
  XNOR2_X1 U19363 ( .A(n17401), .B(n17419), .ZN(n20730) );
  OAI22_X1 U19364 ( .A1(n17403), .A2(n17402), .B1(n20730), .B2(n17522), .ZN(
        P3_U2673) );
  AOI22_X1 U19365 ( .A1(n17547), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n17539), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n17407) );
  AOI22_X1 U19366 ( .A1(n17546), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17548), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n17406) );
  AOI22_X1 U19367 ( .A1(n17540), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n14589), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n17405) );
  AOI22_X1 U19368 ( .A1(n10968), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n20216), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n17404) );
  NAND4_X1 U19369 ( .A1(n17407), .A2(n17406), .A3(n17405), .A4(n17404), .ZN(
        n17413) );
  AOI22_X1 U19370 ( .A1(n10967), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n10971), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n17411) );
  AOI22_X1 U19371 ( .A1(n17505), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10972), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n17410) );
  AOI22_X1 U19372 ( .A1(n17545), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17537), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n17409) );
  AOI22_X1 U19373 ( .A1(n10959), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10975), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n17408) );
  NAND4_X1 U19374 ( .A1(n17411), .A2(n17410), .A3(n17409), .A4(n17408), .ZN(
        n17412) );
  NOR2_X1 U19375 ( .A1(n17413), .A2(n17412), .ZN(n20675) );
  NOR2_X1 U19376 ( .A1(n17526), .A2(n17414), .ZN(n17476) );
  INV_X1 U19377 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n20454) );
  AOI22_X1 U19378 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n17476), .B1(n17445), 
        .B2(n20454), .ZN(n17416) );
  OAI21_X1 U19379 ( .B1(n20675), .B2(n17522), .A(n17416), .ZN(P3_U2682) );
  OAI21_X1 U19380 ( .B1(n17430), .B2(n17417), .A(n17424), .ZN(n20746) );
  INV_X1 U19381 ( .A(P3_EBX_REG_24__SCAN_IN), .ZN(n20488) );
  NAND4_X1 U19382 ( .A1(P3_EBX_REG_23__SCAN_IN), .A2(P3_EBX_REG_22__SCAN_IN), 
        .A3(P3_EBX_REG_21__SCAN_IN), .A4(n17445), .ZN(n17439) );
  NAND2_X1 U19383 ( .A1(P3_EBX_REG_25__SCAN_IN), .A2(n17444), .ZN(n17429) );
  NAND2_X1 U19384 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(n17434), .ZN(n17428) );
  OAI211_X1 U19385 ( .C1(n17434), .C2(P3_EBX_REG_27__SCAN_IN), .A(n17522), .B(
        n17428), .ZN(n17418) );
  OAI21_X1 U19386 ( .B1(n17522), .B2(n20746), .A(n17418), .ZN(P3_U2676) );
  NAND3_X1 U19387 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(P3_EBX_REG_27__SCAN_IN), 
        .A3(n17434), .ZN(n17422) );
  OAI21_X1 U19388 ( .B1(n17423), .B2(n17420), .A(n17419), .ZN(n20734) );
  NAND3_X1 U19389 ( .A1(n17422), .A2(P3_EBX_REG_29__SCAN_IN), .A3(n17522), 
        .ZN(n17421) );
  OAI221_X1 U19390 ( .B1(n17422), .B2(P3_EBX_REG_29__SCAN_IN), .C1(n17522), 
        .C2(n20734), .A(n17421), .ZN(P3_U2674) );
  INV_X1 U19391 ( .A(P3_EBX_REG_28__SCAN_IN), .ZN(n20543) );
  NAND2_X1 U19392 ( .A1(n17522), .A2(n17422), .ZN(n17427) );
  AOI21_X1 U19393 ( .B1(n17425), .B2(n17424), .A(n17423), .ZN(n20735) );
  NAND2_X1 U19394 ( .A1(n20735), .A2(n17526), .ZN(n17426) );
  OAI221_X1 U19395 ( .B1(P3_EBX_REG_28__SCAN_IN), .B2(n17428), .C1(n20543), 
        .C2(n17427), .A(n17426), .ZN(P3_U2675) );
  INV_X1 U19396 ( .A(n17429), .ZN(n17438) );
  AOI21_X1 U19397 ( .B1(P3_EBX_REG_26__SCAN_IN), .B2(n17522), .A(n17438), .ZN(
        n17433) );
  AOI21_X1 U19398 ( .B1(n17431), .B2(n17435), .A(n17430), .ZN(n17432) );
  INV_X1 U19399 ( .A(n17432), .ZN(n20716) );
  OAI22_X1 U19400 ( .A1(n17434), .A2(n17433), .B1(n20716), .B2(n17522), .ZN(
        P3_U2677) );
  AOI21_X1 U19401 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n17522), .A(n17444), .ZN(
        n17437) );
  OAI21_X1 U19402 ( .B1(n17440), .B2(n17436), .A(n17435), .ZN(n20715) );
  OAI22_X1 U19403 ( .A1(n17438), .A2(n17437), .B1(n20715), .B2(n17522), .ZN(
        P3_U2678) );
  INV_X1 U19404 ( .A(n17439), .ZN(n17451) );
  AOI21_X1 U19405 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n17522), .A(n17451), .ZN(
        n17443) );
  AOI21_X1 U19406 ( .B1(n17441), .B2(n17447), .A(n17440), .ZN(n20747) );
  INV_X1 U19407 ( .A(n20747), .ZN(n17442) );
  OAI22_X1 U19408 ( .A1(n17444), .A2(n17443), .B1(n17442), .B2(n17522), .ZN(
        P3_U2679) );
  INV_X1 U19409 ( .A(P3_EBX_REG_22__SCAN_IN), .ZN(n20466) );
  NAND2_X1 U19410 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n17445), .ZN(n17465) );
  NOR2_X1 U19411 ( .A1(n20466), .A2(n17465), .ZN(n17446) );
  AOI21_X1 U19412 ( .B1(P3_EBX_REG_23__SCAN_IN), .B2(n17522), .A(n17446), .ZN(
        n17450) );
  OAI21_X1 U19413 ( .B1(n17449), .B2(n17448), .A(n17447), .ZN(n20757) );
  OAI22_X1 U19414 ( .A1(n17451), .A2(n17450), .B1(n20757), .B2(n17522), .ZN(
        P3_U2680) );
  AOI22_X1 U19415 ( .A1(n10958), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17546), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n17462) );
  AOI22_X1 U19416 ( .A1(n10972), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17537), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n17461) );
  AOI22_X1 U19417 ( .A1(n10966), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n10976), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n17452) );
  OAI21_X1 U19418 ( .B1(n11012), .B2(n17453), .A(n17452), .ZN(n17459) );
  AOI22_X1 U19419 ( .A1(n10961), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17539), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n17457) );
  AOI22_X1 U19420 ( .A1(n17545), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17548), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n17456) );
  AOI22_X1 U19421 ( .A1(n17540), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n14589), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n17455) );
  AOI22_X1 U19422 ( .A1(n10968), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n20216), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n17454) );
  NAND4_X1 U19423 ( .A1(n17457), .A2(n17456), .A3(n17455), .A4(n17454), .ZN(
        n17458) );
  AOI211_X1 U19424 ( .C1(n10967), .C2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A(
        n17459), .B(n17458), .ZN(n17460) );
  NAND3_X1 U19425 ( .A1(n17462), .A2(n17461), .A3(n17460), .ZN(n20685) );
  INV_X1 U19426 ( .A(n20685), .ZN(n17464) );
  NAND3_X1 U19427 ( .A1(n17465), .A2(P3_EBX_REG_22__SCAN_IN), .A3(n17522), 
        .ZN(n17463) );
  OAI221_X1 U19428 ( .B1(n17465), .B2(P3_EBX_REG_22__SCAN_IN), .C1(n17522), 
        .C2(n17464), .A(n17463), .ZN(P3_U2681) );
  AOI22_X1 U19429 ( .A1(n10961), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17546), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n17469) );
  AOI22_X1 U19430 ( .A1(n10958), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n10967), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n17468) );
  AOI22_X1 U19431 ( .A1(n10968), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n20216), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n17467) );
  AOI22_X1 U19432 ( .A1(n17540), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n14589), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n17466) );
  NAND4_X1 U19433 ( .A1(n17469), .A2(n17468), .A3(n17467), .A4(n17466), .ZN(
        n17475) );
  AOI22_X1 U19434 ( .A1(n10971), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n10975), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n17473) );
  AOI22_X1 U19435 ( .A1(n14603), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17537), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n17472) );
  AOI22_X1 U19436 ( .A1(n17547), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n17545), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n17471) );
  AOI22_X1 U19437 ( .A1(n17538), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17539), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n17470) );
  NAND4_X1 U19438 ( .A1(n17473), .A2(n17472), .A3(n17471), .A4(n17470), .ZN(
        n17474) );
  NOR2_X1 U19439 ( .A1(n17475), .A2(n17474), .ZN(n20681) );
  NOR2_X1 U19440 ( .A1(n20711), .A2(n17488), .ZN(n17502) );
  OAI221_X1 U19441 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(P3_EBX_REG_19__SCAN_IN), 
        .C1(P3_EBX_REG_20__SCAN_IN), .C2(n17502), .A(n17476), .ZN(n17477) );
  OAI21_X1 U19442 ( .B1(n20681), .B2(n17522), .A(n17477), .ZN(P3_U2683) );
  AOI22_X1 U19443 ( .A1(n10961), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n14544), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n17481) );
  AOI22_X1 U19444 ( .A1(n10959), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n10967), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n17480) );
  AOI22_X1 U19445 ( .A1(n17540), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n20216), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n17479) );
  AOI22_X1 U19446 ( .A1(n10968), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n14589), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n17478) );
  NAND4_X1 U19447 ( .A1(n17481), .A2(n17480), .A3(n17479), .A4(n17478), .ZN(
        n17487) );
  AOI22_X1 U19448 ( .A1(n17546), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n10971), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n17485) );
  AOI22_X1 U19449 ( .A1(n17545), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17539), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n17484) );
  AOI22_X1 U19450 ( .A1(n17547), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n17548), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n17483) );
  AOI22_X1 U19451 ( .A1(n10972), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n17537), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n17482) );
  NAND4_X1 U19452 ( .A1(n17485), .A2(n17484), .A3(n17483), .A4(n17482), .ZN(
        n17486) );
  NOR2_X1 U19453 ( .A1(n17487), .A2(n17486), .ZN(n20702) );
  AND2_X1 U19454 ( .A1(n17522), .A2(n17488), .ZN(n17503) );
  OAI21_X1 U19455 ( .B1(P3_EBX_REG_18__SCAN_IN), .B2(n17489), .A(n17503), .ZN(
        n17490) );
  OAI21_X1 U19456 ( .B1(n20702), .B2(n17522), .A(n17490), .ZN(P3_U2685) );
  AOI22_X1 U19457 ( .A1(n10958), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17539), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n17494) );
  AOI22_X1 U19458 ( .A1(n17547), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n10966), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n17493) );
  AOI22_X1 U19459 ( .A1(n14589), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n20216), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n17492) );
  AOI22_X1 U19460 ( .A1(n14681), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17540), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n17491) );
  NAND4_X1 U19461 ( .A1(n17494), .A2(n17493), .A3(n17492), .A4(n17491), .ZN(
        n17500) );
  AOI22_X1 U19462 ( .A1(n10961), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17538), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n17498) );
  AOI22_X1 U19463 ( .A1(n10967), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17537), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n17497) );
  AOI22_X1 U19464 ( .A1(n17546), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n10965), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n17496) );
  AOI22_X1 U19465 ( .A1(n17545), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17548), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n17495) );
  NAND4_X1 U19466 ( .A1(n17498), .A2(n17497), .A3(n17496), .A4(n17495), .ZN(
        n17499) );
  NOR2_X1 U19467 ( .A1(n17500), .A2(n17499), .ZN(n20698) );
  AOI22_X1 U19468 ( .A1(P3_EBX_REG_19__SCAN_IN), .A2(n17503), .B1(n17502), 
        .B2(n17501), .ZN(n17504) );
  OAI21_X1 U19469 ( .B1(n20698), .B2(n17522), .A(n17504), .ZN(P3_U2684) );
  AOI22_X1 U19470 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n17505), .B1(
        n17548), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n17509) );
  AOI22_X1 U19471 ( .A1(n10959), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n14544), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n17508) );
  AOI22_X1 U19472 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n10968), .B1(
        P3_INSTQUEUE_REG_10__1__SCAN_IN), .B2(n14589), .ZN(n17507) );
  AOI22_X1 U19473 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n20216), .B1(
        P3_INSTQUEUE_REG_14__1__SCAN_IN), .B2(n17540), .ZN(n17506) );
  NAND4_X1 U19474 ( .A1(n17509), .A2(n17508), .A3(n17507), .A4(n17506), .ZN(
        n17515) );
  AOI22_X1 U19475 ( .A1(n17547), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_12__1__SCAN_IN), .B2(n10967), .ZN(n17513) );
  AOI22_X1 U19476 ( .A1(n17538), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_4__1__SCAN_IN), .B2(n17537), .ZN(n17512) );
  AOI22_X1 U19477 ( .A1(n17545), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n17546), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n17511) );
  AOI22_X1 U19478 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n17539), .B1(
        P3_INSTQUEUE_REG_9__1__SCAN_IN), .B2(n10966), .ZN(n17510) );
  NAND4_X1 U19479 ( .A1(n17513), .A2(n17512), .A3(n17511), .A4(n17510), .ZN(
        n17514) );
  NOR2_X1 U19480 ( .A1(n17515), .A2(n17514), .ZN(n20708) );
  AOI211_X1 U19481 ( .C1(n17518), .C2(n17517), .A(n17516), .B(n17528), .ZN(
        n17519) );
  AOI21_X1 U19482 ( .B1(P3_EBX_REG_17__SCAN_IN), .B2(n17525), .A(n17519), .ZN(
        n17520) );
  OAI21_X1 U19483 ( .B1(n20708), .B2(n17522), .A(n17520), .ZN(P3_U2686) );
  NAND2_X1 U19484 ( .A1(n20179), .A2(n17521), .ZN(n20174) );
  INV_X1 U19485 ( .A(P3_EBX_REG_1__SCAN_IN), .ZN(n20168) );
  OAI222_X1 U19486 ( .A1(n17528), .A2(n20174), .B1(n20168), .B2(n17524), .C1(
        n17523), .C2(n17522), .ZN(P3_U2702) );
  AOI22_X1 U19487 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n17526), .B1(
        P3_EBX_REG_0__SCAN_IN), .B2(n17525), .ZN(n17527) );
  OAI21_X1 U19488 ( .B1(P3_EBX_REG_0__SCAN_IN), .B2(n17528), .A(n17527), .ZN(
        P3_U2703) );
  OAI21_X1 U19489 ( .B1(n21281), .B2(n20112), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n17529) );
  OAI21_X1 U19490 ( .B1(n17530), .B2(n21309), .A(n17529), .ZN(P3_U2634) );
  INV_X1 U19491 ( .A(n17976), .ZN(n17535) );
  OAI21_X1 U19492 ( .B1(P3_FLUSH_REG_SCAN_IN), .B2(n17532), .A(n17531), .ZN(
        n21307) );
  OAI21_X1 U19493 ( .B1(n17533), .B2(n17535), .A(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n17534) );
  OAI221_X1 U19494 ( .B1(n17535), .B2(n21307), .C1(n17535), .C2(n18704), .A(
        n17534), .ZN(P3_U2863) );
  INV_X1 U19495 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n17536) );
  INV_X1 U19496 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n21241) );
  INV_X1 U19497 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n17847) );
  NOR2_X1 U19498 ( .A1(n21241), .A2(n17847), .ZN(n20954) );
  NAND3_X1 U19499 ( .A1(n20954), .A2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n20965) );
  NOR2_X1 U19500 ( .A1(n17536), .A2(n20965), .ZN(n20975) );
  NAND2_X1 U19501 ( .A1(n20975), .A2(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n20977) );
  INV_X1 U19502 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n21172) );
  NOR2_X1 U19503 ( .A1(n20977), .A2(n21172), .ZN(n21168) );
  AOI22_X1 U19504 ( .A1(n17538), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n17537), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n17544) );
  AOI22_X1 U19505 ( .A1(n10971), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n17539), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n17543) );
  AOI22_X1 U19506 ( .A1(n10968), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n14589), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n17542) );
  AOI22_X1 U19507 ( .A1(n17540), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n20216), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n17541) );
  NAND4_X1 U19508 ( .A1(n17544), .A2(n17543), .A3(n17542), .A4(n17541), .ZN(
        n17554) );
  AOI22_X1 U19509 ( .A1(n10959), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n10967), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n17552) );
  AOI22_X1 U19510 ( .A1(n17545), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n10976), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n17551) );
  AOI22_X1 U19511 ( .A1(n17547), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n17546), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n17550) );
  AOI22_X1 U19512 ( .A1(n10961), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n17548), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n17549) );
  NAND4_X1 U19513 ( .A1(n17552), .A2(n17551), .A3(n17550), .A4(n17549), .ZN(
        n17553) );
  NAND2_X1 U19514 ( .A1(n17555), .A2(n20642), .ZN(n17556) );
  NOR2_X1 U19515 ( .A1(n21106), .A2(n17556), .ZN(n17564) );
  XOR2_X1 U19516 ( .A(n21106), .B(n17556), .Z(n17891) );
  NAND2_X1 U19517 ( .A1(n17558), .A2(n17557), .ZN(n17560) );
  INV_X1 U19518 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n20935) );
  NAND2_X1 U19519 ( .A1(n17564), .A2(n17561), .ZN(n17565) );
  NAND2_X1 U19520 ( .A1(n17891), .A2(n17892), .ZN(n17890) );
  NAND2_X1 U19521 ( .A1(n17564), .A2(n17563), .ZN(n17562) );
  OAI211_X1 U19522 ( .C1(n17564), .C2(n17563), .A(n17890), .B(n17562), .ZN(
        n17878) );
  NAND2_X1 U19523 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n17878), .ZN(
        n17877) );
  NAND2_X1 U19524 ( .A1(n17565), .A2(n17877), .ZN(n17576) );
  AOI21_X1 U19525 ( .B1(n21106), .B2(n17568), .A(n17774), .ZN(n17572) );
  NAND2_X1 U19526 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n17569), .ZN(
        n17571) );
  NAND2_X1 U19527 ( .A1(n17572), .A2(n17600), .ZN(n17573) );
  NAND2_X1 U19528 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n17895), .ZN(
        n17894) );
  INV_X1 U19529 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n21232) );
  NOR2_X2 U19530 ( .A1(n17602), .A2(n21232), .ZN(n20950) );
  NAND2_X1 U19531 ( .A1(n21106), .A2(n17577), .ZN(n17829) );
  NAND2_X1 U19532 ( .A1(n21168), .A2(n17872), .ZN(n17820) );
  INV_X1 U19533 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n21198) );
  INV_X1 U19534 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n21191) );
  NOR2_X1 U19535 ( .A1(n21198), .A2(n21191), .ZN(n21170) );
  INV_X1 U19536 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n21183) );
  NAND2_X1 U19537 ( .A1(n21170), .A2(n21183), .ZN(n21189) );
  NAND2_X1 U19538 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n17635) );
  NAND2_X1 U19539 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n17612) );
  INV_X1 U19540 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n20186) );
  NOR2_X1 U19541 ( .A1(n17574), .A2(n20186), .ZN(n17808) );
  AOI21_X1 U19542 ( .B1(n17924), .B2(n17574), .A(n17954), .ZN(n17811) );
  OAI21_X1 U19543 ( .B1(n17808), .B2(n17967), .A(n17811), .ZN(n17592) );
  INV_X1 U19544 ( .A(n19010), .ZN(n18968) );
  INV_X1 U19545 ( .A(n17768), .ZN(n17686) );
  NOR3_X1 U19546 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n17686), .A3(
        n17574), .ZN(n17593) );
  INV_X1 U19547 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n20413) );
  NAND2_X1 U19548 ( .A1(n17588), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n17587) );
  OAI21_X1 U19549 ( .B1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n17808), .A(
        n17587), .ZN(n20409) );
  NAND2_X1 U19550 ( .A1(n21238), .A2(P3_REIP_REG_18__SCAN_IN), .ZN(n21187) );
  OAI21_X1 U19551 ( .B1(n17809), .B2(n20409), .A(n21187), .ZN(n17575) );
  AOI211_X1 U19552 ( .C1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(n17592), .A(
        n17593), .B(n17575), .ZN(n17586) );
  INV_X1 U19553 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n20974) );
  NAND2_X1 U19554 ( .A1(n20975), .A2(n17576), .ZN(n17825) );
  AOI22_X1 U19555 ( .A1(n17885), .A2(n20990), .B1(n17840), .B2(n21174), .ZN(
        n17618) );
  OAI21_X1 U19556 ( .B1(n21170), .B2(n17820), .A(n17618), .ZN(n17817) );
  NAND2_X1 U19557 ( .A1(n21115), .A2(n21183), .ZN(n17644) );
  INV_X1 U19558 ( .A(n17644), .ZN(n17678) );
  AOI21_X1 U19559 ( .B1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n17774), .A(
        n17678), .ZN(n17584) );
  NAND2_X1 U19560 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n21115), .ZN(
        n17578) );
  AOI22_X1 U19561 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n21115), .B1(
        n17774), .B2(n21232), .ZN(n17884) );
  NAND2_X1 U19562 ( .A1(n21168), .A2(n17849), .ZN(n17581) );
  NAND2_X1 U19563 ( .A1(n21241), .A2(n17847), .ZN(n17859) );
  NOR4_X1 U19564 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A4(n17859), .ZN(n17580) );
  AOI21_X1 U19565 ( .B1(n17580), .B2(n17579), .A(n17774), .ZN(n17583) );
  INV_X1 U19566 ( .A(n21170), .ZN(n21175) );
  INV_X1 U19567 ( .A(n17581), .ZN(n17582) );
  NOR2_X1 U19568 ( .A1(n17583), .A2(n17582), .ZN(n17708) );
  OR2_X1 U19569 ( .A1(n21175), .A2(n17708), .ZN(n17594) );
  NAND2_X1 U19570 ( .A1(n17710), .A2(n17594), .ZN(n17645) );
  XNOR2_X1 U19571 ( .A(n17584), .B(n17645), .ZN(n21186) );
  AOI22_X1 U19572 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17817), .B1(
        n17886), .B2(n21186), .ZN(n17585) );
  OAI211_X1 U19573 ( .C1(n17820), .C2(n21189), .A(n17586), .B(n17585), .ZN(
        P3_U2812) );
  INV_X1 U19574 ( .A(n21168), .ZN(n20847) );
  NAND2_X1 U19575 ( .A1(n21170), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n17654) );
  NOR2_X1 U19576 ( .A1(n20847), .A2(n17654), .ZN(n20849) );
  NAND2_X1 U19577 ( .A1(n20849), .A2(n10978), .ZN(n17683) );
  INV_X1 U19578 ( .A(n17587), .ZN(n20424) );
  NAND2_X1 U19579 ( .A1(n17672), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n20423) );
  OAI21_X1 U19580 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n20424), .A(
        n20423), .ZN(n20428) );
  NAND2_X1 U19581 ( .A1(n21238), .A2(P3_REIP_REG_19__SCAN_IN), .ZN(n17590) );
  NAND3_X1 U19582 ( .A1(n17588), .A2(n11228), .A3(n17768), .ZN(n17589) );
  OAI211_X1 U19583 ( .C1(n17809), .C2(n20428), .A(n17590), .B(n17589), .ZN(
        n17591) );
  AOI221_X1 U19584 ( .B1(n17593), .B2(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .C1(
        n17592), .C2(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(n17591), .ZN(
        n17597) );
  INV_X1 U19585 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n21158) );
  NOR3_X1 U19586 ( .A1(n17654), .A2(n21158), .A3(n20990), .ZN(n21150) );
  NOR3_X1 U19587 ( .A1(n17654), .A2(n21158), .A3(n21174), .ZN(n21148) );
  OAI22_X1 U19588 ( .A1(n21150), .A2(n17829), .B1(n21148), .B2(n17971), .ZN(
        n17680) );
  NOR2_X1 U19589 ( .A1(n17644), .A2(n17645), .ZN(n17663) );
  NOR3_X1 U19590 ( .A1(n21115), .A2(n21183), .A3(n17594), .ZN(n17677) );
  NOR2_X1 U19591 ( .A1(n17663), .A2(n17677), .ZN(n17595) );
  XNOR2_X1 U19592 ( .A(n17595), .B(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n21156) );
  AOI22_X1 U19593 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17680), .B1(
        n17886), .B2(n21156), .ZN(n17596) );
  OAI211_X1 U19594 ( .C1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n17683), .A(
        n17597), .B(n17596), .ZN(P3_U2811) );
  NAND2_X1 U19595 ( .A1(n17885), .A2(n20990), .ZN(n17608) );
  NOR2_X1 U19596 ( .A1(n17686), .A2(n17598), .ZN(n17613) );
  INV_X1 U19597 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n20370) );
  NOR2_X1 U19598 ( .A1(n17598), .A2(n20186), .ZN(n17822) );
  AOI21_X1 U19599 ( .B1(n17924), .B2(n17598), .A(n17954), .ZN(n17833) );
  OAI21_X1 U19600 ( .B1(n17822), .B2(n17967), .A(n17833), .ZN(n17611) );
  NAND2_X1 U19601 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n17822), .ZN(
        n17610) );
  OAI21_X1 U19602 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n17822), .A(
        n17610), .ZN(n20368) );
  NAND2_X1 U19603 ( .A1(n21238), .A2(P3_REIP_REG_15__SCAN_IN), .ZN(n21002) );
  OAI21_X1 U19604 ( .B1(n17809), .B2(n20368), .A(n21002), .ZN(n17599) );
  AOI221_X1 U19605 ( .B1(n17613), .B2(n20370), .C1(n17611), .C2(
        P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A(n17599), .ZN(n17607) );
  NAND2_X1 U19606 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n20946) );
  INV_X1 U19607 ( .A(n20946), .ZN(n17601) );
  NAND3_X1 U19608 ( .A1(n17774), .A2(n17601), .A3(n17600), .ZN(n17863) );
  NAND2_X1 U19609 ( .A1(n17602), .A2(n21232), .ZN(n17864) );
  NOR2_X1 U19610 ( .A1(n17859), .A2(n17864), .ZN(n17838) );
  INV_X1 U19611 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n21209) );
  NAND2_X1 U19612 ( .A1(n17838), .A2(n21209), .ZN(n17631) );
  NOR3_X1 U19613 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A3(n17631), .ZN(n17826) );
  NAND2_X1 U19614 ( .A1(n17826), .A2(n20974), .ZN(n17603) );
  OAI21_X1 U19615 ( .B1(n17863), .B2(n20977), .A(n17603), .ZN(n17604) );
  XNOR2_X1 U19616 ( .A(n17604), .B(n21172), .ZN(n21001) );
  NAND2_X1 U19617 ( .A1(n17824), .A2(n21172), .ZN(n21004) );
  OAI22_X1 U19618 ( .A1(n17618), .A2(n21172), .B1(n17971), .B2(n21004), .ZN(
        n17605) );
  AOI21_X1 U19619 ( .B1(n17886), .B2(n21001), .A(n17605), .ZN(n17606) );
  OAI211_X1 U19620 ( .C1(n20994), .C2(n17608), .A(n17607), .B(n17606), .ZN(
        P3_U2815) );
  AOI22_X1 U19621 ( .A1(n17774), .A2(n21198), .B1(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n21115), .ZN(n17609) );
  XNOR2_X1 U19622 ( .A(n17708), .B(n17609), .ZN(n21204) );
  INV_X1 U19623 ( .A(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n20383) );
  AND2_X1 U19624 ( .A1(n17810), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n20392) );
  AOI21_X1 U19625 ( .B1(n20383), .B2(n17610), .A(n20392), .ZN(n20378) );
  AOI22_X1 U19626 ( .A1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n17611), .B1(
        n10962), .B2(n20378), .ZN(n17615) );
  NAND2_X1 U19627 ( .A1(n21238), .A2(P3_REIP_REG_16__SCAN_IN), .ZN(n21205) );
  OAI211_X1 U19628 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(n17613), .B(n17612), .ZN(n17614) );
  NAND3_X1 U19629 ( .A1(n17615), .A2(n21205), .A3(n17614), .ZN(n17616) );
  AOI21_X1 U19630 ( .B1(n17886), .B2(n21204), .A(n17616), .ZN(n17617) );
  OAI221_X1 U19631 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n17820), 
        .C1(n21198), .C2(n17618), .A(n17617), .ZN(P3_U2814) );
  INV_X1 U19632 ( .A(n17630), .ZN(n17620) );
  NAND2_X1 U19633 ( .A1(n20954), .A2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n20967) );
  INV_X1 U19634 ( .A(n20967), .ZN(n17619) );
  NAND3_X1 U19635 ( .A1(n17774), .A2(n17620), .A3(n17619), .ZN(n17621) );
  NAND2_X1 U19636 ( .A1(n17631), .A2(n17621), .ZN(n17622) );
  XNOR2_X1 U19637 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B(n17622), .ZN(
        n20973) );
  NOR2_X1 U19638 ( .A1(n17686), .A2(n17623), .ZN(n17636) );
  INV_X1 U19639 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n20325) );
  NOR2_X1 U19640 ( .A1(n17623), .A2(n20186), .ZN(n17835) );
  AOI21_X1 U19641 ( .B1(n17924), .B2(n17623), .A(n17954), .ZN(n17624) );
  OAI21_X1 U19642 ( .B1(n17835), .B2(n17967), .A(n17624), .ZN(n17640) );
  INV_X1 U19643 ( .A(n17835), .ZN(n17633) );
  AOI22_X1 U19644 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n17633), .B1(
        n17835), .B2(n20325), .ZN(n20322) );
  NAND2_X1 U19645 ( .A1(n21238), .A2(P3_REIP_REG_12__SCAN_IN), .ZN(n20971) );
  OAI21_X1 U19646 ( .B1(n17809), .B2(n20322), .A(n20971), .ZN(n17625) );
  AOI221_X1 U19647 ( .B1(n17636), .B2(n20325), .C1(n17640), .C2(
        P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A(n17625), .ZN(n17628) );
  NOR2_X1 U19648 ( .A1(n21176), .A2(n20965), .ZN(n17629) );
  NOR2_X1 U19649 ( .A1(n20952), .A2(n20965), .ZN(n20961) );
  OAI22_X1 U19650 ( .A1(n17629), .A2(n17829), .B1(n20961), .B2(n17971), .ZN(
        n17641) );
  NOR2_X1 U19651 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n20967), .ZN(
        n17626) );
  AOI22_X1 U19652 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n17641), .B1(
        n17626), .B2(n10978), .ZN(n17627) );
  OAI211_X1 U19653 ( .C1(n20973), .C2(n17876), .A(n17628), .B(n17627), .ZN(
        P3_U2818) );
  INV_X1 U19654 ( .A(n17629), .ZN(n20964) );
  OAI22_X1 U19655 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n17631), .B1(
        n20964), .B2(n17630), .ZN(n17632) );
  XNOR2_X1 U19656 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B(n17632), .ZN(
        n21216) );
  NOR2_X1 U19657 ( .A1(n20325), .A2(n17633), .ZN(n17634) );
  NAND2_X1 U19658 ( .A1(n17821), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n17823) );
  OAI21_X1 U19659 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n17634), .A(
        n17823), .ZN(n20350) );
  OAI211_X1 U19660 ( .C1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A(n17636), .B(n17635), .ZN(n17638) );
  NAND2_X1 U19661 ( .A1(n21238), .A2(P3_REIP_REG_13__SCAN_IN), .ZN(n17637) );
  OAI211_X1 U19662 ( .C1(n17809), .C2(n20350), .A(n17638), .B(n17637), .ZN(
        n17639) );
  AOI21_X1 U19663 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n17640), .A(
        n17639), .ZN(n17643) );
  NOR2_X1 U19664 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n20965), .ZN(
        n21208) );
  AOI22_X1 U19665 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n17641), .B1(
        n21208), .B2(n10978), .ZN(n17642) );
  OAI211_X1 U19666 ( .C1(n21216), .C2(n17876), .A(n17643), .B(n17642), .ZN(
        P3_U2817) );
  INV_X1 U19667 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n21010) );
  NOR4_X1 U19668 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A4(n17644), .ZN(n17689) );
  INV_X1 U19669 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n17669) );
  NOR2_X1 U19670 ( .A1(n17669), .A2(n21158), .ZN(n20861) );
  AND2_X1 U19671 ( .A1(n20861), .A2(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n21031) );
  NAND3_X1 U19672 ( .A1(n21031), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        n17645), .ZN(n17711) );
  INV_X1 U19673 ( .A(n17711), .ZN(n17646) );
  OAI21_X1 U19674 ( .B1(n17689), .B2(n17646), .A(n17710), .ZN(n17690) );
  XNOR2_X1 U19675 ( .A(n21010), .B(n17690), .ZN(n21014) );
  INV_X1 U19676 ( .A(n20423), .ZN(n17671) );
  OAI22_X1 U19677 ( .A1(n17671), .A2(n17967), .B1(n17649), .B2(n17879), .ZN(
        n17647) );
  NOR2_X1 U19678 ( .A1(n17954), .A2(n17647), .ZN(n17674) );
  OAI21_X1 U19679 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n17760), .A(
        n17674), .ZN(n17662) );
  INV_X1 U19680 ( .A(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n17648) );
  INV_X1 U19681 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n17659) );
  NAND2_X1 U19682 ( .A1(n17649), .A2(n17768), .ZN(n17660) );
  AOI221_X1 U19683 ( .B1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .C1(n17648), .C2(n17659), .A(
        n17660), .ZN(n17653) );
  INV_X1 U19684 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n20473) );
  NAND2_X1 U19685 ( .A1(n17649), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n17670) );
  NOR2_X1 U19686 ( .A1(n17659), .A2(n17670), .ZN(n17651) );
  NOR2_X1 U19687 ( .A1(n11038), .A2(n20186), .ZN(n17688) );
  INV_X1 U19688 ( .A(n17688), .ZN(n17650) );
  OAI21_X1 U19689 ( .B1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n17651), .A(
        n17650), .ZN(n20462) );
  OAI22_X1 U19690 ( .A1(n21223), .A2(n20473), .B1(n20462), .B2(n17809), .ZN(
        n17652) );
  AOI211_X1 U19691 ( .C1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .C2(n17662), .A(
        n17653), .B(n17652), .ZN(n17657) );
  INV_X1 U19692 ( .A(n17654), .ZN(n20848) );
  NAND2_X1 U19693 ( .A1(n20848), .A2(n21031), .ZN(n17706) );
  OAI22_X1 U19694 ( .A1(n20856), .A2(n17829), .B1(n20858), .B2(n17971), .ZN(
        n17666) );
  OAI21_X1 U19695 ( .B1(n17706), .B2(n17820), .A(n21010), .ZN(n17655) );
  OAI21_X1 U19696 ( .B1(n21010), .B2(n17666), .A(n17655), .ZN(n17656) );
  OAI211_X1 U19697 ( .C1(n17876), .C2(n21014), .A(n17657), .B(n17656), .ZN(
        P3_U2808) );
  INV_X1 U19698 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n17658) );
  NAND2_X1 U19699 ( .A1(n20861), .A2(n17658), .ZN(n20865) );
  INV_X1 U19700 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n20458) );
  NOR2_X1 U19701 ( .A1(n21223), .A2(n20458), .ZN(n20853) );
  XNOR2_X1 U19702 ( .A(n17659), .B(n17670), .ZN(n20452) );
  OAI22_X1 U19703 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n17660), .B1(
        n17809), .B2(n20452), .ZN(n17661) );
  AOI211_X1 U19704 ( .C1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .C2(n17662), .A(
        n20853), .B(n17661), .ZN(n17668) );
  NOR2_X1 U19705 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n17664) );
  AOI22_X1 U19706 ( .A1(n20861), .A2(n17677), .B1(n17664), .B2(n17663), .ZN(
        n17665) );
  XNOR2_X1 U19707 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .B(n17665), .ZN(
        n20854) );
  AOI22_X1 U19708 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17666), .B1(
        n17886), .B2(n20854), .ZN(n17667) );
  OAI211_X1 U19709 ( .C1(n20865), .C2(n17683), .A(n17668), .B(n17667), .ZN(
        P3_U2809) );
  NAND2_X1 U19710 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17669), .ZN(
        n21167) );
  OAI21_X1 U19711 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n17671), .A(
        n17670), .ZN(n20435) );
  INV_X1 U19712 ( .A(n20435), .ZN(n17676) );
  AOI21_X1 U19713 ( .B1(n17672), .B2(n18884), .A(
        P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n17673) );
  NAND2_X1 U19714 ( .A1(n21238), .A2(P3_REIP_REG_20__SCAN_IN), .ZN(n21165) );
  OAI21_X1 U19715 ( .B1(n17674), .B2(n17673), .A(n21165), .ZN(n17675) );
  AOI221_X1 U19716 ( .B1(n10962), .B2(n17676), .C1(n17759), .C2(n17676), .A(
        n17675), .ZN(n17682) );
  OAI221_X1 U19717 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n17678), 
        .C1(n21158), .C2(n17677), .A(n17710), .ZN(n17679) );
  XNOR2_X1 U19718 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .B(n17679), .ZN(
        n21162) );
  AOI22_X1 U19719 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n17680), .B1(
        n17886), .B2(n21162), .ZN(n17681) );
  OAI211_X1 U19720 ( .C1(n17683), .C2(n21167), .A(n17682), .B(n17681), .ZN(
        P3_U2810) );
  INV_X1 U19721 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n21131) );
  NOR2_X1 U19722 ( .A1(n21010), .A2(n21131), .ZN(n21030) );
  AND2_X1 U19723 ( .A1(n21125), .A2(n17840), .ZN(n17685) );
  NAND2_X1 U19724 ( .A1(n21030), .A2(n20856), .ZN(n21126) );
  AND2_X1 U19725 ( .A1(n21126), .A2(n17885), .ZN(n17684) );
  AOI22_X1 U19726 ( .A1(n20858), .A2(n17685), .B1(n20856), .B2(n17684), .ZN(
        n17697) );
  INV_X1 U19727 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n18066) );
  NOR2_X1 U19728 ( .A1(n21223), .A2(n18066), .ZN(n17695) );
  NOR3_X1 U19729 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n17686), .A3(
        n11038), .ZN(n17694) );
  INV_X1 U19730 ( .A(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n20485) );
  OAI22_X1 U19731 ( .A1(n17688), .A2(n17967), .B1(n17701), .B2(n19009), .ZN(
        n17687) );
  NOR2_X1 U19732 ( .A1(n17954), .A2(n17687), .ZN(n17698) );
  NAND2_X1 U19733 ( .A1(n17701), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n17716) );
  OAI21_X1 U19734 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n17688), .A(
        n17716), .ZN(n20482) );
  OAI22_X1 U19735 ( .A1(n17698), .A2(n20485), .B1(n20482), .B2(n17809), .ZN(
        n17693) );
  AOI22_X1 U19736 ( .A1(n17885), .A2(n21126), .B1(n17840), .B2(n21125), .ZN(
        n17727) );
  NAND2_X1 U19737 ( .A1(n17689), .A2(n21010), .ZN(n17707) );
  AOI221_X1 U19738 ( .B1(n21115), .B2(n17707), .C1(n21010), .C2(n17707), .A(
        n17690), .ZN(n17691) );
  XNOR2_X1 U19739 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B(n17691), .ZN(
        n21136) );
  OAI22_X1 U19740 ( .A1(n17727), .A2(n21131), .B1(n17876), .B2(n21136), .ZN(
        n17692) );
  NOR4_X1 U19741 ( .A1(n17695), .A2(n17694), .A3(n17693), .A4(n17692), .ZN(
        n17696) );
  OAI21_X1 U19742 ( .B1(n17697), .B2(n21010), .A(n17696), .ZN(P3_U2807) );
  INV_X1 U19743 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n21032) );
  XNOR2_X1 U19744 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B(n17735), .ZN(
        n21017) );
  OAI21_X1 U19745 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n17967), .A(
        n17698), .ZN(n17720) );
  INV_X1 U19746 ( .A(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n17699) );
  INV_X1 U19747 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n17700) );
  NAND2_X1 U19748 ( .A1(n17701), .A2(n17768), .ZN(n17717) );
  AOI221_X1 U19749 ( .B1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .C1(n17699), .C2(n17700), .A(
        n17717), .ZN(n17705) );
  INV_X1 U19750 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n20506) );
  NOR2_X1 U19751 ( .A1(n17700), .A2(n17716), .ZN(n17703) );
  NOR2_X1 U19752 ( .A1(n17756), .A2(n20186), .ZN(n17758) );
  INV_X1 U19753 ( .A(n17758), .ZN(n17702) );
  OAI21_X1 U19754 ( .B1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n17703), .A(
        n17702), .ZN(n20503) );
  OAI22_X1 U19755 ( .A1(n21223), .A2(n20506), .B1(n20503), .B2(n17809), .ZN(
        n17704) );
  AOI211_X1 U19756 ( .C1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .C2(n17720), .A(
        n17705), .B(n17704), .ZN(n17715) );
  NOR2_X1 U19757 ( .A1(n21032), .A2(n21126), .ZN(n17734) );
  INV_X1 U19758 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n21033) );
  XNOR2_X1 U19759 ( .A(n17734), .B(n21033), .ZN(n21020) );
  INV_X1 U19760 ( .A(n21030), .ZN(n17712) );
  OR2_X1 U19761 ( .A1(n17712), .A2(n17706), .ZN(n17723) );
  OAI22_X1 U19762 ( .A1(n17708), .A2(n17723), .B1(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n17707), .ZN(n17709) );
  AOI21_X1 U19763 ( .B1(n17774), .B2(n10986), .A(n17753), .ZN(n17713) );
  XNOR2_X1 U19764 ( .A(n17713), .B(n21033), .ZN(n21021) );
  AOI22_X1 U19765 ( .A1(n17885), .A2(n21020), .B1(n17886), .B2(n21021), .ZN(
        n17714) );
  OAI211_X1 U19766 ( .C1(n17971), .C2(n21017), .A(n17715), .B(n17714), .ZN(
        P3_U2805) );
  INV_X1 U19767 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n20505) );
  NOR2_X1 U19768 ( .A1(n21223), .A2(n20505), .ZN(n17719) );
  XOR2_X1 U19769 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .B(n17716), .Z(
        n20493) );
  OAI22_X1 U19770 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n17717), .B1(
        n17809), .B2(n20493), .ZN(n17718) );
  AOI211_X1 U19771 ( .C1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .C2(n17720), .A(
        n17719), .B(n17718), .ZN(n17726) );
  AOI21_X1 U19772 ( .B1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n17722), .A(
        n17721), .ZN(n21144) );
  INV_X1 U19773 ( .A(n21144), .ZN(n17724) );
  NOR2_X1 U19774 ( .A1(n17723), .A2(n17820), .ZN(n17736) );
  AOI22_X1 U19775 ( .A1(n17886), .A2(n17724), .B1(n17736), .B2(n21032), .ZN(
        n17725) );
  OAI211_X1 U19776 ( .C1(n17727), .C2(n21032), .A(n17726), .B(n17725), .ZN(
        P3_U2806) );
  INV_X1 U19777 ( .A(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n20520) );
  AND3_X1 U19778 ( .A1(n11222), .A2(n17768), .A3(n11063), .ZN(n17745) );
  OAI22_X1 U19779 ( .A1(n17758), .A2(n17967), .B1(n11063), .B2(n17879), .ZN(
        n17728) );
  NOR2_X1 U19780 ( .A1(n17954), .A2(n17728), .ZN(n17755) );
  OAI21_X1 U19781 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n17760), .A(
        n17755), .ZN(n17748) );
  NOR2_X1 U19782 ( .A1(n17729), .A2(n20186), .ZN(n17744) );
  NOR2_X1 U19783 ( .A1(n17797), .A2(n20186), .ZN(n17801) );
  INV_X1 U19784 ( .A(n17801), .ZN(n17730) );
  OAI21_X1 U19785 ( .B1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n17744), .A(
        n17730), .ZN(n20548) );
  NAND2_X1 U19786 ( .A1(n21238), .A2(P3_REIP_REG_28__SCAN_IN), .ZN(n21120) );
  INV_X1 U19787 ( .A(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n20542) );
  NAND3_X1 U19788 ( .A1(n17731), .A2(n20542), .A3(n17768), .ZN(n17732) );
  OAI211_X1 U19789 ( .C1(n20548), .C2(n17809), .A(n21120), .B(n17732), .ZN(
        n17733) );
  AOI221_X1 U19790 ( .B1(n17745), .B2(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .C1(
        n17748), .C2(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A(n17733), .ZN(
        n17743) );
  INV_X1 U19791 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n17765) );
  NOR2_X1 U19792 ( .A1(n17765), .A2(n21033), .ZN(n21040) );
  NAND2_X1 U19793 ( .A1(n21040), .A2(n17734), .ZN(n21028) );
  NAND2_X1 U19794 ( .A1(n21040), .A2(n17735), .ZN(n17781) );
  AOI22_X1 U19795 ( .A1(n17885), .A2(n21028), .B1(n17840), .B2(n17781), .ZN(
        n17764) );
  NAND2_X1 U19796 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n17764), .ZN(
        n17749) );
  OAI211_X1 U19797 ( .C1(n17840), .C2(n17885), .A(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B(n17749), .ZN(n17742) );
  NAND3_X1 U19798 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(n17736), .ZN(n17766) );
  NOR2_X1 U19799 ( .A1(n17765), .A2(n17766), .ZN(n17780) );
  INV_X1 U19800 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n21069) );
  NAND3_X1 U19801 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n17780), .A3(
        n21069), .ZN(n17741) );
  NOR2_X1 U19802 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17774), .ZN(
        n17793) );
  AOI21_X1 U19803 ( .B1(n17774), .B2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n17793), .ZN(n21118) );
  AOI21_X1 U19804 ( .B1(n17765), .B2(n21033), .A(n17774), .ZN(n17737) );
  INV_X1 U19805 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n21046) );
  NOR2_X1 U19806 ( .A1(n17738), .A2(n21046), .ZN(n17773) );
  NOR2_X1 U19807 ( .A1(n17792), .A2(n17773), .ZN(n17747) );
  NAND2_X1 U19808 ( .A1(n17774), .A2(n17747), .ZN(n17746) );
  NAND2_X1 U19809 ( .A1(n21119), .A2(n17746), .ZN(n17739) );
  NAND2_X1 U19810 ( .A1(n21118), .A2(n17739), .ZN(n21103) );
  OAI211_X1 U19811 ( .C1(n21118), .C2(n17739), .A(n17886), .B(n21103), .ZN(
        n17740) );
  NAND4_X1 U19812 ( .A1(n17743), .A2(n17742), .A3(n17741), .A4(n17740), .ZN(
        P3_U2802) );
  NAND2_X1 U19813 ( .A1(n11063), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n17757) );
  AOI21_X1 U19814 ( .B1(n11222), .B2(n17757), .A(n17744), .ZN(n20533) );
  AOI21_X1 U19815 ( .B1(n10962), .B2(n20533), .A(n17745), .ZN(n17752) );
  OAI21_X1 U19816 ( .B1(n17774), .B2(n17747), .A(n17746), .ZN(n21039) );
  AOI22_X1 U19817 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n17748), .B1(
        n17886), .B2(n21039), .ZN(n17751) );
  OAI21_X1 U19818 ( .B1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n17780), .A(
        n17749), .ZN(n17750) );
  NAND2_X1 U19819 ( .A1(n21238), .A2(P3_REIP_REG_27__SCAN_IN), .ZN(n21054) );
  NAND4_X1 U19820 ( .A1(n17752), .A2(n17751), .A3(n17750), .A4(n21054), .ZN(
        P3_U2803) );
  AOI221_X1 U19821 ( .B1(n17774), .B2(n21033), .C1(n10986), .C2(
        P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A(n17753), .ZN(n17754) );
  XOR2_X1 U19822 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B(n17754), .Z(
        n21025) );
  AOI221_X1 U19823 ( .B1(n17756), .B2(n20520), .C1(n19009), .C2(n20520), .A(
        n17755), .ZN(n17762) );
  OAI21_X1 U19824 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n17758), .A(
        n17757), .ZN(n20525) );
  INV_X1 U19825 ( .A(n17759), .ZN(n17760) );
  NAND2_X1 U19826 ( .A1(n21238), .A2(P3_REIP_REG_26__SCAN_IN), .ZN(n21036) );
  OAI221_X1 U19827 ( .B1(n20525), .B2(n17809), .C1(n20525), .C2(n17760), .A(
        n21036), .ZN(n17761) );
  AOI211_X1 U19828 ( .C1(n21025), .C2(n17886), .A(n17762), .B(n17761), .ZN(
        n17763) );
  OAI221_X1 U19829 ( .B1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n17766), 
        .C1(n17765), .C2(n17764), .A(n17763), .ZN(P3_U2804) );
  NAND2_X1 U19830 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n21057) );
  NOR2_X1 U19831 ( .A1(n21057), .A2(n21028), .ZN(n21107) );
  NAND3_X1 U19832 ( .A1(n21107), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n17767) );
  XOR2_X1 U19833 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n17767), .Z(
        n21096) );
  INV_X1 U19834 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n20559) );
  XOR2_X2 U19835 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .B(n11039), .Z(
        n20391) );
  INV_X1 U19836 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n20594) );
  NOR2_X1 U19837 ( .A1(n21223), .A2(n20594), .ZN(n21099) );
  NAND2_X1 U19838 ( .A1(n17769), .A2(n17768), .ZN(n17787) );
  INV_X1 U19839 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n17770) );
  XOR2_X1 U19840 ( .A(n17770), .B(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .Z(
        n17771) );
  NOR2_X1 U19841 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n17760), .ZN(
        n17803) );
  OR2_X1 U19842 ( .A1(n19009), .A2(n17769), .ZN(n17798) );
  OAI211_X1 U19843 ( .C1(n17801), .C2(n17967), .A(n17798), .B(n10979), .ZN(
        n17795) );
  NOR2_X1 U19844 ( .A1(n17803), .A2(n17795), .ZN(n17786) );
  OAI22_X1 U19845 ( .A1(n17787), .A2(n17771), .B1(n17786), .B2(n17770), .ZN(
        n17772) );
  AOI211_X1 U19846 ( .C1(n20577), .C2(n10962), .A(n21099), .B(n17772), .ZN(
        n17779) );
  INV_X1 U19847 ( .A(n17773), .ZN(n17776) );
  NAND2_X1 U19848 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17774), .ZN(
        n17775) );
  NOR2_X1 U19849 ( .A1(n17776), .A2(n17775), .ZN(n21105) );
  NAND2_X1 U19850 ( .A1(n21105), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n17782) );
  INV_X1 U19851 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n21082) );
  NAND3_X1 U19852 ( .A1(n17793), .A2(n17792), .A3(n21082), .ZN(n17783) );
  INV_X1 U19853 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n21081) );
  AOI22_X1 U19854 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n17782), .B1(
        n17783), .B2(n21081), .ZN(n17777) );
  XOR2_X1 U19855 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n17777), .Z(
        n21097) );
  NAND2_X1 U19856 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n21089) );
  AOI22_X1 U19857 ( .A1(n17886), .A2(n21097), .B1(n17840), .B2(n21092), .ZN(
        n17778) );
  OAI211_X1 U19858 ( .C1(n21096), .C2(n17829), .A(n17779), .B(n17778), .ZN(
        P3_U2799) );
  NOR2_X1 U19859 ( .A1(n21057), .A2(n21082), .ZN(n21078) );
  NAND2_X1 U19860 ( .A1(n21078), .A2(n17780), .ZN(n17791) );
  INV_X1 U19861 ( .A(n17781), .ZN(n21049) );
  NAND2_X1 U19862 ( .A1(n21049), .A2(n21078), .ZN(n21066) );
  INV_X1 U19863 ( .A(n21028), .ZN(n21044) );
  NAND2_X1 U19864 ( .A1(n21044), .A2(n21078), .ZN(n21067) );
  AOI22_X1 U19865 ( .A1(n17840), .A2(n21066), .B1(n17885), .B2(n21067), .ZN(
        n17807) );
  NAND2_X1 U19866 ( .A1(n17783), .A2(n17782), .ZN(n17784) );
  XNOR2_X1 U19867 ( .A(n17784), .B(n21081), .ZN(n21076) );
  XNOR2_X1 U19868 ( .A(n17785), .B(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n20592) );
  OAI22_X1 U19869 ( .A1(n17786), .A2(n11199), .B1(n20592), .B2(n17809), .ZN(
        n17789) );
  INV_X1 U19870 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n21088) );
  OAI22_X1 U19871 ( .A1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n17787), .B1(
        n21223), .B2(n21088), .ZN(n17788) );
  AOI211_X1 U19872 ( .C1(n17886), .C2(n21076), .A(n17789), .B(n17788), .ZN(
        n17790) );
  OAI221_X1 U19873 ( .B1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n17791), 
        .C1(n21081), .C2(n17807), .A(n17790), .ZN(P3_U2800) );
  AOI211_X1 U19874 ( .C1(n21108), .C2(n17840), .A(
        P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B(n21107), .ZN(n17806) );
  AOI21_X1 U19875 ( .B1(n17793), .B2(n17792), .A(n21105), .ZN(n17794) );
  XNOR2_X1 U19876 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B(n17794), .ZN(
        n21072) );
  NAND2_X1 U19877 ( .A1(n21238), .A2(P3_REIP_REG_29__SCAN_IN), .ZN(n21073) );
  NAND2_X1 U19878 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n17795), .ZN(
        n17796) );
  OAI211_X1 U19879 ( .C1(n17798), .C2(n17797), .A(n21073), .B(n17796), .ZN(
        n17799) );
  AOI21_X1 U19880 ( .B1(n17886), .B2(n21072), .A(n17799), .ZN(n17805) );
  OAI21_X1 U19881 ( .B1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n17801), .A(
        n17800), .ZN(n20567) );
  OAI21_X1 U19882 ( .B1(n17803), .B2(n10962), .A(n11197), .ZN(n17804) );
  OAI211_X1 U19883 ( .C1(n17807), .C2(n17806), .A(n17805), .B(n17804), .ZN(
        P3_U2801) );
  NAND2_X1 U19884 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n21191), .ZN(
        n21197) );
  INV_X1 U19885 ( .A(n17808), .ZN(n20406) );
  OAI21_X1 U19886 ( .B1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n20392), .A(
        n20406), .ZN(n20395) );
  INV_X1 U19887 ( .A(n20395), .ZN(n17814) );
  AOI21_X1 U19888 ( .B1(n17810), .B2(n18884), .A(
        P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n17812) );
  INV_X1 U19889 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n21190) );
  OAI22_X1 U19890 ( .A1(n17812), .A2(n17811), .B1(n21223), .B2(n21190), .ZN(
        n17813) );
  AOI21_X1 U19891 ( .B1(n17814), .B2(n17961), .A(n17813), .ZN(n17819) );
  OAI21_X1 U19892 ( .B1(n17816), .B2(n21191), .A(n17815), .ZN(n21195) );
  AOI22_X1 U19893 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n17817), .B1(
        n17886), .B2(n21195), .ZN(n17818) );
  OAI211_X1 U19894 ( .C1(n17820), .C2(n21197), .A(n17819), .B(n17818), .ZN(
        P3_U2813) );
  AOI21_X1 U19895 ( .B1(n17821), .B2(n18884), .A(
        P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n17834) );
  INV_X1 U19896 ( .A(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n20365) );
  AOI21_X1 U19897 ( .B1(n20365), .B2(n17823), .A(n17822), .ZN(n20353) );
  AOI22_X1 U19898 ( .A1(n21238), .A2(P3_REIP_REG_14__SCAN_IN), .B1(n20353), 
        .B2(n17961), .ZN(n17832) );
  AOI21_X1 U19899 ( .B1(n20974), .B2(n17825), .A(n17824), .ZN(n20984) );
  INV_X1 U19900 ( .A(n17863), .ZN(n17846) );
  AOI21_X1 U19901 ( .B1(n17846), .B2(n20975), .A(n17826), .ZN(n17827) );
  XNOR2_X1 U19902 ( .A(n17827), .B(n20974), .ZN(n20989) );
  OAI21_X1 U19903 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n17828), .A(
        n20994), .ZN(n20983) );
  OAI22_X1 U19904 ( .A1(n20989), .A2(n17876), .B1(n17829), .B2(n20983), .ZN(
        n17830) );
  AOI21_X1 U19905 ( .B1(n17840), .B2(n20984), .A(n17830), .ZN(n17831) );
  OAI211_X1 U19906 ( .C1(n17834), .C2(n17833), .A(n17832), .B(n17831), .ZN(
        P3_U2816) );
  INV_X1 U19907 ( .A(n10978), .ZN(n17845) );
  INV_X1 U19908 ( .A(n20954), .ZN(n17860) );
  NOR2_X1 U19909 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n17860), .ZN(
        n20948) );
  AOI21_X1 U19910 ( .B1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n17860), .A(
        n20948), .ZN(n17844) );
  INV_X1 U19911 ( .A(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n20311) );
  NAND2_X1 U19912 ( .A1(n20310), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n17854) );
  AOI21_X1 U19913 ( .B1(n20311), .B2(n17854), .A(n17835), .ZN(n20314) );
  NAND2_X1 U19914 ( .A1(n20310), .A2(n18884), .ZN(n17852) );
  NAND2_X1 U19915 ( .A1(n10979), .A2(n17879), .ZN(n17962) );
  NAND3_X1 U19916 ( .A1(n17962), .A2(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .A3(
        n17852), .ZN(n17837) );
  NAND2_X1 U19917 ( .A1(n21238), .A2(P3_REIP_REG_11__SCAN_IN), .ZN(n17836) );
  OAI211_X1 U19918 ( .C1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .C2(n17852), .A(
        n17837), .B(n17836), .ZN(n17842) );
  AOI21_X1 U19919 ( .B1(n17846), .B2(n20954), .A(n17838), .ZN(n17839) );
  XNOR2_X1 U19920 ( .A(n17839), .B(n21209), .ZN(n20959) );
  AOI22_X1 U19921 ( .A1(n17840), .A2(n20952), .B1(n17885), .B2(n21176), .ZN(
        n17851) );
  OAI22_X1 U19922 ( .A1(n20959), .A2(n17876), .B1(n17851), .B2(n21209), .ZN(
        n17841) );
  AOI211_X1 U19923 ( .C1(n20314), .C2(n17961), .A(n17842), .B(n17841), .ZN(
        n17843) );
  OAI21_X1 U19924 ( .B1(n17845), .B2(n17844), .A(n17843), .ZN(P3_U2819) );
  OAI221_X1 U19925 ( .B1(n17846), .B2(n21115), .C1(n17846), .C2(n21241), .A(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n17850) );
  OAI221_X1 U19926 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n17864), .C1(
        n21241), .C2(n17863), .A(n17847), .ZN(n17848) );
  OAI221_X1 U19927 ( .B1(n17850), .B2(n21241), .C1(n17850), .C2(n17849), .A(
        n17848), .ZN(n21228) );
  INV_X1 U19928 ( .A(n17851), .ZN(n17873) );
  INV_X1 U19929 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n20306) );
  NOR2_X1 U19930 ( .A1(n21223), .A2(n20306), .ZN(n17858) );
  INV_X1 U19931 ( .A(n17852), .ZN(n17856) );
  INV_X1 U19932 ( .A(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n20284) );
  NAND4_X1 U19933 ( .A1(n20245), .A2(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A4(n18884), .ZN(n17869) );
  NOR2_X1 U19934 ( .A1(n20284), .A2(n17869), .ZN(n17867) );
  AOI21_X1 U19935 ( .B1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n17962), .A(
        n17867), .ZN(n17855) );
  NOR2_X1 U19936 ( .A1(n17853), .A2(n20186), .ZN(n20277) );
  OAI21_X1 U19937 ( .B1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n20277), .A(
        n17854), .ZN(n20291) );
  OAI22_X1 U19938 ( .A1(n17856), .A2(n17855), .B1(n17952), .B2(n20291), .ZN(
        n17857) );
  AOI211_X1 U19939 ( .C1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .C2(n17873), .A(
        n17858), .B(n17857), .ZN(n17862) );
  NAND3_X1 U19940 ( .A1(n17860), .A2(n17859), .A3(n10978), .ZN(n17861) );
  OAI211_X1 U19941 ( .C1(n21228), .C2(n17876), .A(n17862), .B(n17861), .ZN(
        P3_U2820) );
  NAND2_X1 U19942 ( .A1(n17864), .A2(n17863), .ZN(n17865) );
  XNOR2_X1 U19943 ( .A(n17865), .B(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n21247) );
  NAND2_X1 U19944 ( .A1(n17866), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n20279) );
  AOI21_X1 U19945 ( .B1(n20284), .B2(n20279), .A(n20277), .ZN(n20290) );
  INV_X1 U19946 ( .A(n17962), .ZN(n17868) );
  AOI211_X1 U19947 ( .C1(n17869), .C2(n20284), .A(n17868), .B(n17867), .ZN(
        n17871) );
  NAND2_X1 U19948 ( .A1(n21238), .A2(P3_REIP_REG_9__SCAN_IN), .ZN(n21244) );
  INV_X1 U19949 ( .A(n21244), .ZN(n17870) );
  AOI211_X1 U19950 ( .C1(n20290), .C2(n17961), .A(n17871), .B(n17870), .ZN(
        n17875) );
  AOI22_X1 U19951 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n17873), .B1(
        n10978), .B2(n21241), .ZN(n17874) );
  OAI211_X1 U19952 ( .C1(n21247), .C2(n17876), .A(n17875), .B(n17874), .ZN(
        P3_U2821) );
  OAI21_X1 U19953 ( .B1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n17878), .A(
        n17877), .ZN(n20939) );
  OAI21_X1 U19954 ( .B1(n20245), .B2(n17879), .A(n10979), .ZN(n17897) );
  AOI221_X1 U19955 ( .B1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .C1(n17880), .C2(n20264), .A(n19009), .ZN(n17882) );
  NOR2_X1 U19956 ( .A1(n17880), .A2(n20186), .ZN(n20266) );
  OAI21_X1 U19957 ( .B1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n20266), .A(
        n20279), .ZN(n20267) );
  INV_X1 U19958 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n20938) );
  OAI22_X1 U19959 ( .A1(n17952), .A2(n20267), .B1(n21223), .B2(n20938), .ZN(
        n17881) );
  AOI211_X1 U19960 ( .C1(n17897), .C2(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n17882), .B(n17881), .ZN(n17889) );
  XOR2_X1 U19961 ( .A(n17884), .B(n17883), .Z(n17887) );
  INV_X1 U19962 ( .A(n17887), .ZN(n20940) );
  AOI22_X1 U19963 ( .A1(n17887), .A2(n17886), .B1(n17885), .B2(n20940), .ZN(
        n17888) );
  OAI211_X1 U19964 ( .C1(n17971), .C2(n20939), .A(n17889), .B(n17888), .ZN(
        P3_U2822) );
  NAND2_X1 U19965 ( .A1(n20245), .A2(n18884), .ZN(n17900) );
  NAND2_X1 U19966 ( .A1(n20245), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n17901) );
  AOI21_X1 U19967 ( .B1(n11231), .B2(n17901), .A(n20266), .ZN(n20247) );
  AOI22_X1 U19968 ( .A1(n21238), .A2(P3_REIP_REG_7__SCAN_IN), .B1(n20247), 
        .B2(n17961), .ZN(n17899) );
  OAI21_X1 U19969 ( .B1(n17892), .B2(n17891), .A(n17890), .ZN(n17893) );
  XNOR2_X1 U19970 ( .A(n17893), .B(n20935), .ZN(n20927) );
  OAI21_X1 U19971 ( .B1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n17895), .A(
        n17894), .ZN(n20928) );
  OAI22_X1 U19972 ( .A1(n17971), .A2(n20927), .B1(n17970), .B2(n20928), .ZN(
        n17896) );
  AOI21_X1 U19973 ( .B1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n17897), .A(
        n17896), .ZN(n17898) );
  OAI211_X1 U19974 ( .C1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .C2(n17900), .A(
        n17899), .B(n17898), .ZN(P3_U2823) );
  NOR2_X1 U19975 ( .A1(n17903), .A2(n20186), .ZN(n20234) );
  OAI21_X1 U19976 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n20234), .A(
        n17901), .ZN(n20237) );
  NOR2_X1 U19977 ( .A1(n17903), .A2(n19009), .ZN(n17907) );
  OAI22_X1 U19978 ( .A1(n21223), .A2(n20250), .B1(n17971), .B2(n17902), .ZN(
        n17906) );
  OAI21_X1 U19979 ( .B1(n19009), .B2(n17903), .A(n17962), .ZN(n17916) );
  OAI22_X1 U19980 ( .A1(n20233), .A2(n17916), .B1(n17970), .B2(n17904), .ZN(
        n17905) );
  AOI211_X1 U19981 ( .C1(n17907), .C2(n20233), .A(n17906), .B(n17905), .ZN(
        n17908) );
  OAI21_X1 U19982 ( .B1(n17952), .B2(n20237), .A(n17908), .ZN(P3_U2824) );
  OAI21_X1 U19983 ( .B1(n17911), .B2(n17910), .A(n17909), .ZN(n20922) );
  INV_X1 U19984 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n17912) );
  NAND2_X1 U19985 ( .A1(n17913), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n20224) );
  AOI21_X1 U19986 ( .B1(n17912), .B2(n20224), .A(n20234), .ZN(n20226) );
  AOI21_X1 U19987 ( .B1(n17913), .B2(n10979), .A(
        P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n17917) );
  OAI21_X1 U19988 ( .B1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n17915), .A(
        n17914), .ZN(n20917) );
  OAI22_X1 U19989 ( .A1(n17917), .A2(n17916), .B1(n17970), .B2(n20917), .ZN(
        n17918) );
  AOI21_X1 U19990 ( .B1(n20226), .B2(n17961), .A(n17918), .ZN(n17919) );
  NAND2_X1 U19991 ( .A1(n21238), .A2(P3_REIP_REG_5__SCAN_IN), .ZN(n20916) );
  OAI211_X1 U19992 ( .C1(n17971), .C2(n20922), .A(n17919), .B(n20916), .ZN(
        P3_U2825) );
  NOR2_X1 U19993 ( .A1(n17923), .A2(n20186), .ZN(n20207) );
  OAI21_X1 U19994 ( .B1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n20207), .A(
        n20224), .ZN(n20215) );
  NOR3_X1 U19995 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n17923), .A3(
        n19009), .ZN(n17931) );
  INV_X1 U19996 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n20907) );
  OAI21_X1 U19997 ( .B1(n17922), .B2(n17921), .A(n17920), .ZN(n20906) );
  OAI22_X1 U19998 ( .A1(n21223), .A2(n20907), .B1(n17971), .B2(n20906), .ZN(
        n17930) );
  AOI21_X1 U19999 ( .B1(n17924), .B2(n17923), .A(n17954), .ZN(n17941) );
  OAI21_X1 U20000 ( .B1(n17927), .B2(n17926), .A(n17925), .ZN(n20912) );
  OAI22_X1 U20001 ( .A1(n17928), .A2(n17941), .B1(n17970), .B2(n20912), .ZN(
        n17929) );
  NOR3_X1 U20002 ( .A1(n17931), .A2(n17930), .A3(n17929), .ZN(n17932) );
  OAI21_X1 U20003 ( .B1(n17952), .B2(n20215), .A(n17932), .ZN(P3_U2826) );
  OAI21_X1 U20004 ( .B1(n17935), .B2(n17934), .A(n17933), .ZN(n20899) );
  INV_X1 U20005 ( .A(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17936) );
  NAND2_X1 U20006 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n17948) );
  AOI21_X1 U20007 ( .B1(n17936), .B2(n17948), .A(n20207), .ZN(n20197) );
  AOI21_X1 U20008 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n10979), .A(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17942) );
  OAI21_X1 U20009 ( .B1(n17939), .B2(n17938), .A(n17937), .ZN(n17940) );
  XNOR2_X1 U20010 ( .A(n17940), .B(n20915), .ZN(n20900) );
  OAI22_X1 U20011 ( .A1(n17942), .A2(n17941), .B1(n17970), .B2(n20900), .ZN(
        n17943) );
  AOI21_X1 U20012 ( .B1(n20197), .B2(n17961), .A(n17943), .ZN(n17944) );
  NAND2_X1 U20013 ( .A1(n21238), .A2(P3_REIP_REG_3__SCAN_IN), .ZN(n20903) );
  OAI211_X1 U20014 ( .C1(n17971), .C2(n20899), .A(n17944), .B(n20903), .ZN(
        P3_U2827) );
  OAI21_X1 U20015 ( .B1(n17947), .B2(n17946), .A(n17945), .ZN(n20888) );
  INV_X1 U20016 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n20187) );
  OAI21_X1 U20017 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A(n17948), .ZN(n20191) );
  OAI21_X1 U20018 ( .B1(n17951), .B2(n17950), .A(n17949), .ZN(n20889) );
  OAI22_X1 U20019 ( .A1(n17952), .A2(n20191), .B1(n17970), .B2(n20889), .ZN(
        n17953) );
  AOI221_X1 U20020 ( .B1(n17954), .B2(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .C1(
        n18884), .C2(n20187), .A(n17953), .ZN(n17955) );
  NAND2_X1 U20021 ( .A1(n21238), .A2(P3_REIP_REG_2__SCAN_IN), .ZN(n20893) );
  OAI211_X1 U20022 ( .C1(n17971), .C2(n20888), .A(n17955), .B(n20893), .ZN(
        P3_U2828) );
  OAI21_X1 U20023 ( .B1(n17965), .B2(n17959), .A(n17956), .ZN(n20874) );
  AOI21_X1 U20024 ( .B1(n17959), .B2(n17958), .A(n17957), .ZN(n20875) );
  INV_X1 U20025 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n20173) );
  OAI22_X1 U20026 ( .A1(n20875), .A2(n17971), .B1(n21223), .B2(n20173), .ZN(
        n17960) );
  AOI221_X1 U20027 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n17962), .C1(
        n20186), .C2(n17961), .A(n17960), .ZN(n17963) );
  OAI21_X1 U20028 ( .B1(n17970), .B2(n20874), .A(n17963), .ZN(P3_U2829) );
  NOR2_X1 U20029 ( .A1(n17965), .A2(n17964), .ZN(n20870) );
  INV_X1 U20030 ( .A(n20870), .ZN(n20869) );
  NAND3_X1 U20031 ( .A1(n20798), .A2(n17967), .A3(n10979), .ZN(n17968) );
  AOI22_X1 U20032 ( .A1(n21238), .A2(P3_REIP_REG_0__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17968), .ZN(n17969) );
  OAI221_X1 U20033 ( .B1(n20870), .B2(n17971), .C1(n20869), .C2(n17970), .A(
        n17969), .ZN(P3_U2830) );
  INV_X1 U20034 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n21275) );
  NAND2_X1 U20035 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18692), .ZN(
        n18712) );
  INV_X1 U20036 ( .A(n18712), .ZN(n18713) );
  NOR2_X1 U20037 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18692), .ZN(
        n18731) );
  NOR2_X1 U20038 ( .A1(n18713), .A2(n18731), .ZN(n17973) );
  OAI22_X1 U20039 ( .A1(n17974), .A2(n21275), .B1(n17973), .B2(n17972), .ZN(
        P3_U2866) );
  NAND2_X1 U20040 ( .A1(n17976), .A2(n17975), .ZN(n17979) );
  OAI21_X1 U20041 ( .B1(n17977), .B2(n18703), .A(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n17978) );
  OAI21_X1 U20042 ( .B1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n17979), .A(
        n17978), .ZN(P3_U2864) );
  NOR4_X1 U20043 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_12__SCAN_IN), .A3(P3_DATAWIDTH_REG_11__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_10__SCAN_IN), .ZN(n17983) );
  NOR4_X1 U20044 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_16__SCAN_IN), .A3(P3_DATAWIDTH_REG_15__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_14__SCAN_IN), .ZN(n17982) );
  NOR4_X1 U20045 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_4__SCAN_IN), .A3(P3_DATAWIDTH_REG_3__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_2__SCAN_IN), .ZN(n17981) );
  NOR4_X1 U20046 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_8__SCAN_IN), .A3(P3_DATAWIDTH_REG_7__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_6__SCAN_IN), .ZN(n17980) );
  NAND4_X1 U20047 ( .A1(n17983), .A2(n17982), .A3(n17981), .A4(n17980), .ZN(
        n17989) );
  NOR4_X1 U20048 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_28__SCAN_IN), .A3(P3_DATAWIDTH_REG_27__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_26__SCAN_IN), .ZN(n17987) );
  AOI211_X1 U20049 ( .C1(P3_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A(P3_DATAWIDTH_REG_31__SCAN_IN), .B(
        P3_DATAWIDTH_REG_30__SCAN_IN), .ZN(n17986) );
  NOR4_X1 U20050 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_20__SCAN_IN), .A3(P3_DATAWIDTH_REG_19__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_18__SCAN_IN), .ZN(n17985) );
  NOR4_X1 U20051 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_24__SCAN_IN), .A3(P3_DATAWIDTH_REG_23__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_22__SCAN_IN), .ZN(n17984) );
  NAND4_X1 U20052 ( .A1(n17987), .A2(n17986), .A3(n17985), .A4(n17984), .ZN(
        n17988) );
  NOR2_X1 U20053 ( .A1(n17989), .A2(n17988), .ZN(n17997) );
  INV_X1 U20054 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n18079) );
  OAI21_X1 U20055 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(P3_REIP_REG_0__SCAN_IN), 
        .A(n17997), .ZN(n17990) );
  OAI21_X1 U20056 ( .B1(n17997), .B2(n18079), .A(n17990), .ZN(P3_U3293) );
  INV_X1 U20057 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n18083) );
  AOI21_X1 U20058 ( .B1(P3_REIP_REG_0__SCAN_IN), .B2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n17991) );
  OAI221_X1 U20059 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(n17991), .C1(n20173), 
        .C2(P3_REIP_REG_0__SCAN_IN), .A(n17997), .ZN(n17992) );
  OAI21_X1 U20060 ( .B1(n17997), .B2(n18083), .A(n17992), .ZN(P3_U3292) );
  INV_X1 U20061 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n18081) );
  NOR3_X1 U20062 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A3(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n17994) );
  OAI21_X1 U20063 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(n17994), .A(n17997), .ZN(
        n17993) );
  OAI21_X1 U20064 ( .B1(n17997), .B2(n18081), .A(n17993), .ZN(P3_U2638) );
  INV_X1 U20065 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n21702) );
  AOI21_X1 U20066 ( .B1(n20173), .B2(n21702), .A(n17994), .ZN(n17996) );
  INV_X1 U20067 ( .A(P3_BYTEENABLE_REG_3__SCAN_IN), .ZN(n18085) );
  INV_X1 U20068 ( .A(n17997), .ZN(n17995) );
  AOI22_X1 U20069 ( .A1(n17997), .A2(n17996), .B1(n18085), .B2(n17995), .ZN(
        P3_U2639) );
  INV_X1 U20070 ( .A(P3_M_IO_N_REG_SCAN_IN), .ZN(n18086) );
  AOI22_X1 U20071 ( .A1(n21710), .A2(n17998), .B1(n18086), .B2(n21756), .ZN(
        P3_U3297) );
  INV_X1 U20072 ( .A(P3_W_R_N_REG_SCAN_IN), .ZN(n17999) );
  AOI22_X1 U20073 ( .A1(n21710), .A2(P3_READREQUEST_REG_SCAN_IN), .B1(n17999), 
        .B2(n21756), .ZN(P3_U3294) );
  AOI21_X1 U20074 ( .B1(n21758), .B2(n21706), .A(P3_D_C_N_REG_SCAN_IN), .ZN(
        n18000) );
  AOI22_X1 U20075 ( .A1(n21710), .A2(P3_CODEFETCH_REG_SCAN_IN), .B1(n18000), 
        .B2(n21756), .ZN(P3_U2635) );
  INV_X1 U20076 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n20793) );
  AOI22_X1 U20077 ( .A1(n21248), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n18032), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n18001) );
  OAI21_X1 U20078 ( .B1(n20793), .B2(n18018), .A(n18001), .ZN(P3_U2767) );
  INV_X1 U20079 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n20137) );
  AOI22_X1 U20080 ( .A1(n21248), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n18032), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n18002) );
  OAI21_X1 U20081 ( .B1(n20137), .B2(n18018), .A(n18002), .ZN(P3_U2766) );
  INV_X1 U20082 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n20663) );
  AOI22_X1 U20083 ( .A1(n21248), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n18032), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n18003) );
  OAI21_X1 U20084 ( .B1(n20663), .B2(n18018), .A(n18003), .ZN(P3_U2765) );
  INV_X1 U20085 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n20141) );
  AOI22_X1 U20086 ( .A1(n21248), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n18032), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n18004) );
  OAI21_X1 U20087 ( .B1(n20141), .B2(n18018), .A(n18004), .ZN(P3_U2764) );
  INV_X1 U20088 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n20650) );
  AOI22_X1 U20089 ( .A1(n21248), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n18032), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n18005) );
  OAI21_X1 U20090 ( .B1(n20650), .B2(n18018), .A(n18005), .ZN(P3_U2763) );
  INV_X1 U20091 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n18007) );
  AOI22_X1 U20092 ( .A1(n21248), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n18032), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n18006) );
  OAI21_X1 U20093 ( .B1(n18007), .B2(n18018), .A(n18006), .ZN(P3_U2762) );
  INV_X1 U20094 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n20614) );
  AOI22_X1 U20095 ( .A1(n21248), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n18032), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n18008) );
  OAI21_X1 U20096 ( .B1(n20614), .B2(n18018), .A(n18008), .ZN(P3_U2761) );
  INV_X1 U20097 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n20147) );
  AOI22_X1 U20098 ( .A1(n21248), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n18032), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n18009) );
  OAI21_X1 U20099 ( .B1(n20147), .B2(n18018), .A(n18009), .ZN(P3_U2760) );
  INV_X1 U20100 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n20777) );
  AOI22_X1 U20101 ( .A1(n21248), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n18032), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n18010) );
  OAI21_X1 U20102 ( .B1(n20777), .B2(n18018), .A(n18010), .ZN(P3_U2759) );
  INV_X1 U20103 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n20668) );
  AOI22_X1 U20104 ( .A1(n18030), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n18032), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n18011) );
  OAI21_X1 U20105 ( .B1(n20668), .B2(n18018), .A(n18011), .ZN(P3_U2758) );
  INV_X1 U20106 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n20667) );
  AOI22_X1 U20107 ( .A1(n18030), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n18032), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n18012) );
  OAI21_X1 U20108 ( .B1(n20667), .B2(n18018), .A(n18012), .ZN(P3_U2757) );
  INV_X1 U20109 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n20627) );
  AOI22_X1 U20110 ( .A1(n18030), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n18032), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n18013) );
  OAI21_X1 U20111 ( .B1(n20627), .B2(n18018), .A(n18013), .ZN(P3_U2756) );
  INV_X1 U20112 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n20669) );
  AOI22_X1 U20113 ( .A1(n18030), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n18032), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n18014) );
  OAI21_X1 U20114 ( .B1(n20669), .B2(n18018), .A(n18014), .ZN(P3_U2755) );
  INV_X1 U20115 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n20670) );
  AOI22_X1 U20116 ( .A1(n18030), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n18032), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n18015) );
  OAI21_X1 U20117 ( .B1(n20670), .B2(n18018), .A(n18015), .ZN(P3_U2754) );
  INV_X1 U20118 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n20157) );
  AOI22_X1 U20119 ( .A1(n18030), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n18032), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n18016) );
  OAI21_X1 U20120 ( .B1(n20157), .B2(n18018), .A(n18016), .ZN(P3_U2753) );
  INV_X1 U20121 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n20770) );
  AOI22_X1 U20122 ( .A1(n18030), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n18032), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n18017) );
  OAI21_X1 U20123 ( .B1(n20770), .B2(n18018), .A(n18017), .ZN(P3_U2752) );
  INV_X1 U20124 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n18021) );
  NAND2_X1 U20125 ( .A1(n18019), .A2(n20166), .ZN(n18040) );
  AOI22_X1 U20126 ( .A1(n18030), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n18032), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n18020) );
  OAI21_X1 U20127 ( .B1(n18021), .B2(n18040), .A(n18020), .ZN(P3_U2751) );
  INV_X1 U20128 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n20672) );
  AOI22_X1 U20129 ( .A1(n18030), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n18032), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n18022) );
  OAI21_X1 U20130 ( .B1(n20672), .B2(n18040), .A(n18022), .ZN(P3_U2750) );
  INV_X1 U20131 ( .A(P3_EAX_REG_18__SCAN_IN), .ZN(n18024) );
  AOI22_X1 U20132 ( .A1(n18030), .A2(P3_UWORD_REG_2__SCAN_IN), .B1(n18032), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n18023) );
  OAI21_X1 U20133 ( .B1(n18024), .B2(n18040), .A(n18023), .ZN(P3_U2749) );
  INV_X1 U20134 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n20694) );
  AOI22_X1 U20135 ( .A1(n21248), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n18032), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n18025) );
  OAI21_X1 U20136 ( .B1(n20694), .B2(n18040), .A(n18025), .ZN(P3_U2748) );
  INV_X1 U20137 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n20682) );
  AOI22_X1 U20138 ( .A1(n21248), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n18032), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n18026) );
  OAI21_X1 U20139 ( .B1(n20682), .B2(n18040), .A(n18026), .ZN(P3_U2747) );
  INV_X1 U20140 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n20683) );
  AOI22_X1 U20141 ( .A1(n21248), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n18032), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n18027) );
  OAI21_X1 U20142 ( .B1(n20683), .B2(n18040), .A(n18027), .ZN(P3_U2746) );
  INV_X1 U20143 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n20709) );
  AOI22_X1 U20144 ( .A1(n21248), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n18032), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n18028) );
  OAI21_X1 U20145 ( .B1(n20709), .B2(n18040), .A(n18028), .ZN(P3_U2745) );
  INV_X1 U20146 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n20122) );
  AOI22_X1 U20147 ( .A1(n21248), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n18032), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n18029) );
  OAI21_X1 U20148 ( .B1(n20122), .B2(n18040), .A(n18029), .ZN(P3_U2744) );
  INV_X1 U20149 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n20124) );
  AOI22_X1 U20150 ( .A1(n18030), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n18032), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n18031) );
  OAI21_X1 U20151 ( .B1(n20124), .B2(n18040), .A(n18031), .ZN(P3_U2743) );
  INV_X1 U20152 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n18034) );
  AOI22_X1 U20153 ( .A1(n21248), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n18032), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n18033) );
  OAI21_X1 U20154 ( .B1(n18034), .B2(n18040), .A(n18033), .ZN(P3_U2742) );
  INV_X1 U20155 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n20720) );
  AOI22_X1 U20156 ( .A1(n21248), .A2(P3_UWORD_REG_10__SCAN_IN), .B1(n18032), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n18035) );
  OAI21_X1 U20157 ( .B1(n20720), .B2(n18040), .A(n18035), .ZN(P3_U2741) );
  INV_X1 U20158 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n20128) );
  AOI22_X1 U20159 ( .A1(n21248), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n18032), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n18036) );
  OAI21_X1 U20160 ( .B1(n20128), .B2(n18040), .A(n18036), .ZN(P3_U2740) );
  INV_X1 U20161 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n20738) );
  AOI22_X1 U20162 ( .A1(n21248), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n18032), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n18037) );
  OAI21_X1 U20163 ( .B1(n20738), .B2(n18040), .A(n18037), .ZN(P3_U2739) );
  INV_X1 U20164 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n20131) );
  AOI22_X1 U20165 ( .A1(n21248), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n18032), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n18038) );
  OAI21_X1 U20166 ( .B1(n20131), .B2(n18040), .A(n18038), .ZN(P3_U2738) );
  INV_X1 U20167 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n20133) );
  AOI22_X1 U20168 ( .A1(n21248), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(n18032), 
        .B2(P3_DATAO_REG_30__SCAN_IN), .ZN(n18039) );
  OAI21_X1 U20169 ( .B1(n20133), .B2(n18040), .A(n18039), .ZN(P3_U2737) );
  NOR2_X1 U20170 ( .A1(P3_ADS_N_REG_SCAN_IN), .A2(n18041), .ZN(n18042) );
  NOR2_X1 U20171 ( .A1(n21710), .A2(n18042), .ZN(P3_U2633) );
  OR2_X1 U20172 ( .A1(P3_STATE_REG_2__SCAN_IN), .A2(n21756), .ZN(n18073) );
  INV_X1 U20173 ( .A(n18073), .ZN(n18075) );
  AOI22_X1 U20174 ( .A1(n18075), .A2(P3_REIP_REG_2__SCAN_IN), .B1(
        P3_ADDRESS_REG_0__SCAN_IN), .B2(n21756), .ZN(n18043) );
  OAI21_X1 U20175 ( .B1(n18077), .B2(n20173), .A(n18043), .ZN(P3_U3032) );
  INV_X1 U20176 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n20199) );
  AOI22_X1 U20177 ( .A1(P3_REIP_REG_2__SCAN_IN), .A2(n18071), .B1(
        P3_ADDRESS_REG_1__SCAN_IN), .B2(n21756), .ZN(n18044) );
  OAI21_X1 U20178 ( .B1(n20199), .B2(n18073), .A(n18044), .ZN(P3_U3033) );
  AOI22_X1 U20179 ( .A1(n18075), .A2(P3_REIP_REG_4__SCAN_IN), .B1(
        P3_ADDRESS_REG_2__SCAN_IN), .B2(n21756), .ZN(n18045) );
  OAI21_X1 U20180 ( .B1(n18077), .B2(n20199), .A(n18045), .ZN(P3_U3034) );
  AOI22_X1 U20181 ( .A1(n18075), .A2(P3_REIP_REG_5__SCAN_IN), .B1(
        P3_ADDRESS_REG_3__SCAN_IN), .B2(n21756), .ZN(n18046) );
  OAI21_X1 U20182 ( .B1(n18077), .B2(n20907), .A(n18046), .ZN(P3_U3035) );
  AOI22_X1 U20183 ( .A1(P3_REIP_REG_5__SCAN_IN), .A2(n18071), .B1(
        P3_ADDRESS_REG_4__SCAN_IN), .B2(n21756), .ZN(n18047) );
  OAI21_X1 U20184 ( .B1(n20250), .B2(n18073), .A(n18047), .ZN(P3_U3036) );
  AOI22_X1 U20185 ( .A1(n18075), .A2(P3_REIP_REG_7__SCAN_IN), .B1(
        P3_ADDRESS_REG_5__SCAN_IN), .B2(n21756), .ZN(n18048) );
  OAI21_X1 U20186 ( .B1(n18077), .B2(n20250), .A(n18048), .ZN(P3_U3037) );
  INV_X1 U20187 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n20254) );
  AOI22_X1 U20188 ( .A1(n18075), .A2(P3_REIP_REG_8__SCAN_IN), .B1(
        P3_ADDRESS_REG_6__SCAN_IN), .B2(n21756), .ZN(n18049) );
  OAI21_X1 U20189 ( .B1(n18077), .B2(n20254), .A(n18049), .ZN(P3_U3038) );
  AOI22_X1 U20190 ( .A1(n18075), .A2(P3_REIP_REG_9__SCAN_IN), .B1(
        P3_ADDRESS_REG_7__SCAN_IN), .B2(n21756), .ZN(n18050) );
  OAI21_X1 U20191 ( .B1(n18077), .B2(n20938), .A(n18050), .ZN(P3_U3039) );
  INV_X1 U20192 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n20283) );
  AOI22_X1 U20193 ( .A1(n18075), .A2(P3_REIP_REG_10__SCAN_IN), .B1(
        P3_ADDRESS_REG_8__SCAN_IN), .B2(n21756), .ZN(n18051) );
  OAI21_X1 U20194 ( .B1(n18077), .B2(n20283), .A(n18051), .ZN(P3_U3040) );
  AOI22_X1 U20195 ( .A1(n18075), .A2(P3_REIP_REG_11__SCAN_IN), .B1(
        P3_ADDRESS_REG_9__SCAN_IN), .B2(n21756), .ZN(n18052) );
  OAI21_X1 U20196 ( .B1(n18077), .B2(n20306), .A(n18052), .ZN(P3_U3041) );
  INV_X1 U20197 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n20340) );
  AOI22_X1 U20198 ( .A1(P3_REIP_REG_11__SCAN_IN), .A2(n18071), .B1(
        P3_ADDRESS_REG_10__SCAN_IN), .B2(n21756), .ZN(n18053) );
  OAI21_X1 U20199 ( .B1(n20340), .B2(n18073), .A(n18053), .ZN(P3_U3042) );
  AOI22_X1 U20200 ( .A1(n18075), .A2(P3_REIP_REG_13__SCAN_IN), .B1(
        P3_ADDRESS_REG_11__SCAN_IN), .B2(n21756), .ZN(n18054) );
  OAI21_X1 U20201 ( .B1(n18077), .B2(n20340), .A(n18054), .ZN(P3_U3043) );
  INV_X1 U20202 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n20336) );
  AOI22_X1 U20203 ( .A1(n18075), .A2(P3_REIP_REG_14__SCAN_IN), .B1(
        P3_ADDRESS_REG_12__SCAN_IN), .B2(n21756), .ZN(n18055) );
  OAI21_X1 U20204 ( .B1(n18077), .B2(n20336), .A(n18055), .ZN(P3_U3044) );
  INV_X1 U20205 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n20355) );
  AOI22_X1 U20206 ( .A1(n18075), .A2(P3_REIP_REG_15__SCAN_IN), .B1(
        P3_ADDRESS_REG_13__SCAN_IN), .B2(n21756), .ZN(n18056) );
  OAI21_X1 U20207 ( .B1(n18077), .B2(n20355), .A(n18056), .ZN(P3_U3045) );
  INV_X1 U20208 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n20376) );
  AOI22_X1 U20209 ( .A1(n18075), .A2(P3_REIP_REG_16__SCAN_IN), .B1(
        P3_ADDRESS_REG_14__SCAN_IN), .B2(n21756), .ZN(n18057) );
  OAI21_X1 U20210 ( .B1(n18077), .B2(n20376), .A(n18057), .ZN(P3_U3046) );
  INV_X1 U20211 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n20389) );
  AOI22_X1 U20212 ( .A1(n18075), .A2(P3_REIP_REG_17__SCAN_IN), .B1(
        P3_ADDRESS_REG_15__SCAN_IN), .B2(n21756), .ZN(n18058) );
  OAI21_X1 U20213 ( .B1(n18077), .B2(n20389), .A(n18058), .ZN(P3_U3047) );
  AOI22_X1 U20214 ( .A1(n18075), .A2(P3_REIP_REG_18__SCAN_IN), .B1(
        P3_ADDRESS_REG_16__SCAN_IN), .B2(n21756), .ZN(n18059) );
  OAI21_X1 U20215 ( .B1(n18077), .B2(n21190), .A(n18059), .ZN(P3_U3048) );
  INV_X1 U20216 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n20418) );
  AOI22_X1 U20217 ( .A1(n18075), .A2(P3_REIP_REG_19__SCAN_IN), .B1(
        P3_ADDRESS_REG_17__SCAN_IN), .B2(n21756), .ZN(n18060) );
  OAI21_X1 U20218 ( .B1(n18077), .B2(n20418), .A(n18060), .ZN(P3_U3049) );
  INV_X1 U20219 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n20446) );
  AOI22_X1 U20220 ( .A1(P3_REIP_REG_19__SCAN_IN), .A2(n18071), .B1(
        P3_ADDRESS_REG_18__SCAN_IN), .B2(n21756), .ZN(n18061) );
  OAI21_X1 U20221 ( .B1(n20446), .B2(n18073), .A(n18061), .ZN(P3_U3050) );
  AOI22_X1 U20222 ( .A1(n18075), .A2(P3_REIP_REG_21__SCAN_IN), .B1(
        P3_ADDRESS_REG_19__SCAN_IN), .B2(n21756), .ZN(n18062) );
  OAI21_X1 U20223 ( .B1(n18077), .B2(n20446), .A(n18062), .ZN(P3_U3051) );
  AOI22_X1 U20224 ( .A1(n18075), .A2(P3_REIP_REG_22__SCAN_IN), .B1(
        P3_ADDRESS_REG_20__SCAN_IN), .B2(n21756), .ZN(n18063) );
  OAI21_X1 U20225 ( .B1(n18077), .B2(n20458), .A(n18063), .ZN(P3_U3052) );
  AOI22_X1 U20226 ( .A1(n18075), .A2(P3_REIP_REG_23__SCAN_IN), .B1(
        P3_ADDRESS_REG_21__SCAN_IN), .B2(n21756), .ZN(n18064) );
  OAI21_X1 U20227 ( .B1(n18077), .B2(n20473), .A(n18064), .ZN(P3_U3053) );
  AOI22_X1 U20228 ( .A1(n18075), .A2(P3_REIP_REG_24__SCAN_IN), .B1(
        P3_ADDRESS_REG_22__SCAN_IN), .B2(n21756), .ZN(n18065) );
  OAI21_X1 U20229 ( .B1(n18077), .B2(n18066), .A(n18065), .ZN(P3_U3054) );
  AOI22_X1 U20230 ( .A1(n18075), .A2(P3_REIP_REG_25__SCAN_IN), .B1(
        P3_ADDRESS_REG_23__SCAN_IN), .B2(n21756), .ZN(n18067) );
  OAI21_X1 U20231 ( .B1(n18077), .B2(n20505), .A(n18067), .ZN(P3_U3055) );
  AOI22_X1 U20232 ( .A1(n18075), .A2(P3_REIP_REG_26__SCAN_IN), .B1(
        P3_ADDRESS_REG_24__SCAN_IN), .B2(n21756), .ZN(n18068) );
  OAI21_X1 U20233 ( .B1(n18077), .B2(n20506), .A(n18068), .ZN(P3_U3056) );
  INV_X1 U20234 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n20528) );
  AOI22_X1 U20235 ( .A1(n18075), .A2(P3_REIP_REG_27__SCAN_IN), .B1(
        P3_ADDRESS_REG_25__SCAN_IN), .B2(n21756), .ZN(n18069) );
  OAI21_X1 U20236 ( .B1(n18077), .B2(n20528), .A(n18069), .ZN(P3_U3057) );
  INV_X1 U20237 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n20541) );
  AOI22_X1 U20238 ( .A1(n18075), .A2(P3_REIP_REG_28__SCAN_IN), .B1(
        P3_ADDRESS_REG_26__SCAN_IN), .B2(n21756), .ZN(n18070) );
  OAI21_X1 U20239 ( .B1(n18077), .B2(n20541), .A(n18070), .ZN(P3_U3058) );
  INV_X1 U20240 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n20570) );
  AOI22_X1 U20241 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(n18071), .B1(
        P3_ADDRESS_REG_27__SCAN_IN), .B2(n21756), .ZN(n18072) );
  OAI21_X1 U20242 ( .B1(n20570), .B2(n18073), .A(n18072), .ZN(P3_U3059) );
  AOI22_X1 U20243 ( .A1(n18075), .A2(P3_REIP_REG_30__SCAN_IN), .B1(
        P3_ADDRESS_REG_28__SCAN_IN), .B2(n21756), .ZN(n18074) );
  OAI21_X1 U20244 ( .B1(n18077), .B2(n20570), .A(n18074), .ZN(P3_U3060) );
  AOI22_X1 U20245 ( .A1(n18075), .A2(P3_REIP_REG_31__SCAN_IN), .B1(
        P3_ADDRESS_REG_29__SCAN_IN), .B2(n21756), .ZN(n18076) );
  OAI21_X1 U20246 ( .B1(n18077), .B2(n21088), .A(n18076), .ZN(P3_U3061) );
  INV_X1 U20247 ( .A(P3_BE_N_REG_0__SCAN_IN), .ZN(n18078) );
  AOI22_X1 U20248 ( .A1(n21710), .A2(n18079), .B1(n18078), .B2(n21756), .ZN(
        P3_U3277) );
  INV_X1 U20249 ( .A(P3_BE_N_REG_1__SCAN_IN), .ZN(n18080) );
  AOI22_X1 U20250 ( .A1(n21710), .A2(n18081), .B1(n18080), .B2(n21756), .ZN(
        P3_U3276) );
  INV_X1 U20251 ( .A(P3_BE_N_REG_2__SCAN_IN), .ZN(n18082) );
  AOI22_X1 U20252 ( .A1(n21710), .A2(n18083), .B1(n18082), .B2(n21756), .ZN(
        P3_U3275) );
  INV_X1 U20253 ( .A(P3_BE_N_REG_3__SCAN_IN), .ZN(n18084) );
  AOI22_X1 U20254 ( .A1(n21710), .A2(n18085), .B1(n18084), .B2(n21756), .ZN(
        P3_U3274) );
  NOR4_X1 U20255 ( .A1(P3_BE_N_REG_1__SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(P3_BE_N_REG_2__SCAN_IN), .A4(P3_BE_N_REG_0__SCAN_IN), .ZN(n18088)
         );
  NOR4_X1 U20256 ( .A1(P3_ADS_N_REG_SCAN_IN), .A2(P3_D_C_N_REG_SCAN_IN), .A3(
        P3_W_R_N_REG_SCAN_IN), .A4(n18086), .ZN(n18087) );
  NAND3_X1 U20257 ( .A1(n18088), .A2(n18087), .A3(U215), .ZN(U213) );
  NOR2_X1 U20258 ( .A1(n18630), .A2(n19264), .ZN(n18094) );
  INV_X1 U20259 ( .A(n21735), .ZN(n18089) );
  OAI21_X1 U20260 ( .B1(n18089), .B2(n21695), .A(n12760), .ZN(n18092) );
  NAND3_X1 U20261 ( .A1(n18089), .A2(n19676), .A3(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n18091) );
  MUX2_X1 U20262 ( .A(n18092), .B(n18091), .S(n18090), .Z(n18093) );
  OAI21_X1 U20263 ( .B1(n18094), .B2(n18644), .A(n18093), .ZN(n18101) );
  NAND4_X1 U20264 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_STATE2_REG_2__SCAN_IN), .A3(n13554), .A4(n21729), .ZN(n18097) );
  INV_X1 U20265 ( .A(n18095), .ZN(n18096) );
  OAI211_X1 U20266 ( .C1(n18099), .C2(n18098), .A(n18097), .B(n18096), .ZN(
        n18100) );
  MUX2_X1 U20267 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .B(n18101), .S(n18100), 
        .Z(P2_U3610) );
  NAND2_X1 U20268 ( .A1(n18493), .A2(n10964), .ZN(n18513) );
  NOR2_X1 U20269 ( .A1(n18453), .A2(n18518), .ZN(n18105) );
  OAI22_X1 U20270 ( .A1(n18440), .A2(n18103), .B1(n18502), .B2(n18102), .ZN(
        n18104) );
  AOI211_X1 U20271 ( .C1(n18106), .C2(n18457), .A(n18105), .B(n18104), .ZN(
        n18107) );
  OAI21_X1 U20272 ( .B1(n18108), .B2(n18499), .A(n18107), .ZN(n18109) );
  AOI21_X1 U20273 ( .B1(n19151), .B2(n18119), .A(n18109), .ZN(n18111) );
  NOR2_X1 U20274 ( .A1(n10964), .A2(n18634), .ZN(n18347) );
  OAI21_X1 U20275 ( .B1(n18473), .B2(n18347), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n18110) );
  OAI211_X1 U20276 ( .C1(n18112), .C2(n18513), .A(n18111), .B(n18110), .ZN(
        P2_U2855) );
  INV_X1 U20277 ( .A(n18113), .ZN(n18114) );
  AOI22_X1 U20278 ( .A1(n18471), .A2(n18114), .B1(n18473), .B2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n18115) );
  OAI21_X1 U20279 ( .B1(n18502), .B2(n12779), .A(n18115), .ZN(n18118) );
  OAI22_X1 U20280 ( .A1(n18440), .A2(n12777), .B1(n18453), .B2(n18116), .ZN(
        n18117) );
  AOI211_X1 U20281 ( .C1(n18526), .C2(n18509), .A(n18118), .B(n18117), .ZN(
        n18122) );
  AOI22_X1 U20282 ( .A1(n18347), .A2(n18120), .B1(n19168), .B2(n18119), .ZN(
        n18121) );
  OAI211_X1 U20283 ( .C1(n18634), .C2(n18123), .A(n18122), .B(n18121), .ZN(
        P2_U2854) );
  OAI22_X1 U20284 ( .A1(n18124), .A2(n18486), .B1(n13825), .B2(n18502), .ZN(
        n18131) );
  NAND2_X1 U20285 ( .A1(n18510), .A2(n18579), .ZN(n18129) );
  OR2_X1 U20286 ( .A1(n18440), .A2(n18125), .ZN(n18128) );
  NAND2_X1 U20287 ( .A1(n18457), .A2(n18126), .ZN(n18127) );
  NAND4_X1 U20288 ( .A1(n18129), .A2(n18128), .A3(n18589), .A4(n18127), .ZN(
        n18130) );
  NOR2_X1 U20289 ( .A1(n18131), .A2(n18130), .ZN(n18132) );
  OAI21_X1 U20290 ( .B1(n19405), .B2(n18133), .A(n18132), .ZN(n18134) );
  INV_X1 U20291 ( .A(n18134), .ZN(n18140) );
  NAND2_X1 U20292 ( .A1(n18136), .A2(n18135), .ZN(n18146) );
  AND2_X1 U20293 ( .A1(n10964), .A2(n18146), .ZN(n18138) );
  AOI21_X1 U20294 ( .B1(n18147), .B2(n18138), .A(n18634), .ZN(n18137) );
  OAI21_X1 U20295 ( .B1(n18147), .B2(n18138), .A(n18137), .ZN(n18139) );
  OAI211_X1 U20296 ( .C1(n18581), .C2(n18499), .A(n18140), .B(n18139), .ZN(
        P2_U2851) );
  INV_X1 U20297 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n18154) );
  NAND2_X1 U20298 ( .A1(n18331), .A2(P2_REIP_REG_5__SCAN_IN), .ZN(n18145) );
  INV_X1 U20299 ( .A(n18141), .ZN(n18142) );
  NAND2_X1 U20300 ( .A1(n18457), .A2(n18142), .ZN(n18144) );
  OR2_X1 U20301 ( .A1(n18440), .A2(n13848), .ZN(n18143) );
  AND4_X1 U20302 ( .A1(n18145), .A2(n18589), .A3(n18144), .A4(n18143), .ZN(
        n18153) );
  NOR2_X1 U20303 ( .A1(n18147), .A2(n18146), .ZN(n18159) );
  NOR2_X1 U20304 ( .A1(n16641), .A2(n18159), .ZN(n18148) );
  XNOR2_X1 U20305 ( .A(n18158), .B(n18148), .ZN(n18151) );
  OAI22_X1 U20306 ( .A1(n18453), .A2(n19409), .B1(n18499), .B2(n18149), .ZN(
        n18150) );
  AOI21_X1 U20307 ( .B1(n18151), .B2(n18493), .A(n18150), .ZN(n18152) );
  OAI211_X1 U20308 ( .C1(n18154), .C2(n18486), .A(n18153), .B(n18152), .ZN(
        P2_U2850) );
  OAI21_X1 U20309 ( .B1(n18502), .B2(n13834), .A(n18589), .ZN(n18157) );
  NOR2_X1 U20310 ( .A1(n18155), .A2(n18504), .ZN(n18156) );
  AOI211_X1 U20311 ( .C1(n18250), .C2(P2_EBX_REG_6__SCAN_IN), .A(n18157), .B(
        n18156), .ZN(n18166) );
  NAND2_X1 U20312 ( .A1(n18159), .A2(n18158), .ZN(n18168) );
  NAND2_X1 U20313 ( .A1(n10964), .A2(n18168), .ZN(n18160) );
  XNOR2_X1 U20314 ( .A(n18169), .B(n18160), .ZN(n18164) );
  OAI22_X1 U20315 ( .A1(n18453), .A2(n18162), .B1(n18499), .B2(n18161), .ZN(
        n18163) );
  AOI21_X1 U20316 ( .B1(n18261), .B2(n18164), .A(n18163), .ZN(n18165) );
  OAI211_X1 U20317 ( .C1(n18167), .C2(n18486), .A(n18166), .B(n18165), .ZN(
        P2_U2849) );
  NOR2_X1 U20318 ( .A1(n18169), .A2(n18168), .ZN(n18187) );
  NOR2_X1 U20319 ( .A1(n16641), .A2(n18187), .ZN(n18170) );
  XOR2_X1 U20320 ( .A(n18186), .B(n18170), .Z(n18180) );
  NOR2_X1 U20321 ( .A1(n18440), .A2(n18171), .ZN(n18172) );
  AOI211_X1 U20322 ( .C1(P2_REIP_REG_7__SCAN_IN), .C2(n18331), .A(n18572), .B(
        n18172), .ZN(n18173) );
  OAI21_X1 U20323 ( .B1(n18174), .B2(n18504), .A(n18173), .ZN(n18178) );
  OAI22_X1 U20324 ( .A1(n18453), .A2(n18176), .B1(n18499), .B2(n18175), .ZN(
        n18177) );
  AOI211_X1 U20325 ( .C1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .C2(n18507), .A(
        n18178), .B(n18177), .ZN(n18179) );
  OAI21_X1 U20326 ( .B1(n18634), .B2(n18180), .A(n18179), .ZN(P2_U2848) );
  INV_X1 U20327 ( .A(n18181), .ZN(n18185) );
  AOI22_X1 U20328 ( .A1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n18507), .B1(
        P2_REIP_REG_8__SCAN_IN), .B2(n18331), .ZN(n18182) );
  OAI211_X1 U20329 ( .C1(n18440), .C2(n18183), .A(n18182), .B(n18589), .ZN(
        n18184) );
  AOI21_X1 U20330 ( .B1(n18185), .B2(n18471), .A(n18184), .ZN(n18191) );
  NAND2_X1 U20331 ( .A1(n18187), .A2(n18186), .ZN(n18193) );
  NAND2_X1 U20332 ( .A1(n10964), .A2(n18193), .ZN(n18188) );
  XNOR2_X1 U20333 ( .A(n18194), .B(n18188), .ZN(n18189) );
  AOI22_X1 U20334 ( .A1(n18493), .A2(n18189), .B1(n18510), .B2(n18566), .ZN(
        n18190) );
  OAI211_X1 U20335 ( .C1(n18499), .C2(n18192), .A(n18191), .B(n18190), .ZN(
        P2_U2847) );
  NOR2_X1 U20336 ( .A1(n18194), .A2(n18193), .ZN(n18213) );
  NOR2_X1 U20337 ( .A1(n16641), .A2(n18213), .ZN(n18195) );
  XNOR2_X1 U20338 ( .A(n18195), .B(n18211), .ZN(n18206) );
  INV_X1 U20339 ( .A(n18196), .ZN(n18200) );
  NOR2_X1 U20340 ( .A1(n18440), .A2(n18197), .ZN(n18198) );
  AOI211_X1 U20341 ( .C1(P2_REIP_REG_9__SCAN_IN), .C2(n18331), .A(n18572), .B(
        n18198), .ZN(n18199) );
  OAI21_X1 U20342 ( .B1(n18200), .B2(n18504), .A(n18199), .ZN(n18204) );
  OAI22_X1 U20343 ( .A1(n18202), .A2(n18499), .B1(n18201), .B2(n18453), .ZN(
        n18203) );
  AOI211_X1 U20344 ( .C1(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .C2(n18473), .A(
        n18204), .B(n18203), .ZN(n18205) );
  OAI21_X1 U20345 ( .B1(n18634), .B2(n18206), .A(n18205), .ZN(P2_U2846) );
  INV_X1 U20346 ( .A(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n18220) );
  NAND2_X1 U20347 ( .A1(n18250), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n18207) );
  OAI211_X1 U20348 ( .C1(n13922), .C2(n18502), .A(n18207), .B(n18589), .ZN(
        n18208) );
  AOI21_X1 U20349 ( .B1(n18209), .B2(n18457), .A(n18208), .ZN(n18219) );
  INV_X1 U20350 ( .A(n18210), .ZN(n18222) );
  INV_X1 U20351 ( .A(n18211), .ZN(n18212) );
  NAND2_X1 U20352 ( .A1(n18213), .A2(n18212), .ZN(n18221) );
  NAND2_X1 U20353 ( .A1(n10964), .A2(n18221), .ZN(n18214) );
  XNOR2_X1 U20354 ( .A(n18222), .B(n18214), .ZN(n18217) );
  OAI22_X1 U20355 ( .A1(n18215), .A2(n18499), .B1(n19132), .B2(n18453), .ZN(
        n18216) );
  AOI21_X1 U20356 ( .B1(n18261), .B2(n18217), .A(n18216), .ZN(n18218) );
  OAI211_X1 U20357 ( .C1(n18220), .C2(n18486), .A(n18219), .B(n18218), .ZN(
        P2_U2845) );
  NOR2_X1 U20358 ( .A1(n18222), .A2(n18221), .ZN(n18243) );
  NOR2_X1 U20359 ( .A1(n16641), .A2(n18243), .ZN(n18223) );
  XNOR2_X1 U20360 ( .A(n18223), .B(n18241), .ZN(n18234) );
  INV_X1 U20361 ( .A(n18224), .ZN(n18228) );
  NOR2_X1 U20362 ( .A1(n18440), .A2(n18225), .ZN(n18226) );
  AOI211_X1 U20363 ( .C1(P2_REIP_REG_11__SCAN_IN), .C2(n18331), .A(n18572), 
        .B(n18226), .ZN(n18227) );
  OAI21_X1 U20364 ( .B1(n18228), .B2(n18504), .A(n18227), .ZN(n18232) );
  OAI22_X1 U20365 ( .A1(n18230), .A2(n18499), .B1(n18229), .B2(n18453), .ZN(
        n18231) );
  AOI211_X1 U20366 ( .C1(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .C2(n18473), .A(
        n18232), .B(n18231), .ZN(n18233) );
  OAI21_X1 U20367 ( .B1(n18634), .B2(n18234), .A(n18233), .ZN(P2_U2844) );
  INV_X1 U20368 ( .A(n18235), .ZN(n18239) );
  AOI22_X1 U20369 ( .A1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n18473), .B1(
        P2_REIP_REG_12__SCAN_IN), .B2(n18331), .ZN(n18236) );
  OAI211_X1 U20370 ( .C1(n18440), .C2(n18237), .A(n18236), .B(n18589), .ZN(
        n18238) );
  AOI21_X1 U20371 ( .B1(n18239), .B2(n18471), .A(n18238), .ZN(n18248) );
  INV_X1 U20372 ( .A(n18240), .ZN(n18256) );
  INV_X1 U20373 ( .A(n18241), .ZN(n18242) );
  NAND2_X1 U20374 ( .A1(n18243), .A2(n18242), .ZN(n18255) );
  NAND2_X1 U20375 ( .A1(n10964), .A2(n18255), .ZN(n18244) );
  XNOR2_X1 U20376 ( .A(n18256), .B(n18244), .ZN(n18245) );
  AOI22_X1 U20377 ( .A1(n18246), .A2(n18510), .B1(n18493), .B2(n18245), .ZN(
        n18247) );
  OAI211_X1 U20378 ( .C1(n18249), .C2(n18499), .A(n18248), .B(n18247), .ZN(
        P2_U2843) );
  NAND2_X1 U20379 ( .A1(n18250), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n18251) );
  OAI211_X1 U20380 ( .C1(n16391), .C2(n18502), .A(n18251), .B(n18589), .ZN(
        n18252) );
  AOI21_X1 U20381 ( .B1(n18253), .B2(n18471), .A(n18252), .ZN(n18264) );
  INV_X1 U20382 ( .A(n18254), .ZN(n18271) );
  NOR2_X1 U20383 ( .A1(n18256), .A2(n18255), .ZN(n18272) );
  NOR2_X1 U20384 ( .A1(n16641), .A2(n18272), .ZN(n18257) );
  XNOR2_X1 U20385 ( .A(n18271), .B(n18257), .ZN(n18262) );
  OAI22_X1 U20386 ( .A1(n18259), .A2(n18499), .B1(n18258), .B2(n18453), .ZN(
        n18260) );
  AOI21_X1 U20387 ( .B1(n18262), .B2(n18261), .A(n18260), .ZN(n18263) );
  OAI211_X1 U20388 ( .C1(n18265), .C2(n18486), .A(n18264), .B(n18263), .ZN(
        P2_U2842) );
  INV_X1 U20389 ( .A(P2_EBX_REG_14__SCAN_IN), .ZN(n18267) );
  AOI22_X1 U20390 ( .A1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n18473), .B1(
        P2_REIP_REG_14__SCAN_IN), .B2(n18331), .ZN(n18266) );
  OAI211_X1 U20391 ( .C1(n18440), .C2(n18267), .A(n18266), .B(n18589), .ZN(
        n18268) );
  AOI21_X1 U20392 ( .B1(n18269), .B2(n18457), .A(n18268), .ZN(n18276) );
  INV_X1 U20393 ( .A(n18270), .ZN(n18278) );
  NAND2_X1 U20394 ( .A1(n18272), .A2(n18271), .ZN(n18277) );
  NAND2_X1 U20395 ( .A1(n10964), .A2(n18277), .ZN(n18273) );
  XNOR2_X1 U20396 ( .A(n18278), .B(n18273), .ZN(n18274) );
  AOI22_X1 U20397 ( .A1(n18538), .A2(n18510), .B1(n18493), .B2(n18274), .ZN(
        n18275) );
  OAI211_X1 U20398 ( .C1(n18540), .C2(n18499), .A(n18276), .B(n18275), .ZN(
        P2_U2841) );
  NOR2_X1 U20399 ( .A1(n18278), .A2(n18277), .ZN(n18296) );
  NOR2_X1 U20400 ( .A1(n16641), .A2(n18296), .ZN(n18279) );
  XNOR2_X1 U20401 ( .A(n18294), .B(n18279), .ZN(n18289) );
  OAI21_X1 U20402 ( .B1(n18440), .B2(n18280), .A(n18589), .ZN(n18284) );
  OAI22_X1 U20403 ( .A1(n18282), .A2(n18486), .B1(n18281), .B2(n18504), .ZN(
        n18283) );
  AOI211_X1 U20404 ( .C1(P2_REIP_REG_15__SCAN_IN), .C2(n18331), .A(n18284), 
        .B(n18283), .ZN(n18288) );
  AOI22_X1 U20405 ( .A1(n18286), .A2(n18509), .B1(n18285), .B2(n18510), .ZN(
        n18287) );
  OAI211_X1 U20406 ( .C1(n18634), .C2(n18289), .A(n18288), .B(n18287), .ZN(
        P2_U2840) );
  AOI22_X1 U20407 ( .A1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n18473), .B1(
        P2_REIP_REG_16__SCAN_IN), .B2(n18331), .ZN(n18290) );
  OAI211_X1 U20408 ( .C1(n18440), .C2(n18291), .A(n18290), .B(n18589), .ZN(
        n18292) );
  AOI21_X1 U20409 ( .B1(n18293), .B2(n18471), .A(n18292), .ZN(n18300) );
  INV_X1 U20410 ( .A(n18294), .ZN(n18295) );
  NAND2_X1 U20411 ( .A1(n18296), .A2(n18295), .ZN(n18302) );
  NAND2_X1 U20412 ( .A1(n10964), .A2(n18302), .ZN(n18297) );
  XNOR2_X1 U20413 ( .A(n18303), .B(n18297), .ZN(n18298) );
  AOI22_X1 U20414 ( .A1(n19656), .A2(n18510), .B1(n18493), .B2(n18298), .ZN(
        n18299) );
  OAI211_X1 U20415 ( .C1(n18301), .C2(n18499), .A(n18300), .B(n18299), .ZN(
        P2_U2839) );
  NOR2_X1 U20416 ( .A1(n18303), .A2(n18302), .ZN(n18315) );
  NOR2_X1 U20417 ( .A1(n16641), .A2(n18315), .ZN(n18304) );
  XNOR2_X1 U20418 ( .A(n18305), .B(n18304), .ZN(n18313) );
  INV_X1 U20419 ( .A(n18306), .ZN(n18310) );
  INV_X1 U20420 ( .A(P2_EBX_REG_17__SCAN_IN), .ZN(n18308) );
  AOI22_X1 U20421 ( .A1(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n18473), .B1(
        P2_REIP_REG_17__SCAN_IN), .B2(n18331), .ZN(n18307) );
  OAI211_X1 U20422 ( .C1(n18440), .C2(n18308), .A(n18307), .B(n18589), .ZN(
        n18309) );
  AOI21_X1 U20423 ( .B1(n18310), .B2(n18471), .A(n18309), .ZN(n18312) );
  AOI22_X1 U20424 ( .A1(n18554), .A2(n18509), .B1(n18553), .B2(n18510), .ZN(
        n18311) );
  OAI211_X1 U20425 ( .C1(n18634), .C2(n18313), .A(n18312), .B(n18311), .ZN(
        P2_U2838) );
  NAND2_X1 U20426 ( .A1(n18315), .A2(n18314), .ZN(n18327) );
  NAND2_X1 U20427 ( .A1(n10964), .A2(n18327), .ZN(n18316) );
  XNOR2_X1 U20428 ( .A(n18326), .B(n18316), .ZN(n18325) );
  INV_X1 U20429 ( .A(P2_EBX_REG_18__SCAN_IN), .ZN(n18318) );
  AOI22_X1 U20430 ( .A1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n18473), .B1(
        P2_REIP_REG_18__SCAN_IN), .B2(n18331), .ZN(n18317) );
  OAI211_X1 U20431 ( .C1(n18440), .C2(n18318), .A(n18317), .B(n18589), .ZN(
        n18319) );
  AOI21_X1 U20432 ( .B1(n18320), .B2(n18471), .A(n18319), .ZN(n18324) );
  INV_X1 U20433 ( .A(n18321), .ZN(n18322) );
  AOI22_X1 U20434 ( .A1(n18322), .A2(n18509), .B1(n19547), .B2(n18510), .ZN(
        n18323) );
  OAI211_X1 U20435 ( .C1(n18634), .C2(n18325), .A(n18324), .B(n18323), .ZN(
        P2_U2837) );
  INV_X1 U20436 ( .A(n18326), .ZN(n18328) );
  NOR2_X1 U20437 ( .A1(n18328), .A2(n18327), .ZN(n18344) );
  NOR2_X1 U20438 ( .A1(n16641), .A2(n18344), .ZN(n18329) );
  XNOR2_X1 U20439 ( .A(n18342), .B(n18329), .ZN(n18340) );
  INV_X1 U20440 ( .A(n18330), .ZN(n18335) );
  AOI22_X1 U20441 ( .A1(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n18473), .B1(
        P2_REIP_REG_19__SCAN_IN), .B2(n18331), .ZN(n18332) );
  OAI211_X1 U20442 ( .C1(n18440), .C2(n18333), .A(n18332), .B(n18589), .ZN(
        n18334) );
  AOI21_X1 U20443 ( .B1(n18335), .B2(n18457), .A(n18334), .ZN(n18339) );
  AOI22_X1 U20444 ( .A1(n18337), .A2(n18509), .B1(n18336), .B2(n18510), .ZN(
        n18338) );
  OAI211_X1 U20445 ( .C1(n18634), .C2(n18340), .A(n18339), .B(n18338), .ZN(
        P2_U2836) );
  INV_X1 U20446 ( .A(n18341), .ZN(n18348) );
  INV_X1 U20447 ( .A(n18342), .ZN(n18343) );
  NAND2_X1 U20448 ( .A1(n18344), .A2(n18343), .ZN(n18345) );
  OAI21_X1 U20449 ( .B1(n18348), .B2(n18345), .A(n18403), .ZN(n18366) );
  AOI21_X1 U20450 ( .B1(n18348), .B2(n18345), .A(n18366), .ZN(n18346) );
  AOI22_X1 U20451 ( .A1(n18348), .A2(n18347), .B1(n18493), .B2(n18346), .ZN(
        n18357) );
  AOI22_X1 U20452 ( .A1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n18473), .B1(
        n18349), .B2(n18471), .ZN(n18356) );
  OAI22_X1 U20453 ( .A1(n18440), .A2(n18351), .B1(n18502), .B2(n18350), .ZN(
        n18352) );
  INV_X1 U20454 ( .A(n18352), .ZN(n18355) );
  AOI22_X1 U20455 ( .A1(n18353), .A2(n18509), .B1(n19455), .B2(n18510), .ZN(
        n18354) );
  NAND4_X1 U20456 ( .A1(n18357), .A2(n18356), .A3(n18355), .A4(n18354), .ZN(
        P2_U2835) );
  OAI22_X1 U20457 ( .A1(n18440), .A2(n18359), .B1(n18502), .B2(n18358), .ZN(
        n18360) );
  INV_X1 U20458 ( .A(n18360), .ZN(n18370) );
  AOI22_X1 U20459 ( .A1(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n18507), .B1(
        n18361), .B2(n18457), .ZN(n18369) );
  AOI22_X1 U20460 ( .A1(n18363), .A2(n18509), .B1(n18362), .B2(n18510), .ZN(
        n18368) );
  INV_X1 U20461 ( .A(n18364), .ZN(n18365) );
  NAND2_X1 U20462 ( .A1(n18365), .A2(n18366), .ZN(n18376) );
  OAI211_X1 U20463 ( .C1(n18366), .C2(n18365), .A(n18493), .B(n18376), .ZN(
        n18367) );
  NAND4_X1 U20464 ( .A1(n18370), .A2(n18369), .A3(n18368), .A4(n18367), .ZN(
        P2_U2834) );
  INV_X1 U20465 ( .A(P2_EBX_REG_22__SCAN_IN), .ZN(n18372) );
  OAI22_X1 U20466 ( .A1(n18440), .A2(n18372), .B1(n18502), .B2(n18371), .ZN(
        n18373) );
  INV_X1 U20467 ( .A(n18373), .ZN(n18382) );
  AOI22_X1 U20468 ( .A1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n18507), .B1(
        n18374), .B2(n18457), .ZN(n18381) );
  AOI22_X1 U20469 ( .A1(n18375), .A2(n18509), .B1(n19351), .B2(n18510), .ZN(
        n18380) );
  NAND2_X1 U20470 ( .A1(n10964), .A2(n18376), .ZN(n18378) );
  NAND2_X1 U20471 ( .A1(n18377), .A2(n18378), .ZN(n18390) );
  OAI211_X1 U20472 ( .C1(n18378), .C2(n18377), .A(n18493), .B(n18390), .ZN(
        n18379) );
  NAND4_X1 U20473 ( .A1(n18382), .A2(n18381), .A3(n18380), .A4(n18379), .ZN(
        P2_U2833) );
  INV_X1 U20474 ( .A(P2_EBX_REG_23__SCAN_IN), .ZN(n18384) );
  OAI22_X1 U20475 ( .A1(n18440), .A2(n18384), .B1(n18502), .B2(n18383), .ZN(
        n18388) );
  INV_X1 U20476 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n18386) );
  OAI22_X1 U20477 ( .A1(n18386), .A2(n18486), .B1(n18385), .B2(n18504), .ZN(
        n18387) );
  AOI211_X1 U20478 ( .C1(n18389), .C2(n18509), .A(n18388), .B(n18387), .ZN(
        n18394) );
  NAND2_X1 U20479 ( .A1(n10964), .A2(n18390), .ZN(n18392) );
  NAND2_X1 U20480 ( .A1(n18391), .A2(n18392), .ZN(n18402) );
  OAI211_X1 U20481 ( .C1(n18392), .C2(n18391), .A(n18493), .B(n18402), .ZN(
        n18393) );
  OAI211_X1 U20482 ( .C1(n18453), .C2(n18395), .A(n18394), .B(n18393), .ZN(
        P2_U2832) );
  INV_X1 U20483 ( .A(P2_EBX_REG_24__SCAN_IN), .ZN(n18397) );
  OAI22_X1 U20484 ( .A1(n18440), .A2(n18397), .B1(n18502), .B2(n18396), .ZN(
        n18398) );
  INV_X1 U20485 ( .A(n18398), .ZN(n18409) );
  AOI22_X1 U20486 ( .A1(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n18473), .B1(
        n18399), .B2(n18471), .ZN(n18408) );
  AOI22_X1 U20487 ( .A1(n18401), .A2(n18509), .B1(n18400), .B2(n18510), .ZN(
        n18407) );
  NAND2_X1 U20488 ( .A1(n10964), .A2(n18402), .ZN(n18405) );
  NAND2_X1 U20489 ( .A1(n18404), .A2(n18405), .ZN(n18417) );
  OAI211_X1 U20490 ( .C1(n18405), .C2(n18404), .A(n18493), .B(n18417), .ZN(
        n18406) );
  NAND4_X1 U20491 ( .A1(n18409), .A2(n18408), .A3(n18407), .A4(n18406), .ZN(
        P2_U2831) );
  OAI22_X1 U20492 ( .A1(n18440), .A2(n18411), .B1(n18502), .B2(n18410), .ZN(
        n18412) );
  INV_X1 U20493 ( .A(n18412), .ZN(n18424) );
  AOI22_X1 U20494 ( .A1(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n18473), .B1(
        n18413), .B2(n18457), .ZN(n18423) );
  INV_X1 U20495 ( .A(n18414), .ZN(n18415) );
  AOI22_X1 U20496 ( .A1(n18416), .A2(n18509), .B1(n18415), .B2(n18510), .ZN(
        n18422) );
  NAND2_X1 U20497 ( .A1(n10964), .A2(n18417), .ZN(n18420) );
  INV_X1 U20498 ( .A(n18418), .ZN(n18419) );
  NAND2_X1 U20499 ( .A1(n18419), .A2(n18420), .ZN(n18431) );
  OAI211_X1 U20500 ( .C1(n18420), .C2(n18419), .A(n18493), .B(n18431), .ZN(
        n18421) );
  NAND4_X1 U20501 ( .A1(n18424), .A2(n18423), .A3(n18422), .A4(n18421), .ZN(
        P2_U2830) );
  OAI22_X1 U20502 ( .A1(n18440), .A2(n18426), .B1(n18502), .B2(n18425), .ZN(
        n18427) );
  INV_X1 U20503 ( .A(n18427), .ZN(n18437) );
  AOI22_X1 U20504 ( .A1(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n18507), .B1(
        n18428), .B2(n18471), .ZN(n18436) );
  AOI22_X1 U20505 ( .A1(n18430), .A2(n18509), .B1(n18429), .B2(n18510), .ZN(
        n18435) );
  NAND2_X1 U20506 ( .A1(n10964), .A2(n18431), .ZN(n18433) );
  NAND2_X1 U20507 ( .A1(n18432), .A2(n18433), .ZN(n18446) );
  OAI211_X1 U20508 ( .C1(n18433), .C2(n18432), .A(n18493), .B(n18446), .ZN(
        n18434) );
  NAND4_X1 U20509 ( .A1(n18437), .A2(n18436), .A3(n18435), .A4(n18434), .ZN(
        P2_U2829) );
  INV_X1 U20510 ( .A(P2_EBX_REG_27__SCAN_IN), .ZN(n18439) );
  OAI22_X1 U20511 ( .A1(n18440), .A2(n18439), .B1(n18502), .B2(n18438), .ZN(
        n18444) );
  OAI22_X1 U20512 ( .A1(n18442), .A2(n18486), .B1(n18441), .B2(n18504), .ZN(
        n18443) );
  AOI211_X1 U20513 ( .C1(n18445), .C2(n18509), .A(n18444), .B(n18443), .ZN(
        n18451) );
  NAND2_X1 U20514 ( .A1(n10964), .A2(n18446), .ZN(n18449) );
  INV_X1 U20515 ( .A(n18447), .ZN(n18448) );
  NAND2_X1 U20516 ( .A1(n18448), .A2(n18449), .ZN(n18461) );
  OAI211_X1 U20517 ( .C1(n18449), .C2(n18448), .A(n18493), .B(n18461), .ZN(
        n18450) );
  OAI211_X1 U20518 ( .C1(n18453), .C2(n18452), .A(n18451), .B(n18450), .ZN(
        P2_U2828) );
  INV_X1 U20519 ( .A(P2_EBX_REG_28__SCAN_IN), .ZN(n18455) );
  OAI22_X1 U20520 ( .A1(n18440), .A2(n18455), .B1(n18502), .B2(n18454), .ZN(
        n18456) );
  INV_X1 U20521 ( .A(n18456), .ZN(n18467) );
  AOI22_X1 U20522 ( .A1(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n18507), .B1(
        n18458), .B2(n18457), .ZN(n18466) );
  AOI22_X1 U20523 ( .A1(n18460), .A2(n18509), .B1(n18459), .B2(n18510), .ZN(
        n18465) );
  NAND2_X1 U20524 ( .A1(n10964), .A2(n18461), .ZN(n18463) );
  NAND2_X1 U20525 ( .A1(n18462), .A2(n18463), .ZN(n18477) );
  OAI211_X1 U20526 ( .C1(n18463), .C2(n18462), .A(n18493), .B(n18477), .ZN(
        n18464) );
  NAND4_X1 U20527 ( .A1(n18467), .A2(n18466), .A3(n18465), .A4(n18464), .ZN(
        P2_U2827) );
  OAI22_X1 U20528 ( .A1(n18440), .A2(n18469), .B1(n18502), .B2(n18468), .ZN(
        n18470) );
  INV_X1 U20529 ( .A(n18470), .ZN(n18484) );
  AOI22_X1 U20530 ( .A1(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n18473), .B1(
        n18472), .B2(n18471), .ZN(n18483) );
  INV_X1 U20531 ( .A(n18474), .ZN(n18476) );
  AOI22_X1 U20532 ( .A1(n18476), .A2(n18509), .B1(n18475), .B2(n18510), .ZN(
        n18482) );
  NAND2_X1 U20533 ( .A1(n10964), .A2(n18477), .ZN(n18480) );
  INV_X1 U20534 ( .A(n18478), .ZN(n18479) );
  NAND2_X1 U20535 ( .A1(n18479), .A2(n18480), .ZN(n18492) );
  OAI211_X1 U20536 ( .C1(n18480), .C2(n18479), .A(n18493), .B(n18492), .ZN(
        n18481) );
  NAND4_X1 U20537 ( .A1(n18484), .A2(n18483), .A3(n18482), .A4(n18481), .ZN(
        P2_U2826) );
  OAI22_X1 U20538 ( .A1(n18440), .A2(n15414), .B1(n18502), .B2(n18485), .ZN(
        n18490) );
  INV_X1 U20539 ( .A(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n18487) );
  OAI22_X1 U20540 ( .A1(n18488), .A2(n18504), .B1(n18487), .B2(n18486), .ZN(
        n18489) );
  AOI211_X1 U20541 ( .C1(n18491), .C2(n18510), .A(n18490), .B(n18489), .ZN(
        n18497) );
  NAND2_X1 U20542 ( .A1(n10964), .A2(n18492), .ZN(n18495) );
  NAND2_X1 U20543 ( .A1(n18494), .A2(n18495), .ZN(n18514) );
  OAI211_X1 U20544 ( .C1(n18495), .C2(n18494), .A(n18493), .B(n18514), .ZN(
        n18496) );
  OAI211_X1 U20545 ( .C1(n18499), .C2(n18498), .A(n18497), .B(n18496), .ZN(
        P2_U2825) );
  INV_X1 U20546 ( .A(n18500), .ZN(n18503) );
  OAI222_X1 U20547 ( .A1(n18440), .A2(n18505), .B1(n18504), .B2(n18503), .C1(
        n18502), .C2(n18501), .ZN(n18506) );
  AOI21_X1 U20548 ( .B1(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n18507), .A(
        n18506), .ZN(n18512) );
  AOI22_X1 U20549 ( .A1(n18510), .A2(n19113), .B1(n18509), .B2(n18508), .ZN(
        n18511) );
  OAI211_X1 U20550 ( .C1(n18514), .C2(n18513), .A(n18512), .B(n18511), .ZN(
        P2_U2824) );
  AOI22_X1 U20551 ( .A1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n18516), .B1(
        n18568), .B2(n18515), .ZN(n18523) );
  OAI22_X1 U20552 ( .A1(n18594), .A2(n18518), .B1(n18517), .B2(n18606), .ZN(
        n18519) );
  AOI211_X1 U20553 ( .C1(n18591), .C2(n18521), .A(n18520), .B(n18519), .ZN(
        n18522) );
  OAI211_X1 U20554 ( .C1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(n18524), .A(
        n18523), .B(n18522), .ZN(P2_U3046) );
  OR2_X1 U20555 ( .A1(n18525), .A2(n18606), .ZN(n18534) );
  AOI22_X1 U20556 ( .A1(n18527), .A2(n18622), .B1(n18591), .B2(n18526), .ZN(
        n18533) );
  AOI21_X1 U20557 ( .B1(n18537), .B2(n18528), .A(n18613), .ZN(n18529) );
  NAND2_X1 U20558 ( .A1(n18555), .A2(n18529), .ZN(n18532) );
  NAND2_X1 U20559 ( .A1(n18568), .A2(n18530), .ZN(n18531) );
  AND4_X1 U20560 ( .A1(n18534), .A2(n18533), .A3(n18532), .A4(n18531), .ZN(
        n18536) );
  OAI211_X1 U20561 ( .C1(n18625), .C2(n18537), .A(n18536), .B(n18535), .ZN(
        P2_U3045) );
  AOI22_X1 U20562 ( .A1(n18622), .A2(n18538), .B1(P2_REIP_REG_14__SCAN_IN), 
        .B2(n18572), .ZN(n18552) );
  NAND2_X1 U20563 ( .A1(n18539), .A2(n18598), .ZN(n18542) );
  OR2_X1 U20564 ( .A1(n18540), .A2(n18605), .ZN(n18541) );
  OAI211_X1 U20565 ( .C1(n18543), .C2(n18617), .A(n18542), .B(n18541), .ZN(
        n18544) );
  INV_X1 U20566 ( .A(n18544), .ZN(n18551) );
  OAI21_X1 U20567 ( .B1(n18546), .B2(n18545), .A(
        P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n18550) );
  NAND3_X1 U20568 ( .A1(n18548), .A2(n15191), .A3(n18547), .ZN(n18549) );
  NAND4_X1 U20569 ( .A1(n18552), .A2(n18551), .A3(n18550), .A4(n18549), .ZN(
        P2_U3032) );
  AOI22_X1 U20570 ( .A1(n18554), .A2(n18591), .B1(n18622), .B2(n18553), .ZN(
        n18565) );
  NOR2_X1 U20571 ( .A1(n18555), .A2(n18568), .ZN(n18557) );
  OAI21_X1 U20572 ( .B1(n18558), .B2(n18557), .A(n18556), .ZN(n18560) );
  AOI22_X1 U20573 ( .A1(n18560), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .B1(
        n18559), .B2(n18598), .ZN(n18564) );
  OR3_X1 U20574 ( .A1(n18561), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A3(
        n15174), .ZN(n18562) );
  NAND4_X1 U20575 ( .A1(n18565), .A2(n18564), .A3(n18563), .A4(n18562), .ZN(
        P2_U3029) );
  AOI22_X1 U20576 ( .A1(n18567), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .B1(
        n18622), .B2(n18566), .ZN(n18578) );
  AOI222_X1 U20577 ( .A1(n18571), .A2(n18598), .B1(n18591), .B2(n18570), .C1(
        n18569), .C2(n18568), .ZN(n18577) );
  NAND2_X1 U20578 ( .A1(P2_REIP_REG_8__SCAN_IN), .A2(n18572), .ZN(n18576) );
  NAND2_X1 U20579 ( .A1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n18573) );
  OAI211_X1 U20580 ( .C1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(n18574), .B(n18573), .ZN(n18575) );
  NAND4_X1 U20581 ( .A1(n18578), .A2(n18577), .A3(n18576), .A4(n18575), .ZN(
        P2_U3038) );
  AOI22_X1 U20582 ( .A1(n18580), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B1(
        n18622), .B2(n18579), .ZN(n18588) );
  OAI22_X1 U20583 ( .A1(n18582), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B1(
        n18581), .B2(n18605), .ZN(n18586) );
  OAI22_X1 U20584 ( .A1(n18584), .A2(n18606), .B1(n18583), .B2(n18617), .ZN(
        n18585) );
  NOR2_X1 U20585 ( .A1(n18586), .A2(n18585), .ZN(n18587) );
  OAI211_X1 U20586 ( .C1(n13825), .C2(n18589), .A(n18588), .B(n18587), .ZN(
        P2_U3042) );
  NOR2_X1 U20587 ( .A1(n18590), .A2(n18617), .ZN(n18597) );
  NAND2_X1 U20588 ( .A1(n14864), .A2(n18591), .ZN(n18592) );
  OAI211_X1 U20589 ( .C1(n18595), .C2(n18594), .A(n18593), .B(n18592), .ZN(
        n18596) );
  AOI211_X1 U20590 ( .C1(n18599), .C2(n18598), .A(n18597), .B(n18596), .ZN(
        n18600) );
  OAI221_X1 U20591 ( .B1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n18603), .C1(
        n18602), .C2(n18601), .A(n18600), .ZN(P2_U3043) );
  NAND2_X1 U20592 ( .A1(n18614), .A2(n18604), .ZN(n18624) );
  OAI22_X1 U20593 ( .A1(n18607), .A2(n18606), .B1(n18605), .B2(n14807), .ZN(
        n18620) );
  AOI21_X1 U20594 ( .B1(n18610), .B2(n18609), .A(n18608), .ZN(n18612) );
  NOR2_X1 U20595 ( .A1(n18612), .A2(n18611), .ZN(n18616) );
  NAND3_X1 U20596 ( .A1(n18614), .A2(n18626), .A3(n18613), .ZN(n18615) );
  OAI211_X1 U20597 ( .C1(n18618), .C2(n18617), .A(n18616), .B(n18615), .ZN(
        n18619) );
  AOI211_X1 U20598 ( .C1(n18622), .C2(n18621), .A(n18620), .B(n18619), .ZN(
        n18623) );
  OAI221_X1 U20599 ( .B1(n18626), .B2(n18625), .C1(n18626), .C2(n18624), .A(
        n18623), .ZN(P2_U3044) );
  NAND2_X1 U20600 ( .A1(n18641), .A2(n18627), .ZN(n18643) );
  OAI21_X1 U20601 ( .B1(n18629), .B2(n18628), .A(n18649), .ZN(n18633) );
  NAND2_X1 U20602 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(n18630), .ZN(n18631) );
  AOI21_X1 U20603 ( .B1(n18636), .B2(n18643), .A(n18631), .ZN(n18632) );
  AOI21_X1 U20604 ( .B1(n18643), .B2(n18633), .A(n18632), .ZN(n18635) );
  NAND2_X1 U20605 ( .A1(n18635), .A2(n18634), .ZN(P2_U3177) );
  OAI22_X1 U20606 ( .A1(n18638), .A2(n18637), .B1(n21729), .B2(n18636), .ZN(
        n18639) );
  AOI211_X1 U20607 ( .C1(n18641), .C2(P2_STATE2_REG_0__SCAN_IN), .A(n18640), 
        .B(n18639), .ZN(n18647) );
  NOR2_X1 U20608 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n18642), .ZN(n18645) );
  OAI22_X1 U20609 ( .A1(n18645), .A2(n18644), .B1(n21729), .B2(n18643), .ZN(
        n18646) );
  OAI211_X1 U20610 ( .C1(n18648), .C2(n18649), .A(n18647), .B(n18646), .ZN(
        P2_U3176) );
  OR2_X1 U20611 ( .A1(n18650), .A2(n18649), .ZN(n18654) );
  NAND2_X1 U20612 ( .A1(n18654), .A2(P2_MORE_REG_SCAN_IN), .ZN(n18651) );
  OAI21_X1 U20613 ( .B1(n18654), .B2(n18652), .A(n18651), .ZN(P2_U3609) );
  AOI21_X1 U20614 ( .B1(n18654), .B2(P2_FLUSH_REG_SCAN_IN), .A(n18653), .ZN(
        n18655) );
  INV_X1 U20615 ( .A(n18655), .ZN(P2_U2819) );
  INV_X1 U20616 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n20101) );
  INV_X1 U20617 ( .A(BUF2_REG_31__SCAN_IN), .ZN(n18682) );
  AOI22_X1 U20618 ( .A1(n19008), .A2(n20101), .B1(n18682), .B2(U215), .ZN(U282) );
  OAI22_X1 U20619 ( .A1(U215), .A2(P2_DATAO_REG_30__SCAN_IN), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n19008), .ZN(n18656) );
  INV_X1 U20620 ( .A(n18656), .ZN(U281) );
  INV_X1 U20621 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n18658) );
  AOI22_X1 U20622 ( .A1(n19008), .A2(n18658), .B1(n18657), .B2(U215), .ZN(U280) );
  OAI22_X1 U20623 ( .A1(U215), .A2(P2_DATAO_REG_28__SCAN_IN), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n18966), .ZN(n18659) );
  INV_X1 U20624 ( .A(n18659), .ZN(U279) );
  INV_X1 U20625 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n18661) );
  AOI22_X1 U20626 ( .A1(n19008), .A2(n18661), .B1(n18660), .B2(U215), .ZN(U278) );
  OAI22_X1 U20627 ( .A1(U215), .A2(P2_DATAO_REG_26__SCAN_IN), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n18966), .ZN(n18662) );
  INV_X1 U20628 ( .A(n18662), .ZN(U277) );
  OAI22_X1 U20629 ( .A1(U215), .A2(P2_DATAO_REG_25__SCAN_IN), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n19008), .ZN(n18663) );
  INV_X1 U20630 ( .A(n18663), .ZN(U276) );
  INV_X1 U20631 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n18664) );
  AOI22_X1 U20632 ( .A1(n19008), .A2(n18664), .B1(n16212), .B2(U215), .ZN(U275) );
  INV_X1 U20633 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n18665) );
  AOI22_X1 U20634 ( .A1(n19008), .A2(n18665), .B1(n16219), .B2(U215), .ZN(U274) );
  INV_X1 U20635 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n18666) );
  INV_X1 U20636 ( .A(BUF2_REG_22__SCAN_IN), .ZN(n19359) );
  AOI22_X1 U20637 ( .A1(n19008), .A2(n18666), .B1(n19359), .B2(U215), .ZN(U273) );
  INV_X1 U20638 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n18667) );
  AOI22_X1 U20639 ( .A1(n18966), .A2(n18667), .B1(n16232), .B2(U215), .ZN(U272) );
  OAI22_X1 U20640 ( .A1(U215), .A2(P2_DATAO_REG_20__SCAN_IN), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n19008), .ZN(n18668) );
  INV_X1 U20641 ( .A(n18668), .ZN(U271) );
  OAI22_X1 U20642 ( .A1(U215), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n19008), .ZN(n18669) );
  INV_X1 U20643 ( .A(n18669), .ZN(U270) );
  OAI22_X1 U20644 ( .A1(U215), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n19008), .ZN(n18670) );
  INV_X1 U20645 ( .A(n18670), .ZN(U269) );
  INV_X1 U20646 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n18671) );
  INV_X1 U20647 ( .A(BUF2_REG_17__SCAN_IN), .ZN(n19606) );
  AOI22_X1 U20648 ( .A1(n18966), .A2(n18671), .B1(n19606), .B2(U215), .ZN(U268) );
  INV_X1 U20649 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n18672) );
  INV_X1 U20650 ( .A(BUF2_REG_16__SCAN_IN), .ZN(n19680) );
  AOI22_X1 U20651 ( .A1(n19008), .A2(n18672), .B1(n19680), .B2(U215), .ZN(U267) );
  OAI22_X1 U20652 ( .A1(U215), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n19008), .ZN(n18673) );
  INV_X1 U20653 ( .A(n18673), .ZN(U266) );
  OAI22_X1 U20654 ( .A1(U215), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n19008), .ZN(n18674) );
  INV_X1 U20655 ( .A(n18674), .ZN(U265) );
  OAI22_X1 U20656 ( .A1(U215), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(
        BUF2_REG_13__SCAN_IN), .B2(n19008), .ZN(n18675) );
  INV_X1 U20657 ( .A(n18675), .ZN(U264) );
  INV_X1 U20658 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n18676) );
  INV_X1 U20659 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n20624) );
  AOI22_X1 U20660 ( .A1(n18966), .A2(n18676), .B1(n20624), .B2(U215), .ZN(U263) );
  OAI22_X1 U20661 ( .A1(U215), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(
        BUF2_REG_11__SCAN_IN), .B2(n19008), .ZN(n18677) );
  INV_X1 U20662 ( .A(n18677), .ZN(U262) );
  INV_X1 U20663 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n18678) );
  INV_X1 U20664 ( .A(BUF2_REG_10__SCAN_IN), .ZN(n20718) );
  AOI22_X1 U20665 ( .A1(n19008), .A2(n18678), .B1(n20718), .B2(U215), .ZN(U261) );
  INV_X1 U20666 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n18679) );
  INV_X1 U20667 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n20637) );
  AOI22_X1 U20668 ( .A1(n19008), .A2(n18679), .B1(n20637), .B2(U215), .ZN(U260) );
  OAI22_X1 U20669 ( .A1(U215), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n18966), .ZN(n18680) );
  INV_X1 U20670 ( .A(n18680), .ZN(U259) );
  OAI22_X1 U20671 ( .A1(U215), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n18966), .ZN(n18681) );
  INV_X1 U20672 ( .A(n18681), .ZN(U258) );
  NOR3_X1 U20673 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18692), .A3(
        n21275), .ZN(n18683) );
  NAND2_X1 U20674 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18683), .ZN(
        n19112) );
  NAND2_X1 U20675 ( .A1(BUF2_REG_23__SCAN_IN), .A2(n18884), .ZN(n18755) );
  INV_X1 U20676 ( .A(n18683), .ZN(n18691) );
  NOR2_X2 U20677 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18691), .ZN(
        n19029) );
  NAND2_X1 U20678 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n21288), .ZN(n21289) );
  NOR2_X1 U20679 ( .A1(n21275), .A2(n18707), .ZN(n18751) );
  AND2_X1 U20680 ( .A1(n21289), .A2(n18751), .ZN(n19011) );
  AND2_X1 U20681 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n18968), .ZN(n18756) );
  AOI22_X1 U20682 ( .A1(n19029), .A2(n18757), .B1(n19011), .B2(n18756), .ZN(
        n18687) );
  AND2_X1 U20683 ( .A1(n18704), .A2(n18968), .ZN(n18693) );
  AOI22_X1 U20684 ( .A1(n18884), .A2(n18683), .B1(n18751), .B2(n18693), .ZN(
        n19014) );
  NAND2_X1 U20685 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18751), .ZN(
        n19094) );
  INV_X1 U20686 ( .A(n19094), .ZN(n19096) );
  NAND2_X1 U20687 ( .A1(n18685), .A2(n18684), .ZN(n19012) );
  NOR2_X2 U20688 ( .A1(n20687), .A2(n19012), .ZN(n18752) );
  AOI22_X1 U20689 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n19014), .B1(
        n19096), .B2(n18752), .ZN(n18686) );
  OAI211_X1 U20690 ( .C1(n19112), .C2(n18755), .A(n18687), .B(n18686), .ZN(
        P3_U2995) );
  INV_X1 U20691 ( .A(n18757), .ZN(n18720) );
  NOR2_X1 U20692 ( .A1(n21263), .A2(n18712), .ZN(n18701) );
  NAND2_X1 U20693 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18701), .ZN(
        n19021) );
  INV_X1 U20694 ( .A(n18755), .ZN(n18762) );
  INV_X1 U20695 ( .A(n21289), .ZN(n20162) );
  INV_X1 U20696 ( .A(n19112), .ZN(n19023) );
  NAND2_X1 U20697 ( .A1(n21262), .A2(n18751), .ZN(n19101) );
  INV_X1 U20698 ( .A(n19101), .ZN(n19105) );
  NOR2_X1 U20699 ( .A1(n19023), .A2(n19105), .ZN(n18758) );
  NOR2_X1 U20700 ( .A1(n20162), .A2(n18758), .ZN(n19017) );
  AOI22_X1 U20701 ( .A1(n18762), .A2(n19029), .B1(n18756), .B2(n19017), .ZN(
        n18690) );
  NOR2_X1 U20702 ( .A1(n19029), .A2(n19035), .ZN(n18697) );
  OAI22_X1 U20703 ( .A1(n18758), .A2(n19010), .B1(n18697), .B2(n19009), .ZN(
        n18688) );
  OAI21_X1 U20704 ( .B1(n19105), .B2(n21296), .A(n18688), .ZN(n19018) );
  AOI22_X1 U20705 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n19018), .B1(
        n18752), .B2(n19105), .ZN(n18689) );
  OAI211_X1 U20706 ( .C1(n18720), .C2(n19021), .A(n18690), .B(n18689), .ZN(
        P3_U2987) );
  NAND2_X1 U20707 ( .A1(n18701), .A2(n21262), .ZN(n19027) );
  NOR2_X1 U20708 ( .A1(n20162), .A2(n18691), .ZN(n19022) );
  AOI22_X1 U20709 ( .A1(n18762), .A2(n19035), .B1(n18756), .B2(n19022), .ZN(
        n18696) );
  NOR2_X1 U20710 ( .A1(n18692), .A2(n21275), .ZN(n18694) );
  AND2_X1 U20711 ( .A1(n18693), .A2(n21263), .ZN(n18750) );
  AOI22_X1 U20712 ( .A1(n18884), .A2(n18701), .B1(n18694), .B2(n18750), .ZN(
        n19024) );
  AOI22_X1 U20713 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n19024), .B1(
        n19023), .B2(n18752), .ZN(n18695) );
  OAI211_X1 U20714 ( .C1(n18720), .C2(n19027), .A(n18696), .B(n18695), .ZN(
        P3_U2979) );
  NOR2_X1 U20715 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n21262), .ZN(
        n18735) );
  NAND2_X1 U20716 ( .A1(n18713), .A2(n18735), .ZN(n19033) );
  NOR2_X1 U20717 ( .A1(n20162), .A2(n18697), .ZN(n19028) );
  AOI22_X1 U20718 ( .A1(n18762), .A2(n19041), .B1(n18756), .B2(n19028), .ZN(
        n18700) );
  NAND2_X1 U20719 ( .A1(n19027), .A2(n19033), .ZN(n18708) );
  AOI21_X1 U20720 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n19010), .ZN(n18760) );
  INV_X1 U20721 ( .A(n18697), .ZN(n18698) );
  AOI22_X1 U20722 ( .A1(n18884), .A2(n18708), .B1(n18760), .B2(n18698), .ZN(
        n19030) );
  AOI22_X1 U20723 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n19030), .B1(
        n18752), .B2(n19029), .ZN(n18699) );
  OAI211_X1 U20724 ( .C1(n18720), .C2(n19033), .A(n18700), .B(n18699), .ZN(
        P3_U2971) );
  NOR2_X1 U20725 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n21267) );
  NAND2_X1 U20726 ( .A1(n21267), .A2(n18713), .ZN(n19039) );
  INV_X1 U20727 ( .A(n18701), .ZN(n18702) );
  NOR2_X1 U20728 ( .A1(n20162), .A2(n18702), .ZN(n19034) );
  AOI22_X1 U20729 ( .A1(n18757), .A2(n19053), .B1(n18756), .B2(n19034), .ZN(
        n18706) );
  INV_X1 U20730 ( .A(n18703), .ZN(n18726) );
  AOI21_X1 U20731 ( .B1(n21263), .B2(n18726), .A(n19010), .ZN(n18722) );
  AND2_X1 U20732 ( .A1(n18704), .A2(n18722), .ZN(n18741) );
  NAND2_X1 U20733 ( .A1(n18713), .A2(n18741), .ZN(n19036) );
  AOI22_X1 U20734 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19036), .B1(
        n18752), .B2(n19035), .ZN(n18705) );
  OAI211_X1 U20735 ( .C1(n18755), .C2(n19033), .A(n18706), .B(n18705), .ZN(
        P3_U2963) );
  NOR2_X1 U20736 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18707), .ZN(
        n18721) );
  NAND2_X1 U20737 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18721), .ZN(
        n19045) );
  AND2_X1 U20738 ( .A1(n21289), .A2(n18708), .ZN(n19040) );
  AOI22_X1 U20739 ( .A1(n18762), .A2(n19053), .B1(n18756), .B2(n19040), .ZN(
        n18711) );
  NOR2_X1 U20740 ( .A1(n19053), .A2(n19059), .ZN(n18716) );
  OAI22_X1 U20741 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n19033), .B1(n18716), 
        .B2(n18726), .ZN(n18709) );
  OAI21_X1 U20742 ( .B1(n19041), .B2(n18709), .A(n18968), .ZN(n19042) );
  AOI22_X1 U20743 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19042), .B1(
        n18752), .B2(n19041), .ZN(n18710) );
  OAI211_X1 U20744 ( .C1(n18720), .C2(n19045), .A(n18711), .B(n18710), .ZN(
        P3_U2955) );
  NAND2_X1 U20745 ( .A1(n21262), .A2(n18721), .ZN(n19051) );
  INV_X1 U20746 ( .A(n19051), .ZN(n19065) );
  NAND2_X1 U20747 ( .A1(n21263), .A2(n21289), .ZN(n18748) );
  NOR2_X1 U20748 ( .A1(n18712), .A2(n18748), .ZN(n19046) );
  AOI22_X1 U20749 ( .A1(n18757), .A2(n19065), .B1(n18756), .B2(n19046), .ZN(
        n18715) );
  AOI22_X1 U20750 ( .A1(n18884), .A2(n18721), .B1(n18713), .B2(n18750), .ZN(
        n19048) );
  INV_X1 U20751 ( .A(n19033), .ZN(n19047) );
  AOI22_X1 U20752 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19048), .B1(
        n18752), .B2(n19047), .ZN(n18714) );
  OAI211_X1 U20753 ( .C1(n18755), .C2(n19045), .A(n18715), .B(n18714), .ZN(
        P3_U2947) );
  NAND2_X1 U20754 ( .A1(n18735), .A2(n18731), .ZN(n19057) );
  NOR2_X1 U20755 ( .A1(n20162), .A2(n18716), .ZN(n19052) );
  AOI22_X1 U20756 ( .A1(n18762), .A2(n19065), .B1(n18756), .B2(n19052), .ZN(
        n18719) );
  NAND2_X1 U20757 ( .A1(n19051), .A2(n19057), .ZN(n18725) );
  INV_X1 U20758 ( .A(n18716), .ZN(n18717) );
  AOI22_X1 U20759 ( .A1(n18884), .A2(n18725), .B1(n18760), .B2(n18717), .ZN(
        n19054) );
  AOI22_X1 U20760 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19054), .B1(
        n18752), .B2(n19053), .ZN(n18718) );
  OAI211_X1 U20761 ( .C1(n18720), .C2(n19057), .A(n18719), .B(n18718), .ZN(
        P3_U2939) );
  NAND2_X1 U20762 ( .A1(n21267), .A2(n18731), .ZN(n19063) );
  AND2_X1 U20763 ( .A1(n21289), .A2(n18721), .ZN(n19058) );
  AOI22_X1 U20764 ( .A1(n18757), .A2(n19076), .B1(n18756), .B2(n19058), .ZN(
        n18724) );
  OAI211_X1 U20765 ( .C1(n19059), .C2(n21296), .A(n18731), .B(n18722), .ZN(
        n19060) );
  AOI22_X1 U20766 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19060), .B1(
        n18752), .B2(n19059), .ZN(n18723) );
  OAI211_X1 U20767 ( .C1(n18755), .C2(n19057), .A(n18724), .B(n18723), .ZN(
        P3_U2931) );
  NOR2_X1 U20768 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18749) );
  NAND2_X1 U20769 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18749), .ZN(
        n18740) );
  NOR2_X2 U20770 ( .A1(n21262), .A2(n18740), .ZN(n19083) );
  AND2_X1 U20771 ( .A1(n21289), .A2(n18725), .ZN(n19064) );
  AOI22_X1 U20772 ( .A1(n18757), .A2(n19083), .B1(n18756), .B2(n19064), .ZN(
        n18729) );
  NOR2_X1 U20773 ( .A1(n19076), .A2(n19083), .ZN(n18736) );
  OAI22_X1 U20774 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n19057), .B1(n18736), 
        .B2(n18726), .ZN(n18727) );
  OAI21_X1 U20775 ( .B1(n19065), .B2(n18727), .A(n18968), .ZN(n19066) );
  AOI22_X1 U20776 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19066), .B1(
        n18752), .B2(n19065), .ZN(n18728) );
  OAI211_X1 U20777 ( .C1(n18755), .C2(n19063), .A(n18729), .B(n18728), .ZN(
        P3_U2923) );
  INV_X1 U20778 ( .A(n18752), .ZN(n18765) );
  NOR2_X2 U20779 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18740), .ZN(
        n19090) );
  INV_X1 U20780 ( .A(n18731), .ZN(n18730) );
  NOR2_X1 U20781 ( .A1(n18748), .A2(n18730), .ZN(n19070) );
  AOI22_X1 U20782 ( .A1(n18757), .A2(n19090), .B1(n18756), .B2(n19070), .ZN(
        n18734) );
  INV_X1 U20783 ( .A(n18740), .ZN(n18732) );
  AOI22_X1 U20784 ( .A1(n18884), .A2(n18732), .B1(n18750), .B2(n18731), .ZN(
        n19072) );
  AOI22_X1 U20785 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19072), .B1(
        n18762), .B2(n19083), .ZN(n18733) );
  OAI211_X1 U20786 ( .C1(n18765), .C2(n19057), .A(n18734), .B(n18733), .ZN(
        P3_U2915) );
  NAND2_X1 U20787 ( .A1(n18735), .A2(n18749), .ZN(n19088) );
  INV_X1 U20788 ( .A(n19088), .ZN(n19097) );
  NOR2_X1 U20789 ( .A1(n20162), .A2(n18736), .ZN(n19075) );
  AOI22_X1 U20790 ( .A1(n18757), .A2(n19097), .B1(n18756), .B2(n19075), .ZN(
        n18739) );
  NAND2_X1 U20791 ( .A1(n19080), .A2(n19088), .ZN(n18744) );
  INV_X1 U20792 ( .A(n18736), .ZN(n18737) );
  AOI22_X1 U20793 ( .A1(n18884), .A2(n18744), .B1(n18760), .B2(n18737), .ZN(
        n19077) );
  AOI22_X1 U20794 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19077), .B1(
        n18762), .B2(n19090), .ZN(n18738) );
  OAI211_X1 U20795 ( .C1(n18765), .C2(n19063), .A(n18739), .B(n18738), .ZN(
        P3_U2907) );
  NAND2_X1 U20796 ( .A1(n21267), .A2(n18749), .ZN(n18955) );
  INV_X1 U20797 ( .A(n18955), .ZN(n19107) );
  NOR2_X1 U20798 ( .A1(n20162), .A2(n18740), .ZN(n19082) );
  AOI22_X1 U20799 ( .A1(n18757), .A2(n19107), .B1(n18756), .B2(n19082), .ZN(
        n18743) );
  NAND2_X1 U20800 ( .A1(n18741), .A2(n18749), .ZN(n19084) );
  AOI22_X1 U20801 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19084), .B1(
        n18752), .B2(n19083), .ZN(n18742) );
  OAI211_X1 U20802 ( .C1(n18755), .C2(n19088), .A(n18743), .B(n18742), .ZN(
        P3_U2899) );
  AND2_X1 U20803 ( .A1(n21289), .A2(n18744), .ZN(n19089) );
  AOI22_X1 U20804 ( .A1(n19096), .A2(n18757), .B1(n18756), .B2(n19089), .ZN(
        n18746) );
  NAND2_X1 U20805 ( .A1(n19094), .A2(n18955), .ZN(n18759) );
  AOI22_X1 U20806 ( .A1(n18884), .A2(n18759), .B1(n18760), .B2(n18744), .ZN(
        n19091) );
  AOI22_X1 U20807 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19091), .B1(
        n18762), .B2(n19107), .ZN(n18745) );
  OAI211_X1 U20808 ( .C1(n18765), .C2(n19080), .A(n18746), .B(n18745), .ZN(
        P3_U2891) );
  INV_X1 U20809 ( .A(n18749), .ZN(n18747) );
  NOR2_X1 U20810 ( .A1(n18748), .A2(n18747), .ZN(n19095) );
  AOI22_X1 U20811 ( .A1(n18757), .A2(n19105), .B1(n18756), .B2(n19095), .ZN(
        n18754) );
  AOI22_X1 U20812 ( .A1(n18884), .A2(n18751), .B1(n18750), .B2(n18749), .ZN(
        n19098) );
  AOI22_X1 U20813 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19098), .B1(
        n18752), .B2(n19097), .ZN(n18753) );
  OAI211_X1 U20814 ( .C1(n18755), .C2(n19094), .A(n18754), .B(n18753), .ZN(
        P3_U2883) );
  AND2_X1 U20815 ( .A1(n21289), .A2(n18759), .ZN(n19103) );
  AOI22_X1 U20816 ( .A1(n19023), .A2(n18757), .B1(n18756), .B2(n19103), .ZN(
        n18764) );
  INV_X1 U20817 ( .A(n18758), .ZN(n18761) );
  AOI22_X1 U20818 ( .A1(n18884), .A2(n18761), .B1(n18760), .B2(n18759), .ZN(
        n19108) );
  AOI22_X1 U20819 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n19108), .B1(
        n18762), .B2(n19105), .ZN(n18763) );
  OAI211_X1 U20820 ( .C1(n18765), .C2(n18955), .A(n18764), .B(n18763), .ZN(
        P3_U2875) );
  INV_X1 U20821 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n18766) );
  AOI22_X1 U20822 ( .A1(n18966), .A2(n18766), .B1(n20145), .B2(U215), .ZN(U257) );
  OR2_X1 U20823 ( .A1(n19012), .A2(n20674), .ZN(n18802) );
  NOR2_X2 U20824 ( .A1(n19359), .A2(n19009), .ZN(n18798) );
  NOR2_X2 U20825 ( .A1(n20145), .A2(n19010), .ZN(n18797) );
  AOI22_X1 U20826 ( .A1(n19023), .A2(n18798), .B1(n19011), .B2(n18797), .ZN(
        n18768) );
  AND2_X1 U20827 ( .A1(BUF2_REG_30__SCAN_IN), .A2(n18884), .ZN(n18799) );
  AOI22_X1 U20828 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n19014), .B1(
        n19029), .B2(n18799), .ZN(n18767) );
  OAI211_X1 U20829 ( .C1(n19094), .C2(n18802), .A(n18768), .B(n18767), .ZN(
        P3_U2994) );
  AOI22_X1 U20830 ( .A1(n19035), .A2(n18799), .B1(n19017), .B2(n18797), .ZN(
        n18770) );
  AOI22_X1 U20831 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n19018), .B1(
        n19029), .B2(n18798), .ZN(n18769) );
  OAI211_X1 U20832 ( .C1(n19101), .C2(n18802), .A(n18770), .B(n18769), .ZN(
        P3_U2986) );
  AOI22_X1 U20833 ( .A1(n19035), .A2(n18798), .B1(n19022), .B2(n18797), .ZN(
        n18772) );
  AOI22_X1 U20834 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19024), .B1(
        n19041), .B2(n18799), .ZN(n18771) );
  OAI211_X1 U20835 ( .C1(n19112), .C2(n18802), .A(n18772), .B(n18771), .ZN(
        P3_U2978) );
  INV_X1 U20836 ( .A(n19029), .ZN(n18930) );
  AOI22_X1 U20837 ( .A1(n19047), .A2(n18799), .B1(n19028), .B2(n18797), .ZN(
        n18774) );
  AOI22_X1 U20838 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n19030), .B1(
        n19041), .B2(n18798), .ZN(n18773) );
  OAI211_X1 U20839 ( .C1(n18930), .C2(n18802), .A(n18774), .B(n18773), .ZN(
        P3_U2970) );
  AOI22_X1 U20840 ( .A1(n19047), .A2(n18798), .B1(n19034), .B2(n18797), .ZN(
        n18776) );
  AOI22_X1 U20841 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19036), .B1(
        n19053), .B2(n18799), .ZN(n18775) );
  OAI211_X1 U20842 ( .C1(n19021), .C2(n18802), .A(n18776), .B(n18775), .ZN(
        P3_U2962) );
  AOI22_X1 U20843 ( .A1(n19059), .A2(n18799), .B1(n19040), .B2(n18797), .ZN(
        n18778) );
  AOI22_X1 U20844 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19042), .B1(
        n19053), .B2(n18798), .ZN(n18777) );
  OAI211_X1 U20845 ( .C1(n19027), .C2(n18802), .A(n18778), .B(n18777), .ZN(
        P3_U2954) );
  AOI22_X1 U20846 ( .A1(n19065), .A2(n18799), .B1(n19046), .B2(n18797), .ZN(
        n18780) );
  AOI22_X1 U20847 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19048), .B1(
        n19059), .B2(n18798), .ZN(n18779) );
  OAI211_X1 U20848 ( .C1(n19033), .C2(n18802), .A(n18780), .B(n18779), .ZN(
        P3_U2946) );
  INV_X1 U20849 ( .A(n19057), .ZN(n19071) );
  AOI22_X1 U20850 ( .A1(n19071), .A2(n18799), .B1(n19052), .B2(n18797), .ZN(
        n18782) );
  AOI22_X1 U20851 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19054), .B1(
        n19065), .B2(n18798), .ZN(n18781) );
  OAI211_X1 U20852 ( .C1(n19039), .C2(n18802), .A(n18782), .B(n18781), .ZN(
        P3_U2938) );
  AOI22_X1 U20853 ( .A1(n19058), .A2(n18797), .B1(n19076), .B2(n18799), .ZN(
        n18784) );
  AOI22_X1 U20854 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19060), .B1(
        n19071), .B2(n18798), .ZN(n18783) );
  OAI211_X1 U20855 ( .C1(n19045), .C2(n18802), .A(n18784), .B(n18783), .ZN(
        P3_U2930) );
  AOI22_X1 U20856 ( .A1(n19076), .A2(n18798), .B1(n19064), .B2(n18797), .ZN(
        n18786) );
  AOI22_X1 U20857 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19066), .B1(
        n19083), .B2(n18799), .ZN(n18785) );
  OAI211_X1 U20858 ( .C1(n19051), .C2(n18802), .A(n18786), .B(n18785), .ZN(
        P3_U2922) );
  AOI22_X1 U20859 ( .A1(n19090), .A2(n18799), .B1(n19070), .B2(n18797), .ZN(
        n18788) );
  AOI22_X1 U20860 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19072), .B1(
        n19083), .B2(n18798), .ZN(n18787) );
  OAI211_X1 U20861 ( .C1(n19057), .C2(n18802), .A(n18788), .B(n18787), .ZN(
        P3_U2914) );
  AOI22_X1 U20862 ( .A1(n19097), .A2(n18799), .B1(n19075), .B2(n18797), .ZN(
        n18790) );
  AOI22_X1 U20863 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19077), .B1(
        n19090), .B2(n18798), .ZN(n18789) );
  OAI211_X1 U20864 ( .C1(n19063), .C2(n18802), .A(n18790), .B(n18789), .ZN(
        P3_U2906) );
  INV_X1 U20865 ( .A(n19083), .ZN(n19069) );
  AOI22_X1 U20866 ( .A1(n19097), .A2(n18798), .B1(n19082), .B2(n18797), .ZN(
        n18792) );
  AOI22_X1 U20867 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19084), .B1(
        n19107), .B2(n18799), .ZN(n18791) );
  OAI211_X1 U20868 ( .C1(n19069), .C2(n18802), .A(n18792), .B(n18791), .ZN(
        P3_U2898) );
  AOI22_X1 U20869 ( .A1(n19107), .A2(n18798), .B1(n19089), .B2(n18797), .ZN(
        n18794) );
  AOI22_X1 U20870 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19091), .B1(
        n19096), .B2(n18799), .ZN(n18793) );
  OAI211_X1 U20871 ( .C1(n19080), .C2(n18802), .A(n18794), .B(n18793), .ZN(
        P3_U2890) );
  AOI22_X1 U20872 ( .A1(n19096), .A2(n18798), .B1(n19095), .B2(n18797), .ZN(
        n18796) );
  AOI22_X1 U20873 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19098), .B1(
        n19105), .B2(n18799), .ZN(n18795) );
  OAI211_X1 U20874 ( .C1(n19088), .C2(n18802), .A(n18796), .B(n18795), .ZN(
        P3_U2882) );
  AOI22_X1 U20875 ( .A1(n19105), .A2(n18798), .B1(n19103), .B2(n18797), .ZN(
        n18801) );
  AOI22_X1 U20876 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n19108), .B1(
        n19023), .B2(n18799), .ZN(n18800) );
  OAI211_X1 U20877 ( .C1(n18955), .C2(n18802), .A(n18801), .B(n18800), .ZN(
        P3_U2874) );
  INV_X1 U20878 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n18803) );
  INV_X1 U20879 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n20649) );
  AOI22_X1 U20880 ( .A1(n19008), .A2(n18803), .B1(n20649), .B2(U215), .ZN(U256) );
  NAND2_X1 U20881 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n18884), .ZN(n18832) );
  NOR2_X1 U20882 ( .A1(n16232), .A2(n19009), .ZN(n18829) );
  NOR2_X2 U20883 ( .A1(n20649), .A2(n19010), .ZN(n18837) );
  AOI22_X1 U20884 ( .A1(n19023), .A2(n18829), .B1(n19011), .B2(n18837), .ZN(
        n18806) );
  NOR2_X2 U20885 ( .A1(n18804), .A2(n19012), .ZN(n18839) );
  AOI22_X1 U20886 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n19014), .B1(
        n19096), .B2(n18839), .ZN(n18805) );
  OAI211_X1 U20887 ( .C1(n18930), .C2(n18832), .A(n18806), .B(n18805), .ZN(
        P3_U2993) );
  INV_X1 U20888 ( .A(n18829), .ZN(n18842) );
  INV_X1 U20889 ( .A(n18832), .ZN(n18838) );
  AOI22_X1 U20890 ( .A1(n19035), .A2(n18838), .B1(n19017), .B2(n18837), .ZN(
        n18808) );
  AOI22_X1 U20891 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n19018), .B1(
        n19105), .B2(n18839), .ZN(n18807) );
  OAI211_X1 U20892 ( .C1(n18930), .C2(n18842), .A(n18808), .B(n18807), .ZN(
        P3_U2985) );
  AOI22_X1 U20893 ( .A1(n19035), .A2(n18829), .B1(n19022), .B2(n18837), .ZN(
        n18810) );
  AOI22_X1 U20894 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19024), .B1(
        n19023), .B2(n18839), .ZN(n18809) );
  OAI211_X1 U20895 ( .C1(n19027), .C2(n18832), .A(n18810), .B(n18809), .ZN(
        P3_U2977) );
  AOI22_X1 U20896 ( .A1(n19047), .A2(n18838), .B1(n19028), .B2(n18837), .ZN(
        n18812) );
  AOI22_X1 U20897 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19030), .B1(
        n19029), .B2(n18839), .ZN(n18811) );
  OAI211_X1 U20898 ( .C1(n19027), .C2(n18842), .A(n18812), .B(n18811), .ZN(
        P3_U2969) );
  AOI22_X1 U20899 ( .A1(n19034), .A2(n18837), .B1(n19053), .B2(n18838), .ZN(
        n18814) );
  AOI22_X1 U20900 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19036), .B1(
        n19035), .B2(n18839), .ZN(n18813) );
  OAI211_X1 U20901 ( .C1(n19033), .C2(n18842), .A(n18814), .B(n18813), .ZN(
        P3_U2961) );
  AOI22_X1 U20902 ( .A1(n19053), .A2(n18829), .B1(n19040), .B2(n18837), .ZN(
        n18816) );
  AOI22_X1 U20903 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19042), .B1(
        n19041), .B2(n18839), .ZN(n18815) );
  OAI211_X1 U20904 ( .C1(n19045), .C2(n18832), .A(n18816), .B(n18815), .ZN(
        P3_U2953) );
  AOI22_X1 U20905 ( .A1(n19065), .A2(n18838), .B1(n19046), .B2(n18837), .ZN(
        n18818) );
  AOI22_X1 U20906 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19048), .B1(
        n19047), .B2(n18839), .ZN(n18817) );
  OAI211_X1 U20907 ( .C1(n19045), .C2(n18842), .A(n18818), .B(n18817), .ZN(
        P3_U2945) );
  AOI22_X1 U20908 ( .A1(n19065), .A2(n18829), .B1(n19052), .B2(n18837), .ZN(
        n18820) );
  AOI22_X1 U20909 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19054), .B1(
        n19053), .B2(n18839), .ZN(n18819) );
  OAI211_X1 U20910 ( .C1(n19057), .C2(n18832), .A(n18820), .B(n18819), .ZN(
        P3_U2937) );
  AOI22_X1 U20911 ( .A1(n19071), .A2(n18829), .B1(n19058), .B2(n18837), .ZN(
        n18822) );
  AOI22_X1 U20912 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19060), .B1(
        n19059), .B2(n18839), .ZN(n18821) );
  OAI211_X1 U20913 ( .C1(n19063), .C2(n18832), .A(n18822), .B(n18821), .ZN(
        P3_U2929) );
  AOI22_X1 U20914 ( .A1(n19083), .A2(n18838), .B1(n19064), .B2(n18837), .ZN(
        n18824) );
  AOI22_X1 U20915 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19066), .B1(
        n19065), .B2(n18839), .ZN(n18823) );
  OAI211_X1 U20916 ( .C1(n19063), .C2(n18842), .A(n18824), .B(n18823), .ZN(
        P3_U2921) );
  AOI22_X1 U20917 ( .A1(n19083), .A2(n18829), .B1(n19070), .B2(n18837), .ZN(
        n18826) );
  AOI22_X1 U20918 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19072), .B1(
        n19071), .B2(n18839), .ZN(n18825) );
  OAI211_X1 U20919 ( .C1(n19080), .C2(n18832), .A(n18826), .B(n18825), .ZN(
        P3_U2913) );
  AOI22_X1 U20920 ( .A1(n19090), .A2(n18829), .B1(n19075), .B2(n18837), .ZN(
        n18828) );
  AOI22_X1 U20921 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19077), .B1(
        n19076), .B2(n18839), .ZN(n18827) );
  OAI211_X1 U20922 ( .C1(n19088), .C2(n18832), .A(n18828), .B(n18827), .ZN(
        P3_U2905) );
  AOI22_X1 U20923 ( .A1(n19097), .A2(n18829), .B1(n19082), .B2(n18837), .ZN(
        n18831) );
  AOI22_X1 U20924 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19084), .B1(
        n19083), .B2(n18839), .ZN(n18830) );
  OAI211_X1 U20925 ( .C1(n18955), .C2(n18832), .A(n18831), .B(n18830), .ZN(
        P3_U2897) );
  AOI22_X1 U20926 ( .A1(n19096), .A2(n18838), .B1(n19089), .B2(n18837), .ZN(
        n18834) );
  AOI22_X1 U20927 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19091), .B1(
        n19090), .B2(n18839), .ZN(n18833) );
  OAI211_X1 U20928 ( .C1(n18955), .C2(n18842), .A(n18834), .B(n18833), .ZN(
        P3_U2889) );
  AOI22_X1 U20929 ( .A1(n19105), .A2(n18838), .B1(n19095), .B2(n18837), .ZN(
        n18836) );
  AOI22_X1 U20930 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19098), .B1(
        n19097), .B2(n18839), .ZN(n18835) );
  OAI211_X1 U20931 ( .C1(n19094), .C2(n18842), .A(n18836), .B(n18835), .ZN(
        P3_U2881) );
  AOI22_X1 U20932 ( .A1(n19023), .A2(n18838), .B1(n19103), .B2(n18837), .ZN(
        n18841) );
  AOI22_X1 U20933 ( .A1(P3_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n19108), .B1(
        n19107), .B2(n18839), .ZN(n18840) );
  OAI211_X1 U20934 ( .C1(n19101), .C2(n18842), .A(n18841), .B(n18840), .ZN(
        P3_U2873) );
  INV_X1 U20935 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n18843) );
  AOI22_X1 U20936 ( .A1(n19008), .A2(n18843), .B1(n20657), .B2(U215), .ZN(U255) );
  NAND2_X1 U20937 ( .A1(BUF2_REG_20__SCAN_IN), .A2(n18884), .ZN(n18882) );
  NAND2_X1 U20938 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n18884), .ZN(n18874) );
  INV_X1 U20939 ( .A(n18874), .ZN(n18878) );
  NOR2_X2 U20940 ( .A1(n20657), .A2(n19010), .ZN(n18877) );
  AOI22_X1 U20941 ( .A1(n19029), .A2(n18878), .B1(n19011), .B2(n18877), .ZN(
        n18846) );
  NOR2_X2 U20942 ( .A1(n18844), .A2(n19012), .ZN(n18879) );
  AOI22_X1 U20943 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n19014), .B1(
        n19096), .B2(n18879), .ZN(n18845) );
  OAI211_X1 U20944 ( .C1(n19112), .C2(n18882), .A(n18846), .B(n18845), .ZN(
        P3_U2992) );
  INV_X1 U20945 ( .A(n18882), .ZN(n18871) );
  AOI22_X1 U20946 ( .A1(n19029), .A2(n18871), .B1(n19017), .B2(n18877), .ZN(
        n18848) );
  AOI22_X1 U20947 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n19018), .B1(
        n19105), .B2(n18879), .ZN(n18847) );
  OAI211_X1 U20948 ( .C1(n19021), .C2(n18874), .A(n18848), .B(n18847), .ZN(
        P3_U2984) );
  AOI22_X1 U20949 ( .A1(n19035), .A2(n18871), .B1(n19022), .B2(n18877), .ZN(
        n18850) );
  AOI22_X1 U20950 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19024), .B1(
        n19023), .B2(n18879), .ZN(n18849) );
  OAI211_X1 U20951 ( .C1(n19027), .C2(n18874), .A(n18850), .B(n18849), .ZN(
        P3_U2976) );
  AOI22_X1 U20952 ( .A1(n19041), .A2(n18871), .B1(n19028), .B2(n18877), .ZN(
        n18852) );
  AOI22_X1 U20953 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n19030), .B1(
        n19029), .B2(n18879), .ZN(n18851) );
  OAI211_X1 U20954 ( .C1(n19033), .C2(n18874), .A(n18852), .B(n18851), .ZN(
        P3_U2968) );
  AOI22_X1 U20955 ( .A1(n19047), .A2(n18871), .B1(n19034), .B2(n18877), .ZN(
        n18854) );
  AOI22_X1 U20956 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19036), .B1(
        n19035), .B2(n18879), .ZN(n18853) );
  OAI211_X1 U20957 ( .C1(n19039), .C2(n18874), .A(n18854), .B(n18853), .ZN(
        P3_U2960) );
  AOI22_X1 U20958 ( .A1(n19053), .A2(n18871), .B1(n19040), .B2(n18877), .ZN(
        n18856) );
  AOI22_X1 U20959 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19042), .B1(
        n19041), .B2(n18879), .ZN(n18855) );
  OAI211_X1 U20960 ( .C1(n19045), .C2(n18874), .A(n18856), .B(n18855), .ZN(
        P3_U2952) );
  AOI22_X1 U20961 ( .A1(n19059), .A2(n18871), .B1(n19046), .B2(n18877), .ZN(
        n18858) );
  AOI22_X1 U20962 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19048), .B1(
        n19047), .B2(n18879), .ZN(n18857) );
  OAI211_X1 U20963 ( .C1(n19051), .C2(n18874), .A(n18858), .B(n18857), .ZN(
        P3_U2944) );
  AOI22_X1 U20964 ( .A1(n19071), .A2(n18878), .B1(n19052), .B2(n18877), .ZN(
        n18860) );
  AOI22_X1 U20965 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19054), .B1(
        n19053), .B2(n18879), .ZN(n18859) );
  OAI211_X1 U20966 ( .C1(n19051), .C2(n18882), .A(n18860), .B(n18859), .ZN(
        P3_U2936) );
  AOI22_X1 U20967 ( .A1(n19058), .A2(n18877), .B1(n19076), .B2(n18878), .ZN(
        n18862) );
  AOI22_X1 U20968 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19060), .B1(
        n19059), .B2(n18879), .ZN(n18861) );
  OAI211_X1 U20969 ( .C1(n19057), .C2(n18882), .A(n18862), .B(n18861), .ZN(
        P3_U2928) );
  AOI22_X1 U20970 ( .A1(n19076), .A2(n18871), .B1(n19064), .B2(n18877), .ZN(
        n18864) );
  AOI22_X1 U20971 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19066), .B1(
        n19065), .B2(n18879), .ZN(n18863) );
  OAI211_X1 U20972 ( .C1(n19069), .C2(n18874), .A(n18864), .B(n18863), .ZN(
        P3_U2920) );
  AOI22_X1 U20973 ( .A1(n19083), .A2(n18871), .B1(n19070), .B2(n18877), .ZN(
        n18866) );
  AOI22_X1 U20974 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19072), .B1(
        n19071), .B2(n18879), .ZN(n18865) );
  OAI211_X1 U20975 ( .C1(n19080), .C2(n18874), .A(n18866), .B(n18865), .ZN(
        P3_U2912) );
  AOI22_X1 U20976 ( .A1(n19097), .A2(n18878), .B1(n19075), .B2(n18877), .ZN(
        n18868) );
  AOI22_X1 U20977 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19077), .B1(
        n19076), .B2(n18879), .ZN(n18867) );
  OAI211_X1 U20978 ( .C1(n19080), .C2(n18882), .A(n18868), .B(n18867), .ZN(
        P3_U2904) );
  AOI22_X1 U20979 ( .A1(n19097), .A2(n18871), .B1(n19082), .B2(n18877), .ZN(
        n18870) );
  AOI22_X1 U20980 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19084), .B1(
        n19083), .B2(n18879), .ZN(n18869) );
  OAI211_X1 U20981 ( .C1(n18955), .C2(n18874), .A(n18870), .B(n18869), .ZN(
        P3_U2896) );
  AOI22_X1 U20982 ( .A1(n19107), .A2(n18871), .B1(n19089), .B2(n18877), .ZN(
        n18873) );
  AOI22_X1 U20983 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19091), .B1(
        n19090), .B2(n18879), .ZN(n18872) );
  OAI211_X1 U20984 ( .C1(n19094), .C2(n18874), .A(n18873), .B(n18872), .ZN(
        P3_U2888) );
  AOI22_X1 U20985 ( .A1(n19105), .A2(n18878), .B1(n19095), .B2(n18877), .ZN(
        n18876) );
  AOI22_X1 U20986 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19098), .B1(
        n19097), .B2(n18879), .ZN(n18875) );
  OAI211_X1 U20987 ( .C1(n19094), .C2(n18882), .A(n18876), .B(n18875), .ZN(
        P3_U2880) );
  AOI22_X1 U20988 ( .A1(n19023), .A2(n18878), .B1(n19103), .B2(n18877), .ZN(
        n18881) );
  AOI22_X1 U20989 ( .A1(P3_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n19108), .B1(
        n19107), .B2(n18879), .ZN(n18880) );
  OAI211_X1 U20990 ( .C1(n19101), .C2(n18882), .A(n18881), .B(n18880), .ZN(
        P3_U2872) );
  OAI22_X1 U20991 ( .A1(U215), .A2(P2_DATAO_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n18966), .ZN(n18883) );
  INV_X1 U20992 ( .A(n18883), .ZN(U254) );
  NAND2_X1 U20993 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n18884), .ZN(n18923) );
  NAND2_X1 U20994 ( .A1(BUF2_REG_19__SCAN_IN), .A2(n18884), .ZN(n18917) );
  INV_X1 U20995 ( .A(n18917), .ZN(n18919) );
  AND2_X1 U20996 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n18968), .ZN(n18918) );
  AOI22_X1 U20997 ( .A1(n19023), .A2(n18919), .B1(n19011), .B2(n18918), .ZN(
        n18887) );
  NOR2_X2 U20998 ( .A1(n18885), .A2(n19012), .ZN(n18920) );
  AOI22_X1 U20999 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n19014), .B1(
        n19096), .B2(n18920), .ZN(n18886) );
  OAI211_X1 U21000 ( .C1(n18930), .C2(n18923), .A(n18887), .B(n18886), .ZN(
        P3_U2991) );
  AOI22_X1 U21001 ( .A1(n19029), .A2(n18919), .B1(n19017), .B2(n18918), .ZN(
        n18889) );
  AOI22_X1 U21002 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n19018), .B1(
        n19105), .B2(n18920), .ZN(n18888) );
  OAI211_X1 U21003 ( .C1(n19021), .C2(n18923), .A(n18889), .B(n18888), .ZN(
        P3_U2983) );
  AOI22_X1 U21004 ( .A1(n19035), .A2(n18919), .B1(n19022), .B2(n18918), .ZN(
        n18891) );
  AOI22_X1 U21005 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19024), .B1(
        n19023), .B2(n18920), .ZN(n18890) );
  OAI211_X1 U21006 ( .C1(n19027), .C2(n18923), .A(n18891), .B(n18890), .ZN(
        P3_U2975) );
  AOI22_X1 U21007 ( .A1(n19041), .A2(n18919), .B1(n19028), .B2(n18918), .ZN(
        n18893) );
  AOI22_X1 U21008 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n19030), .B1(
        n19029), .B2(n18920), .ZN(n18892) );
  OAI211_X1 U21009 ( .C1(n19033), .C2(n18923), .A(n18893), .B(n18892), .ZN(
        P3_U2967) );
  AOI22_X1 U21010 ( .A1(n19047), .A2(n18919), .B1(n19034), .B2(n18918), .ZN(
        n18895) );
  AOI22_X1 U21011 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19036), .B1(
        n19035), .B2(n18920), .ZN(n18894) );
  OAI211_X1 U21012 ( .C1(n19039), .C2(n18923), .A(n18895), .B(n18894), .ZN(
        P3_U2959) );
  AOI22_X1 U21013 ( .A1(n19053), .A2(n18919), .B1(n19040), .B2(n18918), .ZN(
        n18897) );
  AOI22_X1 U21014 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19042), .B1(
        n19041), .B2(n18920), .ZN(n18896) );
  OAI211_X1 U21015 ( .C1(n19045), .C2(n18923), .A(n18897), .B(n18896), .ZN(
        P3_U2951) );
  AOI22_X1 U21016 ( .A1(n19059), .A2(n18919), .B1(n19046), .B2(n18918), .ZN(
        n18899) );
  AOI22_X1 U21017 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19048), .B1(
        n19047), .B2(n18920), .ZN(n18898) );
  OAI211_X1 U21018 ( .C1(n19051), .C2(n18923), .A(n18899), .B(n18898), .ZN(
        P3_U2943) );
  AOI22_X1 U21019 ( .A1(n19065), .A2(n18919), .B1(n19052), .B2(n18918), .ZN(
        n18901) );
  AOI22_X1 U21020 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19054), .B1(
        n19053), .B2(n18920), .ZN(n18900) );
  OAI211_X1 U21021 ( .C1(n19057), .C2(n18923), .A(n18901), .B(n18900), .ZN(
        P3_U2935) );
  AOI22_X1 U21022 ( .A1(n19071), .A2(n18919), .B1(n19058), .B2(n18918), .ZN(
        n18903) );
  AOI22_X1 U21023 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19060), .B1(
        n19059), .B2(n18920), .ZN(n18902) );
  OAI211_X1 U21024 ( .C1(n19063), .C2(n18923), .A(n18903), .B(n18902), .ZN(
        P3_U2927) );
  INV_X1 U21025 ( .A(n18923), .ZN(n18914) );
  AOI22_X1 U21026 ( .A1(n19083), .A2(n18914), .B1(n19064), .B2(n18918), .ZN(
        n18905) );
  AOI22_X1 U21027 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19066), .B1(
        n19065), .B2(n18920), .ZN(n18904) );
  OAI211_X1 U21028 ( .C1(n19063), .C2(n18917), .A(n18905), .B(n18904), .ZN(
        P3_U2919) );
  AOI22_X1 U21029 ( .A1(n19083), .A2(n18919), .B1(n19070), .B2(n18918), .ZN(
        n18907) );
  AOI22_X1 U21030 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19072), .B1(
        n19071), .B2(n18920), .ZN(n18906) );
  OAI211_X1 U21031 ( .C1(n19080), .C2(n18923), .A(n18907), .B(n18906), .ZN(
        P3_U2911) );
  AOI22_X1 U21032 ( .A1(n19097), .A2(n18914), .B1(n19075), .B2(n18918), .ZN(
        n18909) );
  AOI22_X1 U21033 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19077), .B1(
        n19076), .B2(n18920), .ZN(n18908) );
  OAI211_X1 U21034 ( .C1(n19080), .C2(n18917), .A(n18909), .B(n18908), .ZN(
        P3_U2903) );
  AOI22_X1 U21035 ( .A1(n19082), .A2(n18918), .B1(n19107), .B2(n18914), .ZN(
        n18911) );
  AOI22_X1 U21036 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19084), .B1(
        n19083), .B2(n18920), .ZN(n18910) );
  OAI211_X1 U21037 ( .C1(n19088), .C2(n18917), .A(n18911), .B(n18910), .ZN(
        P3_U2895) );
  AOI22_X1 U21038 ( .A1(n19096), .A2(n18914), .B1(n19089), .B2(n18918), .ZN(
        n18913) );
  AOI22_X1 U21039 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19091), .B1(
        n19090), .B2(n18920), .ZN(n18912) );
  OAI211_X1 U21040 ( .C1(n18955), .C2(n18917), .A(n18913), .B(n18912), .ZN(
        P3_U2887) );
  AOI22_X1 U21041 ( .A1(n19105), .A2(n18914), .B1(n19095), .B2(n18918), .ZN(
        n18916) );
  AOI22_X1 U21042 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19098), .B1(
        n19097), .B2(n18920), .ZN(n18915) );
  OAI211_X1 U21043 ( .C1(n19094), .C2(n18917), .A(n18916), .B(n18915), .ZN(
        P3_U2879) );
  AOI22_X1 U21044 ( .A1(n19105), .A2(n18919), .B1(n19103), .B2(n18918), .ZN(
        n18922) );
  AOI22_X1 U21045 ( .A1(P3_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n19108), .B1(
        n19107), .B2(n18920), .ZN(n18921) );
  OAI211_X1 U21046 ( .C1(n19112), .C2(n18923), .A(n18922), .B(n18921), .ZN(
        P3_U2871) );
  INV_X1 U21047 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n18924) );
  AOI22_X1 U21048 ( .A1(n19008), .A2(n18924), .B1(n20139), .B2(U215), .ZN(U253) );
  NAND2_X1 U21049 ( .A1(BUF2_REG_18__SCAN_IN), .A2(n18884), .ZN(n18965) );
  NAND2_X1 U21050 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n18884), .ZN(n18959) );
  INV_X1 U21051 ( .A(n18959), .ZN(n18961) );
  NOR2_X2 U21052 ( .A1(n20139), .A2(n19010), .ZN(n18960) );
  AOI22_X1 U21053 ( .A1(n19029), .A2(n18961), .B1(n19011), .B2(n18960), .ZN(
        n18927) );
  NOR2_X2 U21054 ( .A1(n18925), .A2(n19012), .ZN(n18962) );
  AOI22_X1 U21055 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n19014), .B1(
        n19096), .B2(n18962), .ZN(n18926) );
  OAI211_X1 U21056 ( .C1(n19112), .C2(n18965), .A(n18927), .B(n18926), .ZN(
        P3_U2990) );
  AOI22_X1 U21057 ( .A1(n19035), .A2(n18961), .B1(n19017), .B2(n18960), .ZN(
        n18929) );
  AOI22_X1 U21058 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n19018), .B1(
        n19105), .B2(n18962), .ZN(n18928) );
  OAI211_X1 U21059 ( .C1(n18930), .C2(n18965), .A(n18929), .B(n18928), .ZN(
        P3_U2982) );
  AOI22_X1 U21060 ( .A1(n19041), .A2(n18961), .B1(n19022), .B2(n18960), .ZN(
        n18932) );
  AOI22_X1 U21061 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19024), .B1(
        n19023), .B2(n18962), .ZN(n18931) );
  OAI211_X1 U21062 ( .C1(n19021), .C2(n18965), .A(n18932), .B(n18931), .ZN(
        P3_U2974) );
  AOI22_X1 U21063 ( .A1(n19047), .A2(n18961), .B1(n19028), .B2(n18960), .ZN(
        n18934) );
  AOI22_X1 U21064 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n19030), .B1(
        n19029), .B2(n18962), .ZN(n18933) );
  OAI211_X1 U21065 ( .C1(n19027), .C2(n18965), .A(n18934), .B(n18933), .ZN(
        P3_U2966) );
  AOI22_X1 U21066 ( .A1(n19034), .A2(n18960), .B1(n19053), .B2(n18961), .ZN(
        n18936) );
  AOI22_X1 U21067 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19036), .B1(
        n19035), .B2(n18962), .ZN(n18935) );
  OAI211_X1 U21068 ( .C1(n19033), .C2(n18965), .A(n18936), .B(n18935), .ZN(
        P3_U2958) );
  AOI22_X1 U21069 ( .A1(n19059), .A2(n18961), .B1(n19040), .B2(n18960), .ZN(
        n18938) );
  AOI22_X1 U21070 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19042), .B1(
        n19041), .B2(n18962), .ZN(n18937) );
  OAI211_X1 U21071 ( .C1(n19039), .C2(n18965), .A(n18938), .B(n18937), .ZN(
        P3_U2950) );
  AOI22_X1 U21072 ( .A1(n19065), .A2(n18961), .B1(n19046), .B2(n18960), .ZN(
        n18940) );
  AOI22_X1 U21073 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19048), .B1(
        n19047), .B2(n18962), .ZN(n18939) );
  OAI211_X1 U21074 ( .C1(n19045), .C2(n18965), .A(n18940), .B(n18939), .ZN(
        P3_U2942) );
  AOI22_X1 U21075 ( .A1(n19071), .A2(n18961), .B1(n19052), .B2(n18960), .ZN(
        n18942) );
  AOI22_X1 U21076 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19054), .B1(
        n19053), .B2(n18962), .ZN(n18941) );
  OAI211_X1 U21077 ( .C1(n19051), .C2(n18965), .A(n18942), .B(n18941), .ZN(
        P3_U2934) );
  INV_X1 U21078 ( .A(n18965), .ZN(n18956) );
  AOI22_X1 U21079 ( .A1(n19071), .A2(n18956), .B1(n19058), .B2(n18960), .ZN(
        n18944) );
  AOI22_X1 U21080 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19060), .B1(
        n19059), .B2(n18962), .ZN(n18943) );
  OAI211_X1 U21081 ( .C1(n19063), .C2(n18959), .A(n18944), .B(n18943), .ZN(
        P3_U2926) );
  AOI22_X1 U21082 ( .A1(n19083), .A2(n18961), .B1(n19064), .B2(n18960), .ZN(
        n18946) );
  AOI22_X1 U21083 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19066), .B1(
        n19065), .B2(n18962), .ZN(n18945) );
  OAI211_X1 U21084 ( .C1(n19063), .C2(n18965), .A(n18946), .B(n18945), .ZN(
        P3_U2918) );
  AOI22_X1 U21085 ( .A1(n19090), .A2(n18961), .B1(n19070), .B2(n18960), .ZN(
        n18948) );
  AOI22_X1 U21086 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19072), .B1(
        n19071), .B2(n18962), .ZN(n18947) );
  OAI211_X1 U21087 ( .C1(n19069), .C2(n18965), .A(n18948), .B(n18947), .ZN(
        P3_U2910) );
  AOI22_X1 U21088 ( .A1(n19097), .A2(n18961), .B1(n19075), .B2(n18960), .ZN(
        n18950) );
  AOI22_X1 U21089 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19077), .B1(
        n19076), .B2(n18962), .ZN(n18949) );
  OAI211_X1 U21090 ( .C1(n19080), .C2(n18965), .A(n18950), .B(n18949), .ZN(
        P3_U2902) );
  AOI22_X1 U21091 ( .A1(n19097), .A2(n18956), .B1(n19082), .B2(n18960), .ZN(
        n18952) );
  AOI22_X1 U21092 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19084), .B1(
        n19083), .B2(n18962), .ZN(n18951) );
  OAI211_X1 U21093 ( .C1(n18955), .C2(n18959), .A(n18952), .B(n18951), .ZN(
        P3_U2894) );
  AOI22_X1 U21094 ( .A1(n19096), .A2(n18961), .B1(n19089), .B2(n18960), .ZN(
        n18954) );
  AOI22_X1 U21095 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19091), .B1(
        n19090), .B2(n18962), .ZN(n18953) );
  OAI211_X1 U21096 ( .C1(n18955), .C2(n18965), .A(n18954), .B(n18953), .ZN(
        P3_U2886) );
  AOI22_X1 U21097 ( .A1(n19096), .A2(n18956), .B1(n19095), .B2(n18960), .ZN(
        n18958) );
  AOI22_X1 U21098 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19098), .B1(
        n19097), .B2(n18962), .ZN(n18957) );
  OAI211_X1 U21099 ( .C1(n19101), .C2(n18959), .A(n18958), .B(n18957), .ZN(
        P3_U2878) );
  AOI22_X1 U21100 ( .A1(n19023), .A2(n18961), .B1(n19103), .B2(n18960), .ZN(
        n18964) );
  AOI22_X1 U21101 ( .A1(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n19108), .B1(
        n19107), .B2(n18962), .ZN(n18963) );
  OAI211_X1 U21102 ( .C1(n19101), .C2(n18965), .A(n18964), .B(n18963), .ZN(
        P3_U2870) );
  OAI22_X1 U21103 ( .A1(U215), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n18966), .ZN(n18967) );
  INV_X1 U21104 ( .A(n18967), .ZN(U252) );
  NAND2_X1 U21105 ( .A1(n18884), .A2(BUF2_REG_17__SCAN_IN), .ZN(n19006) );
  NAND2_X1 U21106 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n18884), .ZN(n18998) );
  AND2_X1 U21107 ( .A1(n18968), .A2(BUF2_REG_1__SCAN_IN), .ZN(n19001) );
  AOI22_X1 U21108 ( .A1(n19029), .A2(n19002), .B1(n19011), .B2(n19001), .ZN(
        n18970) );
  NOR2_X2 U21109 ( .A1(n14680), .A2(n19012), .ZN(n19003) );
  AOI22_X1 U21110 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n19014), .B1(
        n19096), .B2(n19003), .ZN(n18969) );
  OAI211_X1 U21111 ( .C1(n19112), .C2(n19006), .A(n18970), .B(n18969), .ZN(
        P3_U2989) );
  INV_X1 U21112 ( .A(n19006), .ZN(n18995) );
  AOI22_X1 U21113 ( .A1(n19029), .A2(n18995), .B1(n19017), .B2(n19001), .ZN(
        n18972) );
  AOI22_X1 U21114 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n19018), .B1(
        n19105), .B2(n19003), .ZN(n18971) );
  OAI211_X1 U21115 ( .C1(n19021), .C2(n18998), .A(n18972), .B(n18971), .ZN(
        P3_U2981) );
  AOI22_X1 U21116 ( .A1(n19041), .A2(n19002), .B1(n19022), .B2(n19001), .ZN(
        n18974) );
  AOI22_X1 U21117 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19024), .B1(
        n19023), .B2(n19003), .ZN(n18973) );
  OAI211_X1 U21118 ( .C1(n19021), .C2(n19006), .A(n18974), .B(n18973), .ZN(
        P3_U2973) );
  AOI22_X1 U21119 ( .A1(n19041), .A2(n18995), .B1(n19028), .B2(n19001), .ZN(
        n18976) );
  AOI22_X1 U21120 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n19030), .B1(
        n19029), .B2(n19003), .ZN(n18975) );
  OAI211_X1 U21121 ( .C1(n19033), .C2(n18998), .A(n18976), .B(n18975), .ZN(
        P3_U2965) );
  AOI22_X1 U21122 ( .A1(n19034), .A2(n19001), .B1(n19053), .B2(n19002), .ZN(
        n18978) );
  AOI22_X1 U21123 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19036), .B1(
        n19035), .B2(n19003), .ZN(n18977) );
  OAI211_X1 U21124 ( .C1(n19033), .C2(n19006), .A(n18978), .B(n18977), .ZN(
        P3_U2957) );
  AOI22_X1 U21125 ( .A1(n19059), .A2(n19002), .B1(n19040), .B2(n19001), .ZN(
        n18980) );
  AOI22_X1 U21126 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19042), .B1(
        n19041), .B2(n19003), .ZN(n18979) );
  OAI211_X1 U21127 ( .C1(n19039), .C2(n19006), .A(n18980), .B(n18979), .ZN(
        P3_U2949) );
  AOI22_X1 U21128 ( .A1(n19059), .A2(n18995), .B1(n19046), .B2(n19001), .ZN(
        n18982) );
  AOI22_X1 U21129 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19048), .B1(
        n19047), .B2(n19003), .ZN(n18981) );
  OAI211_X1 U21130 ( .C1(n19051), .C2(n18998), .A(n18982), .B(n18981), .ZN(
        P3_U2941) );
  AOI22_X1 U21131 ( .A1(n19071), .A2(n19002), .B1(n19052), .B2(n19001), .ZN(
        n18984) );
  AOI22_X1 U21132 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19054), .B1(
        n19053), .B2(n19003), .ZN(n18983) );
  OAI211_X1 U21133 ( .C1(n19051), .C2(n19006), .A(n18984), .B(n18983), .ZN(
        P3_U2933) );
  AOI22_X1 U21134 ( .A1(n19058), .A2(n19001), .B1(n19076), .B2(n19002), .ZN(
        n18986) );
  AOI22_X1 U21135 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19060), .B1(
        n19059), .B2(n19003), .ZN(n18985) );
  OAI211_X1 U21136 ( .C1(n19057), .C2(n19006), .A(n18986), .B(n18985), .ZN(
        P3_U2925) );
  AOI22_X1 U21137 ( .A1(n19076), .A2(n18995), .B1(n19064), .B2(n19001), .ZN(
        n18988) );
  AOI22_X1 U21138 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19066), .B1(
        n19065), .B2(n19003), .ZN(n18987) );
  OAI211_X1 U21139 ( .C1(n19069), .C2(n18998), .A(n18988), .B(n18987), .ZN(
        P3_U2917) );
  AOI22_X1 U21140 ( .A1(n19083), .A2(n18995), .B1(n19070), .B2(n19001), .ZN(
        n18990) );
  AOI22_X1 U21141 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19072), .B1(
        n19071), .B2(n19003), .ZN(n18989) );
  OAI211_X1 U21142 ( .C1(n19080), .C2(n18998), .A(n18990), .B(n18989), .ZN(
        P3_U2909) );
  AOI22_X1 U21143 ( .A1(n19090), .A2(n18995), .B1(n19075), .B2(n19001), .ZN(
        n18992) );
  AOI22_X1 U21144 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19077), .B1(
        n19076), .B2(n19003), .ZN(n18991) );
  OAI211_X1 U21145 ( .C1(n19088), .C2(n18998), .A(n18992), .B(n18991), .ZN(
        P3_U2901) );
  AOI22_X1 U21146 ( .A1(n19082), .A2(n19001), .B1(n19107), .B2(n19002), .ZN(
        n18994) );
  AOI22_X1 U21147 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19084), .B1(
        n19083), .B2(n19003), .ZN(n18993) );
  OAI211_X1 U21148 ( .C1(n19088), .C2(n19006), .A(n18994), .B(n18993), .ZN(
        P3_U2893) );
  AOI22_X1 U21149 ( .A1(n19107), .A2(n18995), .B1(n19089), .B2(n19001), .ZN(
        n18997) );
  AOI22_X1 U21150 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19091), .B1(
        n19090), .B2(n19003), .ZN(n18996) );
  OAI211_X1 U21151 ( .C1(n19094), .C2(n18998), .A(n18997), .B(n18996), .ZN(
        P3_U2885) );
  AOI22_X1 U21152 ( .A1(n19105), .A2(n19002), .B1(n19095), .B2(n19001), .ZN(
        n19000) );
  AOI22_X1 U21153 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19098), .B1(
        n19097), .B2(n19003), .ZN(n18999) );
  OAI211_X1 U21154 ( .C1(n19094), .C2(n19006), .A(n19000), .B(n18999), .ZN(
        P3_U2877) );
  AOI22_X1 U21155 ( .A1(n19023), .A2(n19002), .B1(n19103), .B2(n19001), .ZN(
        n19005) );
  AOI22_X1 U21156 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n19108), .B1(
        n19107), .B2(n19003), .ZN(n19004) );
  OAI211_X1 U21157 ( .C1(n19101), .C2(n19006), .A(n19005), .B(n19004), .ZN(
        P3_U2869) );
  INV_X1 U21158 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n19007) );
  AOI22_X1 U21159 ( .A1(n19008), .A2(n19007), .B1(n20135), .B2(U215), .ZN(U251) );
  NAND2_X1 U21160 ( .A1(n18884), .A2(BUF2_REG_16__SCAN_IN), .ZN(n19087) );
  NOR2_X1 U21161 ( .A1(n16212), .A2(n19009), .ZN(n19081) );
  NOR2_X2 U21162 ( .A1(n19010), .A2(n20135), .ZN(n19102) );
  AOI22_X1 U21163 ( .A1(n19029), .A2(n19081), .B1(n19011), .B2(n19102), .ZN(
        n19016) );
  NOR2_X2 U21164 ( .A1(n19013), .A2(n19012), .ZN(n19106) );
  AOI22_X1 U21165 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n19014), .B1(
        n19096), .B2(n19106), .ZN(n19015) );
  OAI211_X1 U21166 ( .C1(n19112), .C2(n19087), .A(n19016), .B(n19015), .ZN(
        P3_U2988) );
  INV_X1 U21167 ( .A(n19087), .ZN(n19104) );
  AOI22_X1 U21168 ( .A1(n19029), .A2(n19104), .B1(n19017), .B2(n19102), .ZN(
        n19020) );
  AOI22_X1 U21169 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n19018), .B1(
        n19105), .B2(n19106), .ZN(n19019) );
  OAI211_X1 U21170 ( .C1(n19021), .C2(n19111), .A(n19020), .B(n19019), .ZN(
        P3_U2980) );
  AOI22_X1 U21171 ( .A1(n19035), .A2(n19104), .B1(n19022), .B2(n19102), .ZN(
        n19026) );
  AOI22_X1 U21172 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n19024), .B1(
        n19023), .B2(n19106), .ZN(n19025) );
  OAI211_X1 U21173 ( .C1(n19027), .C2(n19111), .A(n19026), .B(n19025), .ZN(
        P3_U2972) );
  AOI22_X1 U21174 ( .A1(n19041), .A2(n19104), .B1(n19028), .B2(n19102), .ZN(
        n19032) );
  AOI22_X1 U21175 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n19030), .B1(
        n19029), .B2(n19106), .ZN(n19031) );
  OAI211_X1 U21176 ( .C1(n19033), .C2(n19111), .A(n19032), .B(n19031), .ZN(
        P3_U2964) );
  AOI22_X1 U21177 ( .A1(n19047), .A2(n19104), .B1(n19034), .B2(n19102), .ZN(
        n19038) );
  AOI22_X1 U21178 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19036), .B1(
        n19035), .B2(n19106), .ZN(n19037) );
  OAI211_X1 U21179 ( .C1(n19039), .C2(n19111), .A(n19038), .B(n19037), .ZN(
        P3_U2956) );
  AOI22_X1 U21180 ( .A1(n19053), .A2(n19104), .B1(n19040), .B2(n19102), .ZN(
        n19044) );
  AOI22_X1 U21181 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19042), .B1(
        n19041), .B2(n19106), .ZN(n19043) );
  OAI211_X1 U21182 ( .C1(n19045), .C2(n19111), .A(n19044), .B(n19043), .ZN(
        P3_U2948) );
  AOI22_X1 U21183 ( .A1(n19059), .A2(n19104), .B1(n19046), .B2(n19102), .ZN(
        n19050) );
  AOI22_X1 U21184 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n19048), .B1(
        n19047), .B2(n19106), .ZN(n19049) );
  OAI211_X1 U21185 ( .C1(n19051), .C2(n19111), .A(n19050), .B(n19049), .ZN(
        P3_U2940) );
  AOI22_X1 U21186 ( .A1(n19065), .A2(n19104), .B1(n19052), .B2(n19102), .ZN(
        n19056) );
  AOI22_X1 U21187 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19054), .B1(
        n19053), .B2(n19106), .ZN(n19055) );
  OAI211_X1 U21188 ( .C1(n19057), .C2(n19111), .A(n19056), .B(n19055), .ZN(
        P3_U2932) );
  AOI22_X1 U21189 ( .A1(n19071), .A2(n19104), .B1(n19058), .B2(n19102), .ZN(
        n19062) );
  AOI22_X1 U21190 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n19060), .B1(
        n19059), .B2(n19106), .ZN(n19061) );
  OAI211_X1 U21191 ( .C1(n19063), .C2(n19111), .A(n19062), .B(n19061), .ZN(
        P3_U2924) );
  AOI22_X1 U21192 ( .A1(n19076), .A2(n19104), .B1(n19064), .B2(n19102), .ZN(
        n19068) );
  AOI22_X1 U21193 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n19066), .B1(
        n19065), .B2(n19106), .ZN(n19067) );
  OAI211_X1 U21194 ( .C1(n19069), .C2(n19111), .A(n19068), .B(n19067), .ZN(
        P3_U2916) );
  AOI22_X1 U21195 ( .A1(n19083), .A2(n19104), .B1(n19070), .B2(n19102), .ZN(
        n19074) );
  AOI22_X1 U21196 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n19072), .B1(
        n19071), .B2(n19106), .ZN(n19073) );
  OAI211_X1 U21197 ( .C1(n19080), .C2(n19111), .A(n19074), .B(n19073), .ZN(
        P3_U2908) );
  AOI22_X1 U21198 ( .A1(n19097), .A2(n19081), .B1(n19075), .B2(n19102), .ZN(
        n19079) );
  AOI22_X1 U21199 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n19077), .B1(
        n19076), .B2(n19106), .ZN(n19078) );
  OAI211_X1 U21200 ( .C1(n19080), .C2(n19087), .A(n19079), .B(n19078), .ZN(
        P3_U2900) );
  AOI22_X1 U21201 ( .A1(n19082), .A2(n19102), .B1(n19107), .B2(n19081), .ZN(
        n19086) );
  AOI22_X1 U21202 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19084), .B1(
        n19083), .B2(n19106), .ZN(n19085) );
  OAI211_X1 U21203 ( .C1(n19088), .C2(n19087), .A(n19086), .B(n19085), .ZN(
        P3_U2892) );
  AOI22_X1 U21204 ( .A1(n19107), .A2(n19104), .B1(n19089), .B2(n19102), .ZN(
        n19093) );
  AOI22_X1 U21205 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19091), .B1(
        n19090), .B2(n19106), .ZN(n19092) );
  OAI211_X1 U21206 ( .C1(n19094), .C2(n19111), .A(n19093), .B(n19092), .ZN(
        P3_U2884) );
  AOI22_X1 U21207 ( .A1(n19096), .A2(n19104), .B1(n19095), .B2(n19102), .ZN(
        n19100) );
  AOI22_X1 U21208 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19098), .B1(
        n19097), .B2(n19106), .ZN(n19099) );
  OAI211_X1 U21209 ( .C1(n19101), .C2(n19111), .A(n19100), .B(n19099), .ZN(
        P3_U2876) );
  AOI22_X1 U21210 ( .A1(n19105), .A2(n19104), .B1(n19103), .B2(n19102), .ZN(
        n19110) );
  AOI22_X1 U21211 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n19108), .B1(
        n19107), .B2(n19106), .ZN(n19109) );
  OAI211_X1 U21212 ( .C1(n19112), .C2(n19111), .A(n19110), .B(n19109), .ZN(
        P3_U2868) );
  AOI22_X1 U21213 ( .A1(n19654), .A2(BUF1_REG_31__SCAN_IN), .B1(n19548), .B2(
        n19113), .ZN(n19115) );
  AOI22_X1 U21214 ( .A1(P2_EAX_REG_31__SCAN_IN), .A2(n19652), .B1(n19655), 
        .B2(BUF2_REG_31__SCAN_IN), .ZN(n19114) );
  NAND2_X1 U21215 ( .A1(n19115), .A2(n19114), .ZN(P2_U2888) );
  AOI22_X1 U21216 ( .A1(n19556), .A2(P2_UWORD_REG_14__SCAN_IN), .B1(
        P2_EAX_REG_30__SCAN_IN), .B2(n19667), .ZN(n19117) );
  OAI21_X1 U21217 ( .B1(n19119), .B2(n19670), .A(n19117), .ZN(P2_U2966) );
  AOI22_X1 U21218 ( .A1(n19556), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(
        P2_EAX_REG_14__SCAN_IN), .B2(n19667), .ZN(n19118) );
  OAI21_X1 U21219 ( .B1(n19119), .B2(n19670), .A(n19118), .ZN(P2_U2981) );
  AOI22_X1 U21220 ( .A1(n19556), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(
        P2_EAX_REG_29__SCAN_IN), .B2(n19667), .ZN(n19120) );
  OAI21_X1 U21221 ( .B1(n19122), .B2(n19670), .A(n19120), .ZN(P2_U2965) );
  AOI22_X1 U21222 ( .A1(n19556), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(
        P2_EAX_REG_13__SCAN_IN), .B2(n19667), .ZN(n19121) );
  OAI21_X1 U21223 ( .B1(n19122), .B2(n19670), .A(n19121), .ZN(P2_U2980) );
  AOI22_X1 U21224 ( .A1(n19668), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(
        P2_EAX_REG_28__SCAN_IN), .B2(n19667), .ZN(n19123) );
  OAI21_X1 U21225 ( .B1(n19125), .B2(n19670), .A(n19123), .ZN(P2_U2964) );
  AOI22_X1 U21226 ( .A1(n19556), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(
        P2_EAX_REG_12__SCAN_IN), .B2(n19667), .ZN(n19124) );
  OAI21_X1 U21227 ( .B1(n19125), .B2(n19670), .A(n19124), .ZN(P2_U2979) );
  AOI22_X1 U21228 ( .A1(n19556), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(
        P2_EAX_REG_27__SCAN_IN), .B2(n19667), .ZN(n19126) );
  OAI21_X1 U21229 ( .B1(n19128), .B2(n19670), .A(n19126), .ZN(P2_U2963) );
  AOI22_X1 U21230 ( .A1(n19556), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n19667), 
        .B2(P2_EAX_REG_11__SCAN_IN), .ZN(n19127) );
  OAI21_X1 U21231 ( .B1(n19128), .B2(n19670), .A(n19127), .ZN(P2_U2978) );
  AOI22_X1 U21232 ( .A1(n19130), .A2(n19129), .B1(n19652), .B2(
        P2_EAX_REG_10__SCAN_IN), .ZN(n19131) );
  OAI21_X1 U21233 ( .B1(n19410), .B2(n19132), .A(n19131), .ZN(P2_U2909) );
  AOI22_X1 U21234 ( .A1(n19556), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(
        P2_EAX_REG_25__SCAN_IN), .B2(n19667), .ZN(n19133) );
  OAI21_X1 U21235 ( .B1(n19135), .B2(n19670), .A(n19133), .ZN(P2_U2961) );
  AOI22_X1 U21236 ( .A1(n19556), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n19667), 
        .B2(P2_EAX_REG_9__SCAN_IN), .ZN(n19134) );
  OAI21_X1 U21237 ( .B1(n19135), .B2(n19670), .A(n19134), .ZN(P2_U2976) );
  AOI22_X1 U21238 ( .A1(n19556), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(
        P2_EAX_REG_24__SCAN_IN), .B2(n19667), .ZN(n19136) );
  OAI21_X1 U21239 ( .B1(n19138), .B2(n19670), .A(n19136), .ZN(P2_U2960) );
  AOI22_X1 U21240 ( .A1(n19556), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n19667), 
        .B2(P2_EAX_REG_8__SCAN_IN), .ZN(n19137) );
  OAI21_X1 U21241 ( .B1(n19138), .B2(n19670), .A(n19137), .ZN(P2_U2975) );
  AOI22_X1 U21242 ( .A1(n19556), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n19667), 
        .B2(P2_EAX_REG_23__SCAN_IN), .ZN(n19139) );
  OAI21_X1 U21243 ( .B1(n19146), .B2(n19670), .A(n19139), .ZN(P2_U2959) );
  AOI22_X1 U21244 ( .A1(n19556), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n19667), 
        .B2(P2_EAX_REG_7__SCAN_IN), .ZN(n19140) );
  OAI21_X1 U21245 ( .B1(n19146), .B2(n19670), .A(n19140), .ZN(P2_U2974) );
  NAND3_X1 U21246 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19153) );
  OAI21_X1 U21247 ( .B1(n19169), .B2(n19295), .A(n19153), .ZN(n19144) );
  INV_X1 U21248 ( .A(n19334), .ZN(n19251) );
  NAND2_X1 U21249 ( .A1(n14968), .A2(n19251), .ZN(n19142) );
  OAI21_X1 U21250 ( .B1(n19332), .B2(n19677), .A(n19331), .ZN(n19141) );
  NAND2_X1 U21251 ( .A1(n19142), .A2(n19141), .ZN(n19143) );
  OAI21_X1 U21252 ( .B1(n14968), .B2(n19677), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19145) );
  OAI21_X1 U21253 ( .B1(n19153), .B2(n19326), .A(n19145), .ZN(n19678) );
  NOR2_X2 U21254 ( .A1(n19146), .A2(n19673), .ZN(n19345) );
  NOR2_X2 U21255 ( .A1(n13233), .A2(n19675), .ZN(n19342) );
  AOI22_X1 U21256 ( .A1(n19678), .A2(n19345), .B1(n19677), .B2(n19342), .ZN(
        n19149) );
  OAI22_X2 U21257 ( .A1(n20082), .A2(n19681), .B1(n16219), .B2(n19679), .ZN(
        n19344) );
  NOR2_X2 U21258 ( .A1(n19169), .A2(n19293), .ZN(n19687) );
  AOI22_X1 U21259 ( .A1(BUF1_REG_31__SCAN_IN), .A2(n19672), .B1(
        BUF2_REG_31__SCAN_IN), .B2(n19671), .ZN(n19341) );
  INV_X1 U21260 ( .A(n19341), .ZN(n19343) );
  AOI22_X1 U21261 ( .A1(n19784), .A2(n19344), .B1(n19687), .B2(n19343), .ZN(
        n19148) );
  OAI211_X1 U21262 ( .C1(n19610), .C2(n19150), .A(n19149), .B(n19148), .ZN(
        P2_U3175) );
  NOR2_X2 U21263 ( .A1(n19169), .A2(n19306), .ZN(n19695) );
  INV_X1 U21264 ( .A(n19695), .ZN(n19164) );
  NOR2_X1 U21265 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19153), .ZN(
        n19686) );
  AOI22_X1 U21266 ( .A1(n19344), .A2(n19687), .B1(n19686), .B2(n19342), .ZN(
        n19163) );
  NAND2_X1 U21267 ( .A1(n19293), .A2(n19306), .ZN(n19198) );
  NAND2_X1 U21268 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n19198), .ZN(n19314) );
  OAI21_X1 U21269 ( .B1(n19169), .B2(n19314), .A(n19316), .ZN(n19158) );
  INV_X1 U21270 ( .A(n19158), .ZN(n19155) );
  NAND3_X1 U21271 ( .A1(n19296), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19179) );
  NOR2_X1 U21272 ( .A1(n19323), .A2(n19179), .ZN(n19692) );
  INV_X1 U21273 ( .A(n19692), .ZN(n19166) );
  NAND2_X1 U21274 ( .A1(n14960), .A2(n19251), .ZN(n19154) );
  AOI22_X1 U21275 ( .A1(n19155), .A2(n19166), .B1(n19252), .B2(n19154), .ZN(
        n19156) );
  AOI21_X1 U21276 ( .B1(n19686), .B2(n19331), .A(n19156), .ZN(n19688) );
  NOR2_X1 U21277 ( .A1(n19692), .A2(n19686), .ZN(n19157) );
  OR2_X1 U21278 ( .A1(n19158), .A2(n19157), .ZN(n19160) );
  OAI21_X1 U21279 ( .B1(n14960), .B2(n19686), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19159) );
  INV_X1 U21280 ( .A(n19691), .ZN(n19161) );
  AOI22_X1 U21281 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n19688), .B1(
        n19345), .B2(n19161), .ZN(n19162) );
  OAI211_X1 U21282 ( .C1(n19341), .C2(n19164), .A(n19163), .B(n19162), .ZN(
        P2_U3167) );
  OAI21_X1 U21283 ( .B1(n14961), .B2(n19692), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19165) );
  OAI21_X1 U21284 ( .B1(n19179), .B2(n19326), .A(n19165), .ZN(n19693) );
  AOI22_X1 U21285 ( .A1(n19693), .A2(n19345), .B1(n19342), .B2(n19692), .ZN(
        n19174) );
  AOI21_X1 U21286 ( .B1(n19166), .B2(n19326), .A(n19673), .ZN(n19172) );
  INV_X1 U21287 ( .A(n14961), .ZN(n19167) );
  NOR2_X1 U21288 ( .A1(n19167), .A2(n19334), .ZN(n19171) );
  OR2_X1 U21289 ( .A1(n19168), .A2(n21695), .ZN(n19218) );
  OAI21_X1 U21290 ( .B1(n19169), .B2(n19218), .A(n19179), .ZN(n19170) );
  OAI21_X1 U21291 ( .B1(n19172), .B2(n19171), .A(n19170), .ZN(n19694) );
  AOI22_X1 U21292 ( .A1(n19344), .A2(n19695), .B1(
        P2_INSTQUEUE_REG_13__7__SCAN_IN), .B2(n19694), .ZN(n19173) );
  OAI211_X1 U21293 ( .C1(n19341), .C2(n19698), .A(n19174), .B(n19173), .ZN(
        P2_U3159) );
  INV_X1 U21294 ( .A(n19175), .ZN(n19181) );
  INV_X1 U21295 ( .A(n19176), .ZN(n19178) );
  INV_X1 U21296 ( .A(n19248), .ZN(n19177) );
  NAND2_X1 U21297 ( .A1(n19178), .A2(n19177), .ZN(n19282) );
  NOR2_X1 U21298 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19179), .ZN(
        n19699) );
  OAI21_X1 U21299 ( .B1(n14970), .B2(n19699), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19180) );
  OAI21_X1 U21300 ( .B1(n19181), .B2(n19282), .A(n19180), .ZN(n19700) );
  AOI22_X1 U21301 ( .A1(n19700), .A2(n19345), .B1(n19342), .B2(n19699), .ZN(
        n19188) );
  OAI21_X1 U21302 ( .B1(n19701), .B2(n19368), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19182) );
  OAI21_X1 U21303 ( .B1(n19282), .B2(n19200), .A(n19182), .ZN(n19186) );
  INV_X1 U21304 ( .A(n14970), .ZN(n19184) );
  OAI21_X1 U21305 ( .B1(n19316), .B2(n19699), .A(n19331), .ZN(n19183) );
  OAI21_X1 U21306 ( .B1(n19184), .B2(n19334), .A(n19183), .ZN(n19185) );
  NAND2_X1 U21307 ( .A1(n19186), .A2(n19185), .ZN(n19702) );
  AOI22_X1 U21308 ( .A1(n19702), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n19344), .B2(n19701), .ZN(n19187) );
  OAI211_X1 U21309 ( .C1(n19341), .C2(n19710), .A(n19188), .B(n19187), .ZN(
        P2_U3151) );
  NAND3_X1 U21310 ( .A1(n19231), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19199) );
  OAI21_X1 U21311 ( .B1(n19217), .B2(n19295), .A(n19199), .ZN(n19192) );
  NAND2_X1 U21312 ( .A1(n14967), .A2(n19251), .ZN(n19190) );
  NOR2_X1 U21313 ( .A1(n19323), .A2(n19199), .ZN(n19705) );
  NOR2_X1 U21314 ( .A1(n19316), .A2(n19705), .ZN(n19189) );
  AOI21_X1 U21315 ( .B1(n19190), .B2(n19189), .A(n19673), .ZN(n19191) );
  OAI21_X1 U21316 ( .B1(n14967), .B2(n19705), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19193) );
  OAI21_X1 U21317 ( .B1(n19199), .B2(n19326), .A(n19193), .ZN(n19706) );
  AOI22_X1 U21318 ( .A1(n19706), .A2(n19345), .B1(n19342), .B2(n19705), .ZN(
        n19195) );
  NOR2_X2 U21319 ( .A1(n19217), .A2(n19293), .ZN(n19712) );
  AOI22_X1 U21320 ( .A1(n19368), .A2(n19344), .B1(n19712), .B2(n19343), .ZN(
        n19194) );
  OAI211_X1 U21321 ( .C1(n19422), .C2(n19196), .A(n19195), .B(n19194), .ZN(
        P2_U3143) );
  AOI21_X1 U21322 ( .B1(n19198), .B2(n19197), .A(n19326), .ZN(n19207) );
  NOR2_X1 U21323 ( .A1(n19199), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n19711) );
  INV_X1 U21324 ( .A(n19711), .ZN(n19205) );
  NOR3_X1 U21325 ( .A1(n19200), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19229) );
  NAND2_X1 U21326 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19229), .ZN(
        n19221) );
  NAND2_X1 U21327 ( .A1(n19205), .A2(n19221), .ZN(n19209) );
  INV_X1 U21328 ( .A(n19204), .ZN(n19201) );
  AOI21_X1 U21329 ( .B1(n19201), .B2(n19205), .A(n19264), .ZN(n19202) );
  INV_X1 U21330 ( .A(n19345), .ZN(n19277) );
  NOR2_X2 U21331 ( .A1(n19217), .A2(n19306), .ZN(n19718) );
  AOI22_X1 U21332 ( .A1(n19343), .A2(n19718), .B1(n19711), .B2(n19342), .ZN(
        n19212) );
  NAND2_X1 U21333 ( .A1(n19204), .A2(n19203), .ZN(n19206) );
  AOI21_X1 U21334 ( .B1(n19206), .B2(n19205), .A(n19673), .ZN(n19210) );
  INV_X1 U21335 ( .A(n19252), .ZN(n19224) );
  INV_X1 U21336 ( .A(n19207), .ZN(n19208) );
  AOI22_X1 U21337 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19713), .B1(
        n19712), .B2(n19344), .ZN(n19211) );
  OAI211_X1 U21338 ( .C1(n19716), .C2(n19277), .A(n19212), .B(n19211), .ZN(
        P2_U3135) );
  INV_X1 U21339 ( .A(n19229), .ZN(n19213) );
  NOR2_X1 U21340 ( .A1(n19326), .A2(n19213), .ZN(n19216) );
  INV_X1 U21341 ( .A(n19214), .ZN(n19220) );
  AOI21_X1 U21342 ( .B1(n19220), .B2(n19221), .A(n19264), .ZN(n19215) );
  INV_X1 U21343 ( .A(n19221), .ZN(n19717) );
  AOI22_X1 U21344 ( .A1(n19343), .A2(n19724), .B1(n19717), .B2(n19342), .ZN(
        n19228) );
  INV_X1 U21346 ( .A(n19218), .ZN(n19262) );
  NAND2_X1 U21347 ( .A1(n19219), .A2(n19262), .ZN(n19329) );
  NOR2_X1 U21348 ( .A1(n19328), .A2(n19329), .ZN(n19225) );
  NOR2_X1 U21349 ( .A1(n19220), .A2(n19334), .ZN(n19223) );
  NOR2_X1 U21350 ( .A1(n19673), .A2(n19221), .ZN(n19222) );
  OAI33_X1 U21351 ( .A1(1'b0), .A2(n19225), .A3(n19229), .B1(n19224), .B2(
        n19223), .B3(n19222), .ZN(n19719) );
  AOI22_X1 U21352 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n11085), .B1(
        n19718), .B2(n19344), .ZN(n19227) );
  OAI211_X1 U21353 ( .C1(n19722), .C2(n19277), .A(n19228), .B(n19227), .ZN(
        P2_U3127) );
  AND2_X1 U21354 ( .A1(n19323), .A2(n19229), .ZN(n19723) );
  AOI22_X1 U21355 ( .A1(n19344), .A2(n19724), .B1(n19723), .B2(n19342), .ZN(
        n19240) );
  OAI21_X1 U21356 ( .B1(n19724), .B2(n19625), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19230) );
  NAND2_X1 U21357 ( .A1(n19230), .A2(n19332), .ZN(n19238) );
  NOR2_X1 U21358 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19231), .ZN(
        n19257) );
  AND2_X1 U21359 ( .A1(n19232), .A2(n19257), .ZN(n19729) );
  NOR2_X1 U21360 ( .A1(n19238), .A2(n19729), .ZN(n19233) );
  OAI21_X1 U21361 ( .B1(n19723), .B2(n19234), .A(n19331), .ZN(n19726) );
  NOR2_X1 U21362 ( .A1(n19729), .A2(n19723), .ZN(n19237) );
  OAI21_X1 U21363 ( .B1(n19235), .B2(n19723), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19236) );
  AOI22_X1 U21364 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19726), .B1(
        n19345), .B2(n19725), .ZN(n19239) );
  OAI211_X1 U21365 ( .C1(n19341), .C2(n19735), .A(n19240), .B(n19239), .ZN(
        P2_U3119) );
  NAND2_X1 U21366 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19257), .ZN(
        n19250) );
  OAI21_X1 U21367 ( .B1(n15112), .B2(n19729), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19241) );
  OAI21_X1 U21368 ( .B1(n19250), .B2(n19326), .A(n19241), .ZN(n19730) );
  AOI22_X1 U21369 ( .A1(n19730), .A2(n19345), .B1(n19729), .B2(n19342), .ZN(
        n19247) );
  INV_X1 U21370 ( .A(n19250), .ZN(n19244) );
  AOI21_X1 U21371 ( .B1(n15112), .B2(n19251), .A(n19729), .ZN(n19242) );
  OAI21_X1 U21372 ( .B1(n19242), .B2(n19673), .A(n19252), .ZN(n19243) );
  OAI21_X1 U21373 ( .B1(n19245), .B2(n19244), .A(n19243), .ZN(n19732) );
  AOI22_X1 U21374 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19732), .B1(
        n19625), .B2(n19344), .ZN(n19246) );
  OAI211_X1 U21375 ( .C1(n19341), .C2(n19741), .A(n19247), .B(n19246), .ZN(
        P2_U3111) );
  NAND2_X1 U21376 ( .A1(n19248), .A2(n19257), .ZN(n19249) );
  OAI21_X1 U21377 ( .B1(n19267), .B2(n19314), .A(n19249), .ZN(n19256) );
  NOR2_X1 U21378 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19250), .ZN(
        n19736) );
  INV_X1 U21379 ( .A(n19736), .ZN(n19254) );
  NAND2_X1 U21380 ( .A1(n15111), .A2(n19251), .ZN(n19253) );
  OAI211_X1 U21381 ( .C1(n19673), .C2(n19254), .A(n19253), .B(n19252), .ZN(
        n19255) );
  INV_X1 U21382 ( .A(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n19261) );
  INV_X1 U21383 ( .A(n19257), .ZN(n19279) );
  OAI21_X1 U21384 ( .B1(n15111), .B2(n19736), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19258) );
  OAI21_X1 U21385 ( .B1(n19308), .B2(n19279), .A(n19258), .ZN(n19737) );
  AOI22_X1 U21386 ( .A1(n19737), .A2(n19345), .B1(n19342), .B2(n19736), .ZN(
        n19260) );
  NOR2_X2 U21387 ( .A1(n19267), .A2(n19306), .ZN(n19743) );
  AOI22_X1 U21388 ( .A1(n19731), .A2(n19344), .B1(n19743), .B2(n19343), .ZN(
        n19259) );
  OAI211_X1 U21389 ( .C1(n19631), .C2(n19261), .A(n19260), .B(n19259), .ZN(
        P2_U3103) );
  INV_X1 U21390 ( .A(n19267), .ZN(n19263) );
  AOI21_X1 U21391 ( .B1(n19263), .B2(n19262), .A(n19326), .ZN(n19269) );
  NOR2_X1 U21392 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19279), .ZN(
        n19273) );
  INV_X1 U21393 ( .A(n14969), .ZN(n19271) );
  NAND2_X1 U21394 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19273), .ZN(
        n19268) );
  AOI21_X1 U21395 ( .B1(n19271), .B2(n19268), .A(n19264), .ZN(n19265) );
  INV_X1 U21396 ( .A(n19268), .ZN(n19742) );
  AOI22_X1 U21397 ( .A1(n19343), .A2(n19750), .B1(n19742), .B2(n19342), .ZN(
        n19276) );
  INV_X1 U21398 ( .A(n19269), .ZN(n19274) );
  OAI21_X1 U21399 ( .B1(n19316), .B2(n19742), .A(n19331), .ZN(n19270) );
  OAI21_X1 U21400 ( .B1(n19271), .B2(n19334), .A(n19270), .ZN(n19272) );
  AOI22_X1 U21401 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19744), .B1(
        n19743), .B2(n19344), .ZN(n19275) );
  OAI211_X1 U21402 ( .C1(n19748), .C2(n19277), .A(n19276), .B(n19275), .ZN(
        P2_U3095) );
  NOR2_X1 U21403 ( .A1(n19280), .A2(n19279), .ZN(n19749) );
  AOI22_X1 U21404 ( .A1(n19344), .A2(n19750), .B1(n19749), .B2(n19342), .ZN(
        n19292) );
  OAI21_X1 U21405 ( .B1(n19757), .B2(n19750), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19281) );
  NAND2_X1 U21406 ( .A1(n19281), .A2(n19332), .ZN(n19290) );
  NOR2_X1 U21407 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19282), .ZN(
        n19287) );
  INV_X1 U21408 ( .A(n19749), .ZN(n19283) );
  AOI21_X1 U21409 ( .B1(n19283), .B2(n19326), .A(n19673), .ZN(n19286) );
  INV_X1 U21410 ( .A(n14966), .ZN(n19284) );
  NOR2_X1 U21411 ( .A1(n19284), .A2(n19334), .ZN(n19285) );
  INV_X1 U21412 ( .A(n19287), .ZN(n19289) );
  OAI21_X1 U21413 ( .B1(n14966), .B2(n19749), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19288) );
  AOI22_X1 U21414 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19752), .B1(
        n19345), .B2(n19751), .ZN(n19291) );
  OAI211_X1 U21415 ( .C1(n19341), .C2(n19755), .A(n19292), .B(n19291), .ZN(
        P2_U3087) );
  NOR2_X1 U21416 ( .A1(n19294), .A2(n19322), .ZN(n19756) );
  AOI22_X1 U21417 ( .A1(n19344), .A2(n19757), .B1(n19756), .B2(n19342), .ZN(
        n19305) );
  OAI21_X1 U21418 ( .B1(n19315), .B2(n19295), .A(n19316), .ZN(n19303) );
  NOR2_X1 U21419 ( .A1(n19296), .A2(n19322), .ZN(n19300) );
  INV_X1 U21420 ( .A(n19301), .ZN(n19298) );
  OAI21_X1 U21421 ( .B1(n19316), .B2(n19756), .A(n19331), .ZN(n19297) );
  OAI21_X1 U21422 ( .B1(n19298), .B2(n19334), .A(n19297), .ZN(n19299) );
  OAI21_X1 U21423 ( .B1(n19303), .B2(n19300), .A(n19299), .ZN(n19759) );
  INV_X1 U21424 ( .A(n19300), .ZN(n19307) );
  OAI21_X1 U21425 ( .B1(n19301), .B2(n19756), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19302) );
  OAI21_X1 U21426 ( .B1(n19303), .B2(n19307), .A(n19302), .ZN(n19758) );
  AOI22_X1 U21427 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19759), .B1(
        n19345), .B2(n19758), .ZN(n19304) );
  OAI211_X1 U21428 ( .C1(n19341), .C2(n19767), .A(n19305), .B(n19304), .ZN(
        P2_U3079) );
  NOR2_X2 U21429 ( .A1(n19315), .A2(n19306), .ZN(n19771) );
  INV_X1 U21430 ( .A(n19771), .ZN(n19497) );
  NOR2_X1 U21431 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19307), .ZN(
        n19762) );
  OAI21_X1 U21432 ( .B1(n19310), .B2(n19762), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19309) );
  OR2_X1 U21433 ( .A1(n19308), .A2(n19322), .ZN(n19313) );
  NAND2_X1 U21434 ( .A1(n19309), .A2(n19313), .ZN(n19763) );
  AOI22_X1 U21435 ( .A1(n19763), .A2(n19345), .B1(n19342), .B2(n19762), .ZN(
        n19321) );
  INV_X1 U21436 ( .A(n19310), .ZN(n19312) );
  INV_X1 U21437 ( .A(n19762), .ZN(n19311) );
  OAI21_X1 U21438 ( .B1(n19312), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n19311), 
        .ZN(n19318) );
  OAI21_X1 U21439 ( .B1(n19315), .B2(n19314), .A(n19313), .ZN(n19317) );
  MUX2_X1 U21440 ( .A(n19318), .B(n19317), .S(n19316), .Z(n19319) );
  NAND2_X1 U21441 ( .A1(n19319), .A2(n19331), .ZN(n19764) );
  AOI22_X1 U21442 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19764), .B1(
        n19494), .B2(n19344), .ZN(n19320) );
  OAI211_X1 U21443 ( .C1(n19341), .C2(n19497), .A(n19321), .B(n19320), .ZN(
        P2_U3071) );
  NOR2_X1 U21444 ( .A1(n19322), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19337) );
  INV_X1 U21445 ( .A(n19337), .ZN(n19327) );
  NOR2_X1 U21446 ( .A1(n19323), .A2(n19327), .ZN(n19769) );
  OAI21_X1 U21447 ( .B1(n19324), .B2(n19769), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19325) );
  OAI21_X1 U21448 ( .B1(n19327), .B2(n19326), .A(n19325), .ZN(n19770) );
  AOI22_X1 U21449 ( .A1(n19770), .A2(n19345), .B1(n19342), .B2(n19769), .ZN(
        n19340) );
  INV_X1 U21450 ( .A(n19328), .ZN(n19330) );
  NOR2_X1 U21451 ( .A1(n19330), .A2(n19329), .ZN(n19338) );
  OAI21_X1 U21452 ( .B1(n19332), .B2(n19769), .A(n19331), .ZN(n19333) );
  OAI21_X1 U21453 ( .B1(n19335), .B2(n19334), .A(n19333), .ZN(n19336) );
  OAI21_X1 U21454 ( .B1(n19338), .B2(n19337), .A(n19336), .ZN(n19772) );
  AOI22_X1 U21455 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19772), .B1(
        n19771), .B2(n19344), .ZN(n19339) );
  OAI211_X1 U21456 ( .C1(n19341), .C2(n19775), .A(n19340), .B(n19339), .ZN(
        P2_U3063) );
  AOI22_X1 U21457 ( .A1(n19343), .A2(n19784), .B1(n19778), .B2(n19342), .ZN(
        n19347) );
  AOI22_X1 U21458 ( .A1(n19345), .A2(n19781), .B1(n19779), .B2(n19344), .ZN(
        n19346) );
  OAI211_X1 U21459 ( .C1(n19788), .C2(n19348), .A(n19347), .B(n19346), .ZN(
        P2_U3055) );
  AOI22_X1 U21460 ( .A1(n19653), .A2(n19349), .B1(P2_EAX_REG_22__SCAN_IN), 
        .B2(n19652), .ZN(n19355) );
  AOI22_X1 U21461 ( .A1(n19655), .A2(BUF2_REG_22__SCAN_IN), .B1(n19654), .B2(
        BUF1_REG_22__SCAN_IN), .ZN(n19354) );
  INV_X1 U21462 ( .A(n19350), .ZN(n19352) );
  AOI22_X1 U21463 ( .A1(n19352), .A2(n19549), .B1(n19548), .B2(n19351), .ZN(
        n19353) );
  NAND3_X1 U21464 ( .A1(n19355), .A2(n19354), .A3(n19353), .ZN(P2_U2897) );
  AOI22_X1 U21465 ( .A1(n19556), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(
        P2_EAX_REG_22__SCAN_IN), .B2(n19667), .ZN(n19356) );
  OAI21_X1 U21466 ( .B1(n19358), .B2(n19670), .A(n19356), .ZN(P2_U2958) );
  AOI22_X1 U21467 ( .A1(n19556), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n19667), 
        .B2(P2_EAX_REG_6__SCAN_IN), .ZN(n19357) );
  OAI21_X1 U21468 ( .B1(n19358), .B2(n19670), .A(n19357), .ZN(P2_U2973) );
  NOR2_X2 U21469 ( .A1(n19358), .A2(n19673), .ZN(n19396) );
  NOR2_X2 U21470 ( .A1(n12828), .A2(n19675), .ZN(n19394) );
  AOI22_X1 U21471 ( .A1(n19678), .A2(n19396), .B1(n19677), .B2(n19394), .ZN(
        n19361) );
  OAI22_X2 U21472 ( .A1(n20079), .A2(n19681), .B1(n19359), .B2(n19679), .ZN(
        n19395) );
  AOI22_X1 U21473 ( .A1(BUF2_REG_30__SCAN_IN), .A2(n19671), .B1(
        BUF1_REG_30__SCAN_IN), .B2(n19672), .ZN(n19393) );
  INV_X1 U21474 ( .A(n19393), .ZN(n19397) );
  AOI22_X1 U21475 ( .A1(n19784), .A2(n19395), .B1(n19687), .B2(n19397), .ZN(
        n19360) );
  OAI211_X1 U21476 ( .C1(n19610), .C2(n15118), .A(n19361), .B(n19360), .ZN(
        P2_U3174) );
  INV_X1 U21477 ( .A(n19396), .ZN(n19384) );
  AOI22_X1 U21478 ( .A1(n19397), .A2(n19695), .B1(n19686), .B2(n19394), .ZN(
        n19363) );
  AOI22_X1 U21479 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n19688), .B1(
        n19687), .B2(n19395), .ZN(n19362) );
  OAI211_X1 U21480 ( .C1(n19384), .C2(n19691), .A(n19363), .B(n19362), .ZN(
        P2_U3166) );
  AOI22_X1 U21481 ( .A1(n19693), .A2(n19396), .B1(n19394), .B2(n19692), .ZN(
        n19365) );
  AOI22_X1 U21482 ( .A1(n19395), .A2(n19695), .B1(
        P2_INSTQUEUE_REG_13__6__SCAN_IN), .B2(n19694), .ZN(n19364) );
  OAI211_X1 U21483 ( .C1(n19393), .C2(n19698), .A(n19365), .B(n19364), .ZN(
        P2_U3158) );
  AOI22_X1 U21484 ( .A1(n19700), .A2(n19396), .B1(n19394), .B2(n19699), .ZN(
        n19367) );
  AOI22_X1 U21485 ( .A1(n19702), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n19701), .B2(n19395), .ZN(n19366) );
  OAI211_X1 U21486 ( .C1(n19393), .C2(n19710), .A(n19367), .B(n19366), .ZN(
        P2_U3150) );
  AOI22_X1 U21487 ( .A1(n19706), .A2(n19396), .B1(n19394), .B2(n19705), .ZN(
        n19370) );
  AOI22_X1 U21488 ( .A1(n19368), .A2(n19395), .B1(n19712), .B2(n19397), .ZN(
        n19369) );
  OAI211_X1 U21489 ( .C1(n19422), .C2(n13161), .A(n19370), .B(n19369), .ZN(
        P2_U3142) );
  AOI22_X1 U21490 ( .A1(n19397), .A2(n19718), .B1(n19711), .B2(n19394), .ZN(
        n19372) );
  AOI22_X1 U21491 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19713), .B1(
        n19712), .B2(n19395), .ZN(n19371) );
  OAI211_X1 U21492 ( .C1(n19716), .C2(n19384), .A(n19372), .B(n19371), .ZN(
        P2_U3134) );
  AOI22_X1 U21493 ( .A1(n19397), .A2(n19724), .B1(n19717), .B2(n19394), .ZN(
        n19374) );
  AOI22_X1 U21494 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n11085), .B1(
        n19718), .B2(n19395), .ZN(n19373) );
  OAI211_X1 U21495 ( .C1(n19722), .C2(n19384), .A(n19374), .B(n19373), .ZN(
        P2_U3126) );
  AOI22_X1 U21496 ( .A1(n19395), .A2(n19724), .B1(n19723), .B2(n19394), .ZN(
        n19376) );
  AOI22_X1 U21497 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19726), .B1(
        n19396), .B2(n19725), .ZN(n19375) );
  OAI211_X1 U21498 ( .C1(n19393), .C2(n19735), .A(n19376), .B(n19375), .ZN(
        P2_U3118) );
  AOI22_X1 U21499 ( .A1(n19730), .A2(n19396), .B1(n19729), .B2(n19394), .ZN(
        n19378) );
  AOI22_X1 U21500 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19732), .B1(
        n19625), .B2(n19395), .ZN(n19377) );
  OAI211_X1 U21501 ( .C1(n19393), .C2(n19741), .A(n19378), .B(n19377), .ZN(
        P2_U3110) );
  INV_X1 U21502 ( .A(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n19381) );
  AOI22_X1 U21503 ( .A1(n19737), .A2(n19396), .B1(n19394), .B2(n19736), .ZN(
        n19380) );
  AOI22_X1 U21504 ( .A1(n19731), .A2(n19395), .B1(n19743), .B2(n19397), .ZN(
        n19379) );
  OAI211_X1 U21505 ( .C1(n19631), .C2(n19381), .A(n19380), .B(n19379), .ZN(
        P2_U3102) );
  AOI22_X1 U21506 ( .A1(n19397), .A2(n19750), .B1(n19742), .B2(n19394), .ZN(
        n19383) );
  AOI22_X1 U21507 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19744), .B1(
        n19743), .B2(n19395), .ZN(n19382) );
  OAI211_X1 U21508 ( .C1(n19748), .C2(n19384), .A(n19383), .B(n19382), .ZN(
        P2_U3094) );
  AOI22_X1 U21509 ( .A1(n19395), .A2(n19750), .B1(n19749), .B2(n19394), .ZN(
        n19386) );
  AOI22_X1 U21510 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19752), .B1(
        n19396), .B2(n19751), .ZN(n19385) );
  OAI211_X1 U21511 ( .C1(n19393), .C2(n19755), .A(n19386), .B(n19385), .ZN(
        P2_U3086) );
  AOI22_X1 U21512 ( .A1(n19395), .A2(n19757), .B1(n19756), .B2(n19394), .ZN(
        n19388) );
  AOI22_X1 U21513 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19759), .B1(
        n19396), .B2(n19758), .ZN(n19387) );
  OAI211_X1 U21514 ( .C1(n19393), .C2(n19767), .A(n19388), .B(n19387), .ZN(
        P2_U3078) );
  AOI22_X1 U21515 ( .A1(n19763), .A2(n19396), .B1(n19394), .B2(n19762), .ZN(
        n19390) );
  AOI22_X1 U21516 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19764), .B1(
        n19494), .B2(n19395), .ZN(n19389) );
  OAI211_X1 U21517 ( .C1(n19393), .C2(n19497), .A(n19390), .B(n19389), .ZN(
        P2_U3070) );
  AOI22_X1 U21518 ( .A1(n19770), .A2(n19396), .B1(n19394), .B2(n19769), .ZN(
        n19392) );
  AOI22_X1 U21519 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19772), .B1(
        n19771), .B2(n19395), .ZN(n19391) );
  OAI211_X1 U21520 ( .C1(n19393), .C2(n19775), .A(n19392), .B(n19391), .ZN(
        P2_U3062) );
  AOI22_X1 U21521 ( .A1(n19395), .A2(n19779), .B1(n19778), .B2(n19394), .ZN(
        n19399) );
  AOI22_X1 U21522 ( .A1(n19784), .A2(n19397), .B1(n19396), .B2(n19781), .ZN(
        n19398) );
  OAI211_X1 U21523 ( .C1(n19788), .C2(n19400), .A(n19399), .B(n19398), .ZN(
        P2_U3054) );
  OAI22_X1 U21524 ( .A1(n19403), .A2(n19413), .B1(n19402), .B2(n19401), .ZN(
        n19404) );
  INV_X1 U21525 ( .A(n19404), .ZN(n19408) );
  OR3_X1 U21526 ( .A1(n19406), .A2(n19405), .A3(n19659), .ZN(n19407) );
  OAI211_X1 U21527 ( .C1(n19410), .C2(n19409), .A(n19408), .B(n19407), .ZN(
        P2_U2914) );
  AOI22_X1 U21528 ( .A1(n19556), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n19667), 
        .B2(P2_EAX_REG_21__SCAN_IN), .ZN(n19411) );
  OAI21_X1 U21529 ( .B1(n19413), .B2(n19670), .A(n19411), .ZN(P2_U2957) );
  AOI22_X1 U21530 ( .A1(n19556), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n19667), 
        .B2(P2_EAX_REG_5__SCAN_IN), .ZN(n19412) );
  OAI21_X1 U21531 ( .B1(n19413), .B2(n19670), .A(n19412), .ZN(P2_U2972) );
  AOI22_X1 U21532 ( .A1(n19678), .A2(n19448), .B1(n19677), .B2(n19447), .ZN(
        n19415) );
  INV_X1 U21533 ( .A(n19610), .ZN(n19682) );
  AOI22_X1 U21534 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n19682), .B1(
        n19687), .B2(n19437), .ZN(n19414) );
  OAI211_X1 U21535 ( .C1(n19431), .C2(n19562), .A(n19415), .B(n19414), .ZN(
        P2_U3173) );
  INV_X1 U21536 ( .A(n19448), .ZN(n19440) );
  AOI22_X1 U21537 ( .A1(n19437), .A2(n19695), .B1(n19447), .B2(n19686), .ZN(
        n19417) );
  AOI22_X1 U21538 ( .A1(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n19688), .B1(
        n19687), .B2(n19449), .ZN(n19416) );
  OAI211_X1 U21539 ( .C1(n19440), .C2(n19691), .A(n19417), .B(n19416), .ZN(
        P2_U3165) );
  AOI22_X1 U21540 ( .A1(n19693), .A2(n19448), .B1(n19447), .B2(n19692), .ZN(
        n19419) );
  AOI22_X1 U21541 ( .A1(n19449), .A2(n19695), .B1(n19694), .B2(
        P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n19418) );
  OAI211_X1 U21542 ( .C1(n19452), .C2(n19698), .A(n19419), .B(n19418), .ZN(
        P2_U3157) );
  AOI22_X1 U21543 ( .A1(n19700), .A2(n19448), .B1(n19447), .B2(n19699), .ZN(
        n19421) );
  AOI22_X1 U21544 ( .A1(n19702), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n19701), .B2(n19449), .ZN(n19420) );
  OAI211_X1 U21545 ( .C1(n19452), .C2(n19710), .A(n19421), .B(n19420), .ZN(
        P2_U3149) );
  AOI22_X1 U21546 ( .A1(n19706), .A2(n19448), .B1(n19447), .B2(n19705), .ZN(
        n19424) );
  AOI22_X1 U21547 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19707), .B1(
        n19712), .B2(n19437), .ZN(n19423) );
  OAI211_X1 U21548 ( .C1(n19431), .C2(n19710), .A(n19424), .B(n19423), .ZN(
        P2_U3141) );
  AOI22_X1 U21549 ( .A1(n19449), .A2(n19712), .B1(n19447), .B2(n19711), .ZN(
        n19426) );
  AOI22_X1 U21550 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19713), .B1(
        n19718), .B2(n19437), .ZN(n19425) );
  OAI211_X1 U21551 ( .C1(n19716), .C2(n19440), .A(n19426), .B(n19425), .ZN(
        P2_U3133) );
  AOI22_X1 U21552 ( .A1(n19437), .A2(n19724), .B1(n19447), .B2(n19717), .ZN(
        n19428) );
  AOI22_X1 U21553 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n11085), .B1(
        n19718), .B2(n19449), .ZN(n19427) );
  OAI211_X1 U21554 ( .C1(n19722), .C2(n19440), .A(n19428), .B(n19427), .ZN(
        P2_U3125) );
  AOI22_X1 U21555 ( .A1(n19437), .A2(n19625), .B1(n19447), .B2(n19723), .ZN(
        n19430) );
  AOI22_X1 U21556 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19726), .B1(
        n19448), .B2(n19725), .ZN(n19429) );
  OAI211_X1 U21557 ( .C1(n19431), .C2(n19577), .A(n19430), .B(n19429), .ZN(
        P2_U3117) );
  AOI22_X1 U21558 ( .A1(n19730), .A2(n19448), .B1(n19447), .B2(n19729), .ZN(
        n19433) );
  AOI22_X1 U21559 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19732), .B1(
        n19625), .B2(n19449), .ZN(n19432) );
  OAI211_X1 U21560 ( .C1(n19452), .C2(n19741), .A(n19433), .B(n19432), .ZN(
        P2_U3109) );
  AOI22_X1 U21561 ( .A1(n19737), .A2(n19448), .B1(n19447), .B2(n19736), .ZN(
        n19435) );
  AOI22_X1 U21562 ( .A1(n19743), .A2(n19437), .B1(n19731), .B2(n19449), .ZN(
        n19434) );
  OAI211_X1 U21563 ( .C1(n19631), .C2(n19436), .A(n19435), .B(n19434), .ZN(
        P2_U3101) );
  AOI22_X1 U21564 ( .A1(n19437), .A2(n19750), .B1(n19447), .B2(n19742), .ZN(
        n19439) );
  AOI22_X1 U21565 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19744), .B1(
        n19743), .B2(n19449), .ZN(n19438) );
  OAI211_X1 U21566 ( .C1(n19748), .C2(n19440), .A(n19439), .B(n19438), .ZN(
        P2_U3093) );
  AOI22_X1 U21567 ( .A1(n19449), .A2(n19750), .B1(n19447), .B2(n19749), .ZN(
        n19442) );
  AOI22_X1 U21568 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19752), .B1(
        n19448), .B2(n19751), .ZN(n19441) );
  OAI211_X1 U21569 ( .C1(n19452), .C2(n19755), .A(n19442), .B(n19441), .ZN(
        P2_U3085) );
  AOI22_X1 U21570 ( .A1(n19449), .A2(n19757), .B1(n19447), .B2(n19756), .ZN(
        n19444) );
  AOI22_X1 U21571 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19759), .B1(
        n19448), .B2(n19758), .ZN(n19443) );
  OAI211_X1 U21572 ( .C1(n19452), .C2(n19767), .A(n19444), .B(n19443), .ZN(
        P2_U3077) );
  AOI22_X1 U21573 ( .A1(n19763), .A2(n19448), .B1(n19447), .B2(n19762), .ZN(
        n19446) );
  AOI22_X1 U21574 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19764), .B1(
        n19494), .B2(n19449), .ZN(n19445) );
  OAI211_X1 U21575 ( .C1(n19452), .C2(n19497), .A(n19446), .B(n19445), .ZN(
        P2_U3069) );
  AOI22_X1 U21576 ( .A1(n19770), .A2(n19448), .B1(n19447), .B2(n19769), .ZN(
        n19451) );
  AOI22_X1 U21577 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19772), .B1(
        n19771), .B2(n19449), .ZN(n19450) );
  OAI211_X1 U21578 ( .C1(n19452), .C2(n19775), .A(n19451), .B(n19450), .ZN(
        P2_U3061) );
  AOI22_X1 U21579 ( .A1(n19653), .A2(n19453), .B1(n19652), .B2(
        P2_EAX_REG_20__SCAN_IN), .ZN(n19459) );
  AOI22_X1 U21580 ( .A1(n19655), .A2(BUF2_REG_20__SCAN_IN), .B1(n19654), .B2(
        BUF1_REG_20__SCAN_IN), .ZN(n19458) );
  INV_X1 U21581 ( .A(n19454), .ZN(n19456) );
  AOI22_X1 U21582 ( .A1(n19456), .A2(n19549), .B1(n19548), .B2(n19455), .ZN(
        n19457) );
  NAND3_X1 U21583 ( .A1(n19459), .A2(n19458), .A3(n19457), .ZN(P2_U2899) );
  AOI22_X1 U21584 ( .A1(n19556), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(
        P2_EAX_REG_20__SCAN_IN), .B2(n19667), .ZN(n19460) );
  OAI21_X1 U21585 ( .B1(n19462), .B2(n19670), .A(n19460), .ZN(P2_U2956) );
  AOI22_X1 U21586 ( .A1(n19556), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n19667), 
        .B2(P2_EAX_REG_4__SCAN_IN), .ZN(n19461) );
  OAI21_X1 U21587 ( .B1(n19462), .B2(n19670), .A(n19461), .ZN(P2_U2971) );
  INV_X1 U21588 ( .A(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n19467) );
  NOR2_X2 U21589 ( .A1(n19464), .A2(n19675), .ZN(n19501) );
  AOI22_X1 U21590 ( .A1(n19678), .A2(n19463), .B1(n19677), .B2(n19501), .ZN(
        n19466) );
  AOI22_X1 U21591 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n19672), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n19671), .ZN(n19486) );
  AOI22_X1 U21592 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n19671), .B1(
        BUF1_REG_28__SCAN_IN), .B2(n19672), .ZN(n19500) );
  AOI22_X1 U21593 ( .A1(n19784), .A2(n19502), .B1(n19687), .B2(n19503), .ZN(
        n19465) );
  OAI211_X1 U21594 ( .C1(n19610), .C2(n19467), .A(n19466), .B(n19465), .ZN(
        P2_U3172) );
  INV_X1 U21595 ( .A(n19463), .ZN(n19489) );
  AOI22_X1 U21596 ( .A1(n19502), .A2(n19687), .B1(n19686), .B2(n19501), .ZN(
        n19469) );
  AOI22_X1 U21597 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n19688), .B1(
        n19695), .B2(n19503), .ZN(n19468) );
  OAI211_X1 U21598 ( .C1(n19489), .C2(n19691), .A(n19469), .B(n19468), .ZN(
        P2_U3164) );
  AOI22_X1 U21599 ( .A1(n19693), .A2(n19463), .B1(n19501), .B2(n19692), .ZN(
        n19471) );
  AOI22_X1 U21600 ( .A1(n19502), .A2(n19695), .B1(n19694), .B2(
        P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n19470) );
  OAI211_X1 U21601 ( .C1(n19500), .C2(n19698), .A(n19471), .B(n19470), .ZN(
        P2_U3156) );
  AOI22_X1 U21602 ( .A1(n19700), .A2(n19463), .B1(n19501), .B2(n19699), .ZN(
        n19473) );
  AOI22_X1 U21603 ( .A1(n19702), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n19701), .B2(n19502), .ZN(n19472) );
  OAI211_X1 U21604 ( .C1(n19500), .C2(n19710), .A(n19473), .B(n19472), .ZN(
        P2_U3148) );
  AOI22_X1 U21605 ( .A1(n19706), .A2(n19463), .B1(n19501), .B2(n19705), .ZN(
        n19475) );
  AOI22_X1 U21606 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19707), .B1(
        n19712), .B2(n19503), .ZN(n19474) );
  OAI211_X1 U21607 ( .C1(n19486), .C2(n19710), .A(n19475), .B(n19474), .ZN(
        P2_U3140) );
  AOI22_X1 U21608 ( .A1(n19503), .A2(n19718), .B1(n19711), .B2(n19501), .ZN(
        n19477) );
  AOI22_X1 U21609 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19713), .B1(
        n19712), .B2(n19502), .ZN(n19476) );
  OAI211_X1 U21610 ( .C1(n19716), .C2(n19489), .A(n19477), .B(n19476), .ZN(
        P2_U3132) );
  AOI22_X1 U21611 ( .A1(n19503), .A2(n19724), .B1(n19717), .B2(n19501), .ZN(
        n19479) );
  AOI22_X1 U21612 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n11085), .B1(
        n19718), .B2(n19502), .ZN(n19478) );
  OAI211_X1 U21613 ( .C1(n19722), .C2(n19489), .A(n19479), .B(n19478), .ZN(
        P2_U3124) );
  AOI22_X1 U21614 ( .A1(n19503), .A2(n19625), .B1(n19723), .B2(n19501), .ZN(
        n19481) );
  AOI22_X1 U21615 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19726), .B1(
        n19463), .B2(n19725), .ZN(n19480) );
  OAI211_X1 U21616 ( .C1(n19486), .C2(n19577), .A(n19481), .B(n19480), .ZN(
        P2_U3116) );
  AOI22_X1 U21617 ( .A1(n19730), .A2(n19463), .B1(n19729), .B2(n19501), .ZN(
        n19483) );
  AOI22_X1 U21618 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19732), .B1(
        n19625), .B2(n19502), .ZN(n19482) );
  OAI211_X1 U21619 ( .C1(n19500), .C2(n19741), .A(n19483), .B(n19482), .ZN(
        P2_U3108) );
  AOI22_X1 U21620 ( .A1(n19737), .A2(n19463), .B1(n19501), .B2(n19736), .ZN(
        n19485) );
  INV_X1 U21621 ( .A(n19631), .ZN(n19738) );
  AOI22_X1 U21622 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19738), .B1(
        n19743), .B2(n19503), .ZN(n19484) );
  OAI211_X1 U21623 ( .C1(n19486), .C2(n19741), .A(n19485), .B(n19484), .ZN(
        P2_U3100) );
  AOI22_X1 U21624 ( .A1(n19503), .A2(n19750), .B1(n19742), .B2(n19501), .ZN(
        n19488) );
  AOI22_X1 U21625 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19744), .B1(
        n19743), .B2(n19502), .ZN(n19487) );
  OAI211_X1 U21626 ( .C1(n19748), .C2(n19489), .A(n19488), .B(n19487), .ZN(
        P2_U3092) );
  AOI22_X1 U21627 ( .A1(n19502), .A2(n19750), .B1(n19749), .B2(n19501), .ZN(
        n19491) );
  AOI22_X1 U21628 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19752), .B1(
        n19463), .B2(n19751), .ZN(n19490) );
  OAI211_X1 U21629 ( .C1(n19500), .C2(n19755), .A(n19491), .B(n19490), .ZN(
        P2_U3084) );
  AOI22_X1 U21630 ( .A1(n19502), .A2(n19757), .B1(n19756), .B2(n19501), .ZN(
        n19493) );
  AOI22_X1 U21631 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19759), .B1(
        n19463), .B2(n19758), .ZN(n19492) );
  OAI211_X1 U21632 ( .C1(n19500), .C2(n19767), .A(n19493), .B(n19492), .ZN(
        P2_U3076) );
  AOI22_X1 U21633 ( .A1(n19763), .A2(n19463), .B1(n19501), .B2(n19762), .ZN(
        n19496) );
  AOI22_X1 U21634 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19764), .B1(
        n19494), .B2(n19502), .ZN(n19495) );
  OAI211_X1 U21635 ( .C1(n19500), .C2(n19497), .A(n19496), .B(n19495), .ZN(
        P2_U3068) );
  AOI22_X1 U21636 ( .A1(n19770), .A2(n19463), .B1(n19501), .B2(n19769), .ZN(
        n19499) );
  AOI22_X1 U21637 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19772), .B1(
        n19771), .B2(n19502), .ZN(n19498) );
  OAI211_X1 U21638 ( .C1(n19500), .C2(n19775), .A(n19499), .B(n19498), .ZN(
        P2_U3060) );
  AOI22_X1 U21639 ( .A1(n19502), .A2(n19779), .B1(n19778), .B2(n19501), .ZN(
        n19505) );
  AOI22_X1 U21640 ( .A1(n19784), .A2(n19503), .B1(n19463), .B2(n19781), .ZN(
        n19504) );
  OAI211_X1 U21641 ( .C1(n19788), .C2(n19506), .A(n19505), .B(n19504), .ZN(
        P2_U3052) );
  AOI22_X1 U21642 ( .A1(n19556), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n19667), 
        .B2(P2_EAX_REG_19__SCAN_IN), .ZN(n19507) );
  OAI21_X1 U21643 ( .B1(n19509), .B2(n19670), .A(n19507), .ZN(P2_U2955) );
  AOI22_X1 U21644 ( .A1(n19556), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(
        P2_EAX_REG_3__SCAN_IN), .B2(n19667), .ZN(n19508) );
  OAI21_X1 U21645 ( .B1(n19509), .B2(n19670), .A(n19508), .ZN(P2_U2970) );
  AOI22_X1 U21646 ( .A1(n19678), .A2(n16677), .B1(n19677), .B2(n19541), .ZN(
        n19511) );
  AOI22_X1 U21647 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n19682), .B1(
        n19687), .B2(n19537), .ZN(n19510) );
  OAI211_X1 U21648 ( .C1(n19540), .C2(n19562), .A(n19511), .B(n19510), .ZN(
        P2_U3171) );
  AOI22_X1 U21649 ( .A1(n19542), .A2(n19687), .B1(n19541), .B2(n19686), .ZN(
        n19513) );
  AOI22_X1 U21650 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n19688), .B1(
        n19695), .B2(n19537), .ZN(n19512) );
  OAI211_X1 U21651 ( .C1(n19532), .C2(n19691), .A(n19513), .B(n19512), .ZN(
        P2_U3163) );
  AOI22_X1 U21652 ( .A1(n19693), .A2(n16677), .B1(n19541), .B2(n19692), .ZN(
        n19515) );
  AOI22_X1 U21653 ( .A1(n19542), .A2(n19695), .B1(n19694), .B2(
        P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n19514) );
  OAI211_X1 U21654 ( .C1(n19545), .C2(n19698), .A(n19515), .B(n19514), .ZN(
        P2_U3155) );
  AOI22_X1 U21655 ( .A1(n19700), .A2(n16677), .B1(n19541), .B2(n19699), .ZN(
        n19517) );
  AOI22_X1 U21656 ( .A1(n19702), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n19701), .B2(n19542), .ZN(n19516) );
  OAI211_X1 U21657 ( .C1(n19545), .C2(n19710), .A(n19517), .B(n19516), .ZN(
        P2_U3147) );
  AOI22_X1 U21658 ( .A1(n19706), .A2(n16677), .B1(n19541), .B2(n19705), .ZN(
        n19519) );
  AOI22_X1 U21659 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19707), .B1(
        n19712), .B2(n19537), .ZN(n19518) );
  OAI211_X1 U21660 ( .C1(n19540), .C2(n19710), .A(n19519), .B(n19518), .ZN(
        P2_U3139) );
  AOI22_X1 U21661 ( .A1(n19537), .A2(n19718), .B1(n19541), .B2(n19711), .ZN(
        n19521) );
  AOI22_X1 U21662 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19713), .B1(
        n19712), .B2(n19542), .ZN(n19520) );
  OAI211_X1 U21663 ( .C1(n19716), .C2(n19532), .A(n19521), .B(n19520), .ZN(
        P2_U3131) );
  AOI22_X1 U21664 ( .A1(n19537), .A2(n19724), .B1(n19541), .B2(n19717), .ZN(
        n19523) );
  AOI22_X1 U21665 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n11085), .B1(
        n19718), .B2(n19542), .ZN(n19522) );
  OAI211_X1 U21666 ( .C1(n19722), .C2(n19532), .A(n19523), .B(n19522), .ZN(
        P2_U3123) );
  AOI22_X1 U21667 ( .A1(n19537), .A2(n19625), .B1(n19541), .B2(n19723), .ZN(
        n19525) );
  AOI22_X1 U21668 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19726), .B1(
        n16677), .B2(n19725), .ZN(n19524) );
  OAI211_X1 U21669 ( .C1(n19540), .C2(n19577), .A(n19525), .B(n19524), .ZN(
        P2_U3115) );
  AOI22_X1 U21670 ( .A1(n19730), .A2(n16677), .B1(n19541), .B2(n19729), .ZN(
        n19527) );
  AOI22_X1 U21671 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19732), .B1(
        n19625), .B2(n19542), .ZN(n19526) );
  OAI211_X1 U21672 ( .C1(n19545), .C2(n19741), .A(n19527), .B(n19526), .ZN(
        P2_U3107) );
  AOI22_X1 U21673 ( .A1(n19737), .A2(n16677), .B1(n19541), .B2(n19736), .ZN(
        n19529) );
  AOI22_X1 U21674 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19738), .B1(
        n19743), .B2(n19537), .ZN(n19528) );
  OAI211_X1 U21675 ( .C1(n19540), .C2(n19741), .A(n19529), .B(n19528), .ZN(
        P2_U3099) );
  AOI22_X1 U21676 ( .A1(n19537), .A2(n19750), .B1(n19541), .B2(n19742), .ZN(
        n19531) );
  AOI22_X1 U21677 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19744), .B1(
        n19743), .B2(n19542), .ZN(n19530) );
  OAI211_X1 U21678 ( .C1(n19748), .C2(n19532), .A(n19531), .B(n19530), .ZN(
        P2_U3091) );
  AOI22_X1 U21679 ( .A1(n19542), .A2(n19750), .B1(n19541), .B2(n19749), .ZN(
        n19534) );
  AOI22_X1 U21680 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19752), .B1(
        n16677), .B2(n19751), .ZN(n19533) );
  OAI211_X1 U21681 ( .C1(n19545), .C2(n19755), .A(n19534), .B(n19533), .ZN(
        P2_U3083) );
  AOI22_X1 U21682 ( .A1(n19542), .A2(n19757), .B1(n19541), .B2(n19756), .ZN(
        n19536) );
  AOI22_X1 U21683 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19759), .B1(
        n16677), .B2(n19758), .ZN(n19535) );
  OAI211_X1 U21684 ( .C1(n19545), .C2(n19767), .A(n19536), .B(n19535), .ZN(
        P2_U3075) );
  AOI22_X1 U21685 ( .A1(n19763), .A2(n16677), .B1(n19541), .B2(n19762), .ZN(
        n19539) );
  AOI22_X1 U21686 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19764), .B1(
        n19771), .B2(n19537), .ZN(n19538) );
  OAI211_X1 U21687 ( .C1(n19540), .C2(n19767), .A(n19539), .B(n19538), .ZN(
        P2_U3067) );
  AOI22_X1 U21688 ( .A1(n19770), .A2(n16677), .B1(n19541), .B2(n19769), .ZN(
        n19544) );
  AOI22_X1 U21689 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19772), .B1(
        n19771), .B2(n19542), .ZN(n19543) );
  OAI211_X1 U21690 ( .C1(n19545), .C2(n19775), .A(n19544), .B(n19543), .ZN(
        P2_U3059) );
  AOI22_X1 U21691 ( .A1(n19653), .A2(n19554), .B1(n19652), .B2(
        P2_EAX_REG_18__SCAN_IN), .ZN(n19553) );
  AOI22_X1 U21692 ( .A1(n19655), .A2(BUF2_REG_18__SCAN_IN), .B1(n19654), .B2(
        BUF1_REG_18__SCAN_IN), .ZN(n19552) );
  INV_X1 U21693 ( .A(n19546), .ZN(n19550) );
  AOI22_X1 U21694 ( .A1(n19550), .A2(n19549), .B1(n19548), .B2(n19547), .ZN(
        n19551) );
  NAND3_X1 U21695 ( .A1(n19553), .A2(n19552), .A3(n19551), .ZN(P2_U2901) );
  INV_X1 U21696 ( .A(n19554), .ZN(n19558) );
  AOI22_X1 U21697 ( .A1(n19556), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(
        P2_EAX_REG_18__SCAN_IN), .B2(n19667), .ZN(n19555) );
  OAI21_X1 U21698 ( .B1(n19558), .B2(n19670), .A(n19555), .ZN(P2_U2954) );
  AOI22_X1 U21699 ( .A1(n19556), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n19667), 
        .B2(P2_EAX_REG_2__SCAN_IN), .ZN(n19557) );
  OAI21_X1 U21700 ( .B1(n19558), .B2(n19670), .A(n19557), .ZN(P2_U2969) );
  AOI22_X1 U21701 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n19672), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n19671), .ZN(n19591) );
  NOR2_X2 U21702 ( .A1(n19558), .A2(n19673), .ZN(n19597) );
  NOR2_X2 U21703 ( .A1(n19559), .A2(n19675), .ZN(n19595) );
  AOI22_X1 U21704 ( .A1(n19678), .A2(n19597), .B1(n19677), .B2(n19595), .ZN(
        n19561) );
  AOI22_X1 U21705 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n19672), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n19671), .ZN(n19594) );
  AOI22_X1 U21706 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n19682), .B1(
        n19687), .B2(n19598), .ZN(n19560) );
  OAI211_X1 U21707 ( .C1(n19591), .C2(n19562), .A(n19561), .B(n19560), .ZN(
        P2_U3170) );
  INV_X1 U21708 ( .A(n19597), .ZN(n19584) );
  AOI22_X1 U21709 ( .A1(n19596), .A2(n19687), .B1(n19686), .B2(n19595), .ZN(
        n19564) );
  AOI22_X1 U21710 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n19688), .B1(
        n19695), .B2(n19598), .ZN(n19563) );
  OAI211_X1 U21711 ( .C1(n19584), .C2(n19691), .A(n19564), .B(n19563), .ZN(
        P2_U3162) );
  AOI22_X1 U21712 ( .A1(n19693), .A2(n19597), .B1(n19595), .B2(n19692), .ZN(
        n19566) );
  AOI22_X1 U21713 ( .A1(n19596), .A2(n19695), .B1(n19694), .B2(
        P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n19565) );
  OAI211_X1 U21714 ( .C1(n19594), .C2(n19698), .A(n19566), .B(n19565), .ZN(
        P2_U3154) );
  AOI22_X1 U21715 ( .A1(n19700), .A2(n19597), .B1(n19595), .B2(n19699), .ZN(
        n19568) );
  AOI22_X1 U21716 ( .A1(n19702), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n19701), .B2(n19596), .ZN(n19567) );
  OAI211_X1 U21717 ( .C1(n19594), .C2(n19710), .A(n19568), .B(n19567), .ZN(
        P2_U3146) );
  AOI22_X1 U21718 ( .A1(n19706), .A2(n19597), .B1(n19595), .B2(n19705), .ZN(
        n19570) );
  AOI22_X1 U21719 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19707), .B1(
        n19712), .B2(n19598), .ZN(n19569) );
  OAI211_X1 U21720 ( .C1(n19591), .C2(n19710), .A(n19570), .B(n19569), .ZN(
        P2_U3138) );
  AOI22_X1 U21721 ( .A1(n19596), .A2(n19712), .B1(n19711), .B2(n19595), .ZN(
        n19572) );
  AOI22_X1 U21722 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19713), .B1(
        n19718), .B2(n19598), .ZN(n19571) );
  OAI211_X1 U21723 ( .C1(n19716), .C2(n19584), .A(n19572), .B(n19571), .ZN(
        P2_U3130) );
  AOI22_X1 U21724 ( .A1(n19598), .A2(n19724), .B1(n19717), .B2(n19595), .ZN(
        n19574) );
  AOI22_X1 U21725 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n11085), .B1(
        n19718), .B2(n19596), .ZN(n19573) );
  OAI211_X1 U21726 ( .C1(n19722), .C2(n19584), .A(n19574), .B(n19573), .ZN(
        P2_U3122) );
  AOI22_X1 U21727 ( .A1(n19598), .A2(n19625), .B1(n19723), .B2(n19595), .ZN(
        n19576) );
  AOI22_X1 U21728 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19726), .B1(
        n19597), .B2(n19725), .ZN(n19575) );
  OAI211_X1 U21729 ( .C1(n19591), .C2(n19577), .A(n19576), .B(n19575), .ZN(
        P2_U3114) );
  AOI22_X1 U21730 ( .A1(n19730), .A2(n19597), .B1(n19729), .B2(n19595), .ZN(
        n19579) );
  AOI22_X1 U21731 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19732), .B1(
        n19731), .B2(n19598), .ZN(n19578) );
  OAI211_X1 U21732 ( .C1(n19591), .C2(n19735), .A(n19579), .B(n19578), .ZN(
        P2_U3106) );
  AOI22_X1 U21733 ( .A1(n19737), .A2(n19597), .B1(n19595), .B2(n19736), .ZN(
        n19581) );
  AOI22_X1 U21734 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19738), .B1(
        n19743), .B2(n19598), .ZN(n19580) );
  OAI211_X1 U21735 ( .C1(n19591), .C2(n19741), .A(n19581), .B(n19580), .ZN(
        P2_U3098) );
  AOI22_X1 U21736 ( .A1(n19598), .A2(n19750), .B1(n19742), .B2(n19595), .ZN(
        n19583) );
  AOI22_X1 U21737 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19744), .B1(
        n19743), .B2(n19596), .ZN(n19582) );
  OAI211_X1 U21738 ( .C1(n19748), .C2(n19584), .A(n19583), .B(n19582), .ZN(
        P2_U3090) );
  AOI22_X1 U21739 ( .A1(n19596), .A2(n19750), .B1(n19749), .B2(n19595), .ZN(
        n19586) );
  AOI22_X1 U21740 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19752), .B1(
        n19597), .B2(n19751), .ZN(n19585) );
  OAI211_X1 U21741 ( .C1(n19594), .C2(n19755), .A(n19586), .B(n19585), .ZN(
        P2_U3082) );
  AOI22_X1 U21742 ( .A1(n19596), .A2(n19757), .B1(n19756), .B2(n19595), .ZN(
        n19588) );
  AOI22_X1 U21743 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19759), .B1(
        n19597), .B2(n19758), .ZN(n19587) );
  OAI211_X1 U21744 ( .C1(n19594), .C2(n19767), .A(n19588), .B(n19587), .ZN(
        P2_U3074) );
  AOI22_X1 U21745 ( .A1(n19763), .A2(n19597), .B1(n19595), .B2(n19762), .ZN(
        n19590) );
  AOI22_X1 U21746 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19764), .B1(
        n19771), .B2(n19598), .ZN(n19589) );
  OAI211_X1 U21747 ( .C1(n19591), .C2(n19767), .A(n19590), .B(n19589), .ZN(
        P2_U3066) );
  AOI22_X1 U21748 ( .A1(n19770), .A2(n19597), .B1(n19595), .B2(n19769), .ZN(
        n19593) );
  AOI22_X1 U21749 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19772), .B1(
        n19771), .B2(n19596), .ZN(n19592) );
  OAI211_X1 U21750 ( .C1(n19594), .C2(n19775), .A(n19593), .B(n19592), .ZN(
        P2_U3058) );
  AOI22_X1 U21751 ( .A1(n19596), .A2(n19779), .B1(n19778), .B2(n19595), .ZN(
        n19600) );
  AOI22_X1 U21752 ( .A1(n19784), .A2(n19598), .B1(n19597), .B2(n19781), .ZN(
        n19599) );
  OAI211_X1 U21753 ( .C1(n19788), .C2(n19601), .A(n19600), .B(n19599), .ZN(
        P2_U3050) );
  AOI22_X1 U21754 ( .A1(n19668), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n19667), 
        .B2(P2_EAX_REG_17__SCAN_IN), .ZN(n19602) );
  OAI21_X1 U21755 ( .B1(n19604), .B2(n19670), .A(n19602), .ZN(P2_U2953) );
  AOI22_X1 U21756 ( .A1(n19668), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n19667), 
        .B2(P2_EAX_REG_1__SCAN_IN), .ZN(n19603) );
  OAI21_X1 U21757 ( .B1(n19604), .B2(n19670), .A(n19603), .ZN(P2_U2968) );
  NOR2_X2 U21758 ( .A1(n19604), .A2(n19673), .ZN(n19647) );
  NOR2_X2 U21759 ( .A1(n19605), .A2(n19675), .ZN(n19645) );
  AOI22_X1 U21760 ( .A1(n19678), .A2(n19647), .B1(n19677), .B2(n19645), .ZN(
        n19608) );
  OAI22_X2 U21761 ( .A1(n20069), .A2(n19681), .B1(n19606), .B2(n19679), .ZN(
        n19648) );
  AOI22_X1 U21762 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n19672), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n19671), .ZN(n19644) );
  INV_X1 U21763 ( .A(n19644), .ZN(n19646) );
  AOI22_X1 U21764 ( .A1(n19784), .A2(n19648), .B1(n19687), .B2(n19646), .ZN(
        n19607) );
  OAI211_X1 U21765 ( .C1(n19610), .C2(n19609), .A(n19608), .B(n19607), .ZN(
        P2_U3169) );
  INV_X1 U21766 ( .A(n19647), .ZN(n19634) );
  AOI22_X1 U21767 ( .A1(n19646), .A2(n19695), .B1(n19686), .B2(n19645), .ZN(
        n19612) );
  AOI22_X1 U21768 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n19688), .B1(
        n19687), .B2(n19648), .ZN(n19611) );
  OAI211_X1 U21769 ( .C1(n19634), .C2(n19691), .A(n19612), .B(n19611), .ZN(
        P2_U3161) );
  AOI22_X1 U21770 ( .A1(n19693), .A2(n19647), .B1(n19645), .B2(n19692), .ZN(
        n19614) );
  AOI22_X1 U21771 ( .A1(n19648), .A2(n19695), .B1(
        P2_INSTQUEUE_REG_13__1__SCAN_IN), .B2(n19694), .ZN(n19613) );
  OAI211_X1 U21772 ( .C1(n19644), .C2(n19698), .A(n19614), .B(n19613), .ZN(
        P2_U3153) );
  AOI22_X1 U21773 ( .A1(n19700), .A2(n19647), .B1(n19645), .B2(n19699), .ZN(
        n19616) );
  AOI22_X1 U21774 ( .A1(n19702), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n19701), .B2(n19648), .ZN(n19615) );
  OAI211_X1 U21775 ( .C1(n19644), .C2(n19710), .A(n19616), .B(n19615), .ZN(
        P2_U3145) );
  INV_X1 U21776 ( .A(n19648), .ZN(n19641) );
  AOI22_X1 U21777 ( .A1(n19706), .A2(n19647), .B1(n19645), .B2(n19705), .ZN(
        n19618) );
  AOI22_X1 U21778 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19707), .B1(
        n19712), .B2(n19646), .ZN(n19617) );
  OAI211_X1 U21779 ( .C1(n19641), .C2(n19710), .A(n19618), .B(n19617), .ZN(
        P2_U3137) );
  AOI22_X1 U21780 ( .A1(n19648), .A2(n19712), .B1(n19711), .B2(n19645), .ZN(
        n19620) );
  AOI22_X1 U21781 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19713), .B1(
        n19718), .B2(n19646), .ZN(n19619) );
  OAI211_X1 U21782 ( .C1(n19716), .C2(n19634), .A(n19620), .B(n19619), .ZN(
        P2_U3129) );
  AOI22_X1 U21783 ( .A1(n19646), .A2(n19724), .B1(n19717), .B2(n19645), .ZN(
        n19622) );
  AOI22_X1 U21784 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n11085), .B1(
        n19718), .B2(n19648), .ZN(n19621) );
  OAI211_X1 U21785 ( .C1(n19722), .C2(n19634), .A(n19622), .B(n19621), .ZN(
        P2_U3121) );
  AOI22_X1 U21786 ( .A1(n19648), .A2(n19724), .B1(n19723), .B2(n19645), .ZN(
        n19624) );
  AOI22_X1 U21787 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19726), .B1(
        n19647), .B2(n19725), .ZN(n19623) );
  OAI211_X1 U21788 ( .C1(n19644), .C2(n19735), .A(n19624), .B(n19623), .ZN(
        P2_U3113) );
  AOI22_X1 U21789 ( .A1(n19730), .A2(n19647), .B1(n19729), .B2(n19645), .ZN(
        n19627) );
  AOI22_X1 U21790 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19732), .B1(
        n19625), .B2(n19648), .ZN(n19626) );
  OAI211_X1 U21791 ( .C1(n19644), .C2(n19741), .A(n19627), .B(n19626), .ZN(
        P2_U3105) );
  AOI22_X1 U21792 ( .A1(n19737), .A2(n19647), .B1(n19645), .B2(n19736), .ZN(
        n19629) );
  AOI22_X1 U21793 ( .A1(n19731), .A2(n19648), .B1(n19743), .B2(n19646), .ZN(
        n19628) );
  OAI211_X1 U21794 ( .C1(n19631), .C2(n19630), .A(n19629), .B(n19628), .ZN(
        P2_U3097) );
  AOI22_X1 U21795 ( .A1(n19646), .A2(n19750), .B1(n19742), .B2(n19645), .ZN(
        n19633) );
  AOI22_X1 U21796 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19744), .B1(
        n19743), .B2(n19648), .ZN(n19632) );
  OAI211_X1 U21797 ( .C1(n19748), .C2(n19634), .A(n19633), .B(n19632), .ZN(
        P2_U3089) );
  AOI22_X1 U21798 ( .A1(n19648), .A2(n19750), .B1(n19749), .B2(n19645), .ZN(
        n19636) );
  AOI22_X1 U21799 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19752), .B1(
        n19647), .B2(n19751), .ZN(n19635) );
  OAI211_X1 U21800 ( .C1(n19644), .C2(n19755), .A(n19636), .B(n19635), .ZN(
        P2_U3081) );
  AOI22_X1 U21801 ( .A1(n19648), .A2(n19757), .B1(n19756), .B2(n19645), .ZN(
        n19638) );
  AOI22_X1 U21802 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19759), .B1(
        n19647), .B2(n19758), .ZN(n19637) );
  OAI211_X1 U21803 ( .C1(n19644), .C2(n19767), .A(n19638), .B(n19637), .ZN(
        P2_U3073) );
  AOI22_X1 U21804 ( .A1(n19763), .A2(n19647), .B1(n19645), .B2(n19762), .ZN(
        n19640) );
  AOI22_X1 U21805 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19764), .B1(
        n19771), .B2(n19646), .ZN(n19639) );
  OAI211_X1 U21806 ( .C1(n19641), .C2(n19767), .A(n19640), .B(n19639), .ZN(
        P2_U3065) );
  AOI22_X1 U21807 ( .A1(n19770), .A2(n19647), .B1(n19645), .B2(n19769), .ZN(
        n19643) );
  AOI22_X1 U21808 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19772), .B1(
        n19771), .B2(n19648), .ZN(n19642) );
  OAI211_X1 U21809 ( .C1(n19644), .C2(n19775), .A(n19643), .B(n19642), .ZN(
        P2_U3057) );
  AOI22_X1 U21810 ( .A1(n19646), .A2(n19784), .B1(n19778), .B2(n19645), .ZN(
        n19650) );
  AOI22_X1 U21811 ( .A1(n19779), .A2(n19648), .B1(n19647), .B2(n19781), .ZN(
        n19649) );
  OAI211_X1 U21812 ( .C1(n19788), .C2(n19651), .A(n19650), .B(n19649), .ZN(
        P2_U3049) );
  AOI22_X1 U21813 ( .A1(n19653), .A2(n19665), .B1(n19652), .B2(
        P2_EAX_REG_16__SCAN_IN), .ZN(n19664) );
  AOI22_X1 U21814 ( .A1(n19655), .A2(BUF2_REG_16__SCAN_IN), .B1(n19654), .B2(
        BUF1_REG_16__SCAN_IN), .ZN(n19663) );
  INV_X1 U21815 ( .A(n19656), .ZN(n19657) );
  OAI22_X1 U21816 ( .A1(n19660), .A2(n19659), .B1(n19658), .B2(n19657), .ZN(
        n19661) );
  INV_X1 U21817 ( .A(n19661), .ZN(n19662) );
  NAND3_X1 U21818 ( .A1(n19664), .A2(n19663), .A3(n19662), .ZN(P2_U2903) );
  INV_X1 U21819 ( .A(n19665), .ZN(n19674) );
  AOI22_X1 U21820 ( .A1(n19668), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(
        P2_EAX_REG_16__SCAN_IN), .B2(n19667), .ZN(n19666) );
  OAI21_X1 U21821 ( .B1(n19674), .B2(n19670), .A(n19666), .ZN(P2_U2952) );
  AOI22_X1 U21822 ( .A1(n19668), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n19667), 
        .B2(P2_EAX_REG_0__SCAN_IN), .ZN(n19669) );
  OAI21_X1 U21823 ( .B1(n19674), .B2(n19670), .A(n19669), .ZN(P2_U2967) );
  AOI22_X1 U21824 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n19672), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n19671), .ZN(n19776) );
  INV_X1 U21825 ( .A(n19687), .ZN(n19685) );
  NOR2_X2 U21826 ( .A1(n19674), .A2(n19673), .ZN(n19782) );
  NOR2_X2 U21827 ( .A1(n19676), .A2(n19675), .ZN(n19777) );
  AOI22_X1 U21828 ( .A1(n19678), .A2(n19782), .B1(n19677), .B2(n19777), .ZN(
        n19684) );
  OAI22_X2 U21829 ( .A1(n20067), .A2(n19681), .B1(n19680), .B2(n19679), .ZN(
        n19780) );
  AOI22_X1 U21830 ( .A1(P2_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n19682), .B1(
        n19784), .B2(n19780), .ZN(n19683) );
  OAI211_X1 U21831 ( .C1(n19776), .C2(n19685), .A(n19684), .B(n19683), .ZN(
        P2_U3168) );
  INV_X1 U21832 ( .A(n19782), .ZN(n19747) );
  INV_X1 U21833 ( .A(n19776), .ZN(n19783) );
  AOI22_X1 U21834 ( .A1(n19783), .A2(n19695), .B1(n19686), .B2(n19777), .ZN(
        n19690) );
  AOI22_X1 U21835 ( .A1(P2_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n19688), .B1(
        n19687), .B2(n19780), .ZN(n19689) );
  OAI211_X1 U21836 ( .C1(n19747), .C2(n19691), .A(n19690), .B(n19689), .ZN(
        P2_U3160) );
  AOI22_X1 U21837 ( .A1(n19693), .A2(n19782), .B1(n19777), .B2(n19692), .ZN(
        n19697) );
  AOI22_X1 U21838 ( .A1(n19780), .A2(n19695), .B1(
        P2_INSTQUEUE_REG_13__0__SCAN_IN), .B2(n19694), .ZN(n19696) );
  OAI211_X1 U21839 ( .C1(n19776), .C2(n19698), .A(n19697), .B(n19696), .ZN(
        P2_U3152) );
  AOI22_X1 U21840 ( .A1(n19700), .A2(n19782), .B1(n19777), .B2(n19699), .ZN(
        n19704) );
  AOI22_X1 U21841 ( .A1(n19702), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n19701), .B2(n19780), .ZN(n19703) );
  OAI211_X1 U21842 ( .C1(n19776), .C2(n19710), .A(n19704), .B(n19703), .ZN(
        P2_U3144) );
  INV_X1 U21843 ( .A(n19780), .ZN(n19768) );
  AOI22_X1 U21844 ( .A1(n19706), .A2(n19782), .B1(n19777), .B2(n19705), .ZN(
        n19709) );
  AOI22_X1 U21845 ( .A1(P2_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19707), .B1(
        n19712), .B2(n19783), .ZN(n19708) );
  OAI211_X1 U21846 ( .C1(n19768), .C2(n19710), .A(n19709), .B(n19708), .ZN(
        P2_U3136) );
  AOI22_X1 U21847 ( .A1(n19783), .A2(n19718), .B1(n19711), .B2(n19777), .ZN(
        n19715) );
  AOI22_X1 U21848 ( .A1(P2_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19713), .B1(
        n19712), .B2(n19780), .ZN(n19714) );
  OAI211_X1 U21849 ( .C1(n19716), .C2(n19747), .A(n19715), .B(n19714), .ZN(
        P2_U3128) );
  AOI22_X1 U21850 ( .A1(n19783), .A2(n19724), .B1(n19717), .B2(n19777), .ZN(
        n19721) );
  AOI22_X1 U21851 ( .A1(P2_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n11085), .B1(
        n19718), .B2(n19780), .ZN(n19720) );
  OAI211_X1 U21852 ( .C1(n19722), .C2(n19747), .A(n19721), .B(n19720), .ZN(
        P2_U3120) );
  AOI22_X1 U21853 ( .A1(n19780), .A2(n19724), .B1(n19723), .B2(n19777), .ZN(
        n19728) );
  AOI22_X1 U21854 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19726), .B1(
        n19782), .B2(n19725), .ZN(n19727) );
  OAI211_X1 U21855 ( .C1(n19776), .C2(n19735), .A(n19728), .B(n19727), .ZN(
        P2_U3112) );
  AOI22_X1 U21856 ( .A1(n19730), .A2(n19782), .B1(n19729), .B2(n19777), .ZN(
        n19734) );
  AOI22_X1 U21857 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n19732), .B1(
        n19731), .B2(n19783), .ZN(n19733) );
  OAI211_X1 U21858 ( .C1(n19768), .C2(n19735), .A(n19734), .B(n19733), .ZN(
        P2_U3104) );
  AOI22_X1 U21859 ( .A1(n19737), .A2(n19782), .B1(n19777), .B2(n19736), .ZN(
        n19740) );
  AOI22_X1 U21860 ( .A1(P2_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n19738), .B1(
        n19743), .B2(n19783), .ZN(n19739) );
  OAI211_X1 U21861 ( .C1(n19768), .C2(n19741), .A(n19740), .B(n19739), .ZN(
        P2_U3096) );
  AOI22_X1 U21862 ( .A1(n19783), .A2(n19750), .B1(n19742), .B2(n19777), .ZN(
        n19746) );
  AOI22_X1 U21863 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n19744), .B1(
        n19743), .B2(n19780), .ZN(n19745) );
  OAI211_X1 U21864 ( .C1(n19748), .C2(n19747), .A(n19746), .B(n19745), .ZN(
        P2_U3088) );
  AOI22_X1 U21865 ( .A1(n19780), .A2(n19750), .B1(n19777), .B2(n19749), .ZN(
        n19754) );
  AOI22_X1 U21866 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n19752), .B1(
        n19782), .B2(n19751), .ZN(n19753) );
  OAI211_X1 U21867 ( .C1(n19776), .C2(n19755), .A(n19754), .B(n19753), .ZN(
        P2_U3080) );
  AOI22_X1 U21868 ( .A1(n19780), .A2(n19757), .B1(n19756), .B2(n19777), .ZN(
        n19761) );
  AOI22_X1 U21869 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19759), .B1(
        n19782), .B2(n19758), .ZN(n19760) );
  OAI211_X1 U21870 ( .C1(n19776), .C2(n19767), .A(n19761), .B(n19760), .ZN(
        P2_U3072) );
  AOI22_X1 U21871 ( .A1(n19763), .A2(n19782), .B1(n19777), .B2(n19762), .ZN(
        n19766) );
  AOI22_X1 U21872 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19764), .B1(
        n19771), .B2(n19783), .ZN(n19765) );
  OAI211_X1 U21873 ( .C1(n19768), .C2(n19767), .A(n19766), .B(n19765), .ZN(
        P2_U3064) );
  AOI22_X1 U21874 ( .A1(n19770), .A2(n19782), .B1(n19777), .B2(n19769), .ZN(
        n19774) );
  AOI22_X1 U21875 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19772), .B1(
        n19771), .B2(n19780), .ZN(n19773) );
  OAI211_X1 U21876 ( .C1(n19776), .C2(n19775), .A(n19774), .B(n19773), .ZN(
        P2_U3056) );
  AOI22_X1 U21877 ( .A1(n19780), .A2(n19779), .B1(n19778), .B2(n19777), .ZN(
        n19786) );
  AOI22_X1 U21878 ( .A1(n19784), .A2(n19783), .B1(n19782), .B2(n19781), .ZN(
        n19785) );
  OAI211_X1 U21879 ( .C1(n19788), .C2(n19787), .A(n19786), .B(n19785), .ZN(
        P2_U3048) );
  INV_X1 U21880 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n20098) );
  INV_X1 U21881 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n19789) );
  AOI222_X1 U21882 ( .A1(n20098), .A2(P1_DATAO_REG_30__SCAN_IN), .B1(n20101), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .C1(n19789), .C2(
        P3_DATAO_REG_30__SCAN_IN), .ZN(n19790) );
  INV_X2 U21883 ( .A(n19790), .ZN(n19850) );
  INV_X1 U21884 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n19792) );
  AOI22_X1 U21885 ( .A1(n19839), .A2(n19792), .B1(n19791), .B2(n19850), .ZN(
        U376) );
  INV_X1 U21886 ( .A(n19850), .ZN(n19853) );
  INV_X1 U21887 ( .A(P3_ADDRESS_REG_1__SCAN_IN), .ZN(n19794) );
  AOI22_X1 U21888 ( .A1(n19853), .A2(n19794), .B1(n19793), .B2(n19850), .ZN(
        U365) );
  INV_X1 U21889 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n19796) );
  AOI22_X1 U21890 ( .A1(n19839), .A2(n19796), .B1(n19795), .B2(n19850), .ZN(
        U354) );
  INV_X1 U21891 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n19798) );
  AOI22_X1 U21892 ( .A1(n19839), .A2(n19798), .B1(n19797), .B2(n19850), .ZN(
        U353) );
  INV_X1 U21893 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n19800) );
  AOI22_X1 U21894 ( .A1(n19839), .A2(n19800), .B1(n19799), .B2(n19850), .ZN(
        U352) );
  INV_X1 U21895 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n19802) );
  AOI22_X1 U21896 ( .A1(n19839), .A2(n19802), .B1(n19801), .B2(n19850), .ZN(
        U351) );
  INV_X1 U21897 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n19804) );
  AOI22_X1 U21898 ( .A1(n19853), .A2(n19804), .B1(n19803), .B2(n19850), .ZN(
        U350) );
  INV_X1 U21899 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n19806) );
  AOI22_X1 U21900 ( .A1(n19839), .A2(n19806), .B1(n19805), .B2(n19850), .ZN(
        U349) );
  INV_X1 U21901 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n19808) );
  AOI22_X1 U21902 ( .A1(n19839), .A2(n19808), .B1(n19807), .B2(n19850), .ZN(
        U348) );
  INV_X1 U21903 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n19810) );
  AOI22_X1 U21904 ( .A1(n19839), .A2(n19810), .B1(n19809), .B2(n19850), .ZN(
        U347) );
  INV_X1 U21905 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n19812) );
  AOI22_X1 U21906 ( .A1(n19839), .A2(n19812), .B1(n19811), .B2(n19850), .ZN(
        U375) );
  INV_X1 U21907 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n19814) );
  AOI22_X1 U21908 ( .A1(n19839), .A2(n19814), .B1(n19813), .B2(n19850), .ZN(
        U374) );
  INV_X1 U21909 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n19816) );
  AOI22_X1 U21910 ( .A1(n19839), .A2(n19816), .B1(n19815), .B2(n19850), .ZN(
        U373) );
  INV_X1 U21911 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n19818) );
  AOI22_X1 U21912 ( .A1(n19839), .A2(n19818), .B1(n19817), .B2(n19850), .ZN(
        U372) );
  INV_X1 U21913 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n19820) );
  AOI22_X1 U21914 ( .A1(n19839), .A2(n19820), .B1(n19819), .B2(n19850), .ZN(
        U371) );
  INV_X1 U21915 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n19822) );
  AOI22_X1 U21916 ( .A1(n19839), .A2(n19822), .B1(n19821), .B2(n19850), .ZN(
        U370) );
  INV_X1 U21917 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n19824) );
  AOI22_X1 U21918 ( .A1(n19839), .A2(n19824), .B1(n19823), .B2(n19850), .ZN(
        U369) );
  INV_X1 U21919 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n19826) );
  AOI22_X1 U21920 ( .A1(n19839), .A2(n19826), .B1(n19825), .B2(n19850), .ZN(
        U368) );
  INV_X1 U21921 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n19828) );
  AOI22_X1 U21922 ( .A1(n19839), .A2(n19828), .B1(n19827), .B2(n19850), .ZN(
        U367) );
  INV_X1 U21923 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n19830) );
  AOI22_X1 U21924 ( .A1(n19839), .A2(n19830), .B1(n19829), .B2(n19850), .ZN(
        U366) );
  INV_X1 U21925 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n19832) );
  AOI22_X1 U21926 ( .A1(n19839), .A2(n19832), .B1(n19831), .B2(n19850), .ZN(
        U364) );
  INV_X1 U21927 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n19834) );
  AOI22_X1 U21928 ( .A1(n19839), .A2(n19834), .B1(n19833), .B2(n19850), .ZN(
        U363) );
  INV_X1 U21929 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n19836) );
  AOI22_X1 U21930 ( .A1(n19839), .A2(n19836), .B1(n19835), .B2(n19850), .ZN(
        U362) );
  INV_X1 U21931 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n19838) );
  AOI22_X1 U21932 ( .A1(n19839), .A2(n19838), .B1(n19837), .B2(n19850), .ZN(
        U361) );
  INV_X1 U21933 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n19841) );
  AOI22_X1 U21934 ( .A1(n19853), .A2(n19841), .B1(n19840), .B2(n19850), .ZN(
        U360) );
  INV_X1 U21935 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n19843) );
  AOI22_X1 U21936 ( .A1(n19853), .A2(n19843), .B1(n19842), .B2(n19850), .ZN(
        U359) );
  INV_X1 U21937 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n19845) );
  AOI22_X1 U21938 ( .A1(n19853), .A2(n19845), .B1(n19844), .B2(n19850), .ZN(
        U358) );
  INV_X1 U21939 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n19847) );
  AOI22_X1 U21940 ( .A1(n19853), .A2(n19847), .B1(n19846), .B2(n19850), .ZN(
        U357) );
  INV_X1 U21941 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n19849) );
  AOI22_X1 U21942 ( .A1(n19853), .A2(n19849), .B1(n19848), .B2(n19850), .ZN(
        U356) );
  INV_X1 U21943 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n19852) );
  AOI22_X1 U21944 ( .A1(n19853), .A2(n19852), .B1(n19851), .B2(n19850), .ZN(
        U355) );
  AOI22_X1 U21945 ( .A1(n21325), .A2(P1_LWORD_REG_0__SCAN_IN), .B1(n19866), 
        .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n19855) );
  OAI21_X1 U21946 ( .B1(n19856), .B2(n19885), .A(n19855), .ZN(P1_U2936) );
  AOI22_X1 U21947 ( .A1(n19869), .A2(P1_LWORD_REG_1__SCAN_IN), .B1(n19866), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n19857) );
  OAI21_X1 U21948 ( .B1(n19858), .B2(n19885), .A(n19857), .ZN(P1_U2935) );
  AOI22_X1 U21949 ( .A1(n19869), .A2(P1_LWORD_REG_2__SCAN_IN), .B1(n19866), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n19859) );
  OAI21_X1 U21950 ( .B1(n19860), .B2(n19885), .A(n19859), .ZN(P1_U2934) );
  AOI22_X1 U21951 ( .A1(n19869), .A2(P1_LWORD_REG_3__SCAN_IN), .B1(n19866), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n19861) );
  OAI21_X1 U21952 ( .B1(n19862), .B2(n19885), .A(n19861), .ZN(P1_U2933) );
  AOI22_X1 U21953 ( .A1(n19869), .A2(P1_LWORD_REG_4__SCAN_IN), .B1(n19866), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .ZN(n19863) );
  OAI21_X1 U21954 ( .B1(n19864), .B2(n19885), .A(n19863), .ZN(P1_U2932) );
  AOI22_X1 U21955 ( .A1(n19869), .A2(P1_LWORD_REG_5__SCAN_IN), .B1(n19866), 
        .B2(P1_DATAO_REG_5__SCAN_IN), .ZN(n19865) );
  OAI21_X1 U21956 ( .B1(n11769), .B2(n19885), .A(n19865), .ZN(P1_U2931) );
  AOI22_X1 U21957 ( .A1(n19869), .A2(P1_LWORD_REG_6__SCAN_IN), .B1(n19866), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n19867) );
  OAI21_X1 U21958 ( .B1(n11847), .B2(n19885), .A(n19867), .ZN(P1_U2930) );
  AOI22_X1 U21959 ( .A1(n21325), .A2(P1_LWORD_REG_7__SCAN_IN), .B1(n19866), 
        .B2(P1_DATAO_REG_7__SCAN_IN), .ZN(n19868) );
  OAI21_X1 U21960 ( .B1(n11859), .B2(n19885), .A(n19868), .ZN(P1_U2929) );
  AOI22_X1 U21961 ( .A1(n19869), .A2(P1_LWORD_REG_8__SCAN_IN), .B1(n19866), 
        .B2(P1_DATAO_REG_8__SCAN_IN), .ZN(n19870) );
  OAI21_X1 U21962 ( .B1(n19871), .B2(n19885), .A(n19870), .ZN(P1_U2928) );
  AOI22_X1 U21963 ( .A1(n21325), .A2(P1_LWORD_REG_9__SCAN_IN), .B1(n19866), 
        .B2(P1_DATAO_REG_9__SCAN_IN), .ZN(n19872) );
  OAI21_X1 U21964 ( .B1(n19873), .B2(n19885), .A(n19872), .ZN(P1_U2927) );
  AOI22_X1 U21965 ( .A1(n21325), .A2(P1_LWORD_REG_10__SCAN_IN), .B1(n19866), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n19874) );
  OAI21_X1 U21966 ( .B1(n19875), .B2(n19885), .A(n19874), .ZN(P1_U2926) );
  AOI22_X1 U21967 ( .A1(n21325), .A2(P1_LWORD_REG_11__SCAN_IN), .B1(n19866), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n19876) );
  OAI21_X1 U21968 ( .B1(n19877), .B2(n19885), .A(n19876), .ZN(P1_U2925) );
  AOI22_X1 U21969 ( .A1(n21325), .A2(P1_LWORD_REG_12__SCAN_IN), .B1(n19866), 
        .B2(P1_DATAO_REG_12__SCAN_IN), .ZN(n19878) );
  OAI21_X1 U21970 ( .B1(n19879), .B2(n19885), .A(n19878), .ZN(P1_U2924) );
  AOI22_X1 U21971 ( .A1(n21325), .A2(P1_LWORD_REG_13__SCAN_IN), .B1(n19866), 
        .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n19880) );
  OAI21_X1 U21972 ( .B1(n19881), .B2(n19885), .A(n19880), .ZN(P1_U2923) );
  AOI22_X1 U21973 ( .A1(n21325), .A2(P1_LWORD_REG_14__SCAN_IN), .B1(n19866), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n19882) );
  OAI21_X1 U21974 ( .B1(n19883), .B2(n19885), .A(n19882), .ZN(P1_U2922) );
  AOI22_X1 U21975 ( .A1(n21325), .A2(P1_LWORD_REG_15__SCAN_IN), .B1(n19866), 
        .B2(P1_DATAO_REG_15__SCAN_IN), .ZN(n19884) );
  OAI21_X1 U21976 ( .B1(n15702), .B2(n19885), .A(n19884), .ZN(P1_U2921) );
  INV_X2 U21977 ( .A(n22219), .ZN(n22221) );
  INV_X1 U21978 ( .A(n19920), .ZN(n19932) );
  INV_X1 U21979 ( .A(P1_REIP_REG_2__SCAN_IN), .ZN(n19888) );
  NAND2_X1 U21980 ( .A1(n22221), .A2(n21725), .ZN(n19927) );
  INV_X1 U21981 ( .A(n19927), .ZN(n19917) );
  OAI222_X1 U21982 ( .A1(n19932), .A2(n19947), .B1(n19886), .B2(n22221), .C1(
        n19888), .C2(n19928), .ZN(P1_U3197) );
  AOI22_X1 U21983 ( .A1(P1_REIP_REG_3__SCAN_IN), .A2(n19917), .B1(
        P1_ADDRESS_REG_1__SCAN_IN), .B2(n22219), .ZN(n19887) );
  OAI21_X1 U21984 ( .B1(n19888), .B2(n19932), .A(n19887), .ZN(P1_U3198) );
  AOI22_X1 U21985 ( .A1(P1_REIP_REG_3__SCAN_IN), .A2(n19920), .B1(
        P1_ADDRESS_REG_2__SCAN_IN), .B2(n22219), .ZN(n19889) );
  OAI21_X1 U21986 ( .B1(n21437), .B2(n19928), .A(n19889), .ZN(P1_U3199) );
  INV_X1 U21987 ( .A(P1_ADDRESS_REG_3__SCAN_IN), .ZN(n19890) );
  OAI222_X1 U21988 ( .A1(n19928), .A2(n11382), .B1(n19890), .B2(n22221), .C1(
        n21437), .C2(n19932), .ZN(P1_U3200) );
  INV_X1 U21989 ( .A(P1_ADDRESS_REG_4__SCAN_IN), .ZN(n19891) );
  OAI222_X1 U21990 ( .A1(n19927), .A2(n21463), .B1(n19891), .B2(n22221), .C1(
        n11382), .C2(n19932), .ZN(P1_U3201) );
  INV_X1 U21991 ( .A(P1_ADDRESS_REG_5__SCAN_IN), .ZN(n19892) );
  INV_X1 U21992 ( .A(P1_REIP_REG_7__SCAN_IN), .ZN(n21473) );
  OAI222_X1 U21993 ( .A1(n19932), .A2(n21463), .B1(n19892), .B2(n22221), .C1(
        n21473), .C2(n19928), .ZN(P1_U3202) );
  INV_X1 U21994 ( .A(P1_ADDRESS_REG_6__SCAN_IN), .ZN(n19893) );
  OAI222_X1 U21995 ( .A1(n19932), .A2(n21473), .B1(n19893), .B2(n22221), .C1(
        n19895), .C2(n19928), .ZN(P1_U3203) );
  AOI22_X1 U21996 ( .A1(P1_REIP_REG_9__SCAN_IN), .A2(n19917), .B1(
        P1_ADDRESS_REG_7__SCAN_IN), .B2(n22219), .ZN(n19894) );
  OAI21_X1 U21997 ( .B1(n19895), .B2(n19932), .A(n19894), .ZN(P1_U3204) );
  AOI22_X1 U21998 ( .A1(P1_REIP_REG_9__SCAN_IN), .A2(n19920), .B1(
        P1_ADDRESS_REG_8__SCAN_IN), .B2(n22219), .ZN(n19896) );
  OAI21_X1 U21999 ( .B1(n19897), .B2(n19928), .A(n19896), .ZN(P1_U3205) );
  INV_X1 U22000 ( .A(P1_ADDRESS_REG_9__SCAN_IN), .ZN(n19898) );
  OAI222_X1 U22001 ( .A1(n19928), .A2(n21509), .B1(n19898), .B2(n22221), .C1(
        n19897), .C2(n19932), .ZN(P1_U3206) );
  INV_X1 U22002 ( .A(P1_REIP_REG_12__SCAN_IN), .ZN(n21514) );
  INV_X1 U22003 ( .A(P1_ADDRESS_REG_10__SCAN_IN), .ZN(n19899) );
  OAI222_X1 U22004 ( .A1(n19928), .A2(n21514), .B1(n19899), .B2(n22221), .C1(
        n21509), .C2(n19932), .ZN(P1_U3207) );
  INV_X1 U22005 ( .A(P1_ADDRESS_REG_11__SCAN_IN), .ZN(n19900) );
  OAI222_X1 U22006 ( .A1(n19927), .A2(n21522), .B1(n19900), .B2(n22221), .C1(
        n21514), .C2(n19932), .ZN(P1_U3208) );
  AOI22_X1 U22007 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(n19917), .B1(
        P1_ADDRESS_REG_12__SCAN_IN), .B2(n22219), .ZN(n19901) );
  OAI21_X1 U22008 ( .B1(n21522), .B2(n19932), .A(n19901), .ZN(P1_U3209) );
  AOI22_X1 U22009 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(n19920), .B1(
        P1_ADDRESS_REG_13__SCAN_IN), .B2(n22219), .ZN(n19902) );
  OAI21_X1 U22010 ( .B1(n19904), .B2(n19928), .A(n19902), .ZN(P1_U3210) );
  AOI22_X1 U22011 ( .A1(P1_REIP_REG_16__SCAN_IN), .A2(n19917), .B1(
        P1_ADDRESS_REG_14__SCAN_IN), .B2(n22219), .ZN(n19903) );
  OAI21_X1 U22012 ( .B1(n19904), .B2(n19932), .A(n19903), .ZN(P1_U3211) );
  AOI22_X1 U22013 ( .A1(P1_REIP_REG_16__SCAN_IN), .A2(n19920), .B1(
        P1_ADDRESS_REG_15__SCAN_IN), .B2(n22219), .ZN(n19905) );
  OAI21_X1 U22014 ( .B1(n21366), .B2(n19928), .A(n19905), .ZN(P1_U3212) );
  INV_X1 U22015 ( .A(P1_REIP_REG_18__SCAN_IN), .ZN(n21569) );
  INV_X1 U22016 ( .A(P1_ADDRESS_REG_16__SCAN_IN), .ZN(n19906) );
  OAI222_X1 U22017 ( .A1(n19927), .A2(n21569), .B1(n19906), .B2(n22221), .C1(
        n21366), .C2(n19932), .ZN(P1_U3213) );
  INV_X1 U22018 ( .A(P1_ADDRESS_REG_17__SCAN_IN), .ZN(n19907) );
  OAI222_X1 U22019 ( .A1(n19927), .A2(n21582), .B1(n19907), .B2(n22221), .C1(
        n21569), .C2(n19932), .ZN(P1_U3214) );
  INV_X1 U22020 ( .A(P1_ADDRESS_REG_18__SCAN_IN), .ZN(n19908) );
  OAI222_X1 U22021 ( .A1(n19927), .A2(n19909), .B1(n19908), .B2(n22221), .C1(
        n21582), .C2(n19932), .ZN(P1_U3215) );
  INV_X1 U22022 ( .A(P1_ADDRESS_REG_19__SCAN_IN), .ZN(n19910) );
  OAI222_X1 U22023 ( .A1(n19927), .A2(n21601), .B1(n19910), .B2(n22221), .C1(
        n19909), .C2(n19932), .ZN(P1_U3216) );
  INV_X1 U22024 ( .A(P1_ADDRESS_REG_20__SCAN_IN), .ZN(n19911) );
  OAI222_X1 U22025 ( .A1(n19927), .A2(n21615), .B1(n19911), .B2(n22221), .C1(
        n21601), .C2(n19932), .ZN(P1_U3217) );
  INV_X1 U22026 ( .A(P1_ADDRESS_REG_21__SCAN_IN), .ZN(n19912) );
  OAI222_X1 U22027 ( .A1(n19927), .A2(n19913), .B1(n19912), .B2(n22221), .C1(
        n21615), .C2(n19932), .ZN(P1_U3218) );
  INV_X1 U22028 ( .A(P1_ADDRESS_REG_22__SCAN_IN), .ZN(n19914) );
  OAI222_X1 U22029 ( .A1(n19927), .A2(n19915), .B1(n19914), .B2(n22221), .C1(
        n19913), .C2(n19932), .ZN(P1_U3219) );
  INV_X1 U22030 ( .A(P1_ADDRESS_REG_23__SCAN_IN), .ZN(n19916) );
  OAI222_X1 U22031 ( .A1(n19927), .A2(n19919), .B1(n19916), .B2(n22221), .C1(
        n19915), .C2(n19932), .ZN(P1_U3220) );
  AOI22_X1 U22032 ( .A1(P1_REIP_REG_26__SCAN_IN), .A2(n19917), .B1(
        P1_ADDRESS_REG_24__SCAN_IN), .B2(n22219), .ZN(n19918) );
  OAI21_X1 U22033 ( .B1(n19919), .B2(n19932), .A(n19918), .ZN(P1_U3221) );
  AOI22_X1 U22034 ( .A1(P1_REIP_REG_26__SCAN_IN), .A2(n19920), .B1(
        P1_ADDRESS_REG_25__SCAN_IN), .B2(n22219), .ZN(n19921) );
  OAI21_X1 U22035 ( .B1(n21385), .B2(n19928), .A(n19921), .ZN(P1_U3222) );
  INV_X1 U22036 ( .A(P1_ADDRESS_REG_26__SCAN_IN), .ZN(n19922) );
  OAI222_X1 U22037 ( .A1(n19928), .A2(n19924), .B1(n19922), .B2(n22221), .C1(
        n21385), .C2(n19932), .ZN(P1_U3223) );
  INV_X1 U22038 ( .A(P1_ADDRESS_REG_27__SCAN_IN), .ZN(n19923) );
  OAI222_X1 U22039 ( .A1(n19932), .A2(n19924), .B1(n19923), .B2(n22221), .C1(
        n19925), .C2(n19928), .ZN(P1_U3224) );
  INV_X1 U22040 ( .A(P1_ADDRESS_REG_28__SCAN_IN), .ZN(n19926) );
  OAI222_X1 U22041 ( .A1(n19927), .A2(n19931), .B1(n19926), .B2(n22221), .C1(
        n19925), .C2(n19932), .ZN(P1_U3225) );
  INV_X1 U22042 ( .A(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n19930) );
  OAI222_X1 U22043 ( .A1(n19932), .A2(n19931), .B1(n19930), .B2(n22221), .C1(
        n19929), .C2(n19928), .ZN(P1_U3226) );
  INV_X1 U22044 ( .A(P1_BE_N_REG_3__SCAN_IN), .ZN(n19933) );
  AOI22_X1 U22045 ( .A1(n22221), .A2(n19934), .B1(n19933), .B2(n22219), .ZN(
        P1_U3458) );
  AOI221_X1 U22046 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(P1_REIP_REG_1__SCAN_IN), 
        .C1(P1_DATAWIDTH_REG_0__SCAN_IN), .C2(P1_REIP_REG_1__SCAN_IN), .A(
        P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n19945) );
  NOR4_X1 U22047 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_12__SCAN_IN), .A3(P1_DATAWIDTH_REG_11__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_10__SCAN_IN), .ZN(n19938) );
  NOR4_X1 U22048 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_17__SCAN_IN), .A3(P1_DATAWIDTH_REG_16__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_14__SCAN_IN), .ZN(n19937) );
  NOR4_X1 U22049 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_4__SCAN_IN), .A3(P1_DATAWIDTH_REG_3__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_2__SCAN_IN), .ZN(n19936) );
  NOR4_X1 U22050 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_8__SCAN_IN), .A3(P1_DATAWIDTH_REG_7__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_6__SCAN_IN), .ZN(n19935) );
  NAND4_X1 U22051 ( .A1(n19938), .A2(n19937), .A3(n19936), .A4(n19935), .ZN(
        n19944) );
  NOR4_X1 U22052 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_29__SCAN_IN), .A3(P1_DATAWIDTH_REG_28__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_27__SCAN_IN), .ZN(n19942) );
  AOI211_X1 U22053 ( .C1(P1_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_15__SCAN_IN), .B(
        P1_DATAWIDTH_REG_31__SCAN_IN), .ZN(n19941) );
  NOR4_X1 U22054 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_21__SCAN_IN), .A3(P1_DATAWIDTH_REG_20__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_19__SCAN_IN), .ZN(n19940) );
  NOR4_X1 U22055 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_25__SCAN_IN), .A3(P1_DATAWIDTH_REG_24__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_23__SCAN_IN), .ZN(n19939) );
  NAND4_X1 U22056 ( .A1(n19942), .A2(n19941), .A3(n19940), .A4(n19939), .ZN(
        n19943) );
  NOR2_X1 U22057 ( .A1(n19944), .A2(n19943), .ZN(n19958) );
  MUX2_X1 U22058 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .B(n19945), .S(n19958), 
        .Z(P1_U2808) );
  INV_X1 U22059 ( .A(P1_BE_N_REG_2__SCAN_IN), .ZN(n19946) );
  AOI22_X1 U22060 ( .A1(n22221), .A2(n19950), .B1(n19946), .B2(n22219), .ZN(
        P1_U3459) );
  AOI21_X1 U22061 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n19948) );
  OAI221_X1 U22062 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n19948), .C1(n19947), 
        .C2(P1_REIP_REG_0__SCAN_IN), .A(n19958), .ZN(n19949) );
  OAI21_X1 U22063 ( .B1(n19958), .B2(n19950), .A(n19949), .ZN(P1_U3481) );
  INV_X1 U22064 ( .A(P1_BE_N_REG_1__SCAN_IN), .ZN(n19951) );
  AOI22_X1 U22065 ( .A1(n22221), .A2(n19954), .B1(n19951), .B2(n22219), .ZN(
        P1_U3460) );
  NOR3_X1 U22066 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A3(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n19952) );
  OAI21_X1 U22067 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n19952), .A(n19958), .ZN(
        n19953) );
  OAI21_X1 U22068 ( .B1(n19958), .B2(n19954), .A(n19953), .ZN(P1_U2807) );
  INV_X1 U22069 ( .A(P1_BE_N_REG_0__SCAN_IN), .ZN(n19955) );
  AOI22_X1 U22070 ( .A1(n22221), .A2(n19957), .B1(n19955), .B2(n22219), .ZN(
        P1_U3461) );
  OAI21_X1 U22071 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(P1_REIP_REG_0__SCAN_IN), 
        .A(n19958), .ZN(n19956) );
  OAI21_X1 U22072 ( .B1(n19958), .B2(n19957), .A(n19956), .ZN(P1_U3482) );
  INV_X1 U22073 ( .A(n19959), .ZN(n21546) );
  AOI22_X1 U22074 ( .A1(n21547), .A2(n19962), .B1(n19961), .B2(n21546), .ZN(
        n19960) );
  OAI21_X1 U22075 ( .B1(n19969), .B2(n21542), .A(n19960), .ZN(P1_U2857) );
  AOI22_X1 U22076 ( .A1(n21535), .A2(n19962), .B1(n19961), .B2(n21533), .ZN(
        n19963) );
  OAI21_X1 U22077 ( .B1(n19969), .B2(n19964), .A(n19963), .ZN(P1_U2858) );
  OAI22_X1 U22078 ( .A1(n21649), .A2(n19966), .B1(n21647), .B2(n19965), .ZN(
        n19967) );
  INV_X1 U22079 ( .A(n19967), .ZN(n19968) );
  OAI21_X1 U22080 ( .B1(n19969), .B2(n21641), .A(n19968), .ZN(P1_U2846) );
  INV_X1 U22081 ( .A(n19970), .ZN(n19973) );
  INV_X1 U22082 ( .A(n19971), .ZN(n19972) );
  AOI21_X1 U22083 ( .B1(n19973), .B2(n21658), .A(n19972), .ZN(n21411) );
  INV_X1 U22084 ( .A(n21655), .ZN(n20024) );
  OR2_X1 U22085 ( .A1(n20022), .A2(n19974), .ZN(n19975) );
  AOI22_X1 U22086 ( .A1(n21411), .A2(n20024), .B1(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n19975), .ZN(n19976) );
  NAND2_X1 U22087 ( .A1(n10970), .A2(P1_REIP_REG_0__SCAN_IN), .ZN(n21418) );
  OAI211_X1 U22088 ( .C1(n19977), .C2(n20018), .A(n19976), .B(n21418), .ZN(
        P1_U2999) );
  OAI22_X1 U22089 ( .A1(n21445), .A2(n20018), .B1(n21447), .B2(n20028), .ZN(
        n19978) );
  AOI21_X1 U22090 ( .B1(n20024), .B2(n19979), .A(n19978), .ZN(n19981) );
  OAI211_X1 U22091 ( .C1(n19987), .C2(n19982), .A(n19981), .B(n19980), .ZN(
        P1_U2994) );
  INV_X1 U22092 ( .A(n21477), .ZN(n19983) );
  AOI222_X1 U22093 ( .A1(n19984), .A2(n20024), .B1(n20009), .B2(n21474), .C1(
        n19983), .C2(n20005), .ZN(n19986) );
  OAI211_X1 U22094 ( .C1(n19987), .C2(n21467), .A(n19986), .B(n19985), .ZN(
        P1_U2992) );
  AOI22_X1 U22095 ( .A1(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n20022), .B1(
        n10970), .B2(P1_REIP_REG_10__SCAN_IN), .ZN(n19990) );
  INV_X1 U22096 ( .A(n19988), .ZN(n21494) );
  AOI22_X1 U22097 ( .A1(n21495), .A2(n20009), .B1(n21494), .B2(n20005), .ZN(
        n19989) );
  OAI211_X1 U22098 ( .C1(n21655), .C2(n19991), .A(n19990), .B(n19989), .ZN(
        P1_U2989) );
  NOR2_X1 U22099 ( .A1(n21386), .A2(n21509), .ZN(n21341) );
  NAND2_X1 U22100 ( .A1(n19994), .A2(n19992), .ZN(n19993) );
  MUX2_X1 U22101 ( .A(n19994), .B(n19993), .S(n15994), .Z(n19995) );
  OAI22_X1 U22102 ( .A1(n21339), .A2(n21655), .B1(n20028), .B2(n21503), .ZN(
        n19996) );
  OAI21_X1 U22103 ( .B1(n20018), .B2(n21502), .A(n19997), .ZN(P1_U2988) );
  AOI22_X1 U22104 ( .A1(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n20022), .B1(
        n10970), .B2(P1_REIP_REG_12__SCAN_IN), .ZN(n20000) );
  AOI22_X1 U22105 ( .A1(n20005), .A2(n21516), .B1(n20009), .B2(n19998), .ZN(
        n19999) );
  OAI211_X1 U22106 ( .C1(n20001), .C2(n21655), .A(n20000), .B(n19999), .ZN(
        P1_U2987) );
  AOI22_X1 U22107 ( .A1(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n20022), .B1(
        n10970), .B2(P1_REIP_REG_14__SCAN_IN), .ZN(n20003) );
  AOI22_X1 U22108 ( .A1(n21535), .A2(n20009), .B1(n20005), .B2(n21534), .ZN(
        n20002) );
  OAI211_X1 U22109 ( .C1(n20004), .C2(n21655), .A(n20003), .B(n20002), .ZN(
        P1_U2985) );
  AOI22_X1 U22110 ( .A1(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n20022), .B1(
        n10970), .B2(P1_REIP_REG_15__SCAN_IN), .ZN(n20007) );
  AOI22_X1 U22111 ( .A1(n21547), .A2(n20009), .B1(n20005), .B2(n21545), .ZN(
        n20006) );
  OAI211_X1 U22112 ( .C1(n20008), .C2(n21655), .A(n20007), .B(n20006), .ZN(
        P1_U2984) );
  AOI22_X1 U22113 ( .A1(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n20022), .B1(
        n10970), .B2(P1_REIP_REG_16__SCAN_IN), .ZN(n20012) );
  AOI22_X1 U22114 ( .A1(n20010), .A2(n20024), .B1(n20009), .B2(n21554), .ZN(
        n20011) );
  OAI211_X1 U22115 ( .C1(n20028), .C2(n21552), .A(n20012), .B(n20011), .ZN(
        P1_U2983) );
  AOI22_X1 U22116 ( .A1(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n20022), .B1(
        n10970), .B2(P1_REIP_REG_20__SCAN_IN), .ZN(n20016) );
  AOI22_X1 U22117 ( .A1(n20014), .A2(n20009), .B1(n20024), .B2(n20013), .ZN(
        n20015) );
  OAI211_X1 U22118 ( .C1(n20028), .C2(n21590), .A(n20016), .B(n20015), .ZN(
        P1_U2979) );
  AOI22_X1 U22119 ( .A1(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n20022), .B1(
        n10970), .B2(P1_REIP_REG_22__SCAN_IN), .ZN(n20021) );
  OAI22_X1 U22120 ( .A1(n21603), .A2(n20018), .B1(n21655), .B2(n20017), .ZN(
        n20019) );
  INV_X1 U22121 ( .A(n20019), .ZN(n20020) );
  OAI211_X1 U22122 ( .C1(n20028), .C2(n21605), .A(n20021), .B(n20020), .ZN(
        P1_U2977) );
  AOI22_X1 U22123 ( .A1(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n20022), .B1(
        n10970), .B2(P1_REIP_REG_24__SCAN_IN), .ZN(n20027) );
  AOI22_X1 U22124 ( .A1(n20025), .A2(n20009), .B1(n20024), .B2(n20023), .ZN(
        n20026) );
  OAI211_X1 U22125 ( .C1(n20028), .C2(n21619), .A(n20027), .B(n20026), .ZN(
        P1_U2975) );
  AND2_X1 U22126 ( .A1(n20030), .A2(n20029), .ZN(n20032) );
  OAI22_X1 U22127 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20033), .B1(n20032), 
        .B2(n20031), .ZN(P1_U2803) );
  INV_X1 U22128 ( .A(P1_D_C_N_REG_SCAN_IN), .ZN(n20036) );
  OAI21_X1 U22129 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n21725), .A(n20034), 
        .ZN(n20035) );
  AOI22_X1 U22130 ( .A1(n22221), .A2(P1_CODEFETCH_REG_SCAN_IN), .B1(n20036), 
        .B2(n20035), .ZN(P1_U2804) );
  INV_X2 U22131 ( .A(U212), .ZN(n20080) );
  AOI22_X1 U22132 ( .A1(P1_DATAO_REG_0__SCAN_IN), .A2(n20089), .B1(
        P2_DATAO_REG_0__SCAN_IN), .B2(n20080), .ZN(n20038) );
  OAI21_X1 U22133 ( .B1(n20039), .B2(n20100), .A(n20038), .ZN(U247) );
  INV_X1 U22134 ( .A(BUF1_REG_1__SCAN_IN), .ZN(n20041) );
  AOI22_X1 U22135 ( .A1(P1_DATAO_REG_1__SCAN_IN), .A2(n20089), .B1(
        P2_DATAO_REG_1__SCAN_IN), .B2(n20080), .ZN(n20040) );
  OAI21_X1 U22136 ( .B1(n20041), .B2(n20100), .A(n20040), .ZN(U246) );
  AOI22_X1 U22137 ( .A1(P1_DATAO_REG_2__SCAN_IN), .A2(n20089), .B1(
        P2_DATAO_REG_2__SCAN_IN), .B2(n20080), .ZN(n20042) );
  OAI21_X1 U22138 ( .B1(n13789), .B2(n20100), .A(n20042), .ZN(U245) );
  AOI22_X1 U22139 ( .A1(P1_DATAO_REG_3__SCAN_IN), .A2(n20089), .B1(
        P2_DATAO_REG_3__SCAN_IN), .B2(n20080), .ZN(n20043) );
  OAI21_X1 U22140 ( .B1(n13915), .B2(n20100), .A(n20043), .ZN(U244) );
  AOI22_X1 U22141 ( .A1(P1_DATAO_REG_4__SCAN_IN), .A2(n20089), .B1(
        P2_DATAO_REG_4__SCAN_IN), .B2(n20080), .ZN(n20044) );
  OAI21_X1 U22142 ( .B1(n20045), .B2(n20100), .A(n20044), .ZN(U243) );
  AOI22_X1 U22143 ( .A1(P1_DATAO_REG_5__SCAN_IN), .A2(n20089), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n20080), .ZN(n20046) );
  OAI21_X1 U22144 ( .B1(n14164), .B2(n20100), .A(n20046), .ZN(U242) );
  AOI22_X1 U22145 ( .A1(P1_DATAO_REG_6__SCAN_IN), .A2(n20089), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n20080), .ZN(n20047) );
  OAI21_X1 U22146 ( .B1(n20048), .B2(n20100), .A(n20047), .ZN(U241) );
  INV_X1 U22147 ( .A(BUF1_REG_7__SCAN_IN), .ZN(n20050) );
  AOI22_X1 U22148 ( .A1(P1_DATAO_REG_7__SCAN_IN), .A2(n20089), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n20080), .ZN(n20049) );
  OAI21_X1 U22149 ( .B1(n20050), .B2(n20100), .A(n20049), .ZN(U240) );
  INV_X1 U22150 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n20052) );
  AOI22_X1 U22151 ( .A1(P1_DATAO_REG_8__SCAN_IN), .A2(n20089), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n20080), .ZN(n20051) );
  OAI21_X1 U22152 ( .B1(n20052), .B2(n20100), .A(n20051), .ZN(U239) );
  AOI22_X1 U22153 ( .A1(P1_DATAO_REG_9__SCAN_IN), .A2(n20089), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n20080), .ZN(n20053) );
  OAI21_X1 U22154 ( .B1(n13718), .B2(n20100), .A(n20053), .ZN(U238) );
  AOI22_X1 U22155 ( .A1(P1_DATAO_REG_10__SCAN_IN), .A2(n20089), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n20080), .ZN(n20054) );
  OAI21_X1 U22156 ( .B1(n20055), .B2(n20100), .A(n20054), .ZN(U237) );
  INV_X1 U22157 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n20057) );
  AOI22_X1 U22158 ( .A1(P1_DATAO_REG_11__SCAN_IN), .A2(n20089), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n20080), .ZN(n20056) );
  OAI21_X1 U22159 ( .B1(n20057), .B2(n20100), .A(n20056), .ZN(U236) );
  INV_X1 U22160 ( .A(BUF1_REG_12__SCAN_IN), .ZN(n20059) );
  AOI22_X1 U22161 ( .A1(P1_DATAO_REG_12__SCAN_IN), .A2(n20089), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n20080), .ZN(n20058) );
  OAI21_X1 U22162 ( .B1(n20059), .B2(n20100), .A(n20058), .ZN(U235) );
  INV_X1 U22163 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n20061) );
  AOI22_X1 U22164 ( .A1(P1_DATAO_REG_13__SCAN_IN), .A2(n20089), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n20080), .ZN(n20060) );
  OAI21_X1 U22165 ( .B1(n20061), .B2(n20100), .A(n20060), .ZN(U234) );
  INV_X1 U22166 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n20063) );
  AOI22_X1 U22167 ( .A1(P1_DATAO_REG_14__SCAN_IN), .A2(n20089), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n20080), .ZN(n20062) );
  OAI21_X1 U22168 ( .B1(n20063), .B2(n20100), .A(n20062), .ZN(U233) );
  INV_X1 U22169 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n20065) );
  AOI22_X1 U22170 ( .A1(P1_DATAO_REG_15__SCAN_IN), .A2(n20089), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n20080), .ZN(n20064) );
  OAI21_X1 U22171 ( .B1(n20065), .B2(n20100), .A(n20064), .ZN(U232) );
  AOI22_X1 U22172 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n20089), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n20080), .ZN(n20066) );
  OAI21_X1 U22173 ( .B1(n20067), .B2(n20100), .A(n20066), .ZN(U231) );
  AOI22_X1 U22174 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(n20089), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n20080), .ZN(n20068) );
  OAI21_X1 U22175 ( .B1(n20069), .B2(n20100), .A(n20068), .ZN(U230) );
  AOI22_X1 U22176 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(n20089), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n20080), .ZN(n20070) );
  OAI21_X1 U22177 ( .B1(n20071), .B2(n20100), .A(n20070), .ZN(U229) );
  AOI22_X1 U22178 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(n20089), .B1(
        P2_DATAO_REG_19__SCAN_IN), .B2(n20080), .ZN(n20072) );
  OAI21_X1 U22179 ( .B1(n20073), .B2(n20100), .A(n20072), .ZN(U228) );
  AOI22_X1 U22180 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n20089), .B1(
        P2_DATAO_REG_20__SCAN_IN), .B2(n20080), .ZN(n20074) );
  OAI21_X1 U22181 ( .B1(n20075), .B2(n20100), .A(n20074), .ZN(U227) );
  AOI22_X1 U22182 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(n20089), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(n20080), .ZN(n20076) );
  OAI21_X1 U22183 ( .B1(n20077), .B2(n20100), .A(n20076), .ZN(U226) );
  AOI22_X1 U22184 ( .A1(P1_DATAO_REG_22__SCAN_IN), .A2(n20089), .B1(
        P2_DATAO_REG_22__SCAN_IN), .B2(n20080), .ZN(n20078) );
  OAI21_X1 U22185 ( .B1(n20079), .B2(n20100), .A(n20078), .ZN(U225) );
  AOI22_X1 U22186 ( .A1(P1_DATAO_REG_23__SCAN_IN), .A2(n20089), .B1(
        P2_DATAO_REG_23__SCAN_IN), .B2(n20080), .ZN(n20081) );
  OAI21_X1 U22187 ( .B1(n20082), .B2(n20100), .A(n20081), .ZN(U224) );
  AOI22_X1 U22188 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n20089), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(n20080), .ZN(n20083) );
  OAI21_X1 U22189 ( .B1(n20084), .B2(n20100), .A(n20083), .ZN(U223) );
  AOI22_X1 U22190 ( .A1(P1_DATAO_REG_25__SCAN_IN), .A2(n20089), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(n20080), .ZN(n20085) );
  OAI21_X1 U22191 ( .B1(n20086), .B2(n20100), .A(n20085), .ZN(U222) );
  AOI22_X1 U22192 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(n20089), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(n20080), .ZN(n20087) );
  OAI21_X1 U22193 ( .B1(n20088), .B2(n20100), .A(n20087), .ZN(U221) );
  AOI22_X1 U22194 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(n20089), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(n20080), .ZN(n20090) );
  OAI21_X1 U22195 ( .B1(n20091), .B2(n20100), .A(n20090), .ZN(U220) );
  AOI22_X1 U22196 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(n20089), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(n20080), .ZN(n20092) );
  OAI21_X1 U22197 ( .B1(n20093), .B2(n20100), .A(n20092), .ZN(U219) );
  AOI22_X1 U22198 ( .A1(P1_DATAO_REG_29__SCAN_IN), .A2(n20089), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n20080), .ZN(n20094) );
  OAI21_X1 U22199 ( .B1(n20095), .B2(n20100), .A(n20094), .ZN(U218) );
  AOI22_X1 U22200 ( .A1(P1_DATAO_REG_30__SCAN_IN), .A2(n20089), .B1(
        P2_DATAO_REG_30__SCAN_IN), .B2(n20080), .ZN(n20096) );
  OAI21_X1 U22201 ( .B1(n20097), .B2(n20100), .A(n20096), .ZN(U217) );
  OAI222_X1 U22202 ( .A1(U212), .A2(n20101), .B1(n20100), .B2(n20099), .C1(
        U214), .C2(n20098), .ZN(U216) );
  AOI22_X1 U22203 ( .A1(n22221), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n20102), 
        .B2(n22219), .ZN(P1_U3483) );
  OAI21_X1 U22204 ( .B1(P3_STATEBS16_REG_SCAN_IN), .B2(n20171), .A(n20164), 
        .ZN(n20103) );
  AOI211_X1 U22205 ( .C1(n20104), .C2(n20103), .A(n21707), .B(n21288), .ZN(
        n20106) );
  INV_X1 U22206 ( .A(n21301), .ZN(n20105) );
  OAI21_X1 U22207 ( .B1(n20106), .B2(n21309), .A(n20105), .ZN(n20110) );
  AOI21_X1 U22208 ( .B1(n21755), .B2(n21248), .A(n20165), .ZN(n20107) );
  OAI21_X1 U22209 ( .B1(n20108), .B2(n21305), .A(n20107), .ZN(n20109) );
  MUX2_X1 U22210 ( .A(P3_REQUESTPENDING_REG_SCAN_IN), .B(n20110), .S(n20109), 
        .Z(P3_U3296) );
  NOR2_X4 U22211 ( .A1(n20159), .A2(n20152), .ZN(n20158) );
  AOI22_X1 U22212 ( .A1(P3_EAX_REG_16__SCAN_IN), .A2(n20152), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n20158), .ZN(n20114) );
  OAI21_X1 U22213 ( .B1(n20135), .B2(n20154), .A(n20114), .ZN(P3_U2768) );
  AOI22_X1 U22214 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n20159), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n20158), .ZN(n20115) );
  OAI21_X1 U22215 ( .B1(n20672), .B2(n20161), .A(n20115), .ZN(P3_U2769) );
  AOI22_X1 U22216 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n20152), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n20158), .ZN(n20116) );
  OAI21_X1 U22217 ( .B1(n20139), .B2(n20154), .A(n20116), .ZN(P3_U2770) );
  AOI22_X1 U22218 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n20159), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n20158), .ZN(n20117) );
  OAI21_X1 U22219 ( .B1(n20694), .B2(n20161), .A(n20117), .ZN(P3_U2771) );
  AOI22_X1 U22220 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n20152), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n20158), .ZN(n20118) );
  OAI21_X1 U22221 ( .B1(n20657), .B2(n20154), .A(n20118), .ZN(P3_U2772) );
  AOI22_X1 U22222 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(n20152), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n20158), .ZN(n20119) );
  OAI21_X1 U22223 ( .B1(n20649), .B2(n20154), .A(n20119), .ZN(P3_U2773) );
  AOI22_X1 U22224 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(n20152), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n20158), .ZN(n20120) );
  OAI21_X1 U22225 ( .B1(n20145), .B2(n20154), .A(n20120), .ZN(P3_U2774) );
  AOI22_X1 U22226 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n20159), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n20158), .ZN(n20121) );
  OAI21_X1 U22227 ( .B1(n20122), .B2(n20161), .A(n20121), .ZN(P3_U2775) );
  AOI22_X1 U22228 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n20159), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n20158), .ZN(n20123) );
  OAI21_X1 U22229 ( .B1(n20124), .B2(n20161), .A(n20123), .ZN(P3_U2776) );
  AOI22_X1 U22230 ( .A1(P3_EAX_REG_25__SCAN_IN), .A2(n20152), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n20158), .ZN(n20125) );
  OAI21_X1 U22231 ( .B1(n20637), .B2(n20154), .A(n20125), .ZN(P3_U2777) );
  AOI22_X1 U22232 ( .A1(P3_EAX_REG_26__SCAN_IN), .A2(n20152), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n20158), .ZN(n20126) );
  OAI21_X1 U22233 ( .B1(n20718), .B2(n20154), .A(n20126), .ZN(P3_U2778) );
  AOI22_X1 U22234 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n20159), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n20158), .ZN(n20127) );
  OAI21_X1 U22235 ( .B1(n20128), .B2(n20161), .A(n20127), .ZN(P3_U2779) );
  AOI22_X1 U22236 ( .A1(P3_EAX_REG_28__SCAN_IN), .A2(n20152), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n20158), .ZN(n20129) );
  OAI21_X1 U22237 ( .B1(n20624), .B2(n20154), .A(n20129), .ZN(P3_U2780) );
  AOI22_X1 U22238 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n20159), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n20158), .ZN(n20130) );
  OAI21_X1 U22239 ( .B1(n20131), .B2(n20161), .A(n20130), .ZN(P3_U2781) );
  AOI22_X1 U22240 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n20159), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n20158), .ZN(n20132) );
  OAI21_X1 U22241 ( .B1(n20133), .B2(n20161), .A(n20132), .ZN(P3_U2782) );
  AOI22_X1 U22242 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(n20152), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n20158), .ZN(n20134) );
  OAI21_X1 U22243 ( .B1(n20135), .B2(n20154), .A(n20134), .ZN(P3_U2783) );
  AOI22_X1 U22244 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n20159), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n20158), .ZN(n20136) );
  OAI21_X1 U22245 ( .B1(n20137), .B2(n20161), .A(n20136), .ZN(P3_U2784) );
  AOI22_X1 U22246 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(n20152), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n20158), .ZN(n20138) );
  OAI21_X1 U22247 ( .B1(n20139), .B2(n20154), .A(n20138), .ZN(P3_U2785) );
  AOI22_X1 U22248 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n20159), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n20158), .ZN(n20140) );
  OAI21_X1 U22249 ( .B1(n20141), .B2(n20161), .A(n20140), .ZN(P3_U2786) );
  AOI22_X1 U22250 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(n20152), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n20158), .ZN(n20142) );
  OAI21_X1 U22251 ( .B1(n20657), .B2(n20154), .A(n20142), .ZN(P3_U2787) );
  AOI22_X1 U22252 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n20152), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n20158), .ZN(n20143) );
  OAI21_X1 U22253 ( .B1(n20649), .B2(n20154), .A(n20143), .ZN(P3_U2788) );
  AOI22_X1 U22254 ( .A1(P3_EAX_REG_6__SCAN_IN), .A2(n20152), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n20158), .ZN(n20144) );
  OAI21_X1 U22255 ( .B1(n20145), .B2(n20154), .A(n20144), .ZN(P3_U2789) );
  AOI22_X1 U22256 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n20159), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n20158), .ZN(n20146) );
  OAI21_X1 U22257 ( .B1(n20147), .B2(n20161), .A(n20146), .ZN(P3_U2790) );
  AOI22_X1 U22258 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n20159), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n20158), .ZN(n20148) );
  OAI21_X1 U22259 ( .B1(n20777), .B2(n20161), .A(n20148), .ZN(P3_U2791) );
  AOI22_X1 U22260 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(n20152), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n20158), .ZN(n20149) );
  OAI21_X1 U22261 ( .B1(n20637), .B2(n20154), .A(n20149), .ZN(P3_U2792) );
  AOI22_X1 U22262 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n20152), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n20158), .ZN(n20150) );
  OAI21_X1 U22263 ( .B1(n20718), .B2(n20154), .A(n20150), .ZN(P3_U2793) );
  AOI22_X1 U22264 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n20159), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n20158), .ZN(n20151) );
  OAI21_X1 U22265 ( .B1(n20627), .B2(n20161), .A(n20151), .ZN(P3_U2794) );
  AOI22_X1 U22266 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n20152), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n20158), .ZN(n20153) );
  OAI21_X1 U22267 ( .B1(n20624), .B2(n20154), .A(n20153), .ZN(P3_U2795) );
  AOI22_X1 U22268 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n20159), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n20158), .ZN(n20155) );
  OAI21_X1 U22269 ( .B1(n20670), .B2(n20161), .A(n20155), .ZN(P3_U2796) );
  AOI22_X1 U22270 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n20159), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n20158), .ZN(n20156) );
  OAI21_X1 U22271 ( .B1(n20157), .B2(n20161), .A(n20156), .ZN(P3_U2797) );
  AOI22_X1 U22272 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n20159), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n20158), .ZN(n20160) );
  OAI21_X1 U22273 ( .B1(n20770), .B2(n20161), .A(n20160), .ZN(P3_U2798) );
  INV_X1 U22274 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n20276) );
  NOR4_X1 U22275 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(P3_STATE2_REG_2__SCAN_IN), .A3(P3_STATEBS16_REG_SCAN_IN), .A4(n20798), .ZN(n20450) );
  OAI21_X1 U22276 ( .B1(n20391), .B2(n20276), .A(n20450), .ZN(n20278) );
  INV_X1 U22277 ( .A(n20450), .ZN(n21293) );
  AND2_X1 U22278 ( .A1(n21290), .A2(n20162), .ZN(n21303) );
  NOR4_X4 U22279 ( .A1(n21238), .A2(n20165), .A3(n20579), .A4(n21303), .ZN(
        n20513) );
  AOI21_X1 U22280 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n20593), .A(
        n20585), .ZN(n20178) );
  INV_X1 U22281 ( .A(n20163), .ZN(n20801) );
  NOR2_X1 U22282 ( .A1(n20801), .A2(n20180), .ZN(n20800) );
  OAI211_X1 U22283 ( .C1(n20171), .C2(n20164), .A(n21755), .B(n21700), .ZN(
        n20167) );
  INV_X1 U22284 ( .A(n20167), .ZN(n21287) );
  AOI211_X4 U22285 ( .C1(P3_EBX_REG_31__SCAN_IN), .C2(n20171), .A(n21287), .B(
        n20169), .ZN(n20604) );
  OAI22_X1 U22286 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n20600), .B1(n20561), 
        .B2(n20168), .ZN(n20176) );
  INV_X1 U22287 ( .A(n20169), .ZN(n20172) );
  NAND2_X1 U22288 ( .A1(n21755), .A2(n21700), .ZN(n20170) );
  INV_X1 U22289 ( .A(n20513), .ZN(n20605) );
  OAI22_X1 U22290 ( .A1(n20554), .A2(n20174), .B1(n20173), .B2(n20605), .ZN(
        n20175) );
  AOI211_X1 U22291 ( .C1(n20800), .C2(n20601), .A(n20176), .B(n20175), .ZN(
        n20177) );
  OAI221_X1 U22292 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n20278), .C1(
        n20186), .C2(n20178), .A(n20177), .ZN(P3_U2670) );
  NAND2_X1 U22293 ( .A1(n20579), .A2(n20391), .ZN(n20427) );
  NOR2_X1 U22294 ( .A1(n20179), .A2(P3_EBX_REG_2__SCAN_IN), .ZN(n20194) );
  AOI211_X1 U22295 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n20179), .A(n20194), .B(
        n20554), .ZN(n20185) );
  INV_X1 U22296 ( .A(n20180), .ZN(n20810) );
  NAND2_X1 U22297 ( .A1(n20822), .A2(n20810), .ZN(n20827) );
  INV_X1 U22298 ( .A(n20827), .ZN(n20826) );
  NOR2_X1 U22299 ( .A1(n20181), .A2(n20826), .ZN(n20814) );
  AOI22_X1 U22300 ( .A1(P3_REIP_REG_2__SCAN_IN), .A2(n20513), .B1(n20814), 
        .B2(n20601), .ZN(n20183) );
  NAND2_X1 U22301 ( .A1(P3_REIP_REG_2__SCAN_IN), .A2(P3_REIP_REG_1__SCAN_IN), 
        .ZN(n20205) );
  OAI211_X1 U22302 ( .C1(P3_REIP_REG_2__SCAN_IN), .C2(P3_REIP_REG_1__SCAN_IN), 
        .A(n20530), .B(n20205), .ZN(n20182) );
  OAI211_X1 U22303 ( .C1(n20558), .C2(n20187), .A(n20183), .B(n20182), .ZN(
        n20184) );
  AOI211_X1 U22304 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n20604), .A(n20185), .B(
        n20184), .ZN(n20190) );
  NOR2_X1 U22305 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n20186), .ZN(
        n20309) );
  INV_X1 U22306 ( .A(n20309), .ZN(n20188) );
  OAI221_X1 U22307 ( .B1(n20309), .B2(n20191), .C1(n20188), .C2(n20187), .A(
        n20593), .ZN(n20189) );
  OAI211_X1 U22308 ( .C1(n20191), .C2(n20427), .A(n20190), .B(n20189), .ZN(
        P3_U2669) );
  NAND3_X1 U22309 ( .A1(P3_REIP_REG_3__SCAN_IN), .A2(P3_REIP_REG_2__SCAN_IN), 
        .A3(P3_REIP_REG_1__SCAN_IN), .ZN(n20222) );
  NAND2_X1 U22310 ( .A1(n20507), .A2(n20222), .ZN(n20204) );
  OAI21_X1 U22311 ( .B1(n20829), .B2(n20192), .A(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n20832) );
  NAND2_X1 U22312 ( .A1(n20832), .A2(n20193), .ZN(n20840) );
  AOI22_X1 U22313 ( .A1(n20604), .A2(P3_EBX_REG_3__SCAN_IN), .B1(n20601), .B2(
        n20840), .ZN(n20203) );
  INV_X1 U22314 ( .A(n20194), .ZN(n20195) );
  NOR2_X1 U22315 ( .A1(P3_EBX_REG_3__SCAN_IN), .A2(n20195), .ZN(n20210) );
  AOI211_X1 U22316 ( .C1(P3_EBX_REG_3__SCAN_IN), .C2(n20195), .A(n20210), .B(
        n20554), .ZN(n20201) );
  AOI21_X1 U22317 ( .B1(n20530), .B2(n20222), .A(n20513), .ZN(n20212) );
  AOI21_X1 U22318 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n20309), .A(
        n20391), .ZN(n20196) );
  XNOR2_X1 U22319 ( .A(n20197), .B(n20196), .ZN(n20198) );
  OAI22_X1 U22320 ( .A1(n20212), .A2(n20199), .B1(n21293), .B2(n20198), .ZN(
        n20200) );
  AOI211_X1 U22321 ( .C1(n20585), .C2(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .A(
        n20201), .B(n20200), .ZN(n20202) );
  OAI211_X1 U22322 ( .C1(n20205), .C2(n20204), .A(n20203), .B(n20202), .ZN(
        P3_U2668) );
  NOR3_X1 U22323 ( .A1(P3_REIP_REG_4__SCAN_IN), .A2(n20600), .A3(n20222), .ZN(
        n20206) );
  AOI211_X1 U22324 ( .C1(n20604), .C2(P3_EBX_REG_4__SCAN_IN), .A(n21238), .B(
        n20206), .ZN(n20220) );
  INV_X1 U22325 ( .A(n20207), .ZN(n20208) );
  AOI211_X1 U22326 ( .C1(n20577), .C2(n20208), .A(n20278), .B(n20215), .ZN(
        n20214) );
  INV_X1 U22327 ( .A(P3_EBX_REG_4__SCAN_IN), .ZN(n20209) );
  NAND2_X1 U22328 ( .A1(n20210), .A2(n20209), .ZN(n20221) );
  OAI211_X1 U22329 ( .C1(n20210), .C2(n20209), .A(n20603), .B(n20221), .ZN(
        n20211) );
  OAI21_X1 U22330 ( .B1(n20212), .B2(n20907), .A(n20211), .ZN(n20213) );
  AOI211_X1 U22331 ( .C1(n20585), .C2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n20214), .B(n20213), .ZN(n20219) );
  OAI211_X1 U22332 ( .C1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .C2(n20224), .A(
        n20593), .B(n20215), .ZN(n20218) );
  OAI21_X1 U22333 ( .B1(n20216), .B2(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(
        n20601), .ZN(n20217) );
  NAND4_X1 U22334 ( .A1(n20220), .A2(n20219), .A3(n20218), .A4(n20217), .ZN(
        P3_U2667) );
  INV_X1 U22335 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n20232) );
  NOR2_X1 U22336 ( .A1(P3_EBX_REG_5__SCAN_IN), .A2(n20221), .ZN(n20242) );
  AOI211_X1 U22337 ( .C1(P3_EBX_REG_5__SCAN_IN), .C2(n20221), .A(n20242), .B(
        n20554), .ZN(n20230) );
  NOR2_X1 U22338 ( .A1(n20907), .A2(n20222), .ZN(n20223) );
  AOI21_X1 U22339 ( .B1(n20530), .B2(n20223), .A(P3_REIP_REG_5__SCAN_IN), .ZN(
        n20228) );
  NAND2_X1 U22340 ( .A1(P3_REIP_REG_5__SCAN_IN), .A2(n20223), .ZN(n20249) );
  AOI21_X1 U22341 ( .B1(n20530), .B2(n20249), .A(n20513), .ZN(n20256) );
  OAI21_X1 U22342 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n20224), .A(
        n20577), .ZN(n20225) );
  XOR2_X1 U22343 ( .A(n20226), .B(n20225), .Z(n20227) );
  OAI22_X1 U22344 ( .A1(n20228), .A2(n20256), .B1(n21293), .B2(n20227), .ZN(
        n20229) );
  AOI211_X1 U22345 ( .C1(n20585), .C2(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .A(
        n20230), .B(n20229), .ZN(n20231) );
  OAI211_X1 U22346 ( .C1(n20561), .C2(n20232), .A(n20231), .B(n21223), .ZN(
        P3_U2666) );
  OAI22_X1 U22347 ( .A1(n20233), .A2(n20558), .B1(n20250), .B2(n20256), .ZN(
        n20240) );
  NOR2_X1 U22348 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n21293), .ZN(
        n20335) );
  INV_X1 U22349 ( .A(n20427), .ZN(n20333) );
  AOI21_X1 U22350 ( .B1(n20234), .B2(n20335), .A(n20333), .ZN(n20238) );
  NAND2_X1 U22351 ( .A1(n20245), .A2(n20309), .ZN(n20235) );
  NAND3_X1 U22352 ( .A1(n20593), .A2(n20235), .A3(n20237), .ZN(n20236) );
  OAI21_X1 U22353 ( .B1(n20238), .B2(n20237), .A(n20236), .ZN(n20239) );
  AOI211_X1 U22354 ( .C1(n20604), .C2(P3_EBX_REG_6__SCAN_IN), .A(n20240), .B(
        n20239), .ZN(n20244) );
  OR3_X1 U22355 ( .A1(P3_REIP_REG_6__SCAN_IN), .A2(n20600), .A3(n20249), .ZN(
        n20255) );
  INV_X1 U22356 ( .A(P3_EBX_REG_6__SCAN_IN), .ZN(n20241) );
  NAND2_X1 U22357 ( .A1(n20242), .A2(n20241), .ZN(n20248) );
  OAI211_X1 U22358 ( .C1(n20242), .C2(n20241), .A(n20603), .B(n20248), .ZN(
        n20243) );
  NAND4_X1 U22359 ( .A1(n20244), .A2(n21223), .A3(n20255), .A4(n20243), .ZN(
        P3_U2665) );
  AOI21_X1 U22360 ( .B1(n20245), .B2(n20309), .A(n20391), .ZN(n20246) );
  XNOR2_X1 U22361 ( .A(n20247), .B(n20246), .ZN(n20260) );
  NOR2_X1 U22362 ( .A1(P3_EBX_REG_7__SCAN_IN), .A2(n20248), .ZN(n20272) );
  AOI211_X1 U22363 ( .C1(P3_EBX_REG_7__SCAN_IN), .C2(n20248), .A(n20272), .B(
        n20554), .ZN(n20253) );
  NOR2_X1 U22364 ( .A1(n20250), .A2(n20249), .ZN(n20261) );
  NAND3_X1 U22365 ( .A1(n20507), .A2(n20261), .A3(n20254), .ZN(n20251) );
  OAI211_X1 U22366 ( .C1(n11231), .C2(n20558), .A(n21223), .B(n20251), .ZN(
        n20252) );
  AOI211_X1 U22367 ( .C1(P3_EBX_REG_7__SCAN_IN), .C2(n20604), .A(n20253), .B(
        n20252), .ZN(n20259) );
  AOI21_X1 U22368 ( .B1(n20256), .B2(n20255), .A(n20254), .ZN(n20257) );
  INV_X1 U22369 ( .A(n20257), .ZN(n20258) );
  OAI211_X1 U22370 ( .C1(n21293), .C2(n20260), .A(n20259), .B(n20258), .ZN(
        P3_U2664) );
  NAND2_X1 U22371 ( .A1(P3_REIP_REG_7__SCAN_IN), .A2(n20261), .ZN(n20263) );
  NOR2_X1 U22372 ( .A1(n20938), .A2(n20263), .ZN(n20294) );
  NOR2_X1 U22373 ( .A1(n20600), .A2(n20294), .ZN(n20265) );
  INV_X1 U22374 ( .A(n20265), .ZN(n20262) );
  OAI22_X1 U22375 ( .A1(n20264), .A2(n20558), .B1(n20263), .B2(n20262), .ZN(
        n20271) );
  NOR2_X1 U22376 ( .A1(n20513), .A2(n20265), .ZN(n20304) );
  AOI21_X1 U22377 ( .B1(n20266), .B2(n20276), .A(n20391), .ZN(n20268) );
  XOR2_X1 U22378 ( .A(n20268), .B(n20267), .Z(n20269) );
  OAI22_X1 U22379 ( .A1(n20304), .A2(n20938), .B1(n21293), .B2(n20269), .ZN(
        n20270) );
  NOR3_X1 U22380 ( .A1(n21238), .A2(n20271), .A3(n20270), .ZN(n20274) );
  NAND2_X1 U22381 ( .A1(n20272), .A2(n20275), .ZN(n20280) );
  OAI211_X1 U22382 ( .C1(n20272), .C2(n20275), .A(n20603), .B(n20280), .ZN(
        n20273) );
  OAI211_X1 U22383 ( .C1(n20275), .C2(n20561), .A(n20274), .B(n20273), .ZN(
        P3_U2663) );
  AOI21_X1 U22384 ( .B1(n20277), .B2(n20276), .A(n20391), .ZN(n20292) );
  NAND2_X1 U22385 ( .A1(n20579), .A2(n20292), .ZN(n20289) );
  AOI21_X1 U22386 ( .B1(n20577), .B2(n20279), .A(n20278), .ZN(n20287) );
  NOR2_X1 U22387 ( .A1(P3_EBX_REG_9__SCAN_IN), .A2(n20280), .ZN(n20296) );
  AOI21_X1 U22388 ( .B1(n20280), .B2(P3_EBX_REG_9__SCAN_IN), .A(n20554), .ZN(
        n20281) );
  AOI21_X1 U22389 ( .B1(P3_EBX_REG_9__SCAN_IN), .B2(n20604), .A(n20281), .ZN(
        n20282) );
  OAI22_X1 U22390 ( .A1(n20296), .A2(n20282), .B1(n20304), .B2(n20283), .ZN(
        n20286) );
  NAND3_X1 U22391 ( .A1(n20507), .A2(n20294), .A3(n20283), .ZN(n20303) );
  OAI211_X1 U22392 ( .C1(n20284), .C2(n20558), .A(n21223), .B(n20303), .ZN(
        n20285) );
  AOI211_X1 U22393 ( .C1(n20290), .C2(n20287), .A(n20286), .B(n20285), .ZN(
        n20288) );
  OAI21_X1 U22394 ( .B1(n20290), .B2(n20289), .A(n20288), .ZN(P3_U2662) );
  XNOR2_X1 U22395 ( .A(n20292), .B(n20291), .ZN(n20301) );
  OAI22_X1 U22396 ( .A1(n20561), .A2(n20295), .B1(n20293), .B2(n20558), .ZN(
        n20300) );
  NAND2_X1 U22397 ( .A1(P3_REIP_REG_9__SCAN_IN), .A2(n20294), .ZN(n20305) );
  NAND2_X1 U22398 ( .A1(n20507), .A2(n20306), .ZN(n20298) );
  NAND2_X1 U22399 ( .A1(n20296), .A2(n20295), .ZN(n20308) );
  OAI211_X1 U22400 ( .C1(n20296), .C2(n20295), .A(n20603), .B(n20308), .ZN(
        n20297) );
  OAI211_X1 U22401 ( .C1(n20305), .C2(n20298), .A(n21223), .B(n20297), .ZN(
        n20299) );
  AOI211_X1 U22402 ( .C1(n20579), .C2(n20301), .A(n20300), .B(n20299), .ZN(
        n20302) );
  OAI221_X1 U22403 ( .B1(n20306), .B2(n20304), .C1(n20306), .C2(n20303), .A(
        n20302), .ZN(P3_U2661) );
  NOR2_X1 U22404 ( .A1(n20306), .A2(n20305), .ZN(n20307) );
  AOI21_X1 U22405 ( .B1(n20507), .B2(n20307), .A(P3_REIP_REG_11__SCAN_IN), 
        .ZN(n20320) );
  NAND2_X1 U22406 ( .A1(P3_REIP_REG_11__SCAN_IN), .A2(n20307), .ZN(n20339) );
  AOI21_X1 U22407 ( .B1(n20339), .B2(n20530), .A(n20513), .ZN(n20338) );
  NOR2_X1 U22408 ( .A1(P3_EBX_REG_11__SCAN_IN), .A2(n20308), .ZN(n20330) );
  AOI211_X1 U22409 ( .C1(P3_EBX_REG_11__SCAN_IN), .C2(n20308), .A(n20330), .B(
        n20554), .ZN(n20318) );
  NAND2_X1 U22410 ( .A1(n20310), .A2(n20309), .ZN(n20312) );
  NOR2_X1 U22411 ( .A1(n20311), .A2(n20312), .ZN(n20347) );
  NOR2_X1 U22412 ( .A1(n20347), .A2(n20391), .ZN(n20323) );
  AOI21_X1 U22413 ( .B1(n20314), .B2(n20312), .A(n21293), .ZN(n20313) );
  OAI22_X1 U22414 ( .A1(n20314), .A2(n20323), .B1(n20333), .B2(n20313), .ZN(
        n20315) );
  OAI211_X1 U22415 ( .C1(n20561), .C2(n20316), .A(n21223), .B(n20315), .ZN(
        n20317) );
  AOI211_X1 U22416 ( .C1(n20585), .C2(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .A(
        n20318), .B(n20317), .ZN(n20319) );
  OAI21_X1 U22417 ( .B1(n20320), .B2(n20338), .A(n20319), .ZN(P3_U2660) );
  INV_X1 U22418 ( .A(n20338), .ZN(n20328) );
  INV_X1 U22419 ( .A(n20322), .ZN(n20324) );
  INV_X1 U22420 ( .A(n20323), .ZN(n20321) );
  AOI221_X1 U22421 ( .B1(n20324), .B2(n20323), .C1(n20322), .C2(n20321), .A(
        n21293), .ZN(n20327) );
  INV_X1 U22422 ( .A(P3_EBX_REG_12__SCAN_IN), .ZN(n20329) );
  OAI22_X1 U22423 ( .A1(n20561), .A2(n20329), .B1(n20325), .B2(n20558), .ZN(
        n20326) );
  AOI211_X1 U22424 ( .C1(n20328), .C2(P3_REIP_REG_12__SCAN_IN), .A(n20327), 
        .B(n20326), .ZN(n20332) );
  OR3_X1 U22425 ( .A1(n20600), .A2(n20339), .A3(P3_REIP_REG_12__SCAN_IN), .ZN(
        n20337) );
  NAND2_X1 U22426 ( .A1(n20330), .A2(n20329), .ZN(n20341) );
  OAI211_X1 U22427 ( .C1(n20330), .C2(n20329), .A(n20603), .B(n20341), .ZN(
        n20331) );
  NAND4_X1 U22428 ( .A1(n20332), .A2(n21223), .A3(n20337), .A4(n20331), .ZN(
        P3_U2659) );
  INV_X1 U22429 ( .A(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n20334) );
  AOI21_X1 U22430 ( .B1(n20335), .B2(n20334), .A(n20333), .ZN(n20351) );
  AOI21_X1 U22431 ( .B1(n20338), .B2(n20337), .A(n20336), .ZN(n20346) );
  NOR2_X1 U22432 ( .A1(n20340), .A2(n20339), .ZN(n20363) );
  NAND2_X1 U22433 ( .A1(n20530), .A2(n20363), .ZN(n20344) );
  NOR2_X1 U22434 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(n20341), .ZN(n20356) );
  AOI211_X1 U22435 ( .C1(P3_EBX_REG_13__SCAN_IN), .C2(n20341), .A(n20356), .B(
        n20554), .ZN(n20342) );
  AOI211_X1 U22436 ( .C1(n20604), .C2(P3_EBX_REG_13__SCAN_IN), .A(n21238), .B(
        n20342), .ZN(n20343) );
  OAI21_X1 U22437 ( .B1(P3_REIP_REG_13__SCAN_IN), .B2(n20344), .A(n20343), 
        .ZN(n20345) );
  AOI211_X1 U22438 ( .C1(n20585), .C2(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A(
        n20346), .B(n20345), .ZN(n20349) );
  NAND3_X1 U22439 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A3(n20347), .ZN(n20364) );
  NAND3_X1 U22440 ( .A1(n20593), .A2(n20364), .A3(n20350), .ZN(n20348) );
  OAI211_X1 U22441 ( .C1(n20351), .C2(n20350), .A(n20349), .B(n20348), .ZN(
        P3_U2658) );
  NAND2_X1 U22442 ( .A1(n20577), .A2(n20364), .ZN(n20352) );
  XNOR2_X1 U22443 ( .A(n20353), .B(n20352), .ZN(n20360) );
  NAND3_X1 U22444 ( .A1(n20530), .A2(P3_REIP_REG_13__SCAN_IN), .A3(n20363), 
        .ZN(n20354) );
  NAND3_X1 U22445 ( .A1(P3_REIP_REG_13__SCAN_IN), .A2(P3_REIP_REG_14__SCAN_IN), 
        .A3(n20363), .ZN(n20396) );
  AOI21_X1 U22446 ( .B1(n20530), .B2(n20396), .A(n20513), .ZN(n20390) );
  AOI21_X1 U22447 ( .B1(n20355), .B2(n20354), .A(n20390), .ZN(n20359) );
  NAND2_X1 U22448 ( .A1(n20356), .A2(n20362), .ZN(n20369) );
  OAI211_X1 U22449 ( .C1(n20356), .C2(n20362), .A(n20603), .B(n20369), .ZN(
        n20357) );
  OAI21_X1 U22450 ( .B1(n20558), .B2(n20365), .A(n20357), .ZN(n20358) );
  AOI211_X1 U22451 ( .C1(n20579), .C2(n20360), .A(n20359), .B(n20358), .ZN(
        n20361) );
  OAI211_X1 U22452 ( .C1(n20561), .C2(n20362), .A(n20361), .B(n21223), .ZN(
        P3_U2657) );
  NAND4_X1 U22453 ( .A1(n20530), .A2(P3_REIP_REG_13__SCAN_IN), .A3(
        P3_REIP_REG_14__SCAN_IN), .A4(n20363), .ZN(n20404) );
  NOR2_X1 U22454 ( .A1(n20365), .A2(n20364), .ZN(n20393) );
  OR2_X1 U22455 ( .A1(n20391), .A2(n20393), .ZN(n20367) );
  OAI21_X1 U22456 ( .B1(n20368), .B2(n20367), .A(n20579), .ZN(n20366) );
  AOI21_X1 U22457 ( .B1(n20368), .B2(n20367), .A(n20366), .ZN(n20374) );
  NOR2_X1 U22458 ( .A1(P3_EBX_REG_15__SCAN_IN), .A2(n20369), .ZN(n20381) );
  AOI211_X1 U22459 ( .C1(P3_EBX_REG_15__SCAN_IN), .C2(n20369), .A(n20381), .B(
        n20554), .ZN(n20373) );
  OAI22_X1 U22460 ( .A1(n20561), .A2(n20371), .B1(n20370), .B2(n20558), .ZN(
        n20372) );
  NOR4_X1 U22461 ( .A1(n21238), .A2(n20374), .A3(n20373), .A4(n20372), .ZN(
        n20375) );
  OAI221_X1 U22462 ( .B1(P3_REIP_REG_15__SCAN_IN), .B2(n20404), .C1(n20376), 
        .C2(n20390), .A(n20375), .ZN(P3_U2656) );
  NAND2_X1 U22463 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n20393), .ZN(
        n20422) );
  INV_X1 U22464 ( .A(n20422), .ZN(n20425) );
  NOR2_X1 U22465 ( .A1(n20425), .A2(n20391), .ZN(n20379) );
  OAI21_X1 U22466 ( .B1(n20379), .B2(n20378), .A(n20579), .ZN(n20377) );
  AOI21_X1 U22467 ( .B1(n20379), .B2(n20378), .A(n20377), .ZN(n20385) );
  INV_X1 U22468 ( .A(P3_EBX_REG_16__SCAN_IN), .ZN(n20380) );
  NAND2_X1 U22469 ( .A1(n20381), .A2(n20380), .ZN(n20398) );
  OAI211_X1 U22470 ( .C1(n20381), .C2(n20380), .A(n20603), .B(n20398), .ZN(
        n20382) );
  OAI211_X1 U22471 ( .C1(n20383), .C2(n20558), .A(n21223), .B(n20382), .ZN(
        n20384) );
  AOI211_X1 U22472 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n20604), .A(n20385), .B(
        n20384), .ZN(n20388) );
  INV_X1 U22473 ( .A(n20404), .ZN(n20386) );
  NAND2_X1 U22474 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(P3_REIP_REG_15__SCAN_IN), 
        .ZN(n20405) );
  OAI211_X1 U22475 ( .C1(P3_REIP_REG_16__SCAN_IN), .C2(P3_REIP_REG_15__SCAN_IN), .A(n20386), .B(n20405), .ZN(n20387) );
  OAI211_X1 U22476 ( .C1(n20390), .C2(n20389), .A(n20388), .B(n20387), .ZN(
        P3_U2655) );
  AOI21_X1 U22477 ( .B1(n20393), .B2(n20392), .A(n20391), .ZN(n20394) );
  XOR2_X1 U22478 ( .A(n20395), .B(n20394), .Z(n20403) );
  AOI21_X1 U22479 ( .B1(n20604), .B2(P3_EBX_REG_17__SCAN_IN), .A(n21238), .ZN(
        n20402) );
  NOR3_X1 U22480 ( .A1(n21190), .A2(n20396), .A3(n20405), .ZN(n20420) );
  INV_X1 U22481 ( .A(n20420), .ZN(n20397) );
  AOI21_X1 U22482 ( .B1(n20530), .B2(n20397), .A(n20513), .ZN(n20417) );
  AOI221_X1 U22483 ( .B1(n20405), .B2(n21190), .C1(n20404), .C2(n21190), .A(
        n20417), .ZN(n20400) );
  NOR2_X1 U22484 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n20398), .ZN(n20411) );
  AOI211_X1 U22485 ( .C1(P3_EBX_REG_17__SCAN_IN), .C2(n20398), .A(n20411), .B(
        n20554), .ZN(n20399) );
  AOI211_X1 U22486 ( .C1(n20585), .C2(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .A(
        n20400), .B(n20399), .ZN(n20401) );
  OAI211_X1 U22487 ( .C1(n21293), .C2(n20403), .A(n20402), .B(n20401), .ZN(
        P3_U2654) );
  NOR3_X1 U22488 ( .A1(n21190), .A2(n20405), .A3(n20404), .ZN(n20421) );
  INV_X1 U22489 ( .A(n20421), .ZN(n20419) );
  OAI21_X1 U22490 ( .B1(n20422), .B2(n20406), .A(n20577), .ZN(n20408) );
  OAI21_X1 U22491 ( .B1(n20409), .B2(n20408), .A(n20579), .ZN(n20407) );
  AOI21_X1 U22492 ( .B1(n20409), .B2(n20408), .A(n20407), .ZN(n20415) );
  INV_X1 U22493 ( .A(P3_EBX_REG_18__SCAN_IN), .ZN(n20410) );
  NAND2_X1 U22494 ( .A1(n20411), .A2(n20410), .ZN(n20429) );
  OAI211_X1 U22495 ( .C1(n20411), .C2(n20410), .A(n20603), .B(n20429), .ZN(
        n20412) );
  OAI211_X1 U22496 ( .C1(n20413), .C2(n20558), .A(n21223), .B(n20412), .ZN(
        n20414) );
  AOI211_X1 U22497 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n20604), .A(n20415), .B(
        n20414), .ZN(n20416) );
  OAI221_X1 U22498 ( .B1(P3_REIP_REG_18__SCAN_IN), .B2(n20419), .C1(n20418), 
        .C2(n20417), .A(n20416), .ZN(P3_U2653) );
  NAND3_X1 U22499 ( .A1(P3_REIP_REG_18__SCAN_IN), .A2(P3_REIP_REG_19__SCAN_IN), 
        .A3(n20420), .ZN(n20445) );
  AOI21_X1 U22500 ( .B1(n20530), .B2(n20445), .A(n20513), .ZN(n20444) );
  AOI21_X1 U22501 ( .B1(P3_REIP_REG_18__SCAN_IN), .B2(n20421), .A(
        P3_REIP_REG_19__SCAN_IN), .ZN(n20434) );
  AOI21_X1 U22502 ( .B1(n20604), .B2(P3_EBX_REG_19__SCAN_IN), .A(n21238), .ZN(
        n20433) );
  OAI21_X1 U22503 ( .B1(n20423), .B2(n20422), .A(n20577), .ZN(n20436) );
  OAI221_X1 U22504 ( .B1(n20428), .B2(n20425), .C1(n20428), .C2(n20424), .A(
        n20450), .ZN(n20426) );
  AOI22_X1 U22505 ( .A1(n20436), .A2(n20428), .B1(n20427), .B2(n20426), .ZN(
        n20431) );
  NOR2_X1 U22506 ( .A1(P3_EBX_REG_19__SCAN_IN), .A2(n20429), .ZN(n20437) );
  AOI211_X1 U22507 ( .C1(P3_EBX_REG_19__SCAN_IN), .C2(n20429), .A(n20437), .B(
        n20554), .ZN(n20430) );
  AOI211_X1 U22508 ( .C1(n20585), .C2(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n20431), .B(n20430), .ZN(n20432) );
  OAI211_X1 U22509 ( .C1(n20444), .C2(n20434), .A(n20433), .B(n20432), .ZN(
        P3_U2652) );
  NOR3_X1 U22510 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(n20600), .A3(n20445), 
        .ZN(n20442) );
  NAND2_X1 U22511 ( .A1(n20436), .A2(n20435), .ZN(n20449) );
  OAI211_X1 U22512 ( .C1(n20436), .C2(n20435), .A(n20579), .B(n20449), .ZN(
        n20439) );
  NAND2_X1 U22513 ( .A1(n20437), .A2(n20440), .ZN(n20448) );
  OAI211_X1 U22514 ( .C1(n20437), .C2(n20440), .A(n20603), .B(n20448), .ZN(
        n20438) );
  OAI211_X1 U22515 ( .C1(n20440), .C2(n20561), .A(n20439), .B(n20438), .ZN(
        n20441) );
  AOI211_X1 U22516 ( .C1(n20585), .C2(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n20442), .B(n20441), .ZN(n20443) );
  OAI21_X1 U22517 ( .B1(n20444), .B2(n20446), .A(n20443), .ZN(P3_U2651) );
  NOR2_X1 U22518 ( .A1(n20446), .A2(n20445), .ZN(n20459) );
  INV_X1 U22519 ( .A(n20459), .ZN(n20447) );
  AOI21_X1 U22520 ( .B1(n20507), .B2(n20447), .A(n20513), .ZN(n20470) );
  NOR2_X1 U22521 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n20448), .ZN(n20463) );
  AOI211_X1 U22522 ( .C1(P3_EBX_REG_21__SCAN_IN), .C2(n20448), .A(n20463), .B(
        n20554), .ZN(n20456) );
  NAND3_X1 U22523 ( .A1(n20530), .A2(n20459), .A3(n20458), .ZN(n20471) );
  OAI211_X1 U22524 ( .C1(n20452), .C2(n20451), .A(n20450), .B(n20460), .ZN(
        n20453) );
  OAI211_X1 U22525 ( .C1(n20454), .C2(n20561), .A(n20471), .B(n20453), .ZN(
        n20455) );
  AOI211_X1 U22526 ( .C1(n20585), .C2(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A(
        n20456), .B(n20455), .ZN(n20457) );
  OAI21_X1 U22527 ( .B1(n20458), .B2(n20470), .A(n20457), .ZN(P3_U2650) );
  NAND2_X1 U22528 ( .A1(P3_REIP_REG_21__SCAN_IN), .A2(n20459), .ZN(n20472) );
  NOR3_X1 U22529 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(n20600), .A3(n20472), 
        .ZN(n20468) );
  OAI211_X1 U22530 ( .C1(n20462), .C2(n20461), .A(n20579), .B(n20480), .ZN(
        n20465) );
  NAND2_X1 U22531 ( .A1(n20463), .A2(n20466), .ZN(n20477) );
  OAI211_X1 U22532 ( .C1(n20463), .C2(n20466), .A(n20603), .B(n20477), .ZN(
        n20464) );
  OAI211_X1 U22533 ( .C1(n20466), .C2(n20561), .A(n20465), .B(n20464), .ZN(
        n20467) );
  AOI211_X1 U22534 ( .C1(n20585), .C2(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n20468), .B(n20467), .ZN(n20469) );
  OAI221_X1 U22535 ( .B1(n20473), .B2(n20471), .C1(n20473), .C2(n20470), .A(
        n20469), .ZN(P3_U2649) );
  NOR2_X1 U22536 ( .A1(n20473), .A2(n20472), .ZN(n20474) );
  AOI21_X1 U22537 ( .B1(n20474), .B2(n20507), .A(P3_REIP_REG_23__SCAN_IN), 
        .ZN(n20476) );
  NAND2_X1 U22538 ( .A1(P3_REIP_REG_23__SCAN_IN), .A2(n20474), .ZN(n20504) );
  INV_X1 U22539 ( .A(n20504), .ZN(n20486) );
  OAI21_X1 U22540 ( .B1(n20486), .B2(n20600), .A(n20605), .ZN(n20499) );
  INV_X1 U22541 ( .A(n20499), .ZN(n20475) );
  NOR2_X1 U22542 ( .A1(n20476), .A2(n20475), .ZN(n20479) );
  NOR2_X1 U22543 ( .A1(P3_EBX_REG_23__SCAN_IN), .A2(n20477), .ZN(n20487) );
  AOI211_X1 U22544 ( .C1(P3_EBX_REG_23__SCAN_IN), .C2(n20477), .A(n20487), .B(
        n20554), .ZN(n20478) );
  AOI211_X1 U22545 ( .C1(P3_EBX_REG_23__SCAN_IN), .C2(n20604), .A(n20479), .B(
        n20478), .ZN(n20484) );
  NAND2_X1 U22546 ( .A1(n20577), .A2(n20480), .ZN(n20481) );
  NAND2_X1 U22547 ( .A1(n20482), .A2(n20481), .ZN(n20491) );
  OAI211_X1 U22548 ( .C1(n20482), .C2(n20481), .A(n20579), .B(n20491), .ZN(
        n20483) );
  OAI211_X1 U22549 ( .C1(n20558), .C2(n20485), .A(n20484), .B(n20483), .ZN(
        P3_U2648) );
  NOR2_X1 U22550 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n20600), .ZN(n20500) );
  AOI22_X1 U22551 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n20585), .B1(
        n20486), .B2(n20500), .ZN(n20496) );
  NAND2_X1 U22552 ( .A1(n20487), .A2(n20488), .ZN(n20497) );
  NOR2_X1 U22553 ( .A1(n20487), .A2(n20488), .ZN(n20489) );
  OAI22_X1 U22554 ( .A1(n20554), .A2(n20489), .B1(n20561), .B2(n20488), .ZN(
        n20490) );
  AOI22_X1 U22555 ( .A1(n20499), .A2(P3_REIP_REG_24__SCAN_IN), .B1(n20497), 
        .B2(n20490), .ZN(n20495) );
  NAND2_X1 U22556 ( .A1(n20577), .A2(n20491), .ZN(n20492) );
  NAND2_X1 U22557 ( .A1(n20493), .A2(n20492), .ZN(n20501) );
  OAI211_X1 U22558 ( .C1(n20493), .C2(n20492), .A(n20579), .B(n20501), .ZN(
        n20494) );
  NAND3_X1 U22559 ( .A1(n20496), .A2(n20495), .A3(n20494), .ZN(P3_U2647) );
  AOI22_X1 U22560 ( .A1(n20604), .A2(P3_EBX_REG_25__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n20585), .ZN(n20511) );
  NOR2_X1 U22561 ( .A1(P3_EBX_REG_25__SCAN_IN), .A2(n20497), .ZN(n20514) );
  AOI211_X1 U22562 ( .C1(P3_EBX_REG_25__SCAN_IN), .C2(n20497), .A(n20514), .B(
        n20554), .ZN(n20498) );
  AOI221_X1 U22563 ( .B1(n20500), .B2(P3_REIP_REG_25__SCAN_IN), .C1(n20499), 
        .C2(P3_REIP_REG_25__SCAN_IN), .A(n20498), .ZN(n20510) );
  NAND2_X1 U22564 ( .A1(n20577), .A2(n20501), .ZN(n20502) );
  OAI211_X1 U22565 ( .C1(n20503), .C2(n20502), .A(n20579), .B(n20523), .ZN(
        n20509) );
  NOR2_X1 U22566 ( .A1(n20505), .A2(n20504), .ZN(n20512) );
  NAND3_X1 U22567 ( .A1(n20507), .A2(n20512), .A3(n20506), .ZN(n20508) );
  NAND4_X1 U22568 ( .A1(n20511), .A2(n20510), .A3(n20509), .A4(n20508), .ZN(
        P3_U2646) );
  NAND2_X1 U22569 ( .A1(P3_REIP_REG_25__SCAN_IN), .A2(n20512), .ZN(n20519) );
  NOR2_X1 U22570 ( .A1(n20528), .A2(n20519), .ZN(n20529) );
  NOR2_X1 U22571 ( .A1(n20529), .A2(n20600), .ZN(n20517) );
  NOR2_X1 U22572 ( .A1(n20513), .A2(n20517), .ZN(n20553) );
  NAND2_X1 U22573 ( .A1(n20514), .A2(n20515), .ZN(n20531) );
  OAI211_X1 U22574 ( .C1(n20515), .C2(n20514), .A(n20531), .B(n20603), .ZN(
        n20516) );
  INV_X1 U22575 ( .A(n20516), .ZN(n20522) );
  INV_X1 U22576 ( .A(n20517), .ZN(n20518) );
  OAI22_X1 U22577 ( .A1(n20520), .A2(n20558), .B1(n20519), .B2(n20518), .ZN(
        n20521) );
  AOI211_X1 U22578 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n20604), .A(n20522), .B(
        n20521), .ZN(n20527) );
  OAI211_X1 U22579 ( .C1(n20525), .C2(n20524), .A(n20579), .B(n20534), .ZN(
        n20526) );
  OAI211_X1 U22580 ( .C1(n20553), .C2(n20528), .A(n20527), .B(n20526), .ZN(
        P3_U2645) );
  AOI22_X1 U22581 ( .A1(n20604), .A2(P3_EBX_REG_27__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n20585), .ZN(n20539) );
  NAND2_X1 U22582 ( .A1(n20530), .A2(n20529), .ZN(n20556) );
  OAI21_X1 U22583 ( .B1(P3_REIP_REG_27__SCAN_IN), .B2(n20556), .A(n20553), 
        .ZN(n20546) );
  INV_X1 U22584 ( .A(n20556), .ZN(n20580) );
  NOR2_X1 U22585 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(n20531), .ZN(n20540) );
  AOI211_X1 U22586 ( .C1(P3_EBX_REG_27__SCAN_IN), .C2(n20531), .A(n20540), .B(
        n20554), .ZN(n20532) );
  AOI221_X1 U22587 ( .B1(P3_REIP_REG_27__SCAN_IN), .B2(n20546), .C1(n20580), 
        .C2(n20546), .A(n20532), .ZN(n20538) );
  INV_X1 U22588 ( .A(n20533), .ZN(n20536) );
  NAND2_X1 U22589 ( .A1(n20536), .A2(n20535), .ZN(n20547) );
  OAI211_X1 U22590 ( .C1(n20536), .C2(n20535), .A(n20579), .B(n20547), .ZN(
        n20537) );
  NAND3_X1 U22591 ( .A1(n20539), .A2(n20538), .A3(n20537), .ZN(P3_U2644) );
  NAND2_X1 U22592 ( .A1(n20540), .A2(n20543), .ZN(n20555) );
  OAI21_X1 U22593 ( .B1(n20540), .B2(n20543), .A(n20555), .ZN(n20552) );
  NOR3_X1 U22594 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(n20541), .A3(n20556), 
        .ZN(n20545) );
  OAI22_X1 U22595 ( .A1(n20561), .A2(n20543), .B1(n20542), .B2(n20558), .ZN(
        n20544) );
  AOI211_X1 U22596 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(n20546), .A(n20545), 
        .B(n20544), .ZN(n20551) );
  NAND2_X1 U22597 ( .A1(n20577), .A2(n20547), .ZN(n20549) );
  OAI211_X1 U22598 ( .C1(n20549), .C2(n20548), .A(n20579), .B(n20565), .ZN(
        n20550) );
  OAI211_X1 U22599 ( .C1(n20552), .C2(n20554), .A(n20551), .B(n20550), .ZN(
        P3_U2643) );
  NAND2_X1 U22600 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .ZN(n20557) );
  NOR2_X1 U22601 ( .A1(n20570), .A2(n20557), .ZN(n20581) );
  OAI21_X1 U22602 ( .B1(n20581), .B2(n20600), .A(n20553), .ZN(n20571) );
  INV_X1 U22603 ( .A(n20571), .ZN(n20587) );
  NOR2_X1 U22604 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n20555), .ZN(n20573) );
  NOR2_X1 U22605 ( .A1(n20573), .A2(n20554), .ZN(n20572) );
  NAND2_X1 U22606 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n20555), .ZN(n20564) );
  NOR3_X1 U22607 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(n20557), .A3(n20556), 
        .ZN(n20563) );
  OAI22_X1 U22608 ( .A1(n20561), .A2(n20560), .B1(n20559), .B2(n20558), .ZN(
        n20562) );
  AOI211_X1 U22609 ( .C1(n20572), .C2(n20564), .A(n20563), .B(n20562), .ZN(
        n20569) );
  OAI211_X1 U22610 ( .C1(n20567), .C2(n20566), .A(n20579), .B(n20576), .ZN(
        n20568) );
  OAI211_X1 U22611 ( .C1(n20587), .C2(n20570), .A(n20569), .B(n20568), .ZN(
        P3_U2642) );
  AOI22_X1 U22612 ( .A1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n20585), .B1(
        P3_REIP_REG_30__SCAN_IN), .B2(n20571), .ZN(n20584) );
  INV_X1 U22613 ( .A(n20572), .ZN(n20575) );
  AND2_X1 U22614 ( .A1(n20603), .A2(n20573), .ZN(n20590) );
  NOR2_X1 U22615 ( .A1(n20604), .A2(n20590), .ZN(n20574) );
  MUX2_X1 U22616 ( .A(n20575), .B(n20574), .S(P3_EBX_REG_30__SCAN_IN), .Z(
        n20583) );
  NAND2_X1 U22617 ( .A1(n20592), .A2(n20591), .ZN(n20578) );
  OAI211_X1 U22618 ( .C1(n20592), .C2(n20591), .A(n20579), .B(n20578), .ZN(
        n20582) );
  NAND2_X1 U22619 ( .A1(n20595), .A2(n21088), .ZN(n20586) );
  NAND4_X1 U22620 ( .A1(n20584), .A2(n20583), .A3(n20582), .A4(n20586), .ZN(
        P3_U2641) );
  AOI22_X1 U22621 ( .A1(P3_EBX_REG_31__SCAN_IN), .A2(n20604), .B1(
        P3_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n20585), .ZN(n20599) );
  AOI21_X1 U22622 ( .B1(n20587), .B2(n20586), .A(n20594), .ZN(n20588) );
  AOI21_X1 U22623 ( .B1(n20590), .B2(n20589), .A(n20588), .ZN(n20598) );
  NAND3_X1 U22624 ( .A1(n20593), .A2(n20592), .A3(n20591), .ZN(n20597) );
  NAND3_X1 U22625 ( .A1(n20595), .A2(P3_REIP_REG_30__SCAN_IN), .A3(n20594), 
        .ZN(n20596) );
  NAND4_X1 U22626 ( .A1(n20599), .A2(n20598), .A3(n20597), .A4(n20596), .ZN(
        P3_U2640) );
  NAND2_X1 U22627 ( .A1(n20600), .A2(n20605), .ZN(n20602) );
  AOI22_X1 U22628 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(n20602), .B1(n20601), 
        .B2(n20829), .ZN(n20608) );
  OAI21_X1 U22629 ( .B1(n20604), .B2(n20603), .A(P3_EBX_REG_0__SCAN_IN), .ZN(
        n20607) );
  NAND3_X1 U22630 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n20605), .A3(
        n20802), .ZN(n20606) );
  NAND3_X1 U22631 ( .A1(n20608), .A2(n20607), .A3(n20606), .ZN(P3_U2671) );
  NOR2_X2 U22632 ( .A1(n20615), .A2(n20793), .ZN(n20794) );
  NAND2_X2 U22633 ( .A1(n20794), .A2(P3_EAX_REG_1__SCAN_IN), .ZN(n20784) );
  NOR2_X4 U22634 ( .A1(n20784), .A2(n20663), .ZN(n20662) );
  NOR2_X2 U22635 ( .A1(n20641), .A2(n20614), .ZN(n20638) );
  NOR2_X4 U22636 ( .A1(n20778), .A2(n20777), .ZN(n20775) );
  NAND2_X1 U22637 ( .A1(n20687), .A2(n20775), .ZN(n20632) );
  NAND2_X1 U22638 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n20636), .ZN(n20628) );
  NOR2_X1 U22639 ( .A1(n20627), .A2(n20628), .ZN(n20621) );
  NAND2_X1 U22640 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n20621), .ZN(n20620) );
  NAND2_X1 U22641 ( .A1(n20620), .A2(P3_EAX_REG_13__SCAN_IN), .ZN(n20619) );
  NAND2_X1 U22642 ( .A1(n20616), .A2(n20686), .ZN(n20656) );
  AOI22_X1 U22643 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n20790), .B1(n20789), .B2(
        n20617), .ZN(n20618) );
  OAI221_X1 U22644 ( .B1(n20620), .B2(P3_EAX_REG_13__SCAN_IN), .C1(n20619), 
        .C2(n20776), .A(n20618), .ZN(P3_U2722) );
  INV_X1 U22645 ( .A(n20620), .ZN(n20764) );
  AOI21_X1 U22646 ( .B1(P3_EAX_REG_12__SCAN_IN), .B2(n20785), .A(n20621), .ZN(
        n20623) );
  OAI222_X1 U22647 ( .A1(n20656), .A2(n20624), .B1(n20764), .B2(n20623), .C1(
        n20781), .C2(n20622), .ZN(P3_U2723) );
  NAND2_X1 U22648 ( .A1(n20785), .A2(n20628), .ZN(n20631) );
  AOI22_X1 U22649 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n20790), .B1(n20789), .B2(
        n20625), .ZN(n20626) );
  OAI221_X1 U22650 ( .B1(P3_EAX_REG_11__SCAN_IN), .B2(n20628), .C1(n20627), 
        .C2(n20631), .A(n20626), .ZN(P3_U2724) );
  NOR2_X1 U22651 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n20636), .ZN(n20630) );
  OAI222_X1 U22652 ( .A1(n20656), .A2(n20718), .B1(n20631), .B2(n20630), .C1(
        n20781), .C2(n20629), .ZN(P3_U2725) );
  INV_X1 U22653 ( .A(n20632), .ZN(n20633) );
  AOI21_X1 U22654 ( .B1(P3_EAX_REG_9__SCAN_IN), .B2(n20785), .A(n20633), .ZN(
        n20635) );
  OAI222_X1 U22655 ( .A1(n20656), .A2(n20637), .B1(n20636), .B2(n20635), .C1(
        n20781), .C2(n20634), .ZN(P3_U2726) );
  NAND2_X1 U22656 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n20790), .ZN(n20640) );
  OAI211_X1 U22657 ( .C1(n20638), .C2(P3_EAX_REG_7__SCAN_IN), .A(n20785), .B(
        n20778), .ZN(n20639) );
  OAI211_X1 U22658 ( .C1(n21106), .C2(n20781), .A(n20640), .B(n20639), .ZN(
        P3_U2728) );
  NOR2_X1 U22659 ( .A1(n20711), .A2(n20641), .ZN(n20648) );
  INV_X1 U22660 ( .A(n20648), .ZN(n20645) );
  NAND2_X1 U22661 ( .A1(n20645), .A2(P3_EAX_REG_6__SCAN_IN), .ZN(n20644) );
  AOI22_X1 U22662 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n20790), .B1(n20789), .B2(
        n20642), .ZN(n20643) );
  OAI221_X1 U22663 ( .B1(n20645), .B2(P3_EAX_REG_6__SCAN_IN), .C1(n20644), 
        .C2(n20776), .A(n20643), .ZN(P3_U2729) );
  NAND3_X1 U22664 ( .A1(n20687), .A2(n20662), .A3(P3_EAX_REG_3__SCAN_IN), .ZN(
        n20658) );
  NOR2_X1 U22665 ( .A1(n20650), .A2(n20658), .ZN(n20655) );
  AOI21_X1 U22666 ( .B1(P3_EAX_REG_5__SCAN_IN), .B2(n20785), .A(n20655), .ZN(
        n20647) );
  OAI222_X1 U22667 ( .A1(n20649), .A2(n20656), .B1(n20648), .B2(n20647), .C1(
        n20781), .C2(n20646), .ZN(P3_U2730) );
  OAI21_X1 U22668 ( .B1(n20650), .B2(n20776), .A(n20658), .ZN(n20651) );
  INV_X1 U22669 ( .A(n20651), .ZN(n20654) );
  INV_X1 U22670 ( .A(n20652), .ZN(n20653) );
  OAI222_X1 U22671 ( .A1(n20657), .A2(n20656), .B1(n20655), .B2(n20654), .C1(
        n20781), .C2(n20653), .ZN(P3_U2731) );
  NAND2_X1 U22672 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n20790), .ZN(n20660) );
  OAI211_X1 U22673 ( .C1(n20662), .C2(P3_EAX_REG_3__SCAN_IN), .A(n20785), .B(
        n20658), .ZN(n20659) );
  OAI211_X1 U22674 ( .C1(n20661), .C2(n20781), .A(n20660), .B(n20659), .ZN(
        P3_U2732) );
  AOI21_X1 U22675 ( .B1(n20663), .B2(n20784), .A(n20662), .ZN(n20664) );
  AOI22_X1 U22676 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n20790), .B1(n20664), .B2(
        n20785), .ZN(n20665) );
  OAI21_X1 U22677 ( .B1(n20666), .B2(n20781), .A(n20665), .ZN(P3_U2733) );
  NOR4_X1 U22678 ( .A1(n20670), .A2(n20669), .A3(n20668), .A4(n20667), .ZN(
        n20671) );
  NAND4_X2 U22679 ( .A1(n20775), .A2(P3_EAX_REG_14__SCAN_IN), .A3(
        P3_EAX_REG_11__SCAN_IN), .A4(n20671), .ZN(n20771) );
  NOR2_X2 U22680 ( .A1(n20771), .A2(n20770), .ZN(n20769) );
  NAND2_X1 U22681 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n20703), .ZN(n20699) );
  NAND2_X1 U22682 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n20693), .ZN(n20678) );
  NAND2_X1 U22683 ( .A1(n20785), .A2(n20678), .ZN(n20688) );
  NOR2_X2 U22684 ( .A1(n20673), .A2(n20785), .ZN(n20759) );
  NOR2_X2 U22685 ( .A1(n20674), .A2(n20785), .ZN(n20758) );
  INV_X1 U22686 ( .A(n20758), .ZN(n20752) );
  OAI22_X1 U22687 ( .A1(n20675), .A2(n20781), .B1(n16232), .B2(n20752), .ZN(
        n20676) );
  AOI21_X1 U22688 ( .B1(BUF2_REG_5__SCAN_IN), .B2(n20759), .A(n20676), .ZN(
        n20677) );
  OAI221_X1 U22689 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n20678), .C1(n20683), 
        .C2(n20688), .A(n20677), .ZN(P3_U2714) );
  AOI22_X1 U22690 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n20759), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n20758), .ZN(n20680) );
  OAI211_X1 U22691 ( .C1(n20693), .C2(P3_EAX_REG_20__SCAN_IN), .A(n20785), .B(
        n20678), .ZN(n20679) );
  OAI211_X1 U22692 ( .C1(n20681), .C2(n20781), .A(n20680), .B(n20679), .ZN(
        P3_U2715) );
  NOR2_X1 U22693 ( .A1(n20683), .A2(n20682), .ZN(n20684) );
  NAND4_X1 U22694 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(P3_EAX_REG_17__SCAN_IN), 
        .A3(P3_EAX_REG_18__SCAN_IN), .A4(n20684), .ZN(n20710) );
  NOR2_X1 U22695 ( .A1(n20711), .A2(n20760), .ZN(n20705) );
  NAND2_X1 U22696 ( .A1(n20705), .A2(n20709), .ZN(n20692) );
  AOI22_X1 U22697 ( .A1(BUF2_REG_22__SCAN_IN), .A2(n20758), .B1(n20789), .B2(
        n20685), .ZN(n20691) );
  NAND2_X1 U22698 ( .A1(n20687), .A2(n20686), .ZN(n20792) );
  OAI21_X1 U22699 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n20792), .A(n20688), .ZN(
        n20689) );
  AOI22_X1 U22700 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n20759), .B1(
        P3_EAX_REG_22__SCAN_IN), .B2(n20689), .ZN(n20690) );
  OAI211_X1 U22701 ( .C1(n20710), .C2(n20692), .A(n20691), .B(n20690), .ZN(
        P3_U2713) );
  AOI22_X1 U22702 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n20759), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n20758), .ZN(n20697) );
  AOI211_X1 U22703 ( .C1(n20694), .C2(n20699), .A(n20693), .B(n20776), .ZN(
        n20695) );
  INV_X1 U22704 ( .A(n20695), .ZN(n20696) );
  OAI211_X1 U22705 ( .C1(n20698), .C2(n20781), .A(n20697), .B(n20696), .ZN(
        P3_U2716) );
  AOI22_X1 U22706 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n20759), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n20758), .ZN(n20701) );
  OAI211_X1 U22707 ( .C1(n20703), .C2(P3_EAX_REG_18__SCAN_IN), .A(n20785), .B(
        n20699), .ZN(n20700) );
  OAI211_X1 U22708 ( .C1(n20702), .C2(n20781), .A(n20701), .B(n20700), .ZN(
        P3_U2717) );
  AOI22_X1 U22709 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n20759), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n20758), .ZN(n20707) );
  INV_X1 U22710 ( .A(n20703), .ZN(n20704) );
  OAI211_X1 U22711 ( .C1(n20705), .C2(P3_EAX_REG_17__SCAN_IN), .A(n20785), .B(
        n20704), .ZN(n20706) );
  OAI211_X1 U22712 ( .C1(n20708), .C2(n20781), .A(n20707), .B(n20706), .ZN(
        P3_U2718) );
  AOI22_X1 U22713 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n20759), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n20758), .ZN(n20714) );
  NOR3_X2 U22714 ( .A1(n20760), .A2(n20710), .A3(n20709), .ZN(n20754) );
  NAND2_X1 U22715 ( .A1(n20754), .A2(P3_EAX_REG_23__SCAN_IN), .ZN(n20753) );
  OAI211_X1 U22716 ( .C1(n20712), .C2(P3_EAX_REG_25__SCAN_IN), .A(n20785), .B(
        n20719), .ZN(n20713) );
  OAI211_X1 U22717 ( .C1(n20715), .C2(n20781), .A(n20714), .B(n20713), .ZN(
        P3_U2710) );
  INV_X1 U22718 ( .A(n20759), .ZN(n20717) );
  OAI22_X1 U22719 ( .A1(n20718), .A2(n20717), .B1(n20781), .B2(n20716), .ZN(
        n20722) );
  AOI211_X1 U22720 ( .C1(n20720), .C2(n20719), .A(n20743), .B(n20776), .ZN(
        n20721) );
  AOI211_X1 U22721 ( .C1(n20758), .C2(BUF2_REG_26__SCAN_IN), .A(n20722), .B(
        n20721), .ZN(n20723) );
  INV_X1 U22722 ( .A(n20723), .ZN(P3_U2709) );
  NAND2_X1 U22723 ( .A1(n20743), .A2(P3_EAX_REG_27__SCAN_IN), .ZN(n20742) );
  NOR2_X2 U22724 ( .A1(n20742), .A2(n20738), .ZN(n20737) );
  NAND2_X1 U22725 ( .A1(n20737), .A2(P3_EAX_REG_29__SCAN_IN), .ZN(n20731) );
  NAND2_X1 U22726 ( .A1(n20727), .A2(P3_EAX_REG_30__SCAN_IN), .ZN(n20726) );
  OAI22_X1 U22727 ( .A1(n20776), .A2(n20727), .B1(P3_EAX_REG_30__SCAN_IN), 
        .B2(n20792), .ZN(n20724) );
  AOI22_X1 U22728 ( .A1(BUF2_REG_31__SCAN_IN), .A2(n20758), .B1(
        P3_EAX_REG_31__SCAN_IN), .B2(n20724), .ZN(n20725) );
  OAI21_X1 U22729 ( .B1(P3_EAX_REG_31__SCAN_IN), .B2(n20726), .A(n20725), .ZN(
        P3_U2704) );
  AOI22_X1 U22730 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n20759), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n20758), .ZN(n20729) );
  OAI211_X1 U22731 ( .C1(n20727), .C2(P3_EAX_REG_30__SCAN_IN), .A(n20785), .B(
        n20726), .ZN(n20728) );
  OAI211_X1 U22732 ( .C1(n20730), .C2(n20781), .A(n20729), .B(n20728), .ZN(
        P3_U2705) );
  AOI22_X1 U22733 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n20759), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n20758), .ZN(n20733) );
  OAI211_X1 U22734 ( .C1(n20737), .C2(P3_EAX_REG_29__SCAN_IN), .A(n20785), .B(
        n20731), .ZN(n20732) );
  OAI211_X1 U22735 ( .C1(n20734), .C2(n20781), .A(n20733), .B(n20732), .ZN(
        P3_U2706) );
  AOI22_X1 U22736 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n20759), .B1(n20789), .B2(
        n20735), .ZN(n20736) );
  INV_X1 U22737 ( .A(n20736), .ZN(n20740) );
  AOI211_X1 U22738 ( .C1(n20738), .C2(n20742), .A(n20737), .B(n20776), .ZN(
        n20739) );
  AOI211_X1 U22739 ( .C1(n20758), .C2(BUF2_REG_28__SCAN_IN), .A(n20740), .B(
        n20739), .ZN(n20741) );
  INV_X1 U22740 ( .A(n20741), .ZN(P3_U2707) );
  AOI22_X1 U22741 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n20759), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n20758), .ZN(n20745) );
  OAI211_X1 U22742 ( .C1(n20743), .C2(P3_EAX_REG_27__SCAN_IN), .A(n20785), .B(
        n20742), .ZN(n20744) );
  OAI211_X1 U22743 ( .C1(n20746), .C2(n20781), .A(n20745), .B(n20744), .ZN(
        P3_U2708) );
  AOI22_X1 U22744 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n20759), .B1(n20789), .B2(
        n20747), .ZN(n20751) );
  OAI211_X1 U22745 ( .C1(n20749), .C2(P3_EAX_REG_24__SCAN_IN), .A(n20785), .B(
        n20748), .ZN(n20750) );
  OAI211_X1 U22746 ( .C1(n20752), .C2(n16212), .A(n20751), .B(n20750), .ZN(
        P3_U2711) );
  AOI22_X1 U22747 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n20759), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n20758), .ZN(n20756) );
  OAI211_X1 U22748 ( .C1(n20754), .C2(P3_EAX_REG_23__SCAN_IN), .A(n20785), .B(
        n20753), .ZN(n20755) );
  OAI211_X1 U22749 ( .C1(n20757), .C2(n20781), .A(n20756), .B(n20755), .ZN(
        P3_U2712) );
  AOI22_X1 U22750 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n20759), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n20758), .ZN(n20762) );
  OAI211_X1 U22751 ( .C1(n20769), .C2(P3_EAX_REG_16__SCAN_IN), .A(n20785), .B(
        n20760), .ZN(n20761) );
  OAI211_X1 U22752 ( .C1(n20763), .C2(n20781), .A(n20762), .B(n20761), .ZN(
        P3_U2719) );
  NAND2_X1 U22753 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(n20764), .ZN(n20768) );
  AOI22_X1 U22754 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n20790), .B1(n20789), .B2(
        n20765), .ZN(n20767) );
  NAND3_X1 U22755 ( .A1(P3_EAX_REG_14__SCAN_IN), .A2(n20785), .A3(n20771), 
        .ZN(n20766) );
  OAI211_X1 U22756 ( .C1(P3_EAX_REG_14__SCAN_IN), .C2(n20768), .A(n20767), .B(
        n20766), .ZN(P3_U2721) );
  AOI211_X1 U22757 ( .C1(n20771), .C2(n20770), .A(n20776), .B(n20769), .ZN(
        n20772) );
  AOI21_X1 U22758 ( .B1(n20790), .B2(BUF2_REG_15__SCAN_IN), .A(n20772), .ZN(
        n20773) );
  OAI21_X1 U22759 ( .B1(n20774), .B2(n20781), .A(n20773), .ZN(P3_U2720) );
  AOI211_X1 U22760 ( .C1(n20778), .C2(n20777), .A(n20776), .B(n20775), .ZN(
        n20779) );
  AOI21_X1 U22761 ( .B1(n20790), .B2(BUF2_REG_8__SCAN_IN), .A(n20779), .ZN(
        n20780) );
  OAI21_X1 U22762 ( .B1(n20782), .B2(n20781), .A(n20780), .ZN(P3_U2727) );
  AOI22_X1 U22763 ( .A1(n20790), .A2(BUF2_REG_1__SCAN_IN), .B1(n20789), .B2(
        n20783), .ZN(n20787) );
  OAI211_X1 U22764 ( .C1(n20794), .C2(P3_EAX_REG_1__SCAN_IN), .A(n20785), .B(
        n20784), .ZN(n20786) );
  NAND2_X1 U22765 ( .A1(n20787), .A2(n20786), .ZN(P3_U2734) );
  AOI22_X1 U22766 ( .A1(n20790), .A2(BUF2_REG_0__SCAN_IN), .B1(n20789), .B2(
        n20788), .ZN(n20791) );
  OAI221_X1 U22767 ( .B1(n20794), .B2(n20793), .C1(n20794), .C2(n20792), .A(
        n20791), .ZN(P3_U2735) );
  INV_X1 U22768 ( .A(n20795), .ZN(n20796) );
  NAND2_X1 U22769 ( .A1(n21006), .A2(n20796), .ZN(n20799) );
  AOI22_X1 U22770 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n21237), .B1(
        n20799), .B2(n20829), .ZN(n21264) );
  INV_X1 U22771 ( .A(n21264), .ZN(n21261) );
  AOI222_X1 U22772 ( .A1(n20881), .A2(P3_STATE2_REG_1__SCAN_IN), .B1(n21261), 
        .B2(n20839), .C1(n20829), .C2(n21300), .ZN(n20797) );
  AOI22_X1 U22773 ( .A1(n20843), .A2(n20829), .B1(n20797), .B2(n20841), .ZN(
        P3_U3290) );
  NOR2_X1 U22774 ( .A1(n20798), .A2(n20881), .ZN(n20818) );
  INV_X1 U22775 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n21102) );
  AOI22_X1 U22776 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n21102), .B1(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n20882), .ZN(n20815) );
  OAI21_X1 U22777 ( .B1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n21237), .A(
        n21229), .ZN(n20823) );
  INV_X1 U22778 ( .A(n20823), .ZN(n20805) );
  AOI22_X1 U22779 ( .A1(n20800), .A2(n20799), .B1(n20805), .B2(n20825), .ZN(
        n21266) );
  NAND2_X1 U22780 ( .A1(n21300), .A2(n20810), .ZN(n20821) );
  OAI22_X1 U22781 ( .A1(n21266), .A2(n20802), .B1(n20801), .B2(n20821), .ZN(
        n20803) );
  AOI21_X1 U22782 ( .B1(n20818), .B2(n20815), .A(n20803), .ZN(n20804) );
  AOI22_X1 U22783 ( .A1(n20843), .A2(n20825), .B1(n20804), .B2(n20841), .ZN(
        P3_U3289) );
  OAI221_X1 U22784 ( .B1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .C1(n20825), .C2(n20822), .A(
        n20805), .ZN(n20813) );
  AOI22_X1 U22785 ( .A1(n20809), .A2(n20808), .B1(n20807), .B2(n20806), .ZN(
        n20833) );
  INV_X1 U22786 ( .A(n20833), .ZN(n20811) );
  OAI211_X1 U22787 ( .C1(n20828), .C2(n20811), .A(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n20810), .ZN(n20812) );
  OAI211_X1 U22788 ( .C1(n20814), .C2(n11276), .A(n20813), .B(n20812), .ZN(
        n21270) );
  INV_X1 U22789 ( .A(n20815), .ZN(n20819) );
  INV_X1 U22790 ( .A(n20816), .ZN(n20817) );
  AOI222_X1 U22791 ( .A1(n21270), .A2(n20839), .B1(n20819), .B2(n20818), .C1(
        n20817), .C2(n21300), .ZN(n20820) );
  OAI222_X1 U22792 ( .A1(n20822), .A2(n20821), .B1(n20822), .B2(n20841), .C1(
        n20843), .C2(n20820), .ZN(P3_U3288) );
  AOI21_X1 U22793 ( .B1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(n21260), .ZN(n20837) );
  NOR3_X1 U22794 ( .A1(n20825), .A2(n20824), .A3(n20823), .ZN(n20835) );
  OAI221_X1 U22795 ( .B1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n20827), 
        .C1(n21260), .C2(n20826), .A(n21256), .ZN(n20831) );
  NAND3_X1 U22796 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n20829), .A3(
        n20828), .ZN(n20830) );
  OAI211_X1 U22797 ( .C1(n20833), .C2(n20832), .A(n20831), .B(n20830), .ZN(
        n20834) );
  AOI211_X1 U22798 ( .C1(n20837), .C2(n20836), .A(n20835), .B(n20834), .ZN(
        n21259) );
  INV_X1 U22799 ( .A(n21259), .ZN(n20838) );
  AOI22_X1 U22800 ( .A1(n21300), .A2(n20840), .B1(n20839), .B2(n20838), .ZN(
        n20842) );
  AOI22_X1 U22801 ( .A1(n20843), .A2(n21260), .B1(n20842), .B2(n20841), .ZN(
        P3_U3285) );
  NAND2_X1 U22802 ( .A1(n21104), .A2(n21106), .ZN(n21149) );
  OAI22_X1 U22803 ( .A1(n21149), .A2(n21176), .B1(n21147), .B2(n20952), .ZN(
        n20947) );
  INV_X1 U22804 ( .A(n20947), .ZN(n20852) );
  INV_X1 U22805 ( .A(n20849), .ZN(n20851) );
  INV_X1 U22806 ( .A(n21006), .ZN(n21231) );
  NOR2_X1 U22807 ( .A1(n20845), .A2(n20844), .ZN(n20924) );
  NAND3_X1 U22808 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n20924), .A3(
        n20897), .ZN(n21236) );
  NOR2_X1 U22809 ( .A1(n21232), .A2(n21236), .ZN(n21218) );
  NAND2_X1 U22810 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n21218), .ZN(
        n21230) );
  NOR2_X1 U22811 ( .A1(n20851), .A2(n21230), .ZN(n20855) );
  NAND4_X1 U22812 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A3(n20924), .A4(n20846), .ZN(
        n20960) );
  NOR2_X1 U22813 ( .A1(n20847), .A2(n20960), .ZN(n21169) );
  AND2_X1 U22814 ( .A1(n20848), .A2(n21169), .ZN(n21015) );
  NAND2_X1 U22815 ( .A1(n20849), .A2(n21218), .ZN(n21005) );
  INV_X1 U22816 ( .A(n21005), .ZN(n20850) );
  AOI222_X1 U22817 ( .A1(n21231), .A2(n20855), .B1(n21015), .B2(n21256), .C1(
        n21237), .C2(n20850), .ZN(n21060) );
  OAI21_X1 U22818 ( .B1(n20852), .B2(n20851), .A(n21060), .ZN(n21050) );
  NAND2_X1 U22819 ( .A1(n21117), .A2(n21050), .ZN(n21166) );
  AOI21_X1 U22820 ( .B1(n21203), .B2(n20854), .A(n20853), .ZN(n20864) );
  OAI21_X1 U22821 ( .B1(n21006), .B2(n20855), .A(n21117), .ZN(n21146) );
  INV_X1 U22822 ( .A(n20856), .ZN(n20860) );
  OAI21_X1 U22823 ( .B1(n21005), .B2(n21158), .A(n21237), .ZN(n20857) );
  OAI21_X1 U22824 ( .B1(n21015), .B2(n11276), .A(n20857), .ZN(n21145) );
  OAI22_X1 U22825 ( .A1(n21222), .A2(n20861), .B1(n20858), .B2(n21147), .ZN(
        n20859) );
  AOI211_X1 U22826 ( .C1(n21177), .C2(n20860), .A(n21145), .B(n20859), .ZN(
        n21008) );
  OAI21_X1 U22827 ( .B1(n21006), .B2(n20861), .A(n21008), .ZN(n20862) );
  OAI211_X1 U22828 ( .C1(n21146), .C2(n20862), .A(
        P3_INSTADDRPOINTER_REG_21__SCAN_IN), .B(n21223), .ZN(n20863) );
  OAI211_X1 U22829 ( .C1(n21166), .C2(n20865), .A(n20864), .B(n20863), .ZN(
        P3_U2841) );
  AND2_X1 U22830 ( .A1(n21238), .A2(P3_REIP_REG_0__SCAN_IN), .ZN(n20867) );
  NOR2_X1 U22831 ( .A1(n21256), .A2(n21231), .ZN(n21161) );
  AOI221_X1 U22832 ( .B1(n21161), .B2(n20881), .C1(n21219), .C2(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(n21234), .ZN(n20866) );
  AOI211_X1 U22833 ( .C1(n21133), .C2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n20867), .B(n20866), .ZN(n20868) );
  OAI221_X1 U22834 ( .B1(n20870), .B2(n21048), .C1(n20869), .C2(n20929), .A(
        n20868), .ZN(P3_U2862) );
  NOR2_X1 U22835 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n21237), .ZN(
        n20871) );
  NOR2_X1 U22836 ( .A1(n21201), .A2(n20871), .ZN(n20873) );
  NOR2_X1 U22837 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n21161), .ZN(
        n20872) );
  MUX2_X1 U22838 ( .A(n20873), .B(n20872), .S(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .Z(n20877) );
  OAI22_X1 U22839 ( .A1(n20875), .A2(n21048), .B1(n20929), .B2(n20874), .ZN(
        n20876) );
  AOI21_X1 U22840 ( .B1(n21117), .B2(n20877), .A(n20876), .ZN(n20879) );
  NAND2_X1 U22841 ( .A1(n21238), .A2(P3_REIP_REG_1__SCAN_IN), .ZN(n20878) );
  OAI211_X1 U22842 ( .C1(n21220), .C2(n20882), .A(n20879), .B(n20878), .ZN(
        P3_U2861) );
  OR2_X1 U22843 ( .A1(n20882), .A2(n20880), .ZN(n20887) );
  NOR2_X1 U22844 ( .A1(n20882), .A2(n20881), .ZN(n20884) );
  INV_X1 U22845 ( .A(n21173), .ZN(n20896) );
  AOI21_X1 U22846 ( .B1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n20896), .A(
        n21184), .ZN(n20883) );
  AOI21_X1 U22847 ( .B1(n20884), .B2(n21256), .A(n20883), .ZN(n20886) );
  NAND2_X1 U22848 ( .A1(n21256), .A2(n20885), .ZN(n20895) );
  OAI221_X1 U22849 ( .B1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n20887), .C1(
        n20894), .C2(n20886), .A(n20895), .ZN(n20891) );
  OAI22_X1 U22850 ( .A1(n21251), .A2(n20889), .B1(n21147), .B2(n20888), .ZN(
        n20890) );
  OAI21_X1 U22851 ( .B1(n20891), .B2(n20890), .A(n21117), .ZN(n20892) );
  OAI211_X1 U22852 ( .C1(n21220), .C2(n20894), .A(n20893), .B(n20892), .ZN(
        P3_U2860) );
  OAI211_X1 U22853 ( .C1(n21184), .C2(n20897), .A(n20896), .B(n20895), .ZN(
        n20898) );
  OAI21_X1 U22854 ( .B1(n20915), .B2(n20898), .A(n21117), .ZN(n20905) );
  OAI21_X1 U22855 ( .B1(n21220), .B2(n20915), .A(n20905), .ZN(n20902) );
  OAI22_X1 U22856 ( .A1(n20929), .A2(n20900), .B1(n21048), .B2(n20899), .ZN(
        n20901) );
  AOI221_X1 U22857 ( .B1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n20902), .C1(
        n20923), .C2(n20902), .A(n20901), .ZN(n20904) );
  NAND2_X1 U22858 ( .A1(n20904), .A2(n20903), .ZN(P3_U2859) );
  OAI21_X1 U22859 ( .B1(n21201), .B2(n20905), .A(n21220), .ZN(n20910) );
  NOR3_X1 U22860 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n20915), .A3(
        n20913), .ZN(n20909) );
  OAI22_X1 U22861 ( .A1(n21223), .A2(n20907), .B1(n21048), .B2(n20906), .ZN(
        n20908) );
  AOI211_X1 U22862 ( .C1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .C2(n20910), .A(
        n20909), .B(n20908), .ZN(n20911) );
  OAI21_X1 U22863 ( .B1(n20929), .B2(n20912), .A(n20911), .ZN(P3_U2858) );
  NOR4_X1 U22864 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n20915), .A3(
        n20914), .A4(n20913), .ZN(n20919) );
  OAI21_X1 U22865 ( .B1(n20917), .B2(n20929), .A(n20916), .ZN(n20918) );
  AOI211_X1 U22866 ( .C1(n20920), .C2(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A(
        n20919), .B(n20918), .ZN(n20921) );
  OAI21_X1 U22867 ( .B1(n21048), .B2(n20922), .A(n20921), .ZN(P3_U2857) );
  NAND2_X1 U22868 ( .A1(n20924), .A2(n20923), .ZN(n20945) );
  OAI211_X1 U22869 ( .C1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .C2(n11276), .A(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .B(n20925), .ZN(n20926) );
  AOI21_X1 U22870 ( .B1(n21236), .B2(n21229), .A(n20926), .ZN(n20934) );
  AOI211_X1 U22871 ( .C1(n20935), .C2(n20945), .A(n20934), .B(n21234), .ZN(
        n20931) );
  OAI22_X1 U22872 ( .A1(n20929), .A2(n20928), .B1(n21048), .B2(n20927), .ZN(
        n20930) );
  NOR2_X1 U22873 ( .A1(n20931), .A2(n20930), .ZN(n20933) );
  NAND2_X1 U22874 ( .A1(n21238), .A2(P3_REIP_REG_7__SCAN_IN), .ZN(n20932) );
  OAI211_X1 U22875 ( .C1(n21220), .C2(n20935), .A(n20933), .B(n20932), .ZN(
        P3_U2855) );
  NOR3_X1 U22876 ( .A1(n21201), .A2(n20934), .A3(n21232), .ZN(n20937) );
  NOR3_X1 U22877 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n20935), .A3(
        n20945), .ZN(n20936) );
  AOI211_X1 U22878 ( .C1(n21177), .C2(n20940), .A(n20937), .B(n20936), .ZN(
        n20944) );
  NOR2_X1 U22879 ( .A1(n21223), .A2(n20938), .ZN(n20942) );
  OAI22_X1 U22880 ( .A1(n21246), .A2(n20940), .B1(n21048), .B2(n20939), .ZN(
        n20941) );
  AOI211_X1 U22881 ( .C1(n21133), .C2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A(
        n20942), .B(n20941), .ZN(n20943) );
  OAI21_X1 U22882 ( .B1(n20944), .B2(n21234), .A(n20943), .ZN(P3_U2854) );
  NOR2_X1 U22883 ( .A1(n20946), .A2(n20945), .ZN(n20993) );
  NOR2_X1 U22884 ( .A1(n20993), .A2(n20947), .ZN(n20968) );
  AOI22_X1 U22885 ( .A1(n21238), .A2(P3_REIP_REG_11__SCAN_IN), .B1(n21242), 
        .B2(n20948), .ZN(n20958) );
  AOI21_X1 U22886 ( .B1(n20954), .B2(n21218), .A(n21219), .ZN(n20963) );
  NOR2_X1 U22887 ( .A1(n21177), .A2(n21254), .ZN(n21179) );
  NAND2_X1 U22888 ( .A1(n21256), .A2(n20960), .ZN(n20949) );
  OAI21_X1 U22889 ( .B1(n20950), .B2(n21149), .A(n20949), .ZN(n20951) );
  AOI21_X1 U22890 ( .B1(n21254), .B2(n20952), .A(n20951), .ZN(n21240) );
  OAI21_X1 U22891 ( .B1(n21241), .B2(n21230), .A(n21231), .ZN(n20953) );
  OAI211_X1 U22892 ( .C1(n20954), .C2(n21179), .A(n21240), .B(n20953), .ZN(
        n21225) );
  AOI211_X1 U22893 ( .C1(n21256), .C2(n20967), .A(n21234), .B(n21225), .ZN(
        n20955) );
  OAI21_X1 U22894 ( .B1(n21006), .B2(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n20955), .ZN(n20956) );
  OAI211_X1 U22895 ( .C1(n20963), .C2(n20956), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n21223), .ZN(n20957) );
  OAI211_X1 U22896 ( .C1(n20959), .C2(n21246), .A(n20958), .B(n20957), .ZN(
        P3_U2851) );
  OAI21_X1 U22897 ( .B1(n20960), .B2(n20967), .A(n21256), .ZN(n20979) );
  OAI21_X1 U22898 ( .B1(n20961), .B2(n21147), .A(n20979), .ZN(n20962) );
  AOI211_X1 U22899 ( .C1(n21177), .C2(n20964), .A(n20963), .B(n20962), .ZN(
        n21211) );
  AOI211_X1 U22900 ( .C1(n21237), .C2(n21209), .A(n21231), .B(n11379), .ZN(
        n20966) );
  NOR2_X1 U22901 ( .A1(n20965), .A2(n21230), .ZN(n20976) );
  AOI211_X1 U22902 ( .C1(n21211), .C2(n20966), .A(n20976), .B(n21234), .ZN(
        n20970) );
  OAI21_X1 U22903 ( .B1(n20968), .B2(n20967), .A(n11379), .ZN(n20969) );
  AOI22_X1 U22904 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n21133), .B1(
        n20970), .B2(n20969), .ZN(n20972) );
  OAI211_X1 U22905 ( .C1(n20973), .C2(n21246), .A(n20972), .B(n20971), .ZN(
        P3_U2850) );
  AOI22_X1 U22906 ( .A1(n21238), .A2(P3_REIP_REG_14__SCAN_IN), .B1(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n21133), .ZN(n20988) );
  NAND3_X1 U22907 ( .A1(n20975), .A2(n20993), .A3(n20974), .ZN(n20982) );
  OAI22_X1 U22908 ( .A1(n21006), .A2(n20976), .B1(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n11276), .ZN(n21213) );
  INV_X1 U22909 ( .A(n20977), .ZN(n20992) );
  NAND2_X1 U22910 ( .A1(n20992), .A2(n21218), .ZN(n21171) );
  NAND2_X1 U22911 ( .A1(n21237), .A2(n21171), .ZN(n20978) );
  OAI211_X1 U22912 ( .C1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .C2(n21161), .A(
        n20979), .B(n20978), .ZN(n20980) );
  OAI21_X1 U22913 ( .B1(n21213), .B2(n20980), .A(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n20981) );
  OAI211_X1 U22914 ( .C1(n21149), .C2(n20983), .A(n20982), .B(n20981), .ZN(
        n20986) );
  INV_X1 U22915 ( .A(n21048), .ZN(n20985) );
  AOI22_X1 U22916 ( .A1(n21117), .A2(n20986), .B1(n20985), .B2(n20984), .ZN(
        n20987) );
  OAI211_X1 U22917 ( .C1(n20989), .C2(n21246), .A(n20988), .B(n20987), .ZN(
        P3_U2848) );
  NAND2_X1 U22918 ( .A1(n21177), .A2(n20990), .ZN(n20997) );
  AOI221_X1 U22919 ( .B1(n21231), .B2(n21171), .C1(n21237), .C2(n21171), .A(
        n21173), .ZN(n20991) );
  OAI211_X1 U22920 ( .C1(n21169), .C2(n11276), .A(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B(n20991), .ZN(n20996) );
  NAND3_X1 U22921 ( .A1(n20993), .A2(n20992), .A3(n20996), .ZN(n20995) );
  AOI221_X1 U22922 ( .B1(n20997), .B2(n20995), .C1(n20994), .C2(n20995), .A(
        n21234), .ZN(n21000) );
  INV_X1 U22923 ( .A(n20996), .ZN(n21199) );
  INV_X1 U22924 ( .A(n20997), .ZN(n20998) );
  AOI211_X1 U22925 ( .C1(n21254), .C2(n21174), .A(n20998), .B(n21234), .ZN(
        n21200) );
  AOI211_X1 U22926 ( .C1(n21199), .C2(n21200), .A(n21238), .B(n21172), .ZN(
        n20999) );
  AOI211_X1 U22927 ( .C1(n21203), .C2(n21001), .A(n21000), .B(n20999), .ZN(
        n21003) );
  OAI211_X1 U22928 ( .C1(n21004), .C2(n21048), .A(n21003), .B(n21002), .ZN(
        P3_U2847) );
  AOI22_X1 U22929 ( .A1(n21238), .A2(P3_REIP_REG_22__SCAN_IN), .B1(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n21133), .ZN(n21013) );
  AND2_X1 U22930 ( .A1(n21050), .A2(n21031), .ZN(n21011) );
  NAND2_X1 U22931 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n21031), .ZN(
        n21059) );
  NOR2_X1 U22932 ( .A1(n21005), .A2(n21059), .ZN(n21063) );
  AOI21_X1 U22933 ( .B1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n21063), .A(
        n21006), .ZN(n21007) );
  INV_X1 U22934 ( .A(n21007), .ZN(n21016) );
  OAI211_X1 U22935 ( .C1(n21222), .C2(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n21008), .B(n21016), .ZN(n21009) );
  OAI221_X1 U22936 ( .B1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n21011), 
        .C1(n21010), .C2(n21009), .A(n21117), .ZN(n21012) );
  OAI211_X1 U22937 ( .C1(n21014), .C2(n21246), .A(n21013), .B(n21012), .ZN(
        P3_U2840) );
  NAND2_X1 U22938 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n21041) );
  NOR4_X1 U22939 ( .A1(n21060), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A3(
        n21059), .A4(n21041), .ZN(n21019) );
  INV_X1 U22940 ( .A(n21059), .ZN(n21051) );
  AOI21_X1 U22941 ( .B1(n21015), .B2(n21051), .A(n11276), .ZN(n21129) );
  OAI21_X1 U22942 ( .B1(n21219), .B2(n21063), .A(n21016), .ZN(n21124) );
  AOI211_X1 U22943 ( .C1(n21141), .C2(n21041), .A(n21129), .B(n21124), .ZN(
        n21026) );
  OAI22_X1 U22944 ( .A1(n21026), .A2(n21033), .B1(n21147), .B2(n21017), .ZN(
        n21018) );
  AOI211_X1 U22945 ( .C1(n21020), .C2(n21177), .A(n21019), .B(n21018), .ZN(
        n21024) );
  AOI22_X1 U22946 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n21133), .B1(
        n21203), .B2(n21021), .ZN(n21023) );
  NAND2_X1 U22947 ( .A1(n21238), .A2(P3_REIP_REG_25__SCAN_IN), .ZN(n21022) );
  OAI211_X1 U22948 ( .C1(n21024), .C2(n21234), .A(n21023), .B(n21022), .ZN(
        P3_U2837) );
  INV_X1 U22949 ( .A(n21025), .ZN(n21038) );
  OAI211_X1 U22950 ( .C1(n21201), .C2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B(n21026), .ZN(n21027) );
  AOI21_X1 U22951 ( .B1(n21177), .B2(n21028), .A(n21027), .ZN(n21029) );
  OAI22_X1 U22952 ( .A1(n21049), .A2(n21048), .B1(n21029), .B2(n21234), .ZN(
        n21035) );
  NAND3_X1 U22953 ( .A1(n21031), .A2(n21030), .A3(n21050), .ZN(n21137) );
  NOR3_X1 U22954 ( .A1(n21033), .A2(n21032), .A3(n21137), .ZN(n21034) );
  AOI222_X1 U22955 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n21035), 
        .B1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n21133), .C1(n21035), 
        .C2(n21034), .ZN(n21037) );
  OAI211_X1 U22956 ( .C1(n21038), .C2(n21246), .A(n21037), .B(n21036), .ZN(
        P3_U2836) );
  INV_X1 U22957 ( .A(n21039), .ZN(n21056) );
  INV_X1 U22958 ( .A(n21040), .ZN(n21042) );
  NOR2_X1 U22959 ( .A1(n21042), .A2(n21041), .ZN(n21112) );
  INV_X1 U22960 ( .A(n21129), .ZN(n21043) );
  OAI21_X1 U22961 ( .B1(n21112), .B2(n11276), .A(n21043), .ZN(n21064) );
  OAI22_X1 U22962 ( .A1(n21112), .A2(n21184), .B1(n21044), .B2(n21149), .ZN(
        n21045) );
  NOR4_X1 U22963 ( .A1(n21046), .A2(n21064), .A3(n21124), .A4(n21045), .ZN(
        n21047) );
  OAI22_X1 U22964 ( .A1(n21049), .A2(n21048), .B1(n21047), .B2(n21234), .ZN(
        n21053) );
  NAND2_X1 U22965 ( .A1(n21051), .A2(n21050), .ZN(n21132) );
  INV_X1 U22966 ( .A(n21112), .ZN(n21058) );
  NOR2_X1 U22967 ( .A1(n21132), .A2(n21058), .ZN(n21052) );
  AOI222_X1 U22968 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n21053), 
        .B1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n21133), .C1(n21053), 
        .C2(n21052), .ZN(n21055) );
  OAI211_X1 U22969 ( .C1(n21056), .C2(n21246), .A(n21055), .B(n21054), .ZN(
        P3_U2835) );
  NOR4_X1 U22970 ( .A1(n21060), .A2(n21059), .A3(n21058), .A4(n21057), .ZN(
        n21090) );
  NOR2_X1 U22971 ( .A1(n21147), .A2(n21061), .ZN(n21062) );
  AOI211_X1 U22972 ( .C1(n21107), .C2(n21177), .A(n21090), .B(n21062), .ZN(
        n21083) );
  NAND2_X1 U22973 ( .A1(n21117), .A2(n21082), .ZN(n21075) );
  NAND3_X1 U22974 ( .A1(n21112), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A3(
        n21063), .ZN(n21065) );
  AOI211_X1 U22975 ( .C1(n21231), .C2(n21065), .A(n21173), .B(n21064), .ZN(
        n21079) );
  NAND2_X1 U22976 ( .A1(n21237), .A2(n21065), .ZN(n21077) );
  OAI211_X1 U22977 ( .C1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n11276), .A(
        n21079), .B(n21077), .ZN(n21110) );
  AOI22_X1 U22978 ( .A1(n21177), .A2(n21067), .B1(n21254), .B2(n21066), .ZN(
        n21068) );
  INV_X1 U22979 ( .A(n21068), .ZN(n21085) );
  AOI211_X1 U22980 ( .C1(n21069), .C2(n21141), .A(n21110), .B(n21085), .ZN(
        n21070) );
  OAI21_X1 U22981 ( .B1(n21070), .B2(n21234), .A(n21220), .ZN(n21071) );
  AOI22_X1 U22982 ( .A1(n21203), .A2(n21072), .B1(
        P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n21071), .ZN(n21074) );
  OAI211_X1 U22983 ( .C1(n21083), .C2(n21075), .A(n21074), .B(n21073), .ZN(
        P3_U2833) );
  AOI22_X1 U22984 ( .A1(n21133), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B1(
        n21203), .B2(n21076), .ZN(n21087) );
  AND2_X1 U22985 ( .A1(n21078), .A2(n21077), .ZN(n21080) );
  OAI211_X1 U22986 ( .C1(n21201), .C2(n21080), .A(n21079), .B(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n21093) );
  OAI21_X1 U22987 ( .B1(n21083), .B2(n21082), .A(n21081), .ZN(n21084) );
  OAI211_X1 U22988 ( .C1(n21093), .C2(n21085), .A(n21117), .B(n21084), .ZN(
        n21086) );
  OAI211_X1 U22989 ( .C1(n21088), .C2(n21223), .A(n21087), .B(n21086), .ZN(
        P3_U2832) );
  NOR2_X1 U22990 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n21089), .ZN(
        n21091) );
  AOI22_X1 U22991 ( .A1(n21254), .A2(n21092), .B1(n21091), .B2(n21090), .ZN(
        n21095) );
  NAND3_X1 U22992 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n21141), .A3(
        n21093), .ZN(n21094) );
  OAI211_X1 U22993 ( .C1(n21096), .C2(n21149), .A(n21095), .B(n21094), .ZN(
        n21098) );
  AOI22_X1 U22994 ( .A1(n21117), .A2(n21098), .B1(n21203), .B2(n21097), .ZN(
        n21101) );
  INV_X1 U22995 ( .A(n21099), .ZN(n21100) );
  OAI211_X1 U22996 ( .C1(n21102), .C2(n21220), .A(n21101), .B(n21100), .ZN(
        P3_U2831) );
  NAND2_X1 U22997 ( .A1(n21104), .A2(n21103), .ZN(n21114) );
  AOI221_X1 U22998 ( .B1(n21106), .B2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), 
        .C1(n21114), .C2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A(n21105), .ZN(
        n21111) );
  OAI22_X1 U22999 ( .A1(n21108), .A2(n21147), .B1(n21107), .B2(n21149), .ZN(
        n21109) );
  NOR4_X1 U23000 ( .A1(n21111), .A2(n21133), .A3(n21110), .A4(n21109), .ZN(
        n21123) );
  NAND2_X1 U23001 ( .A1(n21112), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n21113) );
  OAI22_X1 U23002 ( .A1(n21115), .A2(n21114), .B1(n21132), .B2(n21113), .ZN(
        n21116) );
  OAI221_X1 U23003 ( .B1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n21117), 
        .C1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .C2(n21116), .A(n21223), .ZN(
        n21122) );
  OR3_X1 U23004 ( .A1(n21119), .A2(n21246), .A3(n21118), .ZN(n21121) );
  OAI211_X1 U23005 ( .C1(n21123), .C2(n21122), .A(n21121), .B(n21120), .ZN(
        P3_U2834) );
  INV_X1 U23006 ( .A(n21124), .ZN(n21128) );
  AOI22_X1 U23007 ( .A1(n21177), .A2(n21126), .B1(n21254), .B2(n21125), .ZN(
        n21127) );
  NAND3_X1 U23008 ( .A1(n21128), .A2(n21127), .A3(n21220), .ZN(n21140) );
  NOR3_X1 U23009 ( .A1(n21129), .A2(n21131), .A3(n21140), .ZN(n21130) );
  NOR2_X1 U23010 ( .A1(n21238), .A2(n21130), .ZN(n21139) );
  OAI21_X1 U23011 ( .B1(n21133), .B2(n21132), .A(n21131), .ZN(n21134) );
  AOI22_X1 U23012 ( .A1(n21238), .A2(P3_REIP_REG_23__SCAN_IN), .B1(n21139), 
        .B2(n21134), .ZN(n21135) );
  OAI21_X1 U23013 ( .B1(n21246), .B2(n21136), .A(n21135), .ZN(P3_U2839) );
  NOR3_X1 U23014 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n21234), .A3(
        n21137), .ZN(n21138) );
  AOI21_X1 U23015 ( .B1(P3_REIP_REG_24__SCAN_IN), .B2(n21238), .A(n21138), 
        .ZN(n21143) );
  OAI211_X1 U23016 ( .C1(n21141), .C2(n21140), .A(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B(n21139), .ZN(n21142) );
  OAI211_X1 U23017 ( .C1(n21144), .C2(n21246), .A(n21143), .B(n21142), .ZN(
        P3_U2838) );
  INV_X1 U23018 ( .A(n21145), .ZN(n21154) );
  INV_X1 U23019 ( .A(n21146), .ZN(n21153) );
  OAI22_X1 U23020 ( .A1(n21150), .A2(n21149), .B1(n21148), .B2(n21147), .ZN(
        n21151) );
  INV_X1 U23021 ( .A(n21151), .ZN(n21152) );
  NAND3_X1 U23022 ( .A1(n21154), .A2(n21153), .A3(n21152), .ZN(n21155) );
  NAND2_X1 U23023 ( .A1(n21223), .A2(n21155), .ZN(n21159) );
  AOI22_X1 U23024 ( .A1(n21238), .A2(P3_REIP_REG_19__SCAN_IN), .B1(n21203), 
        .B2(n21156), .ZN(n21157) );
  OAI221_X1 U23025 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n21166), 
        .C1(n21158), .C2(n21159), .A(n21157), .ZN(P3_U2843) );
  NAND2_X1 U23026 ( .A1(n21158), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n21160) );
  OAI21_X1 U23027 ( .B1(n21161), .B2(n21160), .A(n21159), .ZN(n21163) );
  AOI22_X1 U23028 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n21163), .B1(
        n21203), .B2(n21162), .ZN(n21164) );
  OAI211_X1 U23029 ( .C1(n21167), .C2(n21166), .A(n21165), .B(n21164), .ZN(
        P3_U2842) );
  NAND2_X1 U23030 ( .A1(n21168), .A2(n21242), .ZN(n21207) );
  AOI21_X1 U23031 ( .B1(n21170), .B2(n21169), .A(n11276), .ZN(n21182) );
  NOR4_X1 U23032 ( .A1(n21173), .A2(n21198), .A3(n21172), .A4(n21171), .ZN(
        n21180) );
  AOI211_X1 U23033 ( .C1(n21177), .C2(n21176), .A(n21175), .B(n21174), .ZN(
        n21178) );
  OAI22_X1 U23034 ( .A1(n21184), .A2(n21180), .B1(n21179), .B2(n21178), .ZN(
        n21181) );
  NOR3_X1 U23035 ( .A1(n21182), .A2(n21234), .A3(n21181), .ZN(n21192) );
  AOI221_X1 U23036 ( .B1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n21192), 
        .C1(n21184), .C2(n21192), .A(n21183), .ZN(n21185) );
  AOI22_X1 U23037 ( .A1(n21186), .A2(n21203), .B1(n21185), .B2(n21223), .ZN(
        n21188) );
  OAI211_X1 U23038 ( .C1(n21207), .C2(n21189), .A(n21188), .B(n21187), .ZN(
        P3_U2844) );
  NOR2_X1 U23039 ( .A1(n21223), .A2(n21190), .ZN(n21194) );
  NOR3_X1 U23040 ( .A1(n21238), .A2(n21192), .A3(n21191), .ZN(n21193) );
  AOI211_X1 U23041 ( .C1(n21203), .C2(n21195), .A(n21194), .B(n21193), .ZN(
        n21196) );
  OAI21_X1 U23042 ( .B1(n21207), .B2(n21197), .A(n21196), .ZN(P3_U2845) );
  AOI221_X1 U23043 ( .B1(n21201), .B2(n21200), .C1(n21199), .C2(n21200), .A(
        n21198), .ZN(n21202) );
  AOI22_X1 U23044 ( .A1(n21204), .A2(n21203), .B1(n21202), .B2(n21223), .ZN(
        n21206) );
  OAI211_X1 U23045 ( .C1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .C2(n21207), .A(
        n21206), .B(n21205), .ZN(P3_U2846) );
  AOI22_X1 U23046 ( .A1(n21238), .A2(P3_REIP_REG_13__SCAN_IN), .B1(n21242), 
        .B2(n21208), .ZN(n21215) );
  OAI21_X1 U23047 ( .B1(n11379), .B2(n21209), .A(n21237), .ZN(n21210) );
  NAND3_X1 U23048 ( .A1(n21211), .A2(n21220), .A3(n21210), .ZN(n21212) );
  OAI211_X1 U23049 ( .C1(n21213), .C2(n21212), .A(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B(n21223), .ZN(n21214) );
  OAI211_X1 U23050 ( .C1(n21216), .C2(n21246), .A(n21215), .B(n21214), .ZN(
        P3_U2849) );
  NOR2_X1 U23051 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n21241), .ZN(
        n21217) );
  AOI22_X1 U23052 ( .A1(n21238), .A2(P3_REIP_REG_10__SCAN_IN), .B1(n21242), 
        .B2(n21217), .ZN(n21227) );
  OR2_X1 U23053 ( .A1(n21219), .A2(n21218), .ZN(n21221) );
  OAI211_X1 U23054 ( .C1(n21222), .C2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n21221), .B(n21220), .ZN(n21224) );
  OAI211_X1 U23055 ( .C1(n21225), .C2(n21224), .A(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B(n21223), .ZN(n21226) );
  OAI211_X1 U23056 ( .C1(n21228), .C2(n21246), .A(n21227), .B(n21226), .ZN(
        P3_U2852) );
  OAI211_X1 U23057 ( .C1(n21232), .C2(n21231), .A(n21230), .B(n21229), .ZN(
        n21233) );
  INV_X1 U23058 ( .A(n21233), .ZN(n21235) );
  AOI211_X1 U23059 ( .C1(n21237), .C2(n21236), .A(n21235), .B(n21234), .ZN(
        n21239) );
  AOI21_X1 U23060 ( .B1(n21240), .B2(n21239), .A(n21238), .ZN(n21243) );
  AOI22_X1 U23061 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n21243), .B1(
        n21242), .B2(n21241), .ZN(n21245) );
  OAI211_X1 U23062 ( .C1(n21247), .C2(n21246), .A(n21245), .B(n21244), .ZN(
        P3_U2853) );
  NAND2_X1 U23063 ( .A1(n21707), .A2(n21248), .ZN(n21298) );
  OAI22_X1 U23064 ( .A1(n21252), .A2(n21251), .B1(n21250), .B2(n21249), .ZN(
        n21253) );
  AOI221_X1 U23065 ( .B1(n21256), .B2(n21255), .C1(n21254), .C2(n21255), .A(
        n21253), .ZN(n21313) );
  AOI211_X1 U23066 ( .C1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .C2(n21271), .A(
        n21258), .B(n21257), .ZN(n21285) );
  AOI22_X1 U23067 ( .A1(n21271), .A2(n21260), .B1(n21259), .B2(n21269), .ZN(
        n21278) );
  NOR3_X1 U23068 ( .A1(n21263), .A2(n21262), .A3(n21261), .ZN(n21265) );
  OAI22_X1 U23069 ( .A1(n21266), .A2(n21265), .B1(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n21264), .ZN(n21268) );
  AOI21_X1 U23070 ( .B1(n21268), .B2(n21269), .A(n21267), .ZN(n21273) );
  AOI22_X1 U23071 ( .A1(n21271), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n21270), .B2(n21269), .ZN(n21274) );
  OR2_X1 U23072 ( .A1(n21274), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n21272) );
  AOI221_X1 U23073 ( .B1(n21273), .B2(n21272), .C1(n21274), .C2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n21277) );
  OAI21_X1 U23074 ( .B1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(n21274), .ZN(n21276) );
  AOI222_X1 U23075 ( .A1(n21278), .A2(n21277), .B1(n21278), .B2(n21276), .C1(
        n21277), .C2(n21275), .ZN(n21284) );
  INV_X1 U23076 ( .A(n21279), .ZN(n21282) );
  NOR3_X1 U23077 ( .A1(n21282), .A2(n21281), .A3(n21280), .ZN(n21311) );
  OAI21_X1 U23078 ( .B1(P3_FLUSH_REG_SCAN_IN), .B2(P3_MORE_REG_SCAN_IN), .A(
        n21311), .ZN(n21283) );
  NAND4_X1 U23079 ( .A1(n21313), .A2(n21285), .A3(n21284), .A4(n21283), .ZN(
        n21304) );
  AOI211_X1 U23080 ( .C1(n21287), .C2(n21286), .A(n21310), .B(n21304), .ZN(
        n21294) );
  AOI21_X1 U23081 ( .B1(n21707), .B2(n21288), .A(n21294), .ZN(n21308) );
  NAND3_X1 U23082 ( .A1(n21290), .A2(n21308), .A3(n21289), .ZN(n21291) );
  NAND4_X1 U23083 ( .A1(n21293), .A2(n21298), .A3(n21292), .A4(n21291), .ZN(
        P3_U2997) );
  NOR2_X1 U23084 ( .A1(n21294), .A2(n21309), .ZN(n21297) );
  OAI21_X1 U23085 ( .B1(n21297), .B2(n21296), .A(n21295), .ZN(P3_U3282) );
  INV_X1 U23086 ( .A(n21298), .ZN(n21299) );
  AOI211_X1 U23087 ( .C1(n21301), .C2(n21300), .A(P3_STATE2_REG_0__SCAN_IN), 
        .B(n21299), .ZN(n21302) );
  AOI211_X1 U23088 ( .C1(n21305), .C2(n21304), .A(n21303), .B(n21302), .ZN(
        n21306) );
  OAI221_X1 U23089 ( .B1(n21309), .B2(n21308), .C1(n21309), .C2(n21307), .A(
        n21306), .ZN(P3_U2996) );
  NOR2_X1 U23090 ( .A1(n21311), .A2(n21310), .ZN(n21317) );
  INV_X1 U23091 ( .A(n21317), .ZN(n21314) );
  NAND2_X1 U23092 ( .A1(n21314), .A2(P3_MORE_REG_SCAN_IN), .ZN(n21312) );
  OAI21_X1 U23093 ( .B1(n21314), .B2(n21313), .A(n21312), .ZN(P3_U3295) );
  OAI21_X1 U23094 ( .B1(n21317), .B2(n21316), .A(n21315), .ZN(P3_U2637) );
  AOI211_X1 U23095 ( .C1(n21319), .C2(n14152), .A(n21910), .B(n21318), .ZN(
        n21322) );
  OAI21_X1 U23096 ( .B1(n21322), .B2(n21321), .A(n21320), .ZN(n21327) );
  AOI211_X1 U23097 ( .C1(n21325), .C2(n21675), .A(n21324), .B(n21323), .ZN(
        n21326) );
  MUX2_X1 U23098 ( .A(n21327), .B(P1_REQUESTPENDING_REG_SCAN_IN), .S(n21326), 
        .Z(P1_U3485) );
  INV_X1 U23099 ( .A(n21328), .ZN(n21332) );
  NOR2_X1 U23100 ( .A1(n21386), .A2(n21522), .ZN(n21330) );
  AOI211_X1 U23101 ( .C1(n21332), .C2(n21331), .A(n21330), .B(n21329), .ZN(
        n21336) );
  INV_X1 U23102 ( .A(n21333), .ZN(n21334) );
  AOI22_X1 U23103 ( .A1(n21334), .A2(n21410), .B1(n21409), .B2(n21520), .ZN(
        n21335) );
  OAI211_X1 U23104 ( .C1(n21338), .C2(n21337), .A(n21336), .B(n21335), .ZN(
        P1_U3018) );
  INV_X1 U23105 ( .A(n21339), .ZN(n21345) );
  INV_X1 U23106 ( .A(n21340), .ZN(n21499) );
  AOI21_X1 U23107 ( .B1(n21409), .B2(n21499), .A(n21341), .ZN(n21342) );
  OAI21_X1 U23108 ( .B1(n21343), .B2(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n21342), .ZN(n21344) );
  AOI21_X1 U23109 ( .B1(n21345), .B2(n21410), .A(n21344), .ZN(n21346) );
  OAI21_X1 U23110 ( .B1(n21348), .B2(n21347), .A(n21346), .ZN(P1_U3020) );
  OAI21_X1 U23111 ( .B1(n21351), .B2(n21350), .A(n21349), .ZN(n21362) );
  NOR2_X1 U23112 ( .A1(n21386), .A2(n21569), .ZN(n21356) );
  OAI22_X1 U23113 ( .A1(n21354), .A2(n21353), .B1(n21352), .B2(n21559), .ZN(
        n21355) );
  AOI211_X1 U23114 ( .C1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .C2(n21362), .A(
        n21356), .B(n21355), .ZN(n21357) );
  OAI21_X1 U23115 ( .B1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n21358), .A(
        n21357), .ZN(P1_U3013) );
  INV_X1 U23116 ( .A(n21359), .ZN(n21361) );
  AOI22_X1 U23117 ( .A1(n21361), .A2(n21410), .B1(n21409), .B2(n21360), .ZN(
        n21365) );
  OAI21_X1 U23118 ( .B1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n21363), .A(
        n21362), .ZN(n21364) );
  OAI211_X1 U23119 ( .C1(n21366), .C2(n21386), .A(n21365), .B(n21364), .ZN(
        P1_U3014) );
  INV_X1 U23120 ( .A(n21367), .ZN(n21369) );
  INV_X1 U23121 ( .A(n21368), .ZN(n21570) );
  AOI22_X1 U23122 ( .A1(n21369), .A2(n21410), .B1(n21409), .B2(n21570), .ZN(
        n21374) );
  NAND2_X1 U23123 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n21370), .ZN(
        n21371) );
  OAI21_X1 U23124 ( .B1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n21372), .A(
        n21371), .ZN(n21373) );
  OAI211_X1 U23125 ( .C1(n21582), .C2(n21386), .A(n21374), .B(n21373), .ZN(
        P1_U3012) );
  AOI22_X1 U23126 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n21375), .B1(
        n10970), .B2(P1_REIP_REG_21__SCAN_IN), .ZN(n21380) );
  INV_X1 U23127 ( .A(n21376), .ZN(n21377) );
  AOI22_X1 U23128 ( .A1(n21377), .A2(n21410), .B1(n21409), .B2(n21591), .ZN(
        n21379) );
  NAND3_X1 U23129 ( .A1(n21380), .A2(n21379), .A3(n21378), .ZN(P1_U3010) );
  INV_X1 U23130 ( .A(n21381), .ZN(n21384) );
  INV_X1 U23131 ( .A(n21382), .ZN(n21383) );
  AOI22_X1 U23132 ( .A1(n21384), .A2(n21410), .B1(n21409), .B2(n21383), .ZN(
        n21392) );
  INV_X1 U23133 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n21388) );
  NOR2_X1 U23134 ( .A1(n21386), .A2(n21385), .ZN(n21387) );
  AOI221_X1 U23135 ( .B1(n21390), .B2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), 
        .C1(n21389), .C2(n21388), .A(n21387), .ZN(n21391) );
  NAND2_X1 U23136 ( .A1(n21392), .A2(n21391), .ZN(P1_U3004) );
  AOI21_X1 U23137 ( .B1(P1_REIP_REG_25__SCAN_IN), .B2(n10970), .A(n21393), 
        .ZN(n21397) );
  INV_X1 U23138 ( .A(n21394), .ZN(n21395) );
  AOI22_X1 U23139 ( .A1(n21395), .A2(n21410), .B1(n21409), .B2(n21632), .ZN(
        n21396) );
  OAI211_X1 U23140 ( .C1(n21399), .C2(n21398), .A(n21397), .B(n21396), .ZN(
        P1_U3006) );
  AOI22_X1 U23141 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n21400), .B1(
        n10970), .B2(P1_REIP_REG_23__SCAN_IN), .ZN(n21405) );
  INV_X1 U23142 ( .A(n21401), .ZN(n21403) );
  AOI22_X1 U23143 ( .A1(n21403), .A2(n21410), .B1(n21409), .B2(n21402), .ZN(
        n21404) );
  OAI211_X1 U23144 ( .C1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n21406), .A(
        n21405), .B(n21404), .ZN(P1_U3008) );
  INV_X1 U23145 ( .A(n21407), .ZN(n21408) );
  AOI22_X1 U23146 ( .A1(n21411), .A2(n21410), .B1(n21409), .B2(n21408), .ZN(
        n21419) );
  NAND3_X1 U23147 ( .A1(n21658), .A2(n21413), .A3(n21412), .ZN(n21414) );
  OAI21_X1 U23148 ( .B1(n21416), .B2(n21415), .A(n21414), .ZN(n21417) );
  NAND3_X1 U23149 ( .A1(n21419), .A2(n21418), .A3(n21417), .ZN(P1_U3031) );
  OAI22_X1 U23150 ( .A1(n10973), .A2(n21431), .B1(n21439), .B2(
        P1_REIP_REG_1__SCAN_IN), .ZN(n21420) );
  INV_X1 U23151 ( .A(n21420), .ZN(n21421) );
  OAI21_X1 U23152 ( .B1(n21422), .B2(n19947), .A(n21421), .ZN(n21423) );
  AOI21_X1 U23153 ( .B1(n21645), .B2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n21423), .ZN(n21430) );
  INV_X1 U23154 ( .A(n21424), .ZN(n21426) );
  OAI22_X1 U23155 ( .A1(n21426), .A2(n21646), .B1(n21425), .B2(n21640), .ZN(
        n21427) );
  AOI21_X1 U23156 ( .B1(n21428), .B2(n21449), .A(n21427), .ZN(n21429) );
  OAI211_X1 U23157 ( .C1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n21642), .A(
        n21430), .B(n21429), .ZN(P1_U2839) );
  OAI21_X1 U23158 ( .B1(n21432), .B2(n21431), .A(n21571), .ZN(n21436) );
  OAI22_X1 U23159 ( .A1(n21434), .A2(n21640), .B1(n21646), .B2(n21433), .ZN(
        n21435) );
  AOI211_X1 U23160 ( .C1(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .C2(n21645), .A(
        n21436), .B(n21435), .ZN(n21443) );
  NAND3_X1 U23161 ( .A1(P1_REIP_REG_2__SCAN_IN), .A2(P1_REIP_REG_1__SCAN_IN), 
        .A3(P1_REIP_REG_3__SCAN_IN), .ZN(n21438) );
  OAI21_X1 U23162 ( .B1(n21439), .B2(n21438), .A(n21437), .ZN(n21440) );
  AOI22_X1 U23163 ( .A1(n21441), .A2(n21449), .B1(n10994), .B2(n21440), .ZN(
        n21442) );
  OAI211_X1 U23164 ( .C1(n21444), .C2(n21642), .A(n21443), .B(n21442), .ZN(
        P1_U2836) );
  AOI22_X1 U23165 ( .A1(P1_EBX_REG_5__SCAN_IN), .A2(n21626), .B1(
        P1_REIP_REG_5__SCAN_IN), .B2(n10994), .ZN(n21452) );
  INV_X1 U23166 ( .A(n21445), .ZN(n21450) );
  AOI22_X1 U23167 ( .A1(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n21645), .B1(
        n11065), .B2(n11382), .ZN(n21446) );
  OAI211_X1 U23168 ( .C1(n21642), .C2(n21447), .A(n21446), .B(n21571), .ZN(
        n21448) );
  AOI21_X1 U23169 ( .B1(n21450), .B2(n21449), .A(n21448), .ZN(n21451) );
  OAI211_X1 U23170 ( .C1(n21646), .C2(n21453), .A(n21452), .B(n21451), .ZN(
        P1_U2835) );
  OAI22_X1 U23171 ( .A1(n21455), .A2(n21640), .B1(n21646), .B2(n21454), .ZN(
        n21456) );
  AOI211_X1 U23172 ( .C1(n21645), .C2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n21562), .B(n21456), .ZN(n21466) );
  INV_X1 U23173 ( .A(n21457), .ZN(n21464) );
  NOR4_X1 U23174 ( .A1(n21459), .A2(n11382), .A3(n21458), .A4(n21463), .ZN(
        n21489) );
  NOR2_X1 U23175 ( .A1(n21523), .A2(n21489), .ZN(n21472) );
  OAI22_X1 U23176 ( .A1(n21461), .A2(n21648), .B1(n21460), .B2(n21642), .ZN(
        n21462) );
  AOI221_X1 U23177 ( .B1(n21464), .B2(n21463), .C1(n21472), .C2(
        P1_REIP_REG_6__SCAN_IN), .A(n21462), .ZN(n21465) );
  NAND2_X1 U23178 ( .A1(n21466), .A2(n21465), .ZN(P1_U2834) );
  OAI21_X1 U23179 ( .B1(n21636), .B2(n21467), .A(n21571), .ZN(n21471) );
  OAI22_X1 U23180 ( .A1(n21469), .A2(n21640), .B1(n21646), .B2(n21468), .ZN(
        n21470) );
  AOI211_X1 U23181 ( .C1(P1_REIP_REG_7__SCAN_IN), .C2(n21472), .A(n21471), .B(
        n21470), .ZN(n21476) );
  AOI22_X1 U23182 ( .A1(n21474), .A2(n21611), .B1(n21488), .B2(n21473), .ZN(
        n21475) );
  OAI211_X1 U23183 ( .C1(n21477), .C2(n21642), .A(n21476), .B(n21475), .ZN(
        P1_U2833) );
  AOI22_X1 U23184 ( .A1(n21478), .A2(n21627), .B1(P1_EBX_REG_9__SCAN_IN), .B2(
        n21626), .ZN(n21479) );
  OAI211_X1 U23185 ( .C1(n21636), .C2(n21480), .A(n21479), .B(n21571), .ZN(
        n21481) );
  AOI21_X1 U23186 ( .B1(n21633), .B2(n21482), .A(n21481), .ZN(n21486) );
  AND2_X1 U23187 ( .A1(P1_REIP_REG_9__SCAN_IN), .A2(n21487), .ZN(n21483) );
  AOI22_X1 U23188 ( .A1(n21484), .A2(n21611), .B1(n21483), .B2(n21639), .ZN(
        n21485) );
  OAI211_X1 U23189 ( .C1(P1_REIP_REG_9__SCAN_IN), .C2(n21487), .A(n21486), .B(
        n21485), .ZN(P1_U2831) );
  NAND4_X1 U23190 ( .A1(P1_REIP_REG_9__SCAN_IN), .A2(P1_REIP_REG_8__SCAN_IN), 
        .A3(P1_REIP_REG_7__SCAN_IN), .A4(n21488), .ZN(n21498) );
  NAND2_X1 U23191 ( .A1(n21490), .A2(n21489), .ZN(n21508) );
  AND2_X1 U23192 ( .A1(n21639), .A2(n21508), .ZN(n21500) );
  AOI22_X1 U23193 ( .A1(P1_EBX_REG_10__SCAN_IN), .A2(n21626), .B1(
        P1_REIP_REG_10__SCAN_IN), .B2(n21500), .ZN(n21491) );
  OAI21_X1 U23194 ( .B1(n21646), .B2(n21492), .A(n21491), .ZN(n21493) );
  AOI211_X1 U23195 ( .C1(n21645), .C2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n21562), .B(n21493), .ZN(n21497) );
  AOI22_X1 U23196 ( .A1(n21495), .A2(n21611), .B1(n21494), .B2(n21627), .ZN(
        n21496) );
  OAI211_X1 U23197 ( .C1(P1_REIP_REG_10__SCAN_IN), .C2(n21498), .A(n21497), 
        .B(n21496), .ZN(P1_U2830) );
  AOI22_X1 U23198 ( .A1(P1_REIP_REG_11__SCAN_IN), .A2(n21500), .B1(n21633), 
        .B2(n21499), .ZN(n21501) );
  OAI211_X1 U23199 ( .C1(n21636), .C2(n11909), .A(n21501), .B(n21571), .ZN(
        n21505) );
  OAI22_X1 U23200 ( .A1(n21503), .A2(n21642), .B1(n21648), .B2(n21502), .ZN(
        n21504) );
  AOI211_X1 U23201 ( .C1(P1_EBX_REG_11__SCAN_IN), .C2(n21626), .A(n21505), .B(
        n21504), .ZN(n21506) );
  OAI21_X1 U23202 ( .B1(P1_REIP_REG_11__SCAN_IN), .B2(n21507), .A(n21506), 
        .ZN(P1_U2829) );
  NOR2_X1 U23203 ( .A1(n21509), .A2(n21508), .ZN(n21524) );
  NOR3_X1 U23204 ( .A1(n21523), .A2(n21524), .A3(n21514), .ZN(n21510) );
  AOI211_X1 U23205 ( .C1(n21645), .C2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n21562), .B(n21510), .ZN(n21511) );
  OAI21_X1 U23206 ( .B1(n21646), .B2(n21512), .A(n21511), .ZN(n21513) );
  AOI21_X1 U23207 ( .B1(P1_EBX_REG_12__SCAN_IN), .B2(n21626), .A(n21513), .ZN(
        n21518) );
  AOI22_X1 U23208 ( .A1(n21516), .A2(n21627), .B1(n21515), .B2(n21514), .ZN(
        n21517) );
  OAI211_X1 U23209 ( .C1(n21648), .C2(n21519), .A(n21518), .B(n21517), .ZN(
        P1_U2828) );
  AOI22_X1 U23210 ( .A1(n21520), .A2(n21633), .B1(n21626), .B2(
        P1_EBX_REG_13__SCAN_IN), .ZN(n21521) );
  NAND2_X1 U23211 ( .A1(n21521), .A2(n21571), .ZN(n21526) );
  AOI211_X1 U23212 ( .C1(P1_REIP_REG_12__SCAN_IN), .C2(n21524), .A(n21523), 
        .B(n21522), .ZN(n21525) );
  AOI211_X1 U23213 ( .C1(n21645), .C2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .A(
        n21526), .B(n21525), .ZN(n21527) );
  OAI21_X1 U23214 ( .B1(n21528), .B2(n21648), .A(n21527), .ZN(n21529) );
  AOI21_X1 U23215 ( .B1(n21530), .B2(n21627), .A(n21529), .ZN(n21531) );
  OAI21_X1 U23216 ( .B1(P1_REIP_REG_13__SCAN_IN), .B2(n21532), .A(n21531), 
        .ZN(P1_U2827) );
  AOI22_X1 U23217 ( .A1(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n21645), .B1(
        P1_EBX_REG_14__SCAN_IN), .B2(n21626), .ZN(n21540) );
  AOI21_X1 U23218 ( .B1(n21533), .B2(n21633), .A(n21562), .ZN(n21539) );
  AOI22_X1 U23219 ( .A1(n21535), .A2(n21611), .B1(n21627), .B2(n21534), .ZN(
        n21538) );
  OAI211_X1 U23220 ( .C1(n21536), .C2(P1_REIP_REG_14__SCAN_IN), .A(n21639), 
        .B(n21541), .ZN(n21537) );
  NAND4_X1 U23221 ( .A1(n21540), .A2(n21539), .A3(n21538), .A4(n21537), .ZN(
        P1_U2826) );
  AOI21_X1 U23222 ( .B1(P1_REIP_REG_15__SCAN_IN), .B2(n21639), .A(n11366), 
        .ZN(n21550) );
  OAI22_X1 U23223 ( .A1(n21543), .A2(n21636), .B1(n21542), .B2(n21640), .ZN(
        n21544) );
  AOI211_X1 U23224 ( .C1(n21627), .C2(n21545), .A(n21562), .B(n21544), .ZN(
        n21549) );
  AOI22_X1 U23225 ( .A1(n21547), .A2(n21611), .B1(n21633), .B2(n21546), .ZN(
        n21548) );
  OAI211_X1 U23226 ( .C1(n21555), .C2(n21550), .A(n21549), .B(n21548), .ZN(
        P1_U2825) );
  AOI22_X1 U23227 ( .A1(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n21645), .B1(
        P1_EBX_REG_16__SCAN_IN), .B2(n21626), .ZN(n21551) );
  OAI211_X1 U23228 ( .C1(n21642), .C2(n21552), .A(n21551), .B(n21571), .ZN(
        n21553) );
  AOI21_X1 U23229 ( .B1(n21554), .B2(n21611), .A(n21553), .ZN(n21557) );
  OAI211_X1 U23230 ( .C1(n21555), .C2(P1_REIP_REG_16__SCAN_IN), .A(n21639), 
        .B(n11009), .ZN(n21556) );
  OAI211_X1 U23231 ( .C1(n21558), .C2(n21646), .A(n21557), .B(n21556), .ZN(
        P1_U2824) );
  OAI22_X1 U23232 ( .A1(n21560), .A2(n21640), .B1(n21646), .B2(n21559), .ZN(
        n21561) );
  AOI211_X1 U23233 ( .C1(n21645), .C2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n21562), .B(n21561), .ZN(n21564) );
  NAND2_X1 U23234 ( .A1(n21563), .A2(n21569), .ZN(n21580) );
  OAI211_X1 U23235 ( .C1(n21565), .C2(n21642), .A(n21564), .B(n21580), .ZN(
        n21566) );
  AOI21_X1 U23236 ( .B1(n21567), .B2(n21611), .A(n21566), .ZN(n21568) );
  OAI21_X1 U23237 ( .B1(n21569), .B2(n21581), .A(n21568), .ZN(P1_U2822) );
  AOI22_X1 U23238 ( .A1(P1_EBX_REG_19__SCAN_IN), .A2(n21626), .B1(n21633), 
        .B2(n21570), .ZN(n21572) );
  OAI211_X1 U23239 ( .C1(n21636), .C2(n21573), .A(n21572), .B(n21571), .ZN(
        n21577) );
  OAI22_X1 U23240 ( .A1(n21575), .A2(n21648), .B1(P1_REIP_REG_19__SCAN_IN), 
        .B2(n21574), .ZN(n21576) );
  AOI211_X1 U23241 ( .C1(n21578), .C2(n21627), .A(n21577), .B(n21576), .ZN(
        n21579) );
  OAI221_X1 U23242 ( .B1(n21582), .B2(n21581), .C1(n21582), .C2(n21580), .A(
        n21579), .ZN(P1_U2821) );
  AOI22_X1 U23243 ( .A1(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n21645), .B1(
        P1_EBX_REG_20__SCAN_IN), .B2(n21626), .ZN(n21589) );
  NAND2_X1 U23244 ( .A1(n21600), .A2(n21639), .ZN(n21599) );
  INV_X1 U23245 ( .A(n21599), .ZN(n21586) );
  OAI22_X1 U23246 ( .A1(n21584), .A2(n21648), .B1(n21646), .B2(n21583), .ZN(
        n21585) );
  AOI221_X1 U23247 ( .B1(n21587), .B2(n21586), .C1(P1_REIP_REG_20__SCAN_IN), 
        .C2(n21586), .A(n21585), .ZN(n21588) );
  OAI211_X1 U23248 ( .C1(n21590), .C2(n21642), .A(n21589), .B(n21588), .ZN(
        P1_U2820) );
  AOI22_X1 U23249 ( .A1(P1_EBX_REG_21__SCAN_IN), .A2(n21626), .B1(n21633), 
        .B2(n21591), .ZN(n21592) );
  OAI21_X1 U23250 ( .B1(n21593), .B2(n21636), .A(n21592), .ZN(n21596) );
  OAI22_X1 U23251 ( .A1(n21594), .A2(n21648), .B1(P1_REIP_REG_21__SCAN_IN), 
        .B2(n21600), .ZN(n21595) );
  AOI211_X1 U23252 ( .C1(n21597), .C2(n21627), .A(n21596), .B(n21595), .ZN(
        n21598) );
  OAI21_X1 U23253 ( .B1(n21601), .B2(n21599), .A(n21598), .ZN(P1_U2819) );
  AOI22_X1 U23254 ( .A1(n21602), .A2(n21601), .B1(n21600), .B2(n21639), .ZN(
        n21614) );
  INV_X1 U23255 ( .A(n21603), .ZN(n21612) );
  NOR2_X1 U23256 ( .A1(n21604), .A2(n21646), .ZN(n21610) );
  INV_X1 U23257 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n21608) );
  INV_X1 U23258 ( .A(n21605), .ZN(n21606) );
  AOI22_X1 U23259 ( .A1(n21627), .A2(n21606), .B1(n21626), .B2(
        P1_EBX_REG_22__SCAN_IN), .ZN(n21607) );
  OAI21_X1 U23260 ( .B1(n21608), .B2(n21636), .A(n21607), .ZN(n21609) );
  AOI211_X1 U23261 ( .C1(n21612), .C2(n21611), .A(n21610), .B(n21609), .ZN(
        n21613) );
  OAI221_X1 U23262 ( .B1(P1_REIP_REG_22__SCAN_IN), .B2(n11051), .C1(n21615), 
        .C2(n21614), .A(n21613), .ZN(P1_U2818) );
  AOI21_X1 U23263 ( .B1(P1_REIP_REG_24__SCAN_IN), .B2(n21639), .A(n21617), 
        .ZN(n21625) );
  OAI22_X1 U23264 ( .A1(n21619), .A2(n21642), .B1(n21618), .B2(n21640), .ZN(
        n21623) );
  OAI22_X1 U23265 ( .A1(n21621), .A2(n21648), .B1(n21646), .B2(n21620), .ZN(
        n21622) );
  AOI211_X1 U23266 ( .C1(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .C2(n21645), .A(
        n21623), .B(n21622), .ZN(n21624) );
  OAI21_X1 U23267 ( .B1(n11375), .B2(n21625), .A(n21624), .ZN(P1_U2816) );
  AOI22_X1 U23268 ( .A1(n21628), .A2(n21627), .B1(P1_EBX_REG_25__SCAN_IN), 
        .B2(n21626), .ZN(n21635) );
  AOI21_X1 U23269 ( .B1(P1_REIP_REG_25__SCAN_IN), .B2(n21639), .A(n11375), 
        .ZN(n21629) );
  OAI22_X1 U23270 ( .A1(n21630), .A2(n21648), .B1(n21638), .B2(n21629), .ZN(
        n21631) );
  AOI21_X1 U23271 ( .B1(n21633), .B2(n21632), .A(n21631), .ZN(n21634) );
  OAI211_X1 U23272 ( .C1(n21637), .C2(n21636), .A(n21635), .B(n21634), .ZN(
        P1_U2815) );
  AOI21_X1 U23273 ( .B1(P1_REIP_REG_26__SCAN_IN), .B2(n21639), .A(n21638), 
        .ZN(n21653) );
  OAI22_X1 U23274 ( .A1(n21643), .A2(n21642), .B1(n21641), .B2(n21640), .ZN(
        n21644) );
  AOI21_X1 U23275 ( .B1(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n21645), .A(
        n21644), .ZN(n21652) );
  OAI22_X1 U23276 ( .A1(n21649), .A2(n21648), .B1(n21647), .B2(n21646), .ZN(
        n21650) );
  INV_X1 U23277 ( .A(n21650), .ZN(n21651) );
  OAI211_X1 U23278 ( .C1(n21654), .C2(n21653), .A(n21652), .B(n21651), .ZN(
        P1_U2814) );
  OAI21_X1 U23279 ( .B1(n21657), .B2(n21656), .A(n21655), .ZN(P1_U2806) );
  AOI22_X1 U23280 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n21658), .B1(n11448), 
        .B2(n21683), .ZN(n21659) );
  OAI21_X1 U23281 ( .B1(n21660), .B2(n21666), .A(n21659), .ZN(n21662) );
  AOI22_X1 U23282 ( .A1(n21663), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n21662), .B2(n21661), .ZN(n21664) );
  OAI21_X1 U23283 ( .B1(n21666), .B2(n21665), .A(n21664), .ZN(P1_U3474) );
  NOR2_X1 U23284 ( .A1(n21668), .A2(n21667), .ZN(n21687) );
  OAI22_X1 U23285 ( .A1(n21671), .A2(n21915), .B1(n21670), .B2(n21669), .ZN(
        n21672) );
  OAI21_X1 U23286 ( .B1(n21687), .B2(n21672), .A(n21674), .ZN(n21673) );
  OAI21_X1 U23287 ( .B1(n21674), .B2(n21877), .A(n21673), .ZN(P1_U3478) );
  NAND2_X1 U23288 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n21675), .ZN(n21679) );
  NAND2_X1 U23289 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n21910), .ZN(n21678) );
  OAI211_X1 U23290 ( .C1(n21679), .C2(n21678), .A(n21677), .B(n21676), .ZN(
        P1_U3163) );
  OAI221_X1 U23291 ( .B1(n21868), .B2(P1_STATE2_REG_0__SCAN_IN), .C1(n21868), 
        .C2(n21681), .A(n21680), .ZN(P1_U3466) );
  INV_X1 U23292 ( .A(n21681), .ZN(n21682) );
  AOI21_X1 U23293 ( .B1(n21684), .B2(n21683), .A(n21682), .ZN(n21685) );
  OAI22_X1 U23294 ( .A1(n21687), .A2(n21686), .B1(P1_STATE2_REG_0__SCAN_IN), 
        .B2(n21685), .ZN(n21688) );
  OAI21_X1 U23295 ( .B1(n21690), .B2(n21689), .A(n21688), .ZN(P1_U3161) );
  AOI21_X1 U23296 ( .B1(n16736), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n21692), 
        .ZN(n21691) );
  INV_X1 U23297 ( .A(n21691), .ZN(P1_U2805) );
  AOI21_X1 U23298 ( .B1(n16736), .B2(P1_DATAWIDTH_REG_1__SCAN_IN), .A(n21692), 
        .ZN(n21693) );
  INV_X1 U23299 ( .A(n21693), .ZN(P1_U3465) );
  INV_X1 U23300 ( .A(n21694), .ZN(n21696) );
  OAI21_X1 U23301 ( .B1(n21698), .B2(n21695), .A(n21696), .ZN(P2_U2818) );
  OAI21_X1 U23302 ( .B1(n21698), .B2(n21697), .A(n21696), .ZN(P2_U3592) );
  INV_X1 U23303 ( .A(n21699), .ZN(n21701) );
  OAI21_X1 U23304 ( .B1(n21703), .B2(n21700), .A(n21701), .ZN(P3_U2636) );
  OAI21_X1 U23305 ( .B1(n21703), .B2(n21702), .A(n21701), .ZN(P3_U3281) );
  INV_X1 U23306 ( .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n21704) );
  AOI21_X1 U23307 ( .B1(HOLD), .B2(n21705), .A(n21704), .ZN(n21709) );
  AOI21_X1 U23308 ( .B1(n21707), .B2(P3_STATE_REG_1__SCAN_IN), .A(n21706), 
        .ZN(n21763) );
  OAI21_X1 U23309 ( .B1(P3_STATE_REG_1__SCAN_IN), .B2(n21759), .A(
        P3_STATE_REG_2__SCAN_IN), .ZN(n21762) );
  INV_X1 U23310 ( .A(n21762), .ZN(n21708) );
  OAI22_X1 U23311 ( .A1(n21710), .A2(n21709), .B1(n21763), .B2(n21708), .ZN(
        P3_U3029) );
  NAND2_X1 U23312 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(n21712), .ZN(n21719) );
  NAND2_X1 U23313 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n21719), .ZN(n21724) );
  OAI21_X1 U23314 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n21759), .A(n21724), 
        .ZN(n21717) );
  AOI21_X1 U23315 ( .B1(P1_STATE_REG_2__SCAN_IN), .B2(HOLD), .A(n21714), .ZN(
        n21722) );
  AOI21_X1 U23316 ( .B1(n21712), .B2(n21759), .A(n21711), .ZN(n21713) );
  OAI33_X1 U23317 ( .A1(n21714), .A2(NA), .A3(n21719), .B1(n21757), .B2(n21722), .B3(n21713), .ZN(n21715) );
  NAND2_X1 U23318 ( .A1(n21715), .A2(P1_STATE_REG_0__SCAN_IN), .ZN(n21716) );
  OAI21_X1 U23319 ( .B1(n21717), .B2(n21725), .A(n21716), .ZN(P1_U3196) );
  NAND2_X1 U23320 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(HOLD), .ZN(n21721) );
  AOI21_X1 U23321 ( .B1(P1_STATE_REG_0__SCAN_IN), .B2(n21722), .A(n21718), 
        .ZN(n21720) );
  OAI211_X1 U23322 ( .C1(P1_STATE_REG_2__SCAN_IN), .C2(n21721), .A(n21720), 
        .B(n21719), .ZN(P1_U3195) );
  OAI211_X1 U23323 ( .C1(P1_STATE_REG_0__SCAN_IN), .C2(n21759), .A(n21722), 
        .B(n21721), .ZN(n21723) );
  AOI22_X1 U23324 ( .A1(n21725), .A2(n21724), .B1(n22219), .B2(n21723), .ZN(
        n21726) );
  INV_X1 U23325 ( .A(n21726), .ZN(P1_U3194) );
  NAND2_X1 U23326 ( .A1(HOLD), .A2(n21727), .ZN(n21733) );
  NOR2_X1 U23327 ( .A1(n21729), .A2(n21728), .ZN(n21741) );
  NAND2_X1 U23328 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(
        P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n21738) );
  OAI21_X1 U23329 ( .B1(n21734), .B2(P2_REQUESTPENDING_REG_SCAN_IN), .A(
        P2_STATE_REG_2__SCAN_IN), .ZN(n21730) );
  OAI21_X1 U23330 ( .B1(n21741), .B2(n21738), .A(n21730), .ZN(n21732) );
  NAND2_X1 U23331 ( .A1(n21731), .A2(NA), .ZN(n21740) );
  OAI211_X1 U23332 ( .C1(n21734), .C2(n21733), .A(n21732), .B(n21740), .ZN(
        P2_U3209) );
  AOI211_X1 U23333 ( .C1(n21736), .C2(HOLD), .A(n21741), .B(n21735), .ZN(
        n21737) );
  OAI221_X1 U23334 ( .B1(n21738), .B2(HOLD), .C1(n21738), .C2(
        P2_STATE_REG_2__SCAN_IN), .A(n21737), .ZN(P2_U3210) );
  AOI221_X1 U23335 ( .B1(HOLD), .B2(n21740), .C1(n21739), .C2(n21740), .A(
        n21741), .ZN(n21746) );
  INV_X1 U23336 ( .A(n21741), .ZN(n21742) );
  OAI22_X1 U23337 ( .A1(NA), .A2(n21742), .B1(P2_STATE_REG_1__SCAN_IN), .B2(
        P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n21743) );
  OAI211_X1 U23338 ( .C1(HOLD), .C2(P2_REQUESTPENDING_REG_SCAN_IN), .A(
        P2_STATE_REG_0__SCAN_IN), .B(n21743), .ZN(n21744) );
  OAI21_X1 U23339 ( .B1(n21746), .B2(n21745), .A(n21744), .ZN(P2_U3211) );
  NOR2_X1 U23340 ( .A1(HOLD), .A2(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n21765)
         );
  OAI21_X1 U23341 ( .B1(n21758), .B2(n21757), .A(P3_STATE_REG_1__SCAN_IN), 
        .ZN(n21749) );
  NOR2_X1 U23342 ( .A1(n21755), .A2(n21747), .ZN(n21760) );
  INV_X1 U23343 ( .A(n21760), .ZN(n21748) );
  OAI21_X1 U23344 ( .B1(n21765), .B2(n21749), .A(n21748), .ZN(n21752) );
  OAI211_X1 U23345 ( .C1(n21758), .C2(n21757), .A(P3_STATE_REG_0__SCAN_IN), 
        .B(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n21750) );
  AOI21_X1 U23346 ( .B1(n21750), .B2(n21753), .A(P3_STATE_REG_1__SCAN_IN), 
        .ZN(n21751) );
  AOI21_X1 U23347 ( .B1(n21753), .B2(n21752), .A(n21751), .ZN(n21754) );
  OAI221_X1 U23348 ( .B1(n21756), .B2(P3_STATE_REG_2__SCAN_IN), .C1(n21756), 
        .C2(n21755), .A(n21754), .ZN(P3_U3030) );
  OAI22_X1 U23349 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(
        P3_REQUESTPENDING_REG_SCAN_IN), .B1(n21758), .B2(n21757), .ZN(n21761)
         );
  OAI221_X1 U23350 ( .B1(n21761), .B2(n21760), .C1(n21761), .C2(n21759), .A(
        P3_STATE_REG_0__SCAN_IN), .ZN(n21764) );
  OAI22_X1 U23351 ( .A1(n21765), .A2(n21764), .B1(n21763), .B2(n21762), .ZN(
        P3_U3031) );
  NAND2_X1 U23352 ( .A1(n22134), .A2(n21857), .ZN(n21767) );
  NAND2_X1 U23353 ( .A1(n21881), .A2(n14152), .ZN(n21840) );
  OAI21_X1 U23354 ( .B1(n22142), .B2(n21767), .A(n21840), .ZN(n21774) );
  OR2_X1 U23355 ( .A1(n21769), .A2(n21768), .ZN(n21789) );
  NOR2_X1 U23356 ( .A1(n21789), .A2(n21890), .ZN(n21772) );
  NAND3_X1 U23357 ( .A1(n12300), .A2(n11700), .A3(n21864), .ZN(n21780) );
  INV_X1 U23358 ( .A(n21780), .ZN(n21783) );
  NAND2_X1 U23359 ( .A1(n21877), .A2(n21783), .ZN(n22133) );
  INV_X1 U23360 ( .A(n22133), .ZN(n21770) );
  AOI22_X1 U23361 ( .A1(n22213), .A2(n21900), .B1(n21913), .B2(n21770), .ZN(
        n21778) );
  INV_X1 U23362 ( .A(n21772), .ZN(n21773) );
  AOI22_X1 U23363 ( .A1(n21774), .A2(n21773), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n22133), .ZN(n21775) );
  OAI211_X1 U23364 ( .C1(n21776), .C2(n21910), .A(n21852), .B(n21775), .ZN(
        n22136) );
  AOI22_X1 U23365 ( .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n22136), .B1(
        n22142), .B2(n21921), .ZN(n21777) );
  OAI211_X1 U23366 ( .C1(n22139), .C2(n21876), .A(n21778), .B(n21777), .ZN(
        P1_U3033) );
  INV_X1 U23367 ( .A(n21884), .ZN(n21779) );
  INV_X1 U23368 ( .A(n21789), .ZN(n21798) );
  NOR2_X1 U23369 ( .A1(n21877), .A2(n21780), .ZN(n22140) );
  AOI21_X1 U23370 ( .B1(n21798), .B2(n21878), .A(n22140), .ZN(n21781) );
  OAI22_X1 U23371 ( .A1(n21781), .A2(n21915), .B1(n21780), .B2(n21910), .ZN(
        n22141) );
  AOI22_X1 U23372 ( .A1(n22141), .A2(n21914), .B1(n21913), .B2(n22140), .ZN(
        n21785) );
  INV_X1 U23373 ( .A(n21787), .ZN(n21797) );
  OAI211_X1 U23374 ( .C1(n21797), .C2(n14152), .A(n21881), .B(n21781), .ZN(
        n21782) );
  OAI211_X1 U23375 ( .C1(n21857), .C2(n21783), .A(n21918), .B(n21782), .ZN(
        n22143) );
  AOI22_X1 U23376 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n22143), .B1(
        n22142), .B2(n21900), .ZN(n21784) );
  OAI211_X1 U23377 ( .C1(n21903), .C2(n22146), .A(n21785), .B(n21784), .ZN(
        P1_U3041) );
  NAND2_X1 U23378 ( .A1(n22146), .A2(n21857), .ZN(n21788) );
  INV_X1 U23379 ( .A(n21786), .ZN(n21888) );
  OAI21_X1 U23380 ( .B1(n21788), .B2(n22154), .A(n21840), .ZN(n21790) );
  NOR2_X1 U23381 ( .A1(n21789), .A2(n10973), .ZN(n21792) );
  NOR2_X1 U23382 ( .A1(n21823), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n21812) );
  NAND3_X1 U23383 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n12300), .A3(
        n11700), .ZN(n21801) );
  NOR2_X1 U23384 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21801), .ZN(
        n22147) );
  AOI22_X1 U23385 ( .A1(n22154), .A2(n21921), .B1(n21913), .B2(n22147), .ZN(
        n21795) );
  INV_X1 U23386 ( .A(n21790), .ZN(n21793) );
  INV_X1 U23387 ( .A(n22147), .ZN(n22068) );
  NOR2_X1 U23388 ( .A1(n21812), .A2(n21910), .ZN(n21815) );
  AOI21_X1 U23389 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n22068), .A(n21815), 
        .ZN(n21791) );
  INV_X1 U23390 ( .A(n22146), .ZN(n22148) );
  AOI22_X1 U23391 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n22149), .B1(
        n22148), .B2(n21900), .ZN(n21794) );
  OAI211_X1 U23392 ( .C1(n22152), .C2(n21876), .A(n21795), .B(n21794), .ZN(
        P1_U3049) );
  OAI21_X1 U23393 ( .B1(n21797), .B2(n21796), .A(n21857), .ZN(n21800) );
  NOR2_X1 U23394 ( .A1(n21877), .A2(n21801), .ZN(n22153) );
  AOI21_X1 U23395 ( .B1(n21798), .B2(n21904), .A(n22153), .ZN(n21804) );
  OAI22_X1 U23396 ( .A1(n21910), .A2(n21801), .B1(n21800), .B2(n21804), .ZN(
        n21799) );
  AOI22_X1 U23397 ( .A1(n22154), .A2(n21900), .B1(n21913), .B2(n22153), .ZN(
        n21808) );
  INV_X1 U23398 ( .A(n21800), .ZN(n21805) );
  INV_X1 U23399 ( .A(n21801), .ZN(n21802) );
  OAI21_X1 U23400 ( .B1(n21857), .B2(n21802), .A(n21918), .ZN(n21803) );
  AOI21_X1 U23401 ( .B1(n21805), .B2(n21804), .A(n21803), .ZN(n21806) );
  AOI22_X1 U23402 ( .A1(n22156), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n22155), .B2(n21921), .ZN(n21807) );
  OAI211_X1 U23403 ( .C1(n22159), .C2(n21876), .A(n21808), .B(n21807), .ZN(
        P1_U3057) );
  NOR3_X1 U23404 ( .A1(n22161), .A2(n22162), .A3(n21915), .ZN(n21810) );
  INV_X1 U23405 ( .A(n21840), .ZN(n21809) );
  NOR2_X1 U23406 ( .A1(n21810), .A2(n21809), .ZN(n21819) );
  INV_X1 U23407 ( .A(n21819), .ZN(n21813) );
  NOR2_X1 U23408 ( .A1(n21811), .A2(n10973), .ZN(n21818) );
  NOR3_X2 U23409 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A3(n21916), .ZN(n22160) );
  AOI22_X1 U23410 ( .A1(n22162), .A2(n21921), .B1(n21913), .B2(n22160), .ZN(
        n21821) );
  INV_X1 U23411 ( .A(n22160), .ZN(n21816) );
  AOI211_X1 U23412 ( .C1(n21816), .C2(P1_STATE2_REG_3__SCAN_IN), .A(n21815), 
        .B(n21814), .ZN(n21817) );
  OAI21_X1 U23413 ( .B1(n21819), .B2(n21818), .A(n21817), .ZN(n22163) );
  AOI22_X1 U23414 ( .A1(n22163), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n21900), .B2(n22161), .ZN(n21820) );
  OAI211_X1 U23415 ( .C1(n22166), .C2(n21876), .A(n21821), .B(n21820), .ZN(
        P1_U3081) );
  NAND3_X1 U23416 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n11700), .A3(
        n21864), .ZN(n21832) );
  NOR2_X1 U23417 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21832), .ZN(
        n22167) );
  AOI21_X1 U23418 ( .B1(n21842), .B2(n10973), .A(n22167), .ZN(n21827) );
  NAND2_X1 U23419 ( .A1(n21824), .A2(n21823), .ZN(n21870) );
  INV_X1 U23420 ( .A(n21845), .ZN(n21825) );
  OAI22_X1 U23421 ( .A1(n21827), .A2(n21915), .B1(n21870), .B2(n21825), .ZN(
        n22168) );
  AOI22_X1 U23422 ( .A1(n22168), .A2(n21914), .B1(n21913), .B2(n22167), .ZN(
        n21831) );
  INV_X1 U23423 ( .A(n22178), .ZN(n21826) );
  OAI21_X1 U23424 ( .B1(n21826), .B2(n22169), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n21828) );
  NAND2_X1 U23425 ( .A1(n21828), .A2(n21827), .ZN(n21829) );
  AOI22_X1 U23426 ( .A1(n22170), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n21900), .B2(n22169), .ZN(n21830) );
  OAI211_X1 U23427 ( .C1(n21903), .C2(n22178), .A(n21831), .B(n21830), .ZN(
        P1_U3097) );
  INV_X1 U23428 ( .A(n21900), .ZN(n21924) );
  NOR2_X1 U23429 ( .A1(n21877), .A2(n21832), .ZN(n22173) );
  AOI21_X1 U23430 ( .B1(n21842), .B2(n21878), .A(n22173), .ZN(n21833) );
  OAI22_X1 U23431 ( .A1(n21833), .A2(n21915), .B1(n21832), .B2(n21910), .ZN(
        n22174) );
  AOI22_X1 U23432 ( .A1(n22174), .A2(n21914), .B1(n21913), .B2(n22173), .ZN(
        n21838) );
  INV_X1 U23433 ( .A(n21832), .ZN(n21835) );
  OAI21_X1 U23434 ( .B1(n21836), .B2(n14152), .A(n21833), .ZN(n21834) );
  OAI221_X1 U23435 ( .B1(n21857), .B2(n21835), .C1(n21915), .C2(n21834), .A(
        n21918), .ZN(n22175) );
  AOI22_X1 U23436 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n22175), .B1(
        n22181), .B2(n21921), .ZN(n21837) );
  OAI211_X1 U23437 ( .C1(n21924), .C2(n22178), .A(n21838), .B(n21837), .ZN(
        P1_U3105) );
  INV_X1 U23438 ( .A(n22181), .ZN(n21839) );
  NAND2_X1 U23439 ( .A1(n21839), .A2(n21857), .ZN(n21841) );
  OAI21_X1 U23440 ( .B1(n21841), .B2(n22180), .A(n21840), .ZN(n21850) );
  AND2_X1 U23441 ( .A1(n21842), .A2(n21890), .ZN(n21847) );
  NAND2_X1 U23442 ( .A1(n21843), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n21892) );
  INV_X1 U23443 ( .A(n21892), .ZN(n21844) );
  NOR2_X1 U23444 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21846), .ZN(
        n22179) );
  AOI22_X1 U23445 ( .A1(n22180), .A2(n21921), .B1(n21913), .B2(n22179), .ZN(
        n21854) );
  INV_X1 U23446 ( .A(n21847), .ZN(n21849) );
  INV_X1 U23447 ( .A(n22179), .ZN(n21848) );
  AOI22_X1 U23448 ( .A1(n21850), .A2(n21849), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n21848), .ZN(n21851) );
  NAND2_X1 U23449 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n21892), .ZN(n21897) );
  NAND3_X1 U23450 ( .A1(n21852), .A2(n21851), .A3(n21897), .ZN(n22182) );
  AOI22_X1 U23451 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n22182), .B1(
        n22181), .B2(n21900), .ZN(n21853) );
  OAI211_X1 U23452 ( .C1(n22185), .C2(n21876), .A(n21854), .B(n21853), .ZN(
        P1_U3113) );
  INV_X1 U23453 ( .A(n22200), .ZN(n21856) );
  OAI21_X1 U23454 ( .B1(n22189), .B2(n21856), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n21858) );
  NAND2_X1 U23455 ( .A1(n21858), .A2(n21857), .ZN(n21873) );
  INV_X1 U23456 ( .A(n21873), .ZN(n21863) );
  OR2_X1 U23457 ( .A1(n21860), .A2(n21859), .ZN(n21908) );
  NOR2_X1 U23458 ( .A1(n21908), .A2(n21890), .ZN(n21872) );
  INV_X1 U23459 ( .A(n21870), .ZN(n21861) );
  NAND3_X1 U23460 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n21864), .ZN(n21879) );
  NOR2_X1 U23461 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21879), .ZN(
        n21867) );
  INV_X1 U23462 ( .A(n21867), .ZN(n22186) );
  OAI22_X1 U23463 ( .A1(n22200), .A2(n21903), .B1(n21865), .B2(n22186), .ZN(
        n21866) );
  INV_X1 U23464 ( .A(n21866), .ZN(n21875) );
  OAI21_X1 U23465 ( .B1(n21868), .B2(n21867), .A(n21898), .ZN(n21869) );
  AOI21_X1 U23466 ( .B1(n21870), .B2(P1_STATE2_REG_2__SCAN_IN), .A(n21869), 
        .ZN(n21871) );
  AOI22_X1 U23467 ( .A1(n22190), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n21900), .B2(n22189), .ZN(n21874) );
  OAI211_X1 U23468 ( .C1(n22194), .C2(n21876), .A(n21875), .B(n21874), .ZN(
        P1_U3129) );
  INV_X1 U23469 ( .A(n21908), .ZN(n21891) );
  NOR2_X1 U23470 ( .A1(n21877), .A2(n21879), .ZN(n22195) );
  AOI21_X1 U23471 ( .B1(n21891), .B2(n21878), .A(n22195), .ZN(n21880) );
  OAI22_X1 U23472 ( .A1(n21880), .A2(n21915), .B1(n21879), .B2(n21910), .ZN(
        n22196) );
  AOI22_X1 U23473 ( .A1(n22196), .A2(n21914), .B1(n21913), .B2(n22195), .ZN(
        n21887) );
  INV_X1 U23474 ( .A(n21879), .ZN(n21883) );
  OAI211_X1 U23475 ( .C1(n21885), .C2(n14152), .A(n21881), .B(n21880), .ZN(
        n21882) );
  OAI211_X1 U23476 ( .C1(n21857), .C2(n21883), .A(n21918), .B(n21882), .ZN(
        n22197) );
  AOI22_X1 U23477 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n22197), .B1(
        n22204), .B2(n21921), .ZN(n21886) );
  OAI211_X1 U23478 ( .C1(n21924), .C2(n22200), .A(n21887), .B(n21886), .ZN(
        P1_U3137) );
  NAND2_X1 U23479 ( .A1(n21891), .A2(n21890), .ZN(n21895) );
  OAI22_X1 U23480 ( .A1(n21895), .A2(n21915), .B1(n21893), .B2(n21892), .ZN(
        n22202) );
  NOR3_X2 U23481 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n12300), .A3(
        n21916), .ZN(n22201) );
  AOI22_X1 U23482 ( .A1(n21914), .A2(n22202), .B1(n21913), .B2(n22201), .ZN(
        n21902) );
  INV_X1 U23483 ( .A(n22218), .ZN(n21894) );
  OAI21_X1 U23484 ( .B1(n21894), .B2(n22204), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n21896) );
  AOI21_X1 U23485 ( .B1(n21896), .B2(n21895), .A(P1_STATE2_REG_3__SCAN_IN), 
        .ZN(n21899) );
  AOI22_X1 U23486 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n22205), .B1(
        n22204), .B2(n21900), .ZN(n21901) );
  OAI211_X1 U23487 ( .C1(n21903), .C2(n22218), .A(n21902), .B(n21901), .ZN(
        P1_U3145) );
  INV_X1 U23488 ( .A(n21904), .ZN(n21907) );
  NOR2_X1 U23489 ( .A1(n12300), .A2(n21905), .ZN(n22209) );
  INV_X1 U23490 ( .A(n22209), .ZN(n21906) );
  OAI21_X1 U23491 ( .B1(n21908), .B2(n21907), .A(n21906), .ZN(n21919) );
  INV_X1 U23492 ( .A(n21919), .ZN(n21912) );
  NAND2_X1 U23493 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n21909), .ZN(
        n21911) );
  OAI22_X1 U23494 ( .A1(n21912), .A2(n21915), .B1(n21911), .B2(n21910), .ZN(
        n22212) );
  AOI22_X1 U23495 ( .A1(n22212), .A2(n21914), .B1(n21913), .B2(n22209), .ZN(
        n21923) );
  OAI21_X1 U23496 ( .B1(n21916), .B2(n12300), .A(n21915), .ZN(n21917) );
  OAI211_X1 U23497 ( .C1(n21920), .C2(n21919), .A(n21918), .B(n21917), .ZN(
        n22215) );
  AOI22_X1 U23498 ( .A1(n22215), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n21921), .B2(n22213), .ZN(n21922) );
  OAI211_X1 U23499 ( .C1(n21924), .C2(n22218), .A(n21923), .B(n21922), .ZN(
        P1_U3153) );
  OAI22_X1 U23500 ( .A1(n22134), .A2(n21958), .B1(n21942), .B2(n22133), .ZN(
        n21925) );
  INV_X1 U23501 ( .A(n21925), .ZN(n21927) );
  AOI22_X1 U23502 ( .A1(P1_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n22136), .B1(
        n22142), .B2(n21955), .ZN(n21926) );
  OAI211_X1 U23503 ( .C1(n22139), .C2(n21946), .A(n21927), .B(n21926), .ZN(
        P1_U3034) );
  AOI22_X1 U23504 ( .A1(n22141), .A2(n21954), .B1(n21953), .B2(n22140), .ZN(
        n21929) );
  AOI22_X1 U23505 ( .A1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n22143), .B1(
        n22142), .B2(n21949), .ZN(n21928) );
  OAI211_X1 U23506 ( .C1(n21952), .C2(n22146), .A(n21929), .B(n21928), .ZN(
        P1_U3042) );
  AOI22_X1 U23507 ( .A1(n22154), .A2(n21955), .B1(n21953), .B2(n22147), .ZN(
        n21931) );
  AOI22_X1 U23508 ( .A1(P1_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n22149), .B1(
        n22148), .B2(n21949), .ZN(n21930) );
  OAI211_X1 U23509 ( .C1(n22152), .C2(n21946), .A(n21931), .B(n21930), .ZN(
        P1_U3050) );
  AOI22_X1 U23510 ( .A1(n22155), .A2(n21955), .B1(n21953), .B2(n22153), .ZN(
        n21933) );
  AOI22_X1 U23511 ( .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n22156), .B1(
        n22154), .B2(n21949), .ZN(n21932) );
  OAI211_X1 U23512 ( .C1(n22159), .C2(n21946), .A(n21933), .B(n21932), .ZN(
        P1_U3058) );
  AOI22_X1 U23513 ( .A1(n22162), .A2(n21955), .B1(n21953), .B2(n22160), .ZN(
        n21935) );
  AOI22_X1 U23514 ( .A1(n22163), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n21949), .B2(n22161), .ZN(n21934) );
  OAI211_X1 U23515 ( .C1(n22166), .C2(n21946), .A(n21935), .B(n21934), .ZN(
        P1_U3082) );
  AOI22_X1 U23516 ( .A1(n22168), .A2(n21954), .B1(n21953), .B2(n22167), .ZN(
        n21937) );
  AOI22_X1 U23517 ( .A1(n22170), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n21949), .B2(n22169), .ZN(n21936) );
  OAI211_X1 U23518 ( .C1(n21952), .C2(n22178), .A(n21937), .B(n21936), .ZN(
        P1_U3098) );
  AOI22_X1 U23519 ( .A1(n22174), .A2(n21954), .B1(n21953), .B2(n22173), .ZN(
        n21939) );
  AOI22_X1 U23520 ( .A1(P1_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n22175), .B1(
        n22181), .B2(n21955), .ZN(n21938) );
  OAI211_X1 U23521 ( .C1(n21958), .C2(n22178), .A(n21939), .B(n21938), .ZN(
        P1_U3106) );
  AOI22_X1 U23522 ( .A1(n22180), .A2(n21955), .B1(n21953), .B2(n22179), .ZN(
        n21941) );
  AOI22_X1 U23523 ( .A1(P1_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n22182), .B1(
        n22181), .B2(n21949), .ZN(n21940) );
  OAI211_X1 U23524 ( .C1(n22185), .C2(n21946), .A(n21941), .B(n21940), .ZN(
        P1_U3114) );
  OAI22_X1 U23525 ( .A1(n22200), .A2(n21952), .B1(n21942), .B2(n22186), .ZN(
        n21943) );
  INV_X1 U23526 ( .A(n21943), .ZN(n21945) );
  AOI22_X1 U23527 ( .A1(n22190), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n21949), .B2(n22189), .ZN(n21944) );
  OAI211_X1 U23528 ( .C1(n22194), .C2(n21946), .A(n21945), .B(n21944), .ZN(
        P1_U3130) );
  AOI22_X1 U23529 ( .A1(n22196), .A2(n21954), .B1(n21953), .B2(n22195), .ZN(
        n21948) );
  AOI22_X1 U23530 ( .A1(P1_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n22197), .B1(
        n22204), .B2(n21955), .ZN(n21947) );
  OAI211_X1 U23531 ( .C1(n21958), .C2(n22200), .A(n21948), .B(n21947), .ZN(
        P1_U3138) );
  AOI22_X1 U23532 ( .A1(n21954), .A2(n22202), .B1(n21953), .B2(n22201), .ZN(
        n21951) );
  AOI22_X1 U23533 ( .A1(P1_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n22205), .B1(
        n22204), .B2(n21949), .ZN(n21950) );
  OAI211_X1 U23534 ( .C1(n21952), .C2(n22218), .A(n21951), .B(n21950), .ZN(
        P1_U3146) );
  AOI22_X1 U23535 ( .A1(n22212), .A2(n21954), .B1(n21953), .B2(n22209), .ZN(
        n21957) );
  AOI22_X1 U23536 ( .A1(n22215), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n21955), .B2(n22213), .ZN(n21956) );
  OAI211_X1 U23537 ( .C1(n21958), .C2(n22218), .A(n21957), .B(n21956), .ZN(
        P1_U3154) );
  OAI22_X1 U23538 ( .A1(n22134), .A2(n21993), .B1(n21977), .B2(n22133), .ZN(
        n21959) );
  INV_X1 U23539 ( .A(n21959), .ZN(n21961) );
  AOI22_X1 U23540 ( .A1(P1_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n22136), .B1(
        n22142), .B2(n21990), .ZN(n21960) );
  OAI211_X1 U23541 ( .C1(n22139), .C2(n21981), .A(n21961), .B(n21960), .ZN(
        P1_U3035) );
  AOI22_X1 U23542 ( .A1(n22141), .A2(n21989), .B1(n21988), .B2(n22140), .ZN(
        n21963) );
  AOI22_X1 U23543 ( .A1(P1_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n22143), .B1(
        n22142), .B2(n21984), .ZN(n21962) );
  OAI211_X1 U23544 ( .C1(n21987), .C2(n22146), .A(n21963), .B(n21962), .ZN(
        P1_U3043) );
  OAI22_X1 U23545 ( .A1(n22146), .A2(n21993), .B1(n21977), .B2(n22068), .ZN(
        n21964) );
  INV_X1 U23546 ( .A(n21964), .ZN(n21966) );
  AOI22_X1 U23547 ( .A1(P1_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n22149), .B1(
        n22154), .B2(n21990), .ZN(n21965) );
  OAI211_X1 U23548 ( .C1(n22152), .C2(n21981), .A(n21966), .B(n21965), .ZN(
        P1_U3051) );
  AOI22_X1 U23549 ( .A1(n22154), .A2(n21984), .B1(n21988), .B2(n22153), .ZN(
        n21968) );
  AOI22_X1 U23550 ( .A1(n22156), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n22155), .B2(n21990), .ZN(n21967) );
  OAI211_X1 U23551 ( .C1(n22159), .C2(n21981), .A(n21968), .B(n21967), .ZN(
        P1_U3059) );
  AOI22_X1 U23552 ( .A1(n22162), .A2(n21990), .B1(n21988), .B2(n22160), .ZN(
        n21970) );
  AOI22_X1 U23553 ( .A1(n22163), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n21984), .B2(n22161), .ZN(n21969) );
  OAI211_X1 U23554 ( .C1(n22166), .C2(n21981), .A(n21970), .B(n21969), .ZN(
        P1_U3083) );
  AOI22_X1 U23555 ( .A1(n22168), .A2(n21989), .B1(n21988), .B2(n22167), .ZN(
        n21972) );
  AOI22_X1 U23556 ( .A1(n22170), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n21984), .B2(n22169), .ZN(n21971) );
  OAI211_X1 U23557 ( .C1(n21987), .C2(n22178), .A(n21972), .B(n21971), .ZN(
        P1_U3099) );
  AOI22_X1 U23558 ( .A1(n22174), .A2(n21989), .B1(n21988), .B2(n22173), .ZN(
        n21974) );
  AOI22_X1 U23559 ( .A1(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n22175), .B1(
        n22181), .B2(n21990), .ZN(n21973) );
  OAI211_X1 U23560 ( .C1(n21993), .C2(n22178), .A(n21974), .B(n21973), .ZN(
        P1_U3107) );
  AOI22_X1 U23561 ( .A1(n22181), .A2(n21984), .B1(n21988), .B2(n22179), .ZN(
        n21976) );
  AOI22_X1 U23562 ( .A1(P1_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n22182), .B1(
        n22180), .B2(n21990), .ZN(n21975) );
  OAI211_X1 U23563 ( .C1(n22185), .C2(n21981), .A(n21976), .B(n21975), .ZN(
        P1_U3115) );
  OAI22_X1 U23564 ( .A1(n22200), .A2(n21987), .B1(n21977), .B2(n22186), .ZN(
        n21978) );
  INV_X1 U23565 ( .A(n21978), .ZN(n21980) );
  AOI22_X1 U23566 ( .A1(n22190), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n21984), .B2(n22189), .ZN(n21979) );
  OAI211_X1 U23567 ( .C1(n22194), .C2(n21981), .A(n21980), .B(n21979), .ZN(
        P1_U3131) );
  AOI22_X1 U23568 ( .A1(n22196), .A2(n21989), .B1(n21988), .B2(n22195), .ZN(
        n21983) );
  AOI22_X1 U23569 ( .A1(P1_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n22197), .B1(
        n22204), .B2(n21990), .ZN(n21982) );
  OAI211_X1 U23570 ( .C1(n21993), .C2(n22200), .A(n21983), .B(n21982), .ZN(
        P1_U3139) );
  AOI22_X1 U23571 ( .A1(n21989), .A2(n22202), .B1(n21988), .B2(n22201), .ZN(
        n21986) );
  AOI22_X1 U23572 ( .A1(P1_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n22205), .B1(
        n22204), .B2(n21984), .ZN(n21985) );
  OAI211_X1 U23573 ( .C1(n21987), .C2(n22218), .A(n21986), .B(n21985), .ZN(
        P1_U3147) );
  AOI22_X1 U23574 ( .A1(n22212), .A2(n21989), .B1(n21988), .B2(n22209), .ZN(
        n21992) );
  AOI22_X1 U23575 ( .A1(n22215), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n21990), .B2(n22213), .ZN(n21991) );
  OAI211_X1 U23576 ( .C1(n21993), .C2(n22218), .A(n21992), .B(n21991), .ZN(
        P1_U3155) );
  OAI22_X1 U23577 ( .A1(n22134), .A2(n22027), .B1(n22011), .B2(n22133), .ZN(
        n21994) );
  INV_X1 U23578 ( .A(n21994), .ZN(n21996) );
  AOI22_X1 U23579 ( .A1(P1_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n22136), .B1(
        n22142), .B2(n22024), .ZN(n21995) );
  OAI211_X1 U23580 ( .C1(n22139), .C2(n22015), .A(n21996), .B(n21995), .ZN(
        P1_U3036) );
  AOI22_X1 U23581 ( .A1(n22141), .A2(n22023), .B1(n22022), .B2(n22140), .ZN(
        n21998) );
  AOI22_X1 U23582 ( .A1(P1_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n22143), .B1(
        n22142), .B2(n22018), .ZN(n21997) );
  OAI211_X1 U23583 ( .C1(n22021), .C2(n22146), .A(n21998), .B(n21997), .ZN(
        P1_U3044) );
  AOI22_X1 U23584 ( .A1(n22154), .A2(n22024), .B1(n22022), .B2(n22147), .ZN(
        n22000) );
  AOI22_X1 U23585 ( .A1(P1_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n22149), .B1(
        n22148), .B2(n22018), .ZN(n21999) );
  OAI211_X1 U23586 ( .C1(n22152), .C2(n22015), .A(n22000), .B(n21999), .ZN(
        P1_U3052) );
  AOI22_X1 U23587 ( .A1(n22154), .A2(n22018), .B1(n22022), .B2(n22153), .ZN(
        n22002) );
  AOI22_X1 U23588 ( .A1(n22156), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n22155), .B2(n22024), .ZN(n22001) );
  OAI211_X1 U23589 ( .C1(n22159), .C2(n22015), .A(n22002), .B(n22001), .ZN(
        P1_U3060) );
  AOI22_X1 U23590 ( .A1(n22161), .A2(n22018), .B1(n22022), .B2(n22160), .ZN(
        n22004) );
  AOI22_X1 U23591 ( .A1(n22163), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n22024), .B2(n22162), .ZN(n22003) );
  OAI211_X1 U23592 ( .C1(n22166), .C2(n22015), .A(n22004), .B(n22003), .ZN(
        P1_U3084) );
  AOI22_X1 U23593 ( .A1(n22168), .A2(n22023), .B1(n22022), .B2(n22167), .ZN(
        n22006) );
  AOI22_X1 U23594 ( .A1(n22170), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n22018), .B2(n22169), .ZN(n22005) );
  OAI211_X1 U23595 ( .C1(n22021), .C2(n22178), .A(n22006), .B(n22005), .ZN(
        P1_U3100) );
  AOI22_X1 U23596 ( .A1(n22174), .A2(n22023), .B1(n22022), .B2(n22173), .ZN(
        n22008) );
  AOI22_X1 U23597 ( .A1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n22175), .B1(
        n22181), .B2(n22024), .ZN(n22007) );
  OAI211_X1 U23598 ( .C1(n22027), .C2(n22178), .A(n22008), .B(n22007), .ZN(
        P1_U3108) );
  AOI22_X1 U23599 ( .A1(n22181), .A2(n22018), .B1(n22022), .B2(n22179), .ZN(
        n22010) );
  AOI22_X1 U23600 ( .A1(P1_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n22182), .B1(
        n22180), .B2(n22024), .ZN(n22009) );
  OAI211_X1 U23601 ( .C1(n22185), .C2(n22015), .A(n22010), .B(n22009), .ZN(
        P1_U3116) );
  OAI22_X1 U23602 ( .A1(n22200), .A2(n22021), .B1(n22011), .B2(n22186), .ZN(
        n22012) );
  INV_X1 U23603 ( .A(n22012), .ZN(n22014) );
  AOI22_X1 U23604 ( .A1(n22190), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n22018), .B2(n22189), .ZN(n22013) );
  OAI211_X1 U23605 ( .C1(n22194), .C2(n22015), .A(n22014), .B(n22013), .ZN(
        P1_U3132) );
  AOI22_X1 U23606 ( .A1(n22196), .A2(n22023), .B1(n22022), .B2(n22195), .ZN(
        n22017) );
  AOI22_X1 U23607 ( .A1(P1_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n22197), .B1(
        n22204), .B2(n22024), .ZN(n22016) );
  OAI211_X1 U23608 ( .C1(n22027), .C2(n22200), .A(n22017), .B(n22016), .ZN(
        P1_U3140) );
  AOI22_X1 U23609 ( .A1(n22023), .A2(n22202), .B1(n22022), .B2(n22201), .ZN(
        n22020) );
  AOI22_X1 U23610 ( .A1(P1_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n22205), .B1(
        n22204), .B2(n22018), .ZN(n22019) );
  OAI211_X1 U23611 ( .C1(n22021), .C2(n22218), .A(n22020), .B(n22019), .ZN(
        P1_U3148) );
  AOI22_X1 U23612 ( .A1(n22212), .A2(n22023), .B1(n22022), .B2(n22209), .ZN(
        n22026) );
  AOI22_X1 U23613 ( .A1(n22215), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n22024), .B2(n22213), .ZN(n22025) );
  OAI211_X1 U23614 ( .C1(n22027), .C2(n22218), .A(n22026), .B(n22025), .ZN(
        P1_U3156) );
  OAI22_X1 U23615 ( .A1(n22134), .A2(n22062), .B1(n22046), .B2(n22133), .ZN(
        n22028) );
  INV_X1 U23616 ( .A(n22028), .ZN(n22030) );
  AOI22_X1 U23617 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n22136), .B1(
        n22142), .B2(n22059), .ZN(n22029) );
  OAI211_X1 U23618 ( .C1(n22139), .C2(n22050), .A(n22030), .B(n22029), .ZN(
        P1_U3037) );
  AOI22_X1 U23619 ( .A1(n22141), .A2(n22058), .B1(n22057), .B2(n22140), .ZN(
        n22032) );
  AOI22_X1 U23620 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n22143), .B1(
        n22142), .B2(n22053), .ZN(n22031) );
  OAI211_X1 U23621 ( .C1(n22056), .C2(n22146), .A(n22032), .B(n22031), .ZN(
        P1_U3045) );
  OAI22_X1 U23622 ( .A1(n22146), .A2(n22062), .B1(n22046), .B2(n22068), .ZN(
        n22033) );
  INV_X1 U23623 ( .A(n22033), .ZN(n22035) );
  AOI22_X1 U23624 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n22149), .B1(
        n22154), .B2(n22059), .ZN(n22034) );
  OAI211_X1 U23625 ( .C1(n22152), .C2(n22050), .A(n22035), .B(n22034), .ZN(
        P1_U3053) );
  AOI22_X1 U23626 ( .A1(n22155), .A2(n22059), .B1(n22057), .B2(n22153), .ZN(
        n22037) );
  AOI22_X1 U23627 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n22156), .B1(
        n22154), .B2(n22053), .ZN(n22036) );
  OAI211_X1 U23628 ( .C1(n22159), .C2(n22050), .A(n22037), .B(n22036), .ZN(
        P1_U3061) );
  AOI22_X1 U23629 ( .A1(n22161), .A2(n22053), .B1(n22057), .B2(n22160), .ZN(
        n22039) );
  AOI22_X1 U23630 ( .A1(n22163), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n22059), .B2(n22162), .ZN(n22038) );
  OAI211_X1 U23631 ( .C1(n22166), .C2(n22050), .A(n22039), .B(n22038), .ZN(
        P1_U3085) );
  AOI22_X1 U23632 ( .A1(n22168), .A2(n22058), .B1(n22057), .B2(n22167), .ZN(
        n22041) );
  AOI22_X1 U23633 ( .A1(n22170), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n22053), .B2(n22169), .ZN(n22040) );
  OAI211_X1 U23634 ( .C1(n22056), .C2(n22178), .A(n22041), .B(n22040), .ZN(
        P1_U3101) );
  AOI22_X1 U23635 ( .A1(n22174), .A2(n22058), .B1(n22057), .B2(n22173), .ZN(
        n22043) );
  AOI22_X1 U23636 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n22175), .B1(
        n22181), .B2(n22059), .ZN(n22042) );
  OAI211_X1 U23637 ( .C1(n22062), .C2(n22178), .A(n22043), .B(n22042), .ZN(
        P1_U3109) );
  AOI22_X1 U23638 ( .A1(n22181), .A2(n22053), .B1(n22057), .B2(n22179), .ZN(
        n22045) );
  AOI22_X1 U23639 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n22182), .B1(
        n22180), .B2(n22059), .ZN(n22044) );
  OAI211_X1 U23640 ( .C1(n22185), .C2(n22050), .A(n22045), .B(n22044), .ZN(
        P1_U3117) );
  OAI22_X1 U23641 ( .A1(n22200), .A2(n22056), .B1(n22046), .B2(n22186), .ZN(
        n22047) );
  INV_X1 U23642 ( .A(n22047), .ZN(n22049) );
  AOI22_X1 U23643 ( .A1(n22190), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n22053), .B2(n22189), .ZN(n22048) );
  OAI211_X1 U23644 ( .C1(n22194), .C2(n22050), .A(n22049), .B(n22048), .ZN(
        P1_U3133) );
  AOI22_X1 U23645 ( .A1(n22196), .A2(n22058), .B1(n22057), .B2(n22195), .ZN(
        n22052) );
  AOI22_X1 U23646 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n22197), .B1(
        n22204), .B2(n22059), .ZN(n22051) );
  OAI211_X1 U23647 ( .C1(n22062), .C2(n22200), .A(n22052), .B(n22051), .ZN(
        P1_U3141) );
  AOI22_X1 U23648 ( .A1(n22058), .A2(n22202), .B1(n22057), .B2(n22201), .ZN(
        n22055) );
  AOI22_X1 U23649 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n22205), .B1(
        n22204), .B2(n22053), .ZN(n22054) );
  OAI211_X1 U23650 ( .C1(n22056), .C2(n22218), .A(n22055), .B(n22054), .ZN(
        P1_U3149) );
  AOI22_X1 U23651 ( .A1(n22212), .A2(n22058), .B1(n22057), .B2(n22209), .ZN(
        n22061) );
  AOI22_X1 U23652 ( .A1(n22215), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n22059), .B2(n22213), .ZN(n22060) );
  OAI211_X1 U23653 ( .C1(n22062), .C2(n22218), .A(n22061), .B(n22060), .ZN(
        P1_U3157) );
  OAI22_X1 U23654 ( .A1(n22134), .A2(n22098), .B1(n22082), .B2(n22133), .ZN(
        n22063) );
  INV_X1 U23655 ( .A(n22063), .ZN(n22065) );
  AOI22_X1 U23656 ( .A1(P1_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n22136), .B1(
        n22142), .B2(n22095), .ZN(n22064) );
  OAI211_X1 U23657 ( .C1(n22139), .C2(n22086), .A(n22065), .B(n22064), .ZN(
        P1_U3038) );
  AOI22_X1 U23658 ( .A1(n22141), .A2(n22094), .B1(n22093), .B2(n22140), .ZN(
        n22067) );
  AOI22_X1 U23659 ( .A1(P1_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n22143), .B1(
        n22142), .B2(n22089), .ZN(n22066) );
  OAI211_X1 U23660 ( .C1(n22092), .C2(n22146), .A(n22067), .B(n22066), .ZN(
        P1_U3046) );
  OAI22_X1 U23661 ( .A1(n22146), .A2(n22098), .B1(n22082), .B2(n22068), .ZN(
        n22069) );
  INV_X1 U23662 ( .A(n22069), .ZN(n22071) );
  AOI22_X1 U23663 ( .A1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n22149), .B1(
        n22154), .B2(n22095), .ZN(n22070) );
  OAI211_X1 U23664 ( .C1(n22152), .C2(n22086), .A(n22071), .B(n22070), .ZN(
        P1_U3054) );
  AOI22_X1 U23665 ( .A1(n22154), .A2(n22089), .B1(n22093), .B2(n22153), .ZN(
        n22073) );
  AOI22_X1 U23666 ( .A1(n22156), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n22155), .B2(n22095), .ZN(n22072) );
  OAI211_X1 U23667 ( .C1(n22159), .C2(n22086), .A(n22073), .B(n22072), .ZN(
        P1_U3062) );
  AOI22_X1 U23668 ( .A1(n22161), .A2(n22089), .B1(n22093), .B2(n22160), .ZN(
        n22075) );
  AOI22_X1 U23669 ( .A1(n22163), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n22095), .B2(n22162), .ZN(n22074) );
  OAI211_X1 U23670 ( .C1(n22166), .C2(n22086), .A(n22075), .B(n22074), .ZN(
        P1_U3086) );
  AOI22_X1 U23671 ( .A1(n22168), .A2(n22094), .B1(n22093), .B2(n22167), .ZN(
        n22077) );
  AOI22_X1 U23672 ( .A1(n22170), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n22089), .B2(n22169), .ZN(n22076) );
  OAI211_X1 U23673 ( .C1(n22092), .C2(n22178), .A(n22077), .B(n22076), .ZN(
        P1_U3102) );
  AOI22_X1 U23674 ( .A1(n22174), .A2(n22094), .B1(n22093), .B2(n22173), .ZN(
        n22079) );
  AOI22_X1 U23675 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n22175), .B1(
        n22181), .B2(n22095), .ZN(n22078) );
  OAI211_X1 U23676 ( .C1(n22098), .C2(n22178), .A(n22079), .B(n22078), .ZN(
        P1_U3110) );
  AOI22_X1 U23677 ( .A1(n22181), .A2(n22089), .B1(n22093), .B2(n22179), .ZN(
        n22081) );
  AOI22_X1 U23678 ( .A1(P1_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n22182), .B1(
        n22180), .B2(n22095), .ZN(n22080) );
  OAI211_X1 U23679 ( .C1(n22185), .C2(n22086), .A(n22081), .B(n22080), .ZN(
        P1_U3118) );
  OAI22_X1 U23680 ( .A1(n22200), .A2(n22092), .B1(n22082), .B2(n22186), .ZN(
        n22083) );
  INV_X1 U23681 ( .A(n22083), .ZN(n22085) );
  AOI22_X1 U23682 ( .A1(n22190), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n22089), .B2(n22189), .ZN(n22084) );
  OAI211_X1 U23683 ( .C1(n22194), .C2(n22086), .A(n22085), .B(n22084), .ZN(
        P1_U3134) );
  AOI22_X1 U23684 ( .A1(n22196), .A2(n22094), .B1(n22093), .B2(n22195), .ZN(
        n22088) );
  AOI22_X1 U23685 ( .A1(P1_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n22197), .B1(
        n22204), .B2(n22095), .ZN(n22087) );
  OAI211_X1 U23686 ( .C1(n22098), .C2(n22200), .A(n22088), .B(n22087), .ZN(
        P1_U3142) );
  AOI22_X1 U23687 ( .A1(n22094), .A2(n22202), .B1(n22093), .B2(n22201), .ZN(
        n22091) );
  AOI22_X1 U23688 ( .A1(P1_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n22205), .B1(
        n22204), .B2(n22089), .ZN(n22090) );
  OAI211_X1 U23689 ( .C1(n22092), .C2(n22218), .A(n22091), .B(n22090), .ZN(
        P1_U3150) );
  AOI22_X1 U23690 ( .A1(n22212), .A2(n22094), .B1(n22093), .B2(n22209), .ZN(
        n22097) );
  AOI22_X1 U23691 ( .A1(n22215), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n22095), .B2(n22213), .ZN(n22096) );
  OAI211_X1 U23692 ( .C1(n22098), .C2(n22218), .A(n22097), .B(n22096), .ZN(
        P1_U3158) );
  OAI22_X1 U23693 ( .A1(n22134), .A2(n22132), .B1(n22116), .B2(n22133), .ZN(
        n22099) );
  INV_X1 U23694 ( .A(n22099), .ZN(n22101) );
  AOI22_X1 U23695 ( .A1(P1_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n22136), .B1(
        n22142), .B2(n22129), .ZN(n22100) );
  OAI211_X1 U23696 ( .C1(n22139), .C2(n22120), .A(n22101), .B(n22100), .ZN(
        P1_U3039) );
  AOI22_X1 U23697 ( .A1(n22141), .A2(n22128), .B1(n22127), .B2(n22140), .ZN(
        n22103) );
  AOI22_X1 U23698 ( .A1(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n22143), .B1(
        n22142), .B2(n22123), .ZN(n22102) );
  OAI211_X1 U23699 ( .C1(n22126), .C2(n22146), .A(n22103), .B(n22102), .ZN(
        P1_U3047) );
  AOI22_X1 U23700 ( .A1(n22154), .A2(n22129), .B1(n22127), .B2(n22147), .ZN(
        n22105) );
  AOI22_X1 U23701 ( .A1(P1_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n22149), .B1(
        n22148), .B2(n22123), .ZN(n22104) );
  OAI211_X1 U23702 ( .C1(n22152), .C2(n22120), .A(n22105), .B(n22104), .ZN(
        P1_U3055) );
  AOI22_X1 U23703 ( .A1(n22154), .A2(n22123), .B1(n22127), .B2(n22153), .ZN(
        n22107) );
  AOI22_X1 U23704 ( .A1(n22156), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n22155), .B2(n22129), .ZN(n22106) );
  OAI211_X1 U23705 ( .C1(n22159), .C2(n22120), .A(n22107), .B(n22106), .ZN(
        P1_U3063) );
  AOI22_X1 U23706 ( .A1(n22161), .A2(n22123), .B1(n22127), .B2(n22160), .ZN(
        n22109) );
  AOI22_X1 U23707 ( .A1(n22163), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n22129), .B2(n22162), .ZN(n22108) );
  OAI211_X1 U23708 ( .C1(n22166), .C2(n22120), .A(n22109), .B(n22108), .ZN(
        P1_U3087) );
  AOI22_X1 U23709 ( .A1(n22168), .A2(n22128), .B1(n22127), .B2(n22167), .ZN(
        n22111) );
  AOI22_X1 U23710 ( .A1(n22170), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n22123), .B2(n22169), .ZN(n22110) );
  OAI211_X1 U23711 ( .C1(n22126), .C2(n22178), .A(n22111), .B(n22110), .ZN(
        P1_U3103) );
  AOI22_X1 U23712 ( .A1(n22174), .A2(n22128), .B1(n22127), .B2(n22173), .ZN(
        n22113) );
  AOI22_X1 U23713 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n22175), .B1(
        n22181), .B2(n22129), .ZN(n22112) );
  OAI211_X1 U23714 ( .C1(n22132), .C2(n22178), .A(n22113), .B(n22112), .ZN(
        P1_U3111) );
  AOI22_X1 U23715 ( .A1(n22181), .A2(n22123), .B1(n22127), .B2(n22179), .ZN(
        n22115) );
  AOI22_X1 U23716 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n22182), .B1(
        n22180), .B2(n22129), .ZN(n22114) );
  OAI211_X1 U23717 ( .C1(n22185), .C2(n22120), .A(n22115), .B(n22114), .ZN(
        P1_U3119) );
  OAI22_X1 U23718 ( .A1(n22200), .A2(n22126), .B1(n22116), .B2(n22186), .ZN(
        n22117) );
  INV_X1 U23719 ( .A(n22117), .ZN(n22119) );
  AOI22_X1 U23720 ( .A1(n22190), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n22123), .B2(n22189), .ZN(n22118) );
  OAI211_X1 U23721 ( .C1(n22194), .C2(n22120), .A(n22119), .B(n22118), .ZN(
        P1_U3135) );
  AOI22_X1 U23722 ( .A1(n22196), .A2(n22128), .B1(n22127), .B2(n22195), .ZN(
        n22122) );
  AOI22_X1 U23723 ( .A1(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n22197), .B1(
        n22204), .B2(n22129), .ZN(n22121) );
  OAI211_X1 U23724 ( .C1(n22132), .C2(n22200), .A(n22122), .B(n22121), .ZN(
        P1_U3143) );
  AOI22_X1 U23725 ( .A1(n22128), .A2(n22202), .B1(n22127), .B2(n22201), .ZN(
        n22125) );
  AOI22_X1 U23726 ( .A1(P1_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n22205), .B1(
        n22204), .B2(n22123), .ZN(n22124) );
  OAI211_X1 U23727 ( .C1(n22126), .C2(n22218), .A(n22125), .B(n22124), .ZN(
        P1_U3151) );
  AOI22_X1 U23728 ( .A1(n22212), .A2(n22128), .B1(n22127), .B2(n22209), .ZN(
        n22131) );
  AOI22_X1 U23729 ( .A1(n22215), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n22129), .B2(n22213), .ZN(n22130) );
  OAI211_X1 U23730 ( .C1(n22132), .C2(n22218), .A(n22131), .B(n22130), .ZN(
        P1_U3159) );
  OAI22_X1 U23731 ( .A1(n22134), .A2(n11083), .B1(n22187), .B2(n22133), .ZN(
        n22135) );
  INV_X1 U23732 ( .A(n22135), .ZN(n22138) );
  AOI22_X1 U23733 ( .A1(P1_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n22136), .B1(
        n22142), .B2(n22214), .ZN(n22137) );
  OAI211_X1 U23734 ( .C1(n22139), .C2(n22193), .A(n22138), .B(n22137), .ZN(
        P1_U3040) );
  AOI22_X1 U23735 ( .A1(n22141), .A2(n22211), .B1(n22210), .B2(n22140), .ZN(
        n22145) );
  AOI22_X1 U23736 ( .A1(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n22143), .B1(
        n22142), .B2(n11084), .ZN(n22144) );
  OAI211_X1 U23737 ( .C1(n22208), .C2(n22146), .A(n22145), .B(n22144), .ZN(
        P1_U3048) );
  AOI22_X1 U23738 ( .A1(n22154), .A2(n22214), .B1(n22210), .B2(n22147), .ZN(
        n22151) );
  AOI22_X1 U23739 ( .A1(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n22149), .B1(
        n22148), .B2(n11084), .ZN(n22150) );
  OAI211_X1 U23740 ( .C1(n22152), .C2(n22193), .A(n22151), .B(n22150), .ZN(
        P1_U3056) );
  AOI22_X1 U23741 ( .A1(n22154), .A2(n11084), .B1(n22210), .B2(n22153), .ZN(
        n22158) );
  AOI22_X1 U23742 ( .A1(n22156), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n22155), .B2(n22214), .ZN(n22157) );
  OAI211_X1 U23743 ( .C1(n22159), .C2(n22193), .A(n22158), .B(n22157), .ZN(
        P1_U3064) );
  AOI22_X1 U23744 ( .A1(n22161), .A2(n11084), .B1(n22210), .B2(n22160), .ZN(
        n22165) );
  AOI22_X1 U23745 ( .A1(n22163), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n22214), .B2(n22162), .ZN(n22164) );
  OAI211_X1 U23746 ( .C1(n22166), .C2(n22193), .A(n22165), .B(n22164), .ZN(
        P1_U3088) );
  AOI22_X1 U23747 ( .A1(n22168), .A2(n22211), .B1(n22210), .B2(n22167), .ZN(
        n22172) );
  AOI22_X1 U23748 ( .A1(n22170), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11084), .B2(n22169), .ZN(n22171) );
  OAI211_X1 U23749 ( .C1(n22208), .C2(n22178), .A(n22172), .B(n22171), .ZN(
        P1_U3104) );
  AOI22_X1 U23750 ( .A1(n22174), .A2(n22211), .B1(n22210), .B2(n22173), .ZN(
        n22177) );
  AOI22_X1 U23751 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n22175), .B1(
        n22181), .B2(n22214), .ZN(n22176) );
  OAI211_X1 U23752 ( .C1(n11083), .C2(n22178), .A(n22177), .B(n22176), .ZN(
        P1_U3112) );
  AOI22_X1 U23753 ( .A1(n22180), .A2(n22214), .B1(n22210), .B2(n22179), .ZN(
        n22184) );
  AOI22_X1 U23754 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n22182), .B1(
        n22181), .B2(n11084), .ZN(n22183) );
  OAI211_X1 U23755 ( .C1(n22185), .C2(n22193), .A(n22184), .B(n22183), .ZN(
        P1_U3120) );
  OAI22_X1 U23756 ( .A1(n22200), .A2(n22208), .B1(n22187), .B2(n22186), .ZN(
        n22188) );
  INV_X1 U23757 ( .A(n22188), .ZN(n22192) );
  AOI22_X1 U23758 ( .A1(n22190), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11084), .B2(n22189), .ZN(n22191) );
  OAI211_X1 U23759 ( .C1(n22194), .C2(n22193), .A(n22192), .B(n22191), .ZN(
        P1_U3136) );
  AOI22_X1 U23760 ( .A1(n22196), .A2(n22211), .B1(n22210), .B2(n22195), .ZN(
        n22199) );
  AOI22_X1 U23761 ( .A1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n22197), .B1(
        n22204), .B2(n22214), .ZN(n22198) );
  OAI211_X1 U23762 ( .C1(n11083), .C2(n22200), .A(n22199), .B(n22198), .ZN(
        P1_U3144) );
  AOI22_X1 U23763 ( .A1(n22211), .A2(n22202), .B1(n22210), .B2(n22201), .ZN(
        n22207) );
  AOI22_X1 U23764 ( .A1(P1_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n22205), .B1(
        n22204), .B2(n11084), .ZN(n22206) );
  OAI211_X1 U23765 ( .C1(n22208), .C2(n22218), .A(n22207), .B(n22206), .ZN(
        P1_U3152) );
  AOI22_X1 U23766 ( .A1(n22212), .A2(n22211), .B1(n22210), .B2(n22209), .ZN(
        n22217) );
  AOI22_X1 U23767 ( .A1(n22215), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n22214), .B2(n22213), .ZN(n22216) );
  OAI211_X1 U23768 ( .C1(n11083), .C2(n22218), .A(n22217), .B(n22216), .ZN(
        P1_U3160) );
  AOI22_X1 U23769 ( .A1(n22221), .A2(n13452), .B1(n22220), .B2(n22219), .ZN(
        P1_U3486) );
  NAND2_X1 U13243 ( .A1(n13979), .A2(n11706), .ZN(n21860) );
  BUF_X2 U11103 ( .A(n12532), .Z(n12613) );
  AND2_X1 U11085 ( .A1(n11803), .A2(n11771), .ZN(n11476) );
  AND2_X1 U11132 ( .A1(n13615), .A2(n11499), .ZN(n11930) );
  CLKBUF_X1 U11141 ( .A(n14112), .Z(n10973) );
  INV_X2 U11150 ( .A(n13747), .ZN(n13905) );
  AND2_X1 U11157 ( .A1(n11115), .A2(n11407), .ZN(n15376) );
  CLKBUF_X1 U12187 ( .A(n17966), .Z(n10979) );
  CLKBUF_X1 U12320 ( .A(n17115), .Z(n17126) );
  CLKBUF_X2 U12581 ( .A(n17802), .Z(n10962) );
  CLKBUF_X1 U12628 ( .A(n18966), .Z(n19008) );
  NAND2_X1 U12712 ( .A1(n20577), .A2(n20449), .ZN(n11208) );
endmodule

