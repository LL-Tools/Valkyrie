

module b20_C_2inp_gates_syn ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, ADD_1068_U4, 
        ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58, ADD_1068_U59, 
        ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63, ADD_1068_U47, 
        ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51, ADD_1068_U52, 
        ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46, U126, U123, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439, P1_U3440, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462, P1_U3465, P1_U3468, 
        P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, 
        P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3509, 
        P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, 
        P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, 
        P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, 
        P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, 
        P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, 
        P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, 
        P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3554, P1_U3555, 
        P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, 
        P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, 
        P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, 
        P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, 
        P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U3973, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376, P2_U3377, P2_U3263, 
        P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, 
        P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, 
        P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, 
        P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, 
        P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399, P2_U3402, P2_U3405, 
        P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420, P2_U3423, P2_U3426, 
        P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441, P2_U3444, P2_U3446, 
        P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451, P2_U3452, P2_U3453, 
        P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458, P2_U3459, P2_U3460, 
        P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465, P2_U3466, P2_U3467, 
        P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472, P2_U3473, P2_U3474, 
        P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479, P2_U3480, P2_U3481, 
        P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486, P2_U3487, P2_U3488, 
        P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, 
        P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, 
        P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, 
        P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3491, P2_U3492, 
        P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, 
        P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, 
        P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, 
        P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, 
        P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180, P2_U3179, P2_U3178, 
        P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, P2_U3171, 
        P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, P2_U3164, 
        P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, P2_U3157, 
        P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151, P2_U3150, P2_U3893, 
        keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, 
        keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, 
        keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, 
        keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, 
        keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, 
        keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, 
        keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, 
        keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, 
        keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, 
        keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, 
        keyinput60, keyinput61, keyinput62, keyinput63 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4277,
         n4278, n4279, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288,
         n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298,
         n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308,
         n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318,
         n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328,
         n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338,
         n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348,
         n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358,
         n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368,
         n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378,
         n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388,
         n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398,
         n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408,
         n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418,
         n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428,
         n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438,
         n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448,
         n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458,
         n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468,
         n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478,
         n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488,
         n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498,
         n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508,
         n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518,
         n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528,
         n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538,
         n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548,
         n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558,
         n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568,
         n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578,
         n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588,
         n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598,
         n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608,
         n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618,
         n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628,
         n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638,
         n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648,
         n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658,
         n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668,
         n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678,
         n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688,
         n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698,
         n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708,
         n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718,
         n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728,
         n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738,
         n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748,
         n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758,
         n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768,
         n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778,
         n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788,
         n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798,
         n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808,
         n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818,
         n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828,
         n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838,
         n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848,
         n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858,
         n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868,
         n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878,
         n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888,
         n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898,
         n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908,
         n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918,
         n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928,
         n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938,
         n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948,
         n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958,
         n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968,
         n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978,
         n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988,
         n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998,
         n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008,
         n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018,
         n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028,
         n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038,
         n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048,
         n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058,
         n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068,
         n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078,
         n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088,
         n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098,
         n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108,
         n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118,
         n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128,
         n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138,
         n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148,
         n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158,
         n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168,
         n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178,
         n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188,
         n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198,
         n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208,
         n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218,
         n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228,
         n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238,
         n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248,
         n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258,
         n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268,
         n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278,
         n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288,
         n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298,
         n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308,
         n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318,
         n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328,
         n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338,
         n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348,
         n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358,
         n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368,
         n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378,
         n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388,
         n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398,
         n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408,
         n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418,
         n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428,
         n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438,
         n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448,
         n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458,
         n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468,
         n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478,
         n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488,
         n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498,
         n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508,
         n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518,
         n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528,
         n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538,
         n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548,
         n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558,
         n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568,
         n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578,
         n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588,
         n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598,
         n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608,
         n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618,
         n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628,
         n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638,
         n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648,
         n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658,
         n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668,
         n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678,
         n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688,
         n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698,
         n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708,
         n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718,
         n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728,
         n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738,
         n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748,
         n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758,
         n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768,
         n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778,
         n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788,
         n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798,
         n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808,
         n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818,
         n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828,
         n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838,
         n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848,
         n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858,
         n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868,
         n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878,
         n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888,
         n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898,
         n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908,
         n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918,
         n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928,
         n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938,
         n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948,
         n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958,
         n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968,
         n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978,
         n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988,
         n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998,
         n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008,
         n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018,
         n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028,
         n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038,
         n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048,
         n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058,
         n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068,
         n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078,
         n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088,
         n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098,
         n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108,
         n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118,
         n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128,
         n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138,
         n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148,
         n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158,
         n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168,
         n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178,
         n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188,
         n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198,
         n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208,
         n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218,
         n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228,
         n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238,
         n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248,
         n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258,
         n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268,
         n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278,
         n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288,
         n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298,
         n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308,
         n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318,
         n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328,
         n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338,
         n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348,
         n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358,
         n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368,
         n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378,
         n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388,
         n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398,
         n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408,
         n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418,
         n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428,
         n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438,
         n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448,
         n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458,
         n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468,
         n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478,
         n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488,
         n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498,
         n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508,
         n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518,
         n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528,
         n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538,
         n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548,
         n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558,
         n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568,
         n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578,
         n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588,
         n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598,
         n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608,
         n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618,
         n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628,
         n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638,
         n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648,
         n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658,
         n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668,
         n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678,
         n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688,
         n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698,
         n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708,
         n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718,
         n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728,
         n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738,
         n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748,
         n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758,
         n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768,
         n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778,
         n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788,
         n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798,
         n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808,
         n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818,
         n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828,
         n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838,
         n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848,
         n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858,
         n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868,
         n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878,
         n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888,
         n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898,
         n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908,
         n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918,
         n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928,
         n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938,
         n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948,
         n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958,
         n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968,
         n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978,
         n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988,
         n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998,
         n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008,
         n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018,
         n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028,
         n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038,
         n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048,
         n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058,
         n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068,
         n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078,
         n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088,
         n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098,
         n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108,
         n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118,
         n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128,
         n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138,
         n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148,
         n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158,
         n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168,
         n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178,
         n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188,
         n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198,
         n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208,
         n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218,
         n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228,
         n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238,
         n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248,
         n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258,
         n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268,
         n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278,
         n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288,
         n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298,
         n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308,
         n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318,
         n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328,
         n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338,
         n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348,
         n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358,
         n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368,
         n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378,
         n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388,
         n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398,
         n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408,
         n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418,
         n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428,
         n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438,
         n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448,
         n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458,
         n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468,
         n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478,
         n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488,
         n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498,
         n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508,
         n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518,
         n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528,
         n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538,
         n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548,
         n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558,
         n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568,
         n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578,
         n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588,
         n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598,
         n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608,
         n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618,
         n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628,
         n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638,
         n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648,
         n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658,
         n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668,
         n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678,
         n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688,
         n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698,
         n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708,
         n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718,
         n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728,
         n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738,
         n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748,
         n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758,
         n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768,
         n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778,
         n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788,
         n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798,
         n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808,
         n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818,
         n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828,
         n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838,
         n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848,
         n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858,
         n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868,
         n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878,
         n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888,
         n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898,
         n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908,
         n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918,
         n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928,
         n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938,
         n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948,
         n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958,
         n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968,
         n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978,
         n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988,
         n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998,
         n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008,
         n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018,
         n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028,
         n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038,
         n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048,
         n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058,
         n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068,
         n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078,
         n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088,
         n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098,
         n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108,
         n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118,
         n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128,
         n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138,
         n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148,
         n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158,
         n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168,
         n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178,
         n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188,
         n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198,
         n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208,
         n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218,
         n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228,
         n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238,
         n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248,
         n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258,
         n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268,
         n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278,
         n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288,
         n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298,
         n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308,
         n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318,
         n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328,
         n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338,
         n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348,
         n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358,
         n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368,
         n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378,
         n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388,
         n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398,
         n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408,
         n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418,
         n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428,
         n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438,
         n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448,
         n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458,
         n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468,
         n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478,
         n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488,
         n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498,
         n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508,
         n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518,
         n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528,
         n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538,
         n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548,
         n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558,
         n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568,
         n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578,
         n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588,
         n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598,
         n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608,
         n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618,
         n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628,
         n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638,
         n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648,
         n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658,
         n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668,
         n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678,
         n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688,
         n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698,
         n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708,
         n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718,
         n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728,
         n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738,
         n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748,
         n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758,
         n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768,
         n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778,
         n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788,
         n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798,
         n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808,
         n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818,
         n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828,
         n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838,
         n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848,
         n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858,
         n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868,
         n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878,
         n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888,
         n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898,
         n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908,
         n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918,
         n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928,
         n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938,
         n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948,
         n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958,
         n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968,
         n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978,
         n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988,
         n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998,
         n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008,
         n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018,
         n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028,
         n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038,
         n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048,
         n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058,
         n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068,
         n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078,
         n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088,
         n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098,
         n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108,
         n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118,
         n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128,
         n9129, n9130, n9131, n9132, n9133, n9135, n9136, n9137, n9138, n9139,
         n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149,
         n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159,
         n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169,
         n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179,
         n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189,
         n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199,
         n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209,
         n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219,
         n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229,
         n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239,
         n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249,
         n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259,
         n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269,
         n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279,
         n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289,
         n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299,
         n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309,
         n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319,
         n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329,
         n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339,
         n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349,
         n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359,
         n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369,
         n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379,
         n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389,
         n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399,
         n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409,
         n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419,
         n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429,
         n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439,
         n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449,
         n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459,
         n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469,
         n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479,
         n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489,
         n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499,
         n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509,
         n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519,
         n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529,
         n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539,
         n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549,
         n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559,
         n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569,
         n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579,
         n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589,
         n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599,
         n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609,
         n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619,
         n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629,
         n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639,
         n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649,
         n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659,
         n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669,
         n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679,
         n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689,
         n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699,
         n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709,
         n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719,
         n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729,
         n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739,
         n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749,
         n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759,
         n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769,
         n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779,
         n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789,
         n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799,
         n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809,
         n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819,
         n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829,
         n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839,
         n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849,
         n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859,
         n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869,
         n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879,
         n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889,
         n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899,
         n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909,
         n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919,
         n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929,
         n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939,
         n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949,
         n9950, n9951, n9952, n9953, n9954, n9956, n9957, n9958, n9959, n9960,
         n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970,
         n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980,
         n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990,
         n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
         n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
         n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
         n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
         n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
         n10265, n10266, n10267;

  AOI21_X1 U4773 ( .B1(n7598), .B2(n8096), .A(n8095), .ZN(n7710) );
  NAND2_X1 U4774 ( .A1(n7181), .A2(n7264), .ZN(n7274) );
  INV_X1 U4775 ( .A(n7056), .ZN(n7930) );
  NAND2_X1 U4776 ( .A1(n8216), .A2(n8229), .ZN(n8158) );
  INV_X1 U4777 ( .A(n7819), .ZN(n6923) );
  BUF_X1 U4778 ( .A(n5613), .Z(n5603) );
  INV_X1 U4779 ( .A(n6986), .ZN(n6991) );
  NAND3_X1 U4780 ( .A1(n5257), .A2(n5256), .A3(n5255), .ZN(n6849) );
  OAI211_X1 U4781 ( .C1(n8232), .C2(n5268), .A(n5267), .B(n5266), .ZN(n10043)
         );
  BUF_X2 U4782 ( .A(n5959), .Z(n8008) );
  OAI211_X1 U4783 ( .C1(n6614), .C2(n4458), .A(n5954), .B(n5953), .ZN(n10189)
         );
  BUF_X1 U4784 ( .A(n5958), .Z(n5980) );
  CLKBUF_X3 U4786 ( .A(n5259), .Z(n6658) );
  INV_X1 U4787 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n5013) );
  INV_X1 U4789 ( .A(P2_RD_REG_SCAN_IN), .ZN(n5014) );
  INV_X2 U4790 ( .A(n4279), .ZN(n6283) );
  NAND2_X1 U4791 ( .A1(n8415), .A2(n8419), .ZN(n8453) );
  INV_X1 U4792 ( .A(n5922), .ZN(n8216) );
  INV_X1 U4793 ( .A(n7056), .ZN(n4289) );
  INV_X1 U4794 ( .A(n6678), .ZN(n5323) );
  INV_X1 U4796 ( .A(n6923), .ZN(n9132) );
  AND2_X2 U4797 ( .A1(n6678), .A2(n8003), .ZN(n5613) );
  NAND2_X1 U4798 ( .A1(n4594), .A2(n9077), .ZN(n7880) );
  AND3_X1 U4799 ( .A1(n5140), .A2(n5141), .A3(n5139), .ZN(n5858) );
  INV_X1 U4800 ( .A(n8397), .ZN(n7782) );
  CLKBUF_X2 U4801 ( .A(n5969), .Z(n8011) );
  INV_X1 U4802 ( .A(n8158), .ZN(n8165) );
  INV_X1 U4803 ( .A(n4288), .ZN(n9129) );
  BUF_X1 U4804 ( .A(n9117), .Z(n9166) );
  NAND2_X1 U4805 ( .A1(n4452), .A2(n9630), .ZN(n6468) );
  INV_X1 U4806 ( .A(n5699), .ZN(n5657) );
  INV_X1 U4807 ( .A(n10042), .ZN(n9816) );
  AND2_X1 U4808 ( .A1(n4560), .A2(n5324), .ZN(n5341) );
  INV_X1 U4809 ( .A(n7043), .ZN(n10066) );
  XNOR2_X1 U4810 ( .A(n5745), .B(P1_IR_REG_22__SCAN_IN), .ZN(n4471) );
  OAI21_X1 U4811 ( .B1(n7720), .B2(n6598), .A(n6597), .ZN(n8732) );
  XNOR2_X1 U4812 ( .A(n5930), .B(P2_IR_REG_30__SCAN_IN), .ZN(n5934) );
  INV_X1 U4814 ( .A(n5933), .ZN(n8907) );
  INV_X1 U4815 ( .A(n9788), .ZN(n9630) );
  XNOR2_X1 U4816 ( .A(n4559), .B(n5150), .ZN(n9389) );
  NAND2_X1 U4817 ( .A1(n5172), .A2(n8255), .ZN(n4685) );
  AOI21_X1 U4818 ( .B1(n8505), .B2(n4313), .A(n8504), .ZN(n8516) );
  AND2_X4 U4819 ( .A1(n9706), .A2(n4859), .ZN(n9649) );
  OAI22_X1 U4820 ( .A1(n7042), .A2(n4909), .B1(n7040), .B2(n7041), .ZN(n7055)
         );
  BUF_X4 U4821 ( .A(n6328), .Z(n4279) );
  OR2_X4 U4822 ( .A1(n9618), .A2(n9839), .ZN(n9619) );
  NAND2_X1 U4823 ( .A1(n6614), .A2(n6658), .ZN(n4267) );
  NAND2_X1 U4824 ( .A1(n6614), .A2(n6658), .ZN(n4268) );
  INV_X4 U4825 ( .A(n8008), .ZN(n6195) );
  OR2_X4 U4826 ( .A1(n10009), .A2(n9157), .ZN(n4986) );
  NAND2_X2 U4827 ( .A1(n10010), .A2(n10091), .ZN(n10009) );
  OAI22_X2 U4828 ( .A1(n8698), .A2(n6560), .B1(n8707), .B2(n8272), .ZN(n8683)
         );
  XNOR2_X2 U4829 ( .A(n5030), .B(SI_3_), .ZN(n5243) );
  AOI211_X2 U4830 ( .C1(n9644), .C2(n10046), .A(n9643), .B(n9642), .ZN(n9645)
         );
  AOI21_X2 U4831 ( .B1(n9764), .B2(n9763), .A(n6451), .ZN(n9749) );
  OR2_X2 U4832 ( .A1(n5929), .A2(n5900), .ZN(n5901) );
  OAI22_X2 U4833 ( .A1(n7231), .A2(n6530), .B1(n10174), .B2(n10205), .ZN(n7257) );
  INV_X1 U4834 ( .A(n9057), .ZN(n4269) );
  INV_X1 U4835 ( .A(n4269), .ZN(n4270) );
  AOI21_X2 U4836 ( .B1(n8446), .B2(n8445), .A(n8444), .ZN(n8483) );
  OAI21_X2 U4837 ( .B1(n5714), .B2(P1_IR_REG_21__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5745) );
  OAI21_X2 U4838 ( .B1(n7601), .B2(n6594), .A(n6593), .ZN(n7720) );
  OR2_X1 U4839 ( .A1(n5959), .A2(n9060), .ZN(n5960) );
  NAND2_X2 U4840 ( .A1(n4887), .A2(n4325), .ZN(n4882) );
  INV_X2 U4841 ( .A(n6468), .ZN(n5708) );
  INV_X1 U4842 ( .A(n10176), .ZN(n6523) );
  NAND4_X1 U4843 ( .A1(n5965), .A2(n5964), .A3(n5963), .A4(n5962), .ZN(n10176)
         );
  NAND2_X1 U4844 ( .A1(n5927), .A2(n8225), .ZN(n6328) );
  INV_X1 U4845 ( .A(n5973), .ZN(n4285) );
  BUF_X4 U4846 ( .A(n5974), .Z(n4271) );
  CLKBUF_X2 U4847 ( .A(n5309), .Z(n5654) );
  INV_X1 U4849 ( .A(n5934), .ZN(n8902) );
  NOR2_X1 U4850 ( .A1(n7586), .A2(n7447), .ZN(n4604) );
  BUF_X1 U4851 ( .A(n5912), .Z(n4284) );
  OR2_X1 U4852 ( .A1(n4804), .A2(n5900), .ZN(n4803) );
  NOR2_X1 U4853 ( .A1(n9857), .A2(n4702), .ZN(n9860) );
  AOI211_X1 U4854 ( .C1(n9882), .C2(n9348), .A(n9175), .B(n9174), .ZN(n9176)
         );
  NAND2_X1 U4855 ( .A1(n4704), .A2(n9668), .ZN(n9857) );
  NOR3_X1 U4856 ( .A1(n5740), .A2(n5850), .A3(n4445), .ZN(n5799) );
  NAND3_X1 U4857 ( .A1(n4891), .A2(n8169), .A3(n4889), .ZN(n8625) );
  AND2_X1 U4858 ( .A1(n5189), .A2(n5188), .ZN(n9330) );
  NAND2_X1 U4859 ( .A1(n9729), .A2(n4991), .ZN(n9726) );
  CLKBUF_X1 U4860 ( .A(n9203), .Z(n4443) );
  OR2_X1 U4861 ( .A1(n9858), .A2(n4703), .ZN(n4702) );
  NAND2_X1 U4862 ( .A1(n4562), .A2(n4561), .ZN(n7504) );
  NAND2_X1 U4863 ( .A1(n7439), .A2(n4565), .ZN(n4561) );
  NAND2_X1 U4864 ( .A1(n4564), .A2(n4324), .ZN(n4562) );
  NAND2_X1 U4865 ( .A1(n7542), .A2(n7541), .ZN(n7544) );
  NAND2_X1 U4866 ( .A1(n6226), .A2(n6225), .ZN(n8866) );
  NAND2_X1 U4867 ( .A1(n5200), .A2(n5199), .ZN(n9908) );
  NAND2_X1 U4868 ( .A1(n8080), .A2(n8081), .ZN(n8187) );
  OR2_X1 U4869 ( .A1(n6536), .A2(n7565), .ZN(n8080) );
  NOR2_X1 U4870 ( .A1(n4928), .A2(n7804), .ZN(n4927) );
  NAND2_X1 U4871 ( .A1(n7095), .A2(n7097), .ZN(n7096) );
  NAND2_X1 U4872 ( .A1(n5397), .A2(n5396), .ZN(n9299) );
  INV_X1 U4873 ( .A(n9191), .ZN(n9928) );
  NAND2_X1 U4874 ( .A1(n6084), .A2(n6083), .ZN(n7770) );
  AND2_X1 U4875 ( .A1(n5427), .A2(n5426), .ZN(n9191) );
  OR2_X1 U4876 ( .A1(n7485), .A2(n6531), .ZN(n7448) );
  CLKBUF_X1 U4877 ( .A(n8380), .Z(n8371) );
  AND2_X1 U4878 ( .A1(n7215), .A2(n6482), .ZN(n4836) );
  XNOR2_X1 U4879 ( .A(n4442), .B(n5394), .ZN(n6736) );
  XOR2_X1 U4880 ( .A(n4278), .B(n7803), .Z(n7804) );
  NAND2_X1 U4881 ( .A1(n8028), .A2(n8027), .ZN(n8031) );
  CLKBUF_X1 U4882 ( .A(n9826), .Z(n10046) );
  NAND2_X1 U4883 ( .A1(n5360), .A2(n5359), .ZN(n9157) );
  BUF_X4 U4884 ( .A(n9132), .Z(n4278) );
  INV_X2 U4885 ( .A(n10108), .ZN(n4272) );
  NAND2_X1 U4886 ( .A1(n6910), .A2(n6516), .ZN(n6581) );
  INV_X1 U4887 ( .A(n5341), .ZN(n6425) );
  NAND2_X1 U4889 ( .A1(n5810), .A2(n5812), .ZN(n6419) );
  INV_X2 U4890 ( .A(n6515), .ZN(n6516) );
  NAND2_X1 U4891 ( .A1(n4707), .A2(n5037), .ZN(n5325) );
  NAND2_X1 U4892 ( .A1(n4708), .A2(n4876), .ZN(n5354) );
  AND4_X1 U4893 ( .A1(n5944), .A2(n5943), .A3(n5942), .A4(n5941), .ZN(n6741)
         );
  NAND2_X1 U4894 ( .A1(n4360), .A2(n5292), .ZN(n9374) );
  OAI21_X1 U4895 ( .B1(n5318), .B2(n4482), .A(n4480), .ZN(n4708) );
  NAND2_X1 U4896 ( .A1(n4441), .A2(n5034), .ZN(n5318) );
  INV_X2 U4897 ( .A(n4286), .ZN(n8012) );
  AND4_X1 U4898 ( .A1(n5241), .A2(n5240), .A3(n5239), .A4(n5238), .ZN(n7038)
         );
  CLKBUF_X1 U4899 ( .A(n6782), .Z(n4452) );
  OAI211_X1 U4900 ( .C1(n5242), .C2(n4866), .A(n4483), .B(n4484), .ZN(n4441)
         );
  CLKBUF_X1 U4901 ( .A(n5973), .Z(n4286) );
  OR2_X1 U4902 ( .A1(n6785), .A2(n6783), .ZN(n10008) );
  INV_X2 U4904 ( .A(n5678), .ZN(n5694) );
  CLKBUF_X1 U4905 ( .A(n5872), .Z(n6464) );
  INV_X1 U4906 ( .A(n7557), .ZN(n4603) );
  NAND2_X1 U4907 ( .A1(n5865), .A2(n5864), .ZN(n7557) );
  INV_X2 U4908 ( .A(n6614), .ZN(n8005) );
  CLKBUF_X1 U4909 ( .A(n7223), .Z(n4469) );
  NAND2_X1 U4910 ( .A1(n6614), .A2(n6658), .ZN(n5959) );
  NAND2_X2 U4911 ( .A1(n6962), .A2(n9057), .ZN(n10152) );
  XNOR2_X1 U4912 ( .A(n5743), .B(n5742), .ZN(n7223) );
  CLKBUF_X1 U4913 ( .A(n6367), .Z(n6726) );
  NAND2_X1 U4914 ( .A1(n5869), .A2(n5868), .ZN(n7447) );
  OR2_X1 U4915 ( .A1(n5741), .A2(n5168), .ZN(n5743) );
  NOR2_X1 U4916 ( .A1(n5405), .A2(n4725), .ZN(n4724) );
  NAND2_X1 U4917 ( .A1(n9956), .A2(n5167), .ZN(n9964) );
  NAND3_X1 U4918 ( .A1(n5906), .A2(n4758), .A3(n5907), .ZN(n4757) );
  XNOR2_X1 U4919 ( .A(n5870), .B(n4936), .ZN(n7586) );
  NAND2_X1 U4920 ( .A1(n5862), .A2(n5861), .ZN(n5869) );
  NAND2_X1 U4921 ( .A1(n5165), .A2(n5149), .ZN(n8232) );
  NAND3_X1 U4922 ( .A1(n6330), .A2(P2_IR_REG_31__SCAN_IN), .A3(
        P2_IR_REG_27__SCAN_IN), .ZN(n5906) );
  INV_X1 U4923 ( .A(n8255), .ZN(n4273) );
  NAND2_X1 U4924 ( .A1(n4908), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5930) );
  OAI21_X1 U4925 ( .B1(n5197), .B2(P1_IR_REG_16__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5475) );
  NAND2_X1 U4926 ( .A1(n4558), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4559) );
  OR2_X1 U4927 ( .A1(n5169), .A2(n5168), .ZN(n5171) );
  NAND2_X2 U4928 ( .A1(n6658), .A2(P1_U3086), .ZN(n9963) );
  AND2_X1 U4929 ( .A1(n4803), .A2(P2_IR_REG_29__SCAN_IN), .ZN(n4802) );
  XNOR2_X1 U4930 ( .A(n4535), .B(n5957), .ZN(n9057) );
  NAND2_X1 U4931 ( .A1(n4536), .A2(n8985), .ZN(n5981) );
  AND2_X1 U4932 ( .A1(n5899), .A2(n5928), .ZN(n4804) );
  OAI211_X1 U4933 ( .C1(n5264), .C2(n4642), .A(n5265), .B(n4641), .ZN(n6823)
         );
  AND3_X1 U4934 ( .A1(n4994), .A2(n4996), .A3(n4995), .ZN(n5146) );
  AND2_X1 U4935 ( .A1(n4997), .A2(n4998), .ZN(n5857) );
  NAND4_X1 U4936 ( .A1(n5888), .A2(n5889), .A3(n6052), .A4(n6054), .ZN(n4808)
         );
  AND3_X1 U4937 ( .A1(n5145), .A2(n5143), .A3(n5144), .ZN(n5856) );
  AND2_X1 U4938 ( .A1(n5896), .A2(n4903), .ZN(n4902) );
  INV_X1 U4939 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n4607) );
  INV_X1 U4940 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n4606) );
  NOR2_X1 U4941 ( .A1(P2_IR_REG_4__SCAN_IN), .A2(P2_IR_REG_5__SCAN_IN), .ZN(
        n5890) );
  NOR2_X1 U4942 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n5891) );
  NOR2_X1 U4943 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), .ZN(
        n5140) );
  NOR2_X1 U4944 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n4996) );
  NOR2_X1 U4945 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .ZN(
        n4995) );
  INV_X4 U4946 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  NOR2_X1 U4947 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n4997) );
  NOR2_X1 U4948 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n4998) );
  NOR2_X1 U4949 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n5894) );
  INV_X1 U4950 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n6052) );
  INV_X1 U4951 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n6054) );
  NOR2_X1 U4952 ( .A1(P2_IR_REG_25__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), .ZN(
        n5902) );
  INV_X1 U4953 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n5889) );
  NOR2_X1 U4954 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n5888) );
  NOR2_X1 U4955 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), .ZN(
        n5895) );
  INV_X1 U4956 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n4605) );
  NOR2_X1 U4957 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5892) );
  INV_X4 U4958 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  AND2_X1 U4959 ( .A1(n8517), .A2(n8533), .ZN(n4463) );
  INV_X1 U4960 ( .A(n6852), .ZN(n4274) );
  INV_X2 U4961 ( .A(n4429), .ZN(n6295) );
  OR2_X1 U4962 ( .A1(n8831), .A2(n8896), .ZN(n4418) );
  OR2_X1 U4963 ( .A1(n8831), .A2(n8747), .ZN(n4417) );
  OR2_X1 U4964 ( .A1(n8831), .A2(n8813), .ZN(n4416) );
  NAND2_X2 U4965 ( .A1(n5244), .A2(n5146), .ZN(n5859) );
  NOR2_X2 U4966 ( .A1(n7880), .A2(n7879), .ZN(n9203) );
  AND2_X4 U4967 ( .A1(n9744), .A2(n9725), .ZN(n9706) );
  XNOR2_X1 U4969 ( .A(n6517), .B(n6328), .ZN(n5939) );
  INV_X1 U4970 ( .A(n4279), .ZN(n4275) );
  NAND3_X1 U4971 ( .A1(n10008), .A2(n6790), .A3(n6784), .ZN(n6852) );
  OAI211_X1 U4972 ( .C1(n6659), .C2(n8003), .A(n8240), .B(n5263), .ZN(n5267)
         );
  NAND2_X1 U4973 ( .A1(n4471), .A2(n9788), .ZN(n6787) );
  NAND2_X1 U4974 ( .A1(n8232), .A2(n9389), .ZN(n4277) );
  OAI21_X2 U4975 ( .B1(n8625), .B2(n8150), .A(n8151), .ZN(n8607) );
  CLKBUF_X1 U4977 ( .A(n9389), .Z(n4281) );
  NAND2_X1 U4978 ( .A1(n5016), .A2(n5015), .ZN(n4282) );
  NAND2_X1 U4979 ( .A1(n5016), .A2(n5015), .ZN(n4283) );
  NAND2_X1 U4980 ( .A1(n8902), .A2(n8907), .ZN(n5974) );
  NOR2_X2 U4981 ( .A1(n10034), .A2(n4833), .ZN(n7029) );
  NAND3_X1 U4982 ( .A1(n10008), .A2(n6790), .A3(n6784), .ZN(n4287) );
  NAND3_X1 U4983 ( .A1(n10008), .A2(n6790), .A3(n6784), .ZN(n4288) );
  INV_X2 U4984 ( .A(n7056), .ZN(n4290) );
  NAND2_X4 U4985 ( .A1(n6781), .A2(n6790), .ZN(n7056) );
  NAND2_X1 U4986 ( .A1(n4552), .A2(n4551), .ZN(n9845) );
  AOI21_X1 U4987 ( .B1(n4554), .B2(n4556), .A(n4363), .ZN(n4551) );
  AND2_X1 U4988 ( .A1(n5646), .A2(n6468), .ZN(n4682) );
  AOI21_X1 U4989 ( .B1(n4742), .B2(n4740), .A(n4349), .ZN(n4739) );
  INV_X1 U4990 ( .A(n6573), .ZN(n4740) );
  INV_X1 U4991 ( .A(n8601), .ZN(n8168) );
  OR2_X1 U4992 ( .A1(n8840), .A2(n8620), .ZN(n8155) );
  INV_X1 U4993 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n4903) );
  INV_X1 U4994 ( .A(n9964), .ZN(n5172) );
  OR2_X1 U4995 ( .A1(n9839), .A2(n7171), .ZN(n5791) );
  CLKBUF_X2 U4996 ( .A(n6024), .Z(n6323) );
  AND2_X1 U4997 ( .A1(n5934), .A2(n5933), .ZN(n6024) );
  NAND2_X1 U4998 ( .A1(n6459), .A2(n4965), .ZN(n4964) );
  NAND2_X1 U4999 ( .A1(n8029), .A2(n8165), .ZN(n4456) );
  NAND2_X1 U5000 ( .A1(n8030), .A2(n8158), .ZN(n4455) );
  NOR2_X1 U5001 ( .A1(n4666), .A2(n4660), .ZN(n4659) );
  AND2_X1 U5002 ( .A1(n4766), .A2(n8120), .ZN(n4454) );
  INV_X1 U5003 ( .A(n8157), .ZN(n4771) );
  AND2_X1 U5004 ( .A1(n4739), .A2(n4366), .ZN(n4738) );
  INV_X1 U5005 ( .A(n5750), .ZN(n4675) );
  NAND2_X1 U5006 ( .A1(n4504), .A2(n4500), .ZN(n4503) );
  INV_X1 U5007 ( .A(n4504), .ZN(n4498) );
  NOR2_X1 U5008 ( .A1(n6404), .A2(n6403), .ZN(n6406) );
  AND2_X1 U5009 ( .A1(n4828), .A2(n4826), .ZN(n6404) );
  NOR2_X1 U5010 ( .A1(n6401), .A2(n4827), .ZN(n4826) );
  NAND2_X1 U5011 ( .A1(n7284), .A2(n7358), .ZN(n6048) );
  OR2_X1 U5012 ( .A1(n6321), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n8246) );
  INV_X1 U5013 ( .A(n4742), .ZN(n4741) );
  AND2_X1 U5014 ( .A1(n4321), .A2(n8159), .ZN(n8597) );
  OR2_X1 U5015 ( .A1(n8853), .A2(n8621), .ZN(n8169) );
  OAI21_X1 U5016 ( .B1(n8199), .B2(n4750), .A(n6568), .ZN(n4749) );
  OR2_X1 U5017 ( .A1(n8878), .A2(n8707), .ZN(n8107) );
  NOR2_X1 U5018 ( .A1(n8721), .A2(n6555), .ZN(n6556) );
  NAND2_X1 U5019 ( .A1(n6551), .A2(n4988), .ZN(n4756) );
  INV_X1 U5020 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n6340) );
  INV_X1 U5021 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5915) );
  OR2_X1 U5022 ( .A1(n6020), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n6051) );
  OR2_X1 U5023 ( .A1(n5981), .A2(P2_IR_REG_3__SCAN_IN), .ZN(n5991) );
  OR2_X1 U5024 ( .A1(n8244), .A2(n9625), .ZN(n5794) );
  NAND2_X1 U5025 ( .A1(n4870), .A2(n5628), .ZN(n4873) );
  NAND2_X1 U5026 ( .A1(n4875), .A2(n4871), .ZN(n4870) );
  INV_X1 U5027 ( .A(n4953), .ZN(n4952) );
  OAI21_X1 U5028 ( .B1(n4955), .B2(n4954), .A(n6449), .ZN(n4953) );
  OR2_X1 U5029 ( .A1(n9893), .A2(n9360), .ZN(n6449) );
  INV_X1 U5030 ( .A(n4960), .ZN(n4570) );
  NAND2_X1 U5031 ( .A1(n5341), .A2(n9373), .ZN(n5819) );
  NAND2_X1 U5032 ( .A1(n7578), .A2(n9083), .ZN(n6483) );
  AND2_X1 U5033 ( .A1(n9951), .A2(n6777), .ZN(n6976) );
  NAND2_X1 U5034 ( .A1(n4710), .A2(n4709), .ZN(n5687) );
  AOI21_X1 U5035 ( .B1(n4712), .B2(n4714), .A(n4383), .ZN(n4709) );
  XNOR2_X1 U5036 ( .A(n5687), .B(n5685), .ZN(n5684) );
  NOR2_X1 U5037 ( .A1(n4380), .A2(P1_IR_REG_26__SCAN_IN), .ZN(n4701) );
  AOI21_X1 U5038 ( .B1(n5573), .B2(n5115), .A(n5114), .ZN(n5590) );
  AND2_X1 U5039 ( .A1(n5120), .A2(n5119), .ZN(n5589) );
  NAND2_X1 U5040 ( .A1(n4502), .A2(n4504), .ZN(n5053) );
  OR2_X1 U5041 ( .A1(n6406), .A2(n6405), .ZN(n4824) );
  NOR2_X1 U5042 ( .A1(n4334), .A2(n4812), .ZN(n4811) );
  INV_X1 U5043 ( .A(n4814), .ZN(n4812) );
  NAND2_X1 U5044 ( .A1(n4329), .A2(n4450), .ZN(n4449) );
  NAND2_X1 U5045 ( .A1(n8763), .A2(n8823), .ZN(n4450) );
  NAND2_X1 U5046 ( .A1(n8216), .A2(n8205), .ZN(n8225) );
  AND3_X1 U5047 ( .A1(n6189), .A2(n6188), .A3(n6187), .ZN(n8313) );
  AND2_X1 U5048 ( .A1(n8902), .A2(n5933), .ZN(n5969) );
  OR2_X1 U5049 ( .A1(n6957), .A2(n6964), .ZN(n4614) );
  OR2_X1 U5050 ( .A1(n7173), .A2(n4621), .ZN(n4620) );
  AND2_X1 U5051 ( .A1(n7174), .A2(n7185), .ZN(n4621) );
  NAND2_X1 U5052 ( .A1(n8465), .A2(n8464), .ZN(n8491) );
  OAI21_X1 U5053 ( .B1(n4880), .B2(n4331), .A(n4291), .ZN(n4879) );
  NAND2_X1 U5054 ( .A1(n6172), .A2(n4588), .ZN(n6214) );
  AND2_X1 U5055 ( .A1(n4304), .A2(n4589), .ZN(n4588) );
  INV_X1 U5056 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n4589) );
  OR2_X1 U5057 ( .A1(n7993), .A2(n8383), .ZN(n8097) );
  OR2_X1 U5058 ( .A1(n6899), .A2(n6898), .ZN(n6908) );
  AND2_X1 U5059 ( .A1(n8853), .A2(n8642), .ZN(n6569) );
  AND2_X1 U5060 ( .A1(n6259), .A2(n6258), .ZN(n8631) );
  OR2_X1 U5061 ( .A1(n6616), .A2(n8158), .ZN(n8739) );
  NAND2_X1 U5062 ( .A1(n6579), .A2(n8225), .ZN(n10178) );
  INV_X4 U5063 ( .A(n5980), .ZN(n8007) );
  INV_X1 U5064 ( .A(n4808), .ZN(n4759) );
  AND2_X1 U5065 ( .A1(n7830), .A2(n4913), .ZN(n4912) );
  AND2_X1 U5066 ( .A1(n9252), .A2(n4973), .ZN(n7830) );
  NAND2_X1 U5067 ( .A1(n4274), .A2(n9377), .ZN(n4467) );
  AOI21_X1 U5068 ( .B1(n7884), .B2(n6986), .A(n4466), .ZN(n4465) );
  AND2_X1 U5069 ( .A1(n6791), .A2(P1_IR_REG_0__SCAN_IN), .ZN(n4466) );
  NAND2_X1 U5070 ( .A1(n7949), .A2(n9237), .ZN(n9239) );
  OAI21_X1 U5071 ( .B1(n9172), .B2(n4312), .A(n4932), .ZN(n7949) );
  INV_X1 U5072 ( .A(n4933), .ZN(n4932) );
  OAI21_X1 U5073 ( .B1(n4312), .B2(n4934), .A(n7939), .ZN(n4933) );
  OR2_X1 U5074 ( .A1(n9654), .A2(n5619), .ZN(n5189) );
  INV_X1 U5075 ( .A(n5654), .ZN(n5619) );
  INV_X1 U5076 ( .A(n5697), .ZN(n5620) );
  AND4_X1 U5077 ( .A1(n5316), .A2(n5315), .A3(n5314), .A4(n5313), .ZN(n7209)
         );
  AND2_X1 U5079 ( .A1(n4555), .A2(n9657), .ZN(n4554) );
  OR2_X1 U5080 ( .A1(n4963), .A2(n4556), .ZN(n4555) );
  AOI21_X1 U5081 ( .B1(n6454), .B2(n4542), .A(n4540), .ZN(n4539) );
  NAND2_X1 U5082 ( .A1(n4541), .A2(n6457), .ZN(n4540) );
  AND2_X1 U5083 ( .A1(n9888), .A2(n9359), .ZN(n6451) );
  NOR2_X1 U5084 ( .A1(n4956), .A2(n6448), .ZN(n4955) );
  NOR2_X1 U5085 ( .A1(n9898), .A2(n9361), .ZN(n6448) );
  INV_X1 U5086 ( .A(n6445), .ZN(n4956) );
  NAND2_X1 U5087 ( .A1(n9820), .A2(n4696), .ZN(n4497) );
  OR2_X1 U5088 ( .A1(n7738), .A2(n4697), .ZN(n4694) );
  AND2_X1 U5089 ( .A1(n9908), .A2(n9363), .ZN(n6442) );
  NOR2_X1 U5090 ( .A1(n6440), .A2(n4962), .ZN(n4961) );
  INV_X1 U5091 ( .A(n6437), .ZN(n4962) );
  NAND2_X1 U5092 ( .A1(n5768), .A2(n5767), .ZN(n7131) );
  NAND2_X1 U5093 ( .A1(n10035), .A2(n9630), .ZN(n6799) );
  INV_X1 U5094 ( .A(n8244), .ZN(n9833) );
  NAND2_X1 U5095 ( .A1(n9844), .A2(n9845), .ZN(n4863) );
  AOI21_X1 U5096 ( .B1(n9629), .B2(n10030), .A(n9628), .ZN(n9846) );
  OR2_X1 U5097 ( .A1(n6748), .A2(n6802), .ZN(n10103) );
  AND2_X1 U5098 ( .A1(n5138), .A2(n5137), .ZN(n5180) );
  OR2_X1 U5099 ( .A1(n6676), .A2(P1_U3086), .ZN(n6675) );
  CLKBUF_X1 U5100 ( .A(n6194), .Z(n8558) );
  NAND2_X1 U5101 ( .A1(n6317), .A2(n6316), .ZN(n8611) );
  AOI21_X1 U5102 ( .B1(n4524), .B2(n4519), .A(n4516), .ZN(n4515) );
  OAI21_X1 U5103 ( .B1(n4525), .B2(n8565), .A(n4517), .ZN(n4516) );
  NOR2_X1 U5104 ( .A1(n4521), .A2(n4520), .ZN(n4519) );
  NOR2_X1 U5105 ( .A1(n4518), .A2(n10133), .ZN(n4517) );
  OR2_X1 U5106 ( .A1(n8837), .A2(n8747), .ZN(n4413) );
  OAI211_X1 U5107 ( .C1(n8049), .C2(n8048), .A(n8047), .B(n8046), .ZN(n8053)
         );
  AND2_X1 U5108 ( .A1(n8034), .A2(n8041), .ZN(n8052) );
  AOI21_X1 U5109 ( .B1(n5768), .B2(n4322), .A(n4671), .ZN(n4670) );
  OAI21_X1 U5110 ( .B1(n5285), .B2(n5708), .A(n5770), .ZN(n4671) );
  INV_X1 U5111 ( .A(n8091), .ZN(n4799) );
  INV_X1 U5112 ( .A(n5826), .ZN(n4405) );
  NAND2_X1 U5113 ( .A1(n8191), .A2(n4347), .ZN(n4796) );
  MUX2_X1 U5114 ( .A(n5444), .B(n5443), .S(n5708), .Z(n5462) );
  NAND2_X1 U5115 ( .A1(n4402), .A2(n5778), .ZN(n5443) );
  INV_X1 U5116 ( .A(n8126), .ZN(n4766) );
  INV_X1 U5117 ( .A(n8663), .ZN(n4764) );
  OAI211_X1 U5118 ( .C1(n4655), .C2(n6468), .A(n4652), .B(n4651), .ZN(n4650)
         );
  INV_X1 U5119 ( .A(n5482), .ZN(n4651) );
  NAND2_X1 U5120 ( .A1(n4654), .A2(n4653), .ZN(n4652) );
  NAND2_X1 U5121 ( .A1(n4399), .A2(n4398), .ZN(n5555) );
  AND2_X1 U5122 ( .A1(n9738), .A2(n5718), .ZN(n4398) );
  NAND2_X1 U5123 ( .A1(n5553), .A2(n4400), .ZN(n4399) );
  NOR2_X1 U5124 ( .A1(n4489), .A2(n4401), .ZN(n4400) );
  INV_X1 U5125 ( .A(SI_16_), .ZN(n5076) );
  NOR2_X1 U5126 ( .A1(n4773), .A2(n4771), .ZN(n4768) );
  NOR2_X1 U5127 ( .A1(n8608), .A2(n4774), .ZN(n4773) );
  INV_X1 U5128 ( .A(n8153), .ZN(n4774) );
  MUX2_X1 U5129 ( .A(n8147), .B(n8146), .S(n8165), .Z(n8154) );
  NAND2_X1 U5130 ( .A1(n8597), .A2(n4770), .ZN(n4769) );
  NOR2_X1 U5131 ( .A1(n8624), .A2(n4771), .ZN(n4770) );
  NAND2_X1 U5132 ( .A1(n7093), .A2(n4882), .ZN(n8028) );
  OR2_X1 U5133 ( .A1(n6541), .A2(n7614), .ZN(n6539) );
  INV_X1 U5134 ( .A(n4871), .ZN(n4868) );
  AND2_X1 U5135 ( .A1(n5220), .A2(n5069), .ZN(n5070) );
  INV_X1 U5136 ( .A(SI_14_), .ZN(n5065) );
  NOR2_X1 U5137 ( .A1(n5326), .A2(n4481), .ZN(n4480) );
  OAI21_X1 U5138 ( .B1(n5035), .B2(n4482), .A(n5041), .ZN(n4481) );
  INV_X1 U5139 ( .A(n5040), .ZN(n4877) );
  NAND2_X1 U5140 ( .A1(n6093), .A2(n4820), .ZN(n4819) );
  INV_X1 U5141 ( .A(n4821), .ZN(n4820) );
  XNOR2_X1 U5142 ( .A(n4275), .B(n10189), .ZN(n5955) );
  OR2_X1 U5143 ( .A1(n6635), .A2(n6577), .ZN(n8167) );
  NOR4_X1 U5144 ( .A1(n8697), .A2(n8194), .A3(n8734), .A4(n8193), .ZN(n8196)
         );
  NOR2_X1 U5145 ( .A1(n8823), .A2(n8017), .ZN(n8219) );
  OAI21_X1 U5146 ( .B1(n4295), .B2(n7756), .A(n4841), .ZN(n4840) );
  NAND2_X1 U5147 ( .A1(n4842), .A2(n7406), .ZN(n4841) );
  INV_X1 U5148 ( .A(n7306), .ZN(n4842) );
  INV_X1 U5149 ( .A(n8499), .ZN(n4632) );
  NOR2_X1 U5150 ( .A1(n8482), .A2(n4632), .ZN(n4631) );
  INV_X1 U5151 ( .A(n8510), .ZN(n4513) );
  INV_X1 U5152 ( .A(n8492), .ZN(n4514) );
  INV_X1 U5153 ( .A(n6173), .ZN(n6172) );
  INV_X1 U5154 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n6112) );
  NAND2_X1 U5155 ( .A1(n4900), .A2(n8183), .ZN(n4899) );
  INV_X1 U5156 ( .A(n8041), .ZN(n4900) );
  INV_X1 U5157 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n4587) );
  INV_X1 U5158 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n6025) );
  INV_X1 U5159 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5996) );
  NAND2_X1 U5160 ( .A1(n6521), .A2(n4746), .ZN(n4743) );
  AND2_X1 U5161 ( .A1(n6524), .A2(n6520), .ZN(n4746) );
  OAI21_X1 U5162 ( .B1(n8683), .B2(n6564), .A(n6563), .ZN(n6566) );
  INV_X1 U5163 ( .A(n6562), .ZN(n6563) );
  OR2_X1 U5164 ( .A1(n8866), .A2(n8346), .ZN(n8128) );
  AND2_X1 U5165 ( .A1(n8694), .A2(n8195), .ZN(n8679) );
  AND2_X1 U5166 ( .A1(n8097), .A2(n8098), .ZN(n8191) );
  OR2_X1 U5167 ( .A1(n7636), .A2(n7626), .ZN(n8088) );
  OR2_X1 U5168 ( .A1(n8182), .A2(n7451), .ZN(n7452) );
  NOR2_X1 U5169 ( .A1(n8401), .A2(n10215), .ZN(n4761) );
  INV_X1 U5170 ( .A(n5905), .ZN(n6330) );
  NAND2_X1 U5171 ( .A1(n4460), .A2(n4459), .ZN(n5925) );
  INV_X1 U5172 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n4459) );
  INV_X1 U5173 ( .A(n5923), .ZN(n4460) );
  OAI21_X1 U5174 ( .B1(n6167), .B2(P2_IR_REG_17__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n6179) );
  NOR2_X1 U5175 ( .A1(n6005), .A2(P2_IR_REG_6__SCAN_IN), .ZN(n6018) );
  NAND2_X1 U5176 ( .A1(n4915), .A2(n7816), .ZN(n4914) );
  INV_X1 U5177 ( .A(n4976), .ZN(n4915) );
  AOI211_X1 U5178 ( .C1(n6475), .C2(n5761), .A(n5760), .B(n5759), .ZN(n5842)
         );
  AOI21_X1 U5179 ( .B1(n5762), .B2(n5757), .A(n6473), .ZN(n5758) );
  OAI211_X1 U5180 ( .C1(n4676), .C2(n4301), .A(n4672), .B(n4678), .ZN(n5666)
         );
  INV_X1 U5181 ( .A(n4673), .ZN(n4672) );
  OAI21_X1 U5182 ( .B1(n5645), .B2(n4683), .A(n4679), .ZN(n4678) );
  AOI211_X1 U5183 ( .C1(n5704), .C2(n5708), .A(n5716), .B(n5703), .ZN(n5706)
         );
  OR2_X1 U5184 ( .A1(n4868), .A2(n4493), .ZN(n4492) );
  NAND2_X1 U5185 ( .A1(n4494), .A2(n4990), .ZN(n4493) );
  INV_X1 U5186 ( .A(n4991), .ZN(n4494) );
  OR2_X1 U5187 ( .A1(n4868), .A2(n4496), .ZN(n4495) );
  INV_X1 U5188 ( .A(n4990), .ZN(n4496) );
  NOR2_X1 U5189 ( .A1(n5618), .A2(n9331), .ZN(n5164) );
  NOR2_X1 U5190 ( .A1(n9873), .A2(n9869), .ZN(n4862) );
  AND2_X1 U5191 ( .A1(n4862), .A2(n9680), .ZN(n4861) );
  NAND2_X1 U5192 ( .A1(n4542), .A2(n4543), .ZN(n4541) );
  INV_X1 U5193 ( .A(n9778), .ZN(n4488) );
  OR2_X1 U5194 ( .A1(n9908), .A2(n9231), .ZN(n5719) );
  NAND2_X1 U5195 ( .A1(n9219), .A2(n10072), .ZN(n5770) );
  NAND2_X1 U5196 ( .A1(n9374), .A2(n7141), .ZN(n5726) );
  NAND2_X1 U5197 ( .A1(n9908), .A2(n9231), .ZN(n9801) );
  OR2_X1 U5198 ( .A1(n7206), .A2(n4691), .ZN(n5776) );
  INV_X1 U5199 ( .A(n5773), .ZN(n4692) );
  OR2_X1 U5200 ( .A1(n6468), .A2(n6796), .ZN(n6989) );
  AND2_X1 U5201 ( .A1(n5126), .A2(n5125), .ZN(n5611) );
  INV_X1 U5202 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n5110) );
  NAND2_X1 U5203 ( .A1(n5098), .A2(n4729), .ZN(n4728) );
  NOR2_X1 U5204 ( .A1(n5105), .A2(n4730), .ZN(n4729) );
  INV_X1 U5205 ( .A(n5097), .ZN(n4730) );
  INV_X1 U5206 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n5001) );
  INV_X1 U5207 ( .A(SI_15_), .ZN(n5191) );
  NAND2_X1 U5208 ( .A1(n4506), .A2(n4715), .ZN(n5446) );
  AOI21_X1 U5209 ( .B1(n4717), .B2(n4297), .A(n4355), .ZN(n4715) );
  OAI211_X1 U5210 ( .C1(n5354), .C2(n4498), .A(n4503), .B(n4716), .ZN(n4506)
         );
  AOI21_X1 U5211 ( .B1(n4719), .B2(n4721), .A(n4718), .ZN(n4717) );
  INV_X1 U5212 ( .A(n5060), .ZN(n4718) );
  INV_X1 U5213 ( .A(n4724), .ZN(n4719) );
  NAND2_X1 U5214 ( .A1(n5318), .A2(n5035), .ZN(n4707) );
  NAND2_X1 U5215 ( .A1(n4428), .A2(n6037), .ZN(n7284) );
  XNOR2_X1 U5216 ( .A(n6283), .B(n6552), .ZN(n8309) );
  OAI21_X1 U5217 ( .B1(n8330), .B2(n4357), .A(n4300), .ZN(n4429) );
  INV_X1 U5218 ( .A(n8399), .ZN(n8322) );
  INV_X1 U5219 ( .A(n8382), .ZN(n8356) );
  NAND2_X1 U5220 ( .A1(n4431), .A2(n4430), .ZN(n8352) );
  INV_X1 U5221 ( .A(n8355), .ZN(n4430) );
  NAND2_X1 U5222 ( .A1(n6139), .A2(n6138), .ZN(n7789) );
  INV_X1 U5223 ( .A(n8231), .ZN(n4788) );
  XNOR2_X1 U5224 ( .A(n5916), .B(P2_IR_REG_19__SCAN_IN), .ZN(n6194) );
  NAND2_X1 U5225 ( .A1(n6181), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5916) );
  INV_X1 U5226 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5893) );
  NOR2_X1 U5227 ( .A1(n4807), .A2(n4808), .ZN(n5912) );
  NOR2_X1 U5228 ( .A1(n4785), .A2(n4786), .ZN(n4782) );
  NOR2_X1 U5229 ( .A1(n4787), .A2(n8573), .ZN(n4786) );
  INV_X1 U5230 ( .A(n4978), .ZN(n4787) );
  AND4_X1 U5231 ( .A1(n6119), .A2(n6118), .A3(n6117), .A4(n6116), .ZN(n7793)
         );
  AND4_X1 U5232 ( .A1(n6033), .A2(n6032), .A3(n6031), .A4(n6030), .ZN(n6531)
         );
  XNOR2_X1 U5233 ( .A(n6872), .B(n6871), .ZN(n6755) );
  OAI21_X1 U5234 ( .B1(n8564), .B2(n4438), .A(n4437), .ZN(n6872) );
  NAND2_X1 U5235 ( .A1(n8564), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n4437) );
  NAND2_X1 U5236 ( .A1(n4509), .A2(n6950), .ZN(n10149) );
  XNOR2_X1 U5237 ( .A(n7265), .B(n7271), .ZN(n7263) );
  AND2_X1 U5238 ( .A1(n7270), .A2(n7271), .ZN(n4618) );
  OAI22_X1 U5239 ( .A1(n7531), .A2(n7530), .B1(n7529), .B2(n7528), .ZN(n7702)
         );
  NAND2_X1 U5240 ( .A1(n4462), .A2(n8438), .ZN(n8416) );
  NAND2_X1 U5241 ( .A1(n8409), .A2(n8408), .ZN(n8435) );
  OAI21_X1 U5242 ( .B1(n8481), .B2(n4632), .A(n4630), .ZN(n4629) );
  INV_X1 U5243 ( .A(n8498), .ZN(n4630) );
  INV_X1 U5244 ( .A(n4631), .ZN(n4627) );
  OAI21_X1 U5245 ( .B1(n8483), .B2(n8482), .A(n8481), .ZN(n8500) );
  INV_X1 U5246 ( .A(n4629), .ZN(n4628) );
  NAND2_X1 U5247 ( .A1(n4302), .A2(n8519), .ZN(n4625) );
  NAND2_X1 U5248 ( .A1(n8246), .A2(n6322), .ZN(n8594) );
  NOR2_X1 U5249 ( .A1(n8134), .A2(n4894), .ZN(n4893) );
  INV_X1 U5250 ( .A(n4893), .ZN(n4890) );
  NAND2_X1 U5251 ( .A1(n6552), .A2(n8357), .ZN(n6557) );
  OR2_X1 U5252 ( .A1(n6162), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n6173) );
  OR2_X1 U5253 ( .A1(n6074), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n6076) );
  NAND2_X1 U5254 ( .A1(n4743), .A2(n4745), .ZN(n6527) );
  NAND2_X1 U5255 ( .A1(n8751), .A2(n8031), .ZN(n6521) );
  INV_X1 U5256 ( .A(n8159), .ZN(n4880) );
  NAND2_X1 U5257 ( .A1(n6622), .A2(n10178), .ZN(n4577) );
  OAI21_X1 U5258 ( .B1(n8610), .B2(n4741), .A(n4739), .ZN(n8587) );
  NAND2_X1 U5259 ( .A1(n8588), .A2(n10173), .ZN(n8590) );
  NAND2_X1 U5260 ( .A1(n6566), .A2(n8199), .ZN(n8649) );
  NAND2_X1 U5261 ( .A1(n4754), .A2(n4346), .ZN(n4753) );
  AND2_X1 U5262 ( .A1(n6556), .A2(n6559), .ZN(n4752) );
  OR2_X1 U5263 ( .A1(n8803), .A2(n8313), .ZN(n8694) );
  INV_X1 U5264 ( .A(n8679), .ZN(n8708) );
  NAND2_X1 U5265 ( .A1(n4756), .A2(n6556), .ZN(n8722) );
  OR2_X1 U5266 ( .A1(n6553), .A2(n8300), .ZN(n8111) );
  AND2_X1 U5267 ( .A1(n4311), .A2(n8677), .ZN(n8721) );
  INV_X1 U5268 ( .A(n8191), .ZN(n7983) );
  AND2_X1 U5269 ( .A1(n8056), .A2(n8067), .ZN(n8182) );
  OR2_X1 U5270 ( .A1(n5958), .A2(n6659), .ZN(n5911) );
  OR2_X1 U5271 ( .A1(n8756), .A2(n4391), .ZN(n10201) );
  NAND2_X1 U5272 ( .A1(n6342), .A2(n6343), .ZN(n6695) );
  NAND2_X1 U5273 ( .A1(n4801), .A2(n4800), .ZN(n5931) );
  AOI21_X1 U5274 ( .B1(n4802), .B2(n5900), .A(n4362), .ZN(n4801) );
  NAND2_X1 U5275 ( .A1(n5905), .A2(n4802), .ZN(n4800) );
  AND2_X1 U5276 ( .A1(n6018), .A2(n4284), .ZN(n6156) );
  AND2_X1 U5277 ( .A1(n6143), .A2(n6129), .ZN(n8467) );
  INV_X1 U5278 ( .A(n6764), .ZN(n4536) );
  NOR2_X1 U5279 ( .A1(n4327), .A2(n4935), .ZN(n4934) );
  INV_X1 U5280 ( .A(n7926), .ZN(n4935) );
  INV_X1 U5281 ( .A(n9355), .ZN(n9095) );
  NAND2_X1 U5282 ( .A1(n4475), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n5416) );
  INV_X1 U5283 ( .A(n5414), .ZN(n4475) );
  AOI21_X1 U5284 ( .B1(n4354), .B2(n7853), .A(n4600), .ZN(n4599) );
  INV_X1 U5285 ( .A(n9182), .ZN(n4600) );
  INV_X1 U5286 ( .A(n7853), .ZN(n4601) );
  NAND2_X1 U5287 ( .A1(n4448), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n5429) );
  INV_X1 U5288 ( .A(n5416), .ZN(n4448) );
  INV_X1 U5289 ( .A(n9374), .ZN(n9219) );
  NAND2_X1 U5290 ( .A1(n4446), .A2(n5160), .ZN(n5478) );
  AND2_X1 U5291 ( .A1(P1_REG3_REG_15__SCAN_IN), .A2(P1_REG3_REG_16__SCAN_IN), 
        .ZN(n5160) );
  INV_X1 U5292 ( .A(n5231), .ZN(n4446) );
  AND2_X1 U5293 ( .A1(n7950), .A2(n7948), .ZN(n9237) );
  NAND2_X1 U5294 ( .A1(n4922), .A2(n4926), .ZN(n4919) );
  INV_X1 U5295 ( .A(n7950), .ZN(n4917) );
  INV_X1 U5296 ( .A(n9354), .ZN(n9328) );
  NAND2_X1 U5297 ( .A1(n4356), .A2(n9836), .ZN(n4445) );
  INV_X1 U5298 ( .A(n5851), .ZN(n5881) );
  NOR2_X1 U5299 ( .A1(n4735), .A2(n8242), .ZN(n5851) );
  INV_X1 U5300 ( .A(n4469), .ZN(n6796) );
  AND2_X1 U5301 ( .A1(n5588), .A2(n5587), .ZN(n9286) );
  OAI21_X1 U5302 ( .B1(n5310), .B2(n5254), .A(n4687), .ZN(n4686) );
  OR2_X1 U5303 ( .A1(n5310), .A2(n5270), .ZN(n4937) );
  INV_X1 U5304 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5224) );
  NAND2_X1 U5305 ( .A1(n9572), .A2(n9573), .ZN(n9588) );
  XNOR2_X1 U5306 ( .A(n9616), .B(P1_REG3_REG_28__SCAN_IN), .ZN(n9639) );
  NAND2_X1 U5307 ( .A1(n9666), .A2(n9665), .ZN(n4706) );
  INV_X1 U5308 ( .A(n4873), .ZN(n9666) );
  NAND2_X1 U5309 ( .A1(n4873), .A2(n4872), .ZN(n4874) );
  AND2_X1 U5310 ( .A1(n5717), .A2(n9690), .ZN(n9713) );
  INV_X1 U5311 ( .A(n6455), .ZN(n4545) );
  NAND2_X1 U5312 ( .A1(n6470), .A2(n6469), .ZN(n9729) );
  OR2_X1 U5313 ( .A1(n9888), .A2(n9123), .ZN(n9738) );
  AOI21_X1 U5314 ( .B1(n4952), .B2(n4954), .A(n4350), .ZN(n4950) );
  AOI21_X1 U5315 ( .B1(n4697), .B2(n4294), .A(n4318), .ZN(n4490) );
  AOI21_X1 U5316 ( .B1(n4570), .B2(n4569), .A(n4319), .ZN(n4568) );
  NAND2_X1 U5317 ( .A1(n7575), .A2(n5781), .ZN(n7738) );
  OR2_X1 U5318 ( .A1(n9299), .A2(n7834), .ZN(n7417) );
  OR2_X1 U5319 ( .A1(n4857), .A2(n9368), .ZN(n4571) );
  NAND2_X1 U5320 ( .A1(n4292), .A2(n7344), .ZN(n4942) );
  AND2_X1 U5321 ( .A1(n4292), .A2(n4947), .ZN(n4943) );
  NAND2_X1 U5322 ( .A1(n9157), .A2(n9069), .ZN(n7322) );
  NAND2_X1 U5323 ( .A1(n7209), .A2(n5341), .ZN(n6426) );
  AND2_X1 U5324 ( .A1(n5771), .A2(n5819), .ZN(n10015) );
  NAND2_X1 U5325 ( .A1(n5769), .A2(n7128), .ZN(n7133) );
  NAND2_X1 U5326 ( .A1(n7129), .A2(n5725), .ZN(n7027) );
  AND3_X1 U5327 ( .A1(n4646), .A2(n5253), .A3(n4643), .ZN(n6420) );
  NAND2_X1 U5328 ( .A1(n5613), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n4646) );
  NAND2_X1 U5329 ( .A1(n4645), .A2(n4644), .ZN(n4643) );
  NOR2_X1 U5330 ( .A1(n9377), .A2(n6991), .ZN(n6993) );
  NAND2_X1 U5331 ( .A1(n9377), .A2(n6986), .ZN(n6990) );
  INV_X1 U5332 ( .A(n9329), .ZN(n9304) );
  AOI21_X1 U5333 ( .B1(n6481), .B2(n10030), .A(n9138), .ZN(n9641) );
  INV_X1 U5334 ( .A(n9849), .ZN(n9852) );
  NAND2_X1 U5335 ( .A1(n5561), .A2(n5560), .ZN(n9878) );
  NAND2_X1 U5336 ( .A1(n5229), .A2(n5228), .ZN(n5461) );
  INV_X1 U5337 ( .A(n10103), .ZN(n10084) );
  NAND4_X1 U5338 ( .A1(n6976), .A2(n6502), .A3(n6501), .A4(n6799), .ZN(n7001)
         );
  INV_X1 U5339 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n4700) );
  XNOR2_X1 U5340 ( .A(n5693), .B(n5692), .ZN(n8252) );
  NAND2_X1 U5341 ( .A1(n5689), .A2(n5688), .ZN(n5693) );
  XNOR2_X1 U5342 ( .A(n5684), .B(n5651), .ZN(n8904) );
  OR2_X1 U5343 ( .A1(n5860), .A2(n5859), .ZN(n5866) );
  NAND2_X1 U5344 ( .A1(n4728), .A2(n4726), .ZN(n5573) );
  NOR2_X1 U5345 ( .A1(n5558), .A2(n4727), .ZN(n4726) );
  INV_X1 U5346 ( .A(n5104), .ZN(n4727) );
  INV_X1 U5347 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n5489) );
  OR2_X1 U5348 ( .A1(n5410), .A2(P1_IR_REG_11__SCAN_IN), .ZN(n5424) );
  NAND2_X1 U5349 ( .A1(n4723), .A2(n5055), .ZN(n4442) );
  NAND2_X1 U5350 ( .A1(n5053), .A2(n4724), .ZN(n4723) );
  XNOR2_X1 U5351 ( .A(n5407), .B(n5406), .ZN(n6712) );
  NAND2_X1 U5352 ( .A1(n6506), .A2(n6505), .ZN(n6507) );
  NAND2_X1 U5353 ( .A1(n6863), .A2(n6862), .ZN(n6861) );
  AND2_X1 U5354 ( .A1(n6246), .A2(n6245), .ZN(n8621) );
  AND2_X1 U5355 ( .A1(n4824), .A2(n6407), .ZN(n4822) );
  AND2_X1 U5357 ( .A1(n6204), .A2(n6203), .ZN(n8707) );
  INV_X1 U5358 ( .A(n8225), .ZN(n4789) );
  OR2_X1 U5359 ( .A1(n8019), .A2(n4449), .ZN(n4780) );
  NAND2_X1 U5360 ( .A1(n6224), .A2(n6223), .ZN(n8671) );
  INV_X1 U5361 ( .A(n8313), .ZN(n8725) );
  AND3_X1 U5362 ( .A1(n6177), .A2(n6176), .A3(n6175), .ZN(n8740) );
  INV_X1 U5363 ( .A(n7793), .ZN(n8394) );
  INV_X1 U5364 ( .A(n6531), .ZN(n8400) );
  AOI21_X1 U5365 ( .B1(n10147), .B2(n4614), .A(n4612), .ZN(n4611) );
  INV_X1 U5366 ( .A(n6958), .ZN(n4612) );
  NOR2_X1 U5367 ( .A1(n7070), .A2(n7071), .ZN(n7173) );
  XNOR2_X1 U5368 ( .A(n8435), .B(n8438), .ZN(n8436) );
  AOI21_X1 U5369 ( .B1(n8543), .B2(P2_REG2_REG_17__SCAN_IN), .A(n4527), .ZN(
        n8555) );
  INV_X1 U5370 ( .A(n10133), .ZN(n10160) );
  NAND2_X1 U5371 ( .A1(n4435), .A2(n4523), .ZN(n4434) );
  OR2_X1 U5372 ( .A1(n8538), .A2(n8570), .ZN(n4435) );
  NAND2_X1 U5373 ( .A1(n8539), .A2(n8562), .ZN(n4436) );
  INV_X1 U5374 ( .A(n8575), .ZN(n4616) );
  NAND2_X1 U5375 ( .A1(n8543), .A2(n4394), .ZN(n4524) );
  INV_X1 U5376 ( .A(n4577), .ZN(n4578) );
  NAND2_X1 U5377 ( .A1(n6282), .A2(n6281), .ZN(n8840) );
  NAND2_X1 U5378 ( .A1(n8659), .A2(n8658), .ZN(n8788) );
  NAND2_X1 U5379 ( .A1(n6213), .A2(n6212), .ZN(n8787) );
  INV_X1 U5380 ( .A(n8581), .ZN(n10181) );
  NAND2_X1 U5381 ( .A1(n10186), .A2(n6901), .ZN(n8747) );
  NAND2_X1 U5382 ( .A1(n6648), .A2(n6696), .ZN(n8655) );
  NAND2_X1 U5383 ( .A1(n6308), .A2(n6307), .ZN(n8834) );
  OR2_X1 U5384 ( .A1(n8837), .A2(n8813), .ZN(n4412) );
  NAND2_X1 U5385 ( .A1(n10229), .A2(n10216), .ZN(n8780) );
  NOR2_X1 U5386 ( .A1(n8006), .A2(n8005), .ZN(n8819) );
  OR2_X1 U5387 ( .A1(n8837), .A2(n8896), .ZN(n4414) );
  OAI21_X1 U5388 ( .B1(n8620), .B2(n8737), .A(n4473), .ZN(n4472) );
  NAND2_X1 U5389 ( .A1(n8601), .A2(n10173), .ZN(n4473) );
  AOI21_X1 U5390 ( .B1(n4427), .B2(n10178), .A(n4424), .ZN(n8838) );
  NAND2_X1 U5391 ( .A1(n4426), .A2(n4425), .ZN(n4424) );
  NAND2_X1 U5392 ( .A1(n8611), .A2(n10173), .ZN(n4425) );
  NAND2_X1 U5393 ( .A1(n6238), .A2(n6237), .ZN(n8853) );
  NAND2_X1 U5394 ( .A1(n6251), .A2(n6250), .ZN(n8859) );
  OR2_X1 U5395 ( .A1(n10219), .A2(n10210), .ZN(n8896) );
  INV_X1 U5396 ( .A(n8845), .ZN(n8893) );
  XNOR2_X1 U5397 ( .A(n5748), .B(n5747), .ZN(n6676) );
  NAND2_X1 U5398 ( .A1(n5746), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5748) );
  NAND2_X1 U5399 ( .A1(n5182), .A2(n5181), .ZN(n9850) );
  NAND2_X1 U5400 ( .A1(n5153), .A2(n5152), .ZN(n9636) );
  AND2_X1 U5401 ( .A1(n7917), .A2(n9171), .ZN(n7918) );
  INV_X1 U5402 ( .A(n7478), .ZN(n4857) );
  INV_X1 U5403 ( .A(n9343), .ZN(n9332) );
  AND2_X1 U5404 ( .A1(n6803), .A2(n6795), .ZN(n9326) );
  NAND2_X1 U5405 ( .A1(n6803), .A2(n6802), .ZN(n9345) );
  NAND2_X1 U5406 ( .A1(n5568), .A2(n5567), .ZN(n9357) );
  INV_X1 U5407 ( .A(n7834), .ZN(n9368) );
  XNOR2_X1 U5408 ( .A(n6823), .B(P1_REG2_REG_1__SCAN_IN), .ZN(n9385) );
  NAND2_X1 U5409 ( .A1(n9459), .A2(n9460), .ZN(n9458) );
  NOR2_X1 U5410 ( .A1(n9524), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n4636) );
  NAND2_X1 U5411 ( .A1(n9537), .A2(n9536), .ZN(n9561) );
  AOI21_X1 U5412 ( .B1(n9600), .B2(n9966), .A(n4395), .ZN(n4640) );
  OAI21_X1 U5413 ( .B1(n9995), .B2(n9603), .A(n9602), .ZN(n4638) );
  INV_X1 U5414 ( .A(n9986), .ZN(n9598) );
  OR2_X1 U5415 ( .A1(n8235), .A2(n9833), .ZN(n8238) );
  NAND2_X1 U5416 ( .A1(n4550), .A2(n4554), .ZN(n4970) );
  NAND2_X1 U5417 ( .A1(n4964), .A2(n4963), .ZN(n4553) );
  NAND2_X1 U5418 ( .A1(n5494), .A2(n5493), .ZN(n9898) );
  INV_X1 U5419 ( .A(n6420), .ZN(n4833) );
  INV_X1 U5420 ( .A(n9806), .ZN(n10041) );
  OR2_X1 U5421 ( .A1(n6800), .A2(n6799), .ZN(n9806) );
  NAND2_X1 U5422 ( .A1(n6985), .A2(n9806), .ZN(n9996) );
  NAND2_X1 U5423 ( .A1(n9846), .A2(n4299), .ZN(n9934) );
  AND2_X1 U5424 ( .A1(n9843), .A2(n9842), .ZN(n4575) );
  NOR2_X1 U5425 ( .A1(n7668), .A2(n7667), .ZN(n10243) );
  NAND2_X1 U5426 ( .A1(n4410), .A2(n4409), .ZN(n4408) );
  AOI21_X1 U5427 ( .B1(n8025), .B2(n8165), .A(n8031), .ZN(n4409) );
  NAND2_X1 U5428 ( .A1(n8026), .A2(n8158), .ZN(n4410) );
  MUX2_X1 U5429 ( .A(n8055), .B(n8054), .S(n8158), .Z(n8060) );
  NOR2_X1 U5430 ( .A1(n4670), .A2(n5298), .ZN(n5301) );
  NAND2_X1 U5431 ( .A1(n4664), .A2(n4665), .ZN(n4657) );
  OR2_X1 U5432 ( .A1(n4296), .A2(n5387), .ZN(n4664) );
  AND2_X1 U5433 ( .A1(n4660), .A2(n4663), .ZN(n4658) );
  NAND2_X1 U5434 ( .A1(n4385), .A2(n6429), .ZN(n4663) );
  NOR2_X1 U5435 ( .A1(n4661), .A2(n4668), .ZN(n4660) );
  NOR2_X1 U5436 ( .A1(n5387), .A2(n4662), .ZN(n4661) );
  NAND2_X1 U5437 ( .A1(n4669), .A2(n5386), .ZN(n4668) );
  AND2_X1 U5438 ( .A1(n6431), .A2(n6468), .ZN(n4669) );
  NOR2_X1 U5439 ( .A1(n4296), .A2(n4667), .ZN(n4666) );
  INV_X1 U5440 ( .A(n5771), .ZN(n4667) );
  AND2_X1 U5441 ( .A1(n4799), .A2(n8158), .ZN(n4791) );
  AOI21_X1 U5442 ( .B1(n8084), .B2(n8078), .A(n8077), .ZN(n8086) );
  NOR2_X1 U5443 ( .A1(n8091), .A2(n8158), .ZN(n4795) );
  NOR2_X1 U5444 ( .A1(n4405), .A2(n4404), .ZN(n4403) );
  INV_X1 U5445 ( .A(n5722), .ZN(n4404) );
  NAND2_X1 U5446 ( .A1(n5464), .A2(n5779), .ZN(n4654) );
  AND2_X1 U5447 ( .A1(n5465), .A2(n6468), .ZN(n4653) );
  INV_X1 U5448 ( .A(n5839), .ZN(n4401) );
  NAND2_X1 U5449 ( .A1(n10027), .A2(n5812), .ZN(n5297) );
  NOR2_X1 U5450 ( .A1(n8131), .A2(n8199), .ZN(n4765) );
  NAND2_X1 U5451 ( .A1(n4766), .A2(n4764), .ZN(n4763) );
  NOR2_X1 U5452 ( .A1(n8170), .A2(n4407), .ZN(n4406) );
  MUX2_X1 U5453 ( .A(n5557), .B(n5556), .S(n5708), .Z(n5571) );
  OR2_X1 U5454 ( .A1(n5468), .A2(n5236), .ZN(n5830) );
  INV_X1 U5455 ( .A(n8267), .ZN(n4827) );
  NOR4_X1 U5456 ( .A1(n8180), .A2(n8179), .A3(n8178), .A4(n10171), .ZN(n8181)
         );
  NOR2_X1 U5457 ( .A1(n4336), .A2(n6572), .ZN(n4742) );
  INV_X1 U5458 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5904) );
  NOR4_X1 U5459 ( .A1(n7342), .A2(n5823), .A3(n5772), .A4(n5730), .ZN(n5731)
         );
  OR4_X1 U5460 ( .A1(n5729), .A2(n4662), .A3(n10020), .A4(n5773), .ZN(n5730)
         );
  AND2_X1 U5461 ( .A1(n9778), .A2(n9820), .ZN(n4478) );
  NAND2_X1 U5462 ( .A1(n5636), .A2(n5790), .ZN(n4683) );
  INV_X1 U5463 ( .A(n4682), .ZN(n4679) );
  OR2_X1 U5464 ( .A1(n5637), .A2(n4682), .ZN(n4681) );
  AND2_X1 U5465 ( .A1(n6471), .A2(n6474), .ZN(n4871) );
  NAND2_X1 U5466 ( .A1(n7244), .A2(n7322), .ZN(n5773) );
  INV_X1 U5467 ( .A(n5138), .ZN(n4714) );
  INV_X1 U5468 ( .A(n4713), .ZN(n4712) );
  OAI21_X1 U5469 ( .B1(n5180), .B2(n4714), .A(n5647), .ZN(n4713) );
  INV_X1 U5470 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5004) );
  INV_X1 U5471 ( .A(SI_19_), .ZN(n5086) );
  AND2_X1 U5472 ( .A1(n4717), .A2(n5422), .ZN(n4716) );
  NOR2_X1 U5473 ( .A1(n5394), .A2(n4722), .ZN(n4721) );
  INV_X1 U5474 ( .A(n5055), .ZN(n4722) );
  INV_X1 U5475 ( .A(SI_11_), .ZN(n5056) );
  NOR2_X1 U5476 ( .A1(n4499), .A2(n4505), .ZN(n4504) );
  INV_X1 U5477 ( .A(n4979), .ZN(n4505) );
  INV_X1 U5478 ( .A(n5353), .ZN(n4501) );
  AND2_X1 U5479 ( .A1(n8319), .A2(n6050), .ZN(n4821) );
  NAND2_X1 U5480 ( .A1(n4768), .A2(n8597), .ZN(n4767) );
  NAND4_X1 U5481 ( .A1(n5938), .A2(n5937), .A3(n5936), .A4(n5935), .ZN(n6515)
         );
  OR2_X1 U5482 ( .A1(n4271), .A2(n5932), .ZN(n5937) );
  NAND2_X1 U5483 ( .A1(n4523), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n4522) );
  NAND2_X1 U5484 ( .A1(n6272), .A2(n4579), .ZN(n6321) );
  AND2_X1 U5485 ( .A1(n4306), .A2(n6309), .ZN(n4579) );
  INV_X1 U5486 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n4590) );
  INV_X1 U5487 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n6171) );
  AND2_X1 U5488 ( .A1(n4745), .A2(n7162), .ZN(n4744) );
  AND2_X1 U5489 ( .A1(n6345), .A2(n6697), .ZN(n6645) );
  AND2_X1 U5490 ( .A1(n6344), .A2(n6700), .ZN(n6642) );
  NAND2_X1 U5491 ( .A1(n4738), .A2(n4741), .ZN(n4736) );
  NAND2_X1 U5492 ( .A1(n6559), .A2(n4755), .ZN(n4754) );
  INV_X1 U5493 ( .A(n6557), .ZN(n4755) );
  AND2_X1 U5494 ( .A1(n4311), .A2(n8111), .ZN(n4904) );
  NAND2_X1 U5495 ( .A1(n6614), .A2(n8003), .ZN(n5958) );
  AND3_X1 U5496 ( .A1(n6895), .A2(n6894), .A3(n6639), .ZN(n6381) );
  OR2_X1 U5497 ( .A1(n6094), .A2(P2_IR_REG_11__SCAN_IN), .ZN(n6109) );
  OR3_X1 U5498 ( .A1(n6066), .A2(P2_IR_REG_9__SCAN_IN), .A3(
        P2_IR_REG_10__SCAN_IN), .ZN(n6094) );
  INV_X1 U5499 ( .A(n7802), .ZN(n4930) );
  OR2_X1 U5500 ( .A1(n9150), .A2(n9152), .ZN(n4973) );
  NAND2_X1 U5501 ( .A1(n4914), .A2(n7823), .ZN(n4913) );
  NOR2_X1 U5502 ( .A1(n5562), .A2(n9287), .ZN(n4476) );
  INV_X1 U5503 ( .A(n7058), .ZN(n4921) );
  OR2_X1 U5504 ( .A1(n5312), .A2(n5248), .ZN(n5283) );
  OR2_X1 U5505 ( .A1(n5295), .A2(P1_IR_REG_3__SCAN_IN), .ZN(n5327) );
  INV_X1 U5506 ( .A(n6462), .ZN(n4969) );
  INV_X1 U5507 ( .A(n6461), .ZN(n4556) );
  OR2_X1 U5508 ( .A1(n9850), .A2(n9330), .ZN(n5761) );
  OR2_X1 U5509 ( .A1(n9863), .A2(n9328), .ZN(n6474) );
  OR2_X1 U5510 ( .A1(n9882), .A2(n9285), .ZN(n5753) );
  INV_X1 U5511 ( .A(n4316), .ZN(n4954) );
  NOR2_X1 U5512 ( .A1(n5514), .A2(n5513), .ZN(n4451) );
  NOR2_X1 U5513 ( .A1(n5478), .A2(n9233), .ZN(n4477) );
  INV_X1 U5514 ( .A(n5782), .ZN(n4696) );
  NOR2_X1 U5515 ( .A1(n4308), .A2(n4959), .ZN(n4957) );
  AND2_X1 U5516 ( .A1(n9083), .A2(n9365), .ZN(n5780) );
  OR2_X1 U5517 ( .A1(n9914), .A2(n6441), .ZN(n5720) );
  AOI21_X1 U5518 ( .B1(n7438), .B2(n4571), .A(n4567), .ZN(n4566) );
  AND2_X1 U5519 ( .A1(n4324), .A2(n4571), .ZN(n4565) );
  NOR2_X1 U5520 ( .A1(n9928), .A2(n4857), .ZN(n4858) );
  INV_X1 U5521 ( .A(n5678), .ZN(n4645) );
  INV_X1 U5522 ( .A(n6667), .ZN(n4644) );
  NAND2_X1 U5523 ( .A1(n5821), .A2(n5823), .ZN(n4867) );
  AND2_X1 U5524 ( .A1(n4452), .A2(n7239), .ZN(n6797) );
  INV_X1 U5525 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n8945) );
  NAND2_X1 U5526 ( .A1(n5127), .A2(n5126), .ZN(n5602) );
  AND2_X1 U5527 ( .A1(n5132), .A2(n5131), .ZN(n5601) );
  XNOR2_X1 U5528 ( .A(n5715), .B(P1_IR_REG_21__SCAN_IN), .ZN(n5872) );
  NAND2_X1 U5529 ( .A1(n5714), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5715) );
  INV_X1 U5530 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5742) );
  NAND2_X1 U5531 ( .A1(n4733), .A2(n4731), .ZN(n5502) );
  NOR2_X1 U5532 ( .A1(n4734), .A2(n4732), .ZN(n4731) );
  INV_X1 U5533 ( .A(n5071), .ZN(n4732) );
  INV_X1 U5534 ( .A(n4721), .ZN(n4720) );
  INV_X1 U5535 ( .A(n5052), .ZN(n4725) );
  AOI21_X1 U5536 ( .B1(n5041), .B2(n4877), .A(n4353), .ZN(n4876) );
  OAI21_X1 U5537 ( .B1(n4282), .B2(P1_DATAO_REG_2__SCAN_IN), .A(n5025), .ZN(
        n5026) );
  INV_X1 U5538 ( .A(n8398), .ZN(n7767) );
  NAND2_X1 U5539 ( .A1(n4819), .A2(n4818), .ZN(n4817) );
  INV_X1 U5540 ( .A(n6092), .ZN(n4818) );
  NAND2_X1 U5541 ( .A1(n6280), .A2(n8289), .ZN(n8292) );
  NAND2_X1 U5542 ( .A1(n4815), .A2(n8300), .ZN(n4814) );
  NAND3_X1 U5543 ( .A1(n7096), .A2(n5956), .A3(n5966), .ZN(n7003) );
  NAND2_X1 U5544 ( .A1(n8352), .A2(n4829), .ZN(n4828) );
  NOR2_X1 U5545 ( .A1(n8266), .A2(n4830), .ZN(n4829) );
  INV_X1 U5546 ( .A(n6193), .ZN(n4830) );
  INV_X1 U5547 ( .A(n10189), .ZN(n7093) );
  OAI211_X1 U5548 ( .C1(n6295), .C2(n6298), .A(n6297), .B(n6296), .ZN(n8366)
         );
  NAND2_X1 U5549 ( .A1(n8366), .A2(n8620), .ZN(n8365) );
  NOR4_X1 U5550 ( .A1(n8218), .A2(n8586), .A3(n8599), .A4(n8202), .ZN(n8204)
         );
  AOI21_X1 U5551 ( .B1(n8674), .B2(n6323), .A(n6233), .ZN(n8346) );
  AND4_X1 U5552 ( .A1(n6105), .A2(n6104), .A3(n6103), .A4(n6102), .ZN(n7626)
         );
  AND4_X1 U5553 ( .A1(n6073), .A2(n6072), .A3(n6071), .A4(n6070), .ZN(n7565)
         );
  NAND2_X1 U5554 ( .A1(n6024), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n4885) );
  NAND2_X1 U5555 ( .A1(n5969), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n4883) );
  NAND2_X1 U5556 ( .A1(n5995), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n4884) );
  AOI21_X1 U5557 ( .B1(n6954), .B2(n4458), .A(n6953), .ZN(n10141) );
  XNOR2_X1 U5558 ( .A(n6949), .B(n4269), .ZN(n10131) );
  NAND2_X1 U5559 ( .A1(n4510), .A2(n7300), .ZN(n7407) );
  NAND2_X1 U5560 ( .A1(n7307), .A2(n4295), .ZN(n4846) );
  OAI21_X1 U5561 ( .B1(n7307), .B2(n4843), .A(n4839), .ZN(n7397) );
  NOR2_X1 U5562 ( .A1(n7406), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n4843) );
  INV_X1 U5563 ( .A(n4840), .ZN(n4839) );
  NAND2_X1 U5564 ( .A1(n7307), .A2(n7306), .ZN(n4838) );
  OR2_X1 U5565 ( .A1(n4845), .A2(n4844), .ZN(n7401) );
  NAND2_X1 U5566 ( .A1(n4846), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n4845) );
  INV_X1 U5567 ( .A(n7399), .ZN(n4844) );
  AOI21_X1 U5568 ( .B1(n7702), .B2(n7703), .A(n4444), .ZN(n8418) );
  AND2_X1 U5569 ( .A1(n7533), .A2(n7700), .ZN(n4444) );
  NAND2_X1 U5570 ( .A1(n7524), .A2(n7523), .ZN(n7525) );
  INV_X1 U5571 ( .A(n8455), .ZN(n4850) );
  NAND2_X1 U5572 ( .A1(n8471), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n8505) );
  AOI21_X1 U5573 ( .B1(n4302), .B2(n4624), .A(n8521), .ZN(n4623) );
  NOR2_X1 U5574 ( .A1(n4628), .A2(n8520), .ZN(n4624) );
  AOI21_X1 U5575 ( .B1(n8492), .B2(n8477), .A(n4513), .ZN(n4512) );
  NOR2_X1 U5576 ( .A1(n8565), .A2(n4522), .ZN(n4518) );
  INV_X1 U5577 ( .A(n4525), .ZN(n4521) );
  NAND2_X1 U5578 ( .A1(n8565), .A2(n4522), .ZN(n4520) );
  NAND2_X1 U5579 ( .A1(n4527), .A2(n4526), .ZN(n4525) );
  INV_X1 U5580 ( .A(n8554), .ZN(n4526) );
  AND2_X1 U5581 ( .A1(n8149), .A2(n8148), .ZN(n8624) );
  NOR2_X1 U5582 ( .A1(n8170), .A2(n8199), .ZN(n4892) );
  NAND2_X1 U5583 ( .A1(n6240), .A2(n6239), .ZN(n6273) );
  INV_X1 U5584 ( .A(n6254), .ZN(n6240) );
  OR2_X1 U5585 ( .A1(n6230), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6252) );
  OR2_X1 U5586 ( .A1(n6252), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6254) );
  AND2_X1 U5587 ( .A1(n6216), .A2(n6215), .ZN(n6227) );
  NAND2_X1 U5588 ( .A1(n6227), .A2(n6217), .ZN(n6230) );
  INV_X1 U5589 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n6217) );
  NAND2_X1 U5590 ( .A1(n6172), .A2(n4304), .ZN(n6198) );
  NAND2_X1 U5591 ( .A1(n6172), .A2(n6171), .ZN(n6185) );
  AND2_X1 U5592 ( .A1(n4303), .A2(n4584), .ZN(n4583) );
  INV_X1 U5593 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n4584) );
  NAND2_X1 U5594 ( .A1(n6113), .A2(n4303), .ZN(n6149) );
  NAND2_X1 U5595 ( .A1(n6113), .A2(n6112), .ZN(n6132) );
  NAND2_X1 U5596 ( .A1(n6099), .A2(n6098), .ZN(n6114) );
  INV_X1 U5597 ( .A(n6100), .ZN(n6099) );
  OR2_X1 U5598 ( .A1(n6076), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6100) );
  AND2_X1 U5599 ( .A1(n7590), .A2(n7592), .ZN(n8186) );
  AND2_X1 U5600 ( .A1(n8057), .A2(n8068), .ZN(n8184) );
  AND2_X1 U5601 ( .A1(n4897), .A2(n8067), .ZN(n4896) );
  AND2_X1 U5602 ( .A1(n4323), .A2(n6059), .ZN(n4586) );
  INV_X1 U5603 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n6059) );
  NAND2_X1 U5604 ( .A1(n6026), .A2(n4323), .ZN(n6060) );
  NAND2_X1 U5605 ( .A1(n6585), .A2(n8041), .ZN(n7376) );
  NAND2_X1 U5606 ( .A1(n6026), .A2(n6025), .ZN(n6042) );
  INV_X1 U5607 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n4591) );
  NAND2_X1 U5608 ( .A1(n5970), .A2(n5971), .ZN(n5997) );
  AND4_X1 U5609 ( .A1(n5979), .A2(n5978), .A3(n5977), .A4(n5976), .ZN(n7229)
         );
  INV_X1 U5610 ( .A(n8175), .ZN(n7016) );
  NAND2_X1 U5611 ( .A1(n6902), .A2(n6518), .ZN(n8751) );
  NAND2_X1 U5612 ( .A1(n6891), .A2(n6903), .ZN(n6902) );
  NOR2_X1 U5613 ( .A1(n8578), .A2(n8577), .ZN(n8820) );
  AOI21_X1 U5614 ( .B1(n8610), .B2(n6573), .A(n6572), .ZN(n8600) );
  NAND2_X1 U5615 ( .A1(n8612), .A2(n10175), .ZN(n4426) );
  NAND2_X1 U5616 ( .A1(n6270), .A2(n6269), .ZN(n8286) );
  OAI22_X1 U5617 ( .A1(n6566), .A2(n4747), .B1(n4748), .B2(n4977), .ZN(n8629)
         );
  NAND2_X1 U5618 ( .A1(n4751), .A2(n6567), .ZN(n4747) );
  INV_X1 U5619 ( .A(n4749), .ZN(n4748) );
  AND2_X1 U5620 ( .A1(n8122), .A2(n8663), .ZN(n8684) );
  NAND2_X1 U5621 ( .A1(n6146), .A2(n6145), .ZN(n8814) );
  OR2_X1 U5622 ( .A1(n6537), .A2(n8187), .ZN(n7614) );
  NAND2_X1 U5623 ( .A1(n7376), .A2(n8183), .ZN(n7449) );
  NAND2_X1 U5624 ( .A1(n5922), .A2(n7295), .ZN(n8792) );
  OR2_X1 U5625 ( .A1(n6579), .A2(n8172), .ZN(n6625) );
  AND2_X1 U5626 ( .A1(n6377), .A2(n6696), .ZN(n6627) );
  INV_X1 U5627 ( .A(n8792), .ZN(n10216) );
  AND2_X1 U5628 ( .A1(n6716), .A2(n6702), .ZN(n6696) );
  XNOR2_X1 U5629 ( .A(n6341), .B(n6340), .ZN(n6343) );
  NAND2_X1 U5630 ( .A1(n6330), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6339) );
  INV_X1 U5631 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n6333) );
  NAND2_X1 U5632 ( .A1(n6339), .A2(n6333), .ZN(n6335) );
  XNOR2_X1 U5633 ( .A(n5921), .B(n5920), .ZN(n5922) );
  INV_X1 U5634 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n5920) );
  NAND2_X1 U5635 ( .A1(n5925), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5921) );
  AND2_X1 U5636 ( .A1(n5926), .A2(n5925), .ZN(n8205) );
  INV_X1 U5637 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n5914) );
  AND2_X1 U5638 ( .A1(n6021), .A2(n6051), .ZN(n7271) );
  XNOR2_X1 U5639 ( .A(n6006), .B(P2_IR_REG_6__SCAN_IN), .ZN(n7185) );
  XNOR2_X1 U5640 ( .A(n5982), .B(P2_IR_REG_4__SCAN_IN), .ZN(n6964) );
  INV_X1 U5641 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5744) );
  NAND2_X1 U5642 ( .A1(n9239), .A2(n7950), .ZN(n9193) );
  NOR2_X1 U5643 ( .A1(n9226), .A2(n4310), .ZN(n7887) );
  OR2_X1 U5644 ( .A1(n4468), .A2(n4914), .ZN(n9149) );
  NAND2_X1 U5645 ( .A1(n9263), .A2(n4464), .ZN(n9260) );
  AND2_X1 U5646 ( .A1(n9261), .A2(n9262), .ZN(n4464) );
  INV_X1 U5647 ( .A(n7862), .ZN(n4597) );
  INV_X1 U5648 ( .A(n4476), .ZN(n5581) );
  NAND2_X1 U5649 ( .A1(n9172), .A2(n7926), .ZN(n9089) );
  NAND2_X1 U5650 ( .A1(n9089), .A2(n4989), .ZN(n9090) );
  OR2_X1 U5651 ( .A1(n7849), .A2(n7848), .ZN(n9180) );
  NAND2_X1 U5653 ( .A1(n9193), .A2(n9194), .ZN(n9192) );
  OR2_X1 U5654 ( .A1(n8232), .A2(n6794), .ZN(n9626) );
  INV_X1 U5655 ( .A(n9626), .ZN(n9305) );
  OAI21_X1 U5656 ( .B1(n5713), .B2(n5712), .A(n4985), .ZN(n5877) );
  AND2_X1 U5657 ( .A1(n5530), .A2(n5529), .ZN(n9123) );
  AND3_X1 U5658 ( .A1(n5208), .A2(n5207), .A3(n5206), .ZN(n9231) );
  AND4_X1 U5659 ( .A1(n5404), .A2(n5403), .A3(n5402), .A4(n5401), .ZN(n7834)
         );
  AND4_X1 U5660 ( .A1(n5421), .A2(n5420), .A3(n5419), .A4(n5418), .ZN(n7326)
         );
  AND4_X1 U5661 ( .A1(n5368), .A2(n5367), .A3(n5366), .A4(n5365), .ZN(n9069)
         );
  AND4_X1 U5662 ( .A1(n5385), .A2(n5384), .A3(n5383), .A4(n5382), .ZN(n7208)
         );
  AND4_X1 U5663 ( .A1(n5340), .A2(n5339), .A3(n5338), .A4(n5337), .ZN(n9218)
         );
  OAI21_X1 U5664 ( .B1(n9563), .B2(n9562), .A(n9561), .ZN(n9564) );
  INV_X1 U5665 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n9233) );
  NAND2_X1 U5666 ( .A1(n9588), .A2(n4397), .ZN(n9987) );
  OR2_X1 U5667 ( .A1(n9987), .A2(n9988), .ZN(n9984) );
  AND2_X1 U5668 ( .A1(n5790), .A2(n9621), .ZN(n6478) );
  OR2_X1 U5669 ( .A1(n4964), .A2(n4556), .ZN(n4550) );
  OAI21_X1 U5670 ( .B1(n4491), .B2(n4359), .A(n4869), .ZN(n9658) );
  NAND2_X1 U5671 ( .A1(n9665), .A2(n5627), .ZN(n4869) );
  OAI211_X1 U5672 ( .C1(n9729), .C2(n4495), .A(n4317), .B(n4492), .ZN(n4491)
         );
  NOR2_X1 U5673 ( .A1(n4860), .A2(n9859), .ZN(n4859) );
  INV_X1 U5674 ( .A(n4861), .ZN(n4860) );
  INV_X1 U5675 ( .A(n9850), .ZN(n9652) );
  NOR2_X1 U5676 ( .A1(n4298), .A2(n4968), .ZN(n4963) );
  NAND2_X1 U5677 ( .A1(n9706), .A2(n4862), .ZN(n9696) );
  AND2_X1 U5678 ( .A1(n5628), .A2(n6474), .ZN(n9681) );
  NAND2_X1 U5679 ( .A1(n4293), .A2(n6456), .ZN(n4543) );
  NAND2_X1 U5680 ( .A1(n4364), .A2(n4293), .ZN(n4542) );
  NOR2_X1 U5681 ( .A1(n6455), .A2(n4341), .ZN(n4547) );
  OR2_X1 U5682 ( .A1(n6453), .A2(n4549), .ZN(n4548) );
  NAND2_X1 U5683 ( .A1(n9706), .A2(n9711), .ZN(n9695) );
  AND2_X1 U5684 ( .A1(n9712), .A2(n5638), .ZN(n9727) );
  AND2_X1 U5685 ( .A1(n5753), .A2(n5735), .ZN(n9748) );
  NAND2_X1 U5686 ( .A1(n4451), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n5542) );
  INV_X1 U5687 ( .A(n4451), .ZN(n5524) );
  OAI21_X1 U5688 ( .B1(n4695), .B2(n4489), .A(n4487), .ZN(n9776) );
  AND2_X1 U5689 ( .A1(n4486), .A2(n4485), .ZN(n4487) );
  AOI21_X1 U5690 ( .B1(n4318), .B2(n5789), .A(n4488), .ZN(n4485) );
  NOR2_X1 U5691 ( .A1(n9898), .A2(n4853), .ZN(n4852) );
  INV_X1 U5692 ( .A(n4854), .ZN(n4853) );
  NAND2_X1 U5693 ( .A1(n4477), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n5514) );
  INV_X1 U5694 ( .A(n4477), .ZN(n5496) );
  INV_X1 U5695 ( .A(n5784), .ZN(n9802) );
  NAND2_X1 U5696 ( .A1(n7738), .A2(n5782), .ZN(n9819) );
  NAND2_X1 U5697 ( .A1(n9819), .A2(n9820), .ZN(n9818) );
  NAND2_X1 U5698 ( .A1(n7744), .A2(n7748), .ZN(n9812) );
  INV_X1 U5699 ( .A(n5780), .ZN(n7737) );
  AOI21_X1 U5700 ( .B1(n6438), .B2(n4961), .A(n4351), .ZN(n4960) );
  NAND2_X1 U5701 ( .A1(n4447), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n5231) );
  INV_X1 U5702 ( .A(n5454), .ZN(n4447) );
  NAND2_X1 U5703 ( .A1(n7421), .A2(n4698), .ZN(n7571) );
  NOR2_X1 U5704 ( .A1(n7503), .A2(n4699), .ZN(n4698) );
  INV_X1 U5705 ( .A(n5778), .ZN(n4699) );
  OR2_X1 U5706 ( .A1(n9922), .A2(n9366), .ZN(n6437) );
  NAND2_X1 U5707 ( .A1(n7349), .A2(n4858), .ZN(n7505) );
  NAND2_X1 U5708 ( .A1(n7343), .A2(n5822), .ZN(n7419) );
  NAND2_X1 U5709 ( .A1(n4948), .A2(n7827), .ZN(n4947) );
  NOR2_X1 U5710 ( .A1(n7336), .A2(n4940), .ZN(n4946) );
  NOR2_X1 U5711 ( .A1(n7319), .A2(n4309), .ZN(n4940) );
  NAND2_X1 U5712 ( .A1(n4941), .A2(n4309), .ZN(n4944) );
  INV_X1 U5713 ( .A(n7336), .ZN(n4941) );
  NAND2_X1 U5714 ( .A1(n5345), .A2(n5344), .ZN(n5388) );
  NAND2_X1 U5715 ( .A1(n6431), .A2(n7244), .ZN(n9998) );
  NAND2_X1 U5716 ( .A1(n10014), .A2(n10015), .ZN(n4693) );
  NAND3_X1 U5717 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n5334) );
  INV_X1 U5718 ( .A(n4689), .ZN(n4688) );
  OAI21_X1 U5719 ( .B1(n5278), .B2(n4690), .A(n5810), .ZN(n4689) );
  CLKBUF_X1 U5720 ( .A(n5727), .Z(n6994) );
  NAND2_X1 U5721 ( .A1(n5592), .A2(n5591), .ZN(n9869) );
  NAND2_X1 U5722 ( .A1(n6661), .A2(n5694), .ZN(n4560) );
  NAND2_X1 U5723 ( .A1(n6491), .A2(n6490), .ZN(n9952) );
  INV_X1 U5724 ( .A(n7586), .ZN(n6490) );
  AND2_X1 U5725 ( .A1(n6790), .A2(P1_STATE_REG_SCAN_IN), .ZN(n5871) );
  NOR2_X1 U5726 ( .A1(P1_IR_REG_27__SCAN_IN), .A2(P1_IR_REG_26__SCAN_IN), .ZN(
        n4649) );
  NAND2_X1 U5727 ( .A1(n5168), .A2(P1_IR_REG_28__SCAN_IN), .ZN(n4648) );
  NAND2_X1 U5728 ( .A1(n5147), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5148) );
  XNOR2_X1 U5729 ( .A(n5602), .B(n5601), .ZN(n7584) );
  NAND2_X1 U5730 ( .A1(n4314), .A2(n4980), .ZN(n5864) );
  INV_X1 U5731 ( .A(n5866), .ZN(n5862) );
  INV_X1 U5732 ( .A(n4471), .ZN(n6782) );
  NAND2_X1 U5733 ( .A1(n4728), .A2(n5104), .ZN(n5559) );
  INV_X1 U5734 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n4999) );
  XNOR2_X1 U5735 ( .A(n5196), .B(n5195), .ZN(n7125) );
  INV_X1 U5736 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n5211) );
  XNOR2_X1 U5737 ( .A(n5342), .B(n4979), .ZN(n6708) );
  OAI21_X1 U5738 ( .B1(n5354), .B2(n5353), .A(n5047), .ZN(n5342) );
  OR2_X1 U5739 ( .A1(n5355), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n5371) );
  XNOR2_X1 U5740 ( .A(n5369), .B(n5370), .ZN(n6691) );
  OR3_X1 U5741 ( .A1(n7434), .A2(n7521), .A3(n7685), .ZN(n6716) );
  NAND2_X1 U5742 ( .A1(n7196), .A2(n6017), .ZN(n7286) );
  NAND2_X1 U5743 ( .A1(n6123), .A2(n6122), .ZN(n7788) );
  AND2_X1 U5744 ( .A1(n4823), .A2(n4824), .ZN(n8257) );
  NAND2_X1 U5745 ( .A1(n7096), .A2(n5956), .ZN(n7005) );
  NAND2_X1 U5746 ( .A1(n8352), .A2(n6193), .ZN(n8270) );
  AND2_X1 U5747 ( .A1(n6363), .A2(n8367), .ZN(n6364) );
  NAND2_X1 U5748 ( .A1(n4433), .A2(n4432), .ZN(n4470) );
  INV_X1 U5749 ( .A(n5939), .ZN(n4433) );
  AOI21_X1 U5750 ( .B1(n8691), .B2(n6323), .A(n6211), .ZN(n8282) );
  NAND2_X1 U5751 ( .A1(n7146), .A2(n7147), .ZN(n7145) );
  NAND2_X1 U5752 ( .A1(n4813), .A2(n4814), .ZN(n8311) );
  OR2_X1 U5753 ( .A1(n8303), .A2(n6166), .ZN(n4813) );
  NOR2_X1 U5754 ( .A1(n6376), .A2(n6616), .ZN(n8380) );
  CLKBUF_X1 U5755 ( .A(n7621), .Z(n7622) );
  NAND2_X1 U5756 ( .A1(n4810), .A2(n4809), .ZN(n8354) );
  NAND2_X1 U5757 ( .A1(n7145), .A2(n4825), .ZN(n7196) );
  AND2_X1 U5758 ( .A1(n6004), .A2(n7197), .ZN(n4825) );
  AND2_X1 U5759 ( .A1(n7145), .A2(n6004), .ZN(n7198) );
  AND2_X1 U5760 ( .A1(n6279), .A2(n6278), .ZN(n8632) );
  INV_X1 U5761 ( .A(n8362), .ZN(n8389) );
  NAND2_X1 U5762 ( .A1(n6369), .A2(n6616), .ZN(n8382) );
  NAND2_X1 U5763 ( .A1(n7789), .A2(n4337), .ZN(n8378) );
  INV_X1 U5764 ( .A(n6142), .ZN(n4816) );
  NAND2_X1 U5765 ( .A1(n7789), .A2(n6142), .ZN(n8377) );
  INV_X1 U5766 ( .A(n4782), .ZN(n4781) );
  XNOR2_X1 U5767 ( .A(n6358), .B(P2_IR_REG_22__SCAN_IN), .ZN(n8229) );
  NAND2_X1 U5768 ( .A1(n4778), .A2(n4782), .ZN(n4777) );
  NAND2_X1 U5769 ( .A1(n4582), .A2(n6327), .ZN(n8601) );
  NAND2_X1 U5770 ( .A1(n8594), .A2(n6323), .ZN(n4582) );
  INV_X1 U5771 ( .A(n8632), .ZN(n8612) );
  INV_X1 U5772 ( .A(n8631), .ZN(n8651) );
  INV_X1 U5773 ( .A(n8346), .ZN(n8688) );
  INV_X1 U5774 ( .A(n8707), .ZN(n8687) );
  INV_X1 U5775 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n6734) );
  INV_X1 U5776 ( .A(n7626), .ZN(n8395) );
  INV_X1 U5777 ( .A(n7565), .ZN(n8396) );
  INV_X1 U5778 ( .A(P2_U3893), .ZN(n8403) );
  INV_X1 U5779 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n6763) );
  NOR2_X1 U5780 ( .A1(n4440), .A2(n6767), .ZN(n4439) );
  INV_X1 U5781 ( .A(n6872), .ZN(n4440) );
  XNOR2_X1 U5782 ( .A(n6954), .B(n4458), .ZN(n6873) );
  NAND2_X1 U5783 ( .A1(n4610), .A2(n4614), .ZN(n4613) );
  OR2_X1 U5784 ( .A1(n10146), .A2(n10147), .ZN(n4610) );
  XNOR2_X1 U5785 ( .A(n7074), .B(n7069), .ZN(n7072) );
  OAI21_X1 U5786 ( .B1(n4533), .B2(n7072), .A(n4529), .ZN(n7187) );
  INV_X1 U5787 ( .A(n7075), .ZN(n4533) );
  AOI21_X1 U5788 ( .B1(n7075), .B2(n4532), .A(n4531), .ZN(n4529) );
  INV_X1 U5789 ( .A(n7077), .ZN(n4531) );
  NAND2_X1 U5790 ( .A1(n4530), .A2(n7075), .ZN(n7076) );
  NAND2_X1 U5791 ( .A1(n7072), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n4530) );
  NAND2_X1 U5792 ( .A1(n7067), .A2(n4461), .ZN(n7070) );
  OR2_X1 U5793 ( .A1(n7068), .A2(n7069), .ZN(n4461) );
  AND2_X1 U5794 ( .A1(n4620), .A2(n4619), .ZN(n7269) );
  INV_X1 U5795 ( .A(n7175), .ZN(n4619) );
  INV_X1 U5796 ( .A(n4620), .ZN(n7176) );
  NAND2_X1 U5797 ( .A1(n4835), .A2(n7274), .ZN(n4834) );
  XNOR2_X1 U5798 ( .A(n7407), .B(n7394), .ZN(n7405) );
  AND2_X1 U5799 ( .A1(n6724), .A2(n6723), .ZN(n10164) );
  XNOR2_X1 U5800 ( .A(n7525), .B(n7700), .ZN(n7697) );
  NAND2_X1 U5801 ( .A1(n4382), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n8454) );
  NAND2_X1 U5802 ( .A1(n4534), .A2(n4326), .ZN(n8462) );
  NAND2_X1 U5803 ( .A1(n8436), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n4534) );
  XNOR2_X1 U5804 ( .A(n8491), .B(n8479), .ZN(n8490) );
  NAND2_X1 U5805 ( .A1(n6731), .A2(n6730), .ZN(n10170) );
  NOR2_X1 U5806 ( .A1(n8483), .A2(n4627), .ZN(n4626) );
  NAND2_X1 U5807 ( .A1(n4511), .A2(n8492), .ZN(n8511) );
  NAND2_X1 U5808 ( .A1(n8490), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n4511) );
  OAI21_X1 U5809 ( .B1(n8659), .B2(n4890), .A(n4888), .ZN(n8635) );
  AOI21_X1 U5810 ( .B1(n8199), .B2(n4893), .A(n4407), .ZN(n4888) );
  NAND2_X1 U5811 ( .A1(n8722), .A2(n6557), .ZN(n8705) );
  NAND2_X1 U5812 ( .A1(n6184), .A2(n6183), .ZN(n8803) );
  INV_X1 U5813 ( .A(n6527), .ZN(n10172) );
  INV_X1 U5814 ( .A(n6517), .ZN(n6910) );
  AOI21_X1 U5815 ( .B1(n4881), .B2(n4321), .A(n4880), .ZN(n8585) );
  NAND2_X1 U5816 ( .A1(n8010), .A2(n8009), .ZN(n8823) );
  NAND2_X1 U5817 ( .A1(n8611), .A2(n10175), .ZN(n8589) );
  NAND2_X1 U5818 ( .A1(n8649), .A2(n6567), .ZN(n8641) );
  NAND2_X1 U5819 ( .A1(n8788), .A2(n8139), .ZN(n8639) );
  NAND2_X1 U5820 ( .A1(n6208), .A2(n6207), .ZN(n8872) );
  NAND2_X1 U5821 ( .A1(n6197), .A2(n6196), .ZN(n8878) );
  AND2_X1 U5822 ( .A1(n8727), .A2(n8726), .ZN(n8886) );
  NAND2_X1 U5823 ( .A1(n4905), .A2(n8111), .ZN(n8717) );
  NAND2_X1 U5824 ( .A1(n6131), .A2(n6130), .ZN(n7993) );
  AND2_X1 U5825 ( .A1(n7987), .A2(n7986), .ZN(n7994) );
  NAND2_X1 U5826 ( .A1(n6111), .A2(n6110), .ZN(n8093) );
  NAND2_X1 U5827 ( .A1(n6097), .A2(n6096), .ZN(n7636) );
  NAND2_X1 U5828 ( .A1(n4415), .A2(n6068), .ZN(n6536) );
  NAND2_X1 U5829 ( .A1(n6736), .A2(n8007), .ZN(n4415) );
  AND2_X1 U5830 ( .A1(n7456), .A2(n7455), .ZN(n7464) );
  AND2_X1 U5831 ( .A1(n6718), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6702) );
  AND2_X1 U5832 ( .A1(n4907), .A2(n5899), .ZN(n4906) );
  AND2_X1 U5833 ( .A1(n5928), .A2(n4805), .ZN(n4907) );
  INV_X1 U5834 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n7686) );
  INV_X1 U5835 ( .A(n6343), .ZN(n7685) );
  INV_X1 U5836 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n8983) );
  XNOR2_X1 U5837 ( .A(n6332), .B(n6331), .ZN(n7521) );
  INV_X1 U5838 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n6331) );
  NAND2_X1 U5839 ( .A1(n6335), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6332) );
  NAND2_X1 U5840 ( .A1(n6335), .A2(n6334), .ZN(n7434) );
  OR2_X1 U5841 ( .A1(n6339), .A2(n6333), .ZN(n6334) );
  INV_X1 U5842 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n7375) );
  AND2_X1 U5843 ( .A1(n8003), .A2(P2_U3151), .ZN(n8908) );
  INV_X1 U5844 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7297) );
  INV_X1 U5845 ( .A(n8229), .ZN(n7295) );
  INV_X1 U5846 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n8981) );
  INV_X1 U5847 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7220) );
  INV_X1 U5848 ( .A(n8205), .ZN(n8215) );
  INV_X1 U5849 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7195) );
  INV_X1 U5850 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n7222) );
  INV_X1 U5851 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n7167) );
  INV_X1 U5852 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n7092) );
  INV_X1 U5853 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n9000) );
  INV_X1 U5854 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6869) );
  INV_X1 U5855 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6737) );
  INV_X1 U5856 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6711) );
  INV_X1 U5857 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6703) );
  INV_X1 U5858 ( .A(n7271), .ZN(n7264) );
  NAND2_X1 U5859 ( .A1(n5981), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4535) );
  CLKBUF_X1 U5860 ( .A(n6959), .Z(n4458) );
  INV_X1 U5861 ( .A(n4910), .ZN(n4909) );
  OAI211_X1 U5862 ( .C1(n5678), .C2(n9058), .A(n5247), .B(n5246), .ZN(n7043)
         );
  NAND2_X1 U5863 ( .A1(n5512), .A2(n5511), .ZN(n9893) );
  AND2_X1 U5864 ( .A1(n7968), .A2(n7967), .ZN(n9142) );
  OR2_X1 U5865 ( .A1(n9102), .A2(n4601), .ZN(n4595) );
  CLKBUF_X1 U5866 ( .A(n9228), .Z(n9229) );
  CLKBUF_X1 U5867 ( .A(n9101), .Z(n9102) );
  NAND2_X1 U5868 ( .A1(n5523), .A2(n5522), .ZN(n9888) );
  OR2_X1 U5869 ( .A1(n6780), .A2(n7316), .ZN(n9343) );
  INV_X1 U5870 ( .A(n9194), .ZN(n4918) );
  NAND2_X1 U5871 ( .A1(n9194), .A2(n4917), .ZN(n4916) );
  NOR4_X1 U5872 ( .A1(n5801), .A2(n9630), .A3(n4469), .A4(n6675), .ZN(n5802)
         );
  AOI21_X1 U5873 ( .B1(n5800), .B2(n6677), .A(n5799), .ZN(n5801) );
  OAI21_X1 U5874 ( .B1(n5881), .B2(n9788), .A(n5880), .ZN(n5882) );
  AOI21_X1 U5875 ( .B1(n5853), .B2(n5852), .A(n5851), .ZN(n5855) );
  AND2_X1 U5876 ( .A1(n5662), .A2(n5661), .ZN(n7171) );
  NAND2_X1 U5877 ( .A1(n5178), .A2(n5177), .ZN(n9612) );
  NAND2_X1 U5878 ( .A1(n5625), .A2(n5624), .ZN(n9354) );
  OR2_X1 U5879 ( .A1(n9677), .A2(n5619), .ZN(n5625) );
  NAND2_X1 U5880 ( .A1(n5599), .A2(n5598), .ZN(n9355) );
  INV_X1 U5881 ( .A(n9123), .ZN(n9359) );
  INV_X1 U5882 ( .A(n7864), .ZN(n9366) );
  INV_X1 U5883 ( .A(n7326), .ZN(n6436) );
  INV_X1 U5884 ( .A(n7208), .ZN(n9371) );
  INV_X1 U5885 ( .A(n7209), .ZN(n9373) );
  AND2_X1 U5886 ( .A1(n5291), .A2(n5290), .ZN(n5292) );
  INV_X1 U5887 ( .A(n6854), .ZN(n9375) );
  NAND2_X1 U5888 ( .A1(n5309), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n5255) );
  INV_X1 U5889 ( .A(n4686), .ZN(n5257) );
  NAND2_X1 U5890 ( .A1(n5305), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n4938) );
  NAND2_X1 U5891 ( .A1(n5309), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n5271) );
  INV_X2 U5892 ( .A(P1_U3973), .ZN(n9376) );
  XNOR2_X1 U5893 ( .A(n5252), .B(P1_IR_REG_2__SCAN_IN), .ZN(n9401) );
  NAND2_X1 U5894 ( .A1(n9458), .A2(n4342), .ZN(n9472) );
  NAND2_X1 U5895 ( .A1(n9472), .A2(n9473), .ZN(n9471) );
  NOR2_X1 U5896 ( .A1(n7110), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n4635) );
  NAND2_X1 U5897 ( .A1(n9490), .A2(n4634), .ZN(n9506) );
  NAND2_X1 U5898 ( .A1(n9496), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n4634) );
  NAND2_X1 U5899 ( .A1(n9506), .A2(n9505), .ZN(n9504) );
  NAND2_X1 U5900 ( .A1(n9533), .A2(n4387), .ZN(n9537) );
  AND2_X1 U5901 ( .A1(n5227), .A2(n5226), .ZN(n9550) );
  NOR2_X1 U5902 ( .A1(n9971), .A2(n9972), .ZN(n9970) );
  NAND2_X1 U5903 ( .A1(n5696), .A2(n5695), .ZN(n8244) );
  NAND2_X1 U5904 ( .A1(n5653), .A2(n5652), .ZN(n9839) );
  AND2_X1 U5905 ( .A1(n5607), .A2(n5606), .ZN(n9670) );
  NAND2_X1 U5906 ( .A1(n4705), .A2(n10030), .ZN(n4704) );
  NAND2_X1 U5907 ( .A1(n4706), .A2(n4874), .ZN(n4705) );
  INV_X1 U5908 ( .A(n9869), .ZN(n9702) );
  NAND2_X1 U5909 ( .A1(n6453), .A2(n4545), .ZN(n4544) );
  INV_X1 U5910 ( .A(n6454), .ZN(n4546) );
  NAND2_X1 U5911 ( .A1(n4951), .A2(n4316), .ZN(n9769) );
  NAND2_X1 U5912 ( .A1(n6446), .A2(n4955), .ZN(n4951) );
  NAND2_X1 U5913 ( .A1(n4694), .A2(n4294), .ZN(n5787) );
  NOR2_X1 U5914 ( .A1(n6985), .A2(n9630), .ZN(n9826) );
  INV_X1 U5915 ( .A(n5461), .ZN(n9083) );
  NAND2_X1 U5916 ( .A1(n7421), .A2(n5778), .ZN(n7500) );
  OAI21_X1 U5917 ( .B1(n7439), .B2(n7438), .A(n4571), .ZN(n7416) );
  NAND2_X1 U5918 ( .A1(n5413), .A2(n5412), .ZN(n7841) );
  AOI21_X1 U5919 ( .B1(n7248), .B2(n7319), .A(n4309), .ZN(n7335) );
  NAND2_X1 U5920 ( .A1(n6678), .A2(n9965), .ZN(n5277) );
  NOR2_X1 U5921 ( .A1(n7001), .A2(n7000), .ZN(n10115) );
  INV_X1 U5922 ( .A(n10122), .ZN(n10124) );
  INV_X1 U5923 ( .A(n10115), .ZN(n10122) );
  NOR2_X1 U5924 ( .A1(n9854), .A2(n9853), .ZN(n9855) );
  AND2_X1 U5925 ( .A1(n9952), .A2(n9951), .ZN(n10055) );
  XNOR2_X1 U5926 ( .A(n5677), .B(n5676), .ZN(n9960) );
  INV_X1 U5927 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n5170) );
  MUX2_X1 U5928 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5166), .S(
        P1_IR_REG_29__SCAN_IN), .Z(n5167) );
  XNOR2_X1 U5929 ( .A(n5648), .B(n5647), .ZN(n8909) );
  NAND2_X1 U5930 ( .A1(n4711), .A2(n5138), .ZN(n5648) );
  INV_X1 U5931 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7555) );
  OAI21_X1 U5932 ( .B1(n5578), .B2(n5577), .A(n5576), .ZN(n7372) );
  INV_X1 U5933 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n9026) );
  INV_X1 U5934 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7241) );
  INV_X1 U5935 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7225) );
  AND2_X1 U5936 ( .A1(n5492), .A2(n5491), .ZN(n9991) );
  INV_X1 U5937 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n7049) );
  INV_X1 U5938 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n7013) );
  INV_X1 U5939 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6739) );
  INV_X1 U5940 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n6709) );
  NAND2_X1 U5941 ( .A1(n5168), .A2(n4642), .ZN(n4641) );
  INV_X1 U5942 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n4642) );
  NOR2_X1 U5943 ( .A1(n7666), .A2(n7665), .ZN(n10245) );
  NOR2_X1 U5944 ( .A1(n7670), .A2(n7669), .ZN(n10241) );
  NAND2_X1 U5945 ( .A1(n6507), .A2(n8367), .ZN(n6513) );
  OR2_X1 U5946 ( .A1(n6415), .A2(n6414), .ZN(P2_U3169) );
  NAND2_X1 U5947 ( .A1(n4436), .A2(n4434), .ZN(n8553) );
  NAND2_X1 U5948 ( .A1(n8571), .A2(n10166), .ZN(n4617) );
  OAI21_X1 U5949 ( .B1(n8565), .B2(n4524), .A(n4515), .ZN(n4528) );
  NAND2_X1 U5950 ( .A1(n4419), .A2(n8251), .ZN(P2_U3204) );
  OAI21_X1 U5951 ( .B1(n4578), .B2(n6621), .A(n10186), .ZN(n4419) );
  NAND2_X1 U5952 ( .A1(n8606), .A2(n4338), .ZN(P2_U3206) );
  NAND2_X1 U5953 ( .A1(n8772), .A2(n4344), .ZN(P2_U3486) );
  NAND2_X1 U5954 ( .A1(n8775), .A2(n4422), .ZN(P2_U3485) );
  INV_X1 U5955 ( .A(n4423), .ZN(n4422) );
  OAI21_X1 U5956 ( .B1(n8843), .B2(n8813), .A(n8774), .ZN(n4423) );
  NAND2_X1 U5957 ( .A1(n8836), .A2(n4345), .ZN(P2_U3454) );
  NAND2_X1 U5958 ( .A1(n8842), .A2(n4420), .ZN(P2_U3453) );
  INV_X1 U5959 ( .A(n4421), .ZN(n4420) );
  OAI21_X1 U5960 ( .B1(n8843), .B2(n8896), .A(n8841), .ZN(n4421) );
  NAND2_X1 U5961 ( .A1(n9873), .A2(n9348), .ZN(n4592) );
  AOI21_X1 U5962 ( .B1(n4639), .B2(n9630), .A(n4638), .ZN(n4637) );
  INV_X1 U5963 ( .A(n4832), .ZN(n4831) );
  NAND2_X1 U5964 ( .A1(n4574), .A2(n4572), .ZN(P1_U3551) );
  OR2_X1 U5965 ( .A1(n10124), .A2(n4573), .ZN(n4572) );
  NAND2_X1 U5966 ( .A1(n9934), .A2(n10124), .ZN(n4574) );
  INV_X1 U5967 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n4573) );
  NAND2_X1 U5968 ( .A1(n4508), .A2(n4384), .ZN(P1_U3519) );
  NAND2_X1 U5969 ( .A1(n9934), .A2(n4272), .ZN(n4508) );
  INV_X1 U5970 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n4507) );
  NAND2_X1 U5971 ( .A1(n8601), .A2(n4581), .ZN(n4291) );
  INV_X1 U5972 ( .A(n6429), .ZN(n4662) );
  OR2_X1 U5973 ( .A1(n7841), .A2(n6436), .ZN(n4292) );
  OR2_X1 U5974 ( .A1(n9711), .A2(n9286), .ZN(n4293) );
  AND2_X1 U5975 ( .A1(n5785), .A2(n4497), .ZN(n4294) );
  AND4_X1 U5976 ( .A1(n4314), .A2(n4980), .A3(n4701), .A4(n4700), .ZN(n5169)
         );
  AND2_X1 U5977 ( .A1(n7394), .A2(n7306), .ZN(n4295) );
  NAND2_X1 U5978 ( .A1(n7362), .A2(n4821), .ZN(n7759) );
  NAND2_X1 U5979 ( .A1(n6434), .A2(n5389), .ZN(n4296) );
  AND2_X1 U5980 ( .A1(n5719), .A2(n9801), .ZN(n9820) );
  INV_X1 U5981 ( .A(n9820), .ZN(n4697) );
  INV_X1 U5982 ( .A(n8401), .ZN(n7230) );
  AND2_X1 U5983 ( .A1(n4720), .A2(n5422), .ZN(n4297) );
  NOR2_X1 U5984 ( .A1(n9673), .A2(n9196), .ZN(n4298) );
  INV_X1 U5985 ( .A(n7827), .ZN(n9369) );
  INV_X1 U5986 ( .A(n9836), .ZN(n9838) );
  AND2_X1 U5987 ( .A1(n5791), .A2(n5793), .ZN(n9836) );
  AND2_X1 U5988 ( .A1(n4361), .A2(n4575), .ZN(n4299) );
  OR2_X1 U5989 ( .A1(n4987), .A2(n6268), .ZN(n4300) );
  AND2_X1 U5990 ( .A1(n4680), .A2(n4681), .ZN(n4301) );
  NAND2_X1 U5991 ( .A1(n7349), .A2(n7478), .ZN(n7425) );
  OR2_X1 U5992 ( .A1(n4629), .A2(n4631), .ZN(n4302) );
  AND2_X1 U5993 ( .A1(n6112), .A2(n4585), .ZN(n4303) );
  AND2_X1 U5994 ( .A1(n6171), .A2(n4590), .ZN(n4304) );
  AND2_X1 U5995 ( .A1(n7801), .A2(n4927), .ZN(n4305) );
  NAND2_X1 U5996 ( .A1(n7744), .A2(n4854), .ZN(n4855) );
  NAND2_X1 U5997 ( .A1(n6801), .A2(n9806), .ZN(n9348) );
  AND2_X1 U5998 ( .A1(n6271), .A2(n4580), .ZN(n4306) );
  INV_X1 U5999 ( .A(n8562), .ZN(n4523) );
  INV_X1 U6000 ( .A(n4882), .ZN(n6519) );
  AND2_X2 U6001 ( .A1(n8902), .A2(n8907), .ZN(n5995) );
  INV_X1 U6002 ( .A(n4735), .ZN(n9830) );
  OAI21_X1 U6003 ( .B1(n9960), .B2(n5678), .A(n5679), .ZN(n4735) );
  NAND2_X1 U6004 ( .A1(n5477), .A2(n5476), .ZN(n9903) );
  NAND2_X1 U6005 ( .A1(n6170), .A2(n6169), .ZN(n6552) );
  AND2_X1 U6006 ( .A1(n4467), .A2(n4465), .ZN(n4307) );
  NOR2_X1 U6007 ( .A1(n9914), .A2(n9364), .ZN(n4308) );
  NOR2_X1 U6008 ( .A1(n9157), .A2(n9370), .ZN(n4309) );
  AND2_X1 U6009 ( .A1(n7886), .A2(n7885), .ZN(n4310) );
  OR2_X1 U6010 ( .A1(n6552), .A2(n8740), .ZN(n4311) );
  NAND2_X1 U6011 ( .A1(n9092), .A2(n4975), .ZN(n4312) );
  OR2_X1 U6012 ( .A1(n8470), .A2(n8479), .ZN(n4313) );
  AND4_X2 U6013 ( .A1(n5858), .A2(n5142), .A3(n5857), .A4(n5244), .ZN(n4314)
         );
  AND2_X1 U6014 ( .A1(n9706), .A2(n4861), .ZN(n4315) );
  AOI21_X1 U6015 ( .B1(n9172), .B2(n4934), .A(n4312), .ZN(n4931) );
  INV_X1 U6016 ( .A(n4685), .ZN(n5305) );
  OR2_X1 U6017 ( .A1(n6447), .A2(n9232), .ZN(n4316) );
  INV_X1 U6018 ( .A(n6438), .ZN(n7503) );
  AND2_X1 U6019 ( .A1(n5721), .A2(n5827), .ZN(n6438) );
  NAND2_X1 U6020 ( .A1(n4320), .A2(n5296), .ZN(n10072) );
  AND2_X1 U6021 ( .A1(n8139), .A2(n8132), .ZN(n8658) );
  NAND2_X1 U6022 ( .A1(n5215), .A2(n5214), .ZN(n9914) );
  AND2_X1 U6023 ( .A1(n7417), .A2(n5722), .ZN(n7438) );
  OR2_X1 U6024 ( .A1(n4868), .A2(n6472), .ZN(n4317) );
  NAND2_X1 U6025 ( .A1(n5788), .A2(n5786), .ZN(n4318) );
  NOR2_X1 U6026 ( .A1(n7748), .A2(n6441), .ZN(n4319) );
  OR2_X1 U6027 ( .A1(n6671), .A2(n5678), .ZN(n4320) );
  OR2_X1 U6028 ( .A1(n8834), .A2(n6606), .ZN(n4321) );
  AND2_X1 U6029 ( .A1(n5708), .A2(n5725), .ZN(n4322) );
  AND2_X1 U6030 ( .A1(n6025), .A2(n4587), .ZN(n4323) );
  OR2_X1 U6031 ( .A1(n9928), .A2(n9367), .ZN(n4324) );
  OAI22_X1 U6032 ( .A1(n4546), .A2(n4544), .B1(n6456), .B2(n6455), .ZN(n9705)
         );
  AND2_X1 U6033 ( .A1(n4886), .A2(n4885), .ZN(n4325) );
  OAI21_X1 U6034 ( .B1(n6454), .B2(n4543), .A(n4542), .ZN(n9687) );
  NAND2_X1 U6035 ( .A1(n6454), .A2(n6453), .ZN(n9720) );
  NAND2_X1 U6036 ( .A1(n4553), .A2(n6461), .ZN(n9647) );
  NAND2_X1 U6037 ( .A1(n4964), .A2(n4967), .ZN(n9664) );
  OR2_X1 U6038 ( .A1(n8437), .A2(n8438), .ZN(n4326) );
  AND2_X1 U6039 ( .A1(n4989), .A2(n7938), .ZN(n4327) );
  AND2_X1 U6040 ( .A1(n6446), .A2(n6445), .ZN(n4328) );
  INV_X1 U6041 ( .A(n8197), .ZN(n4407) );
  OR2_X1 U6042 ( .A1(n8819), .A2(n8578), .ZN(n4329) );
  INV_X1 U6043 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n4936) );
  NAND2_X1 U6044 ( .A1(n5450), .A2(n5449), .ZN(n9922) );
  NAND2_X1 U6045 ( .A1(n6320), .A2(n6319), .ZN(n8828) );
  INV_X1 U6046 ( .A(n8828), .ZN(n4581) );
  AND2_X1 U6047 ( .A1(n6093), .A2(n7359), .ZN(n4330) );
  AND2_X1 U6048 ( .A1(n8828), .A2(n8168), .ZN(n4331) );
  OR2_X1 U6049 ( .A1(n5640), .A2(n5641), .ZN(n4332) );
  AND4_X1 U6050 ( .A1(n5858), .A2(n5857), .A3(n4557), .A4(n5244), .ZN(n4333)
         );
  AND2_X1 U6051 ( .A1(n8309), .A2(n8740), .ZN(n4334) );
  OR2_X1 U6052 ( .A1(n4626), .A2(n4629), .ZN(n4335) );
  NOR2_X1 U6053 ( .A1(n6574), .A2(n6606), .ZN(n4336) );
  OR2_X1 U6054 ( .A1(n8787), .A2(n6565), .ZN(n8139) );
  INV_X1 U6055 ( .A(n8139), .ZN(n4894) );
  NOR2_X1 U6056 ( .A1(n8376), .A2(n4816), .ZN(n4337) );
  AND2_X1 U6057 ( .A1(n4413), .A2(n8605), .ZN(n4338) );
  AND2_X1 U6058 ( .A1(n5304), .A2(n5303), .ZN(n4339) );
  AOI21_X1 U6059 ( .B1(n8483), .B2(n4628), .A(n4625), .ZN(n4622) );
  INV_X1 U6060 ( .A(n6456), .ZN(n4549) );
  OR2_X1 U6061 ( .A1(n4690), .A2(n5279), .ZN(n4340) );
  AND2_X1 U6062 ( .A1(n9711), .A2(n9286), .ZN(n4341) );
  OR2_X1 U6063 ( .A1(n6814), .A2(n7213), .ZN(n4342) );
  INV_X1 U6064 ( .A(n4968), .ZN(n4967) );
  INV_X1 U6065 ( .A(n4785), .ZN(n4783) );
  OAI21_X1 U6066 ( .B1(n4978), .B2(n8558), .A(n4788), .ZN(n4785) );
  NOR2_X1 U6067 ( .A1(n9636), .A2(n9612), .ZN(n4343) );
  INV_X1 U6068 ( .A(n9859), .ZN(n9673) );
  NAND2_X1 U6069 ( .A1(n5605), .A2(n5604), .ZN(n9859) );
  AND2_X1 U6070 ( .A1(n4412), .A2(n8771), .ZN(n4344) );
  AND2_X1 U6071 ( .A1(n4414), .A2(n8835), .ZN(n4345) );
  NAND2_X1 U6072 ( .A1(n8803), .A2(n8725), .ZN(n4346) );
  NOR2_X1 U6073 ( .A1(n8094), .A2(n8095), .ZN(n4347) );
  INV_X1 U6074 ( .A(n9665), .ZN(n4872) );
  AND2_X1 U6075 ( .A1(n7960), .A2(n4916), .ZN(n4348) );
  INV_X1 U6076 ( .A(n6567), .ZN(n4750) );
  OR2_X1 U6077 ( .A1(n8787), .A2(n8671), .ZN(n6567) );
  NOR2_X1 U6078 ( .A1(n8834), .A2(n8611), .ZN(n4349) );
  NOR2_X1 U6079 ( .A1(n9775), .A2(n6450), .ZN(n4350) );
  NOR2_X1 U6080 ( .A1(n9083), .A2(n6439), .ZN(n4351) );
  INV_X1 U6081 ( .A(n9215), .ZN(n4926) );
  INV_X1 U6082 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n9110) );
  INV_X1 U6083 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5150) );
  OR2_X1 U6084 ( .A1(n5760), .A2(n5761), .ZN(n4352) );
  INV_X1 U6085 ( .A(n7394), .ZN(n7406) );
  AND2_X1 U6086 ( .A1(n6081), .A2(n6056), .ZN(n7394) );
  INV_X1 U6087 ( .A(n4977), .ZN(n4751) );
  AND2_X1 U6088 ( .A1(n5042), .A2(SI_7_), .ZN(n4353) );
  NAND2_X1 U6089 ( .A1(n7846), .A2(n9180), .ZN(n4354) );
  AND2_X1 U6090 ( .A1(n5062), .A2(SI_12_), .ZN(n4355) );
  NAND2_X1 U6091 ( .A1(n8244), .A2(n9625), .ZN(n4356) );
  OR2_X1 U6092 ( .A1(n6401), .A2(n4987), .ZN(n4357) );
  NAND2_X1 U6093 ( .A1(n4291), .A2(n4321), .ZN(n4358) );
  NAND2_X1 U6094 ( .A1(n5627), .A2(n5628), .ZN(n4359) );
  INV_X1 U6095 ( .A(n9763), .ZN(n4479) );
  AND2_X1 U6096 ( .A1(n5288), .A2(n5287), .ZN(n4360) );
  NAND2_X1 U6097 ( .A1(n9726), .A2(n4990), .ZN(n9689) );
  AND2_X1 U6098 ( .A1(n8541), .A2(n8542), .ZN(n4527) );
  AND2_X1 U6099 ( .A1(n9847), .A2(n4863), .ZN(n4361) );
  AND2_X1 U6100 ( .A1(n8840), .A2(n8602), .ZN(n6572) );
  AND2_X1 U6101 ( .A1(n4805), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4362) );
  OR2_X1 U6102 ( .A1(n4343), .A2(n4969), .ZN(n4363) );
  OR2_X1 U6103 ( .A1(n4682), .A2(n4332), .ZN(n4680) );
  INV_X1 U6104 ( .A(n9747), .ZN(n9882) );
  AND2_X1 U6105 ( .A1(n5540), .A2(n5539), .ZN(n9747) );
  AND2_X1 U6106 ( .A1(n7448), .A2(n8066), .ZN(n8183) );
  INV_X1 U6107 ( .A(n8183), .ZN(n4901) );
  NAND2_X1 U6108 ( .A1(n4548), .A2(n4547), .ZN(n4364) );
  NAND2_X1 U6109 ( .A1(n5615), .A2(n5614), .ZN(n9863) );
  AND2_X1 U6110 ( .A1(n4875), .A2(n6471), .ZN(n4365) );
  OR2_X1 U6111 ( .A1(n8828), .A2(n8601), .ZN(n4366) );
  AND3_X1 U6112 ( .A1(n8099), .A2(n4796), .A3(n8192), .ZN(n4367) );
  AND3_X1 U6113 ( .A1(n5857), .A2(n5141), .A3(n4999), .ZN(n4368) );
  AND2_X1 U6114 ( .A1(n4417), .A2(n8595), .ZN(n4369) );
  NAND2_X1 U6115 ( .A1(n6261), .A2(n8631), .ZN(n4370) );
  AND4_X1 U6116 ( .A1(n5352), .A2(n5351), .A3(n5350), .A4(n5349), .ZN(n7827)
         );
  AND2_X1 U6117 ( .A1(n6178), .A2(n8357), .ZN(n4371) );
  NAND2_X1 U6118 ( .A1(n4930), .A2(n7800), .ZN(n4929) );
  INV_X1 U6119 ( .A(n4929), .ZN(n4928) );
  INV_X1 U6120 ( .A(n8188), .ZN(n8092) );
  AND2_X1 U6121 ( .A1(n4858), .A2(n9281), .ZN(n4372) );
  AND2_X1 U6122 ( .A1(n8853), .A2(n8621), .ZN(n8170) );
  AND2_X1 U6123 ( .A1(n5787), .A2(n5786), .ZN(n4373) );
  AND3_X1 U6124 ( .A1(n4479), .A2(n5788), .A3(n4478), .ZN(n4374) );
  AND2_X1 U6125 ( .A1(n4697), .A2(n5789), .ZN(n4375) );
  AND2_X1 U6126 ( .A1(n6011), .A2(n6012), .ZN(n4376) );
  AND2_X1 U6127 ( .A1(n4418), .A2(n8829), .ZN(n4377) );
  AND2_X1 U6128 ( .A1(n4648), .A2(n5148), .ZN(n4378) );
  OR2_X1 U6129 ( .A1(n6812), .A2(n6813), .ZN(n4379) );
  NAND2_X1 U6130 ( .A1(n5150), .A2(n5147), .ZN(n4380) );
  INV_X1 U6131 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n4805) );
  OR2_X1 U6132 ( .A1(n4581), .A2(n8168), .ZN(n4381) );
  INV_X2 U6133 ( .A(n9996), .ZN(n9768) );
  NAND2_X2 U6134 ( .A1(n6908), .A2(n8655), .ZN(n10186) );
  NOR2_X1 U6135 ( .A1(n9908), .A2(n9914), .ZN(n4854) );
  NAND2_X1 U6136 ( .A1(n4838), .A2(n7406), .ZN(n7399) );
  AND2_X1 U6137 ( .A1(n8416), .A2(n8453), .ZN(n4382) );
  OAI211_X1 U6138 ( .C1(n4271), .C2(n8892), .A(n6165), .B(n6164), .ZN(n8724)
         );
  NAND2_X1 U6139 ( .A1(n5771), .A2(n4693), .ZN(n7206) );
  XNOR2_X1 U6140 ( .A(n6144), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8479) );
  INV_X1 U6141 ( .A(n8479), .ZN(n4856) );
  AND3_X1 U6142 ( .A1(n9799), .A2(n7744), .A3(n4852), .ZN(n9770) );
  INV_X1 U6143 ( .A(n8438), .ZN(n8419) );
  AND2_X1 U6144 ( .A1(n5650), .A2(n5649), .ZN(n4383) );
  OAI21_X1 U6145 ( .B1(n7504), .B2(n6438), .A(n6437), .ZN(n7570) );
  OR2_X1 U6146 ( .A1(n4272), .A2(n4507), .ZN(n4384) );
  NAND2_X1 U6147 ( .A1(n4537), .A2(n6432), .ZN(n7248) );
  NAND2_X1 U6148 ( .A1(n4538), .A2(n6430), .ZN(n9997) );
  AND2_X1 U6149 ( .A1(n5771), .A2(n5770), .ZN(n4385) );
  AOI21_X1 U6150 ( .B1(n7055), .B2(n7054), .A(n7053), .ZN(n7059) );
  INV_X1 U6151 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n6124) );
  AND2_X1 U6152 ( .A1(n5549), .A2(n5548), .ZN(n9285) );
  INV_X1 U6153 ( .A(n9285), .ZN(n9358) );
  AND2_X1 U6154 ( .A1(n4923), .A2(n7804), .ZN(n4386) );
  OR2_X1 U6155 ( .A1(n9535), .A2(n9534), .ZN(n4387) );
  INV_X1 U6156 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n9081) );
  INV_X1 U6157 ( .A(n8620), .ZN(n8602) );
  AND2_X1 U6158 ( .A1(n6305), .A2(n6304), .ZN(n8620) );
  AND2_X1 U6159 ( .A1(n4595), .A2(n4599), .ZN(n4388) );
  NAND2_X1 U6160 ( .A1(n6048), .A2(n7359), .ZN(n7362) );
  AND2_X1 U6161 ( .A1(n7362), .A2(n6050), .ZN(n4389) );
  AND2_X1 U6162 ( .A1(n4867), .A2(n5776), .ZN(n4390) );
  NOR2_X1 U6163 ( .A1(n6900), .A2(n8229), .ZN(n4391) );
  INV_X1 U6164 ( .A(n10229), .ZN(n10227) );
  NAND2_X1 U6165 ( .A1(n6362), .A2(n6361), .ZN(n8367) );
  INV_X1 U6166 ( .A(n5388), .ZN(n4948) );
  NAND2_X1 U6167 ( .A1(n8174), .A2(n6581), .ZN(n6891) );
  NAND2_X1 U6168 ( .A1(n6480), .A2(n6479), .ZN(n10030) );
  OR2_X1 U6169 ( .A1(n7138), .A2(n6425), .ZN(n4392) );
  INV_X1 U6170 ( .A(n6516), .ZN(n4432) );
  NAND2_X1 U6171 ( .A1(n6521), .A2(n6520), .ZN(n7015) );
  NAND2_X1 U6172 ( .A1(n5279), .A2(n5278), .ZN(n10027) );
  AND2_X1 U6173 ( .A1(n9578), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n4393) );
  NOR2_X1 U6174 ( .A1(n8554), .A2(n8728), .ZN(n4394) );
  NOR2_X2 U6175 ( .A1(n6821), .A2(n9390), .ZN(n4395) );
  NAND4_X1 U6176 ( .A1(n4284), .A2(n5917), .A3(n4902), .A4(n5913), .ZN(n4396)
         );
  AND2_X1 U6177 ( .A1(n5580), .A2(n5579), .ZN(n9711) );
  INV_X1 U6178 ( .A(n9711), .ZN(n9873) );
  INV_X1 U6179 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n9096) );
  INV_X1 U6180 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n4580) );
  INV_X1 U6181 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n4585) );
  OR2_X1 U6182 ( .A1(n9592), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n4397) );
  NAND2_X1 U6183 ( .A1(n6008), .A2(n6007), .ZN(n10215) );
  INV_X1 U6184 ( .A(n10215), .ZN(n4806) );
  INV_X1 U6185 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n4532) );
  INV_X1 U6186 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n5971) );
  INV_X1 U6187 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n4438) );
  INV_X1 U6188 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n4851) );
  NAND2_X1 U6189 ( .A1(n5442), .A2(n4403), .ZN(n4402) );
  NAND2_X1 U6190 ( .A1(n8144), .A2(n4406), .ZN(n8145) );
  NAND3_X1 U6191 ( .A1(n4455), .A2(n4408), .A3(n4456), .ZN(n8032) );
  NAND3_X1 U6192 ( .A1(n5886), .A2(n4411), .A3(n5885), .ZN(P1_U3242) );
  NAND2_X1 U6193 ( .A1(n5884), .A2(n5883), .ZN(n4411) );
  INV_X1 U6194 ( .A(n5393), .ZN(n4665) );
  INV_X1 U6195 ( .A(n5639), .ZN(n4676) );
  INV_X1 U6196 ( .A(n5466), .ZN(n4655) );
  NAND2_X1 U6197 ( .A1(n4650), .A2(n9802), .ZN(n5552) );
  NOR2_X1 U6198 ( .A1(n4657), .A2(n4658), .ZN(n4656) );
  NAND2_X1 U6199 ( .A1(n4797), .A2(n4367), .ZN(n8105) );
  AOI21_X1 U6200 ( .B1(n8162), .B2(n8208), .A(n8209), .ZN(n8222) );
  OAI21_X1 U6201 ( .B1(n8114), .B2(n8110), .A(n8109), .ZN(n4453) );
  OAI211_X1 U6202 ( .C1(n8154), .C2(n4769), .A(n8160), .B(n4767), .ZN(n4772)
         );
  AOI21_X2 U6203 ( .B1(n4756), .B2(n4752), .A(n4753), .ZN(n8698) );
  AOI21_X2 U6204 ( .B1(n8618), .B2(n8148), .A(n6571), .ZN(n8610) );
  NAND2_X1 U6205 ( .A1(n6522), .A2(n10176), .ZN(n8045) );
  NAND2_X1 U6206 ( .A1(n6306), .A2(n8365), .ZN(n6506) );
  AOI211_X1 U6207 ( .C1(n8214), .C2(n8213), .A(n8212), .B(n8211), .ZN(n8224)
         );
  OAI22_X2 U6208 ( .A1(n7257), .A2(n4761), .B1(n7230), .B2(n4806), .ZN(n7379)
         );
  AOI21_X2 U6209 ( .B1(n8629), .B2(n6570), .A(n6569), .ZN(n8618) );
  NAND2_X1 U6210 ( .A1(n6548), .A2(n6547), .ZN(n7598) );
  OAI21_X1 U6211 ( .B1(n6651), .B2(n10227), .A(n6653), .ZN(n6654) );
  NAND2_X1 U6212 ( .A1(n8830), .A2(n4377), .ZN(P2_U3455) );
  NAND2_X1 U6213 ( .A1(n8596), .A2(n4369), .ZN(P2_U3205) );
  NAND3_X1 U6214 ( .A1(n8770), .A2(n8769), .A3(n4416), .ZN(P2_U3487) );
  NAND2_X1 U6215 ( .A1(n8768), .A2(n8767), .ZN(n8770) );
  NOR2_X1 U6216 ( .A1(n7871), .A2(n7870), .ZN(n9076) );
  OAI21_X1 U6217 ( .B1(n9117), .B2(n7919), .A(n7918), .ZN(n7921) );
  NAND2_X1 U6218 ( .A1(n8827), .A2(n10229), .ZN(n8768) );
  XNOR2_X1 U6219 ( .A(n8610), .B(n8609), .ZN(n4427) );
  NAND2_X1 U6220 ( .A1(n6535), .A2(n6534), .ZN(n7591) );
  NAND2_X1 U6221 ( .A1(n6605), .A2(n8128), .ZN(n8659) );
  OAI21_X2 U6222 ( .B1(n8598), .B2(n4358), .A(n4879), .ZN(n8015) );
  NAND2_X1 U6223 ( .A1(n7255), .A2(n8040), .ZN(n6585) );
  INV_X1 U6224 ( .A(n7286), .ZN(n4428) );
  NAND2_X1 U6225 ( .A1(n4905), .A2(n4904), .ZN(n8678) );
  NAND2_X2 U6226 ( .A1(n4828), .A2(n8267), .ZN(n8330) );
  NAND2_X1 U6227 ( .A1(n7157), .A2(n5990), .ZN(n7146) );
  INV_X1 U6228 ( .A(n8354), .ZN(n4431) );
  INV_X1 U6229 ( .A(n7788), .ZN(n6139) );
  NAND2_X1 U6230 ( .A1(n6861), .A2(n5950), .ZN(n7095) );
  NAND2_X1 U6231 ( .A1(n5989), .A2(n5988), .ZN(n7157) );
  AOI21_X1 U6232 ( .B1(n4811), .B2(n6166), .A(n4371), .ZN(n4809) );
  OAI21_X1 U6233 ( .B1(n8483), .B2(n4625), .A(n4623), .ZN(n4633) );
  AOI21_X1 U6234 ( .B1(n8533), .B2(n8532), .A(n8531), .ZN(n8536) );
  AOI22_X1 U6235 ( .A1(n7396), .A2(n7395), .B1(n7394), .B2(n7393), .ZN(n7531)
         );
  NOR2_X1 U6236 ( .A1(n6755), .A2(n6756), .ZN(n6870) );
  NOR2_X1 U6237 ( .A1(n6870), .A2(n4439), .ZN(n6874) );
  NOR2_X1 U6238 ( .A1(n8563), .A2(n8537), .ZN(n8538) );
  OAI22_X1 U6239 ( .A1(n7304), .A2(n7303), .B1(n7302), .B2(n7301), .ZN(n7396)
         );
  OAI21_X1 U6240 ( .B1(n6955), .B2(n4270), .A(n10139), .ZN(n10146) );
  OR2_X2 U6241 ( .A1(n9076), .A2(n9079), .ZN(n4594) );
  AOI21_X1 U6242 ( .B1(n4599), .B2(n4601), .A(n4597), .ZN(n4596) );
  NAND2_X1 U6243 ( .A1(n6754), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n6880) );
  NOR2_X2 U6244 ( .A1(n4463), .A2(n8545), .ZN(n8518) );
  NAND2_X2 U6245 ( .A1(n8518), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n8547) );
  NAND2_X1 U6246 ( .A1(n6966), .A2(n7073), .ZN(n7080) );
  NAND2_X1 U6247 ( .A1(n7180), .A2(n7179), .ZN(n7181) );
  OAI21_X1 U6248 ( .B1(n8490), .B2(n4514), .A(n4512), .ZN(n8513) );
  AND2_X1 U6249 ( .A1(n5733), .A2(n4374), .ZN(n5736) );
  XNOR2_X1 U6250 ( .A(n8600), .B(n8599), .ZN(n4474) );
  AOI21_X1 U6251 ( .B1(n4474), .B2(n10178), .A(n4472), .ZN(n8832) );
  NAND3_X1 U6252 ( .A1(n4576), .A2(n6624), .A3(n4577), .ZN(n6651) );
  AOI21_X1 U6253 ( .B1(n8592), .B2(n10178), .A(n8591), .ZN(n8827) );
  NAND2_X1 U6254 ( .A1(n7014), .A2(n8175), .ZN(n6583) );
  NAND2_X1 U6255 ( .A1(n4476), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n5593) );
  INV_X1 U6256 ( .A(n5164), .ZN(n5607) );
  NAND2_X1 U6257 ( .A1(n4677), .A2(n4684), .ZN(n4674) );
  NAND2_X1 U6258 ( .A1(n9442), .A2(n4379), .ZN(n9459) );
  OAI21_X1 U6259 ( .B1(n9599), .B2(n9986), .A(n4640), .ZN(n4639) );
  NOR2_X1 U6260 ( .A1(n7103), .A2(n4635), .ZN(n9492) );
  NAND2_X1 U6261 ( .A1(n9492), .A2(n9491), .ZN(n9490) );
  NOR2_X1 U6262 ( .A1(n9517), .A2(n4636), .ZN(n9520) );
  NAND2_X1 U6263 ( .A1(n9520), .A2(n9519), .ZN(n9533) );
  NOR2_X1 U6264 ( .A1(n9571), .A2(n4393), .ZN(n9572) );
  OAI21_X1 U6265 ( .B1(n9601), .B2(n9630), .A(n4637), .ZN(P1_U3262) );
  AOI21_X2 U6266 ( .B1(n6048), .B2(n4330), .A(n4817), .ZN(n7560) );
  NAND2_X1 U6267 ( .A1(n9273), .A2(n9274), .ZN(n9272) );
  NAND2_X1 U6268 ( .A1(n7921), .A2(n9169), .ZN(n9172) );
  NOR2_X1 U6269 ( .A1(n4307), .A2(n6792), .ZN(n6847) );
  INV_X1 U6270 ( .A(n4927), .ZN(n4922) );
  NAND2_X1 U6271 ( .A1(n9312), .A2(n7823), .ZN(n4911) );
  NAND2_X1 U6272 ( .A1(n5000), .A2(n4368), .ZN(n5197) );
  NAND2_X1 U6273 ( .A1(n5005), .A2(n4971), .ZN(n5008) );
  NOR2_X1 U6274 ( .A1(n9313), .A2(n9314), .ZN(n9312) );
  OAI21_X1 U6275 ( .B1(n7851), .B2(n7850), .A(n9181), .ZN(n7852) );
  NAND3_X1 U6276 ( .A1(n8121), .A2(n4454), .A3(n4453), .ZN(n4762) );
  NAND2_X1 U6277 ( .A1(n4794), .A2(n4795), .ZN(n4793) );
  NOR2_X1 U6278 ( .A1(n4772), .A2(n8161), .ZN(n8209) );
  NAND2_X1 U6279 ( .A1(n4457), .A2(n6850), .ZN(n6851) );
  NAND2_X1 U6280 ( .A1(n7036), .A2(n10043), .ZN(n4457) );
  OR2_X4 U6282 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n6764) );
  NAND2_X1 U6283 ( .A1(n10157), .A2(n6965), .ZN(n6966) );
  AOI21_X1 U6284 ( .B1(n8576), .B2(n10129), .A(n4616), .ZN(n4615) );
  AND2_X1 U6285 ( .A1(n4470), .A2(n5950), .ZN(n6863) );
  NOR2_X1 U6286 ( .A1(n7269), .A2(n4618), .ZN(n7304) );
  NOR2_X1 U6287 ( .A1(n6874), .A2(n6873), .ZN(n6953) );
  NAND2_X2 U6289 ( .A1(n7699), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n7698) );
  INV_X1 U6290 ( .A(n8416), .ZN(n4847) );
  INV_X1 U6291 ( .A(n8415), .ZN(n4462) );
  NOR2_X2 U6292 ( .A1(n8517), .A2(n8533), .ZN(n8545) );
  NAND2_X2 U6293 ( .A1(n7272), .A2(n7273), .ZN(n7307) );
  AOI21_X1 U6294 ( .B1(n6848), .B2(n6923), .A(n6847), .ZN(n6930) );
  NOR2_X2 U6295 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n5251) );
  AND2_X2 U6296 ( .A1(n5913), .A2(n5917), .ZN(n4608) );
  AND3_X2 U6297 ( .A1(n5894), .A2(n5895), .A3(n5893), .ZN(n5917) );
  AND3_X2 U6298 ( .A1(n5892), .A2(n5891), .A3(n5890), .ZN(n5913) );
  AND2_X1 U6299 ( .A1(n8045), .A2(n8033), .ZN(n8175) );
  OAI21_X2 U6300 ( .B1(n8607), .B2(n8608), .A(n8155), .ZN(n8598) );
  NAND2_X1 U6301 ( .A1(n8732), .A2(n8101), .ZN(n4905) );
  NAND2_X1 U6302 ( .A1(n4898), .A2(n4896), .ZN(n7490) );
  OR2_X1 U6303 ( .A1(n4267), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n5910) );
  NAND2_X1 U6304 ( .A1(n6179), .A2(n5915), .ZN(n6181) );
  NOR2_X2 U6305 ( .A1(n5197), .A2(n5002), .ZN(n5741) );
  AND2_X2 U6306 ( .A1(n5905), .A2(n5899), .ZN(n5929) );
  NAND2_X1 U6307 ( .A1(n4598), .A2(n4596), .ZN(n9273) );
  NOR2_X2 U6308 ( .A1(n6506), .A2(n6505), .ZN(n6514) );
  NAND2_X1 U6309 ( .A1(n7059), .A2(n4920), .ZN(n4602) );
  INV_X1 U6310 ( .A(n4680), .ZN(n4677) );
  NAND2_X1 U6311 ( .A1(n5162), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n5616) );
  OAI21_X1 U6312 ( .B1(n4681), .B2(n4675), .A(n4674), .ZN(n4673) );
  NAND2_X1 U6313 ( .A1(n4878), .A2(n5040), .ZN(n5369) );
  NAND4_X1 U6314 ( .A1(n5881), .A2(n9648), .A3(n6478), .A4(n5739), .ZN(n5740)
         );
  INV_X1 U6315 ( .A(n5037), .ZN(n4482) );
  INV_X1 U6316 ( .A(n5294), .ZN(n4483) );
  NAND2_X1 U6317 ( .A1(n4865), .A2(n5032), .ZN(n4484) );
  NAND2_X1 U6318 ( .A1(n5029), .A2(n5028), .ZN(n5242) );
  NAND2_X1 U6319 ( .A1(n4294), .A2(n4375), .ZN(n4486) );
  INV_X1 U6320 ( .A(n5789), .ZN(n4489) );
  NAND2_X1 U6321 ( .A1(n9785), .A2(n5789), .ZN(n9777) );
  NAND2_X1 U6322 ( .A1(n4490), .A2(n4695), .ZN(n9785) );
  NAND2_X1 U6323 ( .A1(n5354), .A2(n5047), .ZN(n4502) );
  NOR2_X1 U6324 ( .A1(n4501), .A2(n4500), .ZN(n4499) );
  INV_X1 U6325 ( .A(n5047), .ZN(n4500) );
  NAND2_X1 U6326 ( .A1(n10150), .A2(n10149), .ZN(n10148) );
  NAND2_X1 U6327 ( .A1(n10131), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n4509) );
  NAND2_X1 U6328 ( .A1(n7405), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n7409) );
  NAND2_X1 U6329 ( .A1(n7299), .A2(n7298), .ZN(n4510) );
  NAND2_X1 U6330 ( .A1(n7697), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n7527) );
  NAND2_X1 U6331 ( .A1(n7410), .A2(n7411), .ZN(n7524) );
  NAND3_X1 U6332 ( .A1(n4528), .A2(n4617), .A3(n4615), .ZN(P2_U3201) );
  NAND2_X1 U6333 ( .A1(n9997), .A2(n9998), .ZN(n4537) );
  NAND2_X1 U6334 ( .A1(n7205), .A2(n7207), .ZN(n4538) );
  INV_X1 U6335 ( .A(n4539), .ZN(n6459) );
  NAND2_X1 U6336 ( .A1(n4964), .A2(n4554), .ZN(n4552) );
  AND2_X1 U6337 ( .A1(n5142), .A2(n4936), .ZN(n4557) );
  NAND2_X1 U6338 ( .A1(n4333), .A2(n4980), .ZN(n4558) );
  NAND2_X1 U6339 ( .A1(n7504), .A2(n4957), .ZN(n4563) );
  INV_X1 U6340 ( .A(n7418), .ZN(n4567) );
  NAND2_X1 U6341 ( .A1(n4563), .A2(n4568), .ZN(n9811) );
  INV_X1 U6342 ( .A(n4566), .ZN(n4564) );
  INV_X1 U6343 ( .A(n4308), .ZN(n4569) );
  INV_X1 U6344 ( .A(n6621), .ZN(n4576) );
  NAND4_X1 U6345 ( .A1(n4577), .A2(n4576), .A3(n6624), .A4(n10217), .ZN(n6634)
         );
  NAND2_X1 U6346 ( .A1(n6272), .A2(n4306), .ZN(n6310) );
  NAND2_X1 U6347 ( .A1(n6272), .A2(n6271), .ZN(n6299) );
  NAND2_X1 U6348 ( .A1(n6113), .A2(n4583), .ZN(n6162) );
  NAND2_X1 U6349 ( .A1(n6026), .A2(n4586), .ZN(n6074) );
  NAND3_X1 U6350 ( .A1(n5970), .A2(n5971), .A3(n5996), .ZN(n6009) );
  NAND4_X1 U6351 ( .A1(n5970), .A2(n5971), .A3(n5996), .A4(n4591), .ZN(n6027)
         );
  NAND3_X1 U6352 ( .A1(n9100), .A2(n9099), .A3(n4592), .ZN(P1_U3216) );
  NAND3_X1 U6353 ( .A1(n7888), .A2(n4593), .A3(n7887), .ZN(n9228) );
  NAND2_X1 U6354 ( .A1(n9203), .A2(n7881), .ZN(n4593) );
  NAND2_X1 U6355 ( .A1(n9101), .A2(n4599), .ZN(n4598) );
  NAND3_X1 U6356 ( .A1(n4602), .A2(n4919), .A3(n4924), .ZN(n9313) );
  AND2_X2 U6357 ( .A1(n5856), .A2(n5146), .ZN(n4980) );
  AND2_X2 U6358 ( .A1(n5251), .A2(n8945), .ZN(n5244) );
  NAND2_X2 U6359 ( .A1(n4604), .A2(n4603), .ZN(n6790) );
  NAND4_X1 U6360 ( .A1(n6124), .A2(n4607), .A3(n4606), .A4(n4605), .ZN(n4807)
         );
  AND4_X4 U6361 ( .A1(n4608), .A2(n4759), .A3(n4760), .A4(n4902), .ZN(n5905)
         );
  NAND2_X1 U6362 ( .A1(n10146), .A2(n4614), .ZN(n4609) );
  NAND2_X1 U6363 ( .A1(n4609), .A2(n4611), .ZN(n7067) );
  OAI211_X1 U6364 ( .C1(n6958), .C2(n4613), .A(n10166), .B(n7067), .ZN(n6974)
         );
  INV_X1 U6365 ( .A(n4633), .ZN(n8531) );
  INV_X2 U6366 ( .A(n8564), .ZN(n8534) );
  MUX2_X1 U6367 ( .A(P2_REG1_REG_2__SCAN_IN), .B(P2_REG2_REG_2__SCAN_IN), .S(
        n8564), .Z(n6954) );
  NAND2_X1 U6368 ( .A1(n10060), .A2(n5284), .ZN(n5812) );
  NAND2_X1 U6369 ( .A1(n4647), .A2(n4378), .ZN(n5149) );
  NAND4_X1 U6370 ( .A1(n4314), .A2(n4980), .A3(P1_IR_REG_28__SCAN_IN), .A4(
        n4649), .ZN(n4647) );
  OAI21_X1 U6371 ( .B1(n4339), .B2(n4659), .A(n4656), .ZN(n5440) );
  NAND2_X1 U6372 ( .A1(n4688), .A2(n4340), .ZN(n5768) );
  INV_X1 U6373 ( .A(n5755), .ZN(n4684) );
  XNOR2_X2 U6374 ( .A(n5171), .B(n5170), .ZN(n8255) );
  NAND3_X1 U6375 ( .A1(n5172), .A2(P1_REG1_REG_1__SCAN_IN), .A3(n8255), .ZN(
        n4687) );
  NAND2_X2 U6376 ( .A1(n4273), .A2(n9964), .ZN(n5310) );
  INV_X1 U6377 ( .A(n5812), .ZN(n4690) );
  NAND3_X1 U6378 ( .A1(n5776), .A2(n4867), .A3(n7344), .ZN(n7343) );
  NAND3_X1 U6379 ( .A1(n4692), .A2(n6434), .A3(n6429), .ZN(n4691) );
  NAND2_X1 U6380 ( .A1(n7738), .A2(n4294), .ZN(n4695) );
  NAND2_X1 U6381 ( .A1(n7571), .A2(n5779), .ZN(n7575) );
  NAND3_X1 U6382 ( .A1(n4314), .A2(n4980), .A3(n4701), .ZN(n5165) );
  AND2_X1 U6383 ( .A1(n9859), .A2(n10084), .ZN(n4703) );
  NAND2_X1 U6384 ( .A1(n5179), .A2(n5180), .ZN(n4711) );
  NAND2_X1 U6385 ( .A1(n5179), .A2(n4712), .ZN(n4710) );
  OAI21_X1 U6386 ( .B1(n5053), .B2(n4720), .A(n4717), .ZN(n5423) );
  NAND2_X1 U6387 ( .A1(n5053), .A2(n5052), .ZN(n5407) );
  NAND2_X1 U6388 ( .A1(n5098), .A2(n5097), .ZN(n5533) );
  NAND2_X1 U6389 ( .A1(n5221), .A2(n5070), .ZN(n4733) );
  NAND2_X1 U6390 ( .A1(n4733), .A2(n5071), .ZN(n5190) );
  INV_X1 U6391 ( .A(n5073), .ZN(n4734) );
  NAND2_X1 U6392 ( .A1(n5133), .A2(n5132), .ZN(n5179) );
  AOI21_X1 U6393 ( .B1(n5571), .B2(n5570), .A(n5569), .ZN(n5639) );
  NOR2_X1 U6394 ( .A1(n5666), .A2(n5665), .ZN(n5713) );
  NAND2_X1 U6395 ( .A1(n5121), .A2(n5120), .ZN(n5612) );
  OAI21_X1 U6396 ( .B1(n5502), .B2(n5096), .A(n5095), .ZN(n5098) );
  NAND2_X1 U6397 ( .A1(n5674), .A2(n5673), .ZN(n5677) );
  XNOR2_X1 U6398 ( .A(n8015), .B(n8162), .ZN(n6623) );
  AND2_X2 U6399 ( .A1(n9621), .A2(n6476), .ZN(n5642) );
  NAND2_X1 U6400 ( .A1(n8610), .A2(n4738), .ZN(n4737) );
  NAND3_X1 U6401 ( .A1(n4737), .A2(n4381), .A3(n4736), .ZN(n6578) );
  NAND2_X1 U6402 ( .A1(n4744), .A2(n4743), .ZN(n6525) );
  NAND3_X1 U6403 ( .A1(n8045), .A2(n6524), .A3(n8033), .ZN(n4745) );
  INV_X2 U6404 ( .A(n4757), .ZN(n8564) );
  NAND2_X4 U6405 ( .A1(n6367), .A2(n4757), .ZN(n6614) );
  MUX2_X1 U6406 ( .A(P2_REG1_REG_0__SCAN_IN), .B(P2_REG2_REG_0__SCAN_IN), .S(
        n8564), .Z(n6727) );
  OR2_X1 U6407 ( .A1(n5909), .A2(n5908), .ZN(n4758) );
  NOR2_X1 U6408 ( .A1(n4807), .A2(P2_IR_REG_23__SCAN_IN), .ZN(n4760) );
  OAI21_X1 U6409 ( .B1(n7379), .B2(n6533), .A(n6532), .ZN(n6535) );
  NAND2_X1 U6410 ( .A1(n8141), .A2(n8142), .ZN(n8144) );
  NAND3_X1 U6411 ( .A1(n4763), .A2(n4762), .A3(n4765), .ZN(n8142) );
  NAND4_X1 U6412 ( .A1(n4777), .A2(n8230), .A3(n4776), .A4(n4775), .ZN(
        P2_U3296) );
  NAND4_X1 U6413 ( .A1(n8224), .A2(n4784), .A3(n8558), .A4(n4783), .ZN(n4775)
         );
  OR2_X1 U6414 ( .A1(n8224), .A2(n4781), .ZN(n4776) );
  INV_X1 U6415 ( .A(n4784), .ZN(n4778) );
  AOI21_X2 U6416 ( .B1(n4780), .B2(n4789), .A(n4779), .ZN(n4784) );
  INV_X1 U6417 ( .A(n8223), .ZN(n4779) );
  NAND4_X1 U6418 ( .A1(n4793), .A2(n4790), .A3(n8191), .A4(n4798), .ZN(n4797)
         );
  NAND2_X1 U6419 ( .A1(n4792), .A2(n4791), .ZN(n4790) );
  INV_X1 U6420 ( .A(n8086), .ZN(n4792) );
  INV_X1 U6421 ( .A(n8085), .ZN(n4794) );
  AOI21_X1 U6422 ( .B1(n4799), .B2(n8188), .A(n8096), .ZN(n4798) );
  NAND2_X1 U6423 ( .A1(n4806), .A2(n8401), .ZN(n8041) );
  NAND3_X1 U6424 ( .A1(n6013), .A2(n4376), .A3(n6014), .ZN(n8401) );
  NAND2_X1 U6425 ( .A1(n8299), .A2(n4811), .ZN(n4810) );
  INV_X1 U6426 ( .A(n8301), .ZN(n4815) );
  NAND2_X1 U6427 ( .A1(n8256), .A2(n4822), .ZN(n6408) );
  NAND3_X1 U6428 ( .A1(n4824), .A2(n4823), .A3(n8631), .ZN(n8256) );
  NAND2_X1 U6429 ( .A1(n6406), .A2(n6405), .ZN(n4823) );
  NAND2_X1 U6430 ( .A1(n4833), .A2(n6854), .ZN(n5810) );
  AOI22_X1 U6431 ( .A1(n7036), .A2(n4833), .B1(n9375), .B2(n7930), .ZN(n6924)
         );
  AOI21_X1 U6432 ( .B1(n10042), .B2(n4833), .A(n4831), .ZN(n10039) );
  AOI22_X1 U6433 ( .A1(n9768), .A2(P1_REG2_REG_2__SCAN_IN), .B1(n10038), .B2(
        n10046), .ZN(n4832) );
  XNOR2_X2 U6434 ( .A(n7544), .B(n7700), .ZN(n7699) );
  NAND2_X1 U6435 ( .A1(n7698), .A2(n7547), .ZN(n7545) );
  NAND2_X1 U6436 ( .A1(n7544), .A2(n7543), .ZN(n7547) );
  NAND2_X1 U6437 ( .A1(n4834), .A2(n7487), .ZN(n7182) );
  OR2_X2 U6438 ( .A1(n7181), .A2(n7264), .ZN(n4835) );
  AND2_X2 U6439 ( .A1(n4836), .A2(n4837), .ZN(n10010) );
  NAND2_X1 U6440 ( .A1(n6482), .A2(n7141), .ZN(n7138) );
  NOR2_X1 U6441 ( .A1(n10072), .A2(n6425), .ZN(n4837) );
  NAND2_X1 U6442 ( .A1(n7399), .A2(n4846), .ZN(n7308) );
  NAND2_X1 U6443 ( .A1(n4847), .A2(n8453), .ZN(n4849) );
  NAND2_X1 U6444 ( .A1(n4849), .A2(n4848), .ZN(n8469) );
  AOI21_X1 U6445 ( .B1(n8453), .B2(n4851), .A(n4850), .ZN(n4848) );
  NAND3_X1 U6446 ( .A1(n9799), .A2(n7744), .A3(n4854), .ZN(n9797) );
  INV_X1 U6447 ( .A(n4855), .ZN(n9795) );
  XNOR2_X1 U6448 ( .A(n8470), .B(n4856), .ZN(n8471) );
  AND2_X2 U6449 ( .A1(n4372), .A2(n7349), .ZN(n7578) );
  NAND2_X1 U6450 ( .A1(n9620), .A2(n9619), .ZN(n9843) );
  NAND2_X1 U6451 ( .A1(n4864), .A2(n5032), .ZN(n5293) );
  NAND2_X1 U6452 ( .A1(n5242), .A2(n5243), .ZN(n4864) );
  INV_X1 U6453 ( .A(n5243), .ZN(n4865) );
  INV_X1 U6454 ( .A(n5032), .ZN(n4866) );
  NAND2_X1 U6455 ( .A1(n9689), .A2(n6472), .ZN(n4875) );
  NAND2_X1 U6456 ( .A1(n5325), .A2(n5038), .ZN(n4878) );
  NAND2_X1 U6457 ( .A1(n6433), .A2(n6435), .ZN(n5774) );
  NAND2_X1 U6458 ( .A1(n5386), .A2(n5773), .ZN(n5775) );
  NAND3_X1 U6459 ( .A1(n5345), .A2(n5344), .A3(n9369), .ZN(n6435) );
  INV_X1 U6460 ( .A(n8598), .ZN(n4881) );
  NAND3_X1 U6461 ( .A1(n4325), .A2(n4887), .A3(n10189), .ZN(n8027) );
  AND2_X1 U6462 ( .A1(n4884), .A2(n4883), .ZN(n4887) );
  NAND2_X1 U6463 ( .A1(n4285), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n4886) );
  NAND3_X1 U6464 ( .A1(n4890), .A2(n8197), .A3(n8143), .ZN(n4889) );
  NAND3_X1 U6465 ( .A1(n8659), .A2(n4892), .A3(n8197), .ZN(n4891) );
  NAND2_X1 U6466 ( .A1(n6585), .A2(n4895), .ZN(n4898) );
  AND2_X1 U6467 ( .A1(n4899), .A2(n8062), .ZN(n4895) );
  NAND3_X1 U6468 ( .A1(n4899), .A2(n8062), .A3(n4901), .ZN(n4897) );
  NAND4_X1 U6469 ( .A1(n5913), .A2(n5917), .A3(n4284), .A4(n5896), .ZN(n6357)
         );
  NAND2_X1 U6470 ( .A1(n5905), .A2(n4906), .ZN(n4908) );
  XNOR2_X1 U6471 ( .A(n7042), .B(n4910), .ZN(n6935) );
  XNOR2_X1 U6472 ( .A(n7040), .B(n7039), .ZN(n4910) );
  NAND2_X1 U6473 ( .A1(n4911), .A2(n4912), .ZN(n9101) );
  NOR2_X1 U6474 ( .A1(n4468), .A2(n4976), .ZN(n9067) );
  OAI21_X2 U6475 ( .B1(n9239), .B2(n4918), .A(n4348), .ZN(n9325) );
  AND2_X2 U6476 ( .A1(n9325), .A2(n7975), .ZN(n9137) );
  NAND2_X1 U6477 ( .A1(n7059), .A2(n7058), .ZN(n7801) );
  NOR2_X1 U6478 ( .A1(n4925), .A2(n4921), .ZN(n4920) );
  NAND2_X1 U6479 ( .A1(n7801), .A2(n4929), .ZN(n4923) );
  NAND2_X1 U6480 ( .A1(n7804), .A2(n4928), .ZN(n4924) );
  NOR2_X1 U6481 ( .A1(n7804), .A2(n4926), .ZN(n4925) );
  NAND4_X2 U6482 ( .A1(n4938), .A2(n5271), .A3(n5272), .A4(n4937), .ZN(n9377)
         );
  NAND2_X1 U6483 ( .A1(n4939), .A2(n4942), .ZN(n7439) );
  NAND3_X1 U6484 ( .A1(n4943), .A2(n4945), .A3(n4944), .ZN(n4939) );
  NAND2_X1 U6485 ( .A1(n7248), .A2(n4946), .ZN(n4945) );
  NAND3_X1 U6486 ( .A1(n4945), .A2(n4944), .A3(n4947), .ZN(n7341) );
  NAND2_X1 U6487 ( .A1(n6446), .A2(n4952), .ZN(n4949) );
  NAND2_X1 U6488 ( .A1(n4949), .A2(n4950), .ZN(n9764) );
  NAND2_X1 U6489 ( .A1(n4958), .A2(n4960), .ZN(n7736) );
  NAND2_X1 U6490 ( .A1(n7504), .A2(n4961), .ZN(n4958) );
  INV_X1 U6491 ( .A(n4961), .ZN(n4959) );
  NAND2_X1 U6492 ( .A1(n6459), .A2(n6458), .ZN(n9676) );
  NOR2_X1 U6493 ( .A1(n4966), .A2(n6460), .ZN(n4965) );
  INV_X1 U6494 ( .A(n6458), .ZN(n4966) );
  NOR2_X1 U6495 ( .A1(n9680), .A2(n9328), .ZN(n4968) );
  NAND2_X1 U6496 ( .A1(n4970), .A2(n6462), .ZN(n9611) );
  NAND2_X1 U6497 ( .A1(n5165), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5166) );
  AND2_X1 U6498 ( .A1(n5876), .A2(n5875), .ZN(n5885) );
  INV_X1 U6499 ( .A(n7030), .ZN(n6482) );
  MUX2_X1 U6500 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5951), .S(
        P2_IR_REG_2__SCAN_IN), .Z(n5952) );
  XNOR2_X1 U6501 ( .A(n5190), .B(n5210), .ZN(n7048) );
  OAI21_X1 U6502 ( .B1(n5190), .B2(n5191), .A(n5209), .ZN(n5193) );
  OAI21_X1 U6503 ( .B1(n6514), .B2(n6513), .A(n4983), .ZN(P2_U3154) );
  CLKBUF_X1 U6504 ( .A(n8299), .Z(n8303) );
  NAND2_X1 U6505 ( .A1(n6295), .A2(n4981), .ZN(n6296) );
  OAI21_X1 U6506 ( .B1(n9856), .B2(n10088), .A(n9855), .ZN(n9935) );
  AND2_X1 U6507 ( .A1(n6614), .A2(n6368), .ZN(n6616) );
  INV_X1 U6508 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n6127) );
  NAND2_X1 U6509 ( .A1(n8238), .A2(n8237), .ZN(n9832) );
  NOR2_X1 U6510 ( .A1(n8516), .A2(n8515), .ZN(n8517) );
  AND2_X1 U6511 ( .A1(n9641), .A2(n6486), .ZN(n6487) );
  CLKBUF_X1 U6512 ( .A(n7560), .Z(n7561) );
  NOR2_X1 U6513 ( .A1(n9604), .A2(n8236), .ZN(n8237) );
  INV_X1 U6514 ( .A(n6849), .ZN(n6853) );
  OR2_X1 U6515 ( .A1(n9845), .A2(n9834), .ZN(n9847) );
  OAI211_X2 U6516 ( .C1(n6614), .C2(n6767), .A(n5910), .B(n5911), .ZN(n6517)
         );
  OR2_X1 U6517 ( .A1(n5310), .A2(n6808), .ZN(n5280) );
  NAND2_X1 U6518 ( .A1(n6523), .A2(n10195), .ZN(n8033) );
  AND2_X2 U6519 ( .A1(n5172), .A2(n4273), .ZN(n5309) );
  NAND2_X1 U6520 ( .A1(n8255), .A2(n9964), .ZN(n5312) );
  INV_X1 U6521 ( .A(n10175), .ZN(n8737) );
  AND2_X1 U6522 ( .A1(n6616), .A2(n8165), .ZN(n10175) );
  AND2_X1 U6523 ( .A1(n5004), .A2(n5489), .ZN(n4971) );
  AND2_X1 U6524 ( .A1(n6791), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n4972) );
  INV_X1 U6525 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5897) );
  INV_X1 U6526 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n8998) );
  NOR3_X1 U6527 ( .A1(n9838), .A2(n10088), .A3(n9837), .ZN(n4974) );
  OR2_X1 U6528 ( .A1(n4989), .A2(n7938), .ZN(n4975) );
  AND2_X1 U6529 ( .A1(n7810), .A2(n7809), .ZN(n4976) );
  AND2_X1 U6530 ( .A1(n8265), .A2(n8631), .ZN(n4977) );
  OR2_X1 U6531 ( .A1(n8763), .A2(n8391), .ZN(n4978) );
  AND2_X1 U6532 ( .A1(n6797), .A2(n4469), .ZN(n10035) );
  INV_X1 U6533 ( .A(n8684), .ZN(n6561) );
  AND2_X1 U6534 ( .A1(n5052), .A2(n5051), .ZN(n4979) );
  AND3_X1 U6535 ( .A1(n6294), .A2(n6293), .A3(n8288), .ZN(n4981) );
  OR2_X1 U6536 ( .A1(n8248), .A2(n8780), .ZN(n4982) );
  AND4_X2 U6537 ( .A1(n6897), .A2(n6898), .A3(n6650), .A4(n6649), .ZN(n10229)
         );
  AND2_X1 U6538 ( .A1(n6512), .A2(n6511), .ZN(n4983) );
  AND2_X1 U6539 ( .A1(n8219), .A2(n8819), .ZN(n4984) );
  AND2_X1 U6540 ( .A1(n5711), .A2(n5710), .ZN(n4985) );
  OR2_X1 U6541 ( .A1(n6407), .A2(n6260), .ZN(n4987) );
  AND3_X1 U6542 ( .A1(n8720), .A2(n6550), .A3(n8718), .ZN(n4988) );
  XOR2_X1 U6543 ( .A(n7929), .B(n4278), .Z(n4989) );
  AND2_X1 U6544 ( .A1(n9713), .A2(n9712), .ZN(n4990) );
  AND2_X1 U6545 ( .A1(n9728), .A2(n9727), .ZN(n4991) );
  INV_X2 U6546 ( .A(n10219), .ZN(n10217) );
  OR2_X1 U6547 ( .A1(n8248), .A2(n8845), .ZN(n4992) );
  OR2_X1 U6548 ( .A1(n9374), .A2(n10072), .ZN(n4993) );
  AOI211_X1 U6549 ( .C1(n5708), .C2(n9665), .A(n5631), .B(n5630), .ZN(n5632)
         );
  AND2_X1 U6550 ( .A1(n7983), .A2(n7714), .ZN(n6549) );
  NOR2_X1 U6551 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), .ZN(
        n5896) );
  INV_X1 U6552 ( .A(n6402), .ZN(n6403) );
  INV_X1 U6553 ( .A(n7890), .ZN(n7891) );
  NAND2_X1 U6554 ( .A1(n5663), .A2(n6468), .ZN(n5664) );
  NOR2_X1 U6555 ( .A1(n7572), .A2(n7573), .ZN(n5779) );
  AND2_X1 U6556 ( .A1(n8514), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n8515) );
  INV_X1 U6557 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n5398) );
  NAND2_X1 U6558 ( .A1(n5161), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n5562) );
  INV_X1 U6559 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n5513) );
  NOR2_X1 U6560 ( .A1(n9840), .A2(n10103), .ZN(n9841) );
  INV_X1 U6561 ( .A(n9784), .ZN(n5788) );
  INV_X1 U6562 ( .A(SI_27_), .ZN(n5134) );
  INV_X1 U6563 ( .A(SI_24_), .ZN(n5116) );
  INV_X1 U6564 ( .A(SI_20_), .ZN(n5532) );
  INV_X1 U6565 ( .A(SI_17_), .ZN(n5075) );
  INV_X1 U6566 ( .A(n7285), .ZN(n6037) );
  INV_X1 U6567 ( .A(n7006), .ZN(n5966) );
  AND2_X1 U6568 ( .A1(n6625), .A2(n6359), .ZN(n6378) );
  INV_X1 U6569 ( .A(n8011), .ZN(n6314) );
  NAND2_X1 U6570 ( .A1(n5934), .A2(n8907), .ZN(n5973) );
  INV_X1 U6571 ( .A(n8161), .ZN(n8162) );
  INV_X1 U6572 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n6239) );
  INV_X1 U6573 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n6098) );
  NAND2_X1 U6574 ( .A1(n6623), .A2(n4391), .ZN(n6624) );
  NAND2_X1 U6575 ( .A1(n8558), .A2(n8215), .ZN(n6900) );
  INV_X1 U6576 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5928) );
  NAND2_X1 U6577 ( .A1(n5163), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n5618) );
  NAND2_X1 U6578 ( .A1(n5305), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n5240) );
  OR2_X1 U6579 ( .A1(n9982), .A2(n9983), .ZN(n9979) );
  NOR2_X1 U6580 ( .A1(n4974), .A2(n9841), .ZN(n9842) );
  INV_X1 U6581 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5147) );
  INV_X1 U6582 ( .A(n5574), .ZN(n5114) );
  AND2_X1 U6583 ( .A1(n5081), .A2(n5080), .ZN(n5473) );
  OR2_X1 U6584 ( .A1(n5424), .A2(P1_IR_REG_12__SCAN_IN), .ZN(n5447) );
  NAND2_X1 U6585 ( .A1(n4283), .A2(n6657), .ZN(n5025) );
  INV_X1 U6586 ( .A(n6510), .ZN(n6511) );
  OR2_X1 U6587 ( .A1(n5973), .A2(n6762), .ZN(n5942) );
  OR2_X1 U6588 ( .A1(n6725), .A2(n8910), .ZN(n6760) );
  INV_X1 U6589 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n6652) );
  AND2_X1 U6590 ( .A1(n6365), .A2(n10216), .ZN(n6648) );
  INV_X1 U6591 ( .A(n6635), .ZN(n8248) );
  NAND2_X1 U6592 ( .A1(n8590), .A2(n8589), .ZN(n8591) );
  INV_X1 U6593 ( .A(n10178), .ZN(n8753) );
  AND2_X1 U6594 ( .A1(n6936), .A2(n6609), .ZN(n8756) );
  AND2_X1 U6595 ( .A1(n7052), .A2(n7051), .ZN(n7053) );
  INV_X1 U6596 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n9287) );
  XNOR2_X1 U6597 ( .A(n6924), .B(n9132), .ZN(n7039) );
  NOR2_X1 U6598 ( .A1(n6793), .A2(n6800), .ZN(n6803) );
  INV_X1 U6599 ( .A(n5312), .ZN(n5269) );
  OR2_X1 U6600 ( .A1(n7119), .A2(n7118), .ZN(n9526) );
  OR2_X1 U6601 ( .A1(n9557), .A2(n9558), .ZN(n9580) );
  INV_X1 U6602 ( .A(n10035), .ZN(n8236) );
  INV_X1 U6603 ( .A(n9893), .ZN(n9775) );
  AND2_X1 U6604 ( .A1(n6435), .A2(n6434), .ZN(n7336) );
  INV_X1 U6605 ( .A(n10072), .ZN(n7141) );
  INV_X1 U6606 ( .A(n9951), .ZN(n6800) );
  NAND2_X1 U6607 ( .A1(n9852), .A2(n9851), .ZN(n9853) );
  INV_X1 U6608 ( .A(n10030), .ZN(n10000) );
  OR2_X1 U6609 ( .A1(n9952), .A2(n6772), .ZN(n6501) );
  INV_X1 U6610 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n5168) );
  INV_X1 U6611 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5861) );
  INV_X1 U6612 ( .A(n8611), .ZN(n6606) );
  NAND2_X1 U6613 ( .A1(n6366), .A2(n8655), .ZN(n8362) );
  INV_X1 U6614 ( .A(n10164), .ZN(n10125) );
  INV_X1 U6615 ( .A(n8570), .ZN(n10166) );
  INV_X1 U6616 ( .A(n10170), .ZN(n10142) );
  INV_X1 U6617 ( .A(n8739), .ZN(n10173) );
  NAND2_X1 U6618 ( .A1(n10227), .A2(n8967), .ZN(n8767) );
  INV_X1 U6619 ( .A(n8780), .ZN(n8810) );
  AND2_X1 U6620 ( .A1(n6639), .A2(n6638), .ZN(n6897) );
  INV_X1 U6621 ( .A(n10201), .ZN(n10210) );
  OR2_X1 U6622 ( .A1(n6630), .A2(n6629), .ZN(n6631) );
  XNOR2_X1 U6623 ( .A(n6356), .B(n5897), .ZN(n6718) );
  AND2_X1 U6624 ( .A1(n6181), .A2(n6182), .ZN(n8562) );
  INV_X1 U6625 ( .A(n8905), .ZN(n8900) );
  INV_X1 U6626 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n5747) );
  INV_X1 U6627 ( .A(n7847), .ZN(n9178) );
  INV_X1 U6628 ( .A(n9167), .ZN(n9302) );
  INV_X1 U6629 ( .A(n9345), .ZN(n9335) );
  AND3_X1 U6630 ( .A1(n5683), .A2(n5682), .A3(n5681), .ZN(n8242) );
  AND4_X1 U6631 ( .A1(n5459), .A2(n5458), .A3(n5457), .A4(n5456), .ZN(n7864)
         );
  AND2_X1 U6632 ( .A1(n6838), .A2(n4281), .ZN(n9966) );
  AND2_X1 U6633 ( .A1(n5718), .A2(n5839), .ZN(n9778) );
  OAI21_X1 U6634 ( .B1(n9952), .B2(P1_D_REG_0__SCAN_IN), .A(n9954), .ZN(n7000)
         );
  AND2_X1 U6635 ( .A1(n7028), .A2(n6989), .ZN(n10088) );
  INV_X1 U6636 ( .A(n10088), .ZN(n10107) );
  AND2_X1 U6637 ( .A1(n6676), .A2(n5871), .ZN(n9951) );
  INV_X1 U6638 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n7649) );
  INV_X1 U6639 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n8977) );
  INV_X1 U6640 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n8955) );
  INV_X1 U6641 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n9539) );
  INV_X1 U6642 ( .A(n6702), .ZN(n6656) );
  INV_X1 U6643 ( .A(n8286), .ZN(n8846) );
  INV_X1 U6644 ( .A(n8367), .ZN(n8375) );
  AND2_X1 U6645 ( .A1(n8014), .A2(n6613), .ZN(n8017) );
  INV_X1 U6646 ( .A(n8621), .ZN(n8642) );
  INV_X1 U6647 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n10169) );
  NAND2_X1 U6648 ( .A1(n6761), .A2(n8564), .ZN(n10133) );
  NAND2_X1 U6649 ( .A1(n6909), .A2(n8757), .ZN(n8581) );
  INV_X1 U6650 ( .A(n8250), .ZN(n7498) );
  INV_X1 U6651 ( .A(n10186), .ZN(n10187) );
  INV_X1 U6652 ( .A(n8819), .ZN(n8763) );
  NAND2_X1 U6653 ( .A1(n10229), .A2(n10201), .ZN(n8813) );
  OR2_X1 U6654 ( .A1(n8711), .A2(n8710), .ZN(n8885) );
  OR2_X1 U6655 ( .A1(n10219), .A2(n8792), .ZN(n8845) );
  AND2_X1 U6656 ( .A1(n6632), .A2(n6631), .ZN(n10219) );
  INV_X1 U6657 ( .A(n6706), .ZN(n6707) );
  NAND2_X1 U6658 ( .A1(n6696), .A2(n6695), .ZN(n6706) );
  INV_X1 U6659 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7433) );
  INV_X1 U6660 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n7169) );
  INV_X1 U6661 ( .A(n9863), .ZN(n9680) );
  INV_X1 U6662 ( .A(n9348), .ZN(n9338) );
  INV_X1 U6663 ( .A(n9326), .ZN(n9350) );
  INV_X1 U6664 ( .A(n9231), .ZN(n9363) );
  OR2_X1 U6665 ( .A1(n6821), .A2(n6820), .ZN(n9986) );
  NAND2_X1 U6666 ( .A1(n6683), .A2(n6681), .ZN(n9995) );
  NAND2_X1 U6667 ( .A1(n9996), .A2(n10033), .ZN(n9828) );
  NAND2_X1 U6668 ( .A1(n10108), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n6503) );
  OR2_X1 U6669 ( .A1(n7001), .A2(n6776), .ZN(n10108) );
  INV_X1 U6670 ( .A(n10055), .ZN(n10056) );
  INV_X1 U6671 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7445) );
  INV_X1 U6672 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7799) );
  INV_X1 U6673 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n6859) );
  INV_X1 U6674 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n6705) );
  NOR2_X1 U6675 ( .A1(n7661), .A2(n7660), .ZN(n10249) );
  NOR2_X1 U6676 ( .A1(n7663), .A2(n7662), .ZN(n10247) );
  NOR2_X2 U6677 ( .A1(n6716), .A2(n6656), .ZN(P2_U3893) );
  AND2_X1 U6678 ( .A1(n6676), .A2(n6655), .ZN(P1_U3973) );
  NOR2_X1 U6679 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n4994) );
  INV_X1 U6680 ( .A(n5859), .ZN(n5000) );
  NOR2_X2 U6681 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n5141) );
  INV_X2 U6682 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5139) );
  NAND4_X1 U6683 ( .A1(n5139), .A2(n5001), .A3(n5004), .A4(n5489), .ZN(n5002)
         );
  NAND2_X1 U6684 ( .A1(n5741), .A2(n5742), .ZN(n5714) );
  NAND2_X1 U6685 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), 
        .ZN(n5003) );
  AND2_X1 U6686 ( .A1(n5003), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5010) );
  AND2_X1 U6687 ( .A1(n5168), .A2(P1_IR_REG_19__SCAN_IN), .ZN(n5009) );
  NAND2_X1 U6688 ( .A1(n5475), .A2(n5139), .ZN(n5488) );
  INV_X1 U6689 ( .A(n5488), .ZN(n5005) );
  AND2_X1 U6690 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), .ZN(
        n5006) );
  NAND2_X1 U6691 ( .A1(n5488), .A2(n5006), .ZN(n5007) );
  OAI211_X2 U6692 ( .C1(n5010), .C2(n5009), .A(n5008), .B(n5007), .ZN(n6783)
         );
  BUF_X4 U6693 ( .A(n6783), .Z(n9788) );
  INV_X2 U6694 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n5012) );
  INV_X2 U6695 ( .A(P1_RD_REG_SCAN_IN), .ZN(n5011) );
  NAND3_X2 U6696 ( .A1(n5013), .A2(n5012), .A3(n5011), .ZN(n5016) );
  NAND3_X2 U6697 ( .A1(n5014), .A2(P1_ADDR_REG_19__SCAN_IN), .A3(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n5015) );
  NAND2_X4 U6698 ( .A1(n5016), .A2(n5015), .ZN(n5259) );
  INV_X1 U6699 ( .A(n5259), .ZN(n5151) );
  AND2_X1 U6700 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n5017) );
  NAND2_X1 U6701 ( .A1(n5151), .A2(n5017), .ZN(n5947) );
  AND2_X1 U6702 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n5018) );
  NAND2_X1 U6703 ( .A1(n4282), .A2(n5018), .ZN(n5275) );
  NAND2_X1 U6704 ( .A1(n5947), .A2(n5275), .ZN(n5258) );
  INV_X1 U6705 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6660) );
  NAND2_X1 U6706 ( .A1(n5259), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n5020) );
  INV_X1 U6707 ( .A(SI_1_), .ZN(n5019) );
  OAI211_X1 U6708 ( .C1(n5259), .C2(n6660), .A(n5020), .B(n5019), .ZN(n5021)
         );
  NAND2_X1 U6709 ( .A1(n5258), .A2(n5021), .ZN(n5024) );
  INV_X1 U6710 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6689) );
  NAND2_X1 U6711 ( .A1(n4282), .A2(n6689), .ZN(n5022) );
  OAI211_X1 U6712 ( .C1(n5259), .C2(P1_DATAO_REG_1__SCAN_IN), .A(n5022), .B(
        SI_1_), .ZN(n5023) );
  NAND2_X1 U6713 ( .A1(n5024), .A2(n5023), .ZN(n5249) );
  INV_X1 U6714 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6668) );
  INV_X1 U6715 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6657) );
  XNOR2_X1 U6716 ( .A(n5026), .B(SI_2_), .ZN(n5250) );
  NAND2_X1 U6717 ( .A1(n5249), .A2(n5250), .ZN(n5029) );
  INV_X1 U6718 ( .A(n5026), .ZN(n5027) );
  NAND2_X1 U6719 ( .A1(n5027), .A2(SI_2_), .ZN(n5028) );
  INV_X1 U6720 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n9060) );
  INV_X1 U6721 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n8922) );
  MUX2_X1 U6722 ( .A(n9060), .B(n8922), .S(n4283), .Z(n5030) );
  INV_X1 U6723 ( .A(n5030), .ZN(n5031) );
  NAND2_X1 U6724 ( .A1(n5031), .A2(SI_3_), .ZN(n5032) );
  MUX2_X1 U6725 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .S(n5259), .Z(n5033) );
  XNOR2_X1 U6726 ( .A(n5033), .B(SI_4_), .ZN(n5294) );
  NAND2_X1 U6727 ( .A1(n5033), .A2(SI_4_), .ZN(n5034) );
  MUX2_X1 U6728 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .S(n4282), .Z(n5036) );
  XNOR2_X1 U6729 ( .A(n5036), .B(SI_5_), .ZN(n5317) );
  INV_X1 U6730 ( .A(n5317), .ZN(n5035) );
  NAND2_X1 U6731 ( .A1(n5036), .A2(SI_5_), .ZN(n5037) );
  MUX2_X1 U6732 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n4283), .Z(n5039) );
  XNOR2_X1 U6733 ( .A(n5039), .B(SI_6_), .ZN(n5326) );
  INV_X1 U6734 ( .A(n5326), .ZN(n5038) );
  NAND2_X1 U6735 ( .A1(n5039), .A2(SI_6_), .ZN(n5040) );
  MUX2_X1 U6736 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n5259), .Z(n5042) );
  XNOR2_X1 U6737 ( .A(n5042), .B(SI_7_), .ZN(n5370) );
  INV_X1 U6738 ( .A(n5370), .ZN(n5041) );
  MUX2_X1 U6739 ( .A(n6703), .B(n6705), .S(n4282), .Z(n5044) );
  INV_X1 U6740 ( .A(SI_8_), .ZN(n5043) );
  NAND2_X1 U6741 ( .A1(n5044), .A2(n5043), .ZN(n5047) );
  INV_X1 U6742 ( .A(n5044), .ZN(n5045) );
  NAND2_X1 U6743 ( .A1(n5045), .A2(SI_8_), .ZN(n5046) );
  NAND2_X1 U6744 ( .A1(n5047), .A2(n5046), .ZN(n5353) );
  MUX2_X1 U6745 ( .A(n6711), .B(n6709), .S(n4283), .Z(n5049) );
  INV_X1 U6746 ( .A(SI_9_), .ZN(n5048) );
  NAND2_X1 U6747 ( .A1(n5049), .A2(n5048), .ZN(n5052) );
  INV_X1 U6748 ( .A(n5049), .ZN(n5050) );
  NAND2_X1 U6749 ( .A1(n5050), .A2(SI_9_), .ZN(n5051) );
  MUX2_X1 U6750 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .S(n5259), .Z(n5054) );
  XNOR2_X1 U6751 ( .A(n5054), .B(SI_10_), .ZN(n5405) );
  NAND2_X1 U6752 ( .A1(n5054), .A2(SI_10_), .ZN(n5055) );
  MUX2_X1 U6753 ( .A(n6737), .B(n6739), .S(n5259), .Z(n5057) );
  NAND2_X1 U6754 ( .A1(n5057), .A2(n5056), .ZN(n5060) );
  INV_X1 U6755 ( .A(n5057), .ZN(n5058) );
  NAND2_X1 U6756 ( .A1(n5058), .A2(SI_11_), .ZN(n5059) );
  NAND2_X1 U6757 ( .A1(n5060), .A2(n5059), .ZN(n5394) );
  MUX2_X1 U6758 ( .A(n6869), .B(n6859), .S(n6658), .Z(n5061) );
  XNOR2_X1 U6759 ( .A(n5061), .B(SI_12_), .ZN(n5422) );
  INV_X1 U6760 ( .A(n5061), .ZN(n5062) );
  MUX2_X1 U6761 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n6658), .Z(n5064) );
  XNOR2_X1 U6762 ( .A(n5064), .B(SI_13_), .ZN(n5445) );
  INV_X1 U6763 ( .A(n5445), .ZN(n5063) );
  NAND2_X1 U6764 ( .A1(n5446), .A2(n5063), .ZN(n5221) );
  NAND2_X1 U6765 ( .A1(n5064), .A2(SI_13_), .ZN(n5220) );
  MUX2_X1 U6766 ( .A(n9000), .B(n7013), .S(n6658), .Z(n5066) );
  NAND2_X1 U6767 ( .A1(n5066), .A2(n5065), .ZN(n5071) );
  INV_X1 U6768 ( .A(n5066), .ZN(n5067) );
  NAND2_X1 U6769 ( .A1(n5067), .A2(SI_14_), .ZN(n5068) );
  NAND2_X1 U6770 ( .A1(n5071), .A2(n5068), .ZN(n5222) );
  INV_X1 U6771 ( .A(n5222), .ZN(n5069) );
  MUX2_X1 U6772 ( .A(n7092), .B(n7049), .S(n6658), .Z(n5209) );
  INV_X1 U6773 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n5072) );
  MUX2_X1 U6774 ( .A(n7167), .B(n5072), .S(n6658), .Z(n5194) );
  AOI22_X1 U6775 ( .A1(n5191), .A2(n5209), .B1(n5194), .B2(n5076), .ZN(n5073)
         );
  INV_X1 U6776 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n5074) );
  MUX2_X1 U6777 ( .A(n7222), .B(n5074), .S(n6658), .Z(n5090) );
  XNOR2_X1 U6778 ( .A(n5090), .B(SI_18_), .ZN(n5486) );
  MUX2_X1 U6779 ( .A(n7169), .B(n6734), .S(n6658), .Z(n5082) );
  NAND2_X1 U6780 ( .A1(n5082), .A2(n5075), .ZN(n5483) );
  NAND2_X1 U6781 ( .A1(n5486), .A2(n5483), .ZN(n5096) );
  OAI21_X1 U6782 ( .B1(n5209), .B2(n5191), .A(n5076), .ZN(n5078) );
  INV_X1 U6783 ( .A(n5194), .ZN(n5077) );
  NAND2_X1 U6784 ( .A1(n5078), .A2(n5077), .ZN(n5081) );
  INV_X1 U6785 ( .A(n5209), .ZN(n5079) );
  NAND3_X1 U6786 ( .A1(n5079), .A2(SI_16_), .A3(SI_15_), .ZN(n5080) );
  INV_X1 U6787 ( .A(n5473), .ZN(n5085) );
  INV_X1 U6788 ( .A(n5082), .ZN(n5083) );
  NAND2_X1 U6789 ( .A1(n5083), .A2(SI_17_), .ZN(n5474) );
  INV_X1 U6790 ( .A(n5474), .ZN(n5084) );
  NOR2_X1 U6791 ( .A1(n5085), .A2(n5084), .ZN(n5503) );
  INV_X1 U6792 ( .A(n5503), .ZN(n5094) );
  INV_X1 U6793 ( .A(n5096), .ZN(n5504) );
  MUX2_X1 U6794 ( .A(n7195), .B(n7799), .S(n6658), .Z(n5087) );
  NAND2_X1 U6795 ( .A1(n5087), .A2(n5086), .ZN(n5097) );
  INV_X1 U6796 ( .A(n5087), .ZN(n5088) );
  NAND2_X1 U6797 ( .A1(n5088), .A2(SI_19_), .ZN(n5089) );
  NAND2_X1 U6798 ( .A1(n5097), .A2(n5089), .ZN(n5508) );
  INV_X1 U6799 ( .A(n5508), .ZN(n5092) );
  INV_X1 U6800 ( .A(n5090), .ZN(n5091) );
  NAND2_X1 U6801 ( .A1(n5091), .A2(SI_18_), .ZN(n5506) );
  NAND2_X1 U6802 ( .A1(n5092), .A2(n5506), .ZN(n5093) );
  AOI21_X1 U6803 ( .B1(n5094), .B2(n5504), .A(n5093), .ZN(n5095) );
  MUX2_X1 U6804 ( .A(n7220), .B(n7225), .S(n6658), .Z(n5531) );
  INV_X1 U6805 ( .A(n5531), .ZN(n5101) );
  MUX2_X1 U6806 ( .A(n8981), .B(n7241), .S(n6658), .Z(n5536) );
  INV_X1 U6807 ( .A(n5536), .ZN(n5102) );
  OAI22_X1 U6808 ( .A1(n5101), .A2(SI_20_), .B1(n5102), .B2(SI_21_), .ZN(n5105) );
  INV_X1 U6809 ( .A(SI_21_), .ZN(n5099) );
  OAI21_X1 U6810 ( .B1(n5531), .B2(n5532), .A(n5099), .ZN(n5103) );
  AND2_X1 U6811 ( .A1(SI_21_), .A2(SI_20_), .ZN(n5100) );
  AOI22_X1 U6812 ( .A1(n5103), .A2(n5102), .B1(n5101), .B2(n5100), .ZN(n5104)
         );
  MUX2_X1 U6813 ( .A(n7297), .B(n9026), .S(n6658), .Z(n5107) );
  INV_X1 U6814 ( .A(SI_22_), .ZN(n5106) );
  NAND2_X1 U6815 ( .A1(n5107), .A2(n5106), .ZN(n5572) );
  INV_X1 U6816 ( .A(n5107), .ZN(n5108) );
  NAND2_X1 U6817 ( .A1(n5108), .A2(SI_22_), .ZN(n5109) );
  NAND2_X1 U6818 ( .A1(n5572), .A2(n5109), .ZN(n5558) );
  MUX2_X1 U6819 ( .A(n7375), .B(n5110), .S(n6658), .Z(n5112) );
  INV_X1 U6820 ( .A(SI_23_), .ZN(n5111) );
  NAND2_X1 U6821 ( .A1(n5112), .A2(n5111), .ZN(n5575) );
  AND2_X1 U6822 ( .A1(n5572), .A2(n5575), .ZN(n5115) );
  INV_X1 U6823 ( .A(n5112), .ZN(n5113) );
  NAND2_X1 U6824 ( .A1(n5113), .A2(SI_23_), .ZN(n5574) );
  MUX2_X1 U6825 ( .A(n7433), .B(n7445), .S(n6658), .Z(n5117) );
  NAND2_X1 U6826 ( .A1(n5117), .A2(n5116), .ZN(n5120) );
  INV_X1 U6827 ( .A(n5117), .ZN(n5118) );
  NAND2_X1 U6828 ( .A1(n5118), .A2(SI_24_), .ZN(n5119) );
  NAND2_X1 U6829 ( .A1(n5590), .A2(n5589), .ZN(n5121) );
  MUX2_X1 U6830 ( .A(n8983), .B(n7555), .S(n6658), .Z(n5123) );
  INV_X1 U6831 ( .A(SI_25_), .ZN(n5122) );
  NAND2_X1 U6832 ( .A1(n5123), .A2(n5122), .ZN(n5126) );
  INV_X1 U6833 ( .A(n5123), .ZN(n5124) );
  NAND2_X1 U6834 ( .A1(n5124), .A2(SI_25_), .ZN(n5125) );
  NAND2_X1 U6835 ( .A1(n5612), .A2(n5611), .ZN(n5127) );
  INV_X1 U6836 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n7585) );
  MUX2_X1 U6837 ( .A(n7686), .B(n7585), .S(n6658), .Z(n5129) );
  INV_X1 U6838 ( .A(SI_26_), .ZN(n5128) );
  NAND2_X1 U6839 ( .A1(n5129), .A2(n5128), .ZN(n5132) );
  INV_X1 U6840 ( .A(n5129), .ZN(n5130) );
  NAND2_X1 U6841 ( .A1(n5130), .A2(SI_26_), .ZN(n5131) );
  NAND2_X1 U6842 ( .A1(n5602), .A2(n5601), .ZN(n5133) );
  INV_X1 U6843 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n7695) );
  INV_X1 U6844 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n8002) );
  MUX2_X1 U6845 ( .A(n7695), .B(n8002), .S(n6658), .Z(n5135) );
  NAND2_X1 U6846 ( .A1(n5135), .A2(n5134), .ZN(n5138) );
  INV_X1 U6847 ( .A(n5135), .ZN(n5136) );
  NAND2_X1 U6848 ( .A1(n5136), .A2(SI_27_), .ZN(n5137) );
  INV_X1 U6849 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n8912) );
  INV_X1 U6850 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n8234) );
  MUX2_X1 U6851 ( .A(n8912), .B(n8234), .S(n6658), .Z(n5650) );
  XNOR2_X1 U6852 ( .A(n5650), .B(SI_28_), .ZN(n5647) );
  NOR2_X1 U6853 ( .A1(P1_IR_REG_25__SCAN_IN), .A2(P1_IR_REG_24__SCAN_IN), .ZN(
        n5142) );
  NOR2_X1 U6854 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .ZN(
        n5145) );
  NOR2_X1 U6855 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_20__SCAN_IN), .ZN(
        n5144) );
  NOR2_X1 U6856 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), .ZN(
        n5143) );
  NAND2_X1 U6858 ( .A1(n8909), .A2(n5694), .ZN(n5153) );
  NAND2_X1 U6859 ( .A1(n5603), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n5152) );
  INV_X1 U6860 ( .A(n5334), .ZN(n5154) );
  NAND2_X1 U6861 ( .A1(n5154), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5378) );
  INV_X1 U6862 ( .A(n5378), .ZN(n5155) );
  NAND2_X1 U6863 ( .A1(n5155), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5380) );
  INV_X1 U6864 ( .A(n5380), .ZN(n5156) );
  NAND2_X1 U6865 ( .A1(n5156), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n5363) );
  INV_X1 U6866 ( .A(n5363), .ZN(n5157) );
  NAND2_X1 U6867 ( .A1(n5157), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n5414) );
  INV_X1 U6868 ( .A(n5429), .ZN(n5158) );
  NAND2_X1 U6869 ( .A1(n5158), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n5452) );
  INV_X1 U6870 ( .A(n5452), .ZN(n5159) );
  NAND2_X1 U6871 ( .A1(n5159), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n5454) );
  INV_X1 U6872 ( .A(n5542), .ZN(n5161) );
  INV_X1 U6873 ( .A(n5593), .ZN(n5162) );
  INV_X1 U6874 ( .A(n5616), .ZN(n5163) );
  INV_X1 U6875 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n9331) );
  NAND2_X1 U6876 ( .A1(n5164), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n9616) );
  INV_X1 U6877 ( .A(n5169), .ZN(n9956) );
  NAND2_X1 U6878 ( .A1(n9639), .A2(n5654), .ZN(n5178) );
  INV_X1 U6879 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n5175) );
  NAND2_X1 U6880 ( .A1(n5620), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n5174) );
  NAND2_X1 U6881 ( .A1(n5657), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n5173) );
  OAI211_X1 U6882 ( .C1(n5175), .C2(n4685), .A(n5174), .B(n5173), .ZN(n5176)
         );
  INV_X1 U6883 ( .A(n5176), .ZN(n5177) );
  INV_X1 U6884 ( .A(n9612), .ZN(n9627) );
  OR2_X1 U6885 ( .A1(n9636), .A2(n9627), .ZN(n5790) );
  XNOR2_X1 U6886 ( .A(n5179), .B(n5180), .ZN(n7694) );
  NAND2_X1 U6887 ( .A1(n7694), .A2(n5694), .ZN(n5182) );
  NAND2_X1 U6888 ( .A1(n5603), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n5181) );
  INV_X1 U6889 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n5183) );
  NAND2_X1 U6890 ( .A1(n5607), .A2(n5183), .ZN(n5184) );
  NAND2_X1 U6891 ( .A1(n9616), .A2(n5184), .ZN(n9654) );
  INV_X1 U6892 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n9653) );
  INV_X2 U6893 ( .A(n4685), .ZN(n5656) );
  NAND2_X1 U6894 ( .A1(n5656), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n5186) );
  NAND2_X1 U6895 ( .A1(n5657), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n5185) );
  OAI211_X1 U6896 ( .C1(n9653), .C2(n5697), .A(n5186), .B(n5185), .ZN(n5187)
         );
  INV_X1 U6897 ( .A(n5187), .ZN(n5188) );
  NAND2_X1 U6898 ( .A1(n5790), .A2(n5761), .ZN(n5646) );
  NAND2_X1 U6899 ( .A1(n5190), .A2(n5191), .ZN(n5192) );
  NAND2_X1 U6900 ( .A1(n5193), .A2(n5192), .ZN(n5196) );
  XNOR2_X1 U6901 ( .A(n5194), .B(SI_16_), .ZN(n5195) );
  NAND2_X1 U6902 ( .A1(n7125), .A2(n5694), .ZN(n5200) );
  NAND2_X1 U6903 ( .A1(n5197), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5198) );
  XNOR2_X1 U6904 ( .A(n5198), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9578) );
  AOI22_X1 U6905 ( .A1(n5603), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n5510), .B2(
        n9578), .ZN(n5199) );
  NAND2_X1 U6906 ( .A1(n5656), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n5202) );
  NAND2_X1 U6907 ( .A1(n5657), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n5201) );
  AND2_X1 U6908 ( .A1(n5202), .A2(n5201), .ZN(n5208) );
  INV_X1 U6909 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n5204) );
  INV_X1 U6910 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n5203) );
  OAI21_X1 U6911 ( .B1(n5231), .B2(n5204), .A(n5203), .ZN(n5205) );
  NAND2_X1 U6912 ( .A1(n5478), .A2(n5205), .ZN(n9813) );
  OR2_X1 U6913 ( .A1(n9813), .A2(n5619), .ZN(n5207) );
  NAND2_X1 U6914 ( .A1(n5620), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n5206) );
  XNOR2_X1 U6915 ( .A(n5209), .B(SI_15_), .ZN(n5210) );
  NAND2_X1 U6916 ( .A1(n7048), .A2(n5694), .ZN(n5215) );
  OR2_X1 U6917 ( .A1(n5859), .A2(P1_IR_REG_9__SCAN_IN), .ZN(n5408) );
  INV_X1 U6918 ( .A(n5408), .ZN(n5212) );
  NAND2_X1 U6919 ( .A1(n5212), .A2(n5211), .ZN(n5410) );
  OAI21_X1 U6920 ( .B1(n5447), .B2(P1_IR_REG_13__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5225) );
  NAND2_X1 U6921 ( .A1(n5225), .A2(n5224), .ZN(n5227) );
  NAND2_X1 U6922 ( .A1(n5227), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5213) );
  XNOR2_X1 U6923 ( .A(n5213), .B(P1_IR_REG_15__SCAN_IN), .ZN(n9975) );
  AOI22_X1 U6924 ( .A1(n9975), .A2(n5510), .B1(n5603), .B2(
        P2_DATAO_REG_15__SCAN_IN), .ZN(n5214) );
  XNOR2_X1 U6925 ( .A(n5231), .B(P1_REG3_REG_15__SCAN_IN), .ZN(n9342) );
  NAND2_X1 U6926 ( .A1(n9342), .A2(n5654), .ZN(n5219) );
  NAND2_X1 U6927 ( .A1(n5656), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n5218) );
  NAND2_X1 U6928 ( .A1(n5620), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n5217) );
  NAND2_X1 U6929 ( .A1(n5657), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n5216) );
  NAND4_X1 U6930 ( .A1(n5219), .A2(n5218), .A3(n5217), .A4(n5216), .ZN(n9364)
         );
  INV_X1 U6931 ( .A(n9364), .ZN(n6441) );
  NAND2_X1 U6932 ( .A1(n9914), .A2(n6441), .ZN(n5782) );
  NAND2_X1 U6933 ( .A1(n9801), .A2(n5782), .ZN(n5468) );
  NAND2_X1 U6934 ( .A1(n5221), .A2(n5220), .ZN(n5223) );
  XNOR2_X1 U6935 ( .A(n5223), .B(n5222), .ZN(n7011) );
  NAND2_X1 U6936 ( .A1(n7011), .A2(n5694), .ZN(n5229) );
  OR2_X1 U6937 ( .A1(n5225), .A2(n5224), .ZN(n5226) );
  AOI22_X1 U6938 ( .A1(n5603), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n9550), .B2(
        n5510), .ZN(n5228) );
  NAND2_X1 U6939 ( .A1(n5656), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n5235) );
  NAND2_X1 U6940 ( .A1(n5620), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n5234) );
  NAND2_X1 U6941 ( .A1(n5454), .A2(n9081), .ZN(n5230) );
  AND2_X1 U6942 ( .A1(n5231), .A2(n5230), .ZN(n9086) );
  NAND2_X1 U6943 ( .A1(n5654), .A2(n9086), .ZN(n5233) );
  NAND2_X1 U6944 ( .A1(n5657), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5232) );
  NAND4_X1 U6945 ( .A1(n5235), .A2(n5234), .A3(n5233), .A4(n5232), .ZN(n9365)
         );
  INV_X1 U6946 ( .A(n9365), .ZN(n6439) );
  NAND2_X1 U6947 ( .A1(n5461), .A2(n6439), .ZN(n5463) );
  INV_X1 U6948 ( .A(n5463), .ZN(n5236) );
  INV_X1 U6949 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n5237) );
  NAND2_X1 U6950 ( .A1(n5309), .A2(n5237), .ZN(n5241) );
  INV_X1 U6951 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n6809) );
  OR2_X1 U6952 ( .A1(n5310), .A2(n6809), .ZN(n5239) );
  NAND2_X1 U6953 ( .A1(n5269), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n5238) );
  XNOR2_X1 U6954 ( .A(n5243), .B(n5242), .ZN(n9058) );
  NAND2_X1 U6955 ( .A1(n5613), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n5247) );
  INV_X1 U6956 ( .A(n5244), .ZN(n5295) );
  NAND2_X1 U6957 ( .A1(n5295), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5245) );
  XNOR2_X1 U6958 ( .A(n5245), .B(P1_IR_REG_3__SCAN_IN), .ZN(n9414) );
  NAND2_X1 U6959 ( .A1(n5323), .A2(n9414), .ZN(n5246) );
  NAND2_X1 U6960 ( .A1(n7038), .A2(n7043), .ZN(n7129) );
  NAND2_X1 U6961 ( .A1(n5305), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5281) );
  NAND2_X1 U6962 ( .A1(n5309), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n5282) );
  INV_X1 U6963 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n6808) );
  INV_X1 U6964 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n5248) );
  AND4_X2 U6965 ( .A1(n5281), .A2(n5282), .A3(n5280), .A4(n5283), .ZN(n6854)
         );
  XNOR2_X1 U6966 ( .A(n5249), .B(n5250), .ZN(n6667) );
  INV_X1 U6967 ( .A(n5251), .ZN(n5265) );
  NAND2_X1 U6968 ( .A1(n5265), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5252) );
  NAND2_X1 U6969 ( .A1(n5323), .A2(n9401), .ZN(n5253) );
  NAND2_X1 U6970 ( .A1(n7129), .A2(n5810), .ZN(n5285) );
  INV_X1 U6971 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n5254) );
  NAND2_X1 U6972 ( .A1(n5269), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n5256) );
  XNOR2_X1 U6973 ( .A(n5258), .B(SI_1_), .ZN(n5261) );
  MUX2_X1 U6974 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .S(n5259), .Z(n5260) );
  XNOR2_X1 U6975 ( .A(n5261), .B(n5260), .ZN(n6659) );
  AND2_X1 U6976 ( .A1(n8003), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n5262) );
  AOI21_X1 U6977 ( .B1(n6659), .B2(n6658), .A(n5262), .ZN(n5268) );
  INV_X1 U6978 ( .A(n9389), .ZN(n8240) );
  NAND2_X1 U6979 ( .A1(n8003), .A2(n6689), .ZN(n5263) );
  NAND2_X1 U6980 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5264) );
  INV_X1 U6981 ( .A(n6823), .ZN(n9380) );
  NAND3_X1 U6982 ( .A1(n8232), .A2(n9380), .A3(n4281), .ZN(n5266) );
  XNOR2_X1 U6983 ( .A(n6849), .B(n10043), .ZN(n5727) );
  NAND2_X1 U6984 ( .A1(n5269), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5272) );
  INV_X1 U6985 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n5270) );
  INV_X1 U6986 ( .A(SI_0_), .ZN(n5274) );
  INV_X1 U6987 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5273) );
  OAI21_X1 U6988 ( .B1(n8003), .B2(n5274), .A(n5273), .ZN(n5276) );
  AND2_X1 U6989 ( .A1(n5276), .A2(n5275), .ZN(n9965) );
  NAND2_X1 U6991 ( .A1(n5727), .A2(n6993), .ZN(n5279) );
  NAND2_X1 U6992 ( .A1(n6853), .A2(n10043), .ZN(n5278) );
  NAND4_X1 U6993 ( .A1(n5283), .A2(n5282), .A3(n5281), .A4(n5280), .ZN(n5284)
         );
  INV_X1 U6994 ( .A(n7038), .ZN(n6931) );
  NAND2_X1 U6995 ( .A1(n6931), .A2(n10066), .ZN(n5725) );
  INV_X1 U6996 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n5286) );
  XNOR2_X1 U6997 ( .A(n5286), .B(P1_REG3_REG_3__SCAN_IN), .ZN(n7139) );
  NAND2_X1 U6998 ( .A1(n5309), .A2(n7139), .ZN(n5288) );
  INV_X1 U6999 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n7137) );
  OR2_X1 U7000 ( .A1(n5697), .A2(n7137), .ZN(n5287) );
  INV_X1 U7001 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n5289) );
  OR2_X1 U7002 ( .A1(n5312), .A2(n5289), .ZN(n5291) );
  NAND2_X1 U7003 ( .A1(n5305), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5290) );
  XNOR2_X1 U7004 ( .A(n5293), .B(n5294), .ZN(n6665) );
  NAND2_X1 U7005 ( .A1(n5327), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5320) );
  XNOR2_X1 U7006 ( .A(n5320), .B(P1_IR_REG_4__SCAN_IN), .ZN(n9427) );
  AOI22_X1 U7007 ( .A1(n5613), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(n5510), .B2(
        n9427), .ZN(n5296) );
  NOR2_X1 U7008 ( .A1(n5297), .A2(n5708), .ZN(n5298) );
  INV_X1 U7009 ( .A(n7129), .ZN(n5299) );
  NAND2_X1 U7010 ( .A1(n5726), .A2(n5725), .ZN(n5815) );
  MUX2_X1 U7011 ( .A(n5299), .B(n5815), .S(n6468), .Z(n5300) );
  OR2_X1 U7012 ( .A1(n5301), .A2(n5300), .ZN(n5304) );
  INV_X1 U7013 ( .A(n5726), .ZN(n5302) );
  NAND2_X1 U7014 ( .A1(n5302), .A2(n5708), .ZN(n5303) );
  NAND2_X1 U7015 ( .A1(n5305), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5316) );
  INV_X1 U7016 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n5307) );
  NAND2_X1 U7017 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n5306) );
  NAND2_X1 U7018 ( .A1(n5307), .A2(n5306), .ZN(n5308) );
  AND2_X1 U7019 ( .A1(n5334), .A2(n5308), .ZN(n10018) );
  NAND2_X1 U7020 ( .A1(n5309), .A2(n10018), .ZN(n5315) );
  INV_X1 U7021 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n6813) );
  OR2_X1 U7022 ( .A1(n5310), .A2(n6813), .ZN(n5314) );
  INV_X1 U7023 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n5311) );
  OR2_X1 U7024 ( .A1(n5312), .A2(n5311), .ZN(n5313) );
  XNOR2_X1 U7025 ( .A(n5318), .B(n5317), .ZN(n6661) );
  INV_X1 U7026 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n5319) );
  NAND2_X1 U7027 ( .A1(n5320), .A2(n5319), .ZN(n5321) );
  NAND2_X1 U7028 ( .A1(n5321), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5322) );
  XNOR2_X1 U7029 ( .A(n5322), .B(P1_IR_REG_5__SCAN_IN), .ZN(n9441) );
  AOI22_X1 U7030 ( .A1(n5613), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n5510), .B2(
        n9441), .ZN(n5324) );
  NAND2_X1 U7031 ( .A1(n7209), .A2(n6425), .ZN(n5771) );
  XNOR2_X1 U7032 ( .A(n5325), .B(n5326), .ZN(n6663) );
  NAND2_X1 U7033 ( .A1(n6663), .A2(n5694), .ZN(n5332) );
  INV_X1 U7034 ( .A(n5327), .ZN(n5329) );
  NOR2_X1 U7035 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .ZN(
        n5328) );
  NAND2_X1 U7036 ( .A1(n5329), .A2(n5328), .ZN(n5355) );
  NAND2_X1 U7037 ( .A1(n5355), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5330) );
  XNOR2_X1 U7038 ( .A(n5330), .B(P1_IR_REG_6__SCAN_IN), .ZN(n9454) );
  AOI22_X1 U7039 ( .A1(n5613), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n5510), .B2(
        n9454), .ZN(n5331) );
  NAND2_X1 U7040 ( .A1(n5332), .A2(n5331), .ZN(n10083) );
  NAND2_X1 U7041 ( .A1(n5656), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n5340) );
  INV_X1 U7042 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n5333) );
  NAND2_X1 U7043 ( .A1(n5334), .A2(n5333), .ZN(n5335) );
  AND2_X1 U7044 ( .A1(n5378), .A2(n5335), .ZN(n9317) );
  NAND2_X1 U7045 ( .A1(n5654), .A2(n9317), .ZN(n5339) );
  INV_X1 U7046 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n5336) );
  OR2_X1 U7047 ( .A1(n5699), .A2(n5336), .ZN(n5338) );
  INV_X1 U7048 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n7213) );
  OR2_X1 U7049 ( .A1(n5697), .A2(n7213), .ZN(n5337) );
  OR2_X1 U7050 ( .A1(n10083), .A2(n9218), .ZN(n7242) );
  AND2_X1 U7051 ( .A1(n7242), .A2(n5819), .ZN(n5387) );
  NAND2_X1 U7052 ( .A1(n10083), .A2(n9218), .ZN(n6429) );
  NAND2_X1 U7053 ( .A1(n6708), .A2(n5694), .ZN(n5345) );
  NAND2_X1 U7054 ( .A1(n5859), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5343) );
  XNOR2_X1 U7055 ( .A(n5343), .B(P1_IR_REG_9__SCAN_IN), .ZN(n7110) );
  AOI22_X1 U7056 ( .A1(n5603), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n5510), .B2(
        n7110), .ZN(n5344) );
  NAND2_X1 U7057 ( .A1(n5656), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n5352) );
  INV_X1 U7058 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n5346) );
  NAND2_X1 U7059 ( .A1(n5363), .A2(n5346), .ZN(n5347) );
  AND2_X1 U7060 ( .A1(n5414), .A2(n5347), .ZN(n9257) );
  NAND2_X1 U7061 ( .A1(n5654), .A2(n9257), .ZN(n5351) );
  INV_X1 U7062 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n5348) );
  OR2_X1 U7063 ( .A1(n5699), .A2(n5348), .ZN(n5350) );
  INV_X1 U7064 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n7337) );
  OR2_X1 U7065 ( .A1(n5697), .A2(n7337), .ZN(n5349) );
  XNOR2_X1 U7066 ( .A(n5354), .B(n5353), .ZN(n6038) );
  NAND2_X1 U7067 ( .A1(n6038), .A2(n5694), .ZN(n5360) );
  INV_X1 U7068 ( .A(n5371), .ZN(n5356) );
  INV_X1 U7069 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n8935) );
  NAND2_X1 U7070 ( .A1(n5356), .A2(n8935), .ZN(n5373) );
  NAND2_X1 U7071 ( .A1(n5373), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5357) );
  MUX2_X1 U7072 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5357), .S(
        P1_IR_REG_8__SCAN_IN), .Z(n5358) );
  AND2_X1 U7073 ( .A1(n5358), .A2(n5859), .ZN(n9483) );
  AOI22_X1 U7074 ( .A1(n5613), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n5510), .B2(
        n9483), .ZN(n5359) );
  NAND2_X1 U7075 ( .A1(n5656), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5368) );
  INV_X1 U7076 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n5361) );
  NAND2_X1 U7077 ( .A1(n5380), .A2(n5361), .ZN(n5362) );
  AND2_X1 U7078 ( .A1(n5363), .A2(n5362), .ZN(n9153) );
  NAND2_X1 U7079 ( .A1(n5654), .A2(n9153), .ZN(n5367) );
  INV_X1 U7080 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n5364) );
  OR2_X1 U7081 ( .A1(n5699), .A2(n5364), .ZN(n5366) );
  INV_X1 U7082 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n6816) );
  OR2_X1 U7083 ( .A1(n5697), .A2(n6816), .ZN(n5365) );
  OR2_X1 U7084 ( .A1(n9157), .A2(n9069), .ZN(n6433) );
  INV_X1 U7085 ( .A(n5774), .ZN(n5386) );
  NAND2_X1 U7086 ( .A1(n6691), .A2(n5694), .ZN(n5376) );
  NAND2_X1 U7087 ( .A1(n5371), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5372) );
  MUX2_X1 U7088 ( .A(n5372), .B(P1_IR_REG_31__SCAN_IN), .S(n8935), .Z(n5374)
         );
  NAND2_X1 U7089 ( .A1(n5374), .A2(n5373), .ZN(n6832) );
  INV_X1 U7090 ( .A(n6832), .ZN(n9467) );
  AOI22_X1 U7091 ( .A1(n5603), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n5510), .B2(
        n9467), .ZN(n5375) );
  NAND2_X1 U7092 ( .A1(n5376), .A2(n5375), .ZN(n10007) );
  NAND2_X1 U7093 ( .A1(n5656), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n5385) );
  INV_X1 U7094 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n5377) );
  NAND2_X1 U7095 ( .A1(n5378), .A2(n5377), .ZN(n5379) );
  AND2_X1 U7096 ( .A1(n5380), .A2(n5379), .ZN(n10006) );
  NAND2_X1 U7097 ( .A1(n5654), .A2(n10006), .ZN(n5384) );
  INV_X1 U7098 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n6815) );
  OR2_X1 U7099 ( .A1(n5697), .A2(n6815), .ZN(n5383) );
  INV_X1 U7100 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n5381) );
  OR2_X1 U7101 ( .A1(n5699), .A2(n5381), .ZN(n5382) );
  OR2_X1 U7102 ( .A1(n10007), .A2(n7208), .ZN(n6431) );
  NAND2_X1 U7103 ( .A1(n5388), .A2(n7827), .ZN(n6434) );
  NAND2_X1 U7104 ( .A1(n10007), .A2(n7208), .ZN(n7244) );
  AND4_X1 U7105 ( .A1(n7322), .A2(n5708), .A3(n7244), .A4(n6429), .ZN(n5389)
         );
  NAND2_X1 U7106 ( .A1(n5773), .A2(n6468), .ZN(n5392) );
  AND2_X1 U7107 ( .A1(n6433), .A2(n6431), .ZN(n5724) );
  INV_X1 U7108 ( .A(n5724), .ZN(n5390) );
  NAND4_X1 U7109 ( .A1(n5390), .A2(n5708), .A3(n7322), .A4(n6434), .ZN(n5391)
         );
  OAI21_X1 U7110 ( .B1(n5774), .B2(n5392), .A(n5391), .ZN(n5393) );
  NAND2_X1 U7111 ( .A1(n6736), .A2(n5694), .ZN(n5397) );
  NAND2_X1 U7112 ( .A1(n5410), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5395) );
  XNOR2_X1 U7113 ( .A(n5395), .B(P1_IR_REG_11__SCAN_IN), .ZN(n9510) );
  AOI22_X1 U7114 ( .A1(n5603), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n5510), .B2(
        n9510), .ZN(n5396) );
  NAND2_X1 U7115 ( .A1(n5656), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n5404) );
  NAND2_X1 U7116 ( .A1(n5416), .A2(n5398), .ZN(n5399) );
  AND2_X1 U7117 ( .A1(n5429), .A2(n5399), .ZN(n9295) );
  NAND2_X1 U7118 ( .A1(n5654), .A2(n9295), .ZN(n5403) );
  INV_X1 U7119 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n7107) );
  OR2_X1 U7120 ( .A1(n5697), .A2(n7107), .ZN(n5402) );
  INV_X1 U7121 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n5400) );
  OR2_X1 U7122 ( .A1(n5699), .A2(n5400), .ZN(n5401) );
  NAND2_X1 U7123 ( .A1(n9299), .A2(n7834), .ZN(n5722) );
  INV_X1 U7124 ( .A(n5405), .ZN(n5406) );
  NAND2_X1 U7125 ( .A1(n6712), .A2(n5694), .ZN(n5413) );
  NAND2_X1 U7126 ( .A1(n5408), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5409) );
  MUX2_X1 U7127 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5409), .S(
        P1_IR_REG_10__SCAN_IN), .Z(n5411) );
  NAND2_X1 U7128 ( .A1(n5411), .A2(n5410), .ZN(n7113) );
  INV_X1 U7129 ( .A(n7113), .ZN(n9496) );
  AOI22_X1 U7130 ( .A1(n5603), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n5510), .B2(
        n9496), .ZN(n5412) );
  NAND2_X1 U7131 ( .A1(n5656), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n5421) );
  NAND2_X1 U7132 ( .A1(n5414), .A2(n9110), .ZN(n5415) );
  AND2_X1 U7133 ( .A1(n5416), .A2(n5415), .ZN(n9114) );
  NAND2_X1 U7134 ( .A1(n5654), .A2(n9114), .ZN(n5420) );
  INV_X1 U7135 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n5417) );
  OR2_X1 U7136 ( .A1(n5699), .A2(n5417), .ZN(n5419) );
  INV_X1 U7137 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n7105) );
  OR2_X1 U7138 ( .A1(n5697), .A2(n7105), .ZN(n5418) );
  NAND2_X1 U7139 ( .A1(n7841), .A2(n7326), .ZN(n7435) );
  AND2_X1 U7140 ( .A1(n5722), .A2(n7435), .ZN(n5822) );
  NAND2_X1 U7141 ( .A1(n5822), .A2(n6434), .ZN(n5437) );
  XNOR2_X1 U7142 ( .A(n5423), .B(n5422), .ZN(n6858) );
  NAND2_X1 U7143 ( .A1(n6858), .A2(n5694), .ZN(n5427) );
  NAND2_X1 U7144 ( .A1(n5424), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5425) );
  XNOR2_X1 U7145 ( .A(n5425), .B(P1_IR_REG_12__SCAN_IN), .ZN(n9524) );
  AOI22_X1 U7146 ( .A1(n5603), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n5510), .B2(
        n9524), .ZN(n5426) );
  NAND2_X1 U7147 ( .A1(n5656), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n5434) );
  NAND2_X1 U7148 ( .A1(n5657), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5433) );
  INV_X1 U7149 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n5428) );
  NAND2_X1 U7150 ( .A1(n5429), .A2(n5428), .ZN(n5430) );
  AND2_X1 U7151 ( .A1(n5452), .A2(n5430), .ZN(n9188) );
  NAND2_X1 U7152 ( .A1(n5654), .A2(n9188), .ZN(n5432) );
  NAND2_X1 U7153 ( .A1(n5620), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n5431) );
  NAND4_X1 U7154 ( .A1(n5434), .A2(n5433), .A3(n5432), .A4(n5431), .ZN(n9367)
         );
  NAND2_X1 U7155 ( .A1(n9191), .A2(n9367), .ZN(n5778) );
  OR2_X1 U7156 ( .A1(n7841), .A2(n7326), .ZN(n5723) );
  INV_X1 U7157 ( .A(n5723), .ZN(n5435) );
  NAND2_X1 U7158 ( .A1(n5822), .A2(n5435), .ZN(n5436) );
  AND3_X1 U7159 ( .A1(n5778), .A2(n5436), .A3(n7417), .ZN(n5806) );
  OAI21_X1 U7160 ( .B1(n5440), .B2(n5437), .A(n5806), .ZN(n5438) );
  INV_X1 U7161 ( .A(n9367), .ZN(n7854) );
  NAND2_X1 U7162 ( .A1(n9928), .A2(n7854), .ZN(n5826) );
  NAND2_X1 U7163 ( .A1(n5438), .A2(n5826), .ZN(n5444) );
  NAND2_X1 U7164 ( .A1(n5723), .A2(n6435), .ZN(n5439) );
  OAI21_X1 U7165 ( .B1(n5440), .B2(n5439), .A(n7435), .ZN(n5441) );
  NAND2_X1 U7166 ( .A1(n5441), .A2(n7417), .ZN(n5442) );
  XNOR2_X1 U7167 ( .A(n5446), .B(n5445), .ZN(n6919) );
  NAND2_X1 U7168 ( .A1(n6919), .A2(n5694), .ZN(n5450) );
  NAND2_X1 U7169 ( .A1(n5447), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5448) );
  XNOR2_X1 U7170 ( .A(n5448), .B(P1_IR_REG_13__SCAN_IN), .ZN(n9541) );
  AOI22_X1 U7171 ( .A1(n5603), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n5510), .B2(
        n9541), .ZN(n5449) );
  NAND2_X1 U7172 ( .A1(n5656), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n5459) );
  INV_X1 U7173 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n5451) );
  NAND2_X1 U7174 ( .A1(n5452), .A2(n5451), .ZN(n5453) );
  AND2_X1 U7175 ( .A1(n5454), .A2(n5453), .ZN(n9278) );
  NAND2_X1 U7176 ( .A1(n5654), .A2(n9278), .ZN(n5458) );
  INV_X1 U7177 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n5455) );
  OR2_X1 U7178 ( .A1(n5699), .A2(n5455), .ZN(n5457) );
  INV_X1 U7179 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n9534) );
  OR2_X1 U7180 ( .A1(n5697), .A2(n9534), .ZN(n5456) );
  NAND2_X1 U7181 ( .A1(n9922), .A2(n7864), .ZN(n5827) );
  NAND2_X1 U7182 ( .A1(n5462), .A2(n5827), .ZN(n5460) );
  OAI21_X1 U7183 ( .B1(n5830), .B2(n5460), .A(n5719), .ZN(n5466) );
  NAND2_X1 U7184 ( .A1(n5719), .A2(n5720), .ZN(n5835) );
  NOR2_X1 U7185 ( .A1(n5835), .A2(n5780), .ZN(n5465) );
  OR2_X1 U7186 ( .A1(n9922), .A2(n7864), .ZN(n5721) );
  NAND2_X1 U7187 ( .A1(n5462), .A2(n5721), .ZN(n5464) );
  NAND2_X1 U7188 ( .A1(n7737), .A2(n5463), .ZN(n7572) );
  INV_X1 U7189 ( .A(n5827), .ZN(n7573) );
  NOR2_X1 U7190 ( .A1(n9914), .A2(n6468), .ZN(n5467) );
  AOI21_X1 U7191 ( .B1(n5468), .B2(n5719), .A(n5467), .ZN(n5472) );
  AOI21_X1 U7192 ( .B1(n9801), .B2(n9364), .A(n6468), .ZN(n5471) );
  INV_X1 U7193 ( .A(n5721), .ZN(n5469) );
  NOR2_X1 U7194 ( .A1(n5780), .A2(n5469), .ZN(n5832) );
  OR3_X1 U7195 ( .A1(n5830), .A2(n5832), .A3(n6468), .ZN(n5470) );
  OAI21_X1 U7196 ( .B1(n5472), .B2(n5471), .A(n5470), .ZN(n5482) );
  NAND2_X1 U7197 ( .A1(n5502), .A2(n5473), .ZN(n5485) );
  NAND2_X1 U7198 ( .A1(n5483), .A2(n5474), .ZN(n5484) );
  XNOR2_X1 U7199 ( .A(n5485), .B(n5484), .ZN(n7155) );
  NAND2_X1 U7200 ( .A1(n7155), .A2(n5694), .ZN(n5477) );
  XNOR2_X1 U7201 ( .A(n5475), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9592) );
  AOI22_X1 U7202 ( .A1(n5603), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n5510), .B2(
        n9592), .ZN(n5476) );
  NAND2_X1 U7203 ( .A1(n5478), .A2(n9233), .ZN(n5479) );
  NAND2_X1 U7204 ( .A1(n5496), .A2(n5479), .ZN(n9807) );
  AOI22_X1 U7205 ( .A1(n5620), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n5656), .B2(
        P1_REG1_REG_17__SCAN_IN), .ZN(n5481) );
  NAND2_X1 U7206 ( .A1(n5657), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n5480) );
  OAI211_X1 U7207 ( .C1(n9807), .C2(n5619), .A(n5481), .B(n5480), .ZN(n9362)
         );
  INV_X1 U7208 ( .A(n9362), .ZN(n6444) );
  OR2_X1 U7209 ( .A1(n9903), .A2(n6444), .ZN(n5786) );
  NAND2_X1 U7210 ( .A1(n9903), .A2(n6444), .ZN(n5501) );
  NAND2_X1 U7211 ( .A1(n5786), .A2(n5501), .ZN(n5784) );
  OAI21_X1 U7212 ( .B1(n5485), .B2(n5484), .A(n5483), .ZN(n5487) );
  XNOR2_X1 U7213 ( .A(n5487), .B(n5486), .ZN(n7192) );
  NAND2_X1 U7214 ( .A1(n7192), .A2(n5694), .ZN(n5494) );
  NAND2_X1 U7215 ( .A1(n5488), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5490) );
  OR2_X1 U7216 ( .A1(n5490), .A2(n5489), .ZN(n5492) );
  NAND2_X1 U7217 ( .A1(n5490), .A2(n5489), .ZN(n5491) );
  AOI22_X1 U7218 ( .A1(n5603), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n5510), .B2(
        n9991), .ZN(n5493) );
  INV_X1 U7219 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n5500) );
  INV_X1 U7220 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n5495) );
  NAND2_X1 U7221 ( .A1(n5496), .A2(n5495), .ZN(n5497) );
  NAND2_X1 U7222 ( .A1(n5514), .A2(n5497), .ZN(n9790) );
  OR2_X1 U7223 ( .A1(n9790), .A2(n5619), .ZN(n5499) );
  AOI22_X1 U7224 ( .A1(n5620), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n5656), .B2(
        P1_REG1_REG_18__SCAN_IN), .ZN(n5498) );
  OAI211_X1 U7225 ( .C1(n5699), .C2(n5500), .A(n5499), .B(n5498), .ZN(n9361)
         );
  INV_X1 U7226 ( .A(n9361), .ZN(n9232) );
  NAND2_X1 U7227 ( .A1(n9898), .A2(n9232), .ZN(n5789) );
  AND2_X1 U7228 ( .A1(n5789), .A2(n5501), .ZN(n5836) );
  OR2_X1 U7229 ( .A1(n9898), .A2(n9232), .ZN(n5734) );
  NAND2_X1 U7230 ( .A1(n5502), .A2(n5503), .ZN(n5505) );
  NAND2_X1 U7231 ( .A1(n5505), .A2(n5504), .ZN(n5507) );
  NAND2_X1 U7232 ( .A1(n5507), .A2(n5506), .ZN(n5509) );
  XNOR2_X1 U7233 ( .A(n5509), .B(n5508), .ZN(n7194) );
  NAND2_X1 U7234 ( .A1(n7194), .A2(n5694), .ZN(n5512) );
  AOI22_X1 U7235 ( .A1(n5603), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n9630), .B2(
        n5510), .ZN(n5511) );
  NAND2_X1 U7236 ( .A1(n5514), .A2(n5513), .ZN(n5515) );
  AND2_X1 U7237 ( .A1(n5524), .A2(n5515), .ZN(n9773) );
  NAND2_X1 U7238 ( .A1(n9773), .A2(n5654), .ZN(n5520) );
  INV_X1 U7239 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n9590) );
  NAND2_X1 U7240 ( .A1(n5656), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n5517) );
  NAND2_X1 U7241 ( .A1(n5657), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n5516) );
  OAI211_X1 U7242 ( .C1(n5697), .C2(n9590), .A(n5517), .B(n5516), .ZN(n5518)
         );
  INV_X1 U7243 ( .A(n5518), .ZN(n5519) );
  NAND2_X1 U7244 ( .A1(n5520), .A2(n5519), .ZN(n9360) );
  INV_X1 U7245 ( .A(n9360), .ZN(n6450) );
  OR2_X1 U7246 ( .A1(n9893), .A2(n6450), .ZN(n5718) );
  NAND2_X1 U7247 ( .A1(n5734), .A2(n5718), .ZN(n5840) );
  AOI21_X1 U7248 ( .B1(n5552), .B2(n5836), .A(n5840), .ZN(n5551) );
  XNOR2_X1 U7249 ( .A(n5531), .B(SI_20_), .ZN(n5521) );
  XNOR2_X1 U7250 ( .A(n5533), .B(n5521), .ZN(n7219) );
  NAND2_X1 U7251 ( .A1(n7219), .A2(n5694), .ZN(n5523) );
  NAND2_X1 U7252 ( .A1(n5603), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n5522) );
  INV_X1 U7253 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n9266) );
  NAND2_X1 U7254 ( .A1(n5524), .A2(n9266), .ZN(n5525) );
  NAND2_X1 U7255 ( .A1(n5542), .A2(n5525), .ZN(n9762) );
  OR2_X1 U7256 ( .A1(n9762), .A2(n5619), .ZN(n5530) );
  INV_X1 U7257 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n9023) );
  NAND2_X1 U7258 ( .A1(n5656), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n5527) );
  NAND2_X1 U7259 ( .A1(n5620), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n5526) );
  OAI211_X1 U7260 ( .C1(n9023), .C2(n5699), .A(n5527), .B(n5526), .ZN(n5528)
         );
  INV_X1 U7261 ( .A(n5528), .ZN(n5529) );
  NAND2_X1 U7262 ( .A1(n9888), .A2(n9123), .ZN(n9737) );
  NAND2_X1 U7263 ( .A1(n9738), .A2(n9737), .ZN(n9763) );
  AOI22_X1 U7264 ( .A1(n4479), .A2(n9775), .B1(n9737), .B2(n9360), .ZN(n5550)
         );
  OAI21_X1 U7265 ( .B1(n5533), .B2(n5532), .A(n5531), .ZN(n5535) );
  NAND2_X1 U7266 ( .A1(n5533), .A2(n5532), .ZN(n5534) );
  NAND2_X1 U7267 ( .A1(n5535), .A2(n5534), .ZN(n5538) );
  XNOR2_X1 U7268 ( .A(n5536), .B(SI_21_), .ZN(n5537) );
  XNOR2_X1 U7269 ( .A(n5538), .B(n5537), .ZN(n7226) );
  NAND2_X1 U7270 ( .A1(n7226), .A2(n5694), .ZN(n5540) );
  NAND2_X1 U7271 ( .A1(n5603), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n5539) );
  INV_X1 U7272 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n5541) );
  NAND2_X1 U7273 ( .A1(n5542), .A2(n5541), .ZN(n5543) );
  NAND2_X1 U7274 ( .A1(n5562), .A2(n5543), .ZN(n9160) );
  OR2_X1 U7275 ( .A1(n9160), .A2(n5619), .ZN(n5549) );
  INV_X1 U7276 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n5546) );
  NAND2_X1 U7277 ( .A1(n5656), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n5545) );
  NAND2_X1 U7278 ( .A1(n5657), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n5544) );
  OAI211_X1 U7279 ( .C1(n5546), .C2(n5697), .A(n5545), .B(n5544), .ZN(n5547)
         );
  INV_X1 U7280 ( .A(n5547), .ZN(n5548) );
  AND2_X1 U7281 ( .A1(n5753), .A2(n9738), .ZN(n6469) );
  OAI21_X1 U7282 ( .B1(n5551), .B2(n5550), .A(n6469), .ZN(n5557) );
  AND2_X1 U7283 ( .A1(n5734), .A2(n5786), .ZN(n5805) );
  NAND2_X1 U7284 ( .A1(n5552), .A2(n5805), .ZN(n5553) );
  NAND2_X1 U7285 ( .A1(n9893), .A2(n6450), .ZN(n5839) );
  NAND2_X1 U7286 ( .A1(n9882), .A2(n9285), .ZN(n5735) );
  NAND2_X1 U7287 ( .A1(n5735), .A2(n9737), .ZN(n5754) );
  INV_X1 U7288 ( .A(n5754), .ZN(n5554) );
  NAND2_X1 U7289 ( .A1(n5555), .A2(n5554), .ZN(n5556) );
  MUX2_X1 U7290 ( .A(n5735), .B(n5753), .S(n5708), .Z(n5570) );
  XNOR2_X1 U7291 ( .A(n5559), .B(n5558), .ZN(n7294) );
  NAND2_X1 U7292 ( .A1(n7294), .A2(n5694), .ZN(n5561) );
  NAND2_X1 U7293 ( .A1(n5613), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n5560) );
  NAND2_X1 U7294 ( .A1(n5562), .A2(n9287), .ZN(n5563) );
  NAND2_X1 U7295 ( .A1(n5581), .A2(n5563), .ZN(n9722) );
  OR2_X1 U7296 ( .A1(n9722), .A2(n5619), .ZN(n5568) );
  INV_X1 U7297 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n9041) );
  NAND2_X1 U7298 ( .A1(n5620), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n5565) );
  NAND2_X1 U7299 ( .A1(n5656), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n5564) );
  OAI211_X1 U7300 ( .C1(n9041), .C2(n5699), .A(n5565), .B(n5564), .ZN(n5566)
         );
  INV_X1 U7301 ( .A(n5566), .ZN(n5567) );
  INV_X1 U7302 ( .A(n9357), .ZN(n9094) );
  OR2_X1 U7303 ( .A1(n9878), .A2(n9094), .ZN(n9712) );
  NAND2_X1 U7304 ( .A1(n9878), .A2(n9094), .ZN(n5638) );
  INV_X1 U7305 ( .A(n9727), .ZN(n5569) );
  NAND2_X1 U7306 ( .A1(n5573), .A2(n5572), .ZN(n5578) );
  AND2_X1 U7307 ( .A1(n5575), .A2(n5574), .ZN(n5577) );
  NAND2_X1 U7308 ( .A1(n5578), .A2(n5577), .ZN(n5576) );
  NAND2_X1 U7309 ( .A1(n7372), .A2(n5694), .ZN(n5580) );
  NAND2_X1 U7310 ( .A1(n5613), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n5579) );
  NAND2_X1 U7311 ( .A1(n5581), .A2(n9096), .ZN(n5582) );
  AND2_X1 U7312 ( .A1(n5593), .A2(n5582), .ZN(n9709) );
  NAND2_X1 U7313 ( .A1(n9709), .A2(n5654), .ZN(n5588) );
  INV_X1 U7314 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n5585) );
  NAND2_X1 U7315 ( .A1(n5656), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n5584) );
  NAND2_X1 U7316 ( .A1(n5657), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n5583) );
  OAI211_X1 U7317 ( .C1(n5585), .C2(n5697), .A(n5584), .B(n5583), .ZN(n5586)
         );
  INV_X1 U7318 ( .A(n5586), .ZN(n5587) );
  OR2_X1 U7319 ( .A1(n9873), .A2(n9286), .ZN(n5717) );
  NAND2_X1 U7320 ( .A1(n5717), .A2(n9712), .ZN(n5750) );
  NAND2_X1 U7321 ( .A1(n9636), .A2(n9627), .ZN(n9621) );
  NAND2_X1 U7322 ( .A1(n9850), .A2(n9330), .ZN(n6476) );
  XNOR2_X1 U7323 ( .A(n5590), .B(n5589), .ZN(n7432) );
  NAND2_X1 U7324 ( .A1(n7432), .A2(n5694), .ZN(n5592) );
  NAND2_X1 U7325 ( .A1(n5613), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n5591) );
  INV_X1 U7326 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n9243) );
  NAND2_X1 U7327 ( .A1(n5593), .A2(n9243), .ZN(n5594) );
  NAND2_X1 U7328 ( .A1(n5616), .A2(n5594), .ZN(n9698) );
  OR2_X1 U7329 ( .A1(n9698), .A2(n5619), .ZN(n5599) );
  INV_X1 U7330 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n8980) );
  NAND2_X1 U7331 ( .A1(n5656), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n5596) );
  NAND2_X1 U7332 ( .A1(n5620), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n5595) );
  OAI211_X1 U7333 ( .C1(n5699), .C2(n8980), .A(n5596), .B(n5595), .ZN(n5597)
         );
  INV_X1 U7334 ( .A(n5597), .ZN(n5598) );
  OR2_X1 U7335 ( .A1(n9869), .A2(n9095), .ZN(n6471) );
  NAND2_X1 U7336 ( .A1(n9869), .A2(n9095), .ZN(n5756) );
  NAND2_X1 U7337 ( .A1(n6471), .A2(n5756), .ZN(n9691) );
  NAND2_X1 U7338 ( .A1(n9873), .A2(n9286), .ZN(n9690) );
  INV_X1 U7339 ( .A(n9690), .ZN(n5600) );
  NOR2_X1 U7340 ( .A1(n9691), .A2(n5600), .ZN(n6472) );
  NAND2_X1 U7341 ( .A1(n7584), .A2(n5694), .ZN(n5605) );
  NAND2_X1 U7342 ( .A1(n5603), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n5604) );
  NAND2_X1 U7343 ( .A1(n5618), .A2(n9331), .ZN(n5606) );
  INV_X1 U7344 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n9017) );
  NAND2_X1 U7345 ( .A1(n5620), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n5609) );
  NAND2_X1 U7346 ( .A1(n5657), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n5608) );
  OAI211_X1 U7347 ( .C1(n4685), .C2(n9017), .A(n5609), .B(n5608), .ZN(n5610)
         );
  AOI21_X2 U7348 ( .B1(n9670), .B2(n5654), .A(n5610), .ZN(n9196) );
  NAND2_X1 U7349 ( .A1(n9859), .A2(n9196), .ZN(n5627) );
  XNOR2_X1 U7350 ( .A(n5612), .B(n5611), .ZN(n7520) );
  NAND2_X1 U7351 ( .A1(n7520), .A2(n5694), .ZN(n5615) );
  NAND2_X1 U7352 ( .A1(n5613), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n5614) );
  INV_X1 U7353 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n9199) );
  NAND2_X1 U7354 ( .A1(n5616), .A2(n9199), .ZN(n5617) );
  NAND2_X1 U7355 ( .A1(n5618), .A2(n5617), .ZN(n9677) );
  INV_X1 U7356 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n9042) );
  NAND2_X1 U7357 ( .A1(n5620), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n5622) );
  NAND2_X1 U7358 ( .A1(n5656), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n5621) );
  OAI211_X1 U7359 ( .C1(n9042), .C2(n5699), .A(n5622), .B(n5621), .ZN(n5623)
         );
  INV_X1 U7360 ( .A(n5623), .ZN(n5624) );
  AND2_X1 U7361 ( .A1(n9863), .A2(n9328), .ZN(n6473) );
  INV_X1 U7362 ( .A(n6473), .ZN(n5628) );
  NAND2_X1 U7363 ( .A1(n5627), .A2(n5628), .ZN(n5626) );
  OR2_X1 U7364 ( .A1(n9859), .A2(n9196), .ZN(n5749) );
  NAND2_X1 U7365 ( .A1(n5626), .A2(n5749), .ZN(n5635) );
  NAND4_X1 U7366 ( .A1(n5642), .A2(n6472), .A3(n5708), .A4(n5635), .ZN(n5637)
         );
  INV_X1 U7367 ( .A(n5627), .ZN(n6475) );
  AOI21_X1 U7368 ( .B1(n6474), .B2(n5749), .A(n6475), .ZN(n5640) );
  NAND2_X1 U7369 ( .A1(n5749), .A2(n5627), .ZN(n9665) );
  INV_X1 U7370 ( .A(n9681), .ZN(n5738) );
  NOR3_X1 U7371 ( .A1(n9702), .A2(n5708), .A3(n9355), .ZN(n5629) );
  NOR3_X1 U7372 ( .A1(n9665), .A2(n5738), .A3(n5629), .ZN(n5633) );
  NOR3_X1 U7373 ( .A1(n9869), .A2(n9095), .A3(n6468), .ZN(n5631) );
  NOR2_X1 U7374 ( .A1(n9681), .A2(n6468), .ZN(n5630) );
  OAI21_X1 U7375 ( .B1(n5640), .B2(n5633), .A(n5632), .ZN(n5634) );
  OAI211_X1 U7376 ( .C1(n6468), .C2(n5635), .A(n5634), .B(n5642), .ZN(n5636)
         );
  AND2_X1 U7377 ( .A1(n9690), .A2(n5638), .ZN(n5755) );
  INV_X1 U7378 ( .A(n9691), .ZN(n9688) );
  NAND3_X1 U7379 ( .A1(n9688), .A2(n6468), .A3(n5717), .ZN(n5641) );
  INV_X1 U7380 ( .A(n5642), .ZN(n5760) );
  INV_X1 U7381 ( .A(n6476), .ZN(n5643) );
  NAND2_X1 U7382 ( .A1(n5643), .A2(n6468), .ZN(n5644) );
  NAND2_X1 U7383 ( .A1(n4352), .A2(n5644), .ZN(n5645) );
  INV_X1 U7384 ( .A(SI_28_), .ZN(n5649) );
  MUX2_X1 U7385 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(P1_DATAO_REG_29__SCAN_IN), 
        .S(n8003), .Z(n5685) );
  INV_X1 U7386 ( .A(SI_29_), .ZN(n5651) );
  NAND2_X1 U7387 ( .A1(n8904), .A2(n5694), .ZN(n5653) );
  NAND2_X1 U7388 ( .A1(n5603), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n5652) );
  NAND2_X1 U7389 ( .A1(n5654), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n5655) );
  OR2_X1 U7390 ( .A1(n9616), .A2(n5655), .ZN(n5662) );
  INV_X1 U7391 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n9614) );
  NAND2_X1 U7392 ( .A1(n5656), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n5659) );
  NAND2_X1 U7393 ( .A1(n5657), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n5658) );
  OAI211_X1 U7394 ( .C1(n9614), .C2(n5697), .A(n5659), .B(n5658), .ZN(n5660)
         );
  INV_X1 U7395 ( .A(n5660), .ZN(n5661) );
  NAND2_X1 U7396 ( .A1(n9839), .A2(n7171), .ZN(n5793) );
  INV_X1 U7397 ( .A(n9621), .ZN(n5663) );
  NAND2_X1 U7398 ( .A1(n9836), .A2(n5664), .ZN(n5665) );
  INV_X1 U7399 ( .A(n5793), .ZN(n5704) );
  MUX2_X1 U7400 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n8003), .Z(n5668) );
  NAND2_X1 U7401 ( .A1(n5668), .A2(SI_30_), .ZN(n5691) );
  NAND2_X1 U7402 ( .A1(n5685), .A2(SI_29_), .ZN(n5667) );
  NAND3_X1 U7403 ( .A1(n5687), .A2(n5691), .A3(n5667), .ZN(n5674) );
  NOR2_X1 U7404 ( .A1(n5685), .A2(SI_29_), .ZN(n5672) );
  INV_X1 U7405 ( .A(n5668), .ZN(n5670) );
  INV_X1 U7406 ( .A(SI_30_), .ZN(n5669) );
  NAND2_X1 U7407 ( .A1(n5670), .A2(n5669), .ZN(n5690) );
  INV_X1 U7408 ( .A(n5690), .ZN(n5671) );
  AOI21_X1 U7409 ( .B1(n5672), .B2(n5691), .A(n5671), .ZN(n5673) );
  MUX2_X1 U7410 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n8003), .Z(n5675) );
  XNOR2_X1 U7411 ( .A(n5675), .B(SI_31_), .ZN(n5676) );
  NAND2_X1 U7412 ( .A1(n5603), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n5679) );
  NAND2_X1 U7413 ( .A1(n5656), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n5683) );
  INV_X1 U7414 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n9606) );
  OR2_X1 U7415 ( .A1(n5697), .A2(n9606), .ZN(n5682) );
  INV_X1 U7416 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n5680) );
  OR2_X1 U7417 ( .A1(n5699), .A2(n5680), .ZN(n5681) );
  AND2_X1 U7418 ( .A1(n4735), .A2(n8242), .ZN(n5716) );
  NAND2_X1 U7419 ( .A1(n5684), .A2(SI_29_), .ZN(n5689) );
  INV_X1 U7420 ( .A(n5685), .ZN(n5686) );
  OR2_X1 U7421 ( .A1(n5687), .A2(n5686), .ZN(n5688) );
  NAND2_X1 U7422 ( .A1(n5691), .A2(n5690), .ZN(n5692) );
  NAND2_X1 U7423 ( .A1(n8252), .A2(n5694), .ZN(n5696) );
  NAND2_X1 U7424 ( .A1(n5603), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n5695) );
  NAND2_X1 U7425 ( .A1(n5656), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n5702) );
  INV_X1 U7426 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n8239) );
  OR2_X1 U7427 ( .A1(n5697), .A2(n8239), .ZN(n5701) );
  INV_X1 U7428 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n5698) );
  OR2_X1 U7429 ( .A1(n5699), .A2(n5698), .ZN(n5700) );
  AND3_X1 U7430 ( .A1(n5702), .A2(n5701), .A3(n5700), .ZN(n9625) );
  NOR3_X1 U7431 ( .A1(n8244), .A2(n9625), .A3(n9830), .ZN(n5703) );
  OAI21_X1 U7432 ( .B1(n9625), .B2(n8242), .A(n8244), .ZN(n5705) );
  OAI211_X1 U7433 ( .C1(n5708), .C2(n5791), .A(n5706), .B(n5705), .ZN(n5712)
         );
  OR4_X1 U7434 ( .A1(n8244), .A2(n9625), .A3(n8242), .A4(n6468), .ZN(n5711) );
  INV_X1 U7435 ( .A(n8242), .ZN(n9352) );
  NAND3_X1 U7436 ( .A1(n9625), .A2(n6468), .A3(n9352), .ZN(n5707) );
  OAI21_X1 U7437 ( .B1(n4735), .B2(n5708), .A(n5707), .ZN(n5709) );
  AOI21_X1 U7438 ( .B1(n8244), .B2(n5709), .A(n5851), .ZN(n5710) );
  OAI21_X1 U7439 ( .B1(n5877), .B2(n4452), .A(n6464), .ZN(n5804) );
  INV_X1 U7440 ( .A(n5716), .ZN(n5879) );
  NAND2_X1 U7441 ( .A1(n5794), .A2(n5879), .ZN(n5850) );
  NAND2_X1 U7442 ( .A1(n5761), .A2(n6476), .ZN(n9657) );
  INV_X1 U7443 ( .A(n9657), .ZN(n9648) );
  NAND2_X1 U7444 ( .A1(n5720), .A2(n5782), .ZN(n7741) );
  NAND2_X1 U7445 ( .A1(n5778), .A2(n5826), .ZN(n7418) );
  NAND2_X1 U7446 ( .A1(n5723), .A2(n7435), .ZN(n7342) );
  NAND3_X1 U7447 ( .A1(n6435), .A2(n5724), .A3(n7242), .ZN(n5823) );
  INV_X1 U7448 ( .A(n6434), .ZN(n5772) );
  AND2_X1 U7449 ( .A1(n9377), .A2(n6991), .ZN(n5807) );
  OR2_X1 U7450 ( .A1(n5807), .A2(n6993), .ZN(n6979) );
  NOR3_X1 U7451 ( .A1(n6979), .A2(n6419), .A3(n6464), .ZN(n5728) );
  INV_X1 U7452 ( .A(n7027), .ZN(n5767) );
  NAND2_X1 U7453 ( .A1(n5770), .A2(n5726), .ZN(n7130) );
  INV_X1 U7454 ( .A(n7130), .ZN(n7128) );
  NAND4_X1 U7455 ( .A1(n5728), .A2(n5767), .A3(n7128), .A4(n6994), .ZN(n5729)
         );
  INV_X1 U7456 ( .A(n10015), .ZN(n10020) );
  NAND4_X1 U7457 ( .A1(n6438), .A2(n4567), .A3(n7438), .A4(n5731), .ZN(n5732)
         );
  NOR4_X1 U7458 ( .A1(n5784), .A2(n7572), .A3(n7741), .A4(n5732), .ZN(n5733)
         );
  NAND2_X1 U7459 ( .A1(n5734), .A2(n5789), .ZN(n9784) );
  NAND4_X1 U7460 ( .A1(n9713), .A2(n9727), .A3(n5736), .A4(n9748), .ZN(n5737)
         );
  NOR4_X1 U7461 ( .A1(n5738), .A2(n9665), .A3(n9691), .A4(n5737), .ZN(n5739)
         );
  NAND2_X1 U7462 ( .A1(n5745), .A2(n5744), .ZN(n5746) );
  NOR4_X1 U7463 ( .A1(n5799), .A2(n4469), .A3(n9788), .A4(n6675), .ZN(n5803)
         );
  NAND2_X1 U7464 ( .A1(n4471), .A2(n6464), .ZN(n6794) );
  INV_X1 U7465 ( .A(n6794), .ZN(n6677) );
  INV_X1 U7466 ( .A(n5761), .ZN(n5766) );
  INV_X1 U7467 ( .A(n5749), .ZN(n5765) );
  NAND3_X1 U7468 ( .A1(n5756), .A2(n9690), .A3(n5750), .ZN(n5751) );
  AND2_X1 U7469 ( .A1(n5751), .A2(n6471), .ZN(n5752) );
  AND2_X1 U7470 ( .A1(n5752), .A2(n6474), .ZN(n5762) );
  NAND2_X1 U7471 ( .A1(n5754), .A2(n5753), .ZN(n9728) );
  NAND3_X1 U7472 ( .A1(n5756), .A2(n5755), .A3(n9728), .ZN(n5757) );
  NOR3_X1 U7473 ( .A1(n5766), .A2(n5765), .A3(n5758), .ZN(n5759) );
  INV_X1 U7474 ( .A(n6469), .ZN(n5764) );
  INV_X1 U7475 ( .A(n5762), .ZN(n5763) );
  NOR4_X1 U7476 ( .A1(n5766), .A2(n5765), .A3(n5764), .A4(n5763), .ZN(n5845)
         );
  NAND2_X1 U7477 ( .A1(n7131), .A2(n7129), .ZN(n5769) );
  NAND2_X1 U7478 ( .A1(n7133), .A2(n5770), .ZN(n10014) );
  AND2_X1 U7479 ( .A1(n5775), .A2(n6434), .ZN(n5821) );
  INV_X1 U7480 ( .A(n7342), .ZN(n7344) );
  NAND2_X1 U7481 ( .A1(n7419), .A2(n7417), .ZN(n5777) );
  NAND2_X1 U7482 ( .A1(n5777), .A2(n4567), .ZN(n7421) );
  NOR2_X1 U7483 ( .A1(n7741), .A2(n5780), .ZN(n5781) );
  INV_X1 U7484 ( .A(n9801), .ZN(n5783) );
  NOR2_X1 U7485 ( .A1(n5784), .A2(n5783), .ZN(n5785) );
  NAND2_X1 U7486 ( .A1(n9776), .A2(n5839), .ZN(n6470) );
  NAND2_X1 U7487 ( .A1(n5845), .A2(n6470), .ZN(n5792) );
  NAND2_X1 U7488 ( .A1(n5791), .A2(n5790), .ZN(n5848) );
  AOI21_X1 U7489 ( .B1(n5842), .B2(n5792), .A(n5848), .ZN(n5797) );
  NAND2_X1 U7490 ( .A1(n4356), .A2(n5793), .ZN(n5846) );
  INV_X1 U7491 ( .A(n5794), .ZN(n5795) );
  OAI21_X1 U7492 ( .B1(n5795), .B2(n8242), .A(n4735), .ZN(n5796) );
  OAI21_X1 U7493 ( .B1(n5797), .B2(n5846), .A(n5796), .ZN(n5798) );
  OAI211_X1 U7494 ( .C1(n9833), .C2(n4735), .A(n5798), .B(n5881), .ZN(n5800)
         );
  AOI21_X1 U7495 ( .B1(n5804), .B2(n5803), .A(n5802), .ZN(n5886) );
  AND2_X2 U7496 ( .A1(n6783), .A2(n7223), .ZN(n6802) );
  INV_X1 U7497 ( .A(n5805), .ZN(n5834) );
  INV_X1 U7498 ( .A(n5806), .ZN(n5829) );
  INV_X1 U7499 ( .A(n5807), .ZN(n5809) );
  INV_X2 U7500 ( .A(n10043), .ZN(n6992) );
  NAND2_X1 U7501 ( .A1(n6849), .A2(n6992), .ZN(n5808) );
  NAND3_X1 U7502 ( .A1(n5809), .A2(n6464), .A3(n5808), .ZN(n5811) );
  NAND2_X1 U7503 ( .A1(n5811), .A2(n5810), .ZN(n5813) );
  NAND2_X1 U7504 ( .A1(n5813), .A2(n5812), .ZN(n5814) );
  NAND3_X1 U7505 ( .A1(n5297), .A2(n7129), .A3(n5814), .ZN(n5817) );
  INV_X1 U7506 ( .A(n5815), .ZN(n5816) );
  NAND2_X1 U7507 ( .A1(n5817), .A2(n5816), .ZN(n5818) );
  NAND2_X1 U7508 ( .A1(n5818), .A2(n4385), .ZN(n5820) );
  AOI21_X1 U7509 ( .B1(n5820), .B2(n5819), .A(n4662), .ZN(n5824) );
  OAI211_X1 U7510 ( .C1(n5824), .C2(n5823), .A(n5822), .B(n5821), .ZN(n5825)
         );
  INV_X1 U7511 ( .A(n5825), .ZN(n5828) );
  OAI211_X1 U7512 ( .C1(n5829), .C2(n5828), .A(n5827), .B(n5826), .ZN(n5831)
         );
  AOI21_X1 U7513 ( .B1(n5832), .B2(n5831), .A(n5830), .ZN(n5833) );
  AOI211_X1 U7514 ( .C1(n9801), .C2(n5835), .A(n5834), .B(n5833), .ZN(n5838)
         );
  INV_X1 U7515 ( .A(n5836), .ZN(n5837) );
  NOR2_X1 U7516 ( .A1(n5838), .A2(n5837), .ZN(n5841) );
  OAI21_X1 U7517 ( .B1(n5841), .B2(n5840), .A(n5839), .ZN(n5844) );
  INV_X1 U7518 ( .A(n5842), .ZN(n5843) );
  AOI21_X1 U7519 ( .B1(n5845), .B2(n5844), .A(n5843), .ZN(n5849) );
  INV_X1 U7520 ( .A(n5846), .ZN(n5847) );
  OAI21_X1 U7521 ( .B1(n5849), .B2(n5848), .A(n5847), .ZN(n5853) );
  INV_X1 U7522 ( .A(n5850), .ZN(n5852) );
  OAI21_X1 U7523 ( .B1(n6796), .B2(n9788), .A(n5855), .ZN(n5854) );
  INV_X1 U7524 ( .A(n6675), .ZN(n7316) );
  OAI211_X1 U7525 ( .C1(n6802), .C2(n5855), .A(n5854), .B(n7316), .ZN(n5876)
         );
  NAND3_X1 U7526 ( .A1(n5858), .A2(n5857), .A3(n5856), .ZN(n5860) );
  NAND2_X1 U7527 ( .A1(n5869), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5863) );
  MUX2_X1 U7528 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5863), .S(
        P1_IR_REG_25__SCAN_IN), .Z(n5865) );
  NAND2_X1 U7529 ( .A1(n5866), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5867) );
  MUX2_X1 U7530 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5867), .S(
        P1_IR_REG_24__SCAN_IN), .Z(n5868) );
  NAND2_X1 U7531 ( .A1(n5864), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5870) );
  INV_X1 U7532 ( .A(n6787), .ZN(n5873) );
  NAND2_X1 U7533 ( .A1(n5872), .A2(n7223), .ZN(n6785) );
  INV_X1 U7534 ( .A(n6785), .ZN(n6781) );
  NOR2_X1 U7535 ( .A1(n8232), .A2(n4281), .ZN(n9393) );
  NAND4_X1 U7536 ( .A1(n9951), .A2(n5873), .A3(n6781), .A4(n9393), .ZN(n5874)
         );
  OAI211_X1 U7537 ( .C1(n4471), .C2(n6675), .A(n5874), .B(P1_B_REG_SCAN_IN), 
        .ZN(n5875) );
  INV_X1 U7538 ( .A(n5877), .ZN(n5878) );
  OAI21_X1 U7539 ( .B1(n6468), .B2(n5879), .A(n5878), .ZN(n5884) );
  NAND2_X1 U7540 ( .A1(n6464), .A2(n6796), .ZN(n6479) );
  NOR3_X1 U7541 ( .A1(n6675), .A2(n4471), .A3(n6479), .ZN(n5880) );
  INV_X1 U7542 ( .A(n5882), .ZN(n5883) );
  NAND2_X1 U7543 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5887) );
  XNOR2_X2 U7544 ( .A(n5887), .B(P2_IR_REG_1__SCAN_IN), .ZN(n6767) );
  NOR2_X1 U7545 ( .A1(P2_IR_REG_26__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), .ZN(
        n5898) );
  AND2_X1 U7546 ( .A1(n5902), .A2(n5898), .ZN(n5899) );
  INV_X1 U7547 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n5900) );
  XNOR2_X2 U7548 ( .A(n5901), .B(n5928), .ZN(n6367) );
  INV_X1 U7549 ( .A(n5902), .ZN(n6337) );
  NAND2_X1 U7550 ( .A1(n6340), .A2(P2_IR_REG_27__SCAN_IN), .ZN(n5903) );
  NOR2_X1 U7551 ( .A1(n6337), .A2(n5903), .ZN(n5909) );
  XNOR2_X1 U7552 ( .A(n5904), .B(P2_IR_REG_31__SCAN_IN), .ZN(n5908) );
  INV_X1 U7553 ( .A(n5929), .ZN(n5907) );
  INV_X1 U7554 ( .A(n5913), .ZN(n6005) );
  NAND2_X1 U7555 ( .A1(n6156), .A2(n5914), .ZN(n6167) );
  INV_X1 U7556 ( .A(n5917), .ZN(n5918) );
  NOR2_X1 U7557 ( .A1(n6005), .A2(n5918), .ZN(n5919) );
  NAND2_X1 U7558 ( .A1(n5919), .A2(n4284), .ZN(n5923) );
  NAND2_X1 U7559 ( .A1(n6194), .A2(n5922), .ZN(n5927) );
  NAND2_X1 U7560 ( .A1(n5923), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5924) );
  MUX2_X1 U7561 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5924), .S(
        P2_IR_REG_20__SCAN_IN), .Z(n5926) );
  AND2_X2 U7562 ( .A1(n4908), .A2(n5931), .ZN(n5933) );
  NAND2_X1 U7563 ( .A1(n5969), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5938) );
  INV_X1 U7564 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n5932) );
  NAND2_X1 U7565 ( .A1(n6024), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n5936) );
  NAND2_X1 U7566 ( .A1(n4285), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n5935) );
  NAND2_X1 U7567 ( .A1(n6516), .A2(n5939), .ZN(n5950) );
  NAND2_X1 U7568 ( .A1(n6024), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n5944) );
  NAND2_X1 U7569 ( .A1(n5969), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5943) );
  INV_X1 U7570 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n6762) );
  INV_X1 U7571 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n5940) );
  OR2_X1 U7572 ( .A1(n5974), .A2(n5940), .ZN(n5941) );
  NAND2_X1 U7573 ( .A1(n8003), .A2(SI_0_), .ZN(n5946) );
  INV_X1 U7574 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5945) );
  NAND2_X1 U7575 ( .A1(n5946), .A2(n5945), .ZN(n5948) );
  AND2_X1 U7576 ( .A1(n5947), .A2(n5948), .ZN(n9063) );
  MUX2_X1 U7577 ( .A(P2_IR_REG_0__SCAN_IN), .B(n9063), .S(n6614), .Z(n6742) );
  NAND2_X1 U7578 ( .A1(n6741), .A2(n6742), .ZN(n8022) );
  INV_X1 U7579 ( .A(n6742), .ZN(n6942) );
  NAND2_X1 U7580 ( .A1(n6942), .A2(n4279), .ZN(n5949) );
  NAND2_X1 U7581 ( .A1(n8022), .A2(n5949), .ZN(n6862) );
  NAND2_X1 U7582 ( .A1(n6764), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5951) );
  INV_X1 U7583 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n8985) );
  NAND2_X2 U7584 ( .A1(n5952), .A2(n5981), .ZN(n6959) );
  OR2_X1 U7585 ( .A1(n5958), .A2(n6667), .ZN(n5954) );
  OR2_X1 U7586 ( .A1(n4268), .A2(n6668), .ZN(n5953) );
  XNOR2_X1 U7587 ( .A(n5955), .B(n4882), .ZN(n7097) );
  NAND2_X1 U7588 ( .A1(n6519), .A2(n5955), .ZN(n5956) );
  INV_X1 U7589 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n5957) );
  OR2_X1 U7590 ( .A1(n9058), .A2(n5980), .ZN(n5961) );
  OAI211_X1 U7591 ( .C1(n6614), .C2(n4270), .A(n5961), .B(n5960), .ZN(n10195)
         );
  XNOR2_X1 U7592 ( .A(n10195), .B(n4279), .ZN(n5967) );
  NAND2_X1 U7593 ( .A1(n6024), .A2(n5971), .ZN(n5965) );
  NAND2_X1 U7594 ( .A1(n4285), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n5964) );
  NAND2_X1 U7595 ( .A1(n5995), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5963) );
  NAND2_X1 U7596 ( .A1(n5969), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5962) );
  XNOR2_X1 U7597 ( .A(n5967), .B(n10176), .ZN(n7006) );
  NAND2_X1 U7598 ( .A1(n5967), .A2(n10176), .ZN(n5968) );
  NAND2_X1 U7599 ( .A1(n7003), .A2(n5968), .ZN(n7160) );
  INV_X1 U7600 ( .A(n7160), .ZN(n5989) );
  NAND2_X1 U7601 ( .A1(n8011), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5979) );
  INV_X1 U7602 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n5970) );
  NAND2_X1 U7603 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n5972) );
  NAND2_X1 U7604 ( .A1(n5997), .A2(n5972), .ZN(n10184) );
  NAND2_X1 U7605 ( .A1(n6323), .A2(n10184), .ZN(n5978) );
  INV_X1 U7606 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n6951) );
  OR2_X1 U7607 ( .A1(n4286), .A2(n6951), .ZN(n5977) );
  INV_X1 U7608 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n5975) );
  OR2_X1 U7609 ( .A1(n4271), .A2(n5975), .ZN(n5976) );
  INV_X1 U7610 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6672) );
  NAND2_X1 U7611 ( .A1(n6665), .A2(n8007), .ZN(n5984) );
  NAND2_X1 U7612 ( .A1(n5991), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5982) );
  NAND2_X1 U7613 ( .A1(n8005), .A2(n6964), .ZN(n5983) );
  OAI211_X1 U7614 ( .C1(n8008), .C2(n6672), .A(n5984), .B(n5983), .ZN(n10200)
         );
  XNOR2_X1 U7615 ( .A(n10200), .B(n6283), .ZN(n5985) );
  NAND2_X1 U7616 ( .A1(n7229), .A2(n5985), .ZN(n5990) );
  INV_X1 U7617 ( .A(n5985), .ZN(n5986) );
  INV_X1 U7618 ( .A(n7229), .ZN(n8402) );
  NAND2_X1 U7619 ( .A1(n5986), .A2(n8402), .ZN(n5987) );
  NAND2_X1 U7620 ( .A1(n5990), .A2(n5987), .ZN(n7159) );
  INV_X1 U7621 ( .A(n7159), .ZN(n5988) );
  NAND2_X1 U7622 ( .A1(n6661), .A2(n8007), .ZN(n5994) );
  OAI21_X1 U7623 ( .B1(n5991), .B2(P2_IR_REG_4__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5992) );
  XNOR2_X1 U7624 ( .A(n5992), .B(P2_IR_REG_5__SCAN_IN), .ZN(n7069) );
  AOI22_X1 U7625 ( .A1(n6195), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n8005), .B2(
        n7069), .ZN(n5993) );
  NAND2_X1 U7626 ( .A1(n5994), .A2(n5993), .ZN(n10205) );
  XNOR2_X1 U7627 ( .A(n10205), .B(n6283), .ZN(n6003) );
  NAND2_X1 U7628 ( .A1(n8012), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n6002) );
  NAND2_X1 U7629 ( .A1(n5995), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n6001) );
  NAND2_X1 U7630 ( .A1(n5997), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5998) );
  NAND2_X1 U7631 ( .A1(n6009), .A2(n5998), .ZN(n7235) );
  NAND2_X1 U7632 ( .A1(n6323), .A2(n7235), .ZN(n6000) );
  NAND2_X1 U7633 ( .A1(n8011), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n5999) );
  NAND4_X1 U7634 ( .A1(n6002), .A2(n6001), .A3(n6000), .A4(n5999), .ZN(n10174)
         );
  XNOR2_X1 U7635 ( .A(n6003), .B(n10174), .ZN(n7147) );
  INV_X1 U7636 ( .A(n10174), .ZN(n7201) );
  NAND2_X1 U7637 ( .A1(n6003), .A2(n7201), .ZN(n6004) );
  NAND2_X1 U7638 ( .A1(n6663), .A2(n8007), .ZN(n6008) );
  NAND2_X1 U7639 ( .A1(n6005), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6006) );
  AOI22_X1 U7640 ( .A1(n6195), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n8005), .B2(
        n7185), .ZN(n6007) );
  XNOR2_X1 U7641 ( .A(n10215), .B(n6283), .ZN(n6015) );
  NAND2_X1 U7642 ( .A1(n8011), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6014) );
  NAND2_X1 U7643 ( .A1(n8012), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n6013) );
  NAND2_X1 U7644 ( .A1(n6009), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n6010) );
  NAND2_X1 U7645 ( .A1(n6027), .A2(n6010), .ZN(n7260) );
  NAND2_X1 U7646 ( .A1(n6024), .A2(n7260), .ZN(n6012) );
  NAND2_X1 U7647 ( .A1(n5995), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n6011) );
  XNOR2_X1 U7648 ( .A(n6015), .B(n8401), .ZN(n7197) );
  INV_X1 U7649 ( .A(n6015), .ZN(n6016) );
  NAND2_X1 U7650 ( .A1(n6016), .A2(n8401), .ZN(n6017) );
  NAND2_X1 U7651 ( .A1(n6691), .A2(n8007), .ZN(n6023) );
  INV_X1 U7652 ( .A(n6018), .ZN(n6020) );
  NAND2_X1 U7653 ( .A1(n6020), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6019) );
  MUX2_X1 U7654 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6019), .S(
        P2_IR_REG_7__SCAN_IN), .Z(n6021) );
  AOI22_X1 U7655 ( .A1(n6195), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n8005), .B2(
        n7271), .ZN(n6022) );
  NAND2_X2 U7656 ( .A1(n6023), .A2(n6022), .ZN(n7485) );
  XNOR2_X1 U7657 ( .A(n7485), .B(n6283), .ZN(n6034) );
  NAND2_X1 U7658 ( .A1(n8011), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6033) );
  INV_X1 U7659 ( .A(n6027), .ZN(n6026) );
  NAND2_X1 U7660 ( .A1(n6027), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n6028) );
  NAND2_X1 U7661 ( .A1(n6042), .A2(n6028), .ZN(n7473) );
  NAND2_X1 U7662 ( .A1(n6323), .A2(n7473), .ZN(n6032) );
  INV_X1 U7663 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n7472) );
  OR2_X1 U7664 ( .A1(n5973), .A2(n7472), .ZN(n6031) );
  INV_X1 U7665 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n6029) );
  OR2_X1 U7666 ( .A1(n4271), .A2(n6029), .ZN(n6030) );
  NAND2_X1 U7667 ( .A1(n6034), .A2(n6531), .ZN(n7358) );
  INV_X1 U7668 ( .A(n6034), .ZN(n6035) );
  NAND2_X1 U7669 ( .A1(n6035), .A2(n8400), .ZN(n6036) );
  NAND2_X1 U7670 ( .A1(n7358), .A2(n6036), .ZN(n7285) );
  NAND2_X1 U7671 ( .A1(n6038), .A2(n8007), .ZN(n6041) );
  NAND2_X1 U7672 ( .A1(n6051), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6039) );
  XNOR2_X1 U7673 ( .A(n6039), .B(P2_IR_REG_8__SCAN_IN), .ZN(n7305) );
  AOI22_X1 U7674 ( .A1(n6195), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n8005), .B2(
        n7305), .ZN(n6040) );
  NAND2_X1 U7675 ( .A1(n6041), .A2(n6040), .ZN(n7465) );
  XNOR2_X1 U7676 ( .A(n7465), .B(n6283), .ZN(n6049) );
  NAND2_X1 U7677 ( .A1(n8011), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n6047) );
  NAND2_X1 U7678 ( .A1(n8012), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n6046) );
  NAND2_X1 U7679 ( .A1(n6042), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n6043) );
  NAND2_X1 U7680 ( .A1(n6060), .A2(n6043), .ZN(n7458) );
  NAND2_X1 U7681 ( .A1(n6323), .A2(n7458), .ZN(n6045) );
  NAND2_X1 U7682 ( .A1(n5995), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n6044) );
  NAND4_X1 U7683 ( .A1(n6047), .A2(n6046), .A3(n6045), .A4(n6044), .ZN(n8399)
         );
  XNOR2_X1 U7684 ( .A(n6049), .B(n8399), .ZN(n7359) );
  NAND2_X1 U7685 ( .A1(n6049), .A2(n8322), .ZN(n6050) );
  NAND2_X1 U7686 ( .A1(n6708), .A2(n8007), .ZN(n6058) );
  INV_X1 U7687 ( .A(n6051), .ZN(n6053) );
  NAND2_X1 U7688 ( .A1(n6053), .A2(n6052), .ZN(n6066) );
  NAND2_X1 U7689 ( .A1(n6066), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6055) );
  NAND2_X1 U7690 ( .A1(n6055), .A2(n6054), .ZN(n6081) );
  OR2_X1 U7691 ( .A1(n6055), .A2(n6054), .ZN(n6056) );
  AOI22_X1 U7692 ( .A1(n6195), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n8005), .B2(
        n7394), .ZN(n6057) );
  NAND2_X1 U7693 ( .A1(n6058), .A2(n6057), .ZN(n8324) );
  XNOR2_X1 U7694 ( .A(n8324), .B(n6283), .ZN(n6085) );
  NAND2_X1 U7695 ( .A1(n8011), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n6065) );
  NAND2_X1 U7696 ( .A1(n8012), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n6064) );
  NAND2_X1 U7697 ( .A1(n6060), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n6061) );
  NAND2_X1 U7698 ( .A1(n6074), .A2(n6061), .ZN(n8325) );
  NAND2_X1 U7699 ( .A1(n6323), .A2(n8325), .ZN(n6063) );
  NAND2_X1 U7700 ( .A1(n5995), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n6062) );
  NAND4_X1 U7701 ( .A1(n6065), .A2(n6064), .A3(n6063), .A4(n6062), .ZN(n8398)
         );
  XNOR2_X1 U7702 ( .A(n6085), .B(n8398), .ZN(n8319) );
  NAND2_X1 U7703 ( .A1(n6094), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6067) );
  XNOR2_X1 U7704 ( .A(n6067), .B(P2_IR_REG_11__SCAN_IN), .ZN(n7700) );
  AOI22_X1 U7705 ( .A1(n6195), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n8005), .B2(
        n7700), .ZN(n6068) );
  NAND2_X1 U7706 ( .A1(n6076), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6069) );
  NAND2_X1 U7707 ( .A1(n6100), .A2(n6069), .ZN(n7784) );
  NAND2_X1 U7708 ( .A1(n6323), .A2(n7784), .ZN(n6073) );
  NAND2_X1 U7709 ( .A1(n8011), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n6072) );
  INV_X1 U7710 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n7696) );
  OR2_X1 U7711 ( .A1(n5973), .A2(n7696), .ZN(n6071) );
  INV_X1 U7712 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n7595) );
  OR2_X1 U7713 ( .A1(n4271), .A2(n7595), .ZN(n6070) );
  NAND2_X1 U7714 ( .A1(n6536), .A2(n7565), .ZN(n8081) );
  XNOR2_X1 U7715 ( .A(n8187), .B(n4279), .ZN(n7779) );
  NAND2_X1 U7716 ( .A1(n8012), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n6080) );
  NAND2_X1 U7717 ( .A1(n8011), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n6079) );
  NAND2_X1 U7718 ( .A1(n6074), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n6075) );
  NAND2_X1 U7719 ( .A1(n6076), .A2(n6075), .ZN(n7769) );
  NAND2_X1 U7720 ( .A1(n6323), .A2(n7769), .ZN(n6078) );
  NAND2_X1 U7721 ( .A1(n5995), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n6077) );
  NAND4_X1 U7722 ( .A1(n6080), .A2(n6079), .A3(n6078), .A4(n6077), .ZN(n8397)
         );
  NAND2_X1 U7723 ( .A1(n6712), .A2(n8007), .ZN(n6084) );
  NAND2_X1 U7724 ( .A1(n6081), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6082) );
  XNOR2_X1 U7725 ( .A(n6082), .B(P2_IR_REG_10__SCAN_IN), .ZN(n7540) );
  AOI22_X1 U7726 ( .A1(n6195), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n8005), .B2(
        n7540), .ZN(n6083) );
  XNOR2_X1 U7727 ( .A(n7770), .B(n4279), .ZN(n7776) );
  INV_X1 U7728 ( .A(n6085), .ZN(n6086) );
  AND2_X1 U7729 ( .A1(n6086), .A2(n8398), .ZN(n7760) );
  AOI21_X1 U7730 ( .B1(n8397), .B2(n7776), .A(n7760), .ZN(n6087) );
  AND2_X1 U7731 ( .A1(n7779), .A2(n6087), .ZN(n6093) );
  NAND3_X1 U7732 ( .A1(n7770), .A2(n7782), .A3(n6283), .ZN(n6088) );
  OAI21_X1 U7733 ( .B1(n6283), .B2(n8396), .A(n6088), .ZN(n6091) );
  NAND2_X1 U7734 ( .A1(n7782), .A2(n4279), .ZN(n6089) );
  OAI22_X1 U7735 ( .A1(n7770), .A2(n6089), .B1(n8396), .B2(n4279), .ZN(n6090)
         );
  MUX2_X1 U7736 ( .A(n6091), .B(n6090), .S(n8187), .Z(n6092) );
  NAND2_X1 U7737 ( .A1(n6858), .A2(n8007), .ZN(n6097) );
  NAND2_X1 U7738 ( .A1(n6109), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6095) );
  XNOR2_X1 U7739 ( .A(n6095), .B(P2_IR_REG_12__SCAN_IN), .ZN(n8412) );
  AOI22_X1 U7740 ( .A1(n6195), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n8005), .B2(
        n8412), .ZN(n6096) );
  XNOR2_X1 U7741 ( .A(n7636), .B(n6283), .ZN(n6106) );
  NAND2_X1 U7742 ( .A1(n8011), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n6105) );
  NAND2_X1 U7743 ( .A1(n6100), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n6101) );
  NAND2_X1 U7744 ( .A1(n6114), .A2(n6101), .ZN(n7632) );
  NAND2_X1 U7745 ( .A1(n6323), .A2(n7632), .ZN(n6104) );
  INV_X1 U7746 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n8407) );
  OR2_X1 U7747 ( .A1(n4286), .A2(n8407), .ZN(n6103) );
  INV_X1 U7748 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n7618) );
  OR2_X1 U7749 ( .A1(n4271), .A2(n7618), .ZN(n6102) );
  NAND2_X1 U7750 ( .A1(n6106), .A2(n7626), .ZN(n7558) );
  NAND2_X1 U7751 ( .A1(n7560), .A2(n7558), .ZN(n6108) );
  INV_X1 U7752 ( .A(n6106), .ZN(n6107) );
  NAND2_X1 U7753 ( .A1(n6107), .A2(n8395), .ZN(n7559) );
  NAND2_X1 U7754 ( .A1(n6108), .A2(n7559), .ZN(n7621) );
  NAND2_X1 U7755 ( .A1(n6919), .A2(n8007), .ZN(n6111) );
  OAI21_X1 U7756 ( .B1(n6109), .B2(P2_IR_REG_12__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n6125) );
  XNOR2_X1 U7757 ( .A(n6125), .B(P2_IR_REG_13__SCAN_IN), .ZN(n8438) );
  AOI22_X1 U7758 ( .A1(n6195), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n8438), .B2(
        n8005), .ZN(n6110) );
  XNOR2_X1 U7759 ( .A(n8093), .B(n6283), .ZN(n7623) );
  NAND2_X1 U7760 ( .A1(n8011), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n6119) );
  INV_X1 U7761 ( .A(n6114), .ZN(n6113) );
  NAND2_X1 U7762 ( .A1(n6114), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n6115) );
  NAND2_X1 U7763 ( .A1(n6132), .A2(n6115), .ZN(n7628) );
  NAND2_X1 U7764 ( .A1(n6323), .A2(n7628), .ZN(n6118) );
  INV_X1 U7765 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n8410) );
  OR2_X1 U7766 ( .A1(n5973), .A2(n8410), .ZN(n6117) );
  INV_X1 U7767 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n7687) );
  OR2_X1 U7768 ( .A1(n4271), .A2(n7687), .ZN(n6116) );
  NAND2_X1 U7769 ( .A1(n7623), .A2(n7793), .ZN(n6120) );
  NAND2_X1 U7770 ( .A1(n7621), .A2(n6120), .ZN(n6123) );
  INV_X1 U7771 ( .A(n7623), .ZN(n6121) );
  NAND2_X1 U7772 ( .A1(n6121), .A2(n8394), .ZN(n6122) );
  NAND2_X1 U7773 ( .A1(n7011), .A2(n8007), .ZN(n6131) );
  NAND2_X1 U7774 ( .A1(n6125), .A2(n6124), .ZN(n6126) );
  NAND2_X1 U7775 ( .A1(n6126), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6128) );
  NAND2_X1 U7776 ( .A1(n6128), .A2(n6127), .ZN(n6143) );
  OR2_X1 U7777 ( .A1(n6128), .A2(n6127), .ZN(n6129) );
  AOI22_X1 U7778 ( .A1(n8467), .A2(n8005), .B1(n6195), .B2(
        P1_DATAO_REG_14__SCAN_IN), .ZN(n6130) );
  XNOR2_X1 U7779 ( .A(n7993), .B(n4279), .ZN(n6140) );
  NAND2_X1 U7780 ( .A1(n8011), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n6137) );
  NAND2_X1 U7781 ( .A1(n8012), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n6136) );
  NAND2_X1 U7782 ( .A1(n6132), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n6133) );
  NAND2_X1 U7783 ( .A1(n6149), .A2(n6133), .ZN(n7997) );
  NAND2_X1 U7784 ( .A1(n6323), .A2(n7997), .ZN(n6135) );
  NAND2_X1 U7785 ( .A1(n5995), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n6134) );
  NAND4_X1 U7786 ( .A1(n6137), .A2(n6136), .A3(n6135), .A4(n6134), .ZN(n8393)
         );
  XNOR2_X1 U7787 ( .A(n6140), .B(n8393), .ZN(n7791) );
  INV_X1 U7788 ( .A(n7791), .ZN(n6138) );
  INV_X1 U7789 ( .A(n6140), .ZN(n6141) );
  INV_X1 U7790 ( .A(n8393), .ZN(n8383) );
  NAND2_X1 U7791 ( .A1(n6141), .A2(n8383), .ZN(n6142) );
  NAND2_X1 U7792 ( .A1(n7048), .A2(n8007), .ZN(n6146) );
  NAND2_X1 U7793 ( .A1(n6143), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6144) );
  AOI22_X1 U7794 ( .A1(n8479), .A2(n8005), .B1(n6195), .B2(
        P1_DATAO_REG_15__SCAN_IN), .ZN(n6145) );
  XNOR2_X1 U7795 ( .A(n8814), .B(n4279), .ZN(n6154) );
  INV_X1 U7796 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n6153) );
  NAND2_X1 U7797 ( .A1(n8012), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n6148) );
  NAND2_X1 U7798 ( .A1(n8011), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n6147) );
  AND2_X1 U7799 ( .A1(n6148), .A2(n6147), .ZN(n6152) );
  NAND2_X1 U7800 ( .A1(n6149), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n6150) );
  NAND2_X1 U7801 ( .A1(n6162), .A2(n6150), .ZN(n8386) );
  NAND2_X1 U7802 ( .A1(n8386), .A2(n6323), .ZN(n6151) );
  OAI211_X1 U7803 ( .C1(n4271), .C2(n6153), .A(n6152), .B(n6151), .ZN(n8392)
         );
  XNOR2_X1 U7804 ( .A(n6154), .B(n8392), .ZN(n8376) );
  NAND2_X1 U7805 ( .A1(n6154), .A2(n8392), .ZN(n6155) );
  NAND2_X1 U7806 ( .A1(n8378), .A2(n6155), .ZN(n8299) );
  NAND2_X1 U7807 ( .A1(n7125), .A2(n8007), .ZN(n6161) );
  INV_X1 U7808 ( .A(n6156), .ZN(n6157) );
  NAND2_X1 U7809 ( .A1(n6157), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6158) );
  MUX2_X1 U7810 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6158), .S(
        P2_IR_REG_16__SCAN_IN), .Z(n6159) );
  NAND2_X1 U7811 ( .A1(n6159), .A2(n6167), .ZN(n8514) );
  INV_X1 U7812 ( .A(n8514), .ZN(n8494) );
  AOI22_X1 U7813 ( .A1(n6195), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n8005), .B2(
        n8494), .ZN(n6160) );
  NAND2_X1 U7814 ( .A1(n6161), .A2(n6160), .ZN(n6553) );
  XNOR2_X1 U7815 ( .A(n6553), .B(n4279), .ZN(n8301) );
  INV_X1 U7816 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n8892) );
  NAND2_X1 U7817 ( .A1(n6162), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n6163) );
  NAND2_X1 U7818 ( .A1(n6173), .A2(n6163), .ZN(n8744) );
  NAND2_X1 U7819 ( .A1(n8744), .A2(n6323), .ZN(n6165) );
  AOI22_X1 U7820 ( .A1(n8011), .A2(P2_REG1_REG_16__SCAN_IN), .B1(n8012), .B2(
        P2_REG2_REG_16__SCAN_IN), .ZN(n6164) );
  AND2_X1 U7821 ( .A1(n8301), .A2(n8724), .ZN(n6166) );
  NAND2_X1 U7822 ( .A1(n7155), .A2(n8007), .ZN(n6170) );
  NAND2_X1 U7823 ( .A1(n6167), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6168) );
  XNOR2_X1 U7824 ( .A(n6168), .B(P2_IR_REG_17__SCAN_IN), .ZN(n8533) );
  AOI22_X1 U7825 ( .A1(n6195), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n8005), .B2(
        n8533), .ZN(n6169) );
  NAND2_X1 U7826 ( .A1(n6173), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n6174) );
  NAND2_X1 U7827 ( .A1(n6185), .A2(n6174), .ZN(n8729) );
  NAND2_X1 U7828 ( .A1(n8729), .A2(n6323), .ZN(n6177) );
  AOI22_X1 U7829 ( .A1(n8011), .A2(P2_REG1_REG_17__SCAN_IN), .B1(n8012), .B2(
        P2_REG2_REG_17__SCAN_IN), .ZN(n6176) );
  NAND2_X1 U7830 ( .A1(n5995), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n6175) );
  INV_X1 U7831 ( .A(n8309), .ZN(n6178) );
  INV_X1 U7832 ( .A(n8740), .ZN(n8357) );
  NAND2_X1 U7833 ( .A1(n7192), .A2(n8007), .ZN(n6184) );
  INV_X1 U7834 ( .A(n6179), .ZN(n6180) );
  NAND2_X1 U7835 ( .A1(n6180), .A2(P2_IR_REG_18__SCAN_IN), .ZN(n6182) );
  AOI22_X1 U7836 ( .A1(n6195), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n8005), .B2(
        n8562), .ZN(n6183) );
  XNOR2_X1 U7837 ( .A(n8803), .B(n6283), .ZN(n6190) );
  NAND2_X1 U7838 ( .A1(n6185), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n6186) );
  NAND2_X1 U7839 ( .A1(n6198), .A2(n6186), .ZN(n8712) );
  NAND2_X1 U7840 ( .A1(n8712), .A2(n6323), .ZN(n6189) );
  AOI22_X1 U7841 ( .A1(n8011), .A2(P2_REG1_REG_18__SCAN_IN), .B1(n8012), .B2(
        P2_REG2_REG_18__SCAN_IN), .ZN(n6188) );
  NAND2_X1 U7842 ( .A1(n5995), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n6187) );
  NAND2_X1 U7843 ( .A1(n6190), .A2(n8313), .ZN(n6193) );
  INV_X1 U7844 ( .A(n6190), .ZN(n6191) );
  NAND2_X1 U7845 ( .A1(n6191), .A2(n8725), .ZN(n6192) );
  NAND2_X1 U7846 ( .A1(n6193), .A2(n6192), .ZN(n8355) );
  NAND2_X1 U7847 ( .A1(n7194), .A2(n8007), .ZN(n6197) );
  AOI22_X1 U7848 ( .A1(n6195), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n8558), .B2(
        n8005), .ZN(n6196) );
  XNOR2_X1 U7849 ( .A(n8878), .B(n6283), .ZN(n6205) );
  NAND2_X1 U7850 ( .A1(n6198), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n6199) );
  NAND2_X1 U7851 ( .A1(n6214), .A2(n6199), .ZN(n8702) );
  NAND2_X1 U7852 ( .A1(n8702), .A2(n6323), .ZN(n6204) );
  INV_X1 U7853 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n9009) );
  NAND2_X1 U7854 ( .A1(n5995), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n6201) );
  NAND2_X1 U7855 ( .A1(n8012), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n6200) );
  OAI211_X1 U7856 ( .C1(n6314), .C2(n9009), .A(n6201), .B(n6200), .ZN(n6202)
         );
  INV_X1 U7857 ( .A(n6202), .ZN(n6203) );
  AND2_X1 U7858 ( .A1(n6205), .A2(n8707), .ZN(n8266) );
  INV_X1 U7859 ( .A(n6205), .ZN(n6206) );
  NAND2_X1 U7860 ( .A1(n6206), .A2(n8687), .ZN(n8267) );
  NAND2_X1 U7861 ( .A1(n7219), .A2(n8007), .ZN(n6208) );
  OR2_X1 U7862 ( .A1(n8008), .A2(n7220), .ZN(n6207) );
  XNOR2_X1 U7863 ( .A(n8872), .B(n6283), .ZN(n6264) );
  XNOR2_X1 U7864 ( .A(n6214), .B(P2_REG3_REG_20__SCAN_IN), .ZN(n8691) );
  INV_X1 U7865 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n8871) );
  NAND2_X1 U7866 ( .A1(n8011), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n6210) );
  NAND2_X1 U7867 ( .A1(n8012), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n6209) );
  OAI211_X1 U7868 ( .C1(n8871), .C2(n4271), .A(n6210), .B(n6209), .ZN(n6211)
         );
  XNOR2_X1 U7869 ( .A(n6264), .B(n8282), .ZN(n8331) );
  NAND2_X1 U7870 ( .A1(n7294), .A2(n8007), .ZN(n6213) );
  OR2_X1 U7871 ( .A1(n8008), .A2(n7297), .ZN(n6212) );
  XNOR2_X1 U7872 ( .A(n8787), .B(n4279), .ZN(n6262) );
  INV_X1 U7873 ( .A(n6214), .ZN(n6216) );
  INV_X1 U7874 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n6215) );
  NAND2_X1 U7875 ( .A1(n6230), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6218) );
  NAND2_X1 U7876 ( .A1(n6252), .A2(n6218), .ZN(n8653) );
  NAND2_X1 U7877 ( .A1(n8653), .A2(n6323), .ZN(n6224) );
  INV_X1 U7878 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n6221) );
  NAND2_X1 U7879 ( .A1(n5995), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n6220) );
  NAND2_X1 U7880 ( .A1(n8012), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n6219) );
  OAI211_X1 U7881 ( .C1(n6314), .C2(n6221), .A(n6220), .B(n6219), .ZN(n6222)
         );
  INV_X1 U7882 ( .A(n6222), .ZN(n6223) );
  NAND2_X1 U7883 ( .A1(n6262), .A2(n8671), .ZN(n8341) );
  NAND2_X1 U7884 ( .A1(n7226), .A2(n8007), .ZN(n6226) );
  OR2_X1 U7885 ( .A1(n8008), .A2(n8981), .ZN(n6225) );
  XNOR2_X1 U7886 ( .A(n8866), .B(n4279), .ZN(n6235) );
  INV_X1 U7887 ( .A(n6235), .ZN(n6234) );
  INV_X1 U7888 ( .A(n6227), .ZN(n6228) );
  NAND2_X1 U7889 ( .A1(n6228), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n6229) );
  NAND2_X1 U7890 ( .A1(n6230), .A2(n6229), .ZN(n8674) );
  INV_X1 U7891 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n8794) );
  NAND2_X1 U7892 ( .A1(n5995), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n6232) );
  NAND2_X1 U7893 ( .A1(n8012), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n6231) );
  OAI211_X1 U7894 ( .C1(n6314), .C2(n8794), .A(n6232), .B(n6231), .ZN(n6233)
         );
  NAND2_X1 U7895 ( .A1(n6234), .A2(n8346), .ZN(n6265) );
  INV_X1 U7896 ( .A(n6265), .ZN(n6236) );
  XNOR2_X1 U7897 ( .A(n6235), .B(n8346), .ZN(n8279) );
  OR2_X1 U7898 ( .A1(n6236), .A2(n8279), .ZN(n8339) );
  NAND2_X1 U7899 ( .A1(n8341), .A2(n8339), .ZN(n6266) );
  OR2_X1 U7900 ( .A1(n8331), .A2(n6266), .ZN(n6401) );
  NAND2_X1 U7901 ( .A1(n7432), .A2(n8007), .ZN(n6238) );
  OR2_X1 U7902 ( .A1(n8008), .A2(n7433), .ZN(n6237) );
  XNOR2_X1 U7903 ( .A(n8853), .B(n6283), .ZN(n6247) );
  NAND2_X1 U7904 ( .A1(n6254), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n6241) );
  NAND2_X1 U7905 ( .A1(n6273), .A2(n6241), .ZN(n8634) );
  NAND2_X1 U7906 ( .A1(n8634), .A2(n6323), .ZN(n6246) );
  INV_X1 U7907 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n8852) );
  NAND2_X1 U7908 ( .A1(n8011), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n6243) );
  NAND2_X1 U7909 ( .A1(n8012), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n6242) );
  OAI211_X1 U7910 ( .C1(n8852), .C2(n4271), .A(n6243), .B(n6242), .ZN(n6244)
         );
  INV_X1 U7911 ( .A(n6244), .ZN(n6245) );
  NAND2_X1 U7912 ( .A1(n6247), .A2(n8621), .ZN(n8288) );
  INV_X1 U7913 ( .A(n6247), .ZN(n6248) );
  NAND2_X1 U7914 ( .A1(n6248), .A2(n8642), .ZN(n6249) );
  NAND2_X1 U7915 ( .A1(n8288), .A2(n6249), .ZN(n6407) );
  NAND2_X1 U7916 ( .A1(n7372), .A2(n8007), .ZN(n6251) );
  OR2_X1 U7917 ( .A1(n8008), .A2(n7375), .ZN(n6250) );
  XNOR2_X1 U7918 ( .A(n8859), .B(n6283), .ZN(n6261) );
  INV_X1 U7919 ( .A(n6261), .ZN(n6405) );
  NAND2_X1 U7920 ( .A1(n6252), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6253) );
  NAND2_X1 U7921 ( .A1(n6254), .A2(n6253), .ZN(n8645) );
  NAND2_X1 U7922 ( .A1(n8645), .A2(n6323), .ZN(n6259) );
  INV_X1 U7923 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n8858) );
  NAND2_X1 U7924 ( .A1(n8011), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n6256) );
  NAND2_X1 U7925 ( .A1(n8012), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n6255) );
  OAI211_X1 U7926 ( .C1(n8858), .C2(n4271), .A(n6256), .B(n6255), .ZN(n6257)
         );
  INV_X1 U7927 ( .A(n6257), .ZN(n6258) );
  AND2_X1 U7928 ( .A1(n6405), .A2(n8651), .ZN(n6260) );
  INV_X1 U7929 ( .A(n6262), .ZN(n6263) );
  INV_X1 U7930 ( .A(n8671), .ZN(n6565) );
  NAND2_X1 U7931 ( .A1(n6263), .A2(n6565), .ZN(n8342) );
  NAND2_X1 U7932 ( .A1(n6264), .A2(n8282), .ZN(n8277) );
  AND2_X1 U7933 ( .A1(n8277), .A2(n6265), .ZN(n8337) );
  OR2_X1 U7934 ( .A1(n6266), .A2(n8337), .ZN(n6267) );
  AND2_X1 U7935 ( .A1(n8342), .A2(n6267), .ZN(n6402) );
  AND2_X1 U7936 ( .A1(n4370), .A2(n6402), .ZN(n6268) );
  NAND2_X1 U7937 ( .A1(n6295), .A2(n8288), .ZN(n6280) );
  NAND2_X1 U7938 ( .A1(n7520), .A2(n8007), .ZN(n6270) );
  OR2_X1 U7939 ( .A1(n8008), .A2(n8983), .ZN(n6269) );
  XNOR2_X1 U7940 ( .A(n8286), .B(n6283), .ZN(n6287) );
  INV_X1 U7941 ( .A(n6273), .ZN(n6272) );
  INV_X1 U7942 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n6271) );
  NAND2_X1 U7943 ( .A1(n6273), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n6274) );
  NAND2_X1 U7944 ( .A1(n6299), .A2(n6274), .ZN(n8623) );
  NAND2_X1 U7945 ( .A1(n8623), .A2(n6323), .ZN(n6279) );
  INV_X1 U7946 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n8965) );
  NAND2_X1 U7947 ( .A1(n8011), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n6276) );
  NAND2_X1 U7948 ( .A1(n8012), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n6275) );
  OAI211_X1 U7949 ( .C1(n8965), .C2(n4271), .A(n6276), .B(n6275), .ZN(n6277)
         );
  INV_X1 U7950 ( .A(n6277), .ZN(n6278) );
  XNOR2_X1 U7951 ( .A(n6287), .B(n8612), .ZN(n8289) );
  NAND2_X1 U7952 ( .A1(n6287), .A2(n8632), .ZN(n6293) );
  NAND2_X1 U7953 ( .A1(n8292), .A2(n6293), .ZN(n6284) );
  NAND2_X1 U7954 ( .A1(n7584), .A2(n8007), .ZN(n6282) );
  OR2_X1 U7955 ( .A1(n8008), .A2(n7686), .ZN(n6281) );
  XNOR2_X1 U7956 ( .A(n8840), .B(n6283), .ZN(n6294) );
  NAND2_X1 U7957 ( .A1(n6284), .A2(n6294), .ZN(n6306) );
  INV_X1 U7958 ( .A(n6294), .ZN(n6289) );
  INV_X1 U7959 ( .A(n6287), .ZN(n6285) );
  NAND2_X1 U7960 ( .A1(n6285), .A2(n8612), .ZN(n6290) );
  NAND2_X1 U7961 ( .A1(n6289), .A2(n6290), .ZN(n6298) );
  NAND2_X1 U7962 ( .A1(n8288), .A2(n8612), .ZN(n6286) );
  NAND2_X1 U7963 ( .A1(n6287), .A2(n6286), .ZN(n6288) );
  OAI211_X1 U7964 ( .C1(n8288), .C2(n8612), .A(n6289), .B(n6288), .ZN(n6292)
         );
  NAND2_X1 U7965 ( .A1(n6294), .A2(n6290), .ZN(n6291) );
  NAND2_X1 U7966 ( .A1(n6292), .A2(n6291), .ZN(n6297) );
  NAND2_X1 U7967 ( .A1(n6299), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n6300) );
  NAND2_X1 U7968 ( .A1(n6310), .A2(n6300), .ZN(n8614) );
  NAND2_X1 U7969 ( .A1(n8614), .A2(n6323), .ZN(n6305) );
  INV_X1 U7970 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n8839) );
  NAND2_X1 U7971 ( .A1(n8011), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n6302) );
  NAND2_X1 U7972 ( .A1(n8012), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n6301) );
  OAI211_X1 U7973 ( .C1(n8839), .C2(n4271), .A(n6302), .B(n6301), .ZN(n6303)
         );
  INV_X1 U7974 ( .A(n6303), .ZN(n6304) );
  NAND2_X1 U7975 ( .A1(n7694), .A2(n8007), .ZN(n6308) );
  OR2_X1 U7976 ( .A1(n8008), .A2(n7695), .ZN(n6307) );
  XNOR2_X1 U7977 ( .A(n8834), .B(n4279), .ZN(n6318) );
  INV_X1 U7978 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n6309) );
  NAND2_X1 U7979 ( .A1(n6310), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n6311) );
  NAND2_X1 U7980 ( .A1(n6321), .A2(n6311), .ZN(n8604) );
  NAND2_X1 U7981 ( .A1(n8604), .A2(n6323), .ZN(n6317) );
  INV_X1 U7982 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n8984) );
  NAND2_X1 U7983 ( .A1(n8012), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n6313) );
  NAND2_X1 U7984 ( .A1(n5995), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n6312) );
  OAI211_X1 U7985 ( .C1(n6314), .C2(n8984), .A(n6313), .B(n6312), .ZN(n6315)
         );
  INV_X1 U7986 ( .A(n6315), .ZN(n6316) );
  XNOR2_X1 U7987 ( .A(n6318), .B(n8611), .ZN(n6505) );
  INV_X1 U7988 ( .A(n6318), .ZN(n6394) );
  NAND2_X1 U7989 ( .A1(n8909), .A2(n8007), .ZN(n6320) );
  OR2_X1 U7990 ( .A1(n8008), .A2(n8912), .ZN(n6319) );
  NAND2_X1 U7991 ( .A1(n6321), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n6322) );
  INV_X1 U7992 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n9028) );
  NAND2_X1 U7993 ( .A1(n8011), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n6325) );
  NAND2_X1 U7994 ( .A1(n8012), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n6324) );
  OAI211_X1 U7995 ( .C1(n9028), .C2(n4271), .A(n6325), .B(n6324), .ZN(n6326)
         );
  INV_X1 U7996 ( .A(n6326), .ZN(n6327) );
  XNOR2_X1 U7997 ( .A(n4279), .B(n8601), .ZN(n6329) );
  XNOR2_X1 U7998 ( .A(n8828), .B(n6329), .ZN(n6363) );
  INV_X1 U7999 ( .A(n6363), .ZN(n6395) );
  XNOR2_X1 U8000 ( .A(n7434), .B(P2_B_REG_SCAN_IN), .ZN(n6336) );
  NAND2_X1 U8001 ( .A1(n7521), .A2(n6336), .ZN(n6342) );
  NAND2_X1 U8002 ( .A1(n6337), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6338) );
  NAND2_X1 U8003 ( .A1(n6339), .A2(n6338), .ZN(n6341) );
  OR2_X1 U8004 ( .A1(n6695), .A2(P2_D_REG_1__SCAN_IN), .ZN(n6344) );
  NAND2_X1 U8005 ( .A1(n7521), .A2(n7685), .ZN(n6700) );
  OR2_X1 U8006 ( .A1(n6695), .A2(P2_D_REG_0__SCAN_IN), .ZN(n6345) );
  NAND2_X1 U8007 ( .A1(n7685), .A2(n7434), .ZN(n6697) );
  NAND2_X1 U8008 ( .A1(n6642), .A2(n6645), .ZN(n6650) );
  NOR2_X1 U8009 ( .A1(P2_D_REG_12__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .ZN(
        n8914) );
  NOR4_X1 U8010 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_7__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n6348) );
  NOR4_X1 U8011 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_28__SCAN_IN), .A3(
        P2_D_REG_27__SCAN_IN), .A4(P2_D_REG_26__SCAN_IN), .ZN(n6347) );
  NOR4_X1 U8012 ( .A1(P2_D_REG_6__SCAN_IN), .A2(P2_D_REG_5__SCAN_IN), .A3(
        P2_D_REG_29__SCAN_IN), .A4(P2_D_REG_30__SCAN_IN), .ZN(n6346) );
  NAND4_X1 U8013 ( .A1(n8914), .A2(n6348), .A3(n6347), .A4(n6346), .ZN(n6354)
         );
  NOR4_X1 U8014 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_18__SCAN_IN), .A3(
        P2_D_REG_15__SCAN_IN), .A4(P2_D_REG_14__SCAN_IN), .ZN(n6352) );
  NOR4_X1 U8015 ( .A1(P2_D_REG_23__SCAN_IN), .A2(P2_D_REG_25__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_9__SCAN_IN), .ZN(n6351) );
  NOR4_X1 U8016 ( .A1(P2_D_REG_10__SCAN_IN), .A2(P2_D_REG_20__SCAN_IN), .A3(
        P2_D_REG_19__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n6350) );
  NOR4_X1 U8017 ( .A1(P2_D_REG_13__SCAN_IN), .A2(P2_D_REG_21__SCAN_IN), .A3(
        P2_D_REG_8__SCAN_IN), .A4(P2_D_REG_11__SCAN_IN), .ZN(n6349) );
  NAND4_X1 U8018 ( .A1(n6352), .A2(n6351), .A3(n6350), .A4(n6349), .ZN(n6353)
         );
  NOR2_X1 U8019 ( .A1(n6354), .A2(n6353), .ZN(n6355) );
  NOR2_X1 U8020 ( .A1(n6695), .A2(n6355), .ZN(n6360) );
  NOR2_X1 U8021 ( .A1(n6650), .A2(n6360), .ZN(n6377) );
  NAND2_X1 U8022 ( .A1(n4396), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6356) );
  NAND2_X1 U8023 ( .A1(n6357), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6358) );
  NAND2_X1 U8024 ( .A1(n8558), .A2(n8229), .ZN(n6579) );
  NAND2_X1 U8025 ( .A1(n5922), .A2(n8205), .ZN(n8172) );
  AND2_X1 U8026 ( .A1(n8158), .A2(n8792), .ZN(n6359) );
  NAND2_X1 U8027 ( .A1(n6627), .A2(n6378), .ZN(n6362) );
  INV_X1 U8028 ( .A(n6642), .ZN(n6895) );
  INV_X1 U8029 ( .A(n6645), .ZN(n6894) );
  INV_X1 U8030 ( .A(n6360), .ZN(n6639) );
  NAND2_X1 U8031 ( .A1(n6381), .A2(n6696), .ZN(n6630) );
  OR2_X1 U8032 ( .A1(n6630), .A2(n6625), .ZN(n6361) );
  OAI211_X1 U8033 ( .C1(n6606), .C2(n6394), .A(n6395), .B(n8367), .ZN(n6400)
         );
  NAND2_X1 U8034 ( .A1(n6514), .A2(n6364), .ZN(n6399) );
  NAND2_X1 U8035 ( .A1(n6627), .A2(n10216), .ZN(n6366) );
  INV_X1 U8036 ( .A(n6900), .ZN(n6365) );
  INV_X1 U8037 ( .A(n8558), .ZN(n8573) );
  NAND2_X1 U8038 ( .A1(n8573), .A2(n8215), .ZN(n6382) );
  OR2_X1 U8039 ( .A1(n6382), .A2(n8158), .ZN(n6936) );
  OR2_X1 U8040 ( .A1(n6630), .A2(n6936), .ZN(n6376) );
  INV_X1 U8041 ( .A(n6376), .ZN(n6369) );
  INV_X1 U8042 ( .A(n6726), .ZN(n8226) );
  NAND2_X1 U8043 ( .A1(n8226), .A2(n8564), .ZN(n6368) );
  INV_X1 U8044 ( .A(n8246), .ZN(n6370) );
  NAND2_X1 U8045 ( .A1(n6370), .A2(n6323), .ZN(n8014) );
  INV_X1 U8046 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n6373) );
  NAND2_X1 U8047 ( .A1(n8012), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n6372) );
  NAND2_X1 U8048 ( .A1(n8011), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n6371) );
  OAI211_X1 U8049 ( .C1(n6373), .C2(n4271), .A(n6372), .B(n6371), .ZN(n6374)
         );
  INV_X1 U8050 ( .A(n6374), .ZN(n6375) );
  NAND2_X1 U8051 ( .A1(n8014), .A2(n6375), .ZN(n8588) );
  NAND2_X1 U8052 ( .A1(n8588), .A2(n8371), .ZN(n6393) );
  INV_X1 U8053 ( .A(n6377), .ZN(n6380) );
  INV_X1 U8054 ( .A(n6378), .ZN(n6379) );
  NAND2_X1 U8055 ( .A1(n6900), .A2(n10216), .ZN(n8628) );
  NAND2_X1 U8056 ( .A1(n6379), .A2(n8628), .ZN(n6628) );
  NAND2_X1 U8057 ( .A1(n6380), .A2(n6628), .ZN(n6386) );
  INV_X1 U8058 ( .A(n6381), .ZN(n6389) );
  INV_X1 U8059 ( .A(n6625), .ZN(n6384) );
  NAND2_X1 U8060 ( .A1(n6382), .A2(n8165), .ZN(n6383) );
  NAND3_X1 U8061 ( .A1(n6383), .A2(n6716), .A3(n6718), .ZN(n6637) );
  AOI21_X1 U8062 ( .B1(n6389), .B2(n6384), .A(n6637), .ZN(n6385) );
  NAND2_X1 U8063 ( .A1(n6386), .A2(n6385), .ZN(n6387) );
  NAND2_X1 U8064 ( .A1(n6387), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6391) );
  INV_X1 U8065 ( .A(n6696), .ZN(n6388) );
  NOR2_X1 U8066 ( .A1(n6388), .A2(n6936), .ZN(n8227) );
  NAND2_X1 U8067 ( .A1(n6389), .A2(n8227), .ZN(n6390) );
  NAND2_X2 U8068 ( .A1(n6391), .A2(n6390), .ZN(n8385) );
  AOI22_X1 U8069 ( .A1(n8594), .A2(n8385), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3151), .ZN(n6392) );
  OAI211_X1 U8070 ( .C1(n6606), .C2(n8382), .A(n6393), .B(n6392), .ZN(n6397)
         );
  NOR4_X1 U8071 ( .A1(n6395), .A2(n6394), .A3(n6606), .A4(n8375), .ZN(n6396)
         );
  AOI211_X1 U8072 ( .C1(n8828), .C2(n8362), .A(n6397), .B(n6396), .ZN(n6398)
         );
  OAI211_X1 U8073 ( .C1(n6514), .C2(n6400), .A(n6399), .B(n6398), .ZN(P2_U3160) );
  AOI21_X1 U8074 ( .B1(n6408), .B2(n8287), .A(n8375), .ZN(n6415) );
  INV_X1 U8075 ( .A(n8380), .ZN(n8360) );
  AOI22_X1 U8076 ( .A1(n8651), .A2(n8356), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3151), .ZN(n6410) );
  NAND2_X1 U8077 ( .A1(n8634), .A2(n8385), .ZN(n6409) );
  OAI211_X1 U8078 ( .C1(n8632), .C2(n8360), .A(n6410), .B(n6409), .ZN(n6411)
         );
  INV_X1 U8079 ( .A(n6411), .ZN(n6413) );
  NAND2_X1 U8080 ( .A1(n8853), .A2(n8362), .ZN(n6412) );
  NAND2_X1 U8081 ( .A1(n6413), .A2(n6412), .ZN(n6414) );
  NAND2_X1 U8082 ( .A1(n6849), .A2(n10043), .ZN(n6416) );
  NAND2_X1 U8083 ( .A1(n6990), .A2(n6416), .ZN(n6418) );
  NAND2_X1 U8084 ( .A1(n6853), .A2(n6992), .ZN(n6417) );
  NAND2_X1 U8085 ( .A1(n6418), .A2(n6417), .ZN(n10032) );
  NAND2_X1 U8086 ( .A1(n10032), .A2(n6419), .ZN(n6422) );
  CLKBUF_X2 U8087 ( .A(n6420), .Z(n10060) );
  NAND2_X1 U8088 ( .A1(n6854), .A2(n10060), .ZN(n6421) );
  NAND2_X1 U8089 ( .A1(n6422), .A2(n6421), .ZN(n7026) );
  NAND2_X1 U8090 ( .A1(n7026), .A2(n7027), .ZN(n6424) );
  NAND2_X1 U8091 ( .A1(n7038), .A2(n10066), .ZN(n6423) );
  NAND2_X1 U8092 ( .A1(n6424), .A2(n6423), .ZN(n7127) );
  NAND2_X1 U8093 ( .A1(n7127), .A2(n7130), .ZN(n10019) );
  OAI21_X1 U8094 ( .B1(n10015), .B2(n4993), .A(n6426), .ZN(n6427) );
  INV_X1 U8095 ( .A(n6427), .ZN(n6428) );
  OAI21_X1 U8096 ( .B1(n10019), .B2(n10015), .A(n6428), .ZN(n7205) );
  NAND2_X1 U8097 ( .A1(n7242), .A2(n6429), .ZN(n7207) );
  INV_X1 U8098 ( .A(n9218), .ZN(n9372) );
  OR2_X1 U8099 ( .A1(n10083), .A2(n9372), .ZN(n6430) );
  OR2_X1 U8100 ( .A1(n10007), .A2(n9371), .ZN(n6432) );
  NAND2_X1 U8101 ( .A1(n6433), .A2(n7322), .ZN(n7319) );
  INV_X1 U8102 ( .A(n9069), .ZN(n9370) );
  INV_X1 U8103 ( .A(n7841), .ZN(n10104) );
  NOR2_X1 U8104 ( .A1(n5461), .A2(n9365), .ZN(n6440) );
  INV_X1 U8105 ( .A(n9914), .ZN(n7748) );
  AOI21_X1 U8106 ( .B1(n9811), .B2(n4697), .A(n6442), .ZN(n9794) );
  NAND2_X1 U8107 ( .A1(n9903), .A2(n9362), .ZN(n6443) );
  NAND2_X1 U8108 ( .A1(n9794), .A2(n6443), .ZN(n6446) );
  INV_X1 U8109 ( .A(n9903), .ZN(n9799) );
  NAND2_X1 U8110 ( .A1(n9799), .A2(n6444), .ZN(n6445) );
  INV_X1 U8111 ( .A(n9898), .ZN(n6447) );
  NAND2_X1 U8112 ( .A1(n9882), .A2(n9358), .ZN(n6452) );
  NAND2_X1 U8113 ( .A1(n9749), .A2(n6452), .ZN(n6454) );
  NAND2_X1 U8114 ( .A1(n9747), .A2(n9285), .ZN(n6453) );
  NAND2_X1 U8115 ( .A1(n9878), .A2(n9357), .ZN(n6456) );
  NOR2_X1 U8116 ( .A1(n9878), .A2(n9357), .ZN(n6455) );
  NAND2_X1 U8117 ( .A1(n9869), .A2(n9355), .ZN(n6457) );
  NAND2_X1 U8118 ( .A1(n9702), .A2(n9095), .ZN(n6458) );
  NOR2_X1 U8119 ( .A1(n9863), .A2(n9354), .ZN(n6460) );
  NAND2_X1 U8120 ( .A1(n9673), .A2(n9196), .ZN(n6461) );
  NAND2_X1 U8121 ( .A1(n9652), .A2(n9330), .ZN(n6462) );
  INV_X1 U8122 ( .A(n6478), .ZN(n6463) );
  XNOR2_X1 U8123 ( .A(n9611), .B(n6463), .ZN(n9635) );
  OR2_X1 U8124 ( .A1(n6787), .A2(n6785), .ZN(n6465) );
  INV_X1 U8125 ( .A(n6464), .ZN(n7239) );
  INV_X1 U8126 ( .A(n6797), .ZN(n6748) );
  AND2_X1 U8127 ( .A1(n6465), .A2(n6748), .ZN(n6978) );
  INV_X1 U8128 ( .A(n6802), .ZN(n6466) );
  NAND2_X1 U8129 ( .A1(n6787), .A2(n6466), .ZN(n6467) );
  NAND2_X1 U8130 ( .A1(n6978), .A2(n6467), .ZN(n7028) );
  NAND2_X1 U8131 ( .A1(n9635), .A2(n10107), .ZN(n6488) );
  OAI21_X1 U8132 ( .B1(n9658), .B2(n9657), .A(n6476), .ZN(n6477) );
  NAND2_X1 U8133 ( .A1(n6477), .A2(n6478), .ZN(n9622) );
  OAI21_X1 U8134 ( .B1(n6478), .B2(n6477), .A(n9622), .ZN(n6481) );
  NAND2_X1 U8135 ( .A1(n4471), .A2(n9630), .ZN(n6480) );
  NAND2_X1 U8136 ( .A1(n6677), .A2(n8232), .ZN(n9329) );
  OAI22_X1 U8137 ( .A1(n9330), .A2(n9626), .B1(n7171), .B2(n9329), .ZN(n9138)
         );
  NAND2_X1 U8138 ( .A1(n6991), .A2(n6992), .ZN(n10034) );
  NAND2_X1 U8139 ( .A1(n7029), .A2(n10066), .ZN(n7030) );
  INV_X1 U8140 ( .A(n10083), .ZN(n7215) );
  INV_X1 U8141 ( .A(n10007), .ZN(n10091) );
  NOR2_X4 U8142 ( .A1(n4986), .A2(n5388), .ZN(n7351) );
  AND2_X2 U8143 ( .A1(n7351), .A2(n10104), .ZN(n7349) );
  INV_X1 U8144 ( .A(n9299), .ZN(n7478) );
  INV_X2 U8145 ( .A(n6483), .ZN(n7744) );
  NAND2_X1 U8146 ( .A1(n9770), .A2(n9775), .ZN(n9757) );
  OR2_X2 U8147 ( .A1(n9757), .A2(n9888), .ZN(n9758) );
  INV_X1 U8148 ( .A(n9878), .ZN(n9725) );
  NAND2_X1 U8149 ( .A1(n9649), .A2(n9652), .ZN(n6484) );
  OR2_X2 U8150 ( .A1(n6484), .A2(n9636), .ZN(n9618) );
  INV_X1 U8151 ( .A(n9618), .ZN(n6485) );
  AOI211_X1 U8152 ( .C1(n9636), .C2(n6484), .A(n8236), .B(n6485), .ZN(n9644)
         );
  AOI21_X1 U8153 ( .B1(n10084), .B2(n9636), .A(n9644), .ZN(n6486) );
  NAND2_X1 U8154 ( .A1(n6488), .A2(n6487), .ZN(n9848) );
  OR2_X1 U8155 ( .A1(n6794), .A2(n6802), .ZN(n6777) );
  NAND2_X1 U8156 ( .A1(n7557), .A2(P1_B_REG_SCAN_IN), .ZN(n6489) );
  MUX2_X1 U8157 ( .A(P1_B_REG_SCAN_IN), .B(n6489), .S(n7447), .Z(n6491) );
  NAND2_X1 U8158 ( .A1(n7557), .A2(n7586), .ZN(n9953) );
  OAI21_X1 U8159 ( .B1(n9952), .B2(P1_D_REG_1__SCAN_IN), .A(n9953), .ZN(n6502)
         );
  NOR4_X1 U8160 ( .A1(P1_D_REG_14__SCAN_IN), .A2(P1_D_REG_16__SCAN_IN), .A3(
        P1_D_REG_19__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n6495) );
  NOR4_X1 U8161 ( .A1(P1_D_REG_11__SCAN_IN), .A2(P1_D_REG_12__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n6494) );
  NOR4_X1 U8162 ( .A1(P1_D_REG_25__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_27__SCAN_IN), .A4(P1_D_REG_28__SCAN_IN), .ZN(n6493) );
  NOR4_X1 U8163 ( .A1(P1_D_REG_21__SCAN_IN), .A2(P1_D_REG_24__SCAN_IN), .A3(
        P1_D_REG_22__SCAN_IN), .A4(P1_D_REG_23__SCAN_IN), .ZN(n6492) );
  NAND4_X1 U8164 ( .A1(n6495), .A2(n6494), .A3(n6493), .A4(n6492), .ZN(n6500)
         );
  NOR2_X1 U8165 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_29__SCAN_IN), .ZN(
        n8915) );
  NOR4_X1 U8166 ( .A1(P1_D_REG_30__SCAN_IN), .A2(P1_D_REG_31__SCAN_IN), .A3(
        P1_D_REG_18__SCAN_IN), .A4(P1_D_REG_2__SCAN_IN), .ZN(n6498) );
  NOR4_X1 U8167 ( .A1(P1_D_REG_7__SCAN_IN), .A2(P1_D_REG_8__SCAN_IN), .A3(
        P1_D_REG_9__SCAN_IN), .A4(P1_D_REG_10__SCAN_IN), .ZN(n6497) );
  NOR4_X1 U8168 ( .A1(P1_D_REG_3__SCAN_IN), .A2(P1_D_REG_4__SCAN_IN), .A3(
        P1_D_REG_5__SCAN_IN), .A4(P1_D_REG_6__SCAN_IN), .ZN(n6496) );
  NAND4_X1 U8169 ( .A1(n8915), .A2(n6498), .A3(n6497), .A4(n6496), .ZN(n6499)
         );
  NOR2_X1 U8170 ( .A1(n6500), .A2(n6499), .ZN(n6772) );
  NAND2_X1 U8171 ( .A1(n7447), .A2(n7586), .ZN(n9954) );
  INV_X1 U8172 ( .A(n7000), .ZN(n6776) );
  NAND2_X1 U8173 ( .A1(n9848), .A2(n4272), .ZN(n6504) );
  NAND2_X1 U8174 ( .A1(n6504), .A2(n6503), .ZN(P1_U3518) );
  NAND2_X1 U8175 ( .A1(n8834), .A2(n8362), .ZN(n6512) );
  NAND2_X1 U8176 ( .A1(n8601), .A2(n8380), .ZN(n6509) );
  AOI22_X1 U8177 ( .A1(n8604), .A2(n8385), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3151), .ZN(n6508) );
  OAI211_X1 U8178 ( .C1(n8620), .C2(n8382), .A(n6509), .B(n6508), .ZN(n6510)
         );
  INV_X1 U8179 ( .A(n6741), .ZN(n8404) );
  NAND2_X1 U8180 ( .A1(n8404), .A2(n6742), .ZN(n6903) );
  NAND2_X1 U8181 ( .A1(n6515), .A2(n6517), .ZN(n8174) );
  NAND2_X1 U8182 ( .A1(n6516), .A2(n6517), .ZN(n6518) );
  NAND2_X1 U8183 ( .A1(n6519), .A2(n7093), .ZN(n6520) );
  INV_X1 U8184 ( .A(n10195), .ZN(n6522) );
  NAND2_X1 U8185 ( .A1(n6523), .A2(n6522), .ZN(n6524) );
  INV_X1 U8186 ( .A(n10200), .ZN(n7162) );
  NAND2_X1 U8187 ( .A1(n6525), .A2(n8402), .ZN(n6529) );
  INV_X1 U8188 ( .A(n7162), .ZN(n6526) );
  NAND2_X1 U8189 ( .A1(n6527), .A2(n6526), .ZN(n6528) );
  NAND2_X1 U8190 ( .A1(n6529), .A2(n6528), .ZN(n7231) );
  AND2_X1 U8191 ( .A1(n10174), .A2(n10205), .ZN(n6530) );
  NAND2_X1 U8192 ( .A1(n7485), .A2(n6531), .ZN(n8066) );
  NAND2_X1 U8193 ( .A1(n7465), .A2(n8399), .ZN(n7727) );
  NAND2_X1 U8194 ( .A1(n4901), .A2(n7727), .ZN(n6533) );
  OR2_X1 U8195 ( .A1(n7465), .A2(n8322), .ZN(n8056) );
  NAND2_X1 U8196 ( .A1(n7465), .A2(n8322), .ZN(n8067) );
  NOR2_X1 U8197 ( .A1(n7485), .A2(n8400), .ZN(n7451) );
  INV_X1 U8198 ( .A(n8324), .ZN(n7758) );
  AOI22_X1 U8199 ( .A1(n7452), .A2(n7727), .B1(n7767), .B2(n7758), .ZN(n6532)
         );
  NAND2_X1 U8200 ( .A1(n8324), .A2(n8398), .ZN(n6534) );
  OR2_X1 U8201 ( .A1(n7770), .A2(n8397), .ZN(n7590) );
  AND2_X1 U8202 ( .A1(n7636), .A2(n8395), .ZN(n6541) );
  NAND2_X1 U8203 ( .A1(n6536), .A2(n8396), .ZN(n6540) );
  INV_X1 U8204 ( .A(n6540), .ZN(n6537) );
  AND2_X1 U8205 ( .A1(n7590), .A2(n6539), .ZN(n6538) );
  NAND2_X1 U8206 ( .A1(n7591), .A2(n6538), .ZN(n6546) );
  INV_X1 U8207 ( .A(n6539), .ZN(n6544) );
  NAND2_X1 U8208 ( .A1(n7770), .A2(n8397), .ZN(n7592) );
  AND2_X1 U8209 ( .A1(n7592), .A2(n6540), .ZN(n7612) );
  INV_X1 U8210 ( .A(n6541), .ZN(n6542) );
  AND2_X1 U8211 ( .A1(n7612), .A2(n6542), .ZN(n6543) );
  OR2_X1 U8212 ( .A1(n6544), .A2(n6543), .ZN(n6545) );
  NAND2_X1 U8213 ( .A1(n6546), .A2(n6545), .ZN(n6548) );
  OR2_X1 U8214 ( .A1(n7636), .A2(n8395), .ZN(n6547) );
  XNOR2_X1 U8215 ( .A(n8093), .B(n7793), .ZN(n8096) );
  NOR2_X1 U8216 ( .A1(n8093), .A2(n8394), .ZN(n8095) );
  AND2_X1 U8217 ( .A1(n7993), .A2(n8383), .ZN(n7721) );
  INV_X1 U8218 ( .A(n7721), .ZN(n8098) );
  OR2_X1 U8219 ( .A1(n8814), .A2(n8392), .ZN(n7714) );
  NAND2_X1 U8220 ( .A1(n7710), .A2(n6549), .ZN(n6551) );
  NAND2_X1 U8221 ( .A1(n6553), .A2(n8724), .ZN(n8720) );
  AND2_X1 U8222 ( .A1(n7993), .A2(n8393), .ZN(n7711) );
  NAND2_X1 U8223 ( .A1(n7714), .A2(n7711), .ZN(n6550) );
  NAND2_X1 U8224 ( .A1(n8814), .A2(n8392), .ZN(n8718) );
  NAND2_X1 U8225 ( .A1(n6552), .A2(n8740), .ZN(n8677) );
  INV_X1 U8226 ( .A(n8724), .ZN(n8300) );
  NAND2_X1 U8227 ( .A1(n6553), .A2(n8300), .ZN(n8101) );
  NAND2_X1 U8228 ( .A1(n8111), .A2(n8101), .ZN(n8734) );
  INV_X1 U8229 ( .A(n8720), .ZN(n6554) );
  NOR2_X1 U8230 ( .A1(n8734), .A2(n6554), .ZN(n6555) );
  INV_X1 U8231 ( .A(n6552), .ZN(n8314) );
  INV_X1 U8232 ( .A(n8803), .ZN(n6558) );
  NAND2_X1 U8233 ( .A1(n6558), .A2(n8313), .ZN(n6559) );
  NAND2_X1 U8234 ( .A1(n8878), .A2(n8707), .ZN(n8680) );
  NAND2_X1 U8235 ( .A1(n8107), .A2(n8680), .ZN(n8697) );
  INV_X1 U8236 ( .A(n8697), .ZN(n6560) );
  INV_X1 U8237 ( .A(n8878), .ZN(n8272) );
  NAND2_X1 U8238 ( .A1(n8866), .A2(n8346), .ZN(n8127) );
  NAND2_X1 U8239 ( .A1(n8128), .A2(n8127), .ZN(n8664) );
  INV_X1 U8240 ( .A(n8664), .ZN(n8668) );
  NOR2_X1 U8241 ( .A1(n8872), .A2(n8282), .ZN(n6602) );
  INV_X1 U8242 ( .A(n6602), .ZN(n8122) );
  NAND2_X1 U8243 ( .A1(n8872), .A2(n8282), .ZN(n8663) );
  NAND2_X1 U8244 ( .A1(n8664), .A2(n6561), .ZN(n6564) );
  INV_X1 U8245 ( .A(n8282), .ZN(n8699) );
  OR2_X1 U8246 ( .A1(n8872), .A2(n8699), .ZN(n8667) );
  OR2_X1 U8247 ( .A1(n8866), .A2(n8688), .ZN(n8648) );
  OAI21_X1 U8248 ( .B1(n8668), .B2(n8667), .A(n8648), .ZN(n6562) );
  NAND2_X1 U8249 ( .A1(n8787), .A2(n6565), .ZN(n8132) );
  INV_X1 U8250 ( .A(n8658), .ZN(n8199) );
  NAND2_X1 U8251 ( .A1(n8859), .A2(n8651), .ZN(n6568) );
  INV_X1 U8252 ( .A(n8859), .ZN(n8265) );
  INV_X1 U8253 ( .A(n8853), .ZN(n8781) );
  NAND2_X1 U8254 ( .A1(n8781), .A2(n8621), .ZN(n6570) );
  NAND2_X1 U8255 ( .A1(n8286), .A2(n8612), .ZN(n8148) );
  OR2_X1 U8256 ( .A1(n8286), .A2(n8612), .ZN(n8149) );
  INV_X1 U8257 ( .A(n8149), .ZN(n6571) );
  INV_X1 U8258 ( .A(n8840), .ZN(n8374) );
  NAND2_X1 U8259 ( .A1(n8374), .A2(n8620), .ZN(n6573) );
  INV_X1 U8260 ( .A(n8834), .ZN(n6574) );
  NAND2_X1 U8261 ( .A1(n8904), .A2(n8007), .ZN(n6576) );
  INV_X1 U8262 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n8906) );
  OR2_X1 U8263 ( .A1(n8008), .A2(n8906), .ZN(n6575) );
  NAND2_X1 U8264 ( .A1(n6576), .A2(n6575), .ZN(n6635) );
  INV_X1 U8265 ( .A(n8588), .ZN(n6577) );
  NAND2_X1 U8266 ( .A1(n6635), .A2(n6577), .ZN(n8016) );
  NAND2_X1 U8267 ( .A1(n8167), .A2(n8016), .ZN(n8161) );
  XNOR2_X1 U8268 ( .A(n6578), .B(n8162), .ZN(n6622) );
  INV_X1 U8269 ( .A(n8022), .ZN(n6580) );
  NAND2_X1 U8270 ( .A1(n6580), .A2(n8174), .ZN(n6893) );
  NAND2_X1 U8271 ( .A1(n6893), .A2(n6581), .ZN(n8749) );
  INV_X1 U8272 ( .A(n8031), .ZN(n8750) );
  NAND2_X1 U8273 ( .A1(n8749), .A2(n8750), .ZN(n6582) );
  NAND2_X1 U8274 ( .A1(n6582), .A2(n8027), .ZN(n7014) );
  NAND2_X1 U8275 ( .A1(n6583), .A2(n8033), .ZN(n10179) );
  OR2_X1 U8276 ( .A1(n7229), .A2(n10200), .ZN(n8035) );
  NAND2_X1 U8277 ( .A1(n10179), .A2(n8035), .ZN(n6584) );
  NAND2_X1 U8278 ( .A1(n7229), .A2(n10200), .ZN(n8046) );
  NAND2_X1 U8279 ( .A1(n6584), .A2(n8046), .ZN(n7227) );
  INV_X1 U8280 ( .A(n10205), .ZN(n7228) );
  NAND2_X1 U8281 ( .A1(n7228), .A2(n10174), .ZN(n8034) );
  NAND2_X1 U8282 ( .A1(n7227), .A2(n8034), .ZN(n7255) );
  NAND2_X1 U8283 ( .A1(n10215), .A2(n7230), .ZN(n8050) );
  NAND2_X1 U8284 ( .A1(n7201), .A2(n10205), .ZN(n8047) );
  AND2_X1 U8285 ( .A1(n8050), .A2(n8047), .ZN(n8040) );
  AND2_X1 U8286 ( .A1(n8056), .A2(n7448), .ZN(n8062) );
  OR2_X1 U8287 ( .A1(n7770), .A2(n7782), .ZN(n8079) );
  OR2_X1 U8288 ( .A1(n8324), .A2(n7767), .ZN(n8057) );
  AND2_X1 U8289 ( .A1(n8079), .A2(n8057), .ZN(n8061) );
  NAND2_X1 U8290 ( .A1(n7490), .A2(n8061), .ZN(n6590) );
  NAND2_X1 U8291 ( .A1(n8324), .A2(n7767), .ZN(n8068) );
  NAND2_X1 U8292 ( .A1(n8068), .A2(n8397), .ZN(n6587) );
  INV_X1 U8293 ( .A(n8068), .ZN(n6586) );
  AOI22_X1 U8294 ( .A1(n7770), .A2(n6587), .B1(n6586), .B2(n7782), .ZN(n6588)
         );
  AND2_X1 U8295 ( .A1(n6588), .A2(n8081), .ZN(n6589) );
  NAND2_X1 U8296 ( .A1(n6590), .A2(n6589), .ZN(n6591) );
  NAND2_X1 U8297 ( .A1(n6591), .A2(n8080), .ZN(n7611) );
  NAND2_X1 U8298 ( .A1(n7636), .A2(n7626), .ZN(n8087) );
  NAND2_X1 U8299 ( .A1(n8088), .A2(n8087), .ZN(n8188) );
  NAND2_X1 U8300 ( .A1(n7611), .A2(n8092), .ZN(n6592) );
  NAND2_X1 U8301 ( .A1(n6592), .A2(n8088), .ZN(n7601) );
  NOR2_X1 U8302 ( .A1(n8093), .A2(n7793), .ZN(n6594) );
  NAND2_X1 U8303 ( .A1(n8093), .A2(n7793), .ZN(n6593) );
  INV_X1 U8304 ( .A(n8392), .ZN(n8738) );
  AND2_X1 U8305 ( .A1(n8814), .A2(n8738), .ZN(n6595) );
  OR2_X1 U8306 ( .A1(n7721), .A2(n6595), .ZN(n6598) );
  OR2_X1 U8307 ( .A1(n8814), .A2(n8738), .ZN(n8100) );
  OR2_X1 U8308 ( .A1(n6595), .A2(n8097), .ZN(n6596) );
  AND2_X1 U8309 ( .A1(n8100), .A2(n6596), .ZN(n6597) );
  NAND2_X1 U8310 ( .A1(n8803), .A2(n8313), .ZN(n8195) );
  NAND2_X1 U8311 ( .A1(n8195), .A2(n8680), .ZN(n6600) );
  INV_X1 U8312 ( .A(n8677), .ZN(n6599) );
  NOR2_X1 U8313 ( .A1(n6600), .A2(n6599), .ZN(n6601) );
  NAND2_X1 U8314 ( .A1(n8678), .A2(n6601), .ZN(n6604) );
  NAND2_X1 U8315 ( .A1(n8694), .A2(n8107), .ZN(n8681) );
  AOI21_X1 U8316 ( .B1(n8680), .B2(n8681), .A(n6602), .ZN(n6603) );
  NAND2_X1 U8317 ( .A1(n6604), .A2(n6603), .ZN(n8662) );
  AND2_X1 U8318 ( .A1(n8127), .A2(n8663), .ZN(n8123) );
  NAND2_X1 U8319 ( .A1(n8662), .A2(n8123), .ZN(n6605) );
  NOR2_X1 U8320 ( .A1(n8859), .A2(n8631), .ZN(n8134) );
  NAND2_X1 U8321 ( .A1(n8859), .A2(n8631), .ZN(n8197) );
  NOR2_X1 U8322 ( .A1(n8286), .A2(n8632), .ZN(n8150) );
  NAND2_X1 U8323 ( .A1(n8286), .A2(n8632), .ZN(n8151) );
  NAND2_X1 U8324 ( .A1(n8840), .A2(n8620), .ZN(n8156) );
  NAND2_X1 U8325 ( .A1(n8155), .A2(n8156), .ZN(n8608) );
  NAND2_X1 U8326 ( .A1(n8834), .A2(n6606), .ZN(n8159) );
  NAND2_X1 U8327 ( .A1(n7295), .A2(n8205), .ZN(n6607) );
  NAND2_X1 U8328 ( .A1(n8792), .A2(n6607), .ZN(n6608) );
  NOR2_X1 U8329 ( .A1(n8558), .A2(n6608), .ZN(n6609) );
  NAND2_X1 U8330 ( .A1(n6623), .A2(n8756), .ZN(n6620) );
  INV_X1 U8331 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n8826) );
  NAND2_X1 U8332 ( .A1(n8011), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n6611) );
  INV_X1 U8333 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n8584) );
  OR2_X1 U8334 ( .A1(n4286), .A2(n8584), .ZN(n6610) );
  OAI211_X1 U8335 ( .C1(n8826), .C2(n4271), .A(n6611), .B(n6610), .ZN(n6612)
         );
  INV_X1 U8336 ( .A(n6612), .ZN(n6613) );
  NAND2_X1 U8337 ( .A1(n6614), .A2(P2_B_REG_SCAN_IN), .ZN(n6615) );
  NAND2_X1 U8338 ( .A1(n10173), .A2(n6615), .ZN(n8577) );
  NAND2_X1 U8339 ( .A1(n8601), .A2(n10175), .ZN(n6617) );
  OAI21_X1 U8340 ( .B1(n8017), .B2(n8577), .A(n6617), .ZN(n6618) );
  INV_X1 U8341 ( .A(n6618), .ZN(n6619) );
  NAND2_X1 U8342 ( .A1(n6620), .A2(n6619), .ZN(n6621) );
  NAND2_X1 U8343 ( .A1(n6936), .A2(n6625), .ZN(n6626) );
  NAND2_X1 U8344 ( .A1(n6627), .A2(n6626), .ZN(n6632) );
  INV_X1 U8345 ( .A(n6628), .ZN(n6629) );
  NAND2_X1 U8346 ( .A1(n10219), .A2(n6373), .ZN(n6633) );
  NAND2_X1 U8347 ( .A1(n6634), .A2(n6633), .ZN(n6636) );
  NAND2_X1 U8348 ( .A1(n6636), .A2(n4992), .ZN(P2_U3456) );
  NOR2_X1 U8349 ( .A1(n6637), .A2(P2_U3151), .ZN(n6638) );
  NAND2_X1 U8350 ( .A1(n8205), .A2(n8229), .ZN(n6640) );
  OR2_X1 U8351 ( .A1(n8558), .A2(n6640), .ZN(n6641) );
  NAND2_X1 U8352 ( .A1(n6641), .A2(n8158), .ZN(n6643) );
  NAND2_X1 U8353 ( .A1(n6642), .A2(n6643), .ZN(n6647) );
  INV_X1 U8354 ( .A(n6643), .ZN(n6644) );
  NAND2_X1 U8355 ( .A1(n6645), .A2(n6644), .ZN(n6646) );
  NAND2_X1 U8356 ( .A1(n6647), .A2(n6646), .ZN(n6898) );
  INV_X1 U8357 ( .A(n6648), .ZN(n6649) );
  NAND2_X1 U8358 ( .A1(n10227), .A2(n6652), .ZN(n6653) );
  NAND2_X1 U8359 ( .A1(n6654), .A2(n4982), .ZN(P2_U3488) );
  NOR2_X1 U8360 ( .A1(n6790), .A2(P1_U3086), .ZN(n6655) );
  NAND2_X2 U8361 ( .A1(n8003), .A2(P1_U3086), .ZN(n8253) );
  INV_X1 U8362 ( .A(n9414), .ZN(n6810) );
  OAI222_X1 U8363 ( .A1(n8253), .A2(n8922), .B1(n9963), .B2(n9058), .C1(
        P1_U3086), .C2(n6810), .ZN(P1_U3352) );
  INV_X1 U8364 ( .A(n9401), .ZN(n6807) );
  OAI222_X1 U8365 ( .A1(n8253), .A2(n6657), .B1(n9963), .B2(n6667), .C1(
        P1_U3086), .C2(n6807), .ZN(P1_U3353) );
  NAND2_X2 U8366 ( .A1(n6658), .A2(P2_U3151), .ZN(n8905) );
  INV_X2 U8367 ( .A(n8908), .ZN(n9059) );
  INV_X1 U8368 ( .A(n6659), .ZN(n6690) );
  INV_X1 U8369 ( .A(n6767), .ZN(n6871) );
  OAI222_X1 U8370 ( .A1(n8905), .A2(n6660), .B1(n9059), .B2(n6690), .C1(
        P2_U3151), .C2(n6871), .ZN(P2_U3294) );
  INV_X1 U8371 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6662) );
  INV_X1 U8372 ( .A(n6661), .ZN(n6673) );
  INV_X1 U8373 ( .A(n9441), .ZN(n6812) );
  OAI222_X1 U8374 ( .A1(n8253), .A2(n6662), .B1(n9963), .B2(n6673), .C1(
        P1_U3086), .C2(n6812), .ZN(P1_U3350) );
  INV_X1 U8375 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6664) );
  INV_X1 U8376 ( .A(n6663), .ZN(n6669) );
  INV_X1 U8377 ( .A(n9454), .ZN(n6814) );
  OAI222_X1 U8378 ( .A1(n8253), .A2(n6664), .B1(n9963), .B2(n6669), .C1(
        P1_U3086), .C2(n6814), .ZN(P1_U3349) );
  INV_X1 U8379 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6666) );
  INV_X1 U8380 ( .A(n6665), .ZN(n6671) );
  INV_X1 U8381 ( .A(n9427), .ZN(n6811) );
  OAI222_X1 U8382 ( .A1(n8253), .A2(n6666), .B1(n9963), .B2(n6671), .C1(
        P1_U3086), .C2(n6811), .ZN(P1_U3351) );
  OAI222_X1 U8383 ( .A1(n8905), .A2(n6668), .B1(n9059), .B2(n6667), .C1(
        P2_U3151), .C2(n4458), .ZN(P2_U3293) );
  INV_X1 U8384 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6670) );
  INV_X1 U8385 ( .A(n7185), .ZN(n7085) );
  OAI222_X1 U8386 ( .A1(n8905), .A2(n6670), .B1(n9059), .B2(n6669), .C1(
        P2_U3151), .C2(n7085), .ZN(P2_U3289) );
  INV_X1 U8387 ( .A(n6964), .ZN(n10163) );
  OAI222_X1 U8388 ( .A1(n8905), .A2(n6672), .B1(n9059), .B2(n6671), .C1(
        P2_U3151), .C2(n10163), .ZN(P2_U3291) );
  INV_X1 U8389 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6674) );
  INV_X1 U8390 ( .A(n7069), .ZN(n7073) );
  OAI222_X1 U8391 ( .A1(n8905), .A2(n6674), .B1(n9059), .B2(n6673), .C1(
        P2_U3151), .C2(n7073), .ZN(P2_U3290) );
  NAND2_X1 U8392 ( .A1(n6800), .A2(n6675), .ZN(n6683) );
  NAND2_X1 U8393 ( .A1(n6677), .A2(n6676), .ZN(n6679) );
  NAND2_X1 U8394 ( .A1(n6679), .A2(n6678), .ZN(n6681) );
  INV_X1 U8395 ( .A(n9995), .ZN(n9576) );
  NOR2_X1 U8396 ( .A1(n9576), .A2(P1_U3973), .ZN(P1_U3085) );
  NAND2_X1 U8397 ( .A1(n9376), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n6680) );
  OAI21_X1 U8398 ( .B1(n9625), .B2(n9376), .A(n6680), .ZN(P1_U3584) );
  INV_X1 U8399 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n6688) );
  INV_X1 U8400 ( .A(n6681), .ZN(n6682) );
  NAND2_X1 U8401 ( .A1(n6683), .A2(n6682), .ZN(n6821) );
  INV_X1 U8402 ( .A(n6821), .ZN(n6838) );
  INV_X1 U8403 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n8934) );
  INV_X1 U8404 ( .A(n8232), .ZN(n9390) );
  OR2_X1 U8405 ( .A1(n4281), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n6684) );
  NAND2_X1 U8406 ( .A1(n9390), .A2(n6684), .ZN(n9392) );
  AOI21_X1 U8407 ( .B1(n4281), .B2(n8934), .A(n9392), .ZN(n6685) );
  INV_X1 U8408 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n9391) );
  XNOR2_X1 U8409 ( .A(n6685), .B(n9391), .ZN(n6686) );
  AOI22_X1 U8410 ( .A1(n6838), .A2(n6686), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        P1_U3086), .ZN(n6687) );
  OAI21_X1 U8411 ( .B1(n9995), .B2(n6688), .A(n6687), .ZN(P1_U3243) );
  OAI222_X1 U8412 ( .A1(n6823), .A2(P1_U3086), .B1(n9963), .B2(n6690), .C1(
        n6689), .C2(n8253), .ZN(P1_U3354) );
  INV_X1 U8413 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6692) );
  INV_X1 U8414 ( .A(n6691), .ZN(n6693) );
  OAI222_X1 U8415 ( .A1(n8253), .A2(n6692), .B1(n9963), .B2(n6693), .C1(
        P1_U3086), .C2(n6832), .ZN(P1_U3348) );
  INV_X1 U8416 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6694) );
  OAI222_X1 U8417 ( .A1(n8905), .A2(n6694), .B1(n9059), .B2(n6693), .C1(
        P2_U3151), .C2(n7264), .ZN(P2_U3288) );
  INV_X1 U8418 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n6699) );
  INV_X1 U8419 ( .A(n6697), .ZN(n6698) );
  AOI22_X1 U8420 ( .A1(n6706), .A2(n6699), .B1(n6702), .B2(n6698), .ZN(
        P2_U3376) );
  INV_X1 U8421 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n8946) );
  INV_X1 U8422 ( .A(n6700), .ZN(n6701) );
  AOI22_X1 U8423 ( .A1(n6706), .A2(n8946), .B1(n6702), .B2(n6701), .ZN(
        P2_U3377) );
  AND2_X1 U8424 ( .A1(n6706), .A2(P2_D_REG_27__SCAN_IN), .ZN(P2_U3238) );
  AND2_X1 U8425 ( .A1(n6706), .A2(P2_D_REG_11__SCAN_IN), .ZN(P2_U3254) );
  AND2_X1 U8426 ( .A1(n6706), .A2(P2_D_REG_28__SCAN_IN), .ZN(P2_U3237) );
  AND2_X1 U8427 ( .A1(n6706), .A2(P2_D_REG_8__SCAN_IN), .ZN(P2_U3257) );
  AND2_X1 U8428 ( .A1(n6706), .A2(P2_D_REG_23__SCAN_IN), .ZN(P2_U3242) );
  AND2_X1 U8429 ( .A1(n6706), .A2(P2_D_REG_13__SCAN_IN), .ZN(P2_U3252) );
  AND2_X1 U8430 ( .A1(n6706), .A2(P2_D_REG_19__SCAN_IN), .ZN(P2_U3246) );
  AND2_X1 U8431 ( .A1(n6706), .A2(P2_D_REG_16__SCAN_IN), .ZN(P2_U3249) );
  AND2_X1 U8432 ( .A1(n6706), .A2(P2_D_REG_10__SCAN_IN), .ZN(P2_U3255) );
  AND2_X1 U8433 ( .A1(n6706), .A2(P2_D_REG_9__SCAN_IN), .ZN(P2_U3256) );
  AND2_X1 U8434 ( .A1(n6706), .A2(P2_D_REG_4__SCAN_IN), .ZN(P2_U3261) );
  AND2_X1 U8435 ( .A1(n6706), .A2(P2_D_REG_2__SCAN_IN), .ZN(P2_U3263) );
  AND2_X1 U8436 ( .A1(n6706), .A2(P2_D_REG_30__SCAN_IN), .ZN(P2_U3235) );
  AND2_X1 U8437 ( .A1(n6706), .A2(P2_D_REG_20__SCAN_IN), .ZN(P2_U3245) );
  AND2_X1 U8438 ( .A1(n6706), .A2(P2_D_REG_14__SCAN_IN), .ZN(P2_U3251) );
  AND2_X1 U8439 ( .A1(n6706), .A2(P2_D_REG_3__SCAN_IN), .ZN(P2_U3262) );
  AND2_X1 U8440 ( .A1(n6706), .A2(P2_D_REG_29__SCAN_IN), .ZN(P2_U3236) );
  AND2_X1 U8441 ( .A1(n6706), .A2(P2_D_REG_26__SCAN_IN), .ZN(P2_U3239) );
  AND2_X1 U8442 ( .A1(n6706), .A2(P2_D_REG_25__SCAN_IN), .ZN(P2_U3240) );
  AND2_X1 U8443 ( .A1(n6706), .A2(P2_D_REG_24__SCAN_IN), .ZN(P2_U3241) );
  AND2_X1 U8444 ( .A1(n6706), .A2(P2_D_REG_18__SCAN_IN), .ZN(P2_U3247) );
  AND2_X1 U8445 ( .A1(n6706), .A2(P2_D_REG_15__SCAN_IN), .ZN(P2_U3250) );
  AND2_X1 U8446 ( .A1(n6706), .A2(P2_D_REG_17__SCAN_IN), .ZN(P2_U3248) );
  AND2_X1 U8447 ( .A1(n6706), .A2(P2_D_REG_21__SCAN_IN), .ZN(P2_U3244) );
  INV_X1 U8448 ( .A(n6038), .ZN(n6704) );
  INV_X1 U8449 ( .A(n7305), .ZN(n7301) );
  OAI222_X1 U8450 ( .A1(n8905), .A2(n6703), .B1(n9059), .B2(n6704), .C1(
        P2_U3151), .C2(n7301), .ZN(P2_U3287) );
  INV_X1 U8451 ( .A(n9483), .ZN(n6817) );
  OAI222_X1 U8452 ( .A1(n8253), .A2(n6705), .B1(n9963), .B2(n6704), .C1(
        P1_U3086), .C2(n6817), .ZN(P1_U3347) );
  INV_X1 U8453 ( .A(P2_D_REG_22__SCAN_IN), .ZN(n9029) );
  NOR2_X1 U8454 ( .A1(n6707), .A2(n9029), .ZN(P2_U3243) );
  INV_X1 U8455 ( .A(P2_D_REG_12__SCAN_IN), .ZN(n9018) );
  NOR2_X1 U8456 ( .A1(n6707), .A2(n9018), .ZN(P2_U3253) );
  INV_X1 U8457 ( .A(P2_D_REG_31__SCAN_IN), .ZN(n8989) );
  NOR2_X1 U8458 ( .A1(n6707), .A2(n8989), .ZN(P2_U3234) );
  INV_X1 U8459 ( .A(P2_D_REG_7__SCAN_IN), .ZN(n8954) );
  NOR2_X1 U8460 ( .A1(n6707), .A2(n8954), .ZN(P2_U3258) );
  INV_X1 U8461 ( .A(P2_D_REG_5__SCAN_IN), .ZN(n9031) );
  NOR2_X1 U8462 ( .A1(n6707), .A2(n9031), .ZN(P2_U3260) );
  INV_X1 U8463 ( .A(P2_D_REG_6__SCAN_IN), .ZN(n9037) );
  NOR2_X1 U8464 ( .A1(n6707), .A2(n9037), .ZN(P2_U3259) );
  INV_X1 U8465 ( .A(n6708), .ZN(n6710) );
  INV_X1 U8466 ( .A(n7110), .ZN(n7104) );
  OAI222_X1 U8467 ( .A1(n8253), .A2(n6709), .B1(n9963), .B2(n6710), .C1(n7104), 
        .C2(P1_U3086), .ZN(P1_U3346) );
  OAI222_X1 U8468 ( .A1(n8905), .A2(n6711), .B1(n7406), .B2(P2_U3151), .C1(
        n9059), .C2(n6710), .ZN(P2_U3286) );
  INV_X1 U8469 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n6713) );
  INV_X1 U8470 ( .A(n6712), .ZN(n6714) );
  OAI222_X1 U8471 ( .A1(n8253), .A2(n6713), .B1(n9963), .B2(n6714), .C1(n7113), 
        .C2(P1_U3086), .ZN(P1_U3345) );
  INV_X1 U8472 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6715) );
  INV_X1 U8473 ( .A(n7540), .ZN(n7528) );
  OAI222_X1 U8474 ( .A1(n8905), .A2(n6715), .B1(n7528), .B2(P2_U3151), .C1(
        n9059), .C2(n6714), .ZN(P2_U3285) );
  INV_X1 U8475 ( .A(n6716), .ZN(n6717) );
  NAND2_X1 U8476 ( .A1(n6717), .A2(n6718), .ZN(n6730) );
  INV_X1 U8477 ( .A(n6718), .ZN(n7373) );
  OR2_X1 U8478 ( .A1(n7373), .A2(n8158), .ZN(n6719) );
  NAND2_X1 U8479 ( .A1(n6730), .A2(n6719), .ZN(n6725) );
  OR2_X1 U8480 ( .A1(n6725), .A2(n8005), .ZN(n6720) );
  NAND2_X1 U8481 ( .A1(n6720), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3150) );
  NOR2_X1 U8482 ( .A1(n8534), .A2(P2_U3151), .ZN(n6721) );
  NAND2_X1 U8483 ( .A1(n6721), .A2(n6726), .ZN(n6722) );
  OR2_X1 U8484 ( .A1(n6725), .A2(n6722), .ZN(n6724) );
  OR2_X1 U8485 ( .A1(n6726), .A2(P2_U3151), .ZN(n8910) );
  OR2_X1 U8486 ( .A1(n6730), .A2(n8910), .ZN(n6723) );
  NAND2_X1 U8487 ( .A1(P2_U3893), .A2(n6726), .ZN(n8570) );
  NOR2_X1 U8488 ( .A1(n6727), .A2(n6763), .ZN(n6756) );
  AOI21_X1 U8489 ( .B1(n6727), .B2(n6763), .A(n6756), .ZN(n6728) );
  AOI21_X1 U8490 ( .B1(n6760), .B2(n8570), .A(n6728), .ZN(n6729) );
  AOI21_X1 U8491 ( .B1(P2_REG3_REG_0__SCAN_IN), .B2(P2_U3151), .A(n6729), .ZN(
        n6733) );
  INV_X1 U8492 ( .A(P2_U3150), .ZN(n6731) );
  NAND2_X1 U8493 ( .A1(n10142), .A2(P2_ADDR_REG_0__SCAN_IN), .ZN(n6732) );
  OAI211_X1 U8494 ( .C1(n10164), .C2(n6763), .A(n6733), .B(n6732), .ZN(
        P2_U3182) );
  MUX2_X1 U8495 ( .A(n6734), .B(n8740), .S(P2_U3893), .Z(n6735) );
  INV_X1 U8496 ( .A(n6735), .ZN(P2_U3508) );
  INV_X1 U8497 ( .A(n6736), .ZN(n6738) );
  INV_X1 U8498 ( .A(n7700), .ZN(n7543) );
  OAI222_X1 U8499 ( .A1(n8905), .A2(n6737), .B1(n9059), .B2(n6738), .C1(
        P2_U3151), .C2(n7543), .ZN(P2_U3284) );
  INV_X1 U8500 ( .A(n9510), .ZN(n7106) );
  OAI222_X1 U8501 ( .A1(n8253), .A2(n6739), .B1(n9963), .B2(n6738), .C1(
        P1_U3086), .C2(n7106), .ZN(P1_U3344) );
  NAND2_X1 U8502 ( .A1(n4432), .A2(n10173), .ZN(n6938) );
  NAND2_X1 U8503 ( .A1(n6742), .A2(n10216), .ZN(n6740) );
  AND2_X1 U8504 ( .A1(n6938), .A2(n6740), .ZN(n6745) );
  OR2_X1 U8505 ( .A1(n6741), .A2(n6742), .ZN(n8020) );
  NAND2_X1 U8506 ( .A1(n8020), .A2(n8022), .ZN(n6937) );
  NAND2_X1 U8507 ( .A1(n10210), .A2(n8753), .ZN(n6743) );
  NAND2_X1 U8508 ( .A1(n6937), .A2(n6743), .ZN(n6744) );
  NAND2_X1 U8509 ( .A1(n6745), .A2(n6744), .ZN(n8818) );
  NAND2_X1 U8510 ( .A1(n10217), .A2(n8818), .ZN(n6746) );
  OAI21_X1 U8511 ( .B1(n10217), .B2(n5940), .A(n6746), .ZN(P2_U3390) );
  INV_X1 U8512 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n6750) );
  OAI21_X1 U8513 ( .B1(n10030), .B2(n10107), .A(n6979), .ZN(n6747) );
  NAND2_X1 U8514 ( .A1(n6849), .A2(n9304), .ZN(n6980) );
  OAI211_X1 U8515 ( .C1(n6991), .C2(n6748), .A(n6747), .B(n6980), .ZN(n9931)
         );
  NAND2_X1 U8516 ( .A1(n9931), .A2(n4272), .ZN(n6749) );
  OAI21_X1 U8517 ( .B1(n4272), .B2(n6750), .A(n6749), .ZN(P1_U3453) );
  INV_X1 U8518 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n6771) );
  NOR2_X2 U8519 ( .A1(n6760), .A2(n8564), .ZN(n10129) );
  NAND2_X1 U8520 ( .A1(n6763), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6751) );
  NAND2_X1 U8521 ( .A1(n6767), .A2(n6751), .ZN(n6753) );
  INV_X1 U8522 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n6752) );
  OR2_X1 U8523 ( .A1(n6764), .A2(n6752), .ZN(n6879) );
  AND2_X1 U8524 ( .A1(n6879), .A2(n6753), .ZN(n6754) );
  OAI21_X1 U8525 ( .B1(P2_REG1_REG_1__SCAN_IN), .B2(n6754), .A(n6880), .ZN(
        n6759) );
  INV_X1 U8526 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n6867) );
  NOR2_X1 U8527 ( .A1(n6867), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6758) );
  AOI211_X1 U8528 ( .C1(n6756), .C2(n6755), .A(n8570), .B(n6870), .ZN(n6757)
         );
  AOI211_X1 U8529 ( .C1(n10129), .C2(n6759), .A(n6758), .B(n6757), .ZN(n6770)
         );
  INV_X1 U8530 ( .A(n6760), .ZN(n6761) );
  OR2_X1 U8531 ( .A1(n6764), .A2(n6762), .ZN(n6876) );
  NAND2_X1 U8532 ( .A1(n6871), .A2(n6876), .ZN(n6766) );
  NAND3_X1 U8533 ( .A1(n6764), .A2(P2_REG2_REG_0__SCAN_IN), .A3(n6763), .ZN(
        n6765) );
  NAND2_X1 U8534 ( .A1(n6766), .A2(n6765), .ZN(n6875) );
  XNOR2_X1 U8535 ( .A(n6875), .B(P2_REG2_REG_1__SCAN_IN), .ZN(n6768) );
  AOI22_X1 U8536 ( .A1(n10160), .A2(n6768), .B1(n10125), .B2(n6767), .ZN(n6769) );
  OAI211_X1 U8537 ( .C1(n10170), .C2(n6771), .A(n6770), .B(n6769), .ZN(
        P2_U3183) );
  INV_X1 U8538 ( .A(n9952), .ZN(n6775) );
  NAND2_X1 U8539 ( .A1(n6772), .A2(P1_D_REG_1__SCAN_IN), .ZN(n6774) );
  INV_X1 U8540 ( .A(n9953), .ZN(n6773) );
  AOI21_X1 U8541 ( .B1(n6775), .B2(n6774), .A(n6773), .ZN(n6977) );
  NAND2_X1 U8542 ( .A1(n6776), .A2(n6977), .ZN(n6793) );
  NAND2_X1 U8543 ( .A1(n6793), .A2(n6799), .ZN(n6779) );
  AND2_X1 U8544 ( .A1(n6777), .A2(n6790), .ZN(n6778) );
  AOI21_X1 U8545 ( .B1(n6779), .B2(n6778), .A(P1_U3086), .ZN(n6780) );
  NAND2_X1 U8546 ( .A1(n9332), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6933) );
  INV_X1 U8547 ( .A(n6933), .ZN(n6806) );
  INV_X1 U8548 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n6982) );
  NAND2_X1 U8549 ( .A1(n9377), .A2(n4289), .ZN(n6789) );
  NAND2_X1 U8550 ( .A1(n6782), .A2(n6802), .ZN(n6784) );
  AND2_X1 U8551 ( .A1(n6785), .A2(n6790), .ZN(n6786) );
  NAND2_X2 U8552 ( .A1(n6787), .A2(n6786), .ZN(n7819) );
  NAND2_X1 U8553 ( .A1(n4287), .A2(n7819), .ZN(n7036) );
  NAND2_X1 U8554 ( .A1(n7036), .A2(n6986), .ZN(n6788) );
  NAND2_X1 U8555 ( .A1(n6789), .A2(n6788), .ZN(n6846) );
  INV_X1 U8556 ( .A(n6790), .ZN(n6791) );
  NOR2_X1 U8557 ( .A1(n6846), .A2(n4972), .ZN(n6792) );
  INV_X2 U8558 ( .A(n7056), .ZN(n7884) );
  AOI21_X1 U8559 ( .B1(n6792), .B2(n4307), .A(n6847), .ZN(n9397) );
  AND2_X1 U8560 ( .A1(n10103), .A2(n6794), .ZN(n6795) );
  NAND2_X1 U8561 ( .A1(n6797), .A2(n6796), .ZN(n6984) );
  INV_X1 U8562 ( .A(n6984), .ZN(n6798) );
  NAND2_X1 U8563 ( .A1(n6803), .A2(n6798), .ZN(n6801) );
  OAI22_X1 U8564 ( .A1(n9338), .A2(n6991), .B1(n9345), .B2(n6980), .ZN(n6804)
         );
  AOI21_X1 U8565 ( .B1(n9397), .B2(n9326), .A(n6804), .ZN(n6805) );
  OAI21_X1 U8566 ( .B1(n6806), .B2(n6982), .A(n6805), .ZN(P1_U3232) );
  XNOR2_X1 U8567 ( .A(n7110), .B(P1_REG2_REG_9__SCAN_IN), .ZN(n6819) );
  MUX2_X1 U8568 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n6808), .S(n9401), .Z(n9404)
         );
  AND2_X1 U8569 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n9394) );
  NAND2_X1 U8570 ( .A1(n9385), .A2(n9394), .ZN(n9384) );
  OAI21_X1 U8571 ( .B1(n5254), .B2(n6823), .A(n9384), .ZN(n9403) );
  NAND2_X1 U8572 ( .A1(n9404), .A2(n9403), .ZN(n9402) );
  OAI21_X1 U8573 ( .B1(n6808), .B2(n6807), .A(n9402), .ZN(n9416) );
  XOR2_X1 U8574 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n9414), .Z(n9417) );
  NAND2_X1 U8575 ( .A1(n9416), .A2(n9417), .ZN(n9415) );
  OAI21_X1 U8576 ( .B1(n6810), .B2(n6809), .A(n9415), .ZN(n9432) );
  MUX2_X1 U8577 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n7137), .S(n9427), .Z(n9433)
         );
  NAND2_X1 U8578 ( .A1(n9432), .A2(n9433), .ZN(n9431) );
  OAI21_X1 U8579 ( .B1(n6811), .B2(n7137), .A(n9431), .ZN(n9443) );
  XOR2_X1 U8580 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n9441), .Z(n9444) );
  NAND2_X1 U8581 ( .A1(n9443), .A2(n9444), .ZN(n9442) );
  MUX2_X1 U8582 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n7213), .S(n9454), .Z(n9460)
         );
  XNOR2_X1 U8583 ( .A(n6832), .B(P1_REG2_REG_7__SCAN_IN), .ZN(n9473) );
  OAI21_X1 U8584 ( .B1(n6815), .B2(n6832), .A(n9471), .ZN(n9479) );
  XOR2_X1 U8585 ( .A(n9483), .B(P1_REG2_REG_8__SCAN_IN), .Z(n9478) );
  NAND2_X1 U8586 ( .A1(n9479), .A2(n9478), .ZN(n9477) );
  OAI21_X1 U8587 ( .B1(n6817), .B2(n6816), .A(n9477), .ZN(n6818) );
  NOR2_X1 U8588 ( .A1(n6818), .A2(n6819), .ZN(n7103) );
  AOI21_X1 U8589 ( .B1(n6819), .B2(n6818), .A(n7103), .ZN(n6843) );
  INV_X1 U8590 ( .A(n9393), .ZN(n6820) );
  INV_X1 U8591 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n6822) );
  NAND2_X1 U8592 ( .A1(P1_U3086), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n9254) );
  OAI21_X1 U8593 ( .B1(n9995), .B2(n6822), .A(n9254), .ZN(n6841) );
  INV_X1 U8594 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n10109) );
  MUX2_X1 U8595 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n10109), .S(n9401), .Z(n9407)
         );
  XNOR2_X1 U8596 ( .A(n6823), .B(P1_REG1_REG_1__SCAN_IN), .ZN(n9383) );
  AND2_X1 U8597 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n9382) );
  NAND2_X1 U8598 ( .A1(n9383), .A2(n9382), .ZN(n9381) );
  NAND2_X1 U8599 ( .A1(n9380), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6824) );
  NAND2_X1 U8600 ( .A1(n9381), .A2(n6824), .ZN(n9406) );
  NAND2_X1 U8601 ( .A1(n9407), .A2(n9406), .ZN(n9405) );
  NAND2_X1 U8602 ( .A1(n9401), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6825) );
  NAND2_X1 U8603 ( .A1(n9405), .A2(n6825), .ZN(n9419) );
  INV_X1 U8604 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6826) );
  XNOR2_X1 U8605 ( .A(n9414), .B(n6826), .ZN(n9420) );
  NAND2_X1 U8606 ( .A1(n9419), .A2(n9420), .ZN(n9418) );
  NAND2_X1 U8607 ( .A1(n9414), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6827) );
  NAND2_X1 U8608 ( .A1(n9418), .A2(n6827), .ZN(n9429) );
  INV_X1 U8609 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n10112) );
  MUX2_X1 U8610 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n10112), .S(n9427), .Z(n9430)
         );
  NAND2_X1 U8611 ( .A1(n9429), .A2(n9430), .ZN(n9428) );
  NAND2_X1 U8612 ( .A1(n9427), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6828) );
  NAND2_X1 U8613 ( .A1(n9428), .A2(n6828), .ZN(n9446) );
  INV_X1 U8614 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n6829) );
  XNOR2_X1 U8615 ( .A(n9441), .B(n6829), .ZN(n9447) );
  NAND2_X1 U8616 ( .A1(n9446), .A2(n9447), .ZN(n9445) );
  NAND2_X1 U8617 ( .A1(n9441), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6830) );
  NAND2_X1 U8618 ( .A1(n9445), .A2(n6830), .ZN(n9456) );
  INV_X1 U8619 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n10116) );
  MUX2_X1 U8620 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n10116), .S(n9454), .Z(n9457)
         );
  NAND2_X1 U8621 ( .A1(n9456), .A2(n9457), .ZN(n9455) );
  NAND2_X1 U8622 ( .A1(n9454), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6831) );
  NAND2_X1 U8623 ( .A1(n9455), .A2(n6831), .ZN(n9469) );
  INV_X1 U8624 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n10118) );
  MUX2_X1 U8625 ( .A(n10118), .B(P1_REG1_REG_7__SCAN_IN), .S(n6832), .Z(n9470)
         );
  NAND2_X1 U8626 ( .A1(n9469), .A2(n9470), .ZN(n9468) );
  NAND2_X1 U8627 ( .A1(n9467), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6833) );
  NAND2_X1 U8628 ( .A1(n9468), .A2(n6833), .ZN(n9485) );
  INV_X1 U8629 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n6834) );
  XNOR2_X1 U8630 ( .A(n9483), .B(n6834), .ZN(n9486) );
  NAND2_X1 U8631 ( .A1(n9485), .A2(n9486), .ZN(n9484) );
  NAND2_X1 U8632 ( .A1(n9483), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6835) );
  NAND2_X1 U8633 ( .A1(n9484), .A2(n6835), .ZN(n6837) );
  INV_X1 U8634 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n10120) );
  MUX2_X1 U8635 ( .A(n10120), .B(P1_REG1_REG_9__SCAN_IN), .S(n7110), .Z(n6836)
         );
  OR2_X1 U8636 ( .A1(n6837), .A2(n6836), .ZN(n7112) );
  NAND2_X1 U8637 ( .A1(n6837), .A2(n6836), .ZN(n6839) );
  INV_X1 U8638 ( .A(n9966), .ZN(n9981) );
  AOI21_X1 U8639 ( .B1(n7112), .B2(n6839), .A(n9981), .ZN(n6840) );
  AOI211_X1 U8640 ( .C1(n4395), .C2(n7110), .A(n6841), .B(n6840), .ZN(n6842)
         );
  OAI21_X1 U8641 ( .B1(n6843), .B2(n9986), .A(n6842), .ZN(P1_U3252) );
  NOR2_X1 U8642 ( .A1(n8385), .A2(P2_U3151), .ZN(n7102) );
  INV_X1 U8643 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n6941) );
  INV_X1 U8644 ( .A(n6937), .ZN(n8176) );
  OAI22_X1 U8645 ( .A1(n8176), .A2(n8375), .B1(n8389), .B2(n6942), .ZN(n6844)
         );
  AOI21_X1 U8646 ( .B1(n8380), .B2(n4432), .A(n6844), .ZN(n6845) );
  OAI21_X1 U8647 ( .B1(n7102), .B2(n6941), .A(n6845), .ZN(P2_U3172) );
  INV_X1 U8648 ( .A(n6846), .ZN(n6848) );
  NAND2_X1 U8649 ( .A1(n6849), .A2(n4290), .ZN(n6850) );
  XNOR2_X1 U8650 ( .A(n6851), .B(n7819), .ZN(n6926) );
  OAI22_X1 U8651 ( .A1(n6853), .A2(n4288), .B1(n6992), .B2(n7056), .ZN(n6925)
         );
  XOR2_X1 U8652 ( .A(n6926), .B(n6925), .Z(n6929) );
  XOR2_X1 U8653 ( .A(n6930), .B(n6929), .Z(n6857) );
  AOI22_X1 U8654 ( .A1(n9375), .A2(n9304), .B1(n9305), .B2(n9377), .ZN(n6995)
         );
  OAI22_X1 U8655 ( .A1(n9338), .A2(n6992), .B1(n6995), .B2(n9345), .ZN(n6855)
         );
  AOI21_X1 U8656 ( .B1(P1_REG3_REG_1__SCAN_IN), .B2(n6933), .A(n6855), .ZN(
        n6856) );
  OAI21_X1 U8657 ( .B1(n6857), .B2(n9350), .A(n6856), .ZN(P1_U3222) );
  INV_X1 U8658 ( .A(n6858), .ZN(n6868) );
  INV_X1 U8659 ( .A(n9524), .ZN(n9518) );
  OAI222_X1 U8660 ( .A1(n8253), .A2(n6859), .B1(n9963), .B2(n6868), .C1(n9518), 
        .C2(P1_U3086), .ZN(P1_U3343) );
  OAI22_X1 U8661 ( .A1(n8389), .A2(n6517), .B1(n6741), .B2(n8382), .ZN(n6860)
         );
  AOI21_X1 U8662 ( .B1(n8380), .B2(n4882), .A(n6860), .ZN(n6866) );
  OAI21_X1 U8663 ( .B1(n6863), .B2(n6862), .A(n6861), .ZN(n6864) );
  NAND2_X1 U8664 ( .A1(n6864), .A2(n8367), .ZN(n6865) );
  OAI211_X1 U8665 ( .C1(n7102), .C2(n6867), .A(n6866), .B(n6865), .ZN(P2_U3162) );
  INV_X1 U8666 ( .A(n8412), .ZN(n7538) );
  OAI222_X1 U8667 ( .A1(n8905), .A2(n6869), .B1(n7538), .B2(P2_U3151), .C1(
        n9059), .C2(n6868), .ZN(P2_U3283) );
  AOI211_X1 U8668 ( .C1(n6874), .C2(n6873), .A(n8570), .B(n6953), .ZN(n6890)
         );
  INV_X1 U8669 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n6888) );
  INV_X1 U8670 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n9008) );
  XNOR2_X1 U8671 ( .A(n6959), .B(n9008), .ZN(n6946) );
  NAND2_X1 U8672 ( .A1(n6875), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n6877) );
  NAND2_X1 U8673 ( .A1(n6877), .A2(n6876), .ZN(n6945) );
  XNOR2_X1 U8674 ( .A(n6946), .B(n6945), .ZN(n6884) );
  INV_X1 U8675 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n6878) );
  XNOR2_X1 U8676 ( .A(n6959), .B(n6878), .ZN(n6882) );
  NAND2_X1 U8677 ( .A1(n6880), .A2(n6879), .ZN(n6881) );
  NAND2_X1 U8678 ( .A1(n6882), .A2(n6881), .ZN(n6961) );
  OAI21_X1 U8679 ( .B1(n6882), .B2(n6881), .A(n6961), .ZN(n6883) );
  AOI22_X1 U8680 ( .A1(n10160), .A2(n6884), .B1(n10129), .B2(n6883), .ZN(n6887) );
  INV_X1 U8681 ( .A(n4458), .ZN(n6885) );
  AOI22_X1 U8682 ( .A1(n10125), .A2(n6885), .B1(P2_U3151), .B2(
        P2_REG3_REG_2__SCAN_IN), .ZN(n6886) );
  OAI211_X1 U8683 ( .C1(n10170), .C2(n6888), .A(n6887), .B(n6886), .ZN(n6889)
         );
  OR2_X1 U8684 ( .A1(n6890), .A2(n6889), .ZN(P2_U3184) );
  INV_X1 U8685 ( .A(n6581), .ZN(n8023) );
  NAND2_X1 U8686 ( .A1(n6891), .A2(n8022), .ZN(n6892) );
  OAI21_X1 U8687 ( .B1(n6893), .B2(n8023), .A(n6892), .ZN(n6915) );
  INV_X1 U8688 ( .A(n6915), .ZN(n6913) );
  NAND2_X1 U8689 ( .A1(n6895), .A2(n6894), .ZN(n6896) );
  NAND2_X1 U8690 ( .A1(n6897), .A2(n6896), .ZN(n6899) );
  NOR2_X1 U8691 ( .A1(n6900), .A2(n5922), .ZN(n8748) );
  OR2_X1 U8692 ( .A1(n8756), .A2(n8748), .ZN(n6901) );
  OAI21_X1 U8693 ( .B1(n6891), .B2(n6903), .A(n6902), .ZN(n6906) );
  NAND2_X1 U8694 ( .A1(n4882), .A2(n10173), .ZN(n6904) );
  OAI21_X1 U8695 ( .B1(n6741), .B2(n8737), .A(n6904), .ZN(n6905) );
  AOI21_X1 U8696 ( .B1(n6906), .B2(n10178), .A(n6905), .ZN(n6916) );
  INV_X1 U8697 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n6907) );
  MUX2_X1 U8698 ( .A(n6916), .B(n6907), .S(n10187), .Z(n6912) );
  INV_X1 U8699 ( .A(n6908), .ZN(n6909) );
  INV_X1 U8700 ( .A(n8628), .ZN(n8757) );
  INV_X2 U8701 ( .A(n8655), .ZN(n10183) );
  AOI22_X1 U8702 ( .A1(n10181), .A2(n6910), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        n10183), .ZN(n6911) );
  OAI211_X1 U8703 ( .C1(n6913), .C2(n8747), .A(n6912), .B(n6911), .ZN(P2_U3232) );
  NOR2_X1 U8704 ( .A1(n6517), .A2(n8792), .ZN(n6914) );
  AOI21_X1 U8705 ( .B1(n6915), .B2(n10201), .A(n6914), .ZN(n6917) );
  AND2_X1 U8706 ( .A1(n6917), .A2(n6916), .ZN(n10188) );
  MUX2_X1 U8707 ( .A(n4438), .B(n10188), .S(n10229), .Z(n6918) );
  INV_X1 U8708 ( .A(n6918), .ZN(P2_U3460) );
  INV_X1 U8709 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6920) );
  INV_X1 U8710 ( .A(n6919), .ZN(n6921) );
  OAI222_X1 U8711 ( .A1(n8905), .A2(n6920), .B1(n9059), .B2(n6921), .C1(
        P2_U3151), .C2(n8419), .ZN(P2_U3282) );
  INV_X1 U8712 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n6922) );
  INV_X1 U8713 ( .A(n9541), .ZN(n9535) );
  OAI222_X1 U8714 ( .A1(n8253), .A2(n6922), .B1(n9963), .B2(n6921), .C1(
        P1_U3086), .C2(n9535), .ZN(P1_U3342) );
  OAI22_X1 U8715 ( .A1(n6852), .A2(n6854), .B1(n10060), .B2(n7056), .ZN(n7040)
         );
  INV_X1 U8716 ( .A(n6925), .ZN(n6928) );
  INV_X1 U8717 ( .A(n6926), .ZN(n6927) );
  AOI22_X1 U8718 ( .A1(n6930), .A2(n6929), .B1(n6928), .B2(n6927), .ZN(n7042)
         );
  AOI22_X1 U8719 ( .A1(n6931), .A2(n9304), .B1(n9305), .B2(n6849), .ZN(n10028)
         );
  OAI22_X1 U8720 ( .A1(n9338), .A2(n10060), .B1(n10028), .B2(n9345), .ZN(n6932) );
  AOI21_X1 U8721 ( .B1(P1_REG3_REG_2__SCAN_IN), .B2(n6933), .A(n6932), .ZN(
        n6934) );
  OAI21_X1 U8722 ( .B1(n6935), .B2(n9350), .A(n6934), .ZN(P1_U3237) );
  NAND3_X1 U8723 ( .A1(n6937), .A2(n6936), .A3(n8792), .ZN(n6939) );
  NAND2_X1 U8724 ( .A1(n6939), .A2(n6938), .ZN(n6940) );
  MUX2_X1 U8725 ( .A(n6940), .B(P2_REG2_REG_0__SCAN_IN), .S(n10187), .Z(n6944)
         );
  OAI22_X1 U8726 ( .A1(n8581), .A2(n6942), .B1(n6941), .B2(n8655), .ZN(n6943)
         );
  OR2_X1 U8727 ( .A1(n6944), .A2(n6943), .ZN(P2_U3233) );
  NAND2_X1 U8728 ( .A1(n6946), .A2(n6945), .ZN(n6948) );
  NAND2_X1 U8729 ( .A1(n6959), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6947) );
  NAND2_X1 U8730 ( .A1(n6948), .A2(n6947), .ZN(n6949) );
  NAND2_X1 U8731 ( .A1(n6949), .A2(n4270), .ZN(n6950) );
  MUX2_X1 U8732 ( .A(n6951), .B(P2_REG2_REG_4__SCAN_IN), .S(n6964), .Z(n10150)
         );
  OR2_X1 U8733 ( .A1(n6964), .A2(n6951), .ZN(n6952) );
  NAND2_X1 U8734 ( .A1(n10148), .A2(n6952), .ZN(n7074) );
  XNOR2_X1 U8735 ( .A(n7072), .B(n4532), .ZN(n6975) );
  MUX2_X1 U8736 ( .A(P2_REG2_REG_3__SCAN_IN), .B(P2_REG1_REG_3__SCAN_IN), .S(
        n8534), .Z(n6955) );
  XOR2_X1 U8737 ( .A(n4270), .B(n6955), .Z(n10140) );
  NAND2_X1 U8738 ( .A1(n10141), .A2(n10140), .ZN(n10139) );
  MUX2_X1 U8739 ( .A(P2_REG2_REG_4__SCAN_IN), .B(P2_REG1_REG_4__SCAN_IN), .S(
        n8534), .Z(n6956) );
  XNOR2_X1 U8740 ( .A(n6956), .B(n10163), .ZN(n10147) );
  INV_X1 U8741 ( .A(n6956), .ZN(n6957) );
  MUX2_X1 U8742 ( .A(P2_REG2_REG_5__SCAN_IN), .B(P2_REG1_REG_5__SCAN_IN), .S(
        n8534), .Z(n7066) );
  XNOR2_X1 U8743 ( .A(n7066), .B(n7069), .ZN(n6958) );
  AND2_X1 U8744 ( .A1(P2_U3151), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n7148) );
  AOI21_X1 U8745 ( .B1(n10125), .B2(n7069), .A(n7148), .ZN(n6971) );
  NAND2_X1 U8746 ( .A1(n6959), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6960) );
  NAND2_X1 U8747 ( .A1(n6961), .A2(n6960), .ZN(n6962) );
  OAI21_X1 U8748 ( .B1(n6962), .B2(n4270), .A(n10152), .ZN(n10126) );
  INV_X1 U8749 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n10221) );
  OR2_X2 U8750 ( .A1(n10126), .A2(n10221), .ZN(n10154) );
  NAND2_X1 U8751 ( .A1(n10154), .A2(n10152), .ZN(n6963) );
  XNOR2_X1 U8752 ( .A(n6964), .B(P2_REG1_REG_4__SCAN_IN), .ZN(n10151) );
  NAND2_X1 U8753 ( .A1(n6963), .A2(n10151), .ZN(n10157) );
  INV_X1 U8754 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n10223) );
  OR2_X1 U8755 ( .A1(n6964), .A2(n10223), .ZN(n6965) );
  OAI21_X1 U8756 ( .B1(n6966), .B2(n7073), .A(n7080), .ZN(n6967) );
  INV_X1 U8757 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n10225) );
  OR2_X2 U8758 ( .A1(n6967), .A2(n10225), .ZN(n7082) );
  NAND2_X1 U8759 ( .A1(n6967), .A2(n10225), .ZN(n6968) );
  NAND2_X1 U8760 ( .A1(n7082), .A2(n6968), .ZN(n6969) );
  NAND2_X1 U8761 ( .A1(n10129), .A2(n6969), .ZN(n6970) );
  OAI211_X1 U8762 ( .C1(n7649), .C2(n10170), .A(n6971), .B(n6970), .ZN(n6972)
         );
  INV_X1 U8763 ( .A(n6972), .ZN(n6973) );
  OAI211_X1 U8764 ( .C1(n6975), .C2(n10133), .A(n6974), .B(n6973), .ZN(
        P2_U3187) );
  NAND3_X1 U8765 ( .A1(n6977), .A2(n6976), .A3(n7000), .ZN(n6985) );
  NAND2_X1 U8766 ( .A1(n6979), .A2(n6978), .ZN(n6981) );
  OAI211_X1 U8767 ( .C1(n9806), .C2(n6982), .A(n6981), .B(n6980), .ZN(n6983)
         );
  NAND2_X1 U8768 ( .A1(n6983), .A2(n9996), .ZN(n6988) );
  NOR2_X2 U8769 ( .A1(n9768), .A2(n6984), .ZN(n10042) );
  AND2_X1 U8770 ( .A1(n9826), .A2(n10035), .ZN(n9752) );
  OAI21_X1 U8771 ( .B1(n10042), .B2(n9752), .A(n6986), .ZN(n6987) );
  OAI211_X1 U8772 ( .C1(n5270), .C2(n9996), .A(n6988), .B(n6987), .ZN(P1_U3293) );
  INV_X1 U8773 ( .A(n6989), .ZN(n10096) );
  XOR2_X1 U8774 ( .A(n6990), .B(n6994), .Z(n10048) );
  OAI211_X1 U8775 ( .C1(n6991), .C2(n6992), .A(n10035), .B(n10034), .ZN(n10044) );
  OAI21_X1 U8776 ( .B1(n6992), .B2(n10103), .A(n10044), .ZN(n6999) );
  INV_X1 U8777 ( .A(n7028), .ZN(n10005) );
  XOR2_X1 U8778 ( .A(n6994), .B(n6993), .Z(n6996) );
  OAI21_X1 U8779 ( .B1(n6996), .B2(n10000), .A(n6995), .ZN(n6997) );
  AOI21_X1 U8780 ( .B1(n10005), .B2(n10048), .A(n6997), .ZN(n10051) );
  INV_X1 U8781 ( .A(n10051), .ZN(n6998) );
  AOI211_X1 U8782 ( .C1(n10096), .C2(n10048), .A(n6999), .B(n6998), .ZN(n10058) );
  NAND2_X1 U8783 ( .A1(n10122), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n7002) );
  OAI21_X1 U8784 ( .B1(n10058), .B2(n10122), .A(n7002), .ZN(P1_U3523) );
  INV_X1 U8785 ( .A(n7003), .ZN(n7004) );
  AOI211_X1 U8786 ( .C1(n7006), .C2(n7005), .A(n8375), .B(n7004), .ZN(n7010)
         );
  INV_X1 U8787 ( .A(n8385), .ZN(n8260) );
  AOI22_X1 U8788 ( .A1(n8356), .A2(n4882), .B1(n8380), .B2(n8402), .ZN(n7008)
         );
  NOR2_X1 U8789 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5971), .ZN(n10134) );
  AOI21_X1 U8790 ( .B1(n8362), .B2(n10195), .A(n10134), .ZN(n7007) );
  OAI211_X1 U8791 ( .C1(P2_REG3_REG_3__SCAN_IN), .C2(n8260), .A(n7008), .B(
        n7007), .ZN(n7009) );
  OR2_X1 U8792 ( .A1(n7010), .A2(n7009), .ZN(P2_U3158) );
  INV_X1 U8793 ( .A(n7011), .ZN(n7012) );
  INV_X1 U8794 ( .A(n8467), .ZN(n8440) );
  OAI222_X1 U8795 ( .A1(n8905), .A2(n9000), .B1(n9059), .B2(n7012), .C1(
        P2_U3151), .C2(n8440), .ZN(P2_U3281) );
  INV_X1 U8796 ( .A(n9550), .ZN(n9563) );
  OAI222_X1 U8797 ( .A1(n8253), .A2(n7013), .B1(n9963), .B2(n7012), .C1(
        P1_U3086), .C2(n9563), .ZN(P1_U3341) );
  XNOR2_X1 U8798 ( .A(n7014), .B(n7016), .ZN(n10194) );
  XNOR2_X1 U8799 ( .A(n7015), .B(n7016), .ZN(n7019) );
  NAND2_X1 U8800 ( .A1(n4882), .A2(n10175), .ZN(n7017) );
  OAI21_X1 U8801 ( .B1(n7229), .B2(n8739), .A(n7017), .ZN(n7018) );
  AOI21_X1 U8802 ( .B1(n7019), .B2(n10178), .A(n7018), .ZN(n10198) );
  INV_X1 U8803 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n10130) );
  MUX2_X1 U8804 ( .A(n10198), .B(n10130), .S(n10187), .Z(n7021) );
  AOI22_X1 U8805 ( .A1(n10181), .A2(n10195), .B1(n5971), .B2(n10183), .ZN(
        n7020) );
  OAI211_X1 U8806 ( .C1(n8747), .C2(n10194), .A(n7021), .B(n7020), .ZN(
        P2_U3230) );
  XNOR2_X1 U8807 ( .A(n7027), .B(n5768), .ZN(n7025) );
  NOR2_X1 U8808 ( .A1(n9219), .A2(n9329), .ZN(n7023) );
  NOR2_X1 U8809 ( .A1(n6854), .A2(n9626), .ZN(n7022) );
  OR2_X1 U8810 ( .A1(n7023), .A2(n7022), .ZN(n7044) );
  INV_X1 U8811 ( .A(n7044), .ZN(n7024) );
  OAI21_X1 U8812 ( .B1(n7025), .B2(n10000), .A(n7024), .ZN(n10067) );
  INV_X1 U8813 ( .A(n10067), .ZN(n7035) );
  XNOR2_X1 U8814 ( .A(n7027), .B(n7026), .ZN(n10069) );
  NAND2_X1 U8815 ( .A1(n7028), .A2(n10008), .ZN(n10033) );
  INV_X1 U8816 ( .A(n9828), .ZN(n10024) );
  OAI211_X1 U8817 ( .C1(n7029), .C2(n10066), .A(n7030), .B(n10035), .ZN(n10065) );
  INV_X1 U8818 ( .A(n9826), .ZN(n9610) );
  NAND2_X1 U8819 ( .A1(n10042), .A2(n7043), .ZN(n7032) );
  AOI22_X1 U8820 ( .A1(n9768), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n10041), .B2(
        n5237), .ZN(n7031) );
  OAI211_X1 U8821 ( .C1(n10065), .C2(n9610), .A(n7032), .B(n7031), .ZN(n7033)
         );
  AOI21_X1 U8822 ( .B1(n10069), .B2(n10024), .A(n7033), .ZN(n7034) );
  OAI21_X1 U8823 ( .B1(n7035), .B2(n9768), .A(n7034), .ZN(P1_U3290) );
  AOI22_X1 U8824 ( .A1(n6931), .A2(n7884), .B1(n7043), .B2(n7904), .ZN(n7037)
         );
  XNOR2_X1 U8825 ( .A(n7037), .B(n4278), .ZN(n7052) );
  OAI22_X1 U8826 ( .A1(n7038), .A2(n4288), .B1(n10066), .B2(n7056), .ZN(n7050)
         );
  XNOR2_X1 U8827 ( .A(n7052), .B(n7050), .ZN(n7054) );
  INV_X1 U8828 ( .A(n7039), .ZN(n7041) );
  XOR2_X1 U8829 ( .A(n7055), .B(n7054), .Z(n7047) );
  AOI22_X1 U8830 ( .A1(n9335), .A2(n7044), .B1(n9348), .B2(n7043), .ZN(n7046)
         );
  MUX2_X1 U8831 ( .A(n9332), .B(P1_STATE_REG_SCAN_IN), .S(
        P1_REG3_REG_3__SCAN_IN), .Z(n7045) );
  OAI211_X1 U8832 ( .C1(n7047), .C2(n9350), .A(n7046), .B(n7045), .ZN(P1_U3218) );
  INV_X1 U8833 ( .A(n7048), .ZN(n7091) );
  INV_X1 U8834 ( .A(n9975), .ZN(n9553) );
  OAI222_X1 U8835 ( .A1(n8253), .A2(n7049), .B1(n9963), .B2(n7091), .C1(n9553), 
        .C2(P1_U3086), .ZN(P1_U3340) );
  INV_X1 U8836 ( .A(n7050), .ZN(n7051) );
  AOI22_X1 U8837 ( .A1(n9374), .A2(n7884), .B1(n10072), .B2(n7904), .ZN(n7057)
         );
  XNOR2_X1 U8838 ( .A(n7057), .B(n4278), .ZN(n7802) );
  OAI22_X1 U8839 ( .A1(n9219), .A2(n4288), .B1(n7141), .B2(n7056), .ZN(n7800)
         );
  XNOR2_X1 U8840 ( .A(n7802), .B(n7800), .ZN(n7058) );
  OAI211_X1 U8841 ( .C1(n7059), .C2(n7058), .A(n7801), .B(n9326), .ZN(n7065)
         );
  NAND2_X1 U8842 ( .A1(n9373), .A2(n9304), .ZN(n7061) );
  NAND2_X1 U8843 ( .A1(n6931), .A2(n9305), .ZN(n7060) );
  AND2_X1 U8844 ( .A1(n7061), .A2(n7060), .ZN(n7134) );
  NAND2_X1 U8845 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n9424) );
  NAND2_X1 U8846 ( .A1(n9348), .A2(n10072), .ZN(n7062) );
  OAI211_X1 U8847 ( .C1(n7134), .C2(n9345), .A(n9424), .B(n7062), .ZN(n7063)
         );
  AOI21_X1 U8848 ( .B1(n7139), .B2(n9343), .A(n7063), .ZN(n7064) );
  NAND2_X1 U8849 ( .A1(n7065), .A2(n7064), .ZN(P1_U3230) );
  MUX2_X1 U8850 ( .A(P2_REG2_REG_6__SCAN_IN), .B(P2_REG1_REG_6__SCAN_IN), .S(
        n8534), .Z(n7172) );
  XOR2_X1 U8851 ( .A(n7185), .B(n7172), .Z(n7071) );
  INV_X1 U8852 ( .A(n7066), .ZN(n7068) );
  AOI21_X1 U8853 ( .B1(n7071), .B2(n7070), .A(n7173), .ZN(n7090) );
  INV_X1 U8854 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n7259) );
  MUX2_X1 U8855 ( .A(n7259), .B(P2_REG2_REG_6__SCAN_IN), .S(n7185), .Z(n7077)
         );
  NAND2_X1 U8856 ( .A1(n7074), .A2(n7073), .ZN(n7075) );
  OAI21_X1 U8857 ( .B1(n7077), .B2(n7076), .A(n7187), .ZN(n7088) );
  NAND2_X1 U8858 ( .A1(n7082), .A2(n7080), .ZN(n7078) );
  XNOR2_X1 U8859 ( .A(n7185), .B(P2_REG1_REG_6__SCAN_IN), .ZN(n7079) );
  NAND2_X1 U8860 ( .A1(n7078), .A2(n7079), .ZN(n7180) );
  INV_X1 U8861 ( .A(n7079), .ZN(n7081) );
  NAND3_X1 U8862 ( .A1(n7082), .A2(n7081), .A3(n7080), .ZN(n7083) );
  INV_X1 U8863 ( .A(n10129), .ZN(n10155) );
  AOI21_X1 U8864 ( .B1(n7180), .B2(n7083), .A(n10155), .ZN(n7087) );
  NAND2_X1 U8865 ( .A1(n10142), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n7084) );
  NAND2_X1 U8866 ( .A1(P2_U3151), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n7199) );
  OAI211_X1 U8867 ( .C1(n10164), .C2(n7085), .A(n7084), .B(n7199), .ZN(n7086)
         );
  AOI211_X1 U8868 ( .C1(n10160), .C2(n7088), .A(n7087), .B(n7086), .ZN(n7089)
         );
  OAI21_X1 U8869 ( .B1(n7090), .B2(n8570), .A(n7089), .ZN(P2_U3188) );
  OAI222_X1 U8870 ( .A1(n8905), .A2(n7092), .B1(n4856), .B2(P2_U3151), .C1(
        n9059), .C2(n7091), .ZN(P2_U3280) );
  INV_X1 U8871 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n7101) );
  OAI22_X1 U8872 ( .A1(n8389), .A2(n7093), .B1(n6516), .B2(n8382), .ZN(n7094)
         );
  AOI21_X1 U8873 ( .B1(n8371), .B2(n10176), .A(n7094), .ZN(n7100) );
  OAI21_X1 U8874 ( .B1(n7097), .B2(n7095), .A(n7096), .ZN(n7098) );
  NAND2_X1 U8875 ( .A1(n7098), .A2(n8367), .ZN(n7099) );
  OAI211_X1 U8876 ( .C1(n7102), .C2(n7101), .A(n7100), .B(n7099), .ZN(P2_U3177) );
  XNOR2_X1 U8877 ( .A(n9524), .B(P1_REG2_REG_12__SCAN_IN), .ZN(n7109) );
  XNOR2_X1 U8878 ( .A(n7113), .B(P1_REG2_REG_10__SCAN_IN), .ZN(n9491) );
  XOR2_X1 U8879 ( .A(P1_REG2_REG_11__SCAN_IN), .B(n9510), .Z(n9505) );
  OAI21_X1 U8880 ( .B1(n7107), .B2(n7106), .A(n9504), .ZN(n7108) );
  NOR2_X1 U8881 ( .A1(n7108), .A2(n7109), .ZN(n9517) );
  AOI21_X1 U8882 ( .B1(n7109), .B2(n7108), .A(n9517), .ZN(n7124) );
  INV_X1 U8883 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n7664) );
  NAND2_X1 U8884 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n9185) );
  OAI21_X1 U8885 ( .B1(n9995), .B2(n7664), .A(n9185), .ZN(n7122) );
  OR2_X1 U8886 ( .A1(n7110), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n7111) );
  NAND2_X1 U8887 ( .A1(n7112), .A2(n7111), .ZN(n9498) );
  INV_X1 U8888 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n7114) );
  MUX2_X1 U8889 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n7114), .S(n7113), .Z(n9497)
         );
  OR2_X1 U8890 ( .A1(n9498), .A2(n9497), .ZN(n9499) );
  NAND2_X1 U8891 ( .A1(n9496), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n7115) );
  NAND2_X1 U8892 ( .A1(n9499), .A2(n7115), .ZN(n9513) );
  INV_X1 U8893 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n7116) );
  XNOR2_X1 U8894 ( .A(n9510), .B(n7116), .ZN(n9512) );
  NAND2_X1 U8895 ( .A1(n9513), .A2(n9512), .ZN(n9511) );
  NAND2_X1 U8896 ( .A1(n9510), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n7117) );
  NAND2_X1 U8897 ( .A1(n9511), .A2(n7117), .ZN(n7119) );
  XNOR2_X1 U8898 ( .A(n9524), .B(P1_REG1_REG_12__SCAN_IN), .ZN(n7118) );
  NAND2_X1 U8899 ( .A1(n7119), .A2(n7118), .ZN(n7120) );
  AOI21_X1 U8900 ( .B1(n9526), .B2(n7120), .A(n9981), .ZN(n7121) );
  AOI211_X1 U8901 ( .C1(n4395), .C2(n9524), .A(n7122), .B(n7121), .ZN(n7123)
         );
  OAI21_X1 U8902 ( .B1(n7124), .B2(n9986), .A(n7123), .ZN(P1_U3255) );
  INV_X1 U8903 ( .A(n7125), .ZN(n7166) );
  INV_X1 U8904 ( .A(n8253), .ZN(n9958) );
  AOI22_X1 U8905 ( .A1(n9578), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n9958), .ZN(n7126) );
  OAI21_X1 U8906 ( .B1(n7166), .B2(n9963), .A(n7126), .ZN(P1_U3339) );
  XNOR2_X1 U8907 ( .A(n7127), .B(n7128), .ZN(n10075) );
  NAND3_X1 U8908 ( .A1(n7131), .A2(n7130), .A3(n7129), .ZN(n7132) );
  AOI21_X1 U8909 ( .B1(n7133), .B2(n7132), .A(n10000), .ZN(n7136) );
  INV_X1 U8910 ( .A(n7134), .ZN(n7135) );
  NOR2_X1 U8911 ( .A1(n7136), .A2(n7135), .ZN(n10074) );
  MUX2_X1 U8912 ( .A(n7137), .B(n10074), .S(n9996), .Z(n7144) );
  INV_X1 U8913 ( .A(n7138), .ZN(n10022) );
  AOI211_X1 U8914 ( .C1(n10072), .C2(n7030), .A(n8236), .B(n10022), .ZN(n10071) );
  INV_X1 U8915 ( .A(n7139), .ZN(n7140) );
  OAI22_X1 U8916 ( .A1(n9816), .A2(n7141), .B1(n7140), .B2(n9806), .ZN(n7142)
         );
  AOI21_X1 U8917 ( .B1(n10071), .B2(n10046), .A(n7142), .ZN(n7143) );
  OAI211_X1 U8918 ( .C1(n10075), .C2(n9828), .A(n7144), .B(n7143), .ZN(
        P1_U3289) );
  OAI21_X1 U8919 ( .B1(n7147), .B2(n7146), .A(n7145), .ZN(n7152) );
  AOI22_X1 U8920 ( .A1(n8362), .A2(n10205), .B1(n8385), .B2(n7235), .ZN(n7150)
         );
  AOI21_X1 U8921 ( .B1(n8356), .B2(n8402), .A(n7148), .ZN(n7149) );
  OAI211_X1 U8922 ( .C1(n7230), .C2(n8360), .A(n7150), .B(n7149), .ZN(n7151)
         );
  AOI21_X1 U8923 ( .B1(n7152), .B2(n8367), .A(n7151), .ZN(n7153) );
  INV_X1 U8924 ( .A(n7153), .ZN(P2_U3167) );
  NAND2_X1 U8925 ( .A1(n9376), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n7154) );
  OAI21_X1 U8926 ( .B1(n9196), .B2(n9376), .A(n7154), .ZN(P1_U3580) );
  INV_X1 U8927 ( .A(n7155), .ZN(n7168) );
  AOI22_X1 U8928 ( .A1(n9592), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n9958), .ZN(n7156) );
  OAI21_X1 U8929 ( .B1(n7168), .B2(n9963), .A(n7156), .ZN(P1_U3338) );
  INV_X1 U8930 ( .A(n7157), .ZN(n7158) );
  AOI21_X1 U8931 ( .B1(n7160), .B2(n7159), .A(n7158), .ZN(n7165) );
  AOI22_X1 U8932 ( .A1(n8356), .A2(n10176), .B1(n8371), .B2(n10174), .ZN(n7161) );
  NAND2_X1 U8933 ( .A1(P2_U3151), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n10161) );
  OAI211_X1 U8934 ( .C1(n7162), .C2(n8389), .A(n7161), .B(n10161), .ZN(n7163)
         );
  AOI21_X1 U8935 ( .B1(n10184), .B2(n8385), .A(n7163), .ZN(n7164) );
  OAI21_X1 U8936 ( .B1(n7165), .B2(n8375), .A(n7164), .ZN(P2_U3170) );
  OAI222_X1 U8937 ( .A1(n8905), .A2(n7167), .B1(n8514), .B2(P2_U3151), .C1(
        n9059), .C2(n7166), .ZN(P2_U3279) );
  INV_X1 U8938 ( .A(n8533), .ZN(n8542) );
  OAI222_X1 U8939 ( .A1(n8905), .A2(n7169), .B1(n9059), .B2(n7168), .C1(
        P2_U3151), .C2(n8542), .ZN(P2_U3278) );
  NAND2_X1 U8940 ( .A1(n9376), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n7170) );
  OAI21_X1 U8941 ( .B1(n7171), .B2(n9376), .A(n7170), .ZN(P1_U3583) );
  INV_X1 U8942 ( .A(n7172), .ZN(n7174) );
  MUX2_X1 U8943 ( .A(P2_REG2_REG_7__SCAN_IN), .B(P2_REG1_REG_7__SCAN_IN), .S(
        n8534), .Z(n7268) );
  XOR2_X1 U8944 ( .A(n7271), .B(n7268), .Z(n7175) );
  AOI21_X1 U8945 ( .B1(n7176), .B2(n7175), .A(n7269), .ZN(n7191) );
  AND2_X1 U8946 ( .A1(P2_U3151), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n7287) );
  INV_X1 U8947 ( .A(n7287), .ZN(n7177) );
  OAI21_X1 U8948 ( .B1(n10164), .B2(n7264), .A(n7177), .ZN(n7184) );
  INV_X1 U8949 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n7178) );
  OR2_X1 U8950 ( .A1(n7185), .A2(n7178), .ZN(n7179) );
  INV_X1 U8951 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n7487) );
  AOI21_X1 U8952 ( .B1(n7276), .B2(n7182), .A(n10155), .ZN(n7183) );
  AOI211_X1 U8953 ( .C1(n10142), .C2(P2_ADDR_REG_7__SCAN_IN), .A(n7184), .B(
        n7183), .ZN(n7190) );
  OR2_X1 U8954 ( .A1(n7185), .A2(n7259), .ZN(n7186) );
  NAND2_X1 U8955 ( .A1(n7187), .A2(n7186), .ZN(n7265) );
  XNOR2_X1 U8956 ( .A(n7263), .B(P2_REG2_REG_7__SCAN_IN), .ZN(n7188) );
  NAND2_X1 U8957 ( .A1(n7188), .A2(n10160), .ZN(n7189) );
  OAI211_X1 U8958 ( .C1(n7191), .C2(n8570), .A(n7190), .B(n7189), .ZN(P2_U3189) );
  INV_X1 U8959 ( .A(n7192), .ZN(n7221) );
  AOI22_X1 U8960 ( .A1(n9991), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n9958), .ZN(n7193) );
  OAI21_X1 U8961 ( .B1(n7221), .B2(n9963), .A(n7193), .ZN(P1_U3337) );
  INV_X1 U8962 ( .A(n7194), .ZN(n7798) );
  OAI222_X1 U8963 ( .A1(n8905), .A2(n7195), .B1(n9059), .B2(n7798), .C1(
        P2_U3151), .C2(n8573), .ZN(P2_U3276) );
  OAI211_X1 U8964 ( .C1(n7198), .C2(n7197), .A(n7196), .B(n8367), .ZN(n7204)
         );
  NAND2_X1 U8965 ( .A1(n8380), .A2(n8400), .ZN(n7200) );
  OAI211_X1 U8966 ( .C1(n7201), .C2(n8382), .A(n7200), .B(n7199), .ZN(n7202)
         );
  AOI21_X1 U8967 ( .B1(n7260), .B2(n8385), .A(n7202), .ZN(n7203) );
  OAI211_X1 U8968 ( .C1(n4806), .C2(n8389), .A(n7204), .B(n7203), .ZN(P2_U3179) );
  XOR2_X1 U8969 ( .A(n7205), .B(n7207), .Z(n10087) );
  XOR2_X1 U8970 ( .A(n7207), .B(n7206), .Z(n7212) );
  NOR2_X1 U8971 ( .A1(n7208), .A2(n9329), .ZN(n7211) );
  NOR2_X1 U8972 ( .A1(n7209), .A2(n9626), .ZN(n7210) );
  OR2_X1 U8973 ( .A1(n7211), .A2(n7210), .ZN(n9316) );
  AOI21_X1 U8974 ( .B1(n7212), .B2(n10030), .A(n9316), .ZN(n10086) );
  MUX2_X1 U8975 ( .A(n7213), .B(n10086), .S(n9996), .Z(n7218) );
  AOI211_X1 U8976 ( .C1(n10083), .C2(n4392), .A(n8236), .B(n10010), .ZN(n10082) );
  INV_X1 U8977 ( .A(n9317), .ZN(n7214) );
  OAI22_X1 U8978 ( .A1(n9816), .A2(n7215), .B1(n9806), .B2(n7214), .ZN(n7216)
         );
  AOI21_X1 U8979 ( .B1(n10082), .B2(n10046), .A(n7216), .ZN(n7217) );
  OAI211_X1 U8980 ( .C1(n10087), .C2(n9828), .A(n7218), .B(n7217), .ZN(
        P1_U3287) );
  INV_X1 U8981 ( .A(n7219), .ZN(n7224) );
  OAI222_X1 U8982 ( .A1(n9059), .A2(n7224), .B1(n8215), .B2(P2_U3151), .C1(
        n7220), .C2(n8905), .ZN(P2_U3275) );
  OAI222_X1 U8983 ( .A1(n8905), .A2(n7222), .B1(n4523), .B2(P2_U3151), .C1(
        n9059), .C2(n7221), .ZN(P2_U3277) );
  OAI222_X1 U8984 ( .A1(n8253), .A2(n7225), .B1(n9963), .B2(n7224), .C1(n4469), 
        .C2(P1_U3086), .ZN(P1_U3335) );
  INV_X1 U8985 ( .A(n7226), .ZN(n7240) );
  OAI222_X1 U8986 ( .A1(n9059), .A2(n7240), .B1(n5922), .B2(P2_U3151), .C1(
        n8981), .C2(n8905), .ZN(P2_U3274) );
  XNOR2_X1 U8987 ( .A(n7228), .B(n10174), .ZN(n8178) );
  XOR2_X1 U8988 ( .A(n7227), .B(n8178), .Z(n10206) );
  INV_X1 U8989 ( .A(n10206), .ZN(n7238) );
  AND2_X1 U8990 ( .A1(n10186), .A2(n8748), .ZN(n8250) );
  OAI22_X1 U8991 ( .A1(n7230), .A2(n8739), .B1(n7229), .B2(n8737), .ZN(n7234)
         );
  XNOR2_X1 U8992 ( .A(n7231), .B(n8178), .ZN(n7232) );
  NOR2_X1 U8993 ( .A1(n7232), .A2(n8753), .ZN(n7233) );
  AOI211_X1 U8994 ( .C1(n8756), .C2(n10206), .A(n7234), .B(n7233), .ZN(n10208)
         );
  MUX2_X1 U8995 ( .A(n4532), .B(n10208), .S(n10186), .Z(n7237) );
  AOI22_X1 U8996 ( .A1(n10181), .A2(n10205), .B1(n10183), .B2(n7235), .ZN(
        n7236) );
  OAI211_X1 U8997 ( .C1(n7238), .C2(n7498), .A(n7237), .B(n7236), .ZN(P2_U3228) );
  OAI222_X1 U8998 ( .A1(n8253), .A2(n7241), .B1(n9963), .B2(n7240), .C1(n7239), 
        .C2(P1_U3086), .ZN(P1_U3334) );
  OR2_X1 U8999 ( .A1(n7206), .A2(n4662), .ZN(n7243) );
  NAND2_X1 U9000 ( .A1(n7243), .A2(n7242), .ZN(n9999) );
  OR2_X1 U9001 ( .A1(n9999), .A2(n9998), .ZN(n10002) );
  NAND2_X1 U9002 ( .A1(n10002), .A2(n7244), .ZN(n7321) );
  XNOR2_X1 U9003 ( .A(n7321), .B(n7319), .ZN(n7247) );
  NAND2_X1 U9004 ( .A1(n9369), .A2(n9304), .ZN(n7246) );
  NAND2_X1 U9005 ( .A1(n9371), .A2(n9305), .ZN(n7245) );
  AND2_X1 U9006 ( .A1(n7246), .A2(n7245), .ZN(n9155) );
  OAI21_X1 U9007 ( .B1(n7247), .B2(n10000), .A(n9155), .ZN(n7386) );
  INV_X1 U9008 ( .A(n7386), .ZN(n7254) );
  XNOR2_X1 U9009 ( .A(n7248), .B(n7319), .ZN(n7388) );
  XOR2_X1 U9010 ( .A(n10009), .B(n9157), .Z(n7249) );
  NAND2_X1 U9011 ( .A1(n7249), .A2(n10035), .ZN(n7384) );
  AOI22_X1 U9012 ( .A1(n9768), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n9153), .B2(
        n10041), .ZN(n7251) );
  NAND2_X1 U9013 ( .A1(n9157), .A2(n10042), .ZN(n7250) );
  OAI211_X1 U9014 ( .C1(n7384), .C2(n9610), .A(n7251), .B(n7250), .ZN(n7252)
         );
  AOI21_X1 U9015 ( .B1(n7388), .B2(n10024), .A(n7252), .ZN(n7253) );
  OAI21_X1 U9016 ( .B1(n7254), .B2(n9768), .A(n7253), .ZN(P1_U3285) );
  NAND2_X1 U9017 ( .A1(n7255), .A2(n8047), .ZN(n7256) );
  NAND2_X1 U9018 ( .A1(n8041), .A2(n8050), .ZN(n8179) );
  XNOR2_X1 U9019 ( .A(n7256), .B(n8179), .ZN(n10211) );
  XNOR2_X1 U9020 ( .A(n7257), .B(n8179), .ZN(n7258) );
  AOI222_X1 U9021 ( .A1(n10178), .A2(n7258), .B1(n8400), .B2(n10173), .C1(
        n10174), .C2(n10175), .ZN(n10212) );
  MUX2_X1 U9022 ( .A(n7259), .B(n10212), .S(n10186), .Z(n7262) );
  AOI22_X1 U9023 ( .A1(n10181), .A2(n10215), .B1(n10183), .B2(n7260), .ZN(
        n7261) );
  OAI211_X1 U9024 ( .C1(n8747), .C2(n10211), .A(n7262), .B(n7261), .ZN(
        P2_U3227) );
  XNOR2_X1 U9025 ( .A(n7305), .B(P2_REG2_REG_8__SCAN_IN), .ZN(n7298) );
  NAND2_X1 U9026 ( .A1(n7263), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n7267) );
  NAND2_X1 U9027 ( .A1(n7265), .A2(n7264), .ZN(n7266) );
  NAND2_X1 U9028 ( .A1(n7267), .A2(n7266), .ZN(n7299) );
  XOR2_X1 U9029 ( .A(n7299), .B(n7298), .Z(n7283) );
  INV_X1 U9030 ( .A(n7268), .ZN(n7270) );
  MUX2_X1 U9031 ( .A(P2_REG2_REG_8__SCAN_IN), .B(P2_REG1_REG_8__SCAN_IN), .S(
        n8534), .Z(n7302) );
  XOR2_X1 U9032 ( .A(n7305), .B(n7302), .Z(n7303) );
  XNOR2_X1 U9033 ( .A(n7304), .B(n7303), .ZN(n7281) );
  NAND2_X1 U9034 ( .A1(n7276), .A2(n7274), .ZN(n7272) );
  XNOR2_X1 U9035 ( .A(n7305), .B(P2_REG1_REG_8__SCAN_IN), .ZN(n7273) );
  INV_X1 U9036 ( .A(n7273), .ZN(n7275) );
  NAND3_X1 U9037 ( .A1(n7276), .A2(n7275), .A3(n7274), .ZN(n7277) );
  AOI21_X1 U9038 ( .B1(n7307), .B2(n7277), .A(n10155), .ZN(n7280) );
  NAND2_X1 U9039 ( .A1(n10142), .A2(P2_ADDR_REG_8__SCAN_IN), .ZN(n7278) );
  NAND2_X1 U9040 ( .A1(P2_U3151), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n7365) );
  OAI211_X1 U9041 ( .C1(n10164), .C2(n7301), .A(n7278), .B(n7365), .ZN(n7279)
         );
  AOI211_X1 U9042 ( .C1(n7281), .C2(n10166), .A(n7280), .B(n7279), .ZN(n7282)
         );
  OAI21_X1 U9043 ( .B1(n7283), .B2(n10133), .A(n7282), .ZN(P2_U3190) );
  INV_X1 U9044 ( .A(n7284), .ZN(n7361) );
  AOI21_X1 U9045 ( .B1(n7286), .B2(n7285), .A(n7361), .ZN(n7293) );
  AOI21_X1 U9046 ( .B1(n8356), .B2(n8401), .A(n7287), .ZN(n7291) );
  NAND2_X1 U9047 ( .A1(n8362), .A2(n7485), .ZN(n7290) );
  NAND2_X1 U9048 ( .A1(n8385), .A2(n7473), .ZN(n7289) );
  NAND2_X1 U9049 ( .A1(n8380), .A2(n8399), .ZN(n7288) );
  AND4_X1 U9050 ( .A1(n7291), .A2(n7290), .A3(n7289), .A4(n7288), .ZN(n7292)
         );
  OAI21_X1 U9051 ( .B1(n7293), .B2(n8375), .A(n7292), .ZN(P2_U3153) );
  INV_X1 U9052 ( .A(n7294), .ZN(n7296) );
  OAI222_X1 U9053 ( .A1(n8253), .A2(n9026), .B1(n9963), .B2(n7296), .C1(
        P1_U3086), .C2(n4452), .ZN(P1_U3333) );
  OAI222_X1 U9054 ( .A1(n8905), .A2(n7297), .B1(n9059), .B2(n7296), .C1(
        P2_U3151), .C2(n7295), .ZN(P2_U3273) );
  NAND2_X1 U9055 ( .A1(n7301), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n7300) );
  INV_X1 U9056 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n7732) );
  XNOR2_X1 U9057 ( .A(n7405), .B(n7732), .ZN(n7315) );
  MUX2_X1 U9058 ( .A(P2_REG2_REG_9__SCAN_IN), .B(P2_REG1_REG_9__SCAN_IN), .S(
        n8534), .Z(n7392) );
  XNOR2_X1 U9059 ( .A(n7392), .B(n7394), .ZN(n7395) );
  XNOR2_X1 U9060 ( .A(n7396), .B(n7395), .ZN(n7313) );
  INV_X1 U9061 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n9024) );
  OR2_X1 U9062 ( .A1(n7305), .A2(n9024), .ZN(n7306) );
  INV_X1 U9063 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n7756) );
  NAND2_X1 U9064 ( .A1(n7308), .A2(n7756), .ZN(n7309) );
  AOI21_X1 U9065 ( .B1(n7401), .B2(n7309), .A(n10155), .ZN(n7312) );
  NAND2_X1 U9066 ( .A1(n10142), .A2(P2_ADDR_REG_9__SCAN_IN), .ZN(n7310) );
  NAND2_X1 U9067 ( .A1(P2_U3151), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n8320) );
  OAI211_X1 U9068 ( .C1(n10164), .C2(n7406), .A(n7310), .B(n8320), .ZN(n7311)
         );
  AOI211_X1 U9069 ( .C1(n7313), .C2(n10166), .A(n7312), .B(n7311), .ZN(n7314)
         );
  OAI21_X1 U9070 ( .B1(n7315), .B2(n10133), .A(n7314), .ZN(P2_U3191) );
  INV_X1 U9071 ( .A(n7372), .ZN(n7318) );
  AOI21_X1 U9072 ( .B1(P2_DATAO_REG_23__SCAN_IN), .B2(n9958), .A(n7316), .ZN(
        n7317) );
  OAI21_X1 U9073 ( .B1(n7318), .B2(n9963), .A(n7317), .ZN(P1_U3332) );
  INV_X1 U9074 ( .A(n7319), .ZN(n7320) );
  NAND2_X1 U9075 ( .A1(n7321), .A2(n7320), .ZN(n7323) );
  NAND2_X1 U9076 ( .A1(n7323), .A2(n7322), .ZN(n7324) );
  XNOR2_X1 U9077 ( .A(n7324), .B(n7336), .ZN(n7325) );
  NAND2_X1 U9078 ( .A1(n7325), .A2(n10030), .ZN(n7333) );
  INV_X1 U9079 ( .A(n7351), .ZN(n7331) );
  AOI21_X1 U9080 ( .B1(n4986), .B2(n5388), .A(n8236), .ZN(n7330) );
  NAND2_X1 U9081 ( .A1(n6436), .A2(n9304), .ZN(n7328) );
  NAND2_X1 U9082 ( .A1(n9370), .A2(n9305), .ZN(n7327) );
  AND2_X1 U9083 ( .A1(n7328), .A2(n7327), .ZN(n9255) );
  INV_X1 U9084 ( .A(n9255), .ZN(n7329) );
  AOI21_X1 U9085 ( .B1(n7331), .B2(n7330), .A(n7329), .ZN(n7332) );
  NAND2_X1 U9086 ( .A1(n7333), .A2(n7332), .ZN(n10100) );
  NAND2_X1 U9087 ( .A1(n7333), .A2(n9630), .ZN(n7334) );
  AOI22_X1 U9088 ( .A1(n10100), .A2(n7334), .B1(n9257), .B2(n10041), .ZN(n7340) );
  XNOR2_X1 U9089 ( .A(n7335), .B(n7336), .ZN(n10097) );
  OAI22_X1 U9090 ( .A1(n4948), .A2(n9816), .B1(n7337), .B2(n9996), .ZN(n7338)
         );
  AOI21_X1 U9091 ( .B1(n10097), .B2(n10024), .A(n7338), .ZN(n7339) );
  OAI21_X1 U9092 ( .B1(n7340), .B2(n9768), .A(n7339), .ZN(P1_U3284) );
  XNOR2_X1 U9093 ( .A(n7341), .B(n7342), .ZN(n10106) );
  INV_X1 U9094 ( .A(n10106), .ZN(n7357) );
  AOI22_X1 U9095 ( .A1(n7841), .A2(n10042), .B1(n9768), .B2(
        P1_REG2_REG_10__SCAN_IN), .ZN(n7356) );
  OAI21_X1 U9096 ( .B1(n7344), .B2(n4390), .A(n7343), .ZN(n7348) );
  NAND2_X1 U9097 ( .A1(n9368), .A2(n9304), .ZN(n7346) );
  NAND2_X1 U9098 ( .A1(n9369), .A2(n9305), .ZN(n7345) );
  AND2_X1 U9099 ( .A1(n7346), .A2(n7345), .ZN(n9111) );
  INV_X1 U9100 ( .A(n9111), .ZN(n7347) );
  AOI21_X1 U9101 ( .B1(n7348), .B2(n10030), .A(n7347), .ZN(n10102) );
  INV_X1 U9102 ( .A(n10102), .ZN(n7354) );
  INV_X1 U9103 ( .A(n7349), .ZN(n7350) );
  OAI211_X1 U9104 ( .C1(n10104), .C2(n7351), .A(n7350), .B(n10035), .ZN(n10101) );
  INV_X1 U9105 ( .A(n9114), .ZN(n7352) );
  OAI22_X1 U9106 ( .A1(n10101), .A2(n9630), .B1(n9806), .B2(n7352), .ZN(n7353)
         );
  OAI21_X1 U9107 ( .B1(n7354), .B2(n7353), .A(n9996), .ZN(n7355) );
  OAI211_X1 U9108 ( .C1(n7357), .C2(n9828), .A(n7356), .B(n7355), .ZN(P1_U3283) );
  INV_X1 U9109 ( .A(n7465), .ZN(n7371) );
  INV_X1 U9110 ( .A(n7358), .ZN(n7360) );
  NOR3_X1 U9111 ( .A1(n7361), .A2(n7360), .A3(n7359), .ZN(n7364) );
  INV_X1 U9112 ( .A(n7362), .ZN(n7363) );
  OAI21_X1 U9113 ( .B1(n7364), .B2(n7363), .A(n8367), .ZN(n7370) );
  INV_X1 U9114 ( .A(n7365), .ZN(n7366) );
  AOI21_X1 U9115 ( .B1(n8356), .B2(n8400), .A(n7366), .ZN(n7367) );
  OAI21_X1 U9116 ( .B1(n7767), .B2(n8360), .A(n7367), .ZN(n7368) );
  AOI21_X1 U9117 ( .B1(n7458), .B2(n8385), .A(n7368), .ZN(n7369) );
  OAI211_X1 U9118 ( .C1(n7371), .C2(n8389), .A(n7370), .B(n7369), .ZN(P2_U3161) );
  NAND2_X1 U9119 ( .A1(n7372), .A2(n8908), .ZN(n7374) );
  NAND2_X1 U9120 ( .A1(n7373), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8231) );
  OAI211_X1 U9121 ( .C1(n7375), .C2(n8905), .A(n7374), .B(n8231), .ZN(P2_U3272) );
  INV_X1 U9122 ( .A(n7376), .ZN(n7378) );
  INV_X1 U9123 ( .A(n7449), .ZN(n7377) );
  AOI21_X1 U9124 ( .B1(n7378), .B2(n4901), .A(n7377), .ZN(n7469) );
  NOR2_X1 U9125 ( .A1(n7379), .A2(n8183), .ZN(n7453) );
  AOI21_X1 U9126 ( .B1(n8183), .B2(n7379), .A(n7453), .ZN(n7382) );
  AOI22_X1 U9127 ( .A1(n10175), .A2(n8401), .B1(n8399), .B2(n10173), .ZN(n7381) );
  NAND2_X1 U9128 ( .A1(n7469), .A2(n8756), .ZN(n7380) );
  OAI211_X1 U9129 ( .C1(n7382), .C2(n8753), .A(n7381), .B(n7380), .ZN(n7470)
         );
  AOI21_X1 U9130 ( .B1(n4391), .B2(n7469), .A(n7470), .ZN(n7486) );
  AOI22_X1 U9131 ( .A1(n8893), .A2(n7485), .B1(P2_REG0_REG_7__SCAN_IN), .B2(
        n10219), .ZN(n7383) );
  OAI21_X1 U9132 ( .B1(n7486), .B2(n10219), .A(n7383), .ZN(P2_U3411) );
  INV_X1 U9133 ( .A(n9157), .ZN(n7385) );
  OAI21_X1 U9134 ( .B1(n7385), .B2(n10103), .A(n7384), .ZN(n7387) );
  AOI211_X1 U9135 ( .C1(n10107), .C2(n7388), .A(n7387), .B(n7386), .ZN(n7391)
         );
  NAND2_X1 U9136 ( .A1(n10122), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n7389) );
  OAI21_X1 U9137 ( .B1(n7391), .B2(n10122), .A(n7389), .ZN(P1_U3530) );
  NAND2_X1 U9138 ( .A1(n10108), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n7390) );
  OAI21_X1 U9139 ( .B1(n7391), .B2(n10108), .A(n7390), .ZN(P1_U3477) );
  MUX2_X1 U9140 ( .A(P2_REG2_REG_10__SCAN_IN), .B(P2_REG1_REG_10__SCAN_IN), 
        .S(n8534), .Z(n7529) );
  XOR2_X1 U9141 ( .A(n7540), .B(n7529), .Z(n7530) );
  INV_X1 U9142 ( .A(n7392), .ZN(n7393) );
  XOR2_X1 U9143 ( .A(n7530), .B(n7531), .Z(n7415) );
  NAND2_X1 U9144 ( .A1(P2_U3151), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n7765) );
  OAI21_X1 U9145 ( .B1(n10164), .B2(n7528), .A(n7765), .ZN(n7404) );
  XNOR2_X1 U9146 ( .A(n7540), .B(P2_REG1_REG_10__SCAN_IN), .ZN(n7398) );
  NAND2_X1 U9147 ( .A1(n7397), .A2(n7398), .ZN(n7542) );
  INV_X1 U9148 ( .A(n7398), .ZN(n7400) );
  NAND3_X1 U9149 ( .A1(n7401), .A2(n7400), .A3(n7399), .ZN(n7402) );
  AOI21_X1 U9150 ( .B1(n7542), .B2(n7402), .A(n10155), .ZN(n7403) );
  AOI211_X1 U9151 ( .C1(n10142), .C2(P2_ADDR_REG_10__SCAN_IN), .A(n7404), .B(
        n7403), .ZN(n7414) );
  INV_X1 U9152 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7522) );
  MUX2_X1 U9153 ( .A(n7522), .B(P2_REG2_REG_10__SCAN_IN), .S(n7540), .Z(n7411)
         );
  NAND2_X1 U9154 ( .A1(n7407), .A2(n7406), .ZN(n7408) );
  NAND2_X1 U9155 ( .A1(n7409), .A2(n7408), .ZN(n7410) );
  OAI21_X1 U9156 ( .B1(n7411), .B2(n7410), .A(n7524), .ZN(n7412) );
  NAND2_X1 U9157 ( .A1(n7412), .A2(n10160), .ZN(n7413) );
  OAI211_X1 U9158 ( .C1(n7415), .C2(n8570), .A(n7414), .B(n7413), .ZN(P2_U3192) );
  XNOR2_X1 U9159 ( .A(n7416), .B(n4567), .ZN(n9930) );
  NAND3_X1 U9160 ( .A1(n7419), .A2(n7418), .A3(n7417), .ZN(n7420) );
  NAND3_X1 U9161 ( .A1(n7421), .A2(n10030), .A3(n7420), .ZN(n7424) );
  NAND2_X1 U9162 ( .A1(n9366), .A2(n9304), .ZN(n7423) );
  NAND2_X1 U9163 ( .A1(n9368), .A2(n9305), .ZN(n7422) );
  AND2_X1 U9164 ( .A1(n7423), .A2(n7422), .ZN(n9186) );
  NAND2_X1 U9165 ( .A1(n7424), .A2(n9186), .ZN(n9927) );
  INV_X1 U9166 ( .A(n7505), .ZN(n7426) );
  AOI211_X1 U9167 ( .C1(n9928), .C2(n7425), .A(n8236), .B(n7426), .ZN(n9926)
         );
  NAND2_X1 U9168 ( .A1(n9926), .A2(n10046), .ZN(n7428) );
  AOI22_X1 U9169 ( .A1(n9768), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n9188), .B2(
        n10041), .ZN(n7427) );
  OAI211_X1 U9170 ( .C1(n9191), .C2(n9816), .A(n7428), .B(n7427), .ZN(n7429)
         );
  AOI21_X1 U9171 ( .B1(n9996), .B2(n9927), .A(n7429), .ZN(n7430) );
  OAI21_X1 U9172 ( .B1(n9930), .B2(n9828), .A(n7430), .ZN(P1_U3281) );
  NAND2_X1 U9173 ( .A1(n8403), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n7431) );
  OAI21_X1 U9174 ( .B1(n8017), .B2(n8403), .A(n7431), .ZN(P2_U3521) );
  INV_X1 U9175 ( .A(n7432), .ZN(n7446) );
  OAI222_X1 U9176 ( .A1(n9059), .A2(n7446), .B1(P2_U3151), .B2(n7434), .C1(
        n7433), .C2(n8905), .ZN(P2_U3271) );
  NAND2_X1 U9177 ( .A1(n7343), .A2(n7435), .ZN(n7436) );
  XOR2_X1 U9178 ( .A(n7438), .B(n7436), .Z(n7437) );
  AOI22_X1 U9179 ( .A1(n6436), .A2(n9305), .B1(n9304), .B2(n9367), .ZN(n9297)
         );
  OAI21_X1 U9180 ( .B1(n7437), .B2(n10000), .A(n9297), .ZN(n7479) );
  INV_X1 U9181 ( .A(n7479), .ZN(n7444) );
  XNOR2_X1 U9182 ( .A(n7439), .B(n7438), .ZN(n7481) );
  OAI211_X1 U9183 ( .C1(n7349), .C2(n7478), .A(n10035), .B(n7425), .ZN(n7477)
         );
  AOI22_X1 U9184 ( .A1(n9768), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n9295), .B2(
        n10041), .ZN(n7441) );
  NAND2_X1 U9185 ( .A1(n9299), .A2(n10042), .ZN(n7440) );
  OAI211_X1 U9186 ( .C1(n7477), .C2(n9610), .A(n7441), .B(n7440), .ZN(n7442)
         );
  AOI21_X1 U9187 ( .B1(n7481), .B2(n10024), .A(n7442), .ZN(n7443) );
  OAI21_X1 U9188 ( .B1(n9768), .B2(n7444), .A(n7443), .ZN(P1_U3282) );
  OAI222_X1 U9189 ( .A1(P1_U3086), .A2(n7447), .B1(n9963), .B2(n7446), .C1(
        n7445), .C2(n8253), .ZN(P1_U3331) );
  NAND2_X1 U9190 ( .A1(n7449), .A2(n7448), .ZN(n7450) );
  XNOR2_X1 U9191 ( .A(n7450), .B(n8182), .ZN(n7468) );
  OAI21_X1 U9192 ( .B1(n7453), .B2(n7451), .A(n8182), .ZN(n7454) );
  OR2_X1 U9193 ( .A1(n7453), .A2(n7452), .ZN(n7728) );
  NAND3_X1 U9194 ( .A1(n7454), .A2(n10178), .A3(n7728), .ZN(n7456) );
  AOI22_X1 U9195 ( .A1(n8400), .A2(n10175), .B1(n10173), .B2(n8398), .ZN(n7455) );
  INV_X1 U9196 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7457) );
  MUX2_X1 U9197 ( .A(n7464), .B(n7457), .S(n10187), .Z(n7460) );
  AOI22_X1 U9198 ( .A1(n10181), .A2(n7465), .B1(n10183), .B2(n7458), .ZN(n7459) );
  OAI211_X1 U9199 ( .C1(n7468), .C2(n8747), .A(n7460), .B(n7459), .ZN(P2_U3225) );
  MUX2_X1 U9200 ( .A(n7464), .B(n9024), .S(n10227), .Z(n7462) );
  NAND2_X1 U9201 ( .A1(n8810), .A2(n7465), .ZN(n7461) );
  OAI211_X1 U9202 ( .C1(n7468), .C2(n8813), .A(n7462), .B(n7461), .ZN(P2_U3467) );
  INV_X1 U9203 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n7463) );
  MUX2_X1 U9204 ( .A(n7464), .B(n7463), .S(n10219), .Z(n7467) );
  NAND2_X1 U9205 ( .A1(n8893), .A2(n7465), .ZN(n7466) );
  OAI211_X1 U9206 ( .C1(n7468), .C2(n8896), .A(n7467), .B(n7466), .ZN(P2_U3414) );
  INV_X1 U9207 ( .A(n7469), .ZN(n7476) );
  INV_X1 U9208 ( .A(n7470), .ZN(n7471) );
  MUX2_X1 U9209 ( .A(n7472), .B(n7471), .S(n10186), .Z(n7475) );
  AOI22_X1 U9210 ( .A1(n10181), .A2(n7485), .B1(n10183), .B2(n7473), .ZN(n7474) );
  OAI211_X1 U9211 ( .C1(n7476), .C2(n7498), .A(n7475), .B(n7474), .ZN(P2_U3226) );
  OAI21_X1 U9212 ( .B1(n7478), .B2(n10103), .A(n7477), .ZN(n7480) );
  AOI211_X1 U9213 ( .C1(n7481), .C2(n10107), .A(n7480), .B(n7479), .ZN(n7484)
         );
  NAND2_X1 U9214 ( .A1(n10108), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n7482) );
  OAI21_X1 U9215 ( .B1(n7484), .B2(n10108), .A(n7482), .ZN(P1_U3486) );
  NAND2_X1 U9216 ( .A1(n10122), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n7483) );
  OAI21_X1 U9217 ( .B1(n7484), .B2(n10122), .A(n7483), .ZN(P1_U3533) );
  INV_X1 U9218 ( .A(n7485), .ZN(n7489) );
  MUX2_X1 U9219 ( .A(n7487), .B(n7486), .S(n10229), .Z(n7488) );
  OAI21_X1 U9220 ( .B1(n7489), .B2(n8780), .A(n7488), .ZN(P2_U3466) );
  INV_X1 U9221 ( .A(n8184), .ZN(n7491) );
  OAI21_X1 U9222 ( .B1(n7490), .B2(n7491), .A(n8057), .ZN(n7588) );
  XNOR2_X1 U9223 ( .A(n7588), .B(n8186), .ZN(n7514) );
  INV_X1 U9224 ( .A(n7514), .ZN(n7499) );
  XNOR2_X1 U9225 ( .A(n7591), .B(n8186), .ZN(n7494) );
  OAI22_X1 U9226 ( .A1(n7767), .A2(n8737), .B1(n7565), .B2(n8739), .ZN(n7492)
         );
  AOI21_X1 U9227 ( .B1(n7514), .B2(n8756), .A(n7492), .ZN(n7493) );
  OAI21_X1 U9228 ( .B1(n8753), .B2(n7494), .A(n7493), .ZN(n7513) );
  INV_X1 U9229 ( .A(n7513), .ZN(n7495) );
  MUX2_X1 U9230 ( .A(n7522), .B(n7495), .S(n10186), .Z(n7497) );
  AOI22_X1 U9231 ( .A1(n7770), .A2(n10181), .B1(n10183), .B2(n7769), .ZN(n7496) );
  OAI211_X1 U9232 ( .C1(n7499), .C2(n7498), .A(n7497), .B(n7496), .ZN(P2_U3223) );
  XNOR2_X1 U9233 ( .A(n7500), .B(n7503), .ZN(n7502) );
  AOI22_X1 U9234 ( .A1(n9305), .A2(n9367), .B1(n9365), .B2(n9304), .ZN(n9276)
         );
  INV_X1 U9235 ( .A(n9276), .ZN(n7501) );
  AOI21_X1 U9236 ( .B1(n7502), .B2(n10030), .A(n7501), .ZN(n9924) );
  XNOR2_X1 U9237 ( .A(n7504), .B(n7503), .ZN(n9925) );
  INV_X1 U9238 ( .A(n9925), .ZN(n7511) );
  INV_X1 U9239 ( .A(n9922), .ZN(n9281) );
  NAND2_X1 U9240 ( .A1(n9922), .A2(n7505), .ZN(n7506) );
  NAND2_X1 U9241 ( .A1(n7506), .A2(n10035), .ZN(n7507) );
  NOR2_X1 U9242 ( .A1(n7578), .A2(n7507), .ZN(n9921) );
  NAND2_X1 U9243 ( .A1(n9921), .A2(n10046), .ZN(n7509) );
  AOI22_X1 U9244 ( .A1(n9768), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n9278), .B2(
        n10041), .ZN(n7508) );
  OAI211_X1 U9245 ( .C1(n9281), .C2(n9816), .A(n7509), .B(n7508), .ZN(n7510)
         );
  AOI21_X1 U9246 ( .B1(n7511), .B2(n10024), .A(n7510), .ZN(n7512) );
  OAI21_X1 U9247 ( .B1(n9768), .B2(n9924), .A(n7512), .ZN(P1_U3280) );
  INV_X1 U9248 ( .A(n7770), .ZN(n7519) );
  INV_X1 U9249 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n7539) );
  AOI21_X1 U9250 ( .B1(n4391), .B2(n7514), .A(n7513), .ZN(n7516) );
  MUX2_X1 U9251 ( .A(n7539), .B(n7516), .S(n10229), .Z(n7515) );
  OAI21_X1 U9252 ( .B1(n7519), .B2(n8780), .A(n7515), .ZN(P2_U3469) );
  INV_X1 U9253 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n7517) );
  MUX2_X1 U9254 ( .A(n7517), .B(n7516), .S(n10217), .Z(n7518) );
  OAI21_X1 U9255 ( .B1(n7519), .B2(n8845), .A(n7518), .ZN(P2_U3420) );
  INV_X1 U9256 ( .A(n7520), .ZN(n7556) );
  OAI222_X1 U9257 ( .A1(n9059), .A2(n7556), .B1(P2_U3151), .B2(n7521), .C1(
        n8983), .C2(n8905), .ZN(P2_U3270) );
  XNOR2_X1 U9258 ( .A(n8412), .B(P2_REG2_REG_12__SCAN_IN), .ZN(n8405) );
  OR2_X1 U9259 ( .A1(n7540), .A2(n7522), .ZN(n7523) );
  NAND2_X1 U9260 ( .A1(n7525), .A2(n7543), .ZN(n7526) );
  NAND2_X1 U9261 ( .A1(n7527), .A2(n7526), .ZN(n8406) );
  XOR2_X1 U9262 ( .A(n8405), .B(n8406), .Z(n7554) );
  MUX2_X1 U9263 ( .A(P2_REG2_REG_11__SCAN_IN), .B(P2_REG1_REG_11__SCAN_IN), 
        .S(n8534), .Z(n7532) );
  XNOR2_X1 U9264 ( .A(n7532), .B(n7700), .ZN(n7703) );
  INV_X1 U9265 ( .A(n7532), .ZN(n7533) );
  INV_X1 U9266 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n8411) );
  MUX2_X1 U9267 ( .A(n8407), .B(n8411), .S(n8534), .Z(n7535) );
  INV_X1 U9268 ( .A(n7535), .ZN(n7534) );
  NAND2_X1 U9269 ( .A1(n7534), .A2(n7538), .ZN(n8422) );
  NAND2_X1 U9270 ( .A1(n7535), .A2(n8412), .ZN(n8417) );
  NAND2_X1 U9271 ( .A1(n8422), .A2(n8417), .ZN(n7536) );
  XNOR2_X1 U9272 ( .A(n8418), .B(n7536), .ZN(n7537) );
  NAND2_X1 U9273 ( .A1(n7537), .A2(n10166), .ZN(n7553) );
  NAND2_X1 U9274 ( .A1(P2_U3151), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n7563) );
  OAI21_X1 U9275 ( .B1(n10164), .B2(n7538), .A(n7563), .ZN(n7551) );
  OR2_X1 U9276 ( .A1(n7540), .A2(n7539), .ZN(n7541) );
  XNOR2_X1 U9277 ( .A(n8412), .B(P2_REG1_REG_12__SCAN_IN), .ZN(n7546) );
  NAND2_X1 U9278 ( .A1(n7545), .A2(n7546), .ZN(n8414) );
  INV_X1 U9279 ( .A(n7546), .ZN(n7548) );
  NAND3_X1 U9280 ( .A1(n7698), .A2(n7548), .A3(n7547), .ZN(n7549) );
  AOI21_X1 U9281 ( .B1(n8414), .B2(n7549), .A(n10155), .ZN(n7550) );
  AOI211_X1 U9282 ( .C1(n10142), .C2(P2_ADDR_REG_12__SCAN_IN), .A(n7551), .B(
        n7550), .ZN(n7552) );
  OAI211_X1 U9283 ( .C1(n7554), .C2(n10133), .A(n7553), .B(n7552), .ZN(
        P2_U3194) );
  OAI222_X1 U9284 ( .A1(P1_U3086), .A2(n7557), .B1(n9963), .B2(n7556), .C1(
        n7555), .C2(n8253), .ZN(P1_U3330) );
  NAND2_X1 U9285 ( .A1(n7559), .A2(n7558), .ZN(n7562) );
  XOR2_X1 U9286 ( .A(n7562), .B(n7561), .Z(n7569) );
  NAND2_X1 U9287 ( .A1(n8380), .A2(n8394), .ZN(n7564) );
  OAI211_X1 U9288 ( .C1(n7565), .C2(n8382), .A(n7564), .B(n7563), .ZN(n7566)
         );
  AOI21_X1 U9289 ( .B1(n7632), .B2(n8385), .A(n7566), .ZN(n7568) );
  NAND2_X1 U9290 ( .A1(n7636), .A2(n8362), .ZN(n7567) );
  OAI211_X1 U9291 ( .C1(n7569), .C2(n8375), .A(n7568), .B(n7567), .ZN(P2_U3164) );
  XOR2_X1 U9292 ( .A(n7572), .B(n7570), .Z(n9920) );
  INV_X1 U9293 ( .A(n7571), .ZN(n7574) );
  OAI21_X1 U9294 ( .B1(n7574), .B2(n7573), .A(n7572), .ZN(n7576) );
  NAND3_X1 U9295 ( .A1(n7576), .A2(n10030), .A3(n7575), .ZN(n7577) );
  AOI22_X1 U9296 ( .A1(n9366), .A2(n9305), .B1(n9304), .B2(n9364), .ZN(n9082)
         );
  NAND2_X1 U9297 ( .A1(n7577), .A2(n9082), .ZN(n9917) );
  INV_X1 U9298 ( .A(n7578), .ZN(n7579) );
  AOI211_X1 U9299 ( .C1(n5461), .C2(n7579), .A(n8236), .B(n7744), .ZN(n9918)
         );
  NAND2_X1 U9300 ( .A1(n9918), .A2(n9826), .ZN(n7581) );
  AOI22_X1 U9301 ( .A1(n9768), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n9086), .B2(
        n10041), .ZN(n7580) );
  OAI211_X1 U9302 ( .C1(n9083), .C2(n9816), .A(n7581), .B(n7580), .ZN(n7582)
         );
  AOI21_X1 U9303 ( .B1(n9996), .B2(n9917), .A(n7582), .ZN(n7583) );
  OAI21_X1 U9304 ( .B1(n9920), .B2(n9828), .A(n7583), .ZN(P1_U3279) );
  INV_X1 U9305 ( .A(n7584), .ZN(n7684) );
  OAI222_X1 U9306 ( .A1(P1_U3086), .A2(n7586), .B1(n9963), .B2(n7684), .C1(
        n7585), .C2(n8253), .ZN(P1_U3329) );
  INV_X1 U9307 ( .A(n8079), .ZN(n7587) );
  NAND2_X1 U9308 ( .A1(n7770), .A2(n7782), .ZN(n8076) );
  OAI21_X1 U9309 ( .B1(n7588), .B2(n7587), .A(n8076), .ZN(n7589) );
  XNOR2_X1 U9310 ( .A(n7589), .B(n8187), .ZN(n7610) );
  NAND2_X1 U9311 ( .A1(n7591), .A2(n7590), .ZN(n7613) );
  NAND2_X1 U9312 ( .A1(n7613), .A2(n7592), .ZN(n7593) );
  XOR2_X1 U9313 ( .A(n8187), .B(n7593), .Z(n7594) );
  AOI222_X1 U9314 ( .A1(n10178), .A2(n7594), .B1(n8397), .B2(n10175), .C1(
        n8395), .C2(n10173), .ZN(n7606) );
  MUX2_X1 U9315 ( .A(n7595), .B(n7606), .S(n10217), .Z(n7597) );
  NAND2_X1 U9316 ( .A1(n6536), .A2(n8893), .ZN(n7596) );
  OAI211_X1 U9317 ( .C1(n7610), .C2(n8896), .A(n7597), .B(n7596), .ZN(P2_U3423) );
  XNOR2_X1 U9318 ( .A(n7598), .B(n8096), .ZN(n7599) );
  AOI222_X1 U9319 ( .A1(n10178), .A2(n7599), .B1(n8395), .B2(n10175), .C1(
        n8393), .C2(n10173), .ZN(n7690) );
  AOI22_X1 U9320 ( .A1(n8093), .A2(n8757), .B1(n10183), .B2(n7628), .ZN(n7600)
         );
  AOI21_X1 U9321 ( .B1(n7690), .B2(n7600), .A(n10187), .ZN(n7603) );
  INV_X1 U9322 ( .A(n8096), .ZN(n8189) );
  XNOR2_X1 U9323 ( .A(n7601), .B(n8189), .ZN(n7693) );
  OAI22_X1 U9324 ( .A1(n7693), .A2(n8747), .B1(n8410), .B2(n10186), .ZN(n7602)
         );
  OR2_X1 U9325 ( .A1(n7603), .A2(n7602), .ZN(P2_U3220) );
  MUX2_X1 U9326 ( .A(n7696), .B(n7606), .S(n10186), .Z(n7605) );
  AOI22_X1 U9327 ( .A1(n6536), .A2(n10181), .B1(n10183), .B2(n7784), .ZN(n7604) );
  OAI211_X1 U9328 ( .C1(n7610), .C2(n8747), .A(n7605), .B(n7604), .ZN(P2_U3222) );
  INV_X1 U9329 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n7607) );
  MUX2_X1 U9330 ( .A(n7607), .B(n7606), .S(n10229), .Z(n7609) );
  NAND2_X1 U9331 ( .A1(n6536), .A2(n8810), .ZN(n7608) );
  OAI211_X1 U9332 ( .C1(n8813), .C2(n7610), .A(n7609), .B(n7608), .ZN(P2_U3470) );
  XNOR2_X1 U9333 ( .A(n7611), .B(n8092), .ZN(n7639) );
  NAND2_X1 U9334 ( .A1(n7613), .A2(n7612), .ZN(n7615) );
  AND2_X1 U9335 ( .A1(n7615), .A2(n7614), .ZN(n7616) );
  XNOR2_X1 U9336 ( .A(n7616), .B(n8092), .ZN(n7617) );
  AOI222_X1 U9337 ( .A1(n10178), .A2(n7617), .B1(n8394), .B2(n10173), .C1(
        n8396), .C2(n10175), .ZN(n7635) );
  MUX2_X1 U9338 ( .A(n7618), .B(n7635), .S(n10217), .Z(n7620) );
  NAND2_X1 U9339 ( .A1(n7636), .A2(n8893), .ZN(n7619) );
  OAI211_X1 U9340 ( .C1(n7639), .C2(n8896), .A(n7620), .B(n7619), .ZN(P2_U3426) );
  XNOR2_X1 U9341 ( .A(n7623), .B(n8394), .ZN(n7624) );
  XNOR2_X1 U9342 ( .A(n7622), .B(n7624), .ZN(n7631) );
  NAND2_X1 U9343 ( .A1(n8371), .A2(n8393), .ZN(n7625) );
  NAND2_X1 U9344 ( .A1(P2_U3151), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n8426) );
  OAI211_X1 U9345 ( .C1(n7626), .C2(n8382), .A(n7625), .B(n8426), .ZN(n7627)
         );
  AOI21_X1 U9346 ( .B1(n7628), .B2(n8385), .A(n7627), .ZN(n7630) );
  NAND2_X1 U9347 ( .A1(n8093), .A2(n8362), .ZN(n7629) );
  OAI211_X1 U9348 ( .C1(n7631), .C2(n8375), .A(n7630), .B(n7629), .ZN(P2_U3174) );
  MUX2_X1 U9349 ( .A(n8407), .B(n7635), .S(n10186), .Z(n7634) );
  AOI22_X1 U9350 ( .A1(n7636), .A2(n10181), .B1(n10183), .B2(n7632), .ZN(n7633) );
  OAI211_X1 U9351 ( .C1(n7639), .C2(n8747), .A(n7634), .B(n7633), .ZN(P2_U3221) );
  MUX2_X1 U9352 ( .A(n8411), .B(n7635), .S(n10229), .Z(n7638) );
  NAND2_X1 U9353 ( .A1(n7636), .A2(n8810), .ZN(n7637) );
  OAI211_X1 U9354 ( .C1(n7639), .C2(n8813), .A(n7638), .B(n7637), .ZN(P2_U3471) );
  NOR2_X1 U9355 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n7679) );
  NOR2_X1 U9356 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n7675) );
  NOR2_X1 U9357 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n7672) );
  NOR2_X1 U9358 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n7670) );
  NOR2_X1 U9359 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n7668) );
  NOR2_X1 U9360 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n7666) );
  NOR2_X1 U9361 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n7663) );
  NOR2_X1 U9362 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n7661) );
  NOR2_X1 U9363 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n7659) );
  NOR2_X1 U9364 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n7657) );
  NOR2_X1 U9365 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n7655) );
  NOR2_X1 U9366 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(P1_ADDR_REG_6__SCAN_IN), 
        .ZN(n7653) );
  NOR2_X1 U9367 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n7651) );
  NOR2_X1 U9368 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n7648) );
  NAND2_X1 U9369 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n7646) );
  INV_X1 U9370 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n9412) );
  XNOR2_X1 U9371 ( .A(n9412), .B(P2_ADDR_REG_3__SCAN_IN), .ZN(n10265) );
  NAND2_X1 U9372 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n7644) );
  AOI21_X1 U9373 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(P2_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10231) );
  INV_X1 U9374 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n7641) );
  NAND2_X1 U9375 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .ZN(n7640) );
  NOR2_X1 U9376 ( .A1(n7641), .A2(n7640), .ZN(n10230) );
  NOR2_X1 U9377 ( .A1(P2_ADDR_REG_1__SCAN_IN), .A2(n10230), .ZN(n7642) );
  NOR2_X1 U9378 ( .A1(n10231), .A2(n7642), .ZN(n10263) );
  XOR2_X1 U9379 ( .A(P2_ADDR_REG_2__SCAN_IN), .B(P1_ADDR_REG_2__SCAN_IN), .Z(
        n10262) );
  NAND2_X1 U9380 ( .A1(n10263), .A2(n10262), .ZN(n7643) );
  NAND2_X1 U9381 ( .A1(n7644), .A2(n7643), .ZN(n10264) );
  NAND2_X1 U9382 ( .A1(n10265), .A2(n10264), .ZN(n7645) );
  NAND2_X1 U9383 ( .A1(n7646), .A2(n7645), .ZN(n10267) );
  XOR2_X1 U9384 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(n10169), .Z(n10266) );
  NOR2_X1 U9385 ( .A1(n10267), .A2(n10266), .ZN(n7647) );
  NOR2_X1 U9386 ( .A1(n7648), .A2(n7647), .ZN(n10255) );
  XOR2_X1 U9387 ( .A(n7649), .B(P1_ADDR_REG_5__SCAN_IN), .Z(n10254) );
  NOR2_X1 U9388 ( .A1(n10255), .A2(n10254), .ZN(n7650) );
  NOR2_X1 U9389 ( .A1(n7651), .A2(n7650), .ZN(n10253) );
  XOR2_X1 U9390 ( .A(n8977), .B(P1_ADDR_REG_6__SCAN_IN), .Z(n10252) );
  NOR2_X1 U9391 ( .A1(n10253), .A2(n10252), .ZN(n7652) );
  NOR2_X1 U9392 ( .A1(n7653), .A2(n7652), .ZN(n10259) );
  INV_X1 U9393 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n9465) );
  XOR2_X1 U9394 ( .A(P2_ADDR_REG_7__SCAN_IN), .B(n9465), .Z(n10258) );
  NOR2_X1 U9395 ( .A1(n10259), .A2(n10258), .ZN(n7654) );
  NOR2_X1 U9396 ( .A1(n7655), .A2(n7654), .ZN(n10261) );
  INV_X1 U9397 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n9481) );
  XOR2_X1 U9398 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(n9481), .Z(n10260) );
  NOR2_X1 U9399 ( .A1(n10261), .A2(n10260), .ZN(n7656) );
  NOR2_X1 U9400 ( .A1(n7657), .A2(n7656), .ZN(n10257) );
  XNOR2_X1 U9401 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n10256) );
  NOR2_X1 U9402 ( .A1(n10257), .A2(n10256), .ZN(n7658) );
  NOR2_X1 U9403 ( .A1(n7659), .A2(n7658), .ZN(n10251) );
  XOR2_X1 U9404 ( .A(n8955), .B(P1_ADDR_REG_10__SCAN_IN), .Z(n10250) );
  NOR2_X1 U9405 ( .A1(n10251), .A2(n10250), .ZN(n7660) );
  XOR2_X1 U9406 ( .A(n8998), .B(P1_ADDR_REG_11__SCAN_IN), .Z(n10248) );
  NOR2_X1 U9407 ( .A1(n10249), .A2(n10248), .ZN(n7662) );
  XOR2_X1 U9408 ( .A(P2_ADDR_REG_12__SCAN_IN), .B(n7664), .Z(n10246) );
  NOR2_X1 U9409 ( .A1(n10247), .A2(n10246), .ZN(n7665) );
  INV_X1 U9410 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n9522) );
  INV_X1 U9411 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n8430) );
  AOI22_X1 U9412 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(n9522), .B1(
        P1_ADDR_REG_13__SCAN_IN), .B2(n8430), .ZN(n10244) );
  NOR2_X1 U9413 ( .A1(n10245), .A2(n10244), .ZN(n7667) );
  XOR2_X1 U9414 ( .A(P2_ADDR_REG_14__SCAN_IN), .B(n9539), .Z(n10242) );
  NOR2_X1 U9415 ( .A1(n10243), .A2(n10242), .ZN(n7669) );
  INV_X1 U9416 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n9978) );
  INV_X1 U9417 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n8474) );
  AOI22_X1 U9418 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(n9978), .B1(
        P1_ADDR_REG_15__SCAN_IN), .B2(n8474), .ZN(n10240) );
  NOR2_X1 U9419 ( .A1(n10241), .A2(n10240), .ZN(n7671) );
  NOR2_X1 U9420 ( .A1(n7672), .A2(n7671), .ZN(n10239) );
  INV_X1 U9421 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n9560) );
  INV_X1 U9422 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n7673) );
  AOI22_X1 U9423 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(n9560), .B1(
        P1_ADDR_REG_16__SCAN_IN), .B2(n7673), .ZN(n10238) );
  NOR2_X1 U9424 ( .A1(n10239), .A2(n10238), .ZN(n7674) );
  NOR2_X1 U9425 ( .A1(n7675), .A2(n7674), .ZN(n10237) );
  INV_X1 U9426 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n7677) );
  INV_X1 U9427 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n7676) );
  AOI22_X1 U9428 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(n7677), .B1(
        P1_ADDR_REG_17__SCAN_IN), .B2(n7676), .ZN(n10236) );
  NOR2_X1 U9429 ( .A1(n10237), .A2(n10236), .ZN(n7678) );
  NOR2_X1 U9430 ( .A1(n7679), .A2(n7678), .ZN(n7680) );
  NOR2_X1 U9431 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n7680), .ZN(n10234) );
  AND2_X1 U9432 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n7680), .ZN(n10233) );
  NOR2_X1 U9433 ( .A1(P2_ADDR_REG_18__SCAN_IN), .A2(n10233), .ZN(n7681) );
  NOR2_X1 U9434 ( .A1(n10234), .A2(n7681), .ZN(n7683) );
  XNOR2_X1 U9435 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(P1_ADDR_REG_19__SCAN_IN), 
        .ZN(n7682) );
  XNOR2_X1 U9436 ( .A(n7683), .B(n7682), .ZN(ADD_1068_U4) );
  OAI222_X1 U9437 ( .A1(n8905), .A2(n7686), .B1(P2_U3151), .B2(n7685), .C1(
        n9059), .C2(n7684), .ZN(P2_U3269) );
  MUX2_X1 U9438 ( .A(n7687), .B(n7690), .S(n10217), .Z(n7689) );
  NAND2_X1 U9439 ( .A1(n8093), .A2(n8893), .ZN(n7688) );
  OAI211_X1 U9440 ( .C1(n7693), .C2(n8896), .A(n7689), .B(n7688), .ZN(P2_U3429) );
  MUX2_X1 U9441 ( .A(n4851), .B(n7690), .S(n10229), .Z(n7692) );
  NAND2_X1 U9442 ( .A1(n8093), .A2(n8810), .ZN(n7691) );
  OAI211_X1 U9443 ( .C1(n8813), .C2(n7693), .A(n7692), .B(n7691), .ZN(P2_U3472) );
  INV_X1 U9444 ( .A(n7694), .ZN(n8001) );
  OAI222_X1 U9445 ( .A1(n9059), .A2(n8001), .B1(n8534), .B2(P2_U3151), .C1(
        n7695), .C2(n8905), .ZN(P2_U3268) );
  XNOR2_X1 U9446 ( .A(n7697), .B(n7696), .ZN(n7709) );
  OAI21_X1 U9447 ( .B1(P2_REG1_REG_11__SCAN_IN), .B2(n7699), .A(n7698), .ZN(
        n7707) );
  NAND2_X1 U9448 ( .A1(P2_U3151), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n7780) );
  NAND2_X1 U9449 ( .A1(n10125), .A2(n7700), .ZN(n7701) );
  OAI211_X1 U9450 ( .C1(n10170), .C2(n8998), .A(n7780), .B(n7701), .ZN(n7706)
         );
  XOR2_X1 U9451 ( .A(n7703), .B(n7702), .Z(n7704) );
  NOR2_X1 U9452 ( .A1(n7704), .A2(n8570), .ZN(n7705) );
  AOI211_X1 U9453 ( .C1(n10129), .C2(n7707), .A(n7706), .B(n7705), .ZN(n7708)
         );
  OAI21_X1 U9454 ( .B1(n7709), .B2(n10133), .A(n7708), .ZN(P2_U3193) );
  INV_X1 U9455 ( .A(n8718), .ZN(n7717) );
  NAND2_X1 U9456 ( .A1(n7710), .A2(n7983), .ZN(n7985) );
  INV_X1 U9457 ( .A(n7711), .ZN(n7712) );
  NAND2_X1 U9458 ( .A1(n7985), .A2(n7712), .ZN(n7713) );
  NAND2_X1 U9459 ( .A1(n7713), .A2(n7714), .ZN(n8719) );
  INV_X1 U9460 ( .A(n7713), .ZN(n7715) );
  NAND2_X1 U9461 ( .A1(n7714), .A2(n8718), .ZN(n8192) );
  AOI21_X1 U9462 ( .B1(n7715), .B2(n8192), .A(n8753), .ZN(n7716) );
  OAI21_X1 U9463 ( .B1(n7717), .B2(n8719), .A(n7716), .ZN(n7719) );
  AOI22_X1 U9464 ( .A1(n8724), .A2(n10173), .B1(n10175), .B2(n8393), .ZN(n7718) );
  AND2_X1 U9465 ( .A1(n7719), .A2(n7718), .ZN(n8817) );
  OR2_X1 U9466 ( .A1(n7720), .A2(n7721), .ZN(n7722) );
  NAND2_X1 U9467 ( .A1(n7722), .A2(n8097), .ZN(n7723) );
  XOR2_X1 U9468 ( .A(n8192), .B(n7723), .Z(n8815) );
  INV_X1 U9469 ( .A(n8747), .ZN(n10182) );
  INV_X1 U9470 ( .A(n8814), .ZN(n8390) );
  AOI22_X1 U9471 ( .A1(n10187), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n10183), 
        .B2(n8386), .ZN(n7724) );
  OAI21_X1 U9472 ( .B1(n8390), .B2(n8581), .A(n7724), .ZN(n7725) );
  AOI21_X1 U9473 ( .B1(n8815), .B2(n10182), .A(n7725), .ZN(n7726) );
  OAI21_X1 U9474 ( .B1(n8817), .B2(n10187), .A(n7726), .ZN(P2_U3218) );
  XNOR2_X1 U9475 ( .A(n7490), .B(n8184), .ZN(n7752) );
  INV_X1 U9476 ( .A(n7752), .ZN(n7735) );
  NAND2_X1 U9477 ( .A1(n7728), .A2(n7727), .ZN(n7729) );
  XOR2_X1 U9478 ( .A(n8184), .B(n7729), .Z(n7730) );
  OAI222_X1 U9479 ( .A1(n8737), .A2(n8322), .B1(n8739), .B2(n7782), .C1(n7730), 
        .C2(n8753), .ZN(n7751) );
  INV_X1 U9480 ( .A(n7751), .ZN(n7731) );
  MUX2_X1 U9481 ( .A(n7732), .B(n7731), .S(n10186), .Z(n7734) );
  AOI22_X1 U9482 ( .A1(n8324), .A2(n10181), .B1(n10183), .B2(n8325), .ZN(n7733) );
  OAI211_X1 U9483 ( .C1(n7735), .C2(n8747), .A(n7734), .B(n7733), .ZN(P2_U3224) );
  XNOR2_X1 U9484 ( .A(n7736), .B(n7741), .ZN(n9916) );
  NAND2_X1 U9485 ( .A1(n7575), .A2(n7737), .ZN(n7740) );
  INV_X1 U9486 ( .A(n7738), .ZN(n7739) );
  AOI21_X1 U9487 ( .B1(n7741), .B2(n7740), .A(n7739), .ZN(n7743) );
  AND2_X1 U9488 ( .A1(n9365), .A2(n9305), .ZN(n7742) );
  AOI21_X1 U9489 ( .B1(n9363), .B2(n9304), .A(n7742), .ZN(n9346) );
  OAI21_X1 U9490 ( .B1(n7743), .B2(n10000), .A(n9346), .ZN(n9912) );
  INV_X1 U9491 ( .A(n9812), .ZN(n7745) );
  AOI211_X1 U9492 ( .C1(n9914), .C2(n6483), .A(n8236), .B(n7745), .ZN(n9913)
         );
  NAND2_X1 U9493 ( .A1(n9913), .A2(n10046), .ZN(n7747) );
  AOI22_X1 U9494 ( .A1(n9768), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n9342), .B2(
        n10041), .ZN(n7746) );
  OAI211_X1 U9495 ( .C1(n7748), .C2(n9816), .A(n7747), .B(n7746), .ZN(n7749)
         );
  AOI21_X1 U9496 ( .B1(n9912), .B2(n9996), .A(n7749), .ZN(n7750) );
  OAI21_X1 U9497 ( .B1(n9916), .B2(n9828), .A(n7750), .ZN(P1_U3278) );
  INV_X1 U9498 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n7753) );
  AOI21_X1 U9499 ( .B1(n7752), .B2(n10201), .A(n7751), .ZN(n7755) );
  MUX2_X1 U9500 ( .A(n7753), .B(n7755), .S(n10217), .Z(n7754) );
  OAI21_X1 U9501 ( .B1(n7758), .B2(n8845), .A(n7754), .ZN(P2_U3417) );
  MUX2_X1 U9502 ( .A(n7756), .B(n7755), .S(n10229), .Z(n7757) );
  OAI21_X1 U9503 ( .B1(n7758), .B2(n8780), .A(n7757), .ZN(P2_U3468) );
  INV_X1 U9504 ( .A(n7760), .ZN(n7761) );
  AND2_X1 U9505 ( .A1(n7759), .A2(n7761), .ZN(n7762) );
  NAND2_X1 U9506 ( .A1(n7762), .A2(n7782), .ZN(n7775) );
  INV_X1 U9507 ( .A(n7762), .ZN(n7763) );
  NAND2_X1 U9508 ( .A1(n7763), .A2(n8397), .ZN(n7774) );
  NAND2_X1 U9509 ( .A1(n7775), .A2(n7774), .ZN(n7764) );
  XOR2_X1 U9510 ( .A(n7776), .B(n7764), .Z(n7773) );
  NAND2_X1 U9511 ( .A1(n8371), .A2(n8396), .ZN(n7766) );
  OAI211_X1 U9512 ( .C1(n7767), .C2(n8382), .A(n7766), .B(n7765), .ZN(n7768)
         );
  AOI21_X1 U9513 ( .B1(n7769), .B2(n8385), .A(n7768), .ZN(n7772) );
  NAND2_X1 U9514 ( .A1(n7770), .A2(n8362), .ZN(n7771) );
  OAI211_X1 U9515 ( .C1(n7773), .C2(n8375), .A(n7772), .B(n7771), .ZN(P2_U3157) );
  INV_X1 U9516 ( .A(n7774), .ZN(n7777) );
  OAI21_X1 U9517 ( .B1(n7777), .B2(n7776), .A(n7775), .ZN(n7778) );
  XOR2_X1 U9518 ( .A(n7779), .B(n7778), .Z(n7787) );
  NAND2_X1 U9519 ( .A1(n8371), .A2(n8395), .ZN(n7781) );
  OAI211_X1 U9520 ( .C1(n7782), .C2(n8382), .A(n7781), .B(n7780), .ZN(n7783)
         );
  AOI21_X1 U9521 ( .B1(n7784), .B2(n8385), .A(n7783), .ZN(n7786) );
  NAND2_X1 U9522 ( .A1(n6536), .A2(n8362), .ZN(n7785) );
  OAI211_X1 U9523 ( .C1(n7787), .C2(n8375), .A(n7786), .B(n7785), .ZN(P2_U3176) );
  INV_X1 U9524 ( .A(n7789), .ZN(n7790) );
  AOI21_X1 U9525 ( .B1(n7791), .B2(n7788), .A(n7790), .ZN(n7797) );
  NAND2_X1 U9526 ( .A1(n8371), .A2(n8392), .ZN(n7792) );
  NAND2_X1 U9527 ( .A1(P2_U3151), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n8439) );
  OAI211_X1 U9528 ( .C1(n7793), .C2(n8382), .A(n7792), .B(n8439), .ZN(n7794)
         );
  AOI21_X1 U9529 ( .B1(n7997), .B2(n8385), .A(n7794), .ZN(n7796) );
  NAND2_X1 U9530 ( .A1(n7993), .A2(n8362), .ZN(n7795) );
  OAI211_X1 U9531 ( .C1(n7797), .C2(n8375), .A(n7796), .B(n7795), .ZN(P2_U3155) );
  OAI222_X1 U9532 ( .A1(n8253), .A2(n7799), .B1(n9963), .B2(n7798), .C1(
        P1_U3086), .C2(n9788), .ZN(P1_U3336) );
  AOI22_X1 U9533 ( .A1(n9373), .A2(n7930), .B1(n6425), .B2(n7904), .ZN(n7803)
         );
  AOI22_X1 U9534 ( .A1(n9373), .A2(n9129), .B1(n7884), .B2(n6425), .ZN(n9215)
         );
  NAND2_X1 U9535 ( .A1(n10083), .A2(n7884), .ZN(n7806) );
  NAND2_X1 U9536 ( .A1(n9372), .A2(n9129), .ZN(n7805) );
  NAND2_X1 U9537 ( .A1(n7806), .A2(n7805), .ZN(n7808) );
  AOI22_X1 U9538 ( .A1(n10083), .A2(n7904), .B1(n9372), .B2(n7930), .ZN(n7807)
         );
  XNOR2_X1 U9539 ( .A(n7807), .B(n4278), .ZN(n7810) );
  XOR2_X1 U9540 ( .A(n7808), .B(n7810), .Z(n9314) );
  INV_X1 U9541 ( .A(n7808), .ZN(n7809) );
  NAND2_X1 U9542 ( .A1(n10007), .A2(n7904), .ZN(n7812) );
  NAND2_X1 U9543 ( .A1(n9371), .A2(n7930), .ZN(n7811) );
  NAND2_X1 U9544 ( .A1(n7812), .A2(n7811), .ZN(n7813) );
  XNOR2_X1 U9545 ( .A(n7813), .B(n4278), .ZN(n9065) );
  NAND2_X1 U9546 ( .A1(n10007), .A2(n4290), .ZN(n7815) );
  NAND2_X1 U9547 ( .A1(n9371), .A2(n9129), .ZN(n7814) );
  NAND2_X1 U9548 ( .A1(n7815), .A2(n7814), .ZN(n9064) );
  OR2_X1 U9549 ( .A1(n9065), .A2(n9064), .ZN(n7816) );
  NAND2_X1 U9550 ( .A1(n9157), .A2(n7904), .ZN(n7818) );
  NAND2_X1 U9551 ( .A1(n9370), .A2(n7884), .ZN(n7817) );
  NAND2_X1 U9552 ( .A1(n7818), .A2(n7817), .ZN(n7820) );
  XNOR2_X1 U9553 ( .A(n7820), .B(n6923), .ZN(n9250) );
  NOR2_X1 U9554 ( .A1(n9069), .A2(n4288), .ZN(n7821) );
  AOI21_X1 U9555 ( .B1(n9157), .B2(n4289), .A(n7821), .ZN(n7829) );
  NAND2_X1 U9556 ( .A1(n9065), .A2(n9064), .ZN(n9148) );
  OAI21_X1 U9557 ( .B1(n9250), .B2(n7829), .A(n9148), .ZN(n7822) );
  INV_X1 U9558 ( .A(n7822), .ZN(n7823) );
  NAND2_X1 U9559 ( .A1(n5388), .A2(n7904), .ZN(n7825) );
  NAND2_X1 U9560 ( .A1(n9369), .A2(n7884), .ZN(n7824) );
  NAND2_X1 U9561 ( .A1(n7825), .A2(n7824), .ZN(n7826) );
  XNOR2_X1 U9562 ( .A(n7826), .B(n4278), .ZN(n7838) );
  NOR2_X1 U9563 ( .A1(n7827), .A2(n4288), .ZN(n7828) );
  AOI21_X1 U9564 ( .B1(n5388), .B2(n4290), .A(n7828), .ZN(n7836) );
  XNOR2_X1 U9565 ( .A(n7838), .B(n7836), .ZN(n9252) );
  INV_X1 U9566 ( .A(n9250), .ZN(n9150) );
  INV_X1 U9567 ( .A(n7829), .ZN(n9152) );
  NAND2_X1 U9568 ( .A1(n9299), .A2(n7904), .ZN(n7832) );
  NAND2_X1 U9569 ( .A1(n9368), .A2(n4290), .ZN(n7831) );
  NAND2_X1 U9570 ( .A1(n7832), .A2(n7831), .ZN(n7833) );
  XNOR2_X1 U9571 ( .A(n7833), .B(n6923), .ZN(n7849) );
  NOR2_X1 U9572 ( .A1(n7834), .A2(n6852), .ZN(n7835) );
  AOI21_X1 U9573 ( .B1(n9299), .B2(n7884), .A(n7835), .ZN(n7848) );
  INV_X1 U9574 ( .A(n7836), .ZN(n7837) );
  NAND2_X1 U9575 ( .A1(n7838), .A2(n7837), .ZN(n7845) );
  INV_X1 U9576 ( .A(n7845), .ZN(n9106) );
  NAND2_X1 U9577 ( .A1(n7841), .A2(n4290), .ZN(n7840) );
  NAND2_X1 U9578 ( .A1(n6436), .A2(n9129), .ZN(n7839) );
  NAND2_X1 U9579 ( .A1(n7840), .A2(n7839), .ZN(n7847) );
  NAND2_X1 U9580 ( .A1(n7841), .A2(n7904), .ZN(n7843) );
  NAND2_X1 U9581 ( .A1(n6436), .A2(n7930), .ZN(n7842) );
  NAND2_X1 U9582 ( .A1(n7843), .A2(n7842), .ZN(n7844) );
  XNOR2_X1 U9583 ( .A(n7844), .B(n6923), .ZN(n9104) );
  NAND2_X1 U9584 ( .A1(n9104), .A2(n7845), .ZN(n9103) );
  OAI21_X1 U9585 ( .B1(n9106), .B2(n7847), .A(n9103), .ZN(n7846) );
  INV_X1 U9586 ( .A(n9180), .ZN(n7851) );
  NAND2_X1 U9587 ( .A1(n9104), .A2(n9178), .ZN(n7850) );
  NAND2_X1 U9588 ( .A1(n7849), .A2(n7848), .ZN(n9181) );
  INV_X1 U9589 ( .A(n7852), .ZN(n7853) );
  INV_X1 U9590 ( .A(n7904), .ZN(n7954) );
  OAI22_X1 U9591 ( .A1(n9191), .A2(n7954), .B1(n7854), .B2(n7056), .ZN(n7855)
         );
  XNOR2_X1 U9592 ( .A(n7855), .B(n6923), .ZN(n7857) );
  AND2_X1 U9593 ( .A1(n9367), .A2(n9129), .ZN(n7856) );
  AOI21_X1 U9594 ( .B1(n9928), .B2(n7930), .A(n7856), .ZN(n7858) );
  NAND2_X1 U9595 ( .A1(n7857), .A2(n7858), .ZN(n7862) );
  INV_X1 U9596 ( .A(n7857), .ZN(n7860) );
  INV_X1 U9597 ( .A(n7858), .ZN(n7859) );
  NAND2_X1 U9598 ( .A1(n7860), .A2(n7859), .ZN(n7861) );
  AND2_X1 U9599 ( .A1(n7862), .A2(n7861), .ZN(n9182) );
  AOI22_X1 U9600 ( .A1(n9922), .A2(n7904), .B1(n7884), .B2(n9366), .ZN(n7863)
         );
  XOR2_X1 U9601 ( .A(n4278), .B(n7863), .Z(n7866) );
  OAI22_X1 U9602 ( .A1(n9281), .A2(n7056), .B1(n7864), .B2(n6852), .ZN(n7865)
         );
  NOR2_X1 U9603 ( .A1(n7866), .A2(n7865), .ZN(n7867) );
  AOI21_X1 U9604 ( .B1(n7866), .B2(n7865), .A(n7867), .ZN(n9274) );
  INV_X1 U9605 ( .A(n7867), .ZN(n7868) );
  AOI22_X1 U9607 ( .A1(n5461), .A2(n7904), .B1(n7930), .B2(n9365), .ZN(n7869)
         );
  XOR2_X1 U9608 ( .A(n4278), .B(n7869), .Z(n7870) );
  AOI22_X1 U9609 ( .A1(n5461), .A2(n7930), .B1(n9129), .B2(n9365), .ZN(n9079)
         );
  NAND2_X1 U9610 ( .A1(n7871), .A2(n7870), .ZN(n9077) );
  AOI22_X1 U9611 ( .A1(n9914), .A2(n7904), .B1(n7884), .B2(n9364), .ZN(n7872)
         );
  XOR2_X1 U9612 ( .A(n4278), .B(n7872), .Z(n7879) );
  NAND2_X1 U9613 ( .A1(n7880), .A2(n7879), .ZN(n9205) );
  AND2_X1 U9614 ( .A1(n9364), .A2(n9129), .ZN(n7873) );
  AOI21_X1 U9615 ( .B1(n9914), .B2(n4290), .A(n7873), .ZN(n9206) );
  NAND2_X1 U9616 ( .A1(n9908), .A2(n7904), .ZN(n7875) );
  NAND2_X1 U9617 ( .A1(n9363), .A2(n4289), .ZN(n7874) );
  NAND2_X1 U9618 ( .A1(n7875), .A2(n7874), .ZN(n7876) );
  XNOR2_X1 U9619 ( .A(n7876), .B(n4278), .ZN(n9208) );
  NAND2_X1 U9620 ( .A1(n9908), .A2(n4290), .ZN(n7878) );
  NAND2_X1 U9621 ( .A1(n9363), .A2(n9129), .ZN(n7877) );
  NAND2_X1 U9622 ( .A1(n7878), .A2(n7877), .ZN(n9207) );
  NAND2_X1 U9623 ( .A1(n9208), .A2(n9207), .ZN(n7881) );
  NAND3_X1 U9624 ( .A1(n9205), .A2(n9206), .A3(n7881), .ZN(n7888) );
  AOI22_X1 U9625 ( .A1(n9903), .A2(n7904), .B1(n4290), .B2(n9362), .ZN(n7882)
         );
  XNOR2_X1 U9626 ( .A(n7882), .B(n4278), .ZN(n7889) );
  AND2_X1 U9627 ( .A1(n9362), .A2(n9129), .ZN(n7883) );
  AOI21_X1 U9628 ( .B1(n9903), .B2(n4289), .A(n7883), .ZN(n7890) );
  XNOR2_X1 U9629 ( .A(n7889), .B(n7890), .ZN(n9226) );
  INV_X1 U9630 ( .A(n9208), .ZN(n7886) );
  INV_X1 U9631 ( .A(n9207), .ZN(n7885) );
  INV_X1 U9632 ( .A(n7889), .ZN(n7892) );
  NAND2_X1 U9633 ( .A1(n7892), .A2(n7891), .ZN(n7893) );
  NAND2_X1 U9634 ( .A1(n9228), .A2(n7893), .ZN(n9117) );
  NAND2_X1 U9635 ( .A1(n9898), .A2(n7904), .ZN(n7895) );
  NAND2_X1 U9636 ( .A1(n9361), .A2(n7884), .ZN(n7894) );
  NAND2_X1 U9637 ( .A1(n7895), .A2(n7894), .ZN(n7896) );
  XNOR2_X1 U9638 ( .A(n7896), .B(n4278), .ZN(n9118) );
  INV_X1 U9639 ( .A(n9118), .ZN(n9162) );
  NAND2_X1 U9640 ( .A1(n9898), .A2(n7884), .ZN(n7898) );
  NAND2_X1 U9641 ( .A1(n9361), .A2(n9129), .ZN(n7897) );
  NAND2_X1 U9642 ( .A1(n7898), .A2(n7897), .ZN(n9167) );
  NAND2_X1 U9643 ( .A1(n9888), .A2(n7904), .ZN(n7900) );
  NAND2_X1 U9644 ( .A1(n9359), .A2(n7930), .ZN(n7899) );
  NAND2_X1 U9645 ( .A1(n7900), .A2(n7899), .ZN(n7901) );
  XNOR2_X1 U9646 ( .A(n7901), .B(n4278), .ZN(n7913) );
  NAND2_X1 U9647 ( .A1(n9888), .A2(n4289), .ZN(n7903) );
  NAND2_X1 U9648 ( .A1(n9359), .A2(n9129), .ZN(n7902) );
  NAND2_X1 U9649 ( .A1(n7903), .A2(n7902), .ZN(n7914) );
  NAND2_X1 U9650 ( .A1(n7913), .A2(n7914), .ZN(n9168) );
  NAND2_X1 U9651 ( .A1(n9893), .A2(n7904), .ZN(n7906) );
  NAND2_X1 U9652 ( .A1(n9360), .A2(n7930), .ZN(n7905) );
  NAND2_X1 U9653 ( .A1(n7906), .A2(n7905), .ZN(n7907) );
  XNOR2_X1 U9654 ( .A(n7907), .B(n4278), .ZN(n9120) );
  NAND2_X1 U9655 ( .A1(n9893), .A2(n7884), .ZN(n7909) );
  NAND2_X1 U9656 ( .A1(n9360), .A2(n9129), .ZN(n7908) );
  NAND2_X1 U9657 ( .A1(n7909), .A2(n7908), .ZN(n9119) );
  NAND2_X1 U9658 ( .A1(n9120), .A2(n9119), .ZN(n9262) );
  OAI211_X1 U9659 ( .C1(n9162), .C2(n9302), .A(n9168), .B(n9262), .ZN(n7919)
         );
  NOR3_X1 U9660 ( .A1(n9118), .A2(n9167), .A3(n9119), .ZN(n7912) );
  NAND2_X1 U9661 ( .A1(n9162), .A2(n9302), .ZN(n7910) );
  AOI21_X1 U9662 ( .B1(n7910), .B2(n9119), .A(n9120), .ZN(n7911) );
  OAI21_X1 U9663 ( .B1(n7912), .B2(n7911), .A(n9168), .ZN(n7917) );
  INV_X1 U9664 ( .A(n7913), .ZN(n7916) );
  INV_X1 U9665 ( .A(n7914), .ZN(n7915) );
  NAND2_X1 U9666 ( .A1(n7916), .A2(n7915), .ZN(n9171) );
  OAI22_X1 U9667 ( .A1(n9747), .A2(n7056), .B1(n9285), .B2(n4288), .ZN(n7923)
         );
  OAI22_X1 U9668 ( .A1(n9747), .A2(n7954), .B1(n9285), .B2(n7056), .ZN(n7920)
         );
  XNOR2_X1 U9669 ( .A(n7920), .B(n4278), .ZN(n7922) );
  XOR2_X1 U9670 ( .A(n7923), .B(n7922), .Z(n9169) );
  INV_X1 U9671 ( .A(n7922), .ZN(n7925) );
  INV_X1 U9672 ( .A(n7923), .ZN(n7924) );
  NAND2_X1 U9673 ( .A1(n7925), .A2(n7924), .ZN(n7926) );
  NAND2_X1 U9674 ( .A1(n9878), .A2(n7904), .ZN(n7928) );
  NAND2_X1 U9675 ( .A1(n9357), .A2(n7930), .ZN(n7927) );
  NAND2_X1 U9676 ( .A1(n7928), .A2(n7927), .ZN(n7929) );
  NAND2_X1 U9677 ( .A1(n9878), .A2(n4290), .ZN(n7932) );
  NAND2_X1 U9678 ( .A1(n9357), .A2(n9129), .ZN(n7931) );
  NAND2_X1 U9679 ( .A1(n7932), .A2(n7931), .ZN(n9284) );
  INV_X1 U9680 ( .A(n9284), .ZN(n7938) );
  OAI22_X1 U9681 ( .A1(n9711), .A2(n7954), .B1(n9286), .B2(n7056), .ZN(n7933)
         );
  XNOR2_X1 U9682 ( .A(n7933), .B(n4278), .ZN(n7937) );
  OR2_X1 U9683 ( .A1(n9711), .A2(n7056), .ZN(n7935) );
  INV_X1 U9684 ( .A(n9286), .ZN(n9356) );
  NAND2_X1 U9685 ( .A1(n9356), .A2(n9129), .ZN(n7934) );
  NAND2_X1 U9686 ( .A1(n7935), .A2(n7934), .ZN(n7936) );
  NOR2_X1 U9687 ( .A1(n7937), .A2(n7936), .ZN(n9238) );
  AOI21_X1 U9688 ( .B1(n7937), .B2(n7936), .A(n9238), .ZN(n9092) );
  INV_X1 U9689 ( .A(n9238), .ZN(n7939) );
  NAND2_X1 U9690 ( .A1(n9869), .A2(n7904), .ZN(n7941) );
  NAND2_X1 U9691 ( .A1(n9355), .A2(n7930), .ZN(n7940) );
  NAND2_X1 U9692 ( .A1(n7941), .A2(n7940), .ZN(n7942) );
  XNOR2_X1 U9693 ( .A(n7942), .B(n6923), .ZN(n7944) );
  AND2_X1 U9694 ( .A1(n9355), .A2(n9129), .ZN(n7943) );
  AOI21_X1 U9695 ( .B1(n9869), .B2(n4289), .A(n7943), .ZN(n7945) );
  NAND2_X1 U9696 ( .A1(n7944), .A2(n7945), .ZN(n7950) );
  INV_X1 U9697 ( .A(n7944), .ZN(n7947) );
  INV_X1 U9698 ( .A(n7945), .ZN(n7946) );
  NAND2_X1 U9699 ( .A1(n7947), .A2(n7946), .ZN(n7948) );
  OAI22_X1 U9700 ( .A1(n9680), .A2(n7056), .B1(n9328), .B2(n6852), .ZN(n7958)
         );
  NAND2_X1 U9701 ( .A1(n9863), .A2(n7904), .ZN(n7952) );
  NAND2_X1 U9702 ( .A1(n9354), .A2(n7884), .ZN(n7951) );
  NAND2_X1 U9703 ( .A1(n7952), .A2(n7951), .ZN(n7953) );
  XNOR2_X1 U9704 ( .A(n7953), .B(n4278), .ZN(n7959) );
  XOR2_X1 U9705 ( .A(n7958), .B(n7959), .Z(n9194) );
  OAI22_X1 U9706 ( .A1(n9673), .A2(n7954), .B1(n9196), .B2(n7056), .ZN(n7955)
         );
  XNOR2_X1 U9707 ( .A(n7955), .B(n4278), .ZN(n7962) );
  OR2_X1 U9708 ( .A1(n9673), .A2(n7056), .ZN(n7957) );
  OR2_X1 U9709 ( .A1(n9196), .A2(n4288), .ZN(n7956) );
  NAND2_X1 U9710 ( .A1(n7957), .A2(n7956), .ZN(n7961) );
  XNOR2_X1 U9711 ( .A(n7962), .B(n7961), .ZN(n9322) );
  NOR2_X1 U9712 ( .A1(n7959), .A2(n7958), .ZN(n9323) );
  NOR2_X1 U9713 ( .A1(n9322), .A2(n9323), .ZN(n7960) );
  NAND2_X1 U9714 ( .A1(n7962), .A2(n7961), .ZN(n7972) );
  NAND2_X1 U9715 ( .A1(n9850), .A2(n7904), .ZN(n7964) );
  INV_X1 U9716 ( .A(n9330), .ZN(n9353) );
  NAND2_X1 U9717 ( .A1(n9353), .A2(n4290), .ZN(n7963) );
  NAND2_X1 U9718 ( .A1(n7964), .A2(n7963), .ZN(n7965) );
  XNOR2_X1 U9719 ( .A(n7965), .B(n6923), .ZN(n7968) );
  INV_X1 U9720 ( .A(n7968), .ZN(n7970) );
  NOR2_X1 U9721 ( .A1(n9330), .A2(n6852), .ZN(n7966) );
  AOI21_X1 U9722 ( .B1(n9850), .B2(n4290), .A(n7966), .ZN(n7967) );
  INV_X1 U9723 ( .A(n7967), .ZN(n7969) );
  AOI21_X1 U9724 ( .B1(n7970), .B2(n7969), .A(n9142), .ZN(n7971) );
  AOI21_X1 U9725 ( .B1(n9325), .B2(n7972), .A(n7971), .ZN(n7976) );
  INV_X1 U9726 ( .A(n7971), .ZN(n7974) );
  INV_X1 U9727 ( .A(n7972), .ZN(n7973) );
  NOR2_X1 U9728 ( .A1(n7974), .A2(n7973), .ZN(n7975) );
  OAI21_X1 U9729 ( .B1(n7976), .B2(n9137), .A(n9326), .ZN(n7982) );
  NOR2_X1 U9730 ( .A1(n9196), .A2(n9626), .ZN(n7977) );
  AOI21_X1 U9731 ( .B1(n9612), .B2(n9304), .A(n7977), .ZN(n9660) );
  INV_X1 U9732 ( .A(n9654), .ZN(n7978) );
  AOI22_X1 U9733 ( .A1(n7978), .A2(n9343), .B1(P1_REG3_REG_27__SCAN_IN), .B2(
        P1_U3086), .ZN(n7979) );
  OAI21_X1 U9734 ( .B1(n9660), .B2(n9345), .A(n7979), .ZN(n7980) );
  AOI21_X1 U9735 ( .B1(n9850), .B2(n9348), .A(n7980), .ZN(n7981) );
  NAND2_X1 U9736 ( .A1(n7982), .A2(n7981), .ZN(P1_U3214) );
  XNOR2_X1 U9737 ( .A(n7720), .B(n7983), .ZN(n8000) );
  INV_X1 U9738 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n7988) );
  OR2_X1 U9739 ( .A1(n7710), .A2(n7983), .ZN(n7984) );
  NAND3_X1 U9740 ( .A1(n7985), .A2(n10178), .A3(n7984), .ZN(n7987) );
  AOI22_X1 U9741 ( .A1(n8394), .A2(n10175), .B1(n10173), .B2(n8392), .ZN(n7986) );
  MUX2_X1 U9742 ( .A(n7988), .B(n7994), .S(n10217), .Z(n7990) );
  NAND2_X1 U9743 ( .A1(n7993), .A2(n8893), .ZN(n7989) );
  OAI211_X1 U9744 ( .C1(n8000), .C2(n8896), .A(n7990), .B(n7989), .ZN(P2_U3432) );
  INV_X1 U9745 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n8466) );
  MUX2_X1 U9746 ( .A(n8466), .B(n7994), .S(n10229), .Z(n7992) );
  NAND2_X1 U9747 ( .A1(n7993), .A2(n8810), .ZN(n7991) );
  OAI211_X1 U9748 ( .C1(n8813), .C2(n8000), .A(n7992), .B(n7991), .ZN(P2_U3473) );
  INV_X1 U9749 ( .A(n7993), .ZN(n7995) );
  OAI21_X1 U9750 ( .B1(n7995), .B2(n8628), .A(n7994), .ZN(n7996) );
  NAND2_X1 U9751 ( .A1(n7996), .A2(n10186), .ZN(n7999) );
  AOI22_X1 U9752 ( .A1(n10187), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n10183), 
        .B2(n7997), .ZN(n7998) );
  OAI211_X1 U9753 ( .C1(n8000), .C2(n8747), .A(n7999), .B(n7998), .ZN(P2_U3219) );
  OAI222_X1 U9754 ( .A1(n8253), .A2(n8002), .B1(n9963), .B2(n8001), .C1(n4281), 
        .C2(P1_U3086), .ZN(P1_U3328) );
  INV_X1 U9755 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n8004) );
  MUX2_X1 U9756 ( .A(n8004), .B(n9960), .S(n8003), .Z(n8006) );
  NAND2_X1 U9757 ( .A1(n8252), .A2(n8007), .ZN(n8010) );
  INV_X1 U9758 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n8978) );
  OR2_X1 U9759 ( .A1(n8008), .A2(n8978), .ZN(n8009) );
  INV_X1 U9760 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n8822) );
  AOI22_X1 U9761 ( .A1(n8012), .A2(P2_REG2_REG_31__SCAN_IN), .B1(n8011), .B2(
        P2_REG1_REG_31__SCAN_IN), .ZN(n8013) );
  OAI211_X1 U9762 ( .C1(n4271), .C2(n8822), .A(n8014), .B(n8013), .ZN(n8391)
         );
  INV_X1 U9763 ( .A(n8391), .ZN(n8578) );
  NAND2_X1 U9764 ( .A1(n8015), .A2(n8167), .ZN(n8018) );
  NAND2_X1 U9765 ( .A1(n8823), .A2(n8017), .ZN(n8164) );
  NAND2_X1 U9766 ( .A1(n8164), .A2(n8016), .ZN(n8206) );
  AOI21_X1 U9767 ( .B1(n8018), .B2(n8163), .A(n4984), .ZN(n8019) );
  MUX2_X1 U9768 ( .A(n8601), .B(n8828), .S(n8158), .Z(n8208) );
  NAND2_X1 U9769 ( .A1(n8174), .A2(n8020), .ZN(n8021) );
  NAND2_X1 U9770 ( .A1(n8021), .A2(n6581), .ZN(n8025) );
  NAND2_X1 U9771 ( .A1(n8022), .A2(n5922), .ZN(n8024) );
  AOI21_X1 U9772 ( .B1(n8025), .B2(n8024), .A(n8023), .ZN(n8026) );
  NAND2_X1 U9773 ( .A1(n8033), .A2(n8027), .ZN(n8030) );
  NAND2_X1 U9774 ( .A1(n8045), .A2(n8028), .ZN(n8029) );
  NAND2_X1 U9775 ( .A1(n8035), .A2(n8046), .ZN(n10171) );
  INV_X1 U9776 ( .A(n10171), .ZN(n10180) );
  NAND2_X1 U9777 ( .A1(n8032), .A2(n10180), .ZN(n8049) );
  INV_X1 U9778 ( .A(n8033), .ZN(n8039) );
  INV_X1 U9779 ( .A(n8052), .ZN(n8037) );
  INV_X1 U9780 ( .A(n8035), .ZN(n8036) );
  NOR2_X1 U9781 ( .A1(n8037), .A2(n8036), .ZN(n8038) );
  OAI21_X1 U9782 ( .B1(n8049), .B2(n8039), .A(n8038), .ZN(n8044) );
  INV_X1 U9783 ( .A(n8040), .ZN(n8042) );
  NAND2_X1 U9784 ( .A1(n8042), .A2(n8041), .ZN(n8043) );
  NAND2_X1 U9785 ( .A1(n8044), .A2(n8043), .ZN(n8055) );
  INV_X1 U9786 ( .A(n8045), .ZN(n8048) );
  INV_X1 U9787 ( .A(n8050), .ZN(n8051) );
  AOI21_X1 U9788 ( .B1(n8053), .B2(n8052), .A(n8051), .ZN(n8054) );
  NAND2_X1 U9789 ( .A1(n8068), .A2(n8067), .ZN(n8063) );
  NAND2_X1 U9790 ( .A1(n8063), .A2(n8158), .ZN(n8059) );
  AND2_X1 U9791 ( .A1(n8057), .A2(n8056), .ZN(n8058) );
  AND2_X1 U9792 ( .A1(n8059), .A2(n8058), .ZN(n8071) );
  NAND3_X1 U9793 ( .A1(n8060), .A2(n8071), .A3(n8183), .ZN(n8075) );
  INV_X1 U9794 ( .A(n8061), .ZN(n8065) );
  NOR2_X1 U9795 ( .A1(n8063), .A2(n8062), .ZN(n8064) );
  NOR2_X1 U9796 ( .A1(n8065), .A2(n8064), .ZN(n8073) );
  NAND2_X1 U9797 ( .A1(n8067), .A2(n8066), .ZN(n8070) );
  NAND2_X1 U9798 ( .A1(n8076), .A2(n8068), .ZN(n8069) );
  AOI21_X1 U9799 ( .B1(n8071), .B2(n8070), .A(n8069), .ZN(n8072) );
  MUX2_X1 U9800 ( .A(n8073), .B(n8072), .S(n8165), .Z(n8074) );
  NAND2_X1 U9801 ( .A1(n8075), .A2(n8074), .ZN(n8084) );
  AND2_X1 U9802 ( .A1(n8081), .A2(n8076), .ZN(n8078) );
  INV_X1 U9803 ( .A(n8080), .ZN(n8077) );
  AND2_X1 U9804 ( .A1(n8080), .A2(n8079), .ZN(n8083) );
  INV_X1 U9805 ( .A(n8081), .ZN(n8082) );
  AOI21_X1 U9806 ( .B1(n8084), .B2(n8083), .A(n8082), .ZN(n8085) );
  INV_X1 U9807 ( .A(n8087), .ZN(n8090) );
  INV_X1 U9808 ( .A(n8088), .ZN(n8089) );
  MUX2_X1 U9809 ( .A(n8090), .B(n8089), .S(n8165), .Z(n8091) );
  MUX2_X1 U9810 ( .A(n8394), .B(n8093), .S(n8165), .Z(n8094) );
  MUX2_X1 U9811 ( .A(n8098), .B(n8097), .S(n8165), .Z(n8099) );
  INV_X1 U9812 ( .A(n8100), .ZN(n8102) );
  INV_X1 U9813 ( .A(n8101), .ZN(n8110) );
  OAI22_X1 U9814 ( .A1(n8734), .A2(n8102), .B1(n8110), .B2(n8158), .ZN(n8104)
         );
  NAND3_X1 U9815 ( .A1(n8814), .A2(n8738), .A3(n8165), .ZN(n8103) );
  NAND3_X1 U9816 ( .A1(n8105), .A2(n8104), .A3(n8103), .ZN(n8106) );
  NAND2_X1 U9817 ( .A1(n8106), .A2(n8721), .ZN(n8114) );
  AND2_X1 U9818 ( .A1(n4311), .A2(n8158), .ZN(n8108) );
  AND4_X1 U9819 ( .A1(n8694), .A2(n8122), .A3(n8108), .A4(n8107), .ZN(n8109)
         );
  INV_X1 U9820 ( .A(n8111), .ZN(n8113) );
  AND4_X1 U9821 ( .A1(n8195), .A2(n8165), .A3(n8677), .A4(n8680), .ZN(n8112)
         );
  OAI21_X1 U9822 ( .B1(n8114), .B2(n8113), .A(n8112), .ZN(n8121) );
  NAND3_X1 U9823 ( .A1(n8195), .A2(n8158), .A3(n8687), .ZN(n8115) );
  AND2_X1 U9824 ( .A1(n8115), .A2(n8122), .ZN(n8119) );
  OAI211_X1 U9825 ( .C1(n8694), .C2(n8707), .A(n8165), .B(n8878), .ZN(n8118)
         );
  OAI211_X1 U9826 ( .C1(n8195), .C2(n8687), .A(n8272), .B(n8158), .ZN(n8117)
         );
  NAND3_X1 U9827 ( .A1(n8694), .A2(n8707), .A3(n8165), .ZN(n8116) );
  NAND4_X1 U9828 ( .A1(n8119), .A2(n8118), .A3(n8117), .A4(n8116), .ZN(n8120)
         );
  NAND2_X1 U9829 ( .A1(n8128), .A2(n8122), .ZN(n8125) );
  INV_X1 U9830 ( .A(n8123), .ZN(n8124) );
  MUX2_X1 U9831 ( .A(n8125), .B(n8124), .S(n8158), .Z(n8126) );
  INV_X1 U9832 ( .A(n8127), .ZN(n8130) );
  INV_X1 U9833 ( .A(n8128), .ZN(n8129) );
  MUX2_X1 U9834 ( .A(n8130), .B(n8129), .S(n8158), .Z(n8131) );
  NAND2_X1 U9835 ( .A1(n8197), .A2(n8132), .ZN(n8133) );
  NAND2_X1 U9836 ( .A1(n8133), .A2(n8158), .ZN(n8135) );
  INV_X1 U9837 ( .A(n8134), .ZN(n8198) );
  AND2_X1 U9838 ( .A1(n8135), .A2(n8198), .ZN(n8138) );
  NAND2_X1 U9839 ( .A1(n8142), .A2(n8138), .ZN(n8136) );
  NAND3_X1 U9840 ( .A1(n8136), .A2(n8198), .A3(n8169), .ZN(n8137) );
  INV_X1 U9841 ( .A(n8170), .ZN(n8143) );
  NAND2_X1 U9842 ( .A1(n8137), .A2(n8143), .ZN(n8147) );
  INV_X1 U9843 ( .A(n8138), .ZN(n8140) );
  NOR2_X1 U9844 ( .A1(n8140), .A2(n4894), .ZN(n8141) );
  NAND2_X1 U9845 ( .A1(n8145), .A2(n8169), .ZN(n8146) );
  INV_X1 U9846 ( .A(n8608), .ZN(n8609) );
  INV_X1 U9847 ( .A(n8150), .ZN(n8152) );
  MUX2_X1 U9848 ( .A(n8152), .B(n8151), .S(n8165), .Z(n8153) );
  MUX2_X1 U9849 ( .A(n8156), .B(n8155), .S(n8165), .Z(n8157) );
  MUX2_X1 U9850 ( .A(n8159), .B(n4321), .S(n8158), .Z(n8160) );
  INV_X1 U9851 ( .A(n8206), .ZN(n8163) );
  OAI21_X1 U9852 ( .B1(n8222), .B2(n8601), .A(n8163), .ZN(n8214) );
  OAI21_X1 U9853 ( .B1(n8219), .B2(n8165), .A(n8164), .ZN(n8166) );
  NAND2_X1 U9854 ( .A1(n8166), .A2(n8215), .ZN(n8210) );
  INV_X1 U9855 ( .A(n8210), .ZN(n8213) );
  INV_X1 U9856 ( .A(n8167), .ZN(n8218) );
  XNOR2_X1 U9857 ( .A(n8828), .B(n8168), .ZN(n8586) );
  INV_X1 U9858 ( .A(n8597), .ZN(n8599) );
  INV_X1 U9859 ( .A(n8169), .ZN(n8171) );
  NOR2_X1 U9860 ( .A1(n8171), .A2(n8170), .ZN(n8636) );
  INV_X1 U9861 ( .A(n8721), .ZN(n8194) );
  INV_X1 U9862 ( .A(n8172), .ZN(n8173) );
  AND3_X1 U9863 ( .A1(n6581), .A2(n8173), .A3(n8174), .ZN(n8177) );
  NAND4_X1 U9864 ( .A1(n8177), .A2(n8176), .A3(n8750), .A4(n8175), .ZN(n8180)
         );
  NAND4_X1 U9865 ( .A1(n8184), .A2(n8183), .A3(n8182), .A4(n8181), .ZN(n8185)
         );
  NOR4_X1 U9866 ( .A1(n8188), .A2(n8187), .A3(n8186), .A4(n8185), .ZN(n8190)
         );
  NAND4_X1 U9867 ( .A1(n8192), .A2(n8191), .A3(n8190), .A4(n8189), .ZN(n8193)
         );
  NAND3_X1 U9868 ( .A1(n8196), .A2(n8679), .A3(n8684), .ZN(n8200) );
  NAND2_X1 U9869 ( .A1(n8198), .A2(n8197), .ZN(n8640) );
  NOR4_X1 U9870 ( .A1(n8200), .A2(n8640), .A3(n8199), .A4(n8664), .ZN(n8201)
         );
  INV_X1 U9871 ( .A(n8624), .ZN(n8617) );
  NAND4_X1 U9872 ( .A1(n8609), .A2(n8636), .A3(n8201), .A4(n8617), .ZN(n8202)
         );
  INV_X1 U9873 ( .A(n8219), .ZN(n8203) );
  NAND3_X1 U9874 ( .A1(n8204), .A2(n8203), .A3(n4329), .ZN(n8207) );
  OAI22_X1 U9875 ( .A1(n8207), .A2(n8206), .B1(n8205), .B2(n4329), .ZN(n8212)
         );
  NAND2_X1 U9876 ( .A1(n8209), .A2(n8208), .ZN(n8220) );
  NOR2_X1 U9877 ( .A1(n8210), .A2(n8220), .ZN(n8211) );
  NAND3_X1 U9878 ( .A1(n8216), .A2(n8229), .A3(n8215), .ZN(n8217) );
  NOR3_X1 U9879 ( .A1(n8219), .A2(n8218), .A3(n8217), .ZN(n8221) );
  OAI211_X1 U9880 ( .C1(n8222), .C2(n8828), .A(n8221), .B(n8220), .ZN(n8223)
         );
  NAND3_X1 U9881 ( .A1(n8227), .A2(n8226), .A3(n8534), .ZN(n8228) );
  OAI211_X1 U9882 ( .C1(n8229), .C2(n8231), .A(n8228), .B(P2_B_REG_SCAN_IN), 
        .ZN(n8230) );
  INV_X1 U9883 ( .A(n8909), .ZN(n8233) );
  OAI222_X1 U9884 ( .A1(n8253), .A2(n8234), .B1(n9963), .B2(n8233), .C1(n8232), 
        .C2(P1_U3086), .ZN(P1_U3327) );
  INV_X1 U9885 ( .A(n9619), .ZN(n8235) );
  NOR2_X2 U9886 ( .A1(n9619), .A2(n8244), .ZN(n9604) );
  NOR2_X1 U9887 ( .A1(n9996), .A2(n8239), .ZN(n8243) );
  AND2_X1 U9888 ( .A1(n8240), .A2(P1_B_REG_SCAN_IN), .ZN(n8241) );
  OR2_X1 U9889 ( .A1(n9329), .A2(n8241), .ZN(n9624) );
  OR2_X1 U9890 ( .A1(n8242), .A2(n9624), .ZN(n9831) );
  NOR2_X1 U9891 ( .A1(n9768), .A2(n9831), .ZN(n9607) );
  AOI211_X1 U9892 ( .C1(n8244), .C2(n10042), .A(n8243), .B(n9607), .ZN(n8245)
         );
  OAI21_X1 U9893 ( .B1(n9832), .B2(n9610), .A(n8245), .ZN(P1_U3264) );
  NOR2_X1 U9894 ( .A1(n8246), .A2(n8655), .ZN(n8579) );
  AOI21_X1 U9895 ( .B1(n10187), .B2(P2_REG2_REG_29__SCAN_IN), .A(n8579), .ZN(
        n8247) );
  OAI21_X1 U9896 ( .B1(n8248), .B2(n8581), .A(n8247), .ZN(n8249) );
  AOI21_X1 U9897 ( .B1(n6623), .B2(n8250), .A(n8249), .ZN(n8251) );
  INV_X1 U9898 ( .A(n8252), .ZN(n8903) );
  INV_X1 U9899 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n8254) );
  OAI222_X1 U9900 ( .A1(P1_U3086), .A2(n8255), .B1(n9963), .B2(n8903), .C1(
        n8254), .C2(n8253), .ZN(P1_U3325) );
  OAI21_X1 U9901 ( .B1(n8631), .B2(n8257), .A(n8256), .ZN(n8258) );
  NAND2_X1 U9902 ( .A1(n8258), .A2(n8367), .ZN(n8264) );
  INV_X1 U9903 ( .A(n8645), .ZN(n8261) );
  AOI22_X1 U9904 ( .A1(n8671), .A2(n8356), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3151), .ZN(n8259) );
  OAI21_X1 U9905 ( .B1(n8261), .B2(n8260), .A(n8259), .ZN(n8262) );
  AOI21_X1 U9906 ( .B1(n8642), .B2(n8380), .A(n8262), .ZN(n8263) );
  OAI211_X1 U9907 ( .C1(n8265), .C2(n8389), .A(n8264), .B(n8263), .ZN(P2_U3156) );
  INV_X1 U9908 ( .A(n8266), .ZN(n8268) );
  NAND2_X1 U9909 ( .A1(n8268), .A2(n8267), .ZN(n8269) );
  XNOR2_X1 U9910 ( .A(n8270), .B(n8269), .ZN(n8276) );
  NAND2_X1 U9911 ( .A1(n8725), .A2(n8356), .ZN(n8271) );
  NAND2_X1 U9912 ( .A1(P2_U3151), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8572) );
  OAI211_X1 U9913 ( .C1(n8282), .C2(n8360), .A(n8271), .B(n8572), .ZN(n8274)
         );
  NOR2_X1 U9914 ( .A1(n8272), .A2(n8389), .ZN(n8273) );
  AOI211_X1 U9915 ( .C1(n8702), .C2(n8385), .A(n8274), .B(n8273), .ZN(n8275)
         );
  OAI21_X1 U9916 ( .B1(n8276), .B2(n8375), .A(n8275), .ZN(P2_U3159) );
  OR2_X1 U9917 ( .A1(n8330), .A2(n8331), .ZN(n8338) );
  NAND2_X1 U9918 ( .A1(n8338), .A2(n8277), .ZN(n8278) );
  XOR2_X1 U9919 ( .A(n8279), .B(n8278), .Z(n8285) );
  AOI22_X1 U9920 ( .A1(n8671), .A2(n8371), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3151), .ZN(n8281) );
  NAND2_X1 U9921 ( .A1(n8674), .A2(n8385), .ZN(n8280) );
  OAI211_X1 U9922 ( .C1(n8282), .C2(n8382), .A(n8281), .B(n8280), .ZN(n8283)
         );
  AOI21_X1 U9923 ( .B1(n8866), .B2(n8362), .A(n8283), .ZN(n8284) );
  OAI21_X1 U9924 ( .B1(n8285), .B2(n8375), .A(n8284), .ZN(P2_U3163) );
  INV_X1 U9925 ( .A(n8287), .ZN(n8291) );
  INV_X1 U9926 ( .A(n8288), .ZN(n8290) );
  NOR3_X1 U9927 ( .A1(n8291), .A2(n8290), .A3(n8289), .ZN(n8294) );
  INV_X1 U9928 ( .A(n8292), .ZN(n8293) );
  OAI21_X1 U9929 ( .B1(n8294), .B2(n8293), .A(n8367), .ZN(n8298) );
  AOI22_X1 U9930 ( .A1(n8623), .A2(n8385), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3151), .ZN(n8295) );
  OAI21_X1 U9931 ( .B1(n8621), .B2(n8382), .A(n8295), .ZN(n8296) );
  AOI21_X1 U9932 ( .B1(n8602), .B2(n8380), .A(n8296), .ZN(n8297) );
  OAI211_X1 U9933 ( .C1(n8846), .C2(n8389), .A(n8298), .B(n8297), .ZN(P2_U3165) );
  XNOR2_X1 U9934 ( .A(n8301), .B(n8300), .ZN(n8302) );
  XNOR2_X1 U9935 ( .A(n8303), .B(n8302), .ZN(n8308) );
  NAND2_X1 U9936 ( .A1(n8357), .A2(n8371), .ZN(n8304) );
  NAND2_X1 U9937 ( .A1(P2_U3151), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8493) );
  OAI211_X1 U9938 ( .C1(n8738), .C2(n8382), .A(n8304), .B(n8493), .ZN(n8305)
         );
  AOI21_X1 U9939 ( .B1(n8744), .B2(n8385), .A(n8305), .ZN(n8307) );
  NAND2_X1 U9940 ( .A1(n6553), .A2(n8362), .ZN(n8306) );
  OAI211_X1 U9941 ( .C1(n8308), .C2(n8375), .A(n8307), .B(n8306), .ZN(P2_U3166) );
  XNOR2_X1 U9942 ( .A(n8309), .B(n8740), .ZN(n8310) );
  XNOR2_X1 U9943 ( .A(n8311), .B(n8310), .ZN(n8318) );
  NAND2_X1 U9944 ( .A1(n8356), .A2(n8724), .ZN(n8312) );
  NAND2_X1 U9945 ( .A1(P2_U3151), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n8522) );
  OAI211_X1 U9946 ( .C1(n8313), .C2(n8360), .A(n8312), .B(n8522), .ZN(n8316)
         );
  NOR2_X1 U9947 ( .A1(n8314), .A2(n8389), .ZN(n8315) );
  AOI211_X1 U9948 ( .C1(n8729), .C2(n8385), .A(n8316), .B(n8315), .ZN(n8317)
         );
  OAI21_X1 U9949 ( .B1(n8318), .B2(n8375), .A(n8317), .ZN(P2_U3168) );
  OAI211_X1 U9950 ( .C1(n8319), .C2(n4389), .A(n7759), .B(n8367), .ZN(n8329)
         );
  NAND2_X1 U9951 ( .A1(n8371), .A2(n8397), .ZN(n8321) );
  OAI211_X1 U9952 ( .C1(n8322), .C2(n8382), .A(n8321), .B(n8320), .ZN(n8323)
         );
  INV_X1 U9953 ( .A(n8323), .ZN(n8328) );
  NAND2_X1 U9954 ( .A1(n8324), .A2(n8362), .ZN(n8327) );
  NAND2_X1 U9955 ( .A1(n8385), .A2(n8325), .ZN(n8326) );
  NAND4_X1 U9956 ( .A1(n8329), .A2(n8328), .A3(n8327), .A4(n8326), .ZN(
        P2_U3171) );
  XOR2_X1 U9957 ( .A(n8331), .B(n8330), .Z(n8336) );
  AOI22_X1 U9958 ( .A1(n8688), .A2(n8371), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3151), .ZN(n8333) );
  NAND2_X1 U9959 ( .A1(n8691), .A2(n8385), .ZN(n8332) );
  OAI211_X1 U9960 ( .C1(n8707), .C2(n8382), .A(n8333), .B(n8332), .ZN(n8334)
         );
  AOI21_X1 U9961 ( .B1(n8872), .B2(n8362), .A(n8334), .ZN(n8335) );
  OAI21_X1 U9962 ( .B1(n8336), .B2(n8375), .A(n8335), .ZN(P2_U3173) );
  NAND2_X1 U9963 ( .A1(n8338), .A2(n8337), .ZN(n8340) );
  AND2_X1 U9964 ( .A1(n8340), .A2(n8339), .ZN(n8344) );
  NAND2_X1 U9965 ( .A1(n8342), .A2(n8341), .ZN(n8343) );
  XNOR2_X1 U9966 ( .A(n8344), .B(n8343), .ZN(n8351) );
  INV_X1 U9967 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n8345) );
  OAI22_X1 U9968 ( .A1(n8346), .A2(n8382), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8345), .ZN(n8348) );
  NOR2_X1 U9969 ( .A1(n8631), .A2(n8360), .ZN(n8347) );
  AOI211_X1 U9970 ( .C1(n8653), .C2(n8385), .A(n8348), .B(n8347), .ZN(n8350)
         );
  NAND2_X1 U9971 ( .A1(n8787), .A2(n8362), .ZN(n8349) );
  OAI211_X1 U9972 ( .C1(n8351), .C2(n8375), .A(n8350), .B(n8349), .ZN(P2_U3175) );
  INV_X1 U9973 ( .A(n8352), .ZN(n8353) );
  AOI21_X1 U9974 ( .B1(n8355), .B2(n8354), .A(n8353), .ZN(n8364) );
  AND2_X1 U9975 ( .A1(P2_U3151), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8540) );
  AOI21_X1 U9976 ( .B1(n8357), .B2(n8356), .A(n8540), .ZN(n8359) );
  NAND2_X1 U9977 ( .A1(n8385), .A2(n8712), .ZN(n8358) );
  OAI211_X1 U9978 ( .C1(n8707), .C2(n8360), .A(n8359), .B(n8358), .ZN(n8361)
         );
  AOI21_X1 U9979 ( .B1(n8803), .B2(n8362), .A(n8361), .ZN(n8363) );
  OAI21_X1 U9980 ( .B1(n8364), .B2(n8375), .A(n8363), .ZN(P2_U3178) );
  OAI21_X1 U9981 ( .B1(n8620), .B2(n8366), .A(n8365), .ZN(n8368) );
  NAND2_X1 U9982 ( .A1(n8368), .A2(n8367), .ZN(n8373) );
  AOI22_X1 U9983 ( .A1(n8614), .A2(n8385), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3151), .ZN(n8369) );
  OAI21_X1 U9984 ( .B1(n8632), .B2(n8382), .A(n8369), .ZN(n8370) );
  AOI21_X1 U9985 ( .B1(n8611), .B2(n8371), .A(n8370), .ZN(n8372) );
  OAI211_X1 U9986 ( .C1(n8374), .C2(n8389), .A(n8373), .B(n8372), .ZN(P2_U3180) );
  AOI21_X1 U9987 ( .B1(n8377), .B2(n8376), .A(n8375), .ZN(n8379) );
  NAND2_X1 U9988 ( .A1(n8379), .A2(n8378), .ZN(n8388) );
  NAND2_X1 U9989 ( .A1(n8380), .A2(n8724), .ZN(n8381) );
  NAND2_X1 U9990 ( .A1(P2_U3151), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8473) );
  OAI211_X1 U9991 ( .C1(n8383), .C2(n8382), .A(n8381), .B(n8473), .ZN(n8384)
         );
  AOI21_X1 U9992 ( .B1(n8386), .B2(n8385), .A(n8384), .ZN(n8387) );
  OAI211_X1 U9993 ( .C1(n8390), .C2(n8389), .A(n8388), .B(n8387), .ZN(P2_U3181) );
  MUX2_X1 U9994 ( .A(n8391), .B(P2_DATAO_REG_31__SCAN_IN), .S(n8403), .Z(
        P2_U3522) );
  MUX2_X1 U9995 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n8588), .S(P2_U3893), .Z(
        P2_U3520) );
  MUX2_X1 U9996 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n8601), .S(P2_U3893), .Z(
        P2_U3519) );
  MUX2_X1 U9997 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8611), .S(P2_U3893), .Z(
        P2_U3518) );
  MUX2_X1 U9998 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n8602), .S(P2_U3893), .Z(
        P2_U3517) );
  MUX2_X1 U9999 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n8612), .S(P2_U3893), .Z(
        P2_U3516) );
  MUX2_X1 U10000 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n8642), .S(P2_U3893), .Z(
        P2_U3515) );
  MUX2_X1 U10001 ( .A(n8651), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8403), .Z(
        P2_U3514) );
  MUX2_X1 U10002 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8671), .S(P2_U3893), .Z(
        P2_U3513) );
  MUX2_X1 U10003 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n8688), .S(P2_U3893), .Z(
        P2_U3512) );
  MUX2_X1 U10004 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8699), .S(P2_U3893), .Z(
        P2_U3511) );
  MUX2_X1 U10005 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n8687), .S(P2_U3893), .Z(
        P2_U3510) );
  MUX2_X1 U10006 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n8725), .S(P2_U3893), .Z(
        P2_U3509) );
  MUX2_X1 U10007 ( .A(n8724), .B(P2_DATAO_REG_16__SCAN_IN), .S(n8403), .Z(
        P2_U3507) );
  MUX2_X1 U10008 ( .A(n8392), .B(P2_DATAO_REG_15__SCAN_IN), .S(n8403), .Z(
        P2_U3506) );
  MUX2_X1 U10009 ( .A(n8393), .B(P2_DATAO_REG_14__SCAN_IN), .S(n8403), .Z(
        P2_U3505) );
  MUX2_X1 U10010 ( .A(n8394), .B(P2_DATAO_REG_13__SCAN_IN), .S(n8403), .Z(
        P2_U3504) );
  MUX2_X1 U10011 ( .A(n8395), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8403), .Z(
        P2_U3503) );
  MUX2_X1 U10012 ( .A(n8396), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8403), .Z(
        P2_U3502) );
  MUX2_X1 U10013 ( .A(n8397), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8403), .Z(
        P2_U3501) );
  MUX2_X1 U10014 ( .A(n8398), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8403), .Z(
        P2_U3500) );
  MUX2_X1 U10015 ( .A(n8399), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8403), .Z(
        P2_U3499) );
  MUX2_X1 U10016 ( .A(n8400), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8403), .Z(
        P2_U3498) );
  MUX2_X1 U10017 ( .A(n8401), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8403), .Z(
        P2_U3497) );
  MUX2_X1 U10018 ( .A(n10174), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8403), .Z(
        P2_U3496) );
  MUX2_X1 U10019 ( .A(n8402), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8403), .Z(
        P2_U3495) );
  MUX2_X1 U10020 ( .A(n10176), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8403), .Z(
        P2_U3494) );
  MUX2_X1 U10021 ( .A(n4882), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8403), .Z(
        P2_U3493) );
  MUX2_X1 U10022 ( .A(n4432), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8403), .Z(
        P2_U3492) );
  MUX2_X1 U10023 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(n8404), .S(P2_U3893), .Z(
        P2_U3491) );
  NAND2_X1 U10024 ( .A1(n8406), .A2(n8405), .ZN(n8409) );
  OR2_X1 U10025 ( .A1(n8412), .A2(n8407), .ZN(n8408) );
  XNOR2_X1 U10026 ( .A(n8436), .B(n8410), .ZN(n8434) );
  OR2_X1 U10027 ( .A1(n8412), .A2(n8411), .ZN(n8413) );
  OAI21_X1 U10028 ( .B1(P2_REG1_REG_13__SCAN_IN), .B2(n4382), .A(n8454), .ZN(
        n8432) );
  NAND2_X1 U10029 ( .A1(n8418), .A2(n8417), .ZN(n8423) );
  MUX2_X1 U10030 ( .A(P2_REG2_REG_13__SCAN_IN), .B(P2_REG1_REG_13__SCAN_IN), 
        .S(n8534), .Z(n8420) );
  NOR2_X1 U10031 ( .A1(n8419), .A2(n8420), .ZN(n8441) );
  AOI21_X1 U10032 ( .B1(n8420), .B2(n8419), .A(n8441), .ZN(n8421) );
  NAND3_X1 U10033 ( .A1(n8423), .A2(n8421), .A3(n8422), .ZN(n8446) );
  INV_X1 U10034 ( .A(n8446), .ZN(n8425) );
  AOI21_X1 U10035 ( .B1(n8423), .B2(n8422), .A(n8421), .ZN(n8424) );
  OAI21_X1 U10036 ( .B1(n8425), .B2(n8424), .A(n10166), .ZN(n8429) );
  INV_X1 U10037 ( .A(n8426), .ZN(n8427) );
  AOI21_X1 U10038 ( .B1(n10125), .B2(n8438), .A(n8427), .ZN(n8428) );
  OAI211_X1 U10039 ( .C1(n8430), .C2(n10170), .A(n8429), .B(n8428), .ZN(n8431)
         );
  AOI21_X1 U10040 ( .B1(n10129), .B2(n8432), .A(n8431), .ZN(n8433) );
  OAI21_X1 U10041 ( .B1(n8434), .B2(n10133), .A(n8433), .ZN(P2_U3195) );
  XNOR2_X1 U10042 ( .A(n8467), .B(P2_REG2_REG_14__SCAN_IN), .ZN(n8461) );
  INV_X1 U10043 ( .A(n8435), .ZN(n8437) );
  XOR2_X1 U10044 ( .A(n8461), .B(n8462), .Z(n8460) );
  OAI21_X1 U10045 ( .B1(n10164), .B2(n8440), .A(n8439), .ZN(n8450) );
  INV_X1 U10046 ( .A(n8441), .ZN(n8445) );
  INV_X1 U10047 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n8463) );
  MUX2_X1 U10048 ( .A(n8463), .B(n8466), .S(n8534), .Z(n8442) );
  NAND2_X1 U10049 ( .A1(n8467), .A2(n8442), .ZN(n8475) );
  OR2_X1 U10050 ( .A1(n8467), .A2(n8442), .ZN(n8443) );
  NAND2_X1 U10051 ( .A1(n8475), .A2(n8443), .ZN(n8444) );
  INV_X1 U10052 ( .A(n8483), .ZN(n8448) );
  NAND3_X1 U10053 ( .A1(n8446), .A2(n8445), .A3(n8444), .ZN(n8447) );
  AOI21_X1 U10054 ( .B1(n8448), .B2(n8447), .A(n8570), .ZN(n8449) );
  AOI211_X1 U10055 ( .C1(n10142), .C2(P2_ADDR_REG_14__SCAN_IN), .A(n8450), .B(
        n8449), .ZN(n8459) );
  INV_X1 U10056 ( .A(n8454), .ZN(n8452) );
  INV_X1 U10057 ( .A(n8453), .ZN(n8451) );
  XNOR2_X1 U10058 ( .A(n8467), .B(P2_REG1_REG_14__SCAN_IN), .ZN(n8455) );
  NOR3_X1 U10059 ( .A1(n8452), .A2(n8451), .A3(n8455), .ZN(n8457) );
  INV_X1 U10060 ( .A(n8469), .ZN(n8456) );
  OAI21_X1 U10061 ( .B1(n8457), .B2(n8456), .A(n10129), .ZN(n8458) );
  OAI211_X1 U10062 ( .C1(n8460), .C2(n10133), .A(n8459), .B(n8458), .ZN(
        P2_U3196) );
  NAND2_X1 U10063 ( .A1(n8462), .A2(n8461), .ZN(n8465) );
  OR2_X1 U10064 ( .A1(n8467), .A2(n8463), .ZN(n8464) );
  INV_X1 U10065 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n8477) );
  XNOR2_X1 U10066 ( .A(n8490), .B(n8477), .ZN(n8489) );
  OR2_X1 U10067 ( .A1(n8467), .A2(n8466), .ZN(n8468) );
  AND2_X2 U10068 ( .A1(n8469), .A2(n8468), .ZN(n8470) );
  OAI21_X1 U10069 ( .B1(P2_REG1_REG_15__SCAN_IN), .B2(n8471), .A(n8505), .ZN(
        n8487) );
  NAND2_X1 U10070 ( .A1(n10125), .A2(n8479), .ZN(n8472) );
  OAI211_X1 U10071 ( .C1(n10170), .C2(n8474), .A(n8473), .B(n8472), .ZN(n8486)
         );
  INV_X1 U10072 ( .A(n8475), .ZN(n8482) );
  INV_X1 U10073 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n8476) );
  MUX2_X1 U10074 ( .A(n8477), .B(n8476), .S(n8534), .Z(n8478) );
  NAND2_X1 U10075 ( .A1(n8479), .A2(n8478), .ZN(n8499) );
  OR2_X1 U10076 ( .A1(n8479), .A2(n8478), .ZN(n8480) );
  AND2_X1 U10077 ( .A1(n8499), .A2(n8480), .ZN(n8481) );
  OR3_X1 U10078 ( .A1(n8483), .A2(n8482), .A3(n8481), .ZN(n8484) );
  AOI21_X1 U10079 ( .B1(n8500), .B2(n8484), .A(n8570), .ZN(n8485) );
  AOI211_X1 U10080 ( .C1(n10129), .C2(n8487), .A(n8486), .B(n8485), .ZN(n8488)
         );
  OAI21_X1 U10081 ( .B1(n8489), .B2(n10133), .A(n8488), .ZN(P2_U3197) );
  INV_X1 U10082 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n9039) );
  XNOR2_X1 U10083 ( .A(n8514), .B(n9039), .ZN(n8510) );
  NAND2_X1 U10084 ( .A1(n8491), .A2(n4856), .ZN(n8492) );
  XOR2_X1 U10085 ( .A(n8510), .B(n8511), .Z(n8509) );
  OAI21_X1 U10086 ( .B1(n10164), .B2(n8514), .A(n8493), .ZN(n8503) );
  INV_X1 U10087 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n8809) );
  MUX2_X1 U10088 ( .A(n9039), .B(n8809), .S(n8534), .Z(n8495) );
  NAND2_X1 U10089 ( .A1(n8495), .A2(n8494), .ZN(n8519) );
  INV_X1 U10090 ( .A(n8495), .ZN(n8496) );
  NAND2_X1 U10091 ( .A1(n8496), .A2(n8514), .ZN(n8497) );
  NAND2_X1 U10092 ( .A1(n8519), .A2(n8497), .ZN(n8498) );
  NAND3_X1 U10093 ( .A1(n8500), .A2(n8499), .A3(n8498), .ZN(n8501) );
  AOI21_X1 U10094 ( .B1(n4335), .B2(n8501), .A(n8570), .ZN(n8502) );
  AOI211_X1 U10095 ( .C1(n10142), .C2(P2_ADDR_REG_16__SCAN_IN), .A(n8503), .B(
        n8502), .ZN(n8508) );
  XNOR2_X1 U10096 ( .A(n8514), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n8504) );
  AND3_X1 U10097 ( .A1(n8505), .A2(n8504), .A3(n4313), .ZN(n8506) );
  OAI21_X1 U10098 ( .B1(n8516), .B2(n8506), .A(n10129), .ZN(n8507) );
  OAI211_X1 U10099 ( .C1(n8509), .C2(n10133), .A(n8508), .B(n8507), .ZN(
        P2_U3198) );
  NAND2_X1 U10100 ( .A1(n8514), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n8512) );
  NAND2_X1 U10101 ( .A1(n8513), .A2(n8512), .ZN(n8541) );
  XNOR2_X1 U10102 ( .A(n8541), .B(n8533), .ZN(n8543) );
  XOR2_X1 U10103 ( .A(P2_REG2_REG_17__SCAN_IN), .B(n8543), .Z(n8529) );
  OAI21_X1 U10104 ( .B1(P2_REG1_REG_17__SCAN_IN), .B2(n8518), .A(n8547), .ZN(
        n8527) );
  INV_X1 U10105 ( .A(n8519), .ZN(n8520) );
  MUX2_X1 U10106 ( .A(P2_REG2_REG_17__SCAN_IN), .B(P2_REG1_REG_17__SCAN_IN), 
        .S(n8534), .Z(n8530) );
  XOR2_X1 U10107 ( .A(n8533), .B(n8530), .Z(n8521) );
  AOI21_X1 U10108 ( .B1(n4622), .B2(n8521), .A(n8531), .ZN(n8525) );
  OAI21_X1 U10109 ( .B1(n10164), .B2(n8542), .A(n8522), .ZN(n8523) );
  AOI21_X1 U10110 ( .B1(n10142), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n8523), .ZN(
        n8524) );
  OAI21_X1 U10111 ( .B1(n8525), .B2(n8570), .A(n8524), .ZN(n8526) );
  AOI21_X1 U10112 ( .B1(n10129), .B2(n8527), .A(n8526), .ZN(n8528) );
  OAI21_X1 U10113 ( .B1(n8529), .B2(n10133), .A(n8528), .ZN(P2_U3199) );
  INV_X1 U10114 ( .A(n8530), .ZN(n8532) );
  MUX2_X1 U10115 ( .A(P2_REG2_REG_18__SCAN_IN), .B(P2_REG1_REG_18__SCAN_IN), 
        .S(n8534), .Z(n8535) );
  NOR2_X1 U10116 ( .A1(n8536), .A2(n8535), .ZN(n8563) );
  NAND2_X1 U10117 ( .A1(n8536), .A2(n8535), .ZN(n8561) );
  INV_X1 U10118 ( .A(n8561), .ZN(n8537) );
  AOI21_X1 U10119 ( .B1(n8538), .B2(P2_U3893), .A(n10125), .ZN(n8539) );
  AOI21_X1 U10120 ( .B1(n10142), .B2(P2_ADDR_REG_18__SCAN_IN), .A(n8540), .ZN(
        n8552) );
  XOR2_X1 U10121 ( .A(P2_REG2_REG_18__SCAN_IN), .B(n8562), .Z(n8554) );
  XNOR2_X1 U10122 ( .A(n8555), .B(n8554), .ZN(n8544) );
  NAND2_X1 U10123 ( .A1(n8544), .A2(n10160), .ZN(n8551) );
  INV_X1 U10124 ( .A(n8545), .ZN(n8546) );
  NAND2_X1 U10125 ( .A1(n8547), .A2(n8546), .ZN(n8557) );
  XNOR2_X1 U10126 ( .A(n8562), .B(P2_REG1_REG_18__SCAN_IN), .ZN(n8548) );
  XNOR2_X1 U10127 ( .A(n8557), .B(n8548), .ZN(n8549) );
  NAND2_X1 U10128 ( .A1(n8549), .A2(n10129), .ZN(n8550) );
  NAND4_X1 U10129 ( .A1(n8553), .A2(n8552), .A3(n8551), .A4(n8550), .ZN(
        P2_U3200) );
  XNOR2_X1 U10130 ( .A(n8558), .B(P2_REG2_REG_19__SCAN_IN), .ZN(n8565) );
  INV_X1 U10131 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8941) );
  INV_X1 U10132 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8804) );
  NAND2_X1 U10133 ( .A1(n8562), .A2(n8804), .ZN(n8556) );
  AOI22_X1 U10134 ( .A1(n8557), .A2(n8556), .B1(P2_REG1_REG_18__SCAN_IN), .B2(
        n4523), .ZN(n8560) );
  XNOR2_X1 U10135 ( .A(n8558), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n8566) );
  INV_X1 U10136 ( .A(n8566), .ZN(n8559) );
  XNOR2_X1 U10137 ( .A(n8560), .B(n8559), .ZN(n8576) );
  OAI21_X1 U10138 ( .B1(n8563), .B2(n8562), .A(n8561), .ZN(n8569) );
  MUX2_X1 U10139 ( .A(n8566), .B(n8565), .S(n8564), .Z(n8567) );
  INV_X1 U10140 ( .A(n8567), .ZN(n8568) );
  XNOR2_X1 U10141 ( .A(n8569), .B(n8568), .ZN(n8571) );
  OAI21_X1 U10142 ( .B1(n10164), .B2(n8573), .A(n8572), .ZN(n8574) );
  AOI21_X1 U10143 ( .B1(n10142), .B2(P2_ADDR_REG_19__SCAN_IN), .A(n8574), .ZN(
        n8575) );
  OAI21_X1 U10144 ( .B1(n8820), .B2(n8579), .A(n10186), .ZN(n8582) );
  NAND2_X1 U10145 ( .A1(n10187), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n8580) );
  OAI211_X1 U10146 ( .C1(n8763), .C2(n8581), .A(n8582), .B(n8580), .ZN(
        P2_U3202) );
  NAND2_X1 U10147 ( .A1(n8823), .A2(n10181), .ZN(n8583) );
  OAI211_X1 U10148 ( .C1(n10186), .C2(n8584), .A(n8583), .B(n8582), .ZN(
        P2_U3203) );
  XOR2_X1 U10149 ( .A(n8585), .B(n8586), .Z(n8831) );
  INV_X1 U10150 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n8593) );
  XNOR2_X1 U10151 ( .A(n8587), .B(n8586), .ZN(n8592) );
  MUX2_X1 U10152 ( .A(n8593), .B(n8827), .S(n10186), .Z(n8596) );
  AOI22_X1 U10153 ( .A1(n8828), .A2(n10181), .B1(n10183), .B2(n8594), .ZN(
        n8595) );
  XNOR2_X1 U10154 ( .A(n8598), .B(n8597), .ZN(n8837) );
  INV_X1 U10155 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n8603) );
  MUX2_X1 U10156 ( .A(n8603), .B(n8832), .S(n10186), .Z(n8606) );
  AOI22_X1 U10157 ( .A1(n8834), .A2(n10181), .B1(n10183), .B2(n8604), .ZN(
        n8605) );
  XNOR2_X1 U10158 ( .A(n8607), .B(n8608), .ZN(n8843) );
  INV_X1 U10159 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n8613) );
  MUX2_X1 U10160 ( .A(n8613), .B(n8838), .S(n10186), .Z(n8616) );
  AOI22_X1 U10161 ( .A1(n8840), .A2(n10181), .B1(n10183), .B2(n8614), .ZN(
        n8615) );
  OAI211_X1 U10162 ( .C1(n8843), .C2(n8747), .A(n8616), .B(n8615), .ZN(
        P2_U3207) );
  NOR2_X1 U10163 ( .A1(n8846), .A2(n8628), .ZN(n8622) );
  XNOR2_X1 U10164 ( .A(n8618), .B(n8617), .ZN(n8619) );
  OAI222_X1 U10165 ( .A1(n8737), .A2(n8621), .B1(n8739), .B2(n8620), .C1(n8753), .C2(n8619), .ZN(n8844) );
  AOI211_X1 U10166 ( .C1(n10183), .C2(n8623), .A(n8622), .B(n8844), .ZN(n8627)
         );
  XNOR2_X1 U10167 ( .A(n8625), .B(n8624), .ZN(n8776) );
  AOI22_X1 U10168 ( .A1(n8776), .A2(n10182), .B1(P2_REG2_REG_25__SCAN_IN), 
        .B2(n10187), .ZN(n8626) );
  OAI21_X1 U10169 ( .B1(n8627), .B2(n10187), .A(n8626), .ZN(P2_U3208) );
  NOR2_X1 U10170 ( .A1(n8781), .A2(n8628), .ZN(n8633) );
  XOR2_X1 U10171 ( .A(n8629), .B(n8636), .Z(n8630) );
  OAI222_X1 U10172 ( .A1(n8739), .A2(n8632), .B1(n8737), .B2(n8631), .C1(n8753), .C2(n8630), .ZN(n8850) );
  AOI211_X1 U10173 ( .C1(n10183), .C2(n8634), .A(n8633), .B(n8850), .ZN(n8638)
         );
  XNOR2_X1 U10174 ( .A(n8635), .B(n8636), .ZN(n8779) );
  AOI22_X1 U10175 ( .A1(n8779), .A2(n10182), .B1(P2_REG2_REG_24__SCAN_IN), 
        .B2(n10187), .ZN(n8637) );
  OAI21_X1 U10176 ( .B1(n8638), .B2(n10187), .A(n8637), .ZN(P2_U3209) );
  XOR2_X1 U10177 ( .A(n8640), .B(n8639), .Z(n8862) );
  INV_X1 U10178 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n8644) );
  XNOR2_X1 U10179 ( .A(n8641), .B(n8640), .ZN(n8643) );
  AOI222_X1 U10180 ( .A1(n10178), .A2(n8643), .B1(n8642), .B2(n10173), .C1(
        n8671), .C2(n10175), .ZN(n8857) );
  MUX2_X1 U10181 ( .A(n8644), .B(n8857), .S(n10186), .Z(n8647) );
  AOI22_X1 U10182 ( .A1(n8859), .A2(n10181), .B1(n10183), .B2(n8645), .ZN(
        n8646) );
  OAI211_X1 U10183 ( .C1(n8862), .C2(n8747), .A(n8647), .B(n8646), .ZN(
        P2_U3210) );
  OR2_X1 U10184 ( .A1(n8683), .A2(n8684), .ZN(n8685) );
  AOI21_X1 U10185 ( .B1(n8685), .B2(n8667), .A(n8668), .ZN(n8666) );
  NAND2_X1 U10186 ( .A1(n8658), .A2(n8648), .ZN(n8650) );
  OAI21_X1 U10187 ( .B1(n8666), .B2(n8650), .A(n8649), .ZN(n8652) );
  AOI222_X1 U10188 ( .A1(n10178), .A2(n8652), .B1(n8688), .B2(n10175), .C1(
        n8651), .C2(n10173), .ZN(n8791) );
  INV_X1 U10189 ( .A(n8653), .ZN(n8656) );
  INV_X1 U10190 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n8654) );
  OAI22_X1 U10191 ( .A1(n8656), .A2(n8655), .B1(n10186), .B2(n8654), .ZN(n8657) );
  AOI21_X1 U10192 ( .B1(n8787), .B2(n10181), .A(n8657), .ZN(n8661) );
  OR2_X1 U10193 ( .A1(n8659), .A2(n8658), .ZN(n8789) );
  NAND3_X1 U10194 ( .A1(n8789), .A2(n10182), .A3(n8788), .ZN(n8660) );
  OAI211_X1 U10195 ( .C1(n8791), .C2(n10187), .A(n8661), .B(n8660), .ZN(
        P2_U3211) );
  NAND2_X1 U10196 ( .A1(n8662), .A2(n8663), .ZN(n8665) );
  XNOR2_X1 U10197 ( .A(n8665), .B(n8664), .ZN(n8869) );
  INV_X1 U10198 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n8673) );
  INV_X1 U10199 ( .A(n8666), .ZN(n8670) );
  NAND3_X1 U10200 ( .A1(n8685), .A2(n8668), .A3(n8667), .ZN(n8669) );
  NAND2_X1 U10201 ( .A1(n8670), .A2(n8669), .ZN(n8672) );
  AOI222_X1 U10202 ( .A1(n10178), .A2(n8672), .B1(n8699), .B2(n10175), .C1(
        n8671), .C2(n10173), .ZN(n8864) );
  MUX2_X1 U10203 ( .A(n8673), .B(n8864), .S(n10186), .Z(n8676) );
  AOI22_X1 U10204 ( .A1(n8866), .A2(n10181), .B1(n10183), .B2(n8674), .ZN(
        n8675) );
  OAI211_X1 U10205 ( .C1(n8869), .C2(n8747), .A(n8676), .B(n8675), .ZN(
        P2_U3212) );
  NAND2_X1 U10206 ( .A1(n8678), .A2(n8677), .ZN(n8709) );
  NOR2_X1 U10207 ( .A1(n8709), .A2(n8708), .ZN(n8711) );
  OAI21_X1 U10208 ( .B1(n8711), .B2(n8681), .A(n8680), .ZN(n8682) );
  XOR2_X1 U10209 ( .A(n8684), .B(n8682), .Z(n8875) );
  INV_X1 U10210 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n8690) );
  INV_X1 U10211 ( .A(n8683), .ZN(n8686) );
  OAI21_X1 U10212 ( .B1(n8686), .B2(n6561), .A(n8685), .ZN(n8689) );
  AOI222_X1 U10213 ( .A1(n10178), .A2(n8689), .B1(n8688), .B2(n10173), .C1(
        n8687), .C2(n10175), .ZN(n8870) );
  MUX2_X1 U10214 ( .A(n8690), .B(n8870), .S(n10186), .Z(n8693) );
  AOI22_X1 U10215 ( .A1(n8872), .A2(n10181), .B1(n8691), .B2(n10183), .ZN(
        n8692) );
  OAI211_X1 U10216 ( .C1(n8875), .C2(n8747), .A(n8693), .B(n8692), .ZN(
        P2_U3213) );
  INV_X1 U10217 ( .A(n8694), .ZN(n8695) );
  NOR2_X1 U10218 ( .A1(n8711), .A2(n8695), .ZN(n8696) );
  XNOR2_X1 U10219 ( .A(n8696), .B(n8697), .ZN(n8881) );
  INV_X1 U10220 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n8701) );
  XNOR2_X1 U10221 ( .A(n8698), .B(n8697), .ZN(n8700) );
  AOI222_X1 U10222 ( .A1(n10178), .A2(n8700), .B1(n8699), .B2(n10173), .C1(
        n8725), .C2(n10175), .ZN(n8876) );
  MUX2_X1 U10223 ( .A(n8701), .B(n8876), .S(n10186), .Z(n8704) );
  AOI22_X1 U10224 ( .A1(n8878), .A2(n10181), .B1(n10183), .B2(n8702), .ZN(
        n8703) );
  OAI211_X1 U10225 ( .C1(n8881), .C2(n8747), .A(n8704), .B(n8703), .ZN(
        P2_U3214) );
  XNOR2_X1 U10226 ( .A(n8705), .B(n8708), .ZN(n8706) );
  OAI222_X1 U10227 ( .A1(n8737), .A2(n8740), .B1(n8739), .B2(n8707), .C1(n8706), .C2(n8753), .ZN(n8802) );
  AND2_X1 U10228 ( .A1(n8709), .A2(n8708), .ZN(n8710) );
  AOI22_X1 U10229 ( .A1(n10187), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n10183), 
        .B2(n8712), .ZN(n8714) );
  NAND2_X1 U10230 ( .A1(n8803), .A2(n10181), .ZN(n8713) );
  OAI211_X1 U10231 ( .C1(n8885), .C2(n8747), .A(n8714), .B(n8713), .ZN(n8715)
         );
  AOI21_X1 U10232 ( .B1(n8802), .B2(n10186), .A(n8715), .ZN(n8716) );
  INV_X1 U10233 ( .A(n8716), .ZN(P2_U3215) );
  XNOR2_X1 U10234 ( .A(n8717), .B(n8721), .ZN(n8890) );
  INV_X1 U10235 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8728) );
  NAND2_X1 U10236 ( .A1(n8719), .A2(n8718), .ZN(n8733) );
  NAND2_X1 U10237 ( .A1(n8733), .A2(n8734), .ZN(n8742) );
  NAND3_X1 U10238 ( .A1(n8742), .A2(n8721), .A3(n8720), .ZN(n8723) );
  NAND3_X1 U10239 ( .A1(n8723), .A2(n10178), .A3(n8722), .ZN(n8727) );
  AOI22_X1 U10240 ( .A1(n8725), .A2(n10173), .B1(n10175), .B2(n8724), .ZN(
        n8726) );
  MUX2_X1 U10241 ( .A(n8728), .B(n8886), .S(n10186), .Z(n8731) );
  AOI22_X1 U10242 ( .A1(n6552), .A2(n10181), .B1(n10183), .B2(n8729), .ZN(
        n8730) );
  OAI211_X1 U10243 ( .C1(n8890), .C2(n8747), .A(n8731), .B(n8730), .ZN(
        P2_U3216) );
  XOR2_X1 U10244 ( .A(n8732), .B(n8734), .Z(n8897) );
  INV_X1 U10245 ( .A(n8733), .ZN(n8736) );
  INV_X1 U10246 ( .A(n8734), .ZN(n8735) );
  AOI21_X1 U10247 ( .B1(n8736), .B2(n8735), .A(n8753), .ZN(n8743) );
  OAI22_X1 U10248 ( .A1(n8740), .A2(n8739), .B1(n8738), .B2(n8737), .ZN(n8741)
         );
  AOI21_X1 U10249 ( .B1(n8743), .B2(n8742), .A(n8741), .ZN(n8891) );
  MUX2_X1 U10250 ( .A(n9039), .B(n8891), .S(n10186), .Z(n8746) );
  AOI22_X1 U10251 ( .A1(n6553), .A2(n10181), .B1(n10183), .B2(n8744), .ZN(
        n8745) );
  OAI211_X1 U10252 ( .C1(n8897), .C2(n8747), .A(n8746), .B(n8745), .ZN(
        P2_U3217) );
  INV_X1 U10253 ( .A(n8748), .ZN(n8760) );
  XNOR2_X1 U10254 ( .A(n8749), .B(n8750), .ZN(n10190) );
  INV_X1 U10255 ( .A(n10190), .ZN(n8759) );
  XNOR2_X1 U10256 ( .A(n8751), .B(n8750), .ZN(n8754) );
  AOI22_X1 U10257 ( .A1(n4432), .A2(n10175), .B1(n10173), .B2(n10176), .ZN(
        n8752) );
  OAI21_X1 U10258 ( .B1(n8754), .B2(n8753), .A(n8752), .ZN(n8755) );
  AOI21_X1 U10259 ( .B1(n8756), .B2(n10190), .A(n8755), .ZN(n10192) );
  AOI22_X1 U10260 ( .A1(n10183), .A2(P2_REG3_REG_2__SCAN_IN), .B1(n8757), .B2(
        n10189), .ZN(n8758) );
  OAI211_X1 U10261 ( .C1(n8760), .C2(n8759), .A(n10192), .B(n8758), .ZN(n8761)
         );
  MUX2_X1 U10262 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n8761), .S(n10186), .Z(
        P2_U3231) );
  NAND2_X1 U10263 ( .A1(n8820), .A2(n10229), .ZN(n8765) );
  NAND2_X1 U10264 ( .A1(n10227), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n8762) );
  OAI211_X1 U10265 ( .C1(n8763), .C2(n8780), .A(n8765), .B(n8762), .ZN(
        P2_U3490) );
  INV_X1 U10266 ( .A(n8823), .ZN(n8766) );
  NAND2_X1 U10267 ( .A1(n10227), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n8764) );
  OAI211_X1 U10268 ( .C1(n8766), .C2(n8780), .A(n8765), .B(n8764), .ZN(
        P2_U3489) );
  INV_X1 U10269 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n8967) );
  NAND2_X1 U10270 ( .A1(n8828), .A2(n8810), .ZN(n8769) );
  MUX2_X1 U10271 ( .A(n8984), .B(n8832), .S(n10229), .Z(n8772) );
  NAND2_X1 U10272 ( .A1(n8834), .A2(n8810), .ZN(n8771) );
  INV_X1 U10273 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n8773) );
  MUX2_X1 U10274 ( .A(n8773), .B(n8838), .S(n10229), .Z(n8775) );
  NAND2_X1 U10275 ( .A1(n8840), .A2(n8810), .ZN(n8774) );
  MUX2_X1 U10276 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n8844), .S(n10229), .Z(
        n8778) );
  INV_X1 U10277 ( .A(n8776), .ZN(n8847) );
  OAI22_X1 U10278 ( .A1(n8847), .A2(n8813), .B1(n8846), .B2(n8780), .ZN(n8777)
         );
  OR2_X1 U10279 ( .A1(n8778), .A2(n8777), .ZN(P2_U3484) );
  MUX2_X1 U10280 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n8850), .S(n10229), .Z(
        n8783) );
  INV_X1 U10281 ( .A(n8779), .ZN(n8856) );
  OAI22_X1 U10282 ( .A1(n8856), .A2(n8813), .B1(n8781), .B2(n8780), .ZN(n8782)
         );
  OR2_X1 U10283 ( .A1(n8783), .A2(n8782), .ZN(P2_U3483) );
  INV_X1 U10284 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n8784) );
  MUX2_X1 U10285 ( .A(n8784), .B(n8857), .S(n10229), .Z(n8786) );
  NAND2_X1 U10286 ( .A1(n8859), .A2(n8810), .ZN(n8785) );
  OAI211_X1 U10287 ( .C1(n8862), .C2(n8813), .A(n8786), .B(n8785), .ZN(
        P2_U3482) );
  INV_X1 U10288 ( .A(n8787), .ZN(n8793) );
  NAND3_X1 U10289 ( .A1(n8789), .A2(n8788), .A3(n10201), .ZN(n8790) );
  OAI211_X1 U10290 ( .C1(n8793), .C2(n8792), .A(n8791), .B(n8790), .ZN(n8863)
         );
  MUX2_X1 U10291 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n8863), .S(n10229), .Z(
        P2_U3481) );
  MUX2_X1 U10292 ( .A(n8794), .B(n8864), .S(n10229), .Z(n8796) );
  NAND2_X1 U10293 ( .A1(n8866), .A2(n8810), .ZN(n8795) );
  OAI211_X1 U10294 ( .C1(n8813), .C2(n8869), .A(n8796), .B(n8795), .ZN(
        P2_U3480) );
  INV_X1 U10295 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n8797) );
  MUX2_X1 U10296 ( .A(n8797), .B(n8870), .S(n10229), .Z(n8799) );
  NAND2_X1 U10297 ( .A1(n8872), .A2(n8810), .ZN(n8798) );
  OAI211_X1 U10298 ( .C1(n8813), .C2(n8875), .A(n8799), .B(n8798), .ZN(
        P2_U3479) );
  MUX2_X1 U10299 ( .A(n9009), .B(n8876), .S(n10229), .Z(n8801) );
  NAND2_X1 U10300 ( .A1(n8878), .A2(n8810), .ZN(n8800) );
  OAI211_X1 U10301 ( .C1(n8881), .C2(n8813), .A(n8801), .B(n8800), .ZN(
        P2_U3478) );
  AOI21_X1 U10302 ( .B1(n10216), .B2(n8803), .A(n8802), .ZN(n8882) );
  MUX2_X1 U10303 ( .A(n8804), .B(n8882), .S(n10229), .Z(n8805) );
  OAI21_X1 U10304 ( .B1(n8813), .B2(n8885), .A(n8805), .ZN(P2_U3477) );
  INV_X1 U10305 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n8806) );
  MUX2_X1 U10306 ( .A(n8806), .B(n8886), .S(n10229), .Z(n8808) );
  NAND2_X1 U10307 ( .A1(n6552), .A2(n8810), .ZN(n8807) );
  OAI211_X1 U10308 ( .C1(n8890), .C2(n8813), .A(n8808), .B(n8807), .ZN(
        P2_U3476) );
  MUX2_X1 U10309 ( .A(n8809), .B(n8891), .S(n10229), .Z(n8812) );
  NAND2_X1 U10310 ( .A1(n6553), .A2(n8810), .ZN(n8811) );
  OAI211_X1 U10311 ( .C1(n8897), .C2(n8813), .A(n8812), .B(n8811), .ZN(
        P2_U3475) );
  AOI22_X1 U10312 ( .A1(n8815), .A2(n10201), .B1(n10216), .B2(n8814), .ZN(
        n8816) );
  NAND2_X1 U10313 ( .A1(n8817), .A2(n8816), .ZN(n8898) );
  MUX2_X1 U10314 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n8898), .S(n10229), .Z(
        P2_U3474) );
  MUX2_X1 U10315 ( .A(n8818), .B(P2_REG1_REG_0__SCAN_IN), .S(n10227), .Z(
        P2_U3459) );
  NAND2_X1 U10316 ( .A1(n8819), .A2(n8893), .ZN(n8821) );
  NAND2_X1 U10317 ( .A1(n8820), .A2(n10217), .ZN(n8824) );
  OAI211_X1 U10318 ( .C1(n10217), .C2(n8822), .A(n8821), .B(n8824), .ZN(
        P2_U3458) );
  NAND2_X1 U10319 ( .A1(n8823), .A2(n8893), .ZN(n8825) );
  OAI211_X1 U10320 ( .C1(n10217), .C2(n8826), .A(n8825), .B(n8824), .ZN(
        P2_U3457) );
  MUX2_X1 U10321 ( .A(n9028), .B(n8827), .S(n10217), .Z(n8830) );
  NAND2_X1 U10322 ( .A1(n8828), .A2(n8893), .ZN(n8829) );
  INV_X1 U10323 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n8833) );
  MUX2_X1 U10324 ( .A(n8833), .B(n8832), .S(n10217), .Z(n8836) );
  NAND2_X1 U10325 ( .A1(n8834), .A2(n8893), .ZN(n8835) );
  MUX2_X1 U10326 ( .A(n8839), .B(n8838), .S(n10217), .Z(n8842) );
  NAND2_X1 U10327 ( .A1(n8840), .A2(n8893), .ZN(n8841) );
  MUX2_X1 U10328 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n8844), .S(n10217), .Z(
        n8849) );
  OAI22_X1 U10329 ( .A1(n8847), .A2(n8896), .B1(n8846), .B2(n8845), .ZN(n8848)
         );
  OR2_X1 U10330 ( .A1(n8849), .A2(n8848), .ZN(P2_U3452) );
  INV_X1 U10331 ( .A(n8850), .ZN(n8851) );
  MUX2_X1 U10332 ( .A(n8852), .B(n8851), .S(n10217), .Z(n8855) );
  NAND2_X1 U10333 ( .A1(n8853), .A2(n8893), .ZN(n8854) );
  OAI211_X1 U10334 ( .C1(n8856), .C2(n8896), .A(n8855), .B(n8854), .ZN(
        P2_U3451) );
  MUX2_X1 U10335 ( .A(n8858), .B(n8857), .S(n10217), .Z(n8861) );
  NAND2_X1 U10336 ( .A1(n8859), .A2(n8893), .ZN(n8860) );
  OAI211_X1 U10337 ( .C1(n8862), .C2(n8896), .A(n8861), .B(n8860), .ZN(
        P2_U3450) );
  MUX2_X1 U10338 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n8863), .S(n10217), .Z(
        P2_U3449) );
  INV_X1 U10339 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n8865) );
  MUX2_X1 U10340 ( .A(n8865), .B(n8864), .S(n10217), .Z(n8868) );
  NAND2_X1 U10341 ( .A1(n8866), .A2(n8893), .ZN(n8867) );
  OAI211_X1 U10342 ( .C1(n8869), .C2(n8896), .A(n8868), .B(n8867), .ZN(
        P2_U3448) );
  MUX2_X1 U10343 ( .A(n8871), .B(n8870), .S(n10217), .Z(n8874) );
  NAND2_X1 U10344 ( .A1(n8872), .A2(n8893), .ZN(n8873) );
  OAI211_X1 U10345 ( .C1(n8875), .C2(n8896), .A(n8874), .B(n8873), .ZN(
        P2_U3447) );
  INV_X1 U10346 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n8877) );
  MUX2_X1 U10347 ( .A(n8877), .B(n8876), .S(n10217), .Z(n8880) );
  NAND2_X1 U10348 ( .A1(n8878), .A2(n8893), .ZN(n8879) );
  OAI211_X1 U10349 ( .C1(n8881), .C2(n8896), .A(n8880), .B(n8879), .ZN(
        P2_U3446) );
  INV_X1 U10350 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n8883) );
  MUX2_X1 U10351 ( .A(n8883), .B(n8882), .S(n10217), .Z(n8884) );
  OAI21_X1 U10352 ( .B1(n8885), .B2(n8896), .A(n8884), .ZN(P2_U3444) );
  INV_X1 U10353 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n8887) );
  MUX2_X1 U10354 ( .A(n8887), .B(n8886), .S(n10217), .Z(n8889) );
  NAND2_X1 U10355 ( .A1(n6552), .A2(n8893), .ZN(n8888) );
  OAI211_X1 U10356 ( .C1(n8890), .C2(n8896), .A(n8889), .B(n8888), .ZN(
        P2_U3441) );
  MUX2_X1 U10357 ( .A(n8892), .B(n8891), .S(n10217), .Z(n8895) );
  NAND2_X1 U10358 ( .A1(n6553), .A2(n8893), .ZN(n8894) );
  OAI211_X1 U10359 ( .C1(n8897), .C2(n8896), .A(n8895), .B(n8894), .ZN(
        P2_U3438) );
  MUX2_X1 U10360 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n8898), .S(n10217), .Z(
        P2_U3435) );
  NOR4_X1 U10361 ( .A1(n4908), .A2(P2_IR_REG_30__SCAN_IN), .A3(P2_U3151), .A4(
        n5900), .ZN(n8899) );
  AOI21_X1 U10362 ( .B1(n8900), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n8899), .ZN(
        n8901) );
  OAI21_X1 U10363 ( .B1(n9960), .B2(n9059), .A(n8901), .ZN(P2_U3264) );
  OAI222_X1 U10364 ( .A1(n8905), .A2(n8978), .B1(n9059), .B2(n8903), .C1(
        P2_U3151), .C2(n8902), .ZN(P2_U3265) );
  INV_X1 U10365 ( .A(n8904), .ZN(n9962) );
  OAI222_X1 U10366 ( .A1(n9059), .A2(n9962), .B1(n8907), .B2(P2_U3151), .C1(
        n8906), .C2(n8905), .ZN(P2_U3266) );
  NAND2_X1 U10367 ( .A1(n8909), .A2(n8908), .ZN(n8911) );
  OAI211_X1 U10368 ( .C1(n8912), .C2(n8905), .A(n8911), .B(n8910), .ZN(
        P2_U3267) );
  NAND4_X1 U10369 ( .A1(P2_D_REG_1__SCAN_IN), .A2(P1_REG2_REG_26__SCAN_IN), 
        .A3(P2_ADDR_REG_6__SCAN_IN), .A4(n8941), .ZN(n8930) );
  NAND4_X1 U10370 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_REG3_REG_27__SCAN_IN), .A4(P2_REG1_REG_22__SCAN_IN), .ZN(n8929) );
  NOR3_X1 U10371 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(P1_REG1_REG_17__SCAN_IN), 
        .A3(P2_REG2_REG_7__SCAN_IN), .ZN(n8913) );
  NAND4_X1 U10372 ( .A1(n8915), .A2(P1_REG2_REG_22__SCAN_IN), .A3(n8914), .A4(
        n8913), .ZN(n8928) );
  NAND3_X1 U10373 ( .A1(P1_REG2_REG_7__SCAN_IN), .A2(P2_REG0_REG_5__SCAN_IN), 
        .A3(n9039), .ZN(n8918) );
  NAND4_X1 U10374 ( .A1(P1_REG1_REG_13__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), 
        .A3(n9042), .A4(n9041), .ZN(n8917) );
  NAND4_X1 U10375 ( .A1(P2_D_REG_5__SCAN_IN), .A2(P1_REG0_REG_20__SCAN_IN), 
        .A3(P2_REG1_REG_8__SCAN_IN), .A4(n9028), .ZN(n8916) );
  NOR4_X1 U10376 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(n8918), .A3(n8917), .A4(
        n8916), .ZN(n8926) );
  NAND4_X1 U10377 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P1_REG0_REG_24__SCAN_IN), 
        .A3(n8989), .A4(n8978), .ZN(n8921) );
  NAND4_X1 U10378 ( .A1(P1_ADDR_REG_19__SCAN_IN), .A2(P1_D_REG_18__SCAN_IN), 
        .A3(P1_DATAO_REG_14__SCAN_IN), .A4(n9017), .ZN(n8920) );
  NAND4_X1 U10379 ( .A1(P2_DATAO_REG_0__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), 
        .A3(P2_REG3_REG_14__SCAN_IN), .A4(P2_REG0_REG_1__SCAN_IN), .ZN(n8919)
         );
  NOR3_X1 U10380 ( .A1(n8921), .A2(n8920), .A3(n8919), .ZN(n8925) );
  NOR4_X1 U10381 ( .A1(n9008), .A2(P2_REG3_REG_26__SCAN_IN), .A3(
        P2_DATAO_REG_22__SCAN_IN), .A4(P2_REG1_REG_19__SCAN_IN), .ZN(n8924) );
  NOR4_X1 U10382 ( .A1(n8922), .A2(P2_REG1_REG_21__SCAN_IN), .A3(
        P1_REG3_REG_6__SCAN_IN), .A4(P1_REG3_REG_21__SCAN_IN), .ZN(n8923) );
  NAND4_X1 U10383 ( .A1(n8926), .A2(n8925), .A3(n8924), .A4(n8923), .ZN(n8927)
         );
  NOR4_X1 U10384 ( .A1(n8930), .A2(n8929), .A3(n8928), .A4(n8927), .ZN(n9056)
         );
  NAND4_X1 U10385 ( .A1(P1_DATAO_REG_25__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), 
        .A3(P2_REG1_REG_27__SCAN_IN), .A4(n8981), .ZN(n8931) );
  NOR3_X1 U10386 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(n8931), .A3(
        P2_ADDR_REG_10__SCAN_IN), .ZN(n8932) );
  NAND3_X1 U10387 ( .A1(n8932), .A2(SI_10_), .A3(n8967), .ZN(n8938) );
  INV_X1 U10388 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n8933) );
  NAND4_X1 U10389 ( .A1(n8934), .A2(n8933), .A3(P1_REG2_REG_0__SCAN_IN), .A4(
        P2_REG3_REG_20__SCAN_IN), .ZN(n8937) );
  NAND4_X1 U10390 ( .A1(n8935), .A2(n8965), .A3(P2_REG1_REG_31__SCAN_IN), .A4(
        P1_REG2_REG_20__SCAN_IN), .ZN(n8936) );
  NOR3_X1 U10391 ( .A1(n8938), .A2(n8937), .A3(n8936), .ZN(n9055) );
  AOI22_X1 U10392 ( .A1(n7472), .A2(keyinput9), .B1(n5139), .B2(keyinput1), 
        .ZN(n8939) );
  OAI221_X1 U10393 ( .B1(n7472), .B2(keyinput9), .C1(n5139), .C2(keyinput1), 
        .A(n8939), .ZN(n8952) );
  INV_X1 U10394 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n8942) );
  AOI22_X1 U10395 ( .A1(n8942), .A2(keyinput3), .B1(keyinput11), .B2(n8941), 
        .ZN(n8940) );
  OAI221_X1 U10396 ( .B1(n8942), .B2(keyinput3), .C1(n8941), .C2(keyinput11), 
        .A(n8940), .ZN(n8951) );
  INV_X1 U10397 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n8944) );
  INV_X1 U10398 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n9577) );
  AOI22_X1 U10399 ( .A1(n8944), .A2(keyinput22), .B1(keyinput7), .B2(n9577), 
        .ZN(n8943) );
  OAI221_X1 U10400 ( .B1(n8944), .B2(keyinput22), .C1(n9577), .C2(keyinput7), 
        .A(n8943), .ZN(n8949) );
  XNOR2_X1 U10401 ( .A(keyinput29), .B(n8945), .ZN(n8948) );
  XNOR2_X1 U10402 ( .A(n8946), .B(keyinput17), .ZN(n8947) );
  OR3_X1 U10403 ( .A1(n8949), .A2(n8948), .A3(n8947), .ZN(n8950) );
  NOR3_X1 U10404 ( .A1(n8952), .A2(n8951), .A3(n8950), .ZN(n8996) );
  AOI22_X1 U10405 ( .A1(n6309), .A2(keyinput60), .B1(n8954), .B2(keyinput5), 
        .ZN(n8953) );
  OAI221_X1 U10406 ( .B1(n6309), .B2(keyinput60), .C1(n8954), .C2(keyinput5), 
        .A(n8953), .ZN(n8963) );
  XOR2_X1 U10407 ( .A(P2_REG1_REG_31__SCAN_IN), .B(keyinput21), .Z(n8962) );
  XNOR2_X1 U10408 ( .A(n8955), .B(keyinput46), .ZN(n8961) );
  XNOR2_X1 U10409 ( .A(P2_REG1_REG_22__SCAN_IN), .B(keyinput59), .ZN(n8959) );
  XNOR2_X1 U10410 ( .A(SI_10_), .B(keyinput18), .ZN(n8958) );
  XNOR2_X1 U10411 ( .A(P1_REG1_REG_0__SCAN_IN), .B(keyinput27), .ZN(n8957) );
  XNOR2_X1 U10412 ( .A(P1_IR_REG_7__SCAN_IN), .B(keyinput47), .ZN(n8956) );
  NAND4_X1 U10413 ( .A1(n8959), .A2(n8958), .A3(n8957), .A4(n8956), .ZN(n8960)
         );
  NOR4_X1 U10414 ( .A1(n8963), .A2(n8962), .A3(n8961), .A4(n8960), .ZN(n8995)
         );
  INV_X1 U10415 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n8966) );
  AOI22_X1 U10416 ( .A1(n8966), .A2(keyinput10), .B1(keyinput50), .B2(n8965), 
        .ZN(n8964) );
  OAI221_X1 U10417 ( .B1(n8966), .B2(keyinput10), .C1(n8965), .C2(keyinput50), 
        .A(n8964), .ZN(n8975) );
  XNOR2_X1 U10418 ( .A(keyinput35), .B(n8967), .ZN(n8974) );
  XNOR2_X1 U10419 ( .A(P2_IR_REG_20__SCAN_IN), .B(keyinput61), .ZN(n8971) );
  XNOR2_X1 U10420 ( .A(P2_REG3_REG_20__SCAN_IN), .B(keyinput28), .ZN(n8970) );
  XNOR2_X1 U10421 ( .A(P2_IR_REG_7__SCAN_IN), .B(keyinput32), .ZN(n8969) );
  XNOR2_X1 U10422 ( .A(P1_REG1_REG_1__SCAN_IN), .B(keyinput2), .ZN(n8968) );
  NAND4_X1 U10423 ( .A1(n8971), .A2(n8970), .A3(n8969), .A4(n8968), .ZN(n8973)
         );
  XNOR2_X1 U10424 ( .A(n5270), .B(keyinput8), .ZN(n8972) );
  NOR4_X1 U10425 ( .A1(n8975), .A2(n8974), .A3(n8973), .A4(n8972), .ZN(n8994)
         );
  AOI22_X1 U10426 ( .A1(n8978), .A2(keyinput36), .B1(keyinput12), .B2(n8977), 
        .ZN(n8976) );
  OAI221_X1 U10427 ( .B1(n8978), .B2(keyinput36), .C1(n8977), .C2(keyinput12), 
        .A(n8976), .ZN(n8992) );
  AOI22_X1 U10428 ( .A1(n8981), .A2(keyinput54), .B1(keyinput58), .B2(n8980), 
        .ZN(n8979) );
  OAI221_X1 U10429 ( .B1(n8981), .B2(keyinput54), .C1(n8980), .C2(keyinput58), 
        .A(n8979), .ZN(n8988) );
  AOI22_X1 U10430 ( .A1(n8984), .A2(keyinput51), .B1(n8983), .B2(keyinput26), 
        .ZN(n8982) );
  OAI221_X1 U10431 ( .B1(n8984), .B2(keyinput51), .C1(n8983), .C2(keyinput26), 
        .A(n8982), .ZN(n8987) );
  XNOR2_X1 U10432 ( .A(keyinput6), .B(n8985), .ZN(n8986) );
  OR3_X1 U10433 ( .A1(n8988), .A2(n8987), .A3(n8986), .ZN(n8991) );
  XNOR2_X1 U10434 ( .A(n8989), .B(keyinput30), .ZN(n8990) );
  NOR3_X1 U10435 ( .A1(n8992), .A2(n8991), .A3(n8990), .ZN(n8993) );
  NAND4_X1 U10436 ( .A1(n8996), .A2(n8995), .A3(n8994), .A4(n8993), .ZN(n9054)
         );
  AOI22_X1 U10437 ( .A1(n6815), .A2(keyinput39), .B1(keyinput20), .B2(n8998), 
        .ZN(n8997) );
  OAI221_X1 U10438 ( .B1(n6815), .B2(keyinput39), .C1(n8998), .C2(keyinput20), 
        .A(n8997), .ZN(n9007) );
  AOI22_X1 U10439 ( .A1(n9000), .A2(keyinput13), .B1(keyinput37), .B2(n5932), 
        .ZN(n8999) );
  OAI221_X1 U10440 ( .B1(n9000), .B2(keyinput13), .C1(n5932), .C2(keyinput37), 
        .A(n8999), .ZN(n9006) );
  INV_X1 U10441 ( .A(P1_D_REG_17__SCAN_IN), .ZN(n10054) );
  AOI22_X1 U10442 ( .A1(n10054), .A2(keyinput42), .B1(keyinput53), .B2(n4585), 
        .ZN(n9001) );
  OAI221_X1 U10443 ( .B1(n10054), .B2(keyinput42), .C1(n4585), .C2(keyinput53), 
        .A(n9001), .ZN(n9005) );
  XNOR2_X1 U10444 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(keyinput40), .ZN(n9003) );
  XNOR2_X1 U10445 ( .A(P2_IR_REG_16__SCAN_IN), .B(keyinput43), .ZN(n9002) );
  NAND2_X1 U10446 ( .A1(n9003), .A2(n9002), .ZN(n9004) );
  NOR4_X1 U10447 ( .A1(n9007), .A2(n9006), .A3(n9005), .A4(n9004), .ZN(n9052)
         );
  INV_X1 U10448 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n9603) );
  XNOR2_X1 U10449 ( .A(n9603), .B(keyinput49), .ZN(n9012) );
  XNOR2_X1 U10450 ( .A(n9008), .B(keyinput19), .ZN(n9011) );
  XNOR2_X1 U10451 ( .A(n9009), .B(keyinput16), .ZN(n9010) );
  NOR3_X1 U10452 ( .A1(n9012), .A2(n9011), .A3(n9010), .ZN(n9015) );
  XNOR2_X1 U10453 ( .A(P1_REG3_REG_21__SCAN_IN), .B(keyinput0), .ZN(n9014) );
  XNOR2_X1 U10454 ( .A(P1_REG3_REG_6__SCAN_IN), .B(keyinput57), .ZN(n9013) );
  NAND3_X1 U10455 ( .A1(n9015), .A2(n9014), .A3(n9013), .ZN(n9021) );
  INV_X1 U10456 ( .A(P1_D_REG_18__SCAN_IN), .ZN(n10053) );
  AOI22_X1 U10457 ( .A1(n9017), .A2(keyinput4), .B1(n10053), .B2(keyinput33), 
        .ZN(n9016) );
  OAI221_X1 U10458 ( .B1(n9017), .B2(keyinput4), .C1(n10053), .C2(keyinput33), 
        .A(n9016), .ZN(n9020) );
  XNOR2_X1 U10459 ( .A(n9018), .B(keyinput63), .ZN(n9019) );
  NOR3_X1 U10460 ( .A1(n9021), .A2(n9020), .A3(n9019), .ZN(n9051) );
  AOI22_X1 U10461 ( .A1(n9024), .A2(keyinput48), .B1(n9023), .B2(keyinput14), 
        .ZN(n9022) );
  OAI221_X1 U10462 ( .B1(n9024), .B2(keyinput48), .C1(n9023), .C2(keyinput14), 
        .A(n9022), .ZN(n9035) );
  AOI22_X1 U10463 ( .A1(n4580), .A2(keyinput41), .B1(n9026), .B2(keyinput44), 
        .ZN(n9025) );
  OAI221_X1 U10464 ( .B1(n4580), .B2(keyinput41), .C1(n9026), .C2(keyinput44), 
        .A(n9025), .ZN(n9034) );
  AOI22_X1 U10465 ( .A1(n9029), .A2(keyinput31), .B1(keyinput34), .B2(n9028), 
        .ZN(n9027) );
  OAI221_X1 U10466 ( .B1(n9029), .B2(keyinput31), .C1(n9028), .C2(keyinput34), 
        .A(n9027), .ZN(n9033) );
  INV_X1 U10467 ( .A(P1_D_REG_29__SCAN_IN), .ZN(n10052) );
  AOI22_X1 U10468 ( .A1(n10052), .A2(keyinput55), .B1(keyinput56), .B2(n9031), 
        .ZN(n9030) );
  OAI221_X1 U10469 ( .B1(n10052), .B2(keyinput55), .C1(n9031), .C2(keyinput56), 
        .A(n9030), .ZN(n9032) );
  NOR4_X1 U10470 ( .A1(n9035), .A2(n9034), .A3(n9033), .A4(n9032), .ZN(n9050)
         );
  INV_X1 U10471 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n9527) );
  AOI22_X1 U10472 ( .A1(n9527), .A2(keyinput62), .B1(keyinput24), .B2(n9037), 
        .ZN(n9036) );
  OAI221_X1 U10473 ( .B1(n9527), .B2(keyinput62), .C1(n9037), .C2(keyinput24), 
        .A(n9036), .ZN(n9048) );
  INV_X1 U10474 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n10209) );
  AOI22_X1 U10475 ( .A1(n10209), .A2(keyinput38), .B1(n9039), .B2(keyinput52), 
        .ZN(n9038) );
  OAI221_X1 U10476 ( .B1(n10209), .B2(keyinput38), .C1(n9039), .C2(keyinput52), 
        .A(n9038), .ZN(n9047) );
  AOI22_X1 U10477 ( .A1(n9042), .A2(keyinput15), .B1(keyinput25), .B2(n9041), 
        .ZN(n9040) );
  OAI221_X1 U10478 ( .B1(n9042), .B2(keyinput15), .C1(n9041), .C2(keyinput25), 
        .A(n9040), .ZN(n9046) );
  XNOR2_X1 U10479 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(keyinput23), .ZN(n9044) );
  XNOR2_X1 U10480 ( .A(P2_REG1_REG_21__SCAN_IN), .B(keyinput45), .ZN(n9043) );
  NAND2_X1 U10481 ( .A1(n9044), .A2(n9043), .ZN(n9045) );
  NOR4_X1 U10482 ( .A1(n9048), .A2(n9047), .A3(n9046), .A4(n9045), .ZN(n9049)
         );
  NAND4_X1 U10483 ( .A1(n9052), .A2(n9051), .A3(n9050), .A4(n9049), .ZN(n9053)
         );
  AOI211_X1 U10484 ( .C1(n9056), .C2(n9055), .A(n9054), .B(n9053), .ZN(n9062)
         );
  OAI222_X1 U10485 ( .A1(n8905), .A2(n9060), .B1(n9059), .B2(n9058), .C1(
        P2_U3151), .C2(n4270), .ZN(n9061) );
  XOR2_X1 U10486 ( .A(n9062), .B(n9061), .Z(P2_U3292) );
  MUX2_X1 U10487 ( .A(n9063), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  XNOR2_X1 U10488 ( .A(n9065), .B(n9064), .ZN(n9066) );
  XNOR2_X1 U10489 ( .A(n9067), .B(n9066), .ZN(n9068) );
  NAND2_X1 U10490 ( .A1(n9068), .A2(n9326), .ZN(n9075) );
  NOR2_X1 U10491 ( .A1(n9069), .A2(n9329), .ZN(n9071) );
  NOR2_X1 U10492 ( .A1(n9218), .A2(n9626), .ZN(n9070) );
  OR2_X1 U10493 ( .A1(n9071), .A2(n9070), .ZN(n10004) );
  AOI22_X1 U10494 ( .A1(n9335), .A2(n10004), .B1(P1_REG3_REG_7__SCAN_IN), .B2(
        P1_U3086), .ZN(n9074) );
  NAND2_X1 U10495 ( .A1(n9348), .A2(n10007), .ZN(n9073) );
  NAND2_X1 U10496 ( .A1(n9343), .A2(n10006), .ZN(n9072) );
  NAND4_X1 U10497 ( .A1(n9075), .A2(n9074), .A3(n9073), .A4(n9072), .ZN(
        P1_U3213) );
  INV_X1 U10498 ( .A(n9076), .ZN(n9078) );
  NAND2_X1 U10499 ( .A1(n9078), .A2(n9077), .ZN(n9080) );
  XNOR2_X1 U10500 ( .A(n9080), .B(n9079), .ZN(n9088) );
  OAI22_X1 U10501 ( .A1(n9082), .A2(n9345), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9081), .ZN(n9085) );
  NOR2_X1 U10502 ( .A1(n9083), .A2(n9338), .ZN(n9084) );
  AOI211_X1 U10503 ( .C1(n9086), .C2(n9343), .A(n9085), .B(n9084), .ZN(n9087)
         );
  OAI21_X1 U10504 ( .B1(n9088), .B2(n9350), .A(n9087), .ZN(P1_U3215) );
  OAI21_X1 U10505 ( .B1(n9089), .B2(n4989), .A(n9090), .ZN(n9283) );
  NOR2_X1 U10506 ( .A1(n9283), .A2(n9284), .ZN(n9282) );
  INV_X1 U10507 ( .A(n9090), .ZN(n9091) );
  NOR3_X1 U10508 ( .A1(n9282), .A2(n9092), .A3(n9091), .ZN(n9093) );
  OAI21_X1 U10509 ( .B1(n9093), .B2(n4931), .A(n9326), .ZN(n9100) );
  OAI22_X1 U10510 ( .A1(n9095), .A2(n9329), .B1(n9094), .B2(n9626), .ZN(n9715)
         );
  INV_X1 U10511 ( .A(n9709), .ZN(n9097) );
  OAI22_X1 U10512 ( .A1(n9097), .A2(n9332), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9096), .ZN(n9098) );
  AOI21_X1 U10513 ( .B1(n9715), .B2(n9335), .A(n9098), .ZN(n9099) );
  INV_X1 U10514 ( .A(n9102), .ZN(n9107) );
  NOR2_X1 U10515 ( .A1(n9107), .A2(n9103), .ZN(n9179) );
  INV_X1 U10516 ( .A(n9179), .ZN(n9108) );
  INV_X1 U10517 ( .A(n9104), .ZN(n9105) );
  OAI21_X1 U10518 ( .B1(n9107), .B2(n9106), .A(n9105), .ZN(n9177) );
  NAND2_X1 U10519 ( .A1(n9108), .A2(n9177), .ZN(n9109) );
  XNOR2_X1 U10520 ( .A(n9109), .B(n9178), .ZN(n9116) );
  OAI22_X1 U10521 ( .A1(n9111), .A2(n9345), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9110), .ZN(n9113) );
  NOR2_X1 U10522 ( .A1(n10104), .A2(n9338), .ZN(n9112) );
  AOI211_X1 U10523 ( .C1(n9114), .C2(n9343), .A(n9113), .B(n9112), .ZN(n9115)
         );
  OAI21_X1 U10524 ( .B1(n9116), .B2(n9350), .A(n9115), .ZN(P1_U3217) );
  XNOR2_X1 U10525 ( .A(n9166), .B(n9118), .ZN(n9303) );
  OAI22_X1 U10526 ( .A1(n9303), .A2(n9167), .B1(n9166), .B2(n9118), .ZN(n9122)
         );
  OR2_X1 U10527 ( .A1(n9120), .A2(n9119), .ZN(n9164) );
  NAND2_X1 U10528 ( .A1(n9262), .A2(n9164), .ZN(n9121) );
  XNOR2_X1 U10529 ( .A(n9122), .B(n9121), .ZN(n9128) );
  INV_X1 U10530 ( .A(n9773), .ZN(n9125) );
  OAI22_X1 U10531 ( .A1(n9123), .A2(n9329), .B1(n9232), .B2(n9626), .ZN(n9779)
         );
  AOI22_X1 U10532 ( .A1(n9779), .A2(n9335), .B1(P1_REG3_REG_19__SCAN_IN), .B2(
        P1_U3086), .ZN(n9124) );
  OAI21_X1 U10533 ( .B1(n9332), .B2(n9125), .A(n9124), .ZN(n9126) );
  AOI21_X1 U10534 ( .B1(n9893), .B2(n9348), .A(n9126), .ZN(n9127) );
  OAI21_X1 U10535 ( .B1(n9128), .B2(n9350), .A(n9127), .ZN(P1_U3219) );
  NAND2_X1 U10536 ( .A1(n9636), .A2(n7884), .ZN(n9131) );
  NAND2_X1 U10537 ( .A1(n9612), .A2(n9129), .ZN(n9130) );
  NAND2_X1 U10538 ( .A1(n9131), .A2(n9130), .ZN(n9133) );
  XNOR2_X1 U10539 ( .A(n9133), .B(n4278), .ZN(n9136) );
  AOI22_X1 U10540 ( .A1(n9636), .A2(n7904), .B1(n7930), .B2(n9612), .ZN(n9135)
         );
  XNOR2_X1 U10541 ( .A(n9136), .B(n9135), .ZN(n9143) );
  OR4_X2 U10542 ( .A1(n9137), .A2(n9142), .A3(n9143), .A4(n9350), .ZN(n9147)
         );
  NAND3_X1 U10543 ( .A1(n9137), .A2(n9326), .A3(n9143), .ZN(n9146) );
  INV_X1 U10544 ( .A(n9138), .ZN(n9140) );
  AOI22_X1 U10545 ( .A1(n9639), .A2(n9343), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3086), .ZN(n9139) );
  OAI21_X1 U10546 ( .B1(n9140), .B2(n9345), .A(n9139), .ZN(n9141) );
  AOI21_X1 U10547 ( .B1(n9636), .B2(n9348), .A(n9141), .ZN(n9145) );
  NAND3_X1 U10548 ( .A1(n9143), .A2(n9142), .A3(n9326), .ZN(n9144) );
  NAND4_X1 U10549 ( .A1(n9147), .A2(n9146), .A3(n9145), .A4(n9144), .ZN(
        P1_U3220) );
  NAND2_X1 U10550 ( .A1(n9149), .A2(n9148), .ZN(n9248) );
  XNOR2_X1 U10551 ( .A(n9248), .B(n9150), .ZN(n9151) );
  NOR2_X1 U10552 ( .A1(n9151), .A2(n9152), .ZN(n9249) );
  AOI21_X1 U10553 ( .B1(n9152), .B2(n9151), .A(n9249), .ZN(n9159) );
  NAND2_X1 U10554 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n9480) );
  NAND2_X1 U10555 ( .A1(n9343), .A2(n9153), .ZN(n9154) );
  OAI211_X1 U10556 ( .C1(n9155), .C2(n9345), .A(n9480), .B(n9154), .ZN(n9156)
         );
  AOI21_X1 U10557 ( .B1(n9157), .B2(n9348), .A(n9156), .ZN(n9158) );
  OAI21_X1 U10558 ( .B1(n9159), .B2(n9350), .A(n9158), .ZN(P1_U3221) );
  AOI22_X1 U10559 ( .A1(n9357), .A2(n9304), .B1(n9359), .B2(n9305), .ZN(n9741)
         );
  INV_X1 U10560 ( .A(n9160), .ZN(n9745) );
  AOI22_X1 U10561 ( .A1(n9745), .A2(n9343), .B1(P1_REG3_REG_21__SCAN_IN), .B2(
        P1_U3086), .ZN(n9161) );
  OAI21_X1 U10562 ( .B1(n9741), .B2(n9345), .A(n9161), .ZN(n9175) );
  INV_X1 U10563 ( .A(n9166), .ZN(n9163) );
  OAI21_X1 U10564 ( .B1(n9163), .B2(n9302), .A(n9162), .ZN(n9165) );
  OAI211_X1 U10565 ( .C1(n9167), .C2(n9166), .A(n9165), .B(n9164), .ZN(n9263)
         );
  AND2_X1 U10566 ( .A1(n9168), .A2(n9171), .ZN(n9261) );
  INV_X1 U10567 ( .A(n9169), .ZN(n9170) );
  NAND3_X1 U10568 ( .A1(n9260), .A2(n9171), .A3(n9170), .ZN(n9173) );
  AOI21_X1 U10569 ( .B1(n9173), .B2(n9172), .A(n9350), .ZN(n9174) );
  INV_X1 U10570 ( .A(n9176), .ZN(P1_U3223) );
  OAI21_X1 U10571 ( .B1(n9179), .B2(n9178), .A(n9177), .ZN(n9293) );
  NAND2_X1 U10572 ( .A1(n9180), .A2(n9181), .ZN(n9294) );
  NOR2_X1 U10573 ( .A1(n9293), .A2(n9294), .ZN(n9292) );
  INV_X1 U10574 ( .A(n9181), .ZN(n9183) );
  NOR3_X1 U10575 ( .A1(n9292), .A2(n9183), .A3(n9182), .ZN(n9184) );
  OAI21_X1 U10576 ( .B1(n9184), .B2(n4388), .A(n9326), .ZN(n9190) );
  OAI21_X1 U10577 ( .B1(n9186), .B2(n9345), .A(n9185), .ZN(n9187) );
  AOI21_X1 U10578 ( .B1(n9188), .B2(n9343), .A(n9187), .ZN(n9189) );
  OAI211_X1 U10579 ( .C1(n9191), .C2(n9338), .A(n9190), .B(n9189), .ZN(
        P1_U3224) );
  OAI21_X1 U10580 ( .B1(n9194), .B2(n9193), .A(n9192), .ZN(n9195) );
  NAND2_X1 U10581 ( .A1(n9195), .A2(n9326), .ZN(n9202) );
  OR2_X1 U10582 ( .A1(n9196), .A2(n9329), .ZN(n9198) );
  NAND2_X1 U10583 ( .A1(n9355), .A2(n9305), .ZN(n9197) );
  NAND2_X1 U10584 ( .A1(n9198), .A2(n9197), .ZN(n9682) );
  OAI22_X1 U10585 ( .A1(n9677), .A2(n9332), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9199), .ZN(n9200) );
  AOI21_X1 U10586 ( .B1(n9682), .B2(n9335), .A(n9200), .ZN(n9201) );
  OAI211_X1 U10587 ( .C1(n9680), .C2(n9338), .A(n9202), .B(n9201), .ZN(
        P1_U3225) );
  INV_X1 U10588 ( .A(n4443), .ZN(n9204) );
  NAND2_X1 U10589 ( .A1(n9205), .A2(n9204), .ZN(n9340) );
  INV_X1 U10590 ( .A(n9206), .ZN(n9341) );
  NOR2_X1 U10591 ( .A1(n9340), .A2(n9341), .ZN(n9339) );
  NOR2_X1 U10592 ( .A1(n9339), .A2(n4443), .ZN(n9210) );
  XNOR2_X1 U10593 ( .A(n9208), .B(n9207), .ZN(n9209) );
  NOR2_X1 U10594 ( .A1(n9210), .A2(n9209), .ZN(n9227) );
  AOI21_X1 U10595 ( .B1(n9210), .B2(n9209), .A(n9227), .ZN(n9214) );
  NOR2_X1 U10596 ( .A1(n9332), .A2(n9813), .ZN(n9212) );
  AOI22_X1 U10597 ( .A1(n9362), .A2(n9304), .B1(n9305), .B2(n9364), .ZN(n9821)
         );
  NAND2_X1 U10598 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9559) );
  OAI21_X1 U10599 ( .B1(n9821), .B2(n9345), .A(n9559), .ZN(n9211) );
  AOI211_X1 U10600 ( .C1(n9908), .C2(n9348), .A(n9212), .B(n9211), .ZN(n9213)
         );
  OAI21_X1 U10601 ( .B1(n9214), .B2(n9350), .A(n9213), .ZN(P1_U3226) );
  NOR2_X1 U10602 ( .A1(n4305), .A2(n4386), .ZN(n9216) );
  XNOR2_X1 U10603 ( .A(n9216), .B(n9215), .ZN(n9217) );
  NAND2_X1 U10604 ( .A1(n9217), .A2(n9326), .ZN(n9225) );
  NOR2_X1 U10605 ( .A1(n9218), .A2(n9329), .ZN(n9221) );
  NOR2_X1 U10606 ( .A1(n9219), .A2(n9626), .ZN(n9220) );
  OR2_X1 U10607 ( .A1(n9221), .A2(n9220), .ZN(n10016) );
  AOI22_X1 U10608 ( .A1(n9335), .A2(n10016), .B1(P1_REG3_REG_5__SCAN_IN), .B2(
        P1_U3086), .ZN(n9224) );
  NAND2_X1 U10609 ( .A1(n9348), .A2(n6425), .ZN(n9223) );
  NAND2_X1 U10610 ( .A1(n9343), .A2(n10018), .ZN(n9222) );
  NAND4_X1 U10611 ( .A1(n9225), .A2(n9224), .A3(n9223), .A4(n9222), .ZN(
        P1_U3227) );
  OAI21_X1 U10612 ( .B1(n9227), .B2(n4310), .A(n9226), .ZN(n9230) );
  NAND3_X1 U10613 ( .A1(n9230), .A2(n9326), .A3(n9229), .ZN(n9236) );
  OAI22_X1 U10614 ( .A1(n9232), .A2(n9329), .B1(n9231), .B2(n9626), .ZN(n9804)
         );
  NOR2_X1 U10615 ( .A1(n9233), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9575) );
  NOR2_X1 U10616 ( .A1(n9332), .A2(n9807), .ZN(n9234) );
  AOI211_X1 U10617 ( .C1(n9335), .C2(n9804), .A(n9575), .B(n9234), .ZN(n9235)
         );
  OAI211_X1 U10618 ( .C1(n9799), .C2(n9338), .A(n9236), .B(n9235), .ZN(
        P1_U3228) );
  NOR3_X1 U10619 ( .A1(n4931), .A2(n9238), .A3(n9237), .ZN(n9241) );
  INV_X1 U10620 ( .A(n9239), .ZN(n9240) );
  OAI21_X1 U10621 ( .B1(n9241), .B2(n9240), .A(n9326), .ZN(n9247) );
  NOR2_X1 U10622 ( .A1(n9286), .A2(n9626), .ZN(n9242) );
  AOI21_X1 U10623 ( .B1(n9354), .B2(n9304), .A(n9242), .ZN(n9693) );
  INV_X1 U10624 ( .A(n9693), .ZN(n9245) );
  OAI22_X1 U10625 ( .A1(n9698), .A2(n9332), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9243), .ZN(n9244) );
  AOI21_X1 U10626 ( .B1(n9245), .B2(n9335), .A(n9244), .ZN(n9246) );
  OAI211_X1 U10627 ( .C1(n9702), .C2(n9338), .A(n9247), .B(n9246), .ZN(
        P1_U3229) );
  INV_X1 U10628 ( .A(n9248), .ZN(n9251) );
  AOI21_X1 U10629 ( .B1(n9251), .B2(n9250), .A(n9249), .ZN(n9253) );
  OAI211_X1 U10630 ( .C1(n9253), .C2(n9252), .A(n9326), .B(n9102), .ZN(n9259)
         );
  OAI21_X1 U10631 ( .B1(n9255), .B2(n9345), .A(n9254), .ZN(n9256) );
  AOI21_X1 U10632 ( .B1(n9257), .B2(n9343), .A(n9256), .ZN(n9258) );
  OAI211_X1 U10633 ( .C1(n4948), .C2(n9338), .A(n9259), .B(n9258), .ZN(
        P1_U3231) );
  INV_X1 U10634 ( .A(n9888), .ZN(n9271) );
  INV_X1 U10635 ( .A(n9260), .ZN(n9265) );
  AOI21_X1 U10636 ( .B1(n9263), .B2(n9262), .A(n9261), .ZN(n9264) );
  OAI21_X1 U10637 ( .B1(n9265), .B2(n9264), .A(n9326), .ZN(n9270) );
  INV_X1 U10638 ( .A(n9762), .ZN(n9268) );
  AOI22_X1 U10639 ( .A1(n9358), .A2(n9304), .B1(n9305), .B2(n9360), .ZN(n9754)
         );
  OAI22_X1 U10640 ( .A1(n9754), .A2(n9345), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9266), .ZN(n9267) );
  AOI21_X1 U10641 ( .B1(n9268), .B2(n9343), .A(n9267), .ZN(n9269) );
  OAI211_X1 U10642 ( .C1(n9271), .C2(n9338), .A(n9270), .B(n9269), .ZN(
        P1_U3233) );
  OAI21_X1 U10643 ( .B1(n9274), .B2(n9273), .A(n9272), .ZN(n9275) );
  NAND2_X1 U10644 ( .A1(n9275), .A2(n9326), .ZN(n9280) );
  NAND2_X1 U10645 ( .A1(P1_U3086), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n9521) );
  OAI21_X1 U10646 ( .B1(n9276), .B2(n9345), .A(n9521), .ZN(n9277) );
  AOI21_X1 U10647 ( .B1(n9278), .B2(n9343), .A(n9277), .ZN(n9279) );
  OAI211_X1 U10648 ( .C1(n9281), .C2(n9338), .A(n9280), .B(n9279), .ZN(
        P1_U3234) );
  AOI21_X1 U10649 ( .B1(n9284), .B2(n9283), .A(n9282), .ZN(n9291) );
  OAI22_X1 U10650 ( .A1(n9286), .A2(n9329), .B1(n9285), .B2(n9626), .ZN(n9732)
         );
  OAI22_X1 U10651 ( .A1(n9722), .A2(n9332), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9287), .ZN(n9289) );
  NOR2_X1 U10652 ( .A1(n9725), .A2(n9338), .ZN(n9288) );
  AOI211_X1 U10653 ( .C1(n9335), .C2(n9732), .A(n9289), .B(n9288), .ZN(n9290)
         );
  OAI21_X1 U10654 ( .B1(n9291), .B2(n9350), .A(n9290), .ZN(P1_U3235) );
  AOI21_X1 U10655 ( .B1(n9294), .B2(n9293), .A(n9292), .ZN(n9301) );
  NAND2_X1 U10656 ( .A1(P1_U3086), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n9507) );
  NAND2_X1 U10657 ( .A1(n9343), .A2(n9295), .ZN(n9296) );
  OAI211_X1 U10658 ( .C1(n9297), .C2(n9345), .A(n9507), .B(n9296), .ZN(n9298)
         );
  AOI21_X1 U10659 ( .B1(n4857), .B2(n9348), .A(n9298), .ZN(n9300) );
  OAI21_X1 U10660 ( .B1(n9301), .B2(n9350), .A(n9300), .ZN(P1_U3236) );
  XNOR2_X1 U10661 ( .A(n9303), .B(n9302), .ZN(n9311) );
  NAND2_X1 U10662 ( .A1(n9360), .A2(n9304), .ZN(n9307) );
  NAND2_X1 U10663 ( .A1(n9362), .A2(n9305), .ZN(n9306) );
  NAND2_X1 U10664 ( .A1(n9307), .A2(n9306), .ZN(n9786) );
  AOI22_X1 U10665 ( .A1(n9786), .A2(n9335), .B1(P1_REG3_REG_18__SCAN_IN), .B2(
        P1_U3086), .ZN(n9308) );
  OAI21_X1 U10666 ( .B1(n9332), .B2(n9790), .A(n9308), .ZN(n9309) );
  AOI21_X1 U10667 ( .B1(n9898), .B2(n9348), .A(n9309), .ZN(n9310) );
  OAI21_X1 U10668 ( .B1(n9311), .B2(n9350), .A(n9310), .ZN(P1_U3238) );
  AOI21_X1 U10669 ( .B1(n9314), .B2(n9313), .A(n4468), .ZN(n9315) );
  OR2_X1 U10670 ( .A1(n9315), .A2(n9350), .ZN(n9321) );
  AOI22_X1 U10671 ( .A1(n9335), .A2(n9316), .B1(P1_REG3_REG_6__SCAN_IN), .B2(
        P1_U3086), .ZN(n9320) );
  NAND2_X1 U10672 ( .A1(n9348), .A2(n10083), .ZN(n9319) );
  NAND2_X1 U10673 ( .A1(n9343), .A2(n9317), .ZN(n9318) );
  NAND4_X1 U10674 ( .A1(n9321), .A2(n9320), .A3(n9319), .A4(n9318), .ZN(
        P1_U3239) );
  INV_X1 U10675 ( .A(n9192), .ZN(n9324) );
  OAI21_X1 U10676 ( .B1(n9324), .B2(n9323), .A(n9322), .ZN(n9327) );
  NAND3_X1 U10677 ( .A1(n9327), .A2(n9326), .A3(n9325), .ZN(n9337) );
  OAI22_X1 U10678 ( .A1(n9330), .A2(n9329), .B1(n9328), .B2(n9626), .ZN(n9667)
         );
  INV_X1 U10679 ( .A(n9670), .ZN(n9333) );
  OAI22_X1 U10680 ( .A1(n9333), .A2(n9332), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9331), .ZN(n9334) );
  AOI21_X1 U10681 ( .B1(n9667), .B2(n9335), .A(n9334), .ZN(n9336) );
  OAI211_X1 U10682 ( .C1(n9673), .C2(n9338), .A(n9337), .B(n9336), .ZN(
        P1_U3240) );
  AOI21_X1 U10683 ( .B1(n9341), .B2(n9340), .A(n9339), .ZN(n9351) );
  NAND2_X1 U10684 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9976) );
  NAND2_X1 U10685 ( .A1(n9343), .A2(n9342), .ZN(n9344) );
  OAI211_X1 U10686 ( .C1(n9346), .C2(n9345), .A(n9976), .B(n9344), .ZN(n9347)
         );
  AOI21_X1 U10687 ( .B1(n9914), .B2(n9348), .A(n9347), .ZN(n9349) );
  OAI21_X1 U10688 ( .B1(n9351), .B2(n9350), .A(n9349), .ZN(P1_U3241) );
  MUX2_X1 U10689 ( .A(n9352), .B(P1_DATAO_REG_31__SCAN_IN), .S(n9376), .Z(
        P1_U3585) );
  MUX2_X1 U10690 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9612), .S(P1_U3973), .Z(
        P1_U3582) );
  MUX2_X1 U10691 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9353), .S(P1_U3973), .Z(
        P1_U3581) );
  MUX2_X1 U10692 ( .A(n9354), .B(P1_DATAO_REG_25__SCAN_IN), .S(n9376), .Z(
        P1_U3579) );
  MUX2_X1 U10693 ( .A(n9355), .B(P1_DATAO_REG_24__SCAN_IN), .S(n9376), .Z(
        P1_U3578) );
  MUX2_X1 U10694 ( .A(n9356), .B(P1_DATAO_REG_23__SCAN_IN), .S(n9376), .Z(
        P1_U3577) );
  MUX2_X1 U10695 ( .A(n9357), .B(P1_DATAO_REG_22__SCAN_IN), .S(n9376), .Z(
        P1_U3576) );
  MUX2_X1 U10696 ( .A(n9358), .B(P1_DATAO_REG_21__SCAN_IN), .S(n9376), .Z(
        P1_U3575) );
  MUX2_X1 U10697 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9359), .S(P1_U3973), .Z(
        P1_U3574) );
  MUX2_X1 U10698 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9360), .S(P1_U3973), .Z(
        P1_U3573) );
  MUX2_X1 U10699 ( .A(n9361), .B(P1_DATAO_REG_18__SCAN_IN), .S(n9376), .Z(
        P1_U3572) );
  MUX2_X1 U10700 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9362), .S(P1_U3973), .Z(
        P1_U3571) );
  MUX2_X1 U10701 ( .A(n9363), .B(P1_DATAO_REG_16__SCAN_IN), .S(n9376), .Z(
        P1_U3570) );
  MUX2_X1 U10702 ( .A(n9364), .B(P1_DATAO_REG_15__SCAN_IN), .S(n9376), .Z(
        P1_U3569) );
  MUX2_X1 U10703 ( .A(n9365), .B(P1_DATAO_REG_14__SCAN_IN), .S(n9376), .Z(
        P1_U3568) );
  MUX2_X1 U10704 ( .A(n9366), .B(P1_DATAO_REG_13__SCAN_IN), .S(n9376), .Z(
        P1_U3567) );
  MUX2_X1 U10705 ( .A(n9367), .B(P1_DATAO_REG_12__SCAN_IN), .S(n9376), .Z(
        P1_U3566) );
  MUX2_X1 U10706 ( .A(n9368), .B(P1_DATAO_REG_11__SCAN_IN), .S(n9376), .Z(
        P1_U3565) );
  MUX2_X1 U10707 ( .A(n6436), .B(P1_DATAO_REG_10__SCAN_IN), .S(n9376), .Z(
        P1_U3564) );
  MUX2_X1 U10708 ( .A(n9369), .B(P1_DATAO_REG_9__SCAN_IN), .S(n9376), .Z(
        P1_U3563) );
  MUX2_X1 U10709 ( .A(n9370), .B(P1_DATAO_REG_8__SCAN_IN), .S(n9376), .Z(
        P1_U3562) );
  MUX2_X1 U10710 ( .A(n9371), .B(P1_DATAO_REG_7__SCAN_IN), .S(n9376), .Z(
        P1_U3561) );
  MUX2_X1 U10711 ( .A(n9372), .B(P1_DATAO_REG_6__SCAN_IN), .S(n9376), .Z(
        P1_U3560) );
  MUX2_X1 U10712 ( .A(n9373), .B(P1_DATAO_REG_5__SCAN_IN), .S(n9376), .Z(
        P1_U3559) );
  MUX2_X1 U10713 ( .A(n9374), .B(P1_DATAO_REG_4__SCAN_IN), .S(n9376), .Z(
        P1_U3558) );
  MUX2_X1 U10714 ( .A(n6931), .B(P1_DATAO_REG_3__SCAN_IN), .S(n9376), .Z(
        P1_U3557) );
  MUX2_X1 U10715 ( .A(n9375), .B(P1_DATAO_REG_2__SCAN_IN), .S(n9376), .Z(
        P1_U3556) );
  MUX2_X1 U10716 ( .A(n6849), .B(P1_DATAO_REG_1__SCAN_IN), .S(n9376), .Z(
        P1_U3555) );
  MUX2_X1 U10717 ( .A(n9377), .B(P1_DATAO_REG_0__SCAN_IN), .S(n9376), .Z(
        P1_U3554) );
  INV_X1 U10718 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n9378) );
  OAI22_X1 U10719 ( .A1(n9995), .A2(n7641), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9378), .ZN(n9379) );
  AOI21_X1 U10720 ( .B1(n9380), .B2(n4395), .A(n9379), .ZN(n9388) );
  OAI211_X1 U10721 ( .C1(n9383), .C2(n9382), .A(n9966), .B(n9381), .ZN(n9387)
         );
  OAI211_X1 U10722 ( .C1(n9385), .C2(n9394), .A(n9598), .B(n9384), .ZN(n9386)
         );
  NAND3_X1 U10723 ( .A1(n9388), .A2(n9387), .A3(n9386), .ZN(P1_U3244) );
  NAND2_X1 U10724 ( .A1(n9390), .A2(n4281), .ZN(n9396) );
  AOI22_X1 U10725 ( .A1(n9394), .A2(n9393), .B1(n9392), .B2(n9391), .ZN(n9395)
         );
  OAI211_X1 U10726 ( .C1(n9397), .C2(n9396), .A(P1_U3973), .B(n9395), .ZN(
        n9437) );
  INV_X1 U10727 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n9399) );
  INV_X1 U10728 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n9398) );
  OAI22_X1 U10729 ( .A1(n9995), .A2(n9399), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9398), .ZN(n9400) );
  AOI21_X1 U10730 ( .B1(n9401), .B2(n4395), .A(n9400), .ZN(n9410) );
  OAI211_X1 U10731 ( .C1(n9404), .C2(n9403), .A(n9598), .B(n9402), .ZN(n9409)
         );
  OAI211_X1 U10732 ( .C1(n9407), .C2(n9406), .A(n9966), .B(n9405), .ZN(n9408)
         );
  NAND4_X1 U10733 ( .A1(n9437), .A2(n9410), .A3(n9409), .A4(n9408), .ZN(
        P1_U3245) );
  NAND2_X1 U10734 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_U3086), .ZN(n9411) );
  OAI21_X1 U10735 ( .B1(n9995), .B2(n9412), .A(n9411), .ZN(n9413) );
  AOI21_X1 U10736 ( .B1(n9414), .B2(n4395), .A(n9413), .ZN(n9423) );
  OAI211_X1 U10737 ( .C1(n9417), .C2(n9416), .A(n9598), .B(n9415), .ZN(n9422)
         );
  OAI211_X1 U10738 ( .C1(n9420), .C2(n9419), .A(n9966), .B(n9418), .ZN(n9421)
         );
  NAND3_X1 U10739 ( .A1(n9423), .A2(n9422), .A3(n9421), .ZN(P1_U3246) );
  INV_X1 U10740 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n9425) );
  OAI21_X1 U10741 ( .B1(n9995), .B2(n9425), .A(n9424), .ZN(n9426) );
  AOI21_X1 U10742 ( .B1(n9427), .B2(n4395), .A(n9426), .ZN(n9436) );
  OAI211_X1 U10743 ( .C1(n9430), .C2(n9429), .A(n9966), .B(n9428), .ZN(n9435)
         );
  OAI211_X1 U10744 ( .C1(n9433), .C2(n9432), .A(n9598), .B(n9431), .ZN(n9434)
         );
  NAND4_X1 U10745 ( .A1(n9437), .A2(n9436), .A3(n9435), .A4(n9434), .ZN(
        P1_U3247) );
  INV_X1 U10746 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n9439) );
  NAND2_X1 U10747 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n9438) );
  OAI21_X1 U10748 ( .B1(n9995), .B2(n9439), .A(n9438), .ZN(n9440) );
  AOI21_X1 U10749 ( .B1(n9441), .B2(n4395), .A(n9440), .ZN(n9450) );
  OAI211_X1 U10750 ( .C1(n9444), .C2(n9443), .A(n9598), .B(n9442), .ZN(n9449)
         );
  OAI211_X1 U10751 ( .C1(n9447), .C2(n9446), .A(n9966), .B(n9445), .ZN(n9448)
         );
  NAND3_X1 U10752 ( .A1(n9450), .A2(n9449), .A3(n9448), .ZN(P1_U3248) );
  INV_X1 U10753 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n9452) );
  NAND2_X1 U10754 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_U3086), .ZN(n9451) );
  OAI21_X1 U10755 ( .B1(n9995), .B2(n9452), .A(n9451), .ZN(n9453) );
  AOI21_X1 U10756 ( .B1(n9454), .B2(n4395), .A(n9453), .ZN(n9463) );
  OAI211_X1 U10757 ( .C1(n9457), .C2(n9456), .A(n9966), .B(n9455), .ZN(n9462)
         );
  OAI211_X1 U10758 ( .C1(n9460), .C2(n9459), .A(n9598), .B(n9458), .ZN(n9461)
         );
  NAND3_X1 U10759 ( .A1(n9463), .A2(n9462), .A3(n9461), .ZN(P1_U3249) );
  NAND2_X1 U10760 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3086), .ZN(n9464) );
  OAI21_X1 U10761 ( .B1(n9995), .B2(n9465), .A(n9464), .ZN(n9466) );
  AOI21_X1 U10762 ( .B1(n9467), .B2(n4395), .A(n9466), .ZN(n9476) );
  OAI211_X1 U10763 ( .C1(n9470), .C2(n9469), .A(n9966), .B(n9468), .ZN(n9475)
         );
  OAI211_X1 U10764 ( .C1(n9473), .C2(n9472), .A(n9598), .B(n9471), .ZN(n9474)
         );
  NAND3_X1 U10765 ( .A1(n9476), .A2(n9475), .A3(n9474), .ZN(P1_U3250) );
  OAI211_X1 U10766 ( .C1(n9479), .C2(n9478), .A(n9477), .B(n9598), .ZN(n9489)
         );
  OAI21_X1 U10767 ( .B1(n9995), .B2(n9481), .A(n9480), .ZN(n9482) );
  AOI21_X1 U10768 ( .B1(n9483), .B2(n4395), .A(n9482), .ZN(n9488) );
  OAI211_X1 U10769 ( .C1(n9486), .C2(n9485), .A(n9966), .B(n9484), .ZN(n9487)
         );
  NAND3_X1 U10770 ( .A1(n9489), .A2(n9488), .A3(n9487), .ZN(P1_U3251) );
  OAI211_X1 U10771 ( .C1(n9492), .C2(n9491), .A(n9490), .B(n9598), .ZN(n9503)
         );
  INV_X1 U10772 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n9494) );
  NAND2_X1 U10773 ( .A1(P1_REG3_REG_10__SCAN_IN), .A2(P1_U3086), .ZN(n9493) );
  OAI21_X1 U10774 ( .B1(n9995), .B2(n9494), .A(n9493), .ZN(n9495) );
  AOI21_X1 U10775 ( .B1(n9496), .B2(n4395), .A(n9495), .ZN(n9502) );
  AOI21_X1 U10776 ( .B1(n9498), .B2(n9497), .A(n9981), .ZN(n9500) );
  NAND2_X1 U10777 ( .A1(n9500), .A2(n9499), .ZN(n9501) );
  NAND3_X1 U10778 ( .A1(n9503), .A2(n9502), .A3(n9501), .ZN(P1_U3253) );
  OAI211_X1 U10779 ( .C1(n9506), .C2(n9505), .A(n9504), .B(n9598), .ZN(n9516)
         );
  INV_X1 U10780 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n9508) );
  OAI21_X1 U10781 ( .B1(n9995), .B2(n9508), .A(n9507), .ZN(n9509) );
  AOI21_X1 U10782 ( .B1(n9510), .B2(n4395), .A(n9509), .ZN(n9515) );
  OAI211_X1 U10783 ( .C1(n9513), .C2(n9512), .A(n9511), .B(n9966), .ZN(n9514)
         );
  NAND3_X1 U10784 ( .A1(n9516), .A2(n9515), .A3(n9514), .ZN(P1_U3254) );
  XOR2_X1 U10785 ( .A(P1_REG2_REG_13__SCAN_IN), .B(n9541), .Z(n9519) );
  OAI211_X1 U10786 ( .C1(n9520), .C2(n9519), .A(n9533), .B(n9598), .ZN(n9532)
         );
  OAI21_X1 U10787 ( .B1(n9995), .B2(n9522), .A(n9521), .ZN(n9523) );
  AOI21_X1 U10788 ( .B1(n9541), .B2(n4395), .A(n9523), .ZN(n9531) );
  OR2_X1 U10789 ( .A1(n9524), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n9525) );
  AND2_X1 U10790 ( .A1(n9526), .A2(n9525), .ZN(n9529) );
  XNOR2_X1 U10791 ( .A(n9541), .B(n9527), .ZN(n9528) );
  NAND2_X1 U10792 ( .A1(n9529), .A2(n9528), .ZN(n9543) );
  OAI211_X1 U10793 ( .C1(n9529), .C2(n9528), .A(n9543), .B(n9966), .ZN(n9530)
         );
  NAND3_X1 U10794 ( .A1(n9532), .A2(n9531), .A3(n9530), .ZN(P1_U3256) );
  XOR2_X1 U10795 ( .A(P1_REG2_REG_14__SCAN_IN), .B(n9550), .Z(n9536) );
  OAI211_X1 U10796 ( .C1(n9537), .C2(n9536), .A(n9561), .B(n9598), .ZN(n9549)
         );
  NAND2_X1 U10797 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n9538) );
  OAI21_X1 U10798 ( .B1(n9995), .B2(n9539), .A(n9538), .ZN(n9540) );
  AOI21_X1 U10799 ( .B1(n9550), .B2(n4395), .A(n9540), .ZN(n9548) );
  NAND2_X1 U10800 ( .A1(n9541), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n9542) );
  NAND2_X1 U10801 ( .A1(n9543), .A2(n9542), .ZN(n9546) );
  INV_X1 U10802 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n9544) );
  XNOR2_X1 U10803 ( .A(n9550), .B(n9544), .ZN(n9545) );
  NAND2_X1 U10804 ( .A1(n9546), .A2(n9545), .ZN(n9552) );
  OAI211_X1 U10805 ( .C1(n9546), .C2(n9545), .A(n9552), .B(n9966), .ZN(n9547)
         );
  NAND3_X1 U10806 ( .A1(n9549), .A2(n9548), .A3(n9547), .ZN(P1_U3257) );
  XNOR2_X1 U10807 ( .A(n9578), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n9558) );
  NAND2_X1 U10808 ( .A1(n9550), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n9551) );
  NAND2_X1 U10809 ( .A1(n9552), .A2(n9551), .ZN(n9554) );
  XNOR2_X1 U10810 ( .A(n9554), .B(n9553), .ZN(n9968) );
  NAND2_X1 U10811 ( .A1(n9968), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n9967) );
  NAND2_X1 U10812 ( .A1(n9554), .A2(n9975), .ZN(n9555) );
  NAND2_X1 U10813 ( .A1(n9967), .A2(n9555), .ZN(n9557) );
  INV_X1 U10814 ( .A(n9580), .ZN(n9556) );
  AOI21_X1 U10815 ( .B1(n9558), .B2(n9557), .A(n9556), .ZN(n9570) );
  OAI21_X1 U10816 ( .B1(n9995), .B2(n9560), .A(n9559), .ZN(n9568) );
  INV_X1 U10817 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n9562) );
  INV_X1 U10818 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n9971) );
  XNOR2_X1 U10819 ( .A(n9564), .B(n9975), .ZN(n9972) );
  AOI21_X1 U10820 ( .B1(n9564), .B2(n9975), .A(n9970), .ZN(n9566) );
  XNOR2_X1 U10821 ( .A(n9578), .B(P1_REG2_REG_16__SCAN_IN), .ZN(n9565) );
  NOR2_X1 U10822 ( .A1(n9566), .A2(n9565), .ZN(n9571) );
  AOI211_X1 U10823 ( .C1(n9566), .C2(n9565), .A(n9986), .B(n9571), .ZN(n9567)
         );
  AOI211_X1 U10824 ( .C1(n4395), .C2(n9578), .A(n9568), .B(n9567), .ZN(n9569)
         );
  OAI21_X1 U10825 ( .B1(n9570), .B2(n9981), .A(n9569), .ZN(P1_U3259) );
  XOR2_X1 U10826 ( .A(P1_REG2_REG_17__SCAN_IN), .B(n9592), .Z(n9573) );
  OAI21_X1 U10827 ( .B1(n9573), .B2(n9572), .A(n9588), .ZN(n9574) );
  NAND2_X1 U10828 ( .A1(n9574), .A2(n9598), .ZN(n9587) );
  AOI21_X1 U10829 ( .B1(n9576), .B2(P1_ADDR_REG_17__SCAN_IN), .A(n9575), .ZN(
        n9586) );
  XNOR2_X1 U10830 ( .A(n9592), .B(n9577), .ZN(n9582) );
  OR2_X1 U10831 ( .A1(n9578), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n9579) );
  NAND2_X1 U10832 ( .A1(n9580), .A2(n9579), .ZN(n9581) );
  NAND2_X1 U10833 ( .A1(n9581), .A2(n9582), .ZN(n9594) );
  OAI21_X1 U10834 ( .B1(n9582), .B2(n9581), .A(n9594), .ZN(n9583) );
  NAND2_X1 U10835 ( .A1(n9583), .A2(n9966), .ZN(n9585) );
  NAND2_X1 U10836 ( .A1(n4395), .A2(n9592), .ZN(n9584) );
  NAND4_X1 U10837 ( .A1(n9587), .A2(n9586), .A3(n9585), .A4(n9584), .ZN(
        P1_U3260) );
  NAND2_X1 U10838 ( .A1(n9991), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9589) );
  OAI21_X1 U10839 ( .B1(n9991), .B2(P1_REG2_REG_18__SCAN_IN), .A(n9589), .ZN(
        n9988) );
  NAND2_X1 U10840 ( .A1(n9984), .A2(n9589), .ZN(n9591) );
  XNOR2_X1 U10841 ( .A(n9591), .B(n9590), .ZN(n9599) );
  OR2_X1 U10842 ( .A1(n9592), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n9593) );
  NAND2_X1 U10843 ( .A1(n9594), .A2(n9593), .ZN(n9982) );
  NAND2_X1 U10844 ( .A1(n9991), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n9595) );
  OAI21_X1 U10845 ( .B1(n9991), .B2(P1_REG1_REG_18__SCAN_IN), .A(n9595), .ZN(
        n9983) );
  NAND2_X1 U10846 ( .A1(n9979), .A2(n9595), .ZN(n9596) );
  XNOR2_X1 U10847 ( .A(n9596), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n9600) );
  INV_X1 U10848 ( .A(n9600), .ZN(n9597) );
  AOI22_X1 U10849 ( .A1(n9599), .A2(n9598), .B1(n9966), .B2(n9597), .ZN(n9601)
         );
  NAND2_X1 U10850 ( .A1(P1_REG3_REG_19__SCAN_IN), .A2(P1_U3086), .ZN(n9602) );
  XNOR2_X1 U10851 ( .A(n9604), .B(n4735), .ZN(n9605) );
  NAND2_X1 U10852 ( .A1(n9605), .A2(n10035), .ZN(n9829) );
  NOR2_X1 U10853 ( .A1(n9996), .A2(n9606), .ZN(n9608) );
  AOI211_X1 U10854 ( .C1(n4735), .C2(n10042), .A(n9608), .B(n9607), .ZN(n9609)
         );
  OAI21_X1 U10855 ( .B1(n9829), .B2(n9610), .A(n9609), .ZN(P1_U3263) );
  AND2_X1 U10856 ( .A1(n9636), .A2(n9612), .ZN(n9835) );
  INV_X1 U10857 ( .A(n9835), .ZN(n9837) );
  NAND2_X1 U10858 ( .A1(n9845), .A2(n9837), .ZN(n9613) );
  XNOR2_X1 U10859 ( .A(n9613), .B(n9838), .ZN(n9634) );
  NAND2_X1 U10860 ( .A1(n10041), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n9615) );
  OAI22_X1 U10861 ( .A1(n9616), .A2(n9615), .B1(n9614), .B2(n9996), .ZN(n9617)
         );
  AOI21_X1 U10862 ( .B1(n9839), .B2(n10042), .A(n9617), .ZN(n9633) );
  AOI21_X1 U10863 ( .B1(n9839), .B2(n9618), .A(n8236), .ZN(n9620) );
  NAND2_X1 U10864 ( .A1(n9622), .A2(n9621), .ZN(n9623) );
  XNOR2_X1 U10865 ( .A(n9623), .B(n9836), .ZN(n9629) );
  OAI22_X1 U10866 ( .A1(n9627), .A2(n9626), .B1(n9625), .B2(n9624), .ZN(n9628)
         );
  OAI21_X1 U10867 ( .B1(n9630), .B2(n9843), .A(n9846), .ZN(n9631) );
  NAND2_X1 U10868 ( .A1(n9631), .A2(n9996), .ZN(n9632) );
  OAI211_X1 U10869 ( .C1(n9634), .C2(n9828), .A(n9633), .B(n9632), .ZN(
        P1_U3356) );
  INV_X1 U10870 ( .A(n9635), .ZN(n9646) );
  INV_X1 U10871 ( .A(n9636), .ZN(n9638) );
  INV_X1 U10872 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n9637) );
  OAI22_X1 U10873 ( .A1(n9638), .A2(n9816), .B1(n9637), .B2(n9996), .ZN(n9643)
         );
  NAND2_X1 U10874 ( .A1(n9639), .A2(n10041), .ZN(n9640) );
  AOI21_X1 U10875 ( .B1(n9641), .B2(n9640), .A(n9768), .ZN(n9642) );
  OAI21_X1 U10876 ( .B1(n9646), .B2(n9828), .A(n9645), .ZN(P1_U3265) );
  XNOR2_X1 U10877 ( .A(n9647), .B(n9648), .ZN(n9856) );
  INV_X1 U10878 ( .A(n9649), .ZN(n9651) );
  INV_X1 U10879 ( .A(n6484), .ZN(n9650) );
  AOI211_X1 U10880 ( .C1(n9850), .C2(n9651), .A(n8236), .B(n9650), .ZN(n9849)
         );
  NOR2_X1 U10881 ( .A1(n9652), .A2(n9816), .ZN(n9656) );
  OAI22_X1 U10882 ( .A1(n9654), .A2(n9806), .B1(n9653), .B2(n9996), .ZN(n9655)
         );
  AOI211_X1 U10883 ( .C1(n9849), .C2(n9826), .A(n9656), .B(n9655), .ZN(n9663)
         );
  XNOR2_X1 U10884 ( .A(n9658), .B(n9657), .ZN(n9659) );
  NAND2_X1 U10885 ( .A1(n9659), .A2(n10030), .ZN(n9661) );
  NAND2_X1 U10886 ( .A1(n9661), .A2(n9660), .ZN(n9854) );
  NAND2_X1 U10887 ( .A1(n9854), .A2(n9996), .ZN(n9662) );
  OAI211_X1 U10888 ( .C1(n9856), .C2(n9828), .A(n9663), .B(n9662), .ZN(
        P1_U3266) );
  XNOR2_X1 U10889 ( .A(n9664), .B(n9665), .ZN(n9861) );
  INV_X1 U10890 ( .A(n9667), .ZN(n9668) );
  INV_X1 U10891 ( .A(n4315), .ZN(n9669) );
  AOI211_X1 U10892 ( .C1(n9859), .C2(n9669), .A(n8236), .B(n9649), .ZN(n9858)
         );
  NAND2_X1 U10893 ( .A1(n9858), .A2(n9826), .ZN(n9672) );
  AOI22_X1 U10894 ( .A1(n9670), .A2(n10041), .B1(P1_REG2_REG_26__SCAN_IN), 
        .B2(n9768), .ZN(n9671) );
  OAI211_X1 U10895 ( .C1(n9673), .C2(n9816), .A(n9672), .B(n9671), .ZN(n9674)
         );
  AOI21_X1 U10896 ( .B1(n9857), .B2(n9996), .A(n9674), .ZN(n9675) );
  OAI21_X1 U10897 ( .B1(n9861), .B2(n9828), .A(n9675), .ZN(P1_U3267) );
  XNOR2_X1 U10898 ( .A(n9676), .B(n9681), .ZN(n9866) );
  AOI211_X1 U10899 ( .C1(n9863), .C2(n9696), .A(n8236), .B(n4315), .ZN(n9862)
         );
  INV_X1 U10900 ( .A(n9677), .ZN(n9678) );
  AOI22_X1 U10901 ( .A1(n9678), .A2(n10041), .B1(P1_REG2_REG_25__SCAN_IN), 
        .B2(n9768), .ZN(n9679) );
  OAI21_X1 U10902 ( .B1(n9680), .B2(n9816), .A(n9679), .ZN(n9685) );
  XNOR2_X1 U10903 ( .A(n4365), .B(n9681), .ZN(n9683) );
  AOI21_X1 U10904 ( .B1(n9683), .B2(n10030), .A(n9682), .ZN(n9865) );
  NOR2_X1 U10905 ( .A1(n9865), .A2(n9768), .ZN(n9684) );
  AOI211_X1 U10906 ( .C1(n9862), .C2(n9826), .A(n9685), .B(n9684), .ZN(n9686)
         );
  OAI21_X1 U10907 ( .B1(n9866), .B2(n9828), .A(n9686), .ZN(P1_U3268) );
  XNOR2_X1 U10908 ( .A(n9687), .B(n9688), .ZN(n9871) );
  NAND2_X1 U10909 ( .A1(n9689), .A2(n9690), .ZN(n9692) );
  XNOR2_X1 U10910 ( .A(n9692), .B(n9691), .ZN(n9694) );
  OAI21_X1 U10911 ( .B1(n9694), .B2(n10000), .A(n9693), .ZN(n9867) );
  INV_X1 U10912 ( .A(n9696), .ZN(n9697) );
  AOI211_X1 U10913 ( .C1(n9869), .C2(n9695), .A(n8236), .B(n9697), .ZN(n9868)
         );
  NAND2_X1 U10914 ( .A1(n9868), .A2(n9826), .ZN(n9701) );
  INV_X1 U10915 ( .A(n9698), .ZN(n9699) );
  AOI22_X1 U10916 ( .A1(n9699), .A2(n10041), .B1(P1_REG2_REG_24__SCAN_IN), 
        .B2(n9768), .ZN(n9700) );
  OAI211_X1 U10917 ( .C1(n9702), .C2(n9816), .A(n9701), .B(n9700), .ZN(n9703)
         );
  AOI21_X1 U10918 ( .B1(n9996), .B2(n9867), .A(n9703), .ZN(n9704) );
  OAI21_X1 U10919 ( .B1(n9871), .B2(n9828), .A(n9704), .ZN(P1_U3269) );
  XOR2_X1 U10920 ( .A(n9705), .B(n9713), .Z(n9876) );
  INV_X1 U10921 ( .A(n9706), .ZN(n9708) );
  INV_X1 U10922 ( .A(n9695), .ZN(n9707) );
  AOI211_X1 U10923 ( .C1(n9873), .C2(n9708), .A(n8236), .B(n9707), .ZN(n9872)
         );
  AOI22_X1 U10924 ( .A1(n9709), .A2(n10041), .B1(P1_REG2_REG_23__SCAN_IN), 
        .B2(n9768), .ZN(n9710) );
  OAI21_X1 U10925 ( .B1(n9711), .B2(n9816), .A(n9710), .ZN(n9718) );
  AND2_X1 U10926 ( .A1(n9726), .A2(n9712), .ZN(n9714) );
  OAI21_X1 U10927 ( .B1(n9714), .B2(n9713), .A(n9689), .ZN(n9716) );
  AOI21_X1 U10928 ( .B1(n9716), .B2(n10030), .A(n9715), .ZN(n9875) );
  NOR2_X1 U10929 ( .A1(n9875), .A2(n9768), .ZN(n9717) );
  AOI211_X1 U10930 ( .C1(n9872), .C2(n10046), .A(n9718), .B(n9717), .ZN(n9719)
         );
  OAI21_X1 U10931 ( .B1(n9876), .B2(n9828), .A(n9719), .ZN(P1_U3270) );
  XNOR2_X1 U10932 ( .A(n9720), .B(n9727), .ZN(n9881) );
  INV_X1 U10933 ( .A(n9744), .ZN(n9721) );
  AOI211_X1 U10934 ( .C1(n9878), .C2(n9721), .A(n8236), .B(n9706), .ZN(n9877)
         );
  INV_X1 U10935 ( .A(n9722), .ZN(n9723) );
  AOI22_X1 U10936 ( .A1(n9723), .A2(n10041), .B1(P1_REG2_REG_22__SCAN_IN), 
        .B2(n9768), .ZN(n9724) );
  OAI21_X1 U10937 ( .B1(n9725), .B2(n9816), .A(n9724), .ZN(n9735) );
  INV_X1 U10938 ( .A(n9726), .ZN(n9731) );
  AOI21_X1 U10939 ( .B1(n9729), .B2(n9728), .A(n9727), .ZN(n9730) );
  NOR3_X1 U10940 ( .A1(n9731), .A2(n9730), .A3(n10000), .ZN(n9733) );
  NOR2_X1 U10941 ( .A1(n9733), .A2(n9732), .ZN(n9880) );
  NOR2_X1 U10942 ( .A1(n9880), .A2(n9768), .ZN(n9734) );
  AOI211_X1 U10943 ( .C1(n9877), .C2(n9826), .A(n9735), .B(n9734), .ZN(n9736)
         );
  OAI21_X1 U10944 ( .B1(n9881), .B2(n9828), .A(n9736), .ZN(P1_U3271) );
  INV_X1 U10945 ( .A(n9737), .ZN(n9739) );
  OAI21_X1 U10946 ( .B1(n6470), .B2(n9739), .A(n9738), .ZN(n9740) );
  XOR2_X1 U10947 ( .A(n9748), .B(n9740), .Z(n9743) );
  INV_X1 U10948 ( .A(n9741), .ZN(n9742) );
  AOI21_X1 U10949 ( .B1(n9743), .B2(n10030), .A(n9742), .ZN(n9885) );
  AOI21_X1 U10950 ( .B1(n9882), .B2(n9758), .A(n9744), .ZN(n9883) );
  AOI22_X1 U10951 ( .A1(n9745), .A2(n10041), .B1(P1_REG2_REG_21__SCAN_IN), 
        .B2(n9768), .ZN(n9746) );
  OAI21_X1 U10952 ( .B1(n9747), .B2(n9816), .A(n9746), .ZN(n9751) );
  XNOR2_X1 U10953 ( .A(n9749), .B(n9748), .ZN(n9886) );
  NOR2_X1 U10954 ( .A1(n9886), .A2(n9828), .ZN(n9750) );
  AOI211_X1 U10955 ( .C1(n9883), .C2(n9752), .A(n9751), .B(n9750), .ZN(n9753)
         );
  OAI21_X1 U10956 ( .B1(n9768), .B2(n9885), .A(n9753), .ZN(P1_U3272) );
  XNOR2_X1 U10957 ( .A(n6470), .B(n4479), .ZN(n9756) );
  INV_X1 U10958 ( .A(n9754), .ZN(n9755) );
  AOI21_X1 U10959 ( .B1(n9756), .B2(n10030), .A(n9755), .ZN(n9890) );
  AOI21_X1 U10960 ( .B1(n9757), .B2(n9888), .A(n8236), .ZN(n9759) );
  AND2_X1 U10961 ( .A1(n9759), .A2(n9758), .ZN(n9887) );
  NAND2_X1 U10962 ( .A1(n9888), .A2(n10042), .ZN(n9761) );
  NAND2_X1 U10963 ( .A1(n9768), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n9760) );
  OAI211_X1 U10964 ( .C1(n9806), .C2(n9762), .A(n9761), .B(n9760), .ZN(n9766)
         );
  XNOR2_X1 U10965 ( .A(n9764), .B(n9763), .ZN(n9891) );
  NOR2_X1 U10966 ( .A1(n9891), .A2(n9828), .ZN(n9765) );
  AOI211_X1 U10967 ( .C1(n9887), .C2(n10046), .A(n9766), .B(n9765), .ZN(n9767)
         );
  OAI21_X1 U10968 ( .B1(n9768), .B2(n9890), .A(n9767), .ZN(P1_U3273) );
  XOR2_X1 U10969 ( .A(n9769), .B(n9778), .Z(n9896) );
  INV_X1 U10970 ( .A(n9770), .ZN(n9772) );
  INV_X1 U10971 ( .A(n9757), .ZN(n9771) );
  AOI211_X1 U10972 ( .C1(n9893), .C2(n9772), .A(n8236), .B(n9771), .ZN(n9892)
         );
  AOI22_X1 U10973 ( .A1(n9773), .A2(n10041), .B1(P1_REG2_REG_19__SCAN_IN), 
        .B2(n9768), .ZN(n9774) );
  OAI21_X1 U10974 ( .B1(n9775), .B2(n9816), .A(n9774), .ZN(n9782) );
  OAI21_X1 U10975 ( .B1(n9778), .B2(n9777), .A(n9776), .ZN(n9780) );
  AOI21_X1 U10976 ( .B1(n9780), .B2(n10030), .A(n9779), .ZN(n9895) );
  NOR2_X1 U10977 ( .A1(n9895), .A2(n9768), .ZN(n9781) );
  AOI211_X1 U10978 ( .C1(n9892), .C2(n9826), .A(n9782), .B(n9781), .ZN(n9783)
         );
  OAI21_X1 U10979 ( .B1(n9896), .B2(n9828), .A(n9783), .ZN(P1_U3274) );
  XNOR2_X1 U10980 ( .A(n4328), .B(n9784), .ZN(n9901) );
  AOI22_X1 U10981 ( .A1(n9898), .A2(n10042), .B1(P1_REG2_REG_18__SCAN_IN), 
        .B2(n9768), .ZN(n9793) );
  OAI21_X1 U10982 ( .B1(n4373), .B2(n5788), .A(n9785), .ZN(n9787) );
  AOI21_X1 U10983 ( .B1(n9787), .B2(n10030), .A(n9786), .ZN(n9900) );
  AOI211_X1 U10984 ( .C1(n9898), .C2(n9797), .A(n8236), .B(n9770), .ZN(n9897)
         );
  NAND2_X1 U10985 ( .A1(n9897), .A2(n9788), .ZN(n9789) );
  OAI211_X1 U10986 ( .C1(n9806), .C2(n9790), .A(n9900), .B(n9789), .ZN(n9791)
         );
  NAND2_X1 U10987 ( .A1(n9791), .A2(n9996), .ZN(n9792) );
  OAI211_X1 U10988 ( .C1(n9901), .C2(n9828), .A(n9793), .B(n9792), .ZN(
        P1_U3275) );
  XNOR2_X1 U10989 ( .A(n9794), .B(n9802), .ZN(n9906) );
  AOI21_X1 U10990 ( .B1(n4855), .B2(n9903), .A(n8236), .ZN(n9796) );
  AND2_X1 U10991 ( .A1(n9797), .A2(n9796), .ZN(n9902) );
  INV_X1 U10992 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n9798) );
  OAI22_X1 U10993 ( .A1(n9799), .A2(n9816), .B1(n9996), .B2(n9798), .ZN(n9800)
         );
  AOI21_X1 U10994 ( .B1(n9902), .B2(n9826), .A(n9800), .ZN(n9810) );
  NAND2_X1 U10995 ( .A1(n9818), .A2(n9801), .ZN(n9803) );
  XNOR2_X1 U10996 ( .A(n9803), .B(n9802), .ZN(n9805) );
  AOI21_X1 U10997 ( .B1(n9805), .B2(n10030), .A(n9804), .ZN(n9905) );
  OAI21_X1 U10998 ( .B1(n9807), .B2(n9806), .A(n9905), .ZN(n9808) );
  NAND2_X1 U10999 ( .A1(n9808), .A2(n9996), .ZN(n9809) );
  OAI211_X1 U11000 ( .C1(n9906), .C2(n9828), .A(n9810), .B(n9809), .ZN(
        P1_U3276) );
  XNOR2_X1 U11001 ( .A(n9811), .B(n4697), .ZN(n9911) );
  AOI211_X1 U11002 ( .C1(n9908), .C2(n9812), .A(n8236), .B(n9795), .ZN(n9907)
         );
  INV_X1 U11003 ( .A(n9908), .ZN(n9817) );
  INV_X1 U11004 ( .A(n9813), .ZN(n9814) );
  AOI22_X1 U11005 ( .A1(n9768), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n9814), .B2(
        n10041), .ZN(n9815) );
  OAI21_X1 U11006 ( .B1(n9817), .B2(n9816), .A(n9815), .ZN(n9825) );
  OAI21_X1 U11007 ( .B1(n9820), .B2(n9819), .A(n9818), .ZN(n9823) );
  INV_X1 U11008 ( .A(n9821), .ZN(n9822) );
  AOI21_X1 U11009 ( .B1(n9823), .B2(n10030), .A(n9822), .ZN(n9910) );
  NOR2_X1 U11010 ( .A1(n9910), .A2(n9768), .ZN(n9824) );
  AOI211_X1 U11011 ( .C1(n9907), .C2(n9826), .A(n9825), .B(n9824), .ZN(n9827)
         );
  OAI21_X1 U11012 ( .B1(n9911), .B2(n9828), .A(n9827), .ZN(P1_U3277) );
  OAI211_X1 U11013 ( .C1(n9830), .C2(n10103), .A(n9829), .B(n9831), .ZN(n9932)
         );
  MUX2_X1 U11014 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n9932), .S(n10124), .Z(
        P1_U3553) );
  OAI211_X1 U11015 ( .C1(n9833), .C2(n10103), .A(n9832), .B(n9831), .ZN(n9933)
         );
  MUX2_X1 U11016 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n9933), .S(n10124), .Z(
        P1_U3552) );
  NAND2_X1 U11017 ( .A1(n9836), .A2(n10107), .ZN(n9834) );
  NOR3_X1 U11018 ( .A1(n9836), .A2(n10088), .A3(n9835), .ZN(n9844) );
  INV_X1 U11019 ( .A(n9839), .ZN(n9840) );
  MUX2_X1 U11020 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n9848), .S(n10124), .Z(
        P1_U3550) );
  NAND2_X1 U11021 ( .A1(n9850), .A2(n10084), .ZN(n9851) );
  MUX2_X1 U11022 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9935), .S(n10124), .Z(
        P1_U3549) );
  OAI21_X1 U11023 ( .B1(n9861), .B2(n10088), .A(n9860), .ZN(n9936) );
  MUX2_X1 U11024 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9936), .S(n10124), .Z(
        P1_U3548) );
  AOI21_X1 U11025 ( .B1(n10084), .B2(n9863), .A(n9862), .ZN(n9864) );
  OAI211_X1 U11026 ( .C1(n9866), .C2(n10088), .A(n9865), .B(n9864), .ZN(n9937)
         );
  MUX2_X1 U11027 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9937), .S(n10124), .Z(
        P1_U3547) );
  AOI211_X1 U11028 ( .C1(n10084), .C2(n9869), .A(n9868), .B(n9867), .ZN(n9870)
         );
  OAI21_X1 U11029 ( .B1(n9871), .B2(n10088), .A(n9870), .ZN(n9938) );
  MUX2_X1 U11030 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9938), .S(n10124), .Z(
        P1_U3546) );
  AOI21_X1 U11031 ( .B1(n10084), .B2(n9873), .A(n9872), .ZN(n9874) );
  OAI211_X1 U11032 ( .C1(n9876), .C2(n10088), .A(n9875), .B(n9874), .ZN(n9939)
         );
  MUX2_X1 U11033 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9939), .S(n10124), .Z(
        P1_U3545) );
  AOI21_X1 U11034 ( .B1(n10084), .B2(n9878), .A(n9877), .ZN(n9879) );
  OAI211_X1 U11035 ( .C1(n9881), .C2(n10088), .A(n9880), .B(n9879), .ZN(n9940)
         );
  MUX2_X1 U11036 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9940), .S(n10124), .Z(
        P1_U3544) );
  AOI22_X1 U11037 ( .A1(n9883), .A2(n10035), .B1(n10084), .B2(n9882), .ZN(
        n9884) );
  OAI211_X1 U11038 ( .C1(n9886), .C2(n10088), .A(n9885), .B(n9884), .ZN(n9941)
         );
  MUX2_X1 U11039 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9941), .S(n10124), .Z(
        P1_U3543) );
  AOI21_X1 U11040 ( .B1(n10084), .B2(n9888), .A(n9887), .ZN(n9889) );
  OAI211_X1 U11041 ( .C1(n9891), .C2(n10088), .A(n9890), .B(n9889), .ZN(n9942)
         );
  MUX2_X1 U11042 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9942), .S(n10124), .Z(
        P1_U3542) );
  AOI21_X1 U11043 ( .B1(n10084), .B2(n9893), .A(n9892), .ZN(n9894) );
  OAI211_X1 U11044 ( .C1(n9896), .C2(n10088), .A(n9895), .B(n9894), .ZN(n9943)
         );
  MUX2_X1 U11045 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9943), .S(n10115), .Z(
        P1_U3541) );
  AOI21_X1 U11046 ( .B1(n10084), .B2(n9898), .A(n9897), .ZN(n9899) );
  OAI211_X1 U11047 ( .C1(n9901), .C2(n10088), .A(n9900), .B(n9899), .ZN(n9944)
         );
  MUX2_X1 U11048 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9944), .S(n10115), .Z(
        P1_U3540) );
  AOI21_X1 U11049 ( .B1(n10084), .B2(n9903), .A(n9902), .ZN(n9904) );
  OAI211_X1 U11050 ( .C1(n9906), .C2(n10088), .A(n9905), .B(n9904), .ZN(n9945)
         );
  MUX2_X1 U11051 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9945), .S(n10115), .Z(
        P1_U3539) );
  AOI21_X1 U11052 ( .B1(n10084), .B2(n9908), .A(n9907), .ZN(n9909) );
  OAI211_X1 U11053 ( .C1(n9911), .C2(n10088), .A(n9910), .B(n9909), .ZN(n9946)
         );
  MUX2_X1 U11054 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9946), .S(n10115), .Z(
        P1_U3538) );
  AOI211_X1 U11055 ( .C1(n10084), .C2(n9914), .A(n9913), .B(n9912), .ZN(n9915)
         );
  OAI21_X1 U11056 ( .B1(n9916), .B2(n10088), .A(n9915), .ZN(n9947) );
  MUX2_X1 U11057 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n9947), .S(n10115), .Z(
        P1_U3537) );
  AOI211_X1 U11058 ( .C1(n10084), .C2(n5461), .A(n9918), .B(n9917), .ZN(n9919)
         );
  OAI21_X1 U11059 ( .B1(n9920), .B2(n10088), .A(n9919), .ZN(n9948) );
  MUX2_X1 U11060 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n9948), .S(n10115), .Z(
        P1_U3536) );
  AOI21_X1 U11061 ( .B1(n10084), .B2(n9922), .A(n9921), .ZN(n9923) );
  OAI211_X1 U11062 ( .C1(n9925), .C2(n10088), .A(n9924), .B(n9923), .ZN(n9949)
         );
  MUX2_X1 U11063 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n9949), .S(n10115), .Z(
        P1_U3535) );
  AOI211_X1 U11064 ( .C1(n10084), .C2(n9928), .A(n9927), .B(n9926), .ZN(n9929)
         );
  OAI21_X1 U11065 ( .B1(n9930), .B2(n10088), .A(n9929), .ZN(n9950) );
  MUX2_X1 U11066 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n9950), .S(n10124), .Z(
        P1_U3534) );
  MUX2_X1 U11067 ( .A(n9931), .B(P1_REG1_REG_0__SCAN_IN), .S(n10122), .Z(
        P1_U3522) );
  MUX2_X1 U11068 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n9932), .S(n4272), .Z(
        P1_U3521) );
  MUX2_X1 U11069 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n9933), .S(n4272), .Z(
        P1_U3520) );
  MUX2_X1 U11070 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9935), .S(n4272), .Z(
        P1_U3517) );
  MUX2_X1 U11071 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9936), .S(n4272), .Z(
        P1_U3516) );
  MUX2_X1 U11072 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9937), .S(n4272), .Z(
        P1_U3515) );
  MUX2_X1 U11073 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9938), .S(n4272), .Z(
        P1_U3514) );
  MUX2_X1 U11074 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9939), .S(n4272), .Z(
        P1_U3513) );
  MUX2_X1 U11075 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9940), .S(n4272), .Z(
        P1_U3512) );
  MUX2_X1 U11076 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9941), .S(n4272), .Z(
        P1_U3511) );
  MUX2_X1 U11077 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9942), .S(n4272), .Z(
        P1_U3510) );
  MUX2_X1 U11078 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9943), .S(n4272), .Z(
        P1_U3509) );
  MUX2_X1 U11079 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9944), .S(n4272), .Z(
        P1_U3507) );
  MUX2_X1 U11080 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9945), .S(n4272), .Z(
        P1_U3504) );
  MUX2_X1 U11081 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n9946), .S(n4272), .Z(
        P1_U3501) );
  MUX2_X1 U11082 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n9947), .S(n4272), .Z(
        P1_U3498) );
  MUX2_X1 U11083 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n9948), .S(n4272), .Z(
        P1_U3495) );
  MUX2_X1 U11084 ( .A(P1_REG0_REG_13__SCAN_IN), .B(n9949), .S(n4272), .Z(
        P1_U3492) );
  MUX2_X1 U11085 ( .A(P1_REG0_REG_12__SCAN_IN), .B(n9950), .S(n4272), .Z(
        P1_U3489) );
  MUX2_X1 U11086 ( .A(P1_D_REG_1__SCAN_IN), .B(n9953), .S(n10055), .Z(P1_U3440) );
  MUX2_X1 U11087 ( .A(P1_D_REG_0__SCAN_IN), .B(n9954), .S(n10055), .Z(P1_U3439) );
  NOR4_X1 U11088 ( .A1(n9956), .A2(P1_IR_REG_30__SCAN_IN), .A3(n5168), .A4(
        P1_U3086), .ZN(n9957) );
  AOI21_X1 U11089 ( .B1(n9958), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9957), .ZN(
        n9959) );
  OAI21_X1 U11090 ( .B1(n9960), .B2(n9963), .A(n9959), .ZN(P1_U3324) );
  INV_X1 U11091 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n9961) );
  OAI222_X1 U11092 ( .A1(n9964), .A2(P1_U3086), .B1(n9963), .B2(n9962), .C1(
        n9961), .C2(n8253), .ZN(P1_U3326) );
  MUX2_X1 U11093 ( .A(n9965), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  XNOR2_X1 U11094 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U11095 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  OAI211_X1 U11096 ( .C1(n9968), .C2(P1_REG1_REG_15__SCAN_IN), .A(n9967), .B(
        n9966), .ZN(n9969) );
  INV_X1 U11097 ( .A(n9969), .ZN(n9974) );
  AOI211_X1 U11098 ( .C1(n9972), .C2(n9971), .A(n9970), .B(n9986), .ZN(n9973)
         );
  AOI211_X1 U11099 ( .C1(n4395), .C2(n9975), .A(n9974), .B(n9973), .ZN(n9977)
         );
  OAI211_X1 U11100 ( .C1(n9995), .C2(n9978), .A(n9977), .B(n9976), .ZN(
        P1_U3258) );
  INV_X1 U11101 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n9994) );
  INV_X1 U11102 ( .A(n9979), .ZN(n9980) );
  AOI211_X1 U11103 ( .C1(n9983), .C2(n9982), .A(n9981), .B(n9980), .ZN(n9990)
         );
  INV_X1 U11104 ( .A(n9984), .ZN(n9985) );
  AOI211_X1 U11105 ( .C1(n9988), .C2(n9987), .A(n9986), .B(n9985), .ZN(n9989)
         );
  AOI211_X1 U11106 ( .C1(n4395), .C2(n9991), .A(n9990), .B(n9989), .ZN(n9993)
         );
  NAND2_X1 U11107 ( .A1(P1_REG3_REG_18__SCAN_IN), .A2(P1_U3086), .ZN(n9992) );
  OAI211_X1 U11108 ( .C1(n9995), .C2(n9994), .A(n9993), .B(n9992), .ZN(
        P1_U3261) );
  XNOR2_X1 U11109 ( .A(n9997), .B(n9998), .ZN(n10095) );
  NAND2_X1 U11110 ( .A1(n9999), .A2(n9998), .ZN(n10001) );
  AOI21_X1 U11111 ( .B1(n10002), .B2(n10001), .A(n10000), .ZN(n10003) );
  AOI211_X1 U11112 ( .C1(n10005), .C2(n10095), .A(n10004), .B(n10003), .ZN(
        n10092) );
  AOI222_X1 U11113 ( .A1(n10007), .A2(n10042), .B1(P1_REG2_REG_7__SCAN_IN), 
        .B2(n9768), .C1(n10041), .C2(n10006), .ZN(n10013) );
  NOR2_X1 U11114 ( .A1(n9768), .A2(n10008), .ZN(n10047) );
  OAI211_X1 U11115 ( .C1(n10010), .C2(n10091), .A(n10035), .B(n10009), .ZN(
        n10090) );
  INV_X1 U11116 ( .A(n10090), .ZN(n10011) );
  AOI22_X1 U11117 ( .A1(n10095), .A2(n10047), .B1(n10046), .B2(n10011), .ZN(
        n10012) );
  OAI211_X1 U11118 ( .C1(n9768), .C2(n10092), .A(n10013), .B(n10012), .ZN(
        P1_U3286) );
  XNOR2_X1 U11119 ( .A(n10014), .B(n10015), .ZN(n10017) );
  AOI21_X1 U11120 ( .B1(n10017), .B2(n10030), .A(n10016), .ZN(n10078) );
  AOI222_X1 U11121 ( .A1(n6425), .A2(n10042), .B1(P1_REG2_REG_5__SCAN_IN), 
        .B2(n9768), .C1(n10041), .C2(n10018), .ZN(n10026) );
  NAND2_X1 U11122 ( .A1(n10019), .A2(n4993), .ZN(n10021) );
  XNOR2_X1 U11123 ( .A(n10021), .B(n10020), .ZN(n10081) );
  OAI211_X1 U11124 ( .C1(n5341), .C2(n10022), .A(n4392), .B(n10035), .ZN(
        n10077) );
  INV_X1 U11125 ( .A(n10077), .ZN(n10023) );
  AOI22_X1 U11126 ( .A1(n10081), .A2(n10024), .B1(n10046), .B2(n10023), .ZN(
        n10025) );
  OAI211_X1 U11127 ( .C1(n9768), .C2(n10078), .A(n10026), .B(n10025), .ZN(
        P1_U3288) );
  XOR2_X1 U11128 ( .A(n10027), .B(n6419), .Z(n10031) );
  INV_X1 U11129 ( .A(n10028), .ZN(n10029) );
  AOI21_X1 U11130 ( .B1(n10031), .B2(n10030), .A(n10029), .ZN(n10061) );
  XNOR2_X1 U11131 ( .A(n6419), .B(n10032), .ZN(n10064) );
  AOI22_X1 U11132 ( .A1(n10064), .A2(n10033), .B1(P1_REG3_REG_2__SCAN_IN), 
        .B2(n10041), .ZN(n10040) );
  INV_X1 U11133 ( .A(n10034), .ZN(n10037) );
  INV_X1 U11134 ( .A(n7029), .ZN(n10036) );
  OAI211_X1 U11135 ( .C1(n10060), .C2(n10037), .A(n10036), .B(n10035), .ZN(
        n10059) );
  INV_X1 U11136 ( .A(n10059), .ZN(n10038) );
  OAI221_X1 U11137 ( .B1(n9768), .B2(n10061), .C1(n9768), .C2(n10040), .A(
        n10039), .ZN(P1_U3291) );
  AOI222_X1 U11138 ( .A1(n10043), .A2(n10042), .B1(P1_REG2_REG_1__SCAN_IN), 
        .B2(n9768), .C1(n10041), .C2(P1_REG3_REG_1__SCAN_IN), .ZN(n10050) );
  INV_X1 U11139 ( .A(n10044), .ZN(n10045) );
  AOI22_X1 U11140 ( .A1(n10048), .A2(n10047), .B1(n10046), .B2(n10045), .ZN(
        n10049) );
  OAI211_X1 U11141 ( .C1(n9768), .C2(n10051), .A(n10050), .B(n10049), .ZN(
        P1_U3292) );
  AND2_X1 U11142 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n10056), .ZN(P1_U3294) );
  AND2_X1 U11143 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n10056), .ZN(P1_U3295) );
  NOR2_X1 U11144 ( .A1(n10055), .A2(n10052), .ZN(P1_U3296) );
  AND2_X1 U11145 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n10056), .ZN(P1_U3297) );
  AND2_X1 U11146 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n10056), .ZN(P1_U3298) );
  AND2_X1 U11147 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n10056), .ZN(P1_U3299) );
  AND2_X1 U11148 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n10056), .ZN(P1_U3300) );
  AND2_X1 U11149 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n10056), .ZN(P1_U3301) );
  AND2_X1 U11150 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n10056), .ZN(P1_U3302) );
  AND2_X1 U11151 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n10056), .ZN(P1_U3303) );
  AND2_X1 U11152 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n10056), .ZN(P1_U3304) );
  AND2_X1 U11153 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n10056), .ZN(P1_U3305) );
  AND2_X1 U11154 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n10056), .ZN(P1_U3306) );
  NOR2_X1 U11155 ( .A1(n10055), .A2(n10053), .ZN(P1_U3307) );
  NOR2_X1 U11156 ( .A1(n10055), .A2(n10054), .ZN(P1_U3308) );
  AND2_X1 U11157 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n10056), .ZN(P1_U3309) );
  AND2_X1 U11158 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n10056), .ZN(P1_U3310) );
  AND2_X1 U11159 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n10056), .ZN(P1_U3311) );
  AND2_X1 U11160 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n10056), .ZN(P1_U3312) );
  AND2_X1 U11161 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n10056), .ZN(P1_U3313) );
  AND2_X1 U11162 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n10056), .ZN(P1_U3314) );
  AND2_X1 U11163 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n10056), .ZN(P1_U3315) );
  AND2_X1 U11164 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n10056), .ZN(P1_U3316) );
  AND2_X1 U11165 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n10056), .ZN(P1_U3317) );
  AND2_X1 U11166 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n10056), .ZN(P1_U3318) );
  AND2_X1 U11167 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n10056), .ZN(P1_U3319) );
  AND2_X1 U11168 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n10056), .ZN(P1_U3320) );
  AND2_X1 U11169 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n10056), .ZN(P1_U3321) );
  AND2_X1 U11170 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n10056), .ZN(P1_U3322) );
  AND2_X1 U11171 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n10056), .ZN(P1_U3323) );
  INV_X1 U11172 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n10057) );
  AOI22_X1 U11173 ( .A1(n4272), .A2(n10058), .B1(n10057), .B2(n10108), .ZN(
        P1_U3456) );
  OAI21_X1 U11174 ( .B1(n10060), .B2(n10103), .A(n10059), .ZN(n10063) );
  INV_X1 U11175 ( .A(n10061), .ZN(n10062) );
  AOI211_X1 U11176 ( .C1(n10107), .C2(n10064), .A(n10063), .B(n10062), .ZN(
        n10110) );
  AOI22_X1 U11177 ( .A1(n4272), .A2(n10110), .B1(n5248), .B2(n10108), .ZN(
        P1_U3459) );
  OAI21_X1 U11178 ( .B1(n10066), .B2(n10103), .A(n10065), .ZN(n10068) );
  AOI211_X1 U11179 ( .C1(n10107), .C2(n10069), .A(n10068), .B(n10067), .ZN(
        n10111) );
  INV_X1 U11180 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n10070) );
  AOI22_X1 U11181 ( .A1(n4272), .A2(n10111), .B1(n10070), .B2(n10108), .ZN(
        P1_U3462) );
  AOI21_X1 U11182 ( .B1(n10084), .B2(n10072), .A(n10071), .ZN(n10073) );
  OAI211_X1 U11183 ( .C1(n10088), .C2(n10075), .A(n10074), .B(n10073), .ZN(
        n10076) );
  INV_X1 U11184 ( .A(n10076), .ZN(n10113) );
  AOI22_X1 U11185 ( .A1(n4272), .A2(n10113), .B1(n5289), .B2(n10108), .ZN(
        P1_U3465) );
  OAI21_X1 U11186 ( .B1(n5341), .B2(n10103), .A(n10077), .ZN(n10080) );
  INV_X1 U11187 ( .A(n10078), .ZN(n10079) );
  AOI211_X1 U11188 ( .C1(n10107), .C2(n10081), .A(n10080), .B(n10079), .ZN(
        n10114) );
  AOI22_X1 U11189 ( .A1(n4272), .A2(n10114), .B1(n5311), .B2(n10108), .ZN(
        P1_U3468) );
  AOI21_X1 U11190 ( .B1(n10084), .B2(n10083), .A(n10082), .ZN(n10085) );
  OAI211_X1 U11191 ( .C1(n10088), .C2(n10087), .A(n10086), .B(n10085), .ZN(
        n10089) );
  INV_X1 U11192 ( .A(n10089), .ZN(n10117) );
  AOI22_X1 U11193 ( .A1(n4272), .A2(n10117), .B1(n5336), .B2(n10108), .ZN(
        P1_U3471) );
  OAI21_X1 U11194 ( .B1(n10091), .B2(n10103), .A(n10090), .ZN(n10094) );
  INV_X1 U11195 ( .A(n10092), .ZN(n10093) );
  AOI211_X1 U11196 ( .C1(n10096), .C2(n10095), .A(n10094), .B(n10093), .ZN(
        n10119) );
  AOI22_X1 U11197 ( .A1(n4272), .A2(n10119), .B1(n5381), .B2(n10108), .ZN(
        P1_U3474) );
  NAND2_X1 U11198 ( .A1(n10097), .A2(n10107), .ZN(n10098) );
  OAI21_X1 U11199 ( .B1(n4948), .B2(n10103), .A(n10098), .ZN(n10099) );
  NOR2_X1 U11200 ( .A1(n10100), .A2(n10099), .ZN(n10121) );
  AOI22_X1 U11201 ( .A1(n4272), .A2(n10121), .B1(n5348), .B2(n10108), .ZN(
        P1_U3480) );
  OAI211_X1 U11202 ( .C1(n10104), .C2(n10103), .A(n10102), .B(n10101), .ZN(
        n10105) );
  AOI21_X1 U11203 ( .B1(n10107), .B2(n10106), .A(n10105), .ZN(n10123) );
  AOI22_X1 U11204 ( .A1(n4272), .A2(n10123), .B1(n5417), .B2(n10108), .ZN(
        P1_U3483) );
  AOI22_X1 U11205 ( .A1(n10124), .A2(n10110), .B1(n10109), .B2(n10122), .ZN(
        P1_U3524) );
  AOI22_X1 U11206 ( .A1(n10124), .A2(n10111), .B1(n6826), .B2(n10122), .ZN(
        P1_U3525) );
  AOI22_X1 U11207 ( .A1(n10115), .A2(n10113), .B1(n10112), .B2(n10122), .ZN(
        P1_U3526) );
  AOI22_X1 U11208 ( .A1(n10115), .A2(n10114), .B1(n6829), .B2(n10122), .ZN(
        P1_U3527) );
  AOI22_X1 U11209 ( .A1(n10124), .A2(n10117), .B1(n10116), .B2(n10122), .ZN(
        P1_U3528) );
  AOI22_X1 U11210 ( .A1(n10124), .A2(n10119), .B1(n10118), .B2(n10122), .ZN(
        P1_U3529) );
  AOI22_X1 U11211 ( .A1(n10124), .A2(n10121), .B1(n10120), .B2(n10122), .ZN(
        P1_U3531) );
  AOI22_X1 U11212 ( .A1(n10124), .A2(n10123), .B1(n7114), .B2(n10122), .ZN(
        P1_U3532) );
  NAND2_X1 U11213 ( .A1(n10125), .A2(n4269), .ZN(n10138) );
  NAND2_X1 U11214 ( .A1(n10126), .A2(n10221), .ZN(n10127) );
  NAND2_X1 U11215 ( .A1(n10154), .A2(n10127), .ZN(n10128) );
  NAND2_X1 U11216 ( .A1(n10129), .A2(n10128), .ZN(n10137) );
  XNOR2_X1 U11217 ( .A(n10131), .B(n10130), .ZN(n10132) );
  OR2_X1 U11218 ( .A1(n10133), .A2(n10132), .ZN(n10136) );
  INV_X1 U11219 ( .A(n10134), .ZN(n10135) );
  AND4_X1 U11220 ( .A1(n10138), .A2(n10137), .A3(n10136), .A4(n10135), .ZN(
        n10145) );
  OAI21_X1 U11221 ( .B1(n10141), .B2(n10140), .A(n10139), .ZN(n10143) );
  AOI22_X1 U11222 ( .A1(n10143), .A2(n10166), .B1(n10142), .B2(
        P2_ADDR_REG_3__SCAN_IN), .ZN(n10144) );
  NAND2_X1 U11223 ( .A1(n10145), .A2(n10144), .ZN(P2_U3185) );
  XOR2_X1 U11224 ( .A(n10146), .B(n10147), .Z(n10167) );
  OAI21_X1 U11225 ( .B1(n10150), .B2(n10149), .A(n10148), .ZN(n10159) );
  INV_X1 U11226 ( .A(n10151), .ZN(n10153) );
  NAND3_X1 U11227 ( .A1(n10154), .A2(n10153), .A3(n10152), .ZN(n10156) );
  AOI21_X1 U11228 ( .B1(n10157), .B2(n10156), .A(n10155), .ZN(n10158) );
  AOI21_X1 U11229 ( .B1(n10160), .B2(n10159), .A(n10158), .ZN(n10162) );
  OAI211_X1 U11230 ( .C1(n10164), .C2(n10163), .A(n10162), .B(n10161), .ZN(
        n10165) );
  AOI21_X1 U11231 ( .B1(n10167), .B2(n10166), .A(n10165), .ZN(n10168) );
  OAI21_X1 U11232 ( .B1(n10170), .B2(n10169), .A(n10168), .ZN(P2_U3186) );
  XNOR2_X1 U11233 ( .A(n10172), .B(n10171), .ZN(n10177) );
  AOI222_X1 U11234 ( .A1(n10178), .A2(n10177), .B1(n10176), .B2(n10175), .C1(
        n10174), .C2(n10173), .ZN(n10204) );
  XNOR2_X1 U11235 ( .A(n10179), .B(n10180), .ZN(n10202) );
  AOI222_X1 U11236 ( .A1(n10184), .A2(n10183), .B1(n10202), .B2(n10182), .C1(
        n10200), .C2(n10181), .ZN(n10185) );
  OAI221_X1 U11237 ( .B1(n10187), .B2(n10204), .C1(n10186), .C2(n6951), .A(
        n10185), .ZN(P2_U3229) );
  AOI22_X1 U11238 ( .A1(n10219), .A2(n5932), .B1(n10188), .B2(n10217), .ZN(
        P2_U3393) );
  INV_X1 U11239 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n10193) );
  AOI22_X1 U11240 ( .A1(n10190), .A2(n4391), .B1(n10216), .B2(n10189), .ZN(
        n10191) );
  AND2_X1 U11241 ( .A1(n10192), .A2(n10191), .ZN(n10220) );
  AOI22_X1 U11242 ( .A1(n10219), .A2(n10193), .B1(n10220), .B2(n10217), .ZN(
        P2_U3396) );
  INV_X1 U11243 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n10199) );
  OR2_X1 U11244 ( .A1(n10194), .A2(n10210), .ZN(n10197) );
  NAND2_X1 U11245 ( .A1(n10195), .A2(n10216), .ZN(n10196) );
  AND3_X1 U11246 ( .A1(n10198), .A2(n10197), .A3(n10196), .ZN(n10222) );
  AOI22_X1 U11247 ( .A1(n10219), .A2(n10199), .B1(n10222), .B2(n10217), .ZN(
        P2_U3399) );
  AOI22_X1 U11248 ( .A1(n10202), .A2(n10201), .B1(n10216), .B2(n10200), .ZN(
        n10203) );
  AND2_X1 U11249 ( .A1(n10204), .A2(n10203), .ZN(n10224) );
  AOI22_X1 U11250 ( .A1(n10219), .A2(n5975), .B1(n10224), .B2(n10217), .ZN(
        P2_U3402) );
  AOI22_X1 U11251 ( .A1(n10206), .A2(n4391), .B1(n10216), .B2(n10205), .ZN(
        n10207) );
  AND2_X1 U11252 ( .A1(n10208), .A2(n10207), .ZN(n10226) );
  AOI22_X1 U11253 ( .A1(n10219), .A2(n10209), .B1(n10226), .B2(n10217), .ZN(
        P2_U3405) );
  INV_X1 U11254 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10218) );
  NOR2_X1 U11255 ( .A1(n10211), .A2(n10210), .ZN(n10214) );
  INV_X1 U11256 ( .A(n10212), .ZN(n10213) );
  AOI211_X1 U11257 ( .C1(n10216), .C2(n10215), .A(n10214), .B(n10213), .ZN(
        n10228) );
  AOI22_X1 U11258 ( .A1(n10219), .A2(n10218), .B1(n10228), .B2(n10217), .ZN(
        P2_U3408) );
  AOI22_X1 U11259 ( .A1(n10229), .A2(n10220), .B1(n6878), .B2(n10227), .ZN(
        P2_U3461) );
  AOI22_X1 U11260 ( .A1(n10229), .A2(n10222), .B1(n10221), .B2(n10227), .ZN(
        P2_U3462) );
  AOI22_X1 U11261 ( .A1(n10229), .A2(n10224), .B1(n10223), .B2(n10227), .ZN(
        P2_U3463) );
  AOI22_X1 U11262 ( .A1(n10229), .A2(n10226), .B1(n10225), .B2(n10227), .ZN(
        P2_U3464) );
  AOI22_X1 U11263 ( .A1(n10229), .A2(n10228), .B1(n7178), .B2(n10227), .ZN(
        P2_U3465) );
  NOR2_X1 U11264 ( .A1(n10231), .A2(n10230), .ZN(n10232) );
  XOR2_X1 U11265 ( .A(P2_ADDR_REG_1__SCAN_IN), .B(n10232), .Z(ADD_1068_U5) );
  XOR2_X1 U11266 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1068_U46) );
  NOR2_X1 U11267 ( .A1(n10234), .A2(n10233), .ZN(n10235) );
  XOR2_X1 U11268 ( .A(P2_ADDR_REG_18__SCAN_IN), .B(n10235), .Z(ADD_1068_U55)
         );
  XNOR2_X1 U11269 ( .A(n10237), .B(n10236), .ZN(ADD_1068_U56) );
  XNOR2_X1 U11270 ( .A(n10239), .B(n10238), .ZN(ADD_1068_U57) );
  XNOR2_X1 U11271 ( .A(n10241), .B(n10240), .ZN(ADD_1068_U58) );
  XNOR2_X1 U11272 ( .A(n10243), .B(n10242), .ZN(ADD_1068_U59) );
  XNOR2_X1 U11273 ( .A(n10245), .B(n10244), .ZN(ADD_1068_U60) );
  XNOR2_X1 U11274 ( .A(n10247), .B(n10246), .ZN(ADD_1068_U61) );
  XNOR2_X1 U11275 ( .A(n10249), .B(n10248), .ZN(ADD_1068_U62) );
  XNOR2_X1 U11276 ( .A(n10251), .B(n10250), .ZN(ADD_1068_U63) );
  XNOR2_X1 U11277 ( .A(n10253), .B(n10252), .ZN(ADD_1068_U50) );
  XNOR2_X1 U11278 ( .A(n10255), .B(n10254), .ZN(ADD_1068_U51) );
  XNOR2_X1 U11279 ( .A(n10257), .B(n10256), .ZN(ADD_1068_U47) );
  XNOR2_X1 U11280 ( .A(n10259), .B(n10258), .ZN(ADD_1068_U49) );
  XNOR2_X1 U11281 ( .A(n10261), .B(n10260), .ZN(ADD_1068_U48) );
  XOR2_X1 U11282 ( .A(n10263), .B(n10262), .Z(ADD_1068_U54) );
  XOR2_X1 U11283 ( .A(n10265), .B(n10264), .Z(ADD_1068_U53) );
  XNOR2_X1 U11284 ( .A(n10267), .B(n10266), .ZN(ADD_1068_U52) );
  BUF_X1 U4785 ( .A(n5151), .Z(n8003) );
  BUF_X2 U4903 ( .A(n5323), .Z(n5510) );
  CLKBUF_X3 U4788 ( .A(n7036), .Z(n7904) );
  NAND2_X1 U4795 ( .A1(n8414), .A2(n8413), .ZN(n8415) );
  AND2_X1 U4813 ( .A1(n9272), .A2(n7868), .ZN(n7871) );
  NAND3_X1 U4848 ( .A1(n4835), .A2(P2_REG1_REG_7__SCAN_IN), .A3(n7274), .ZN(
        n7276) );
  CLKBUF_X1 U4888 ( .A(n9312), .Z(n4468) );
  CLKBUF_X2 U4968 ( .A(n5310), .Z(n5697) );
  NAND2_X1 U4976 ( .A1(n4277), .A2(n6658), .ZN(n5678) );
  NOR2_X2 U5078 ( .A1(n9758), .A2(n9882), .ZN(n9744) );
  NAND2_X1 U5356 ( .A1(n8232), .A2(n9389), .ZN(n6678) );
  CLKBUF_X1 U5652 ( .A(n6295), .Z(n8287) );
  CLKBUF_X1 U6281 ( .A(n5312), .Z(n5699) );
  OAI21_X1 U6288 ( .B1(n6678), .B2(n9391), .A(n5277), .ZN(n6986) );
endmodule

