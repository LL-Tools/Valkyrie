

module b15_C_AntiSAT_k_256_3 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, 
        READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, 
        CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, 
        REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, 
        FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, 
        keyinput128, keyinput129, keyinput130, keyinput131, keyinput132, 
        keyinput133, keyinput134, keyinput135, keyinput136, keyinput137, 
        keyinput138, keyinput139, keyinput140, keyinput141, keyinput142, 
        keyinput143, keyinput144, keyinput145, keyinput146, keyinput147, 
        keyinput148, keyinput149, keyinput150, keyinput151, keyinput152, 
        keyinput153, keyinput154, keyinput155, keyinput156, keyinput157, 
        keyinput158, keyinput159, keyinput160, keyinput161, keyinput162, 
        keyinput163, keyinput164, keyinput165, keyinput166, keyinput167, 
        keyinput168, keyinput169, keyinput170, keyinput171, keyinput172, 
        keyinput173, keyinput174, keyinput175, keyinput176, keyinput177, 
        keyinput178, keyinput179, keyinput180, keyinput181, keyinput182, 
        keyinput183, keyinput184, keyinput185, keyinput186, keyinput187, 
        keyinput188, keyinput189, keyinput190, keyinput191, keyinput192, 
        keyinput193, keyinput194, keyinput195, keyinput196, keyinput197, 
        keyinput198, keyinput199, keyinput200, keyinput201, keyinput202, 
        keyinput203, keyinput204, keyinput205, keyinput206, keyinput207, 
        keyinput208, keyinput209, keyinput210, keyinput211, keyinput212, 
        keyinput213, keyinput214, keyinput215, keyinput216, keyinput217, 
        keyinput218, keyinput219, keyinput220, keyinput221, keyinput222, 
        keyinput223, keyinput224, keyinput225, keyinput226, keyinput227, 
        keyinput228, keyinput229, keyinput230, keyinput231, keyinput232, 
        keyinput233, keyinput234, keyinput235, keyinput236, keyinput237, 
        keyinput238, keyinput239, keyinput240, keyinput241, keyinput242, 
        keyinput243, keyinput244, keyinput245, keyinput246, keyinput247, 
        keyinput248, keyinput249, keyinput250, keyinput251, keyinput252, 
        keyinput253, keyinput254, keyinput255, U3445, U3446, U3447, U3448, 
        U3213, U3212, U3211, U3210, U3209, U3208, U3207, U3206, U3205, U3204, 
        U3203, U3202, U3201, U3200, U3199, U3198, U3197, U3196, U3195, U3194, 
        U3193, U3192, U3191, U3190, U3189, U3188, U3187, U3186, U3185, U3184, 
        U3183, U3182, U3181, U3451, U3452, U3180, U3179, U3178, U3177, U3176, 
        U3175, U3174, U3173, U3172, U3171, U3170, U3169, U3168, U3167, U3166, 
        U3165, U3164, U3163, U3162, U3161, U3160, U3159, U3158, U3157, U3156, 
        U3155, U3154, U3153, U3152, U3151, U3453, U3150, U3149, U3148, U3147, 
        U3146, U3145, U3144, U3143, U3142, U3141, U3140, U3139, U3138, U3137, 
        U3136, U3135, U3134, U3133, U3132, U3131, U3130, U3129, U3128, U3127, 
        U3126, U3125, U3124, U3123, U3122, U3121, U3120, U3119, U3118, U3117, 
        U3116, U3115, U3114, U3113, U3112, U3111, U3110, U3109, U3108, U3107, 
        U3106, U3105, U3104, U3103, U3102, U3101, U3100, U3099, U3098, U3097, 
        U3096, U3095, U3094, U3093, U3092, U3091, U3090, U3089, U3088, U3087, 
        U3086, U3085, U3084, U3083, U3082, U3081, U3080, U3079, U3078, U3077, 
        U3076, U3075, U3074, U3073, U3072, U3071, U3070, U3069, U3068, U3067, 
        U3066, U3065, U3064, U3063, U3062, U3061, U3060, U3059, U3058, U3057, 
        U3056, U3055, U3054, U3053, U3052, U3051, U3050, U3049, U3048, U3047, 
        U3046, U3045, U3044, U3043, U3042, U3041, U3040, U3039, U3038, U3037, 
        U3036, U3035, U3034, U3033, U3032, U3031, U3030, U3029, U3028, U3027, 
        U3026, U3025, U3024, U3023, U3022, U3021, U3020, U3455, U3456, U3459, 
        U3460, U3461, U3019, U3462, U3463, U3464, U3465, U3018, U3017, U3016, 
        U3015, U3014, U3013, U3012, U3011, U3010, U3009, U3008, U3007, U3006, 
        U3005, U3004, U3003, U3002, U3001, U3000, U2999, U2998, U2997, U2996, 
        U2995, U2994, U2993, U2992, U2991, U2990, U2989, U2988, U2987, U2986, 
        U2985, U2984, U2983, U2982, U2981, U2980, U2979, U2978, U2977, U2976, 
        U2975, U2974, U2973, U2972, U2971, U2970, U2969, U2968, U2967, U2966, 
        U2965, U2964, U2963, U2962, U2961, U2960, U2959, U2958, U2957, U2956, 
        U2955, U2954, U2953, U2952, U2951, U2950, U2949, U2948, U2947, U2946, 
        U2945, U2944, U2943, U2942, U2941, U2940, U2939, U2938, U2937, U2936, 
        U2935, U2934, U2933, U2932, U2931, U2930, U2929, U2928, U2927, U2926, 
        U2925, U2924, U2923, U2922, U2921, U2920, U2919, U2918, U2917, U2916, 
        U2915, U2914, U2913, U2912, U2911, U2910, U2909, U2908, U2907, U2906, 
        U2905, U2904, U2903, U2902, U2901, U2900, U2899, U2898, U2897, U2896, 
        U2895, U2894, U2893, U2892, U2891, U2890, U2889, U2888, U2887, U2886, 
        U2885, U2884, U2883, U2882, U2881, U2880, U2879, U2878, U2877, U2876, 
        U2875, U2874, U2873, U2872, U2871, U2870, U2869, U2868, U2867, U2866, 
        U2865, U2864, U2863, U2862, U2861, U2860, U2859, U2858, U2857, U2856, 
        U2855, U2854, U2853, U2852, U2851, U2850, U2849, U2848, U2847, U2846, 
        U2845, U2844, U2843, U2842, U2841, U2840, U2839, U2838, U2837, U2836, 
        U2835, U2834, U2833, U2832, U2831, U2830, U2829, U2828, U2827, U2826, 
        U2825, U2824, U2823, U2822, U2821, U2820, U2819, U2818, U2817, U2816, 
        U2815, U2814, U2813, U2812, U2811, U2810, U2809, U2808, U2807, U2806, 
        U2805, U2804, U2803, U2802, U2801, U2800, U2799, U2798, U2797, U2796, 
        U2795, U3468, U2794, U3469, U3470, U2793, U3471, U2792, U3472, U2791, 
        U3473, U2790, U2789, U3474, U2788 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
         READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
         M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
         STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
         W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput0, keyinput1,
         keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7,
         keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13,
         keyinput14, keyinput15, keyinput16, keyinput17, keyinput18,
         keyinput19, keyinput20, keyinput21, keyinput22, keyinput23,
         keyinput24, keyinput25, keyinput26, keyinput27, keyinput28,
         keyinput29, keyinput30, keyinput31, keyinput32, keyinput33,
         keyinput34, keyinput35, keyinput36, keyinput37, keyinput38,
         keyinput39, keyinput40, keyinput41, keyinput42, keyinput43,
         keyinput44, keyinput45, keyinput46, keyinput47, keyinput48,
         keyinput49, keyinput50, keyinput51, keyinput52, keyinput53,
         keyinput54, keyinput55, keyinput56, keyinput57, keyinput58,
         keyinput59, keyinput60, keyinput61, keyinput62, keyinput63,
         keyinput64, keyinput65, keyinput66, keyinput67, keyinput68,
         keyinput69, keyinput70, keyinput71, keyinput72, keyinput73,
         keyinput74, keyinput75, keyinput76, keyinput77, keyinput78,
         keyinput79, keyinput80, keyinput81, keyinput82, keyinput83,
         keyinput84, keyinput85, keyinput86, keyinput87, keyinput88,
         keyinput89, keyinput90, keyinput91, keyinput92, keyinput93,
         keyinput94, keyinput95, keyinput96, keyinput97, keyinput98,
         keyinput99, keyinput100, keyinput101, keyinput102, keyinput103,
         keyinput104, keyinput105, keyinput106, keyinput107, keyinput108,
         keyinput109, keyinput110, keyinput111, keyinput112, keyinput113,
         keyinput114, keyinput115, keyinput116, keyinput117, keyinput118,
         keyinput119, keyinput120, keyinput121, keyinput122, keyinput123,
         keyinput124, keyinput125, keyinput126, keyinput127, keyinput128,
         keyinput129, keyinput130, keyinput131, keyinput132, keyinput133,
         keyinput134, keyinput135, keyinput136, keyinput137, keyinput138,
         keyinput139, keyinput140, keyinput141, keyinput142, keyinput143,
         keyinput144, keyinput145, keyinput146, keyinput147, keyinput148,
         keyinput149, keyinput150, keyinput151, keyinput152, keyinput153,
         keyinput154, keyinput155, keyinput156, keyinput157, keyinput158,
         keyinput159, keyinput160, keyinput161, keyinput162, keyinput163,
         keyinput164, keyinput165, keyinput166, keyinput167, keyinput168,
         keyinput169, keyinput170, keyinput171, keyinput172, keyinput173,
         keyinput174, keyinput175, keyinput176, keyinput177, keyinput178,
         keyinput179, keyinput180, keyinput181, keyinput182, keyinput183,
         keyinput184, keyinput185, keyinput186, keyinput187, keyinput188,
         keyinput189, keyinput190, keyinput191, keyinput192, keyinput193,
         keyinput194, keyinput195, keyinput196, keyinput197, keyinput198,
         keyinput199, keyinput200, keyinput201, keyinput202, keyinput203,
         keyinput204, keyinput205, keyinput206, keyinput207, keyinput208,
         keyinput209, keyinput210, keyinput211, keyinput212, keyinput213,
         keyinput214, keyinput215, keyinput216, keyinput217, keyinput218,
         keyinput219, keyinput220, keyinput221, keyinput222, keyinput223,
         keyinput224, keyinput225, keyinput226, keyinput227, keyinput228,
         keyinput229, keyinput230, keyinput231, keyinput232, keyinput233,
         keyinput234, keyinput235, keyinput236, keyinput237, keyinput238,
         keyinput239, keyinput240, keyinput241, keyinput242, keyinput243,
         keyinput244, keyinput245, keyinput246, keyinput247, keyinput248,
         keyinput249, keyinput250, keyinput251, keyinput252, keyinput253,
         keyinput254, keyinput255;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185,
         n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195,
         n3196, n3197, n3198, n3199, n3200, n3201, n3203, n3204, n3205, n3206,
         n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216,
         n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226,
         n3227, n3228, n3229, n3232, n3233, n3234, n3235, n3236, n3237, n3238,
         n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248,
         n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258,
         n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268,
         n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278,
         n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288,
         n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298,
         n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308,
         n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318,
         n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328,
         n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338,
         n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348,
         n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358,
         n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368,
         n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378,
         n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388,
         n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398,
         n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408,
         n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418,
         n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428,
         n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438,
         n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448,
         n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458,
         n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468,
         n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478,
         n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488,
         n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498,
         n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508,
         n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518,
         n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528,
         n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538,
         n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548,
         n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558,
         n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568,
         n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578,
         n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588,
         n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598,
         n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608,
         n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618,
         n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628,
         n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638,
         n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648,
         n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658,
         n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668,
         n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678,
         n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688,
         n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698,
         n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708,
         n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718,
         n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728,
         n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738,
         n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748,
         n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758,
         n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768,
         n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778,
         n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788,
         n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798,
         n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808,
         n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818,
         n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828,
         n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838,
         n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848,
         n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858,
         n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868,
         n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878,
         n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888,
         n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898,
         n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908,
         n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918,
         n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928,
         n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938,
         n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948,
         n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958,
         n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968,
         n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978,
         n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988,
         n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998,
         n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008,
         n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018,
         n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028,
         n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038,
         n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048,
         n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058,
         n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068,
         n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078,
         n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088,
         n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098,
         n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108,
         n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118,
         n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128,
         n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138,
         n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148,
         n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158,
         n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168,
         n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178,
         n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188,
         n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198,
         n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208,
         n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218,
         n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228,
         n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238,
         n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248,
         n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258,
         n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268,
         n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278,
         n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288,
         n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298,
         n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308,
         n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318,
         n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328,
         n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338,
         n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348,
         n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358,
         n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368,
         n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378,
         n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388,
         n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398,
         n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408,
         n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418,
         n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428,
         n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438,
         n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448,
         n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458,
         n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468,
         n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478,
         n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488,
         n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498,
         n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508,
         n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518,
         n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528,
         n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538,
         n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548,
         n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558,
         n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568,
         n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578,
         n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588,
         n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598,
         n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608,
         n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4617, n4618, n4619,
         n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629,
         n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639,
         n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649,
         n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659,
         n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669,
         n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679,
         n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689,
         n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699,
         n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709,
         n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719,
         n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729,
         n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739,
         n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749,
         n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759,
         n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769,
         n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779,
         n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789,
         n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799,
         n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809,
         n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819,
         n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829,
         n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839,
         n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849,
         n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859,
         n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869,
         n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879,
         n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889,
         n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899,
         n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909,
         n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919,
         n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929,
         n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939,
         n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949,
         n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959,
         n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969,
         n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979,
         n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989,
         n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999,
         n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009,
         n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019,
         n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029,
         n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039,
         n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049,
         n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059,
         n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069,
         n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079,
         n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089,
         n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099,
         n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109,
         n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119,
         n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129,
         n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139,
         n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149,
         n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159,
         n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169,
         n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179,
         n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189,
         n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199,
         n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209,
         n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219,
         n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229,
         n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239,
         n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249,
         n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259,
         n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269,
         n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279,
         n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289,
         n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299,
         n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309,
         n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319,
         n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329,
         n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339,
         n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349,
         n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359,
         n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369,
         n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379,
         n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389,
         n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399,
         n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409,
         n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419,
         n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429,
         n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439,
         n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449,
         n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459,
         n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469,
         n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479,
         n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489,
         n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499,
         n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509,
         n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519,
         n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529,
         n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539,
         n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549,
         n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559,
         n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569,
         n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579,
         n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589,
         n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599,
         n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609,
         n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619,
         n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629,
         n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639,
         n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649,
         n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659,
         n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669,
         n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679,
         n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689,
         n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699,
         n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709,
         n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719,
         n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729,
         n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739,
         n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749,
         n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759,
         n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769,
         n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779,
         n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789,
         n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799,
         n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809,
         n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819,
         n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829,
         n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839,
         n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849,
         n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859,
         n5860, n5861, n5862, n5863, n5864, n5866, n5867, n5868, n5869, n5870,
         n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880,
         n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890,
         n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900,
         n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910,
         n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920,
         n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930,
         n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940,
         n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950,
         n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960,
         n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970,
         n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980,
         n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990,
         n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000,
         n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010,
         n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020,
         n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030,
         n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040,
         n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050,
         n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060,
         n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070,
         n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080,
         n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090,
         n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100,
         n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110,
         n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120,
         n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130,
         n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140,
         n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150,
         n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160,
         n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170,
         n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180,
         n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190,
         n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200,
         n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210,
         n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220,
         n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230,
         n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240,
         n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250,
         n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260,
         n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270,
         n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280,
         n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290,
         n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300,
         n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310,
         n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320,
         n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330,
         n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340,
         n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350,
         n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360,
         n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370,
         n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380,
         n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390,
         n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400,
         n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410,
         n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420,
         n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430,
         n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440,
         n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450,
         n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460,
         n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470,
         n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480,
         n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490,
         n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500,
         n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510,
         n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520,
         n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530,
         n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540,
         n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550,
         n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560,
         n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570,
         n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580,
         n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590,
         n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600,
         n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610,
         n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620,
         n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630,
         n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640,
         n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650,
         n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660,
         n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670,
         n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680,
         n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690,
         n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700,
         n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710,
         n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720,
         n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730,
         n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740,
         n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750,
         n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760,
         n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770,
         n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780,
         n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790,
         n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800,
         n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810,
         n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820,
         n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830,
         n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840,
         n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850,
         n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860,
         n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870,
         n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880,
         n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890,
         n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900,
         n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910,
         n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920,
         n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930,
         n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940,
         n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950,
         n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960,
         n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970,
         n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980,
         n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990,
         n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000,
         n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010,
         n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020,
         n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030,
         n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038;

  INV_X2 U3624 ( .A(n6476), .ZN(n5989) );
  AND2_X1 U3625 ( .A1(n3507), .A2(n3506), .ZN(n3573) );
  CLKBUF_X2 U3626 ( .A(n3398), .Z(n4192) );
  CLKBUF_X2 U3627 ( .A(n3395), .Z(n3945) );
  CLKBUF_X2 U3628 ( .A(n3523), .Z(n3207) );
  CLKBUF_X2 U3629 ( .A(n3469), .Z(n4186) );
  AND4_X1 U3630 ( .A1(n3376), .A2(n3375), .A3(n3374), .A4(n3373), .ZN(n3214)
         );
  OR2_X2 U3631 ( .A1(n3368), .A2(n3367), .ZN(n3446) );
  AND2_X1 U3632 ( .A1(n3300), .A2(n4887), .ZN(n3469) );
  AND2_X2 U3633 ( .A1(n3297), .A2(n3299), .ZN(n3399) );
  AND2_X1 U3634 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n5032) );
  AND2_X2 U3635 ( .A1(n3299), .A2(n4887), .ZN(n3396) );
  AND2_X2 U3636 ( .A1(n4880), .A2(n5032), .ZN(n3524) );
  AND4_X1 U3637 ( .A1(n3316), .A2(n3315), .A3(n3314), .A4(n3313), .ZN(n3322)
         );
  NAND3_X1 U3638 ( .A1(n5892), .A2(n4999), .A3(n6199), .ZN(n4728) );
  AND2_X1 U3639 ( .A1(n3443), .A2(n3442), .ZN(n4603) );
  CLKBUF_X2 U3640 ( .A(n3388), .Z(n3474) );
  INV_X1 U3641 ( .A(n3444), .ZN(n5234) );
  INV_X1 U3642 ( .A(n6267), .ZN(n6261) );
  NOR2_X1 U3643 ( .A1(n5864), .A2(n4693), .ZN(n5727) );
  INV_X1 U3644 ( .A(n3446), .ZN(n5216) );
  NAND2_X1 U3645 ( .A1(n5567), .A2(n5569), .ZN(n5568) );
  INV_X2 U3646 ( .A(n3179), .ZN(n6523) );
  INV_X1 U3647 ( .A(n6201), .ZN(n6185) );
  AND2_X1 U3649 ( .A1(n4887), .A2(n5032), .ZN(n3388) );
  AND4_X1 U3650 ( .A1(n3240), .A2(n3239), .A3(n3385), .A4(n3238), .ZN(n3176)
         );
  AND2_X2 U3651 ( .A1(n4888), .A2(n5032), .ZN(n3523) );
  INV_X2 U3652 ( .A(n7038), .ZN(n3206) );
  NAND2_X4 U3653 ( .A1(n3679), .A2(n3682), .ZN(n3704) );
  BUF_X8 U3654 ( .A(n3704), .Z(n3211) );
  NAND2_X2 U3655 ( .A1(n5242), .A2(n5243), .ZN(n3689) );
  NAND2_X2 U3656 ( .A1(n3678), .A2(n3677), .ZN(n5242) );
  XNOR2_X2 U3657 ( .A(n5004), .B(n6573), .ZN(n4969) );
  AND2_X2 U3658 ( .A1(n6495), .A2(n3604), .ZN(n4915) );
  NAND2_X2 U3659 ( .A1(n3383), .A2(n3382), .ZN(n3441) );
  NOR2_X2 U3660 ( .A1(n4733), .A2(n4734), .ZN(n3765) );
  NAND2_X1 U3661 ( .A1(n3406), .A2(n3378), .ZN(n3763) );
  XNOR2_X2 U3662 ( .A(n3616), .B(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4906)
         );
  NAND2_X4 U3663 ( .A1(n3597), .A2(n3596), .ZN(n3774) );
  NOR2_X2 U3664 ( .A1(n3647), .A2(n3646), .ZN(n3660) );
  INV_X2 U3665 ( .A(n3211), .ZN(n5633) );
  OR2_X1 U3666 ( .A1(n5550), .A2(n5549), .ZN(n6060) );
  INV_X2 U3667 ( .A(n6365), .ZN(n6358) );
  NAND2_X1 U3668 ( .A1(n4708), .A2(n4635), .ZN(n4710) );
  AND2_X1 U3669 ( .A1(n3712), .A2(n4611), .ZN(n3749) );
  CLKBUF_X1 U3670 ( .A(n4635), .Z(n3205) );
  INV_X1 U3671 ( .A(n7038), .ZN(n3177) );
  INV_X1 U3672 ( .A(n3456), .ZN(n4611) );
  INV_X2 U3673 ( .A(n3429), .ZN(n3714) );
  BUF_X1 U3674 ( .A(n3406), .Z(n3710) );
  AND4_X1 U3675 ( .A1(n3330), .A2(n3329), .A3(n3328), .A4(n3327), .ZN(n3336)
         );
  CLKBUF_X2 U3676 ( .A(n3399), .Z(n4196) );
  NOR2_X1 U3677 ( .A1(n3195), .A2(n4766), .ZN(n4767) );
  CLKBUF_X1 U3678 ( .A(n5797), .Z(n5798) );
  AND2_X2 U3679 ( .A1(n3181), .A2(n3182), .ZN(n3191) );
  NOR2_X2 U3680 ( .A1(n4039), .A2(n4038), .ZN(n4072) );
  CLKBUF_X1 U3681 ( .A(n5853), .Z(n5854) );
  AND2_X1 U3682 ( .A1(n5504), .A2(n3256), .ZN(n5543) );
  AND2_X1 U3683 ( .A1(n5504), .A2(n3256), .ZN(n3192) );
  CLKBUF_X1 U3684 ( .A(n5098), .Z(n5270) );
  AND2_X1 U3685 ( .A1(n3485), .A2(n3484), .ZN(n3510) );
  AND2_X1 U3686 ( .A1(n3414), .A2(n4883), .ZN(n3435) );
  AND3_X1 U3687 ( .A1(n3377), .A2(n3446), .A3(n3431), .ZN(n3383) );
  INV_X1 U3688 ( .A(n4635), .ZN(n6250) );
  NAND2_X1 U3689 ( .A1(n3456), .A2(STATE2_REG_0__SCAN_IN), .ZN(n5259) );
  INV_X1 U3690 ( .A(n3378), .ZN(n3325) );
  BUF_X2 U3691 ( .A(n3834), .Z(n4195) );
  CLKBUF_X2 U3692 ( .A(n3524), .Z(n4184) );
  BUF_X2 U3693 ( .A(n3386), .Z(n3208) );
  BUF_X2 U3694 ( .A(n3396), .Z(n4183) );
  CLKBUF_X3 U3695 ( .A(n3386), .Z(n4182) );
  CLKBUF_X1 U3696 ( .A(n3213), .Z(n3178) );
  CLKBUF_X2 U3697 ( .A(n3397), .Z(n4167) );
  AND2_X2 U3698 ( .A1(n3289), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3297)
         );
  XNOR2_X1 U3699 ( .A(n4234), .B(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n5645)
         );
  XNOR2_X1 U3700 ( .A(n4584), .B(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n4765)
         );
  AOI21_X1 U3701 ( .B1(n4250), .B2(n5989), .A(n4249), .ZN(n4251) );
  CLKBUF_X1 U3702 ( .A(n4241), .Z(n5962) );
  INV_X1 U3703 ( .A(n5790), .ZN(n5931) );
  XNOR2_X1 U3704 ( .A(n5605), .B(n5606), .ZN(n5927) );
  INV_X1 U3705 ( .A(n3191), .ZN(n5737) );
  NOR2_X1 U3706 ( .A1(n4807), .A2(n4806), .ZN(n4808) );
  NAND2_X1 U3707 ( .A1(n3696), .A2(n3695), .ZN(n5513) );
  AND2_X1 U3708 ( .A1(n5669), .A2(n4727), .ZN(n5902) );
  NAND2_X1 U3709 ( .A1(n5685), .A2(n4726), .ZN(n5669) );
  AND2_X1 U3710 ( .A1(n3695), .A2(n3190), .ZN(n3189) );
  OAI21_X1 U3711 ( .B1(n3278), .B2(n3688), .A(n3279), .ZN(n3277) );
  XNOR2_X1 U3712 ( .A(n3687), .B(n5250), .ZN(n5243) );
  NOR2_X1 U3713 ( .A1(n6945), .A2(n6142), .ZN(n6126) );
  OAI21_X1 U3714 ( .B1(n3821), .B2(n3820), .A(n3819), .ZN(n5257) );
  NAND2_X1 U3715 ( .A1(n3815), .A2(n3814), .ZN(n5271) );
  OR2_X1 U3716 ( .A1(n4747), .A2(n6872), .ZN(n4929) );
  AND2_X1 U3717 ( .A1(n4815), .A2(n4810), .ZN(n7036) );
  BUF_X2 U3718 ( .A(n3768), .Z(n4966) );
  OR2_X1 U3719 ( .A1(n4852), .A2(n4851), .ZN(n4854) );
  NAND2_X1 U3720 ( .A1(n3550), .A2(n3549), .ZN(n5042) );
  NAND2_X1 U3721 ( .A1(n3228), .A2(n3227), .ZN(n6179) );
  CLKBUF_X1 U3722 ( .A(n4969), .Z(n6636) );
  NAND2_X1 U3723 ( .A1(n3532), .A2(n3531), .ZN(n3572) );
  INV_X1 U3724 ( .A(n5125), .ZN(n3228) );
  NAND2_X1 U3725 ( .A1(n3229), .A2(n4643), .ZN(n5125) );
  CLKBUF_X1 U3726 ( .A(n4968), .Z(n3210) );
  INV_X1 U3727 ( .A(n4941), .ZN(n3229) );
  AND3_X1 U3728 ( .A1(n3780), .A2(n3779), .A3(n3778), .ZN(n4851) );
  NAND2_X1 U3729 ( .A1(n3420), .A2(n3419), .ZN(n3485) );
  INV_X1 U3730 ( .A(n5124), .ZN(n3227) );
  INV_X1 U3731 ( .A(n4940), .ZN(n4643) );
  NAND2_X1 U3732 ( .A1(n3441), .A2(n6199), .ZN(n3421) );
  NAND2_X1 U3733 ( .A1(n6250), .A2(n3206), .ZN(n4713) );
  NAND2_X1 U3734 ( .A1(n5892), .A2(n3217), .ZN(n5021) );
  NAND2_X1 U3735 ( .A1(n3518), .A2(n5259), .ZN(n3755) );
  MUX2_X1 U3736 ( .A(n3498), .B(n3680), .S(n3501), .Z(n3595) );
  AND2_X1 U3737 ( .A1(n3444), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3712) );
  INV_X1 U3738 ( .A(n3599), .ZN(n3501) );
  AND2_X1 U3740 ( .A1(n4988), .A2(n3426), .ZN(n5892) );
  OR2_X1 U3741 ( .A1(n3467), .A2(n3466), .ZN(n3585) );
  NAND2_X1 U3742 ( .A1(n3714), .A2(n4592), .ZN(n3445) );
  OR2_X1 U3743 ( .A1(n3497), .A2(n3496), .ZN(n3599) );
  OR2_X1 U3744 ( .A1(n3481), .A2(n3480), .ZN(n3683) );
  AND4_X1 U3746 ( .A1(n3357), .A2(n3356), .A3(n3355), .A4(n3354), .ZN(n3423)
         );
  NAND2_X2 U3747 ( .A1(n3215), .A2(n3214), .ZN(n3427) );
  AND4_X1 U3748 ( .A1(n3340), .A2(n3339), .A3(n3338), .A4(n3337), .ZN(n3357)
         );
  AND4_X1 U3749 ( .A1(n3353), .A2(n3352), .A3(n3351), .A4(n3350), .ZN(n3354)
         );
  AND4_X1 U3750 ( .A1(n3344), .A2(n3343), .A3(n3342), .A4(n3341), .ZN(n3356)
         );
  AOI21_X1 U3751 ( .B1(n4076), .B2(INSTQUEUE_REG_1__1__SCAN_IN), .A(n3387), 
        .ZN(n3392) );
  AND4_X1 U3752 ( .A1(n3334), .A2(n3333), .A3(n3332), .A4(n3331), .ZN(n3335)
         );
  AND4_X1 U3753 ( .A1(n3308), .A2(n3307), .A3(n3306), .A4(n3305), .ZN(n3324)
         );
  AND2_X1 U3754 ( .A1(n3234), .A2(n3233), .ZN(n3232) );
  AND4_X1 U3755 ( .A1(n3312), .A2(n3311), .A3(n3310), .A4(n3309), .ZN(n3323)
         );
  AND2_X1 U3756 ( .A1(n3242), .A2(n3384), .ZN(n3241) );
  AND4_X1 U3757 ( .A1(n3348), .A2(n3347), .A3(n3346), .A4(n3345), .ZN(n3355)
         );
  AND4_X1 U3758 ( .A1(n3320), .A2(n3319), .A3(n3318), .A4(n3317), .ZN(n3321)
         );
  BUF_X2 U3759 ( .A(n3349), .Z(n4193) );
  BUF_X2 U3760 ( .A(n3475), .Z(n4185) );
  BUF_X2 U3761 ( .A(n4076), .Z(n4191) );
  NOR2_X1 U3762 ( .A1(n6476), .A2(n5236), .ZN(n6839) );
  INV_X2 U3763 ( .A(n6431), .ZN(n6419) );
  INV_X2 U3764 ( .A(n6216), .ZN(n3179) );
  OR2_X2 U3765 ( .A1(n6907), .A2(n6776), .ZN(n6476) );
  CLKBUF_X1 U3766 ( .A(n3213), .Z(n3180) );
  AND2_X1 U3767 ( .A1(n3397), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3290) );
  INV_X2 U3768 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n6773) );
  NAND2_X1 U3769 ( .A1(n3696), .A2(n3184), .ZN(n3181) );
  OR2_X1 U3770 ( .A1(n3183), .A2(n3199), .ZN(n3182) );
  INV_X1 U3771 ( .A(n3197), .ZN(n3183) );
  AND2_X1 U3772 ( .A1(n3695), .A2(n3197), .ZN(n3184) );
  OR2_X1 U3773 ( .A1(n5973), .A2(n5972), .ZN(n5975) );
  INV_X1 U3774 ( .A(n5256), .ZN(n3251) );
  AND2_X2 U3775 ( .A1(n4898), .A2(n3809), .ZN(n4897) );
  NAND2_X2 U3776 ( .A1(n3792), .A2(n3791), .ZN(n4898) );
  OAI22_X2 U3777 ( .A1(n5930), .A2(n6185), .B1(n6236), .B2(n5781), .ZN(n5782)
         );
  BUF_X2 U3778 ( .A(n5780), .Z(n5930) );
  NAND2_X1 U3779 ( .A1(n3615), .A2(n3614), .ZN(n3616) );
  AND2_X4 U3780 ( .A1(n3297), .A2(n3300), .ZN(n3457) );
  CLKBUF_X1 U3781 ( .A(n5512), .Z(n3185) );
  INV_X2 U3782 ( .A(n5512), .ZN(n3696) );
  OAI21_X2 U3783 ( .B1(n3693), .B2(n3282), .A(n3280), .ZN(n5512) );
  NAND2_X1 U3784 ( .A1(n3696), .A2(n3189), .ZN(n3186) );
  AND2_X2 U3785 ( .A1(n3186), .A2(n3187), .ZN(n5586) );
  OR2_X1 U3786 ( .A1(n3188), .A2(n3199), .ZN(n3187) );
  INV_X1 U3787 ( .A(n3190), .ZN(n3188) );
  AND2_X1 U3788 ( .A1(n6058), .A2(n3197), .ZN(n3190) );
  AND2_X2 U3789 ( .A1(n3192), .A2(n3193), .ZN(n5567) );
  AND2_X1 U3790 ( .A1(n3194), .A2(n5756), .ZN(n3193) );
  INV_X1 U3791 ( .A(n5589), .ZN(n3194) );
  NAND2_X1 U3792 ( .A1(n5797), .A2(n5799), .ZN(n3195) );
  OR2_X2 U3793 ( .A1(n3195), .A2(n3196), .ZN(n5605) );
  OR2_X1 U3794 ( .A1(n4178), .A2(n4766), .ZN(n3196) );
  OR2_X1 U3795 ( .A1(n3198), .A2(n3699), .ZN(n3197) );
  INV_X1 U3796 ( .A(n3701), .ZN(n3198) );
  AND2_X1 U3797 ( .A1(n3697), .A2(n3701), .ZN(n3199) );
  OR2_X2 U3798 ( .A1(n3200), .A2(n3201), .ZN(n3406) );
  NAND4_X1 U3799 ( .A1(n3296), .A2(n3295), .A3(n3294), .A4(n3293), .ZN(n3200)
         );
  NAND4_X1 U3800 ( .A1(n3304), .A2(n3303), .A3(n3302), .A4(n3301), .ZN(n3201)
         );
  INV_X1 U3801 ( .A(n3206), .ZN(n3203) );
  AND2_X1 U3802 ( .A1(n3456), .A2(n3406), .ZN(n3766) );
  AND2_X4 U3803 ( .A1(n3291), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4880)
         );
  OR2_X1 U3804 ( .A1(n3573), .A2(n3572), .ZN(n3574) );
  NOR2_X1 U3805 ( .A1(n3441), .A2(n3440), .ZN(n4586) );
  NAND2_X1 U3806 ( .A1(n3508), .A2(n3511), .ZN(n3535) );
  AOI21_X1 U3807 ( .B1(n3512), .B2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(n3517), 
        .ZN(n3533) );
  AND2_X4 U3808 ( .A1(n3297), .A2(n3298), .ZN(n3349) );
  AND2_X1 U3809 ( .A1(n3297), .A2(n5032), .ZN(n3212) );
  AND2_X1 U3810 ( .A1(n3300), .A2(n4887), .ZN(n3204) );
  AND2_X4 U3811 ( .A1(n3299), .A2(n4888), .ZN(n3394) );
  AND2_X2 U3812 ( .A1(n3416), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3512) );
  BUF_X4 U3813 ( .A(n3457), .Z(n3834) );
  AND4_X2 U3814 ( .A1(n3324), .A2(n3323), .A3(n3322), .A4(n3321), .ZN(n3378)
         );
  NAND2_X2 U3815 ( .A1(n3326), .A2(n3325), .ZN(n3410) );
  OAI21_X2 U3816 ( .B1(n4222), .B2(n4220), .A(n5633), .ZN(n4224) );
  NAND3_X2 U3817 ( .A1(n3272), .A2(n3273), .A3(n3274), .ZN(n4222) );
  NAND2_X2 U3818 ( .A1(n5476), .A2(n5477), .ZN(n3693) );
  XNOR2_X2 U3819 ( .A(n4245), .B(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5667)
         );
  OAI21_X2 U3820 ( .B1(n3689), .B2(n3278), .A(n3276), .ZN(n5458) );
  NAND4_X2 U3821 ( .A1(n3218), .A2(n3391), .A3(n3392), .A4(n3393), .ZN(n3429)
         );
  XNOR2_X2 U3822 ( .A(n3510), .B(n3455), .ZN(n4882) );
  BUF_X4 U3823 ( .A(n3386), .Z(n3209) );
  XNOR2_X2 U3824 ( .A(n3581), .B(n3580), .ZN(n3583) );
  NOR2_X4 U3825 ( .A1(n5505), .A2(n5506), .ZN(n5504) );
  XNOR2_X2 U3826 ( .A(n3583), .B(n3582), .ZN(n3768) );
  AND2_X1 U3827 ( .A1(n3297), .A2(n5032), .ZN(n3213) );
  INV_X1 U3828 ( .A(n4241), .ZN(n4244) );
  NAND2_X1 U3829 ( .A1(n3251), .A2(n3249), .ZN(n3255) );
  NOR2_X1 U3830 ( .A1(n3250), .A2(n5470), .ZN(n3249) );
  INV_X1 U3831 ( .A(n3252), .ZN(n3250) );
  OAI211_X1 U3832 ( .C1(n3660), .C2(n3269), .A(n3267), .B(n3265), .ZN(n3821)
         );
  NAND2_X1 U3833 ( .A1(n3671), .A2(n3268), .ZN(n3267) );
  INV_X1 U3834 ( .A(n3671), .ZN(n3269) );
  NAND2_X1 U3835 ( .A1(n3660), .A2(n3266), .ZN(n3265) );
  OR2_X1 U3836 ( .A1(n3660), .A2(n3286), .ZN(n3826) );
  NAND2_X1 U3837 ( .A1(n4897), .A2(n5271), .ZN(n5098) );
  AND2_X1 U3838 ( .A1(n5261), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3936) );
  INV_X1 U3839 ( .A(n4708), .ZN(n4723) );
  OR2_X1 U3840 ( .A1(n7008), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4044) );
  NAND2_X1 U3841 ( .A1(n5685), .A2(n3225), .ZN(n5671) );
  NOR2_X1 U3842 ( .A1(n5668), .A2(n3226), .ZN(n3225) );
  INV_X1 U3843 ( .A(n4726), .ZN(n3226) );
  NAND2_X1 U3844 ( .A1(n6891), .A2(n5889), .ZN(n5762) );
  AND2_X1 U3845 ( .A1(n3211), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n4242)
         );
  NOR2_X1 U3846 ( .A1(n3681), .A2(n3740), .ZN(n3682) );
  AND2_X1 U3847 ( .A1(n6891), .A2(n4610), .ZN(n6878) );
  OAI22_X1 U3848 ( .A1(n3738), .A2(n3737), .B1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n5603), .ZN(n3745) );
  XNOR2_X1 U3849 ( .A(n3739), .B(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3746)
         );
  NAND2_X1 U3850 ( .A1(n3398), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3239) );
  NAND2_X1 U3851 ( .A1(n4182), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3237) );
  NAND2_X1 U3852 ( .A1(n4076), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3233) );
  NAND2_X1 U3853 ( .A1(n3523), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3234)
         );
  INV_X1 U3854 ( .A(n3645), .ZN(n3646) );
  OAI22_X1 U3855 ( .A1(n4044), .A2(n6638), .B1(n3767), .B2(n6859), .ZN(n3451)
         );
  INV_X1 U3856 ( .A(n3444), .ZN(n3407) );
  NOR2_X2 U3857 ( .A1(n4585), .A2(n6894), .ZN(n4206) );
  INV_X1 U3858 ( .A(n3692), .ZN(n3281) );
  INV_X1 U3859 ( .A(n5515), .ZN(n3695) );
  INV_X1 U3860 ( .A(n5398), .ZN(n3278) );
  NAND2_X1 U3861 ( .A1(n5234), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3518) );
  AND2_X1 U3862 ( .A1(n3580), .A2(n3271), .ZN(n3270) );
  NAND2_X1 U3863 ( .A1(n3468), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3271) );
  NOR2_X1 U3864 ( .A1(n3580), .A2(n3247), .ZN(n3246) );
  NAND2_X1 U3865 ( .A1(n3535), .A2(n3534), .ZN(n5004) );
  INV_X1 U3866 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6859) );
  AND2_X1 U3867 ( .A1(n7002), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3767) );
  INV_X1 U3868 ( .A(n6254), .ZN(n4802) );
  NOR2_X2 U3869 ( .A1(n3444), .A2(n3429), .ZN(n6199) );
  OR2_X1 U3870 ( .A1(n4815), .A2(n4813), .ZN(n6447) );
  XNOR2_X1 U3871 ( .A(n4236), .B(n4329), .ZN(n5576) );
  NOR2_X1 U3872 ( .A1(n4235), .A2(n5769), .ZN(n4236) );
  INV_X1 U3873 ( .A(n3786), .ZN(n4213) );
  NAND2_X1 U3874 ( .A1(n4072), .A2(n3260), .ZN(n5807) );
  NOR2_X1 U3875 ( .A1(n3264), .A2(n3262), .ZN(n3260) );
  INV_X1 U3876 ( .A(n5617), .ZN(n3264) );
  NOR2_X1 U3877 ( .A1(n5545), .A2(n3257), .ZN(n3256) );
  INV_X1 U3878 ( .A(n5533), .ZN(n3257) );
  OR2_X2 U3879 ( .A1(n3255), .A2(n3254), .ZN(n5505) );
  INV_X1 U3880 ( .A(n5478), .ZN(n3254) );
  NOR2_X1 U3881 ( .A1(n5311), .A2(n3253), .ZN(n3252) );
  INV_X1 U3882 ( .A(n5399), .ZN(n3253) );
  XNOR2_X1 U3883 ( .A(n3211), .B(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n5398)
         );
  AND2_X1 U3884 ( .A1(n5257), .A2(n3827), .ZN(n3828) );
  INV_X1 U3885 ( .A(n5098), .ZN(n3829) );
  NOR4_X1 U3886 ( .A1(n4244), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .A3(n3211), 
        .A4(n4758), .ZN(n5608) );
  NOR3_X1 U3887 ( .A1(n6023), .A2(n6010), .A3(n4757), .ZN(n4221) );
  NAND4_X1 U3888 ( .A1(n4219), .A2(n4218), .A3(n5700), .A4(n5716), .ZN(n4220)
         );
  NAND2_X1 U3889 ( .A1(n5564), .A2(n4687), .ZN(n5864) );
  INV_X1 U3890 ( .A(n5880), .ZN(n4687) );
  OAI21_X1 U3891 ( .B1(n4222), .B2(n5980), .A(n3705), .ZN(n5973) );
  NOR2_X2 U3892 ( .A1(n6060), .A2(n6059), .ZN(n6061) );
  NAND2_X1 U3893 ( .A1(n4958), .A2(n4927), .ZN(n4941) );
  NAND2_X1 U3894 ( .A1(n4882), .A2(n6894), .ZN(n3248) );
  INV_X1 U3895 ( .A(n3710), .ZN(n4999) );
  BUF_X1 U3896 ( .A(n3378), .Z(n5261) );
  OR2_X1 U3897 ( .A1(n6075), .A2(n6901), .ZN(n4810) );
  OR2_X1 U3898 ( .A1(n5773), .A2(n6983), .ZN(n4805) );
  NAND2_X1 U3899 ( .A1(n5571), .A2(n4785), .ZN(n6236) );
  AND2_X1 U3900 ( .A1(n5576), .A2(n6903), .ZN(n6201) );
  OAI211_X1 U3901 ( .C1(n5671), .C2(n5658), .A(n5656), .B(n4779), .ZN(n4782)
         );
  OR2_X1 U3902 ( .A1(n6496), .A2(n4041), .ZN(n5640) );
  INV_X1 U3903 ( .A(n6498), .ZN(n6490) );
  AND2_X1 U3904 ( .A1(n5640), .A2(n4850), .ZN(n6498) );
  AND2_X1 U3905 ( .A1(n6878), .A2(n5889), .ZN(n6496) );
  OAI21_X1 U3906 ( .B1(n5681), .B2(n4758), .A(n5673), .ZN(n4233) );
  OR2_X1 U3907 ( .A1(n5687), .A2(n4754), .ZN(n4761) );
  NAND2_X1 U3908 ( .A1(n4581), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n4582) );
  OR2_X1 U3909 ( .A1(n4747), .A2(n4732), .ZN(n6512) );
  INV_X1 U3910 ( .A(n6512), .ZN(n6525) );
  INV_X1 U3911 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6864) );
  AOI22_X1 U3912 ( .A1(n3524), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3475), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3293) );
  AOI21_X1 U3913 ( .B1(n3349), .B2(INSTQUEUE_REG_6__5__SCAN_IN), .A(n3290), 
        .ZN(n3296) );
  AOI22_X1 U3914 ( .A1(n3523), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3388), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3303) );
  NOR2_X1 U3915 ( .A1(n3671), .A2(n3268), .ZN(n3266) );
  OR2_X1 U3916 ( .A1(n3657), .A2(n3656), .ZN(n3664) );
  OR2_X1 U3917 ( .A1(n3563), .A2(n3562), .ZN(n3636) );
  NAND3_X1 U3918 ( .A1(n3446), .A2(n3411), .A3(n3410), .ZN(n4733) );
  NAND2_X1 U3919 ( .A1(n3381), .A2(n3380), .ZN(n3382) );
  NAND2_X1 U3920 ( .A1(n3379), .A2(n3775), .ZN(n3381) );
  AND2_X1 U3921 ( .A1(n3386), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3387) );
  AOI22_X1 U3922 ( .A1(n3396), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3394), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3370) );
  AOI22_X1 U3923 ( .A1(n3395), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3834), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3376) );
  AOI21_X1 U3924 ( .B1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n6864), .A(n3748), 
        .ZN(n3754) );
  AOI21_X1 U3925 ( .B1(n3834), .B2(INSTQUEUE_REG_2__7__SCAN_IN), .A(n3362), 
        .ZN(n3365) );
  AND2_X1 U3926 ( .A1(n3212), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3362) );
  NAND2_X1 U3927 ( .A1(n3394), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3240) );
  NAND2_X1 U3928 ( .A1(n3204), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3238) );
  NAND2_X1 U3929 ( .A1(n3395), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3242) );
  NAND2_X1 U3930 ( .A1(n3399), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3243)
         );
  NAND2_X1 U3931 ( .A1(n3397), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3244) );
  NAND2_X1 U3932 ( .A1(n3349), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3235) );
  NAND2_X1 U3933 ( .A1(n4228), .A2(n3284), .ZN(n4241) );
  NAND2_X1 U3934 ( .A1(n3259), .A2(n3223), .ZN(n5860) );
  INV_X1 U3935 ( .A(n5568), .ZN(n3259) );
  INV_X1 U3936 ( .A(n5988), .ZN(n3258) );
  INV_X1 U3937 ( .A(n3719), .ZN(n3740) );
  NOR2_X1 U3938 ( .A1(n6021), .A2(n6058), .ZN(n3275) );
  NAND2_X1 U3939 ( .A1(n4745), .A2(n4744), .ZN(n6872) );
  NAND2_X1 U3940 ( .A1(n3423), .A2(n3427), .ZN(n4734) );
  AND2_X1 U3941 ( .A1(n3710), .A2(n4812), .ZN(n3719) );
  OR2_X1 U3942 ( .A1(n5259), .A2(n3683), .ZN(n3486) );
  OR2_X1 U3943 ( .A1(n3530), .A2(n3529), .ZN(n3566) );
  INV_X1 U3944 ( .A(n3451), .ZN(n3452) );
  OR2_X1 U3945 ( .A1(n3763), .A2(n3762), .ZN(n4585) );
  NAND2_X1 U3946 ( .A1(n4969), .A2(n6894), .ZN(n3550) );
  NAND2_X1 U3947 ( .A1(n3749), .A2(n3719), .ZN(n3758) );
  NAND2_X1 U3948 ( .A1(REIP_REG_14__SCAN_IN), .A2(n6122), .ZN(n5862) );
  NAND2_X1 U3949 ( .A1(n4723), .A2(n3206), .ZN(n4780) );
  AND2_X1 U3950 ( .A1(n5724), .A2(n5842), .ZN(n5844) );
  NAND2_X1 U3951 ( .A1(n6061), .A2(n6048), .ZN(n6050) );
  OR2_X1 U3952 ( .A1(n4159), .A2(n4158), .ZN(n4235) );
  OR2_X1 U3953 ( .A1(n4767), .A2(n4246), .ZN(n4247) );
  NAND2_X1 U3954 ( .A1(n4110), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n4141)
         );
  INV_X1 U3955 ( .A(n5641), .ZN(n3263) );
  OR2_X1 U3956 ( .A1(n4093), .A2(n5630), .ZN(n4094) );
  NOR2_X1 U3957 ( .A1(n4094), .A2(n4389), .ZN(n4110) );
  NOR2_X1 U3958 ( .A1(n4023), .A2(n4022), .ZN(n4024) );
  NOR2_X1 U3959 ( .A1(n3995), .A2(n5882), .ZN(n3996) );
  AND2_X1 U3960 ( .A1(n3968), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n3969)
         );
  NAND2_X1 U3961 ( .A1(n3969), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n3995)
         );
  NOR2_X1 U3962 ( .A1(n3955), .A2(n6105), .ZN(n3968) );
  NAND2_X1 U3963 ( .A1(n3950), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3955)
         );
  INV_X1 U3964 ( .A(n3923), .ZN(n3924) );
  NOR2_X1 U3965 ( .A1(n3924), .A2(n6118), .ZN(n3950) );
  NOR2_X1 U3966 ( .A1(n6128), .A2(n3900), .ZN(n3923) );
  NAND2_X1 U3967 ( .A1(n3871), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3872)
         );
  NOR2_X1 U3968 ( .A1(n3872), .A2(n6144), .ZN(n3895) );
  OR2_X1 U3969 ( .A1(n3844), .A2(n6170), .ZN(n3845) );
  NOR2_X1 U3970 ( .A1(n3845), .A2(n6164), .ZN(n3871) );
  NOR2_X1 U3971 ( .A1(n3822), .A2(n6192), .ZN(n3816) );
  NAND2_X1 U3972 ( .A1(PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n3816), .ZN(n3844)
         );
  NOR2_X1 U3973 ( .A1(n3818), .A2(n3283), .ZN(n3819) );
  INV_X1 U3974 ( .A(n3817), .ZN(n3818) );
  AOI21_X1 U3975 ( .B1(n3826), .B2(n3936), .A(n3825), .ZN(n5099) );
  NAND2_X1 U3976 ( .A1(n3811), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3822)
         );
  INV_X1 U3977 ( .A(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3794) );
  NOR2_X1 U3978 ( .A1(n3800), .A2(n3794), .ZN(n3811) );
  AND2_X1 U3979 ( .A1(n3808), .A2(n4907), .ZN(n3809) );
  NAND3_X1 U3980 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .A3(PHYADDRPOINTER_REG_3__SCAN_IN), 
        .ZN(n3800) );
  NOR2_X2 U3981 ( .A1(n5809), .A2(n4717), .ZN(n5813) );
  NAND2_X1 U3982 ( .A1(n5844), .A2(n5711), .ZN(n5710) );
  NAND2_X1 U3983 ( .A1(n5633), .A2(n3224), .ZN(n3274) );
  NAND2_X1 U3984 ( .A1(n3191), .A2(n3275), .ZN(n3272) );
  NAND2_X1 U3985 ( .A1(n5586), .A2(n5633), .ZN(n3273) );
  AND2_X1 U3986 ( .A1(n4686), .A2(n4685), .ZN(n5880) );
  NOR2_X1 U3987 ( .A1(n5248), .A2(n4749), .ZN(n5556) );
  NAND2_X1 U3988 ( .A1(n5526), .A2(n4670), .ZN(n5550) );
  AOI21_X1 U3989 ( .B1(n3281), .B2(n5494), .A(n3221), .ZN(n3280) );
  INV_X1 U3990 ( .A(n5494), .ZN(n3282) );
  XNOR2_X1 U3991 ( .A(n3211), .B(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n5494)
         );
  NOR2_X1 U3992 ( .A1(n5556), .A2(n6036), .ZN(n5495) );
  XNOR2_X1 U3993 ( .A(n3704), .B(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n5477)
         );
  INV_X1 U3994 ( .A(n3277), .ZN(n3276) );
  NAND2_X1 U3995 ( .A1(n5633), .A2(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n3279)
         );
  XNOR2_X1 U3996 ( .A(n3211), .B(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n5459)
         );
  AND2_X1 U3997 ( .A1(n4648), .A2(n4647), .ZN(n5124) );
  NAND2_X1 U3998 ( .A1(n4632), .A2(n4631), .ZN(n4957) );
  INV_X1 U3999 ( .A(n4919), .ZN(n4631) );
  NOR2_X2 U4000 ( .A1(n4957), .A2(n4956), .ZN(n4958) );
  NOR2_X1 U4001 ( .A1(n4728), .A2(n5267), .ZN(n4612) );
  AND2_X1 U4002 ( .A1(n4608), .A2(n4607), .ZN(n4747) );
  NAND2_X1 U4003 ( .A1(n3248), .A2(n3246), .ZN(n3506) );
  INV_X1 U4004 ( .A(n4966), .ZN(n5077) );
  OR2_X1 U4005 ( .A1(n6876), .A2(n3714), .ZN(n6851) );
  INV_X1 U4006 ( .A(n5337), .ZN(n5104) );
  AND2_X1 U4007 ( .A1(n6615), .A2(n5077), .ZN(n5145) );
  OR2_X1 U4008 ( .A1(n6676), .A2(n4966), .ZN(n5167) );
  INV_X1 U4009 ( .A(n3427), .ZN(n4988) );
  NAND3_X1 U4010 ( .A1(STATE2_REG_3__SCAN_IN), .A2(n6894), .A3(n4981), .ZN(
        n5322) );
  NAND2_X1 U4011 ( .A1(n6894), .A2(n4981), .ZN(n6646) );
  AOI21_X1 U4012 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n6769), .A(n6646), .ZN(
        n6780) );
  NOR2_X1 U4013 ( .A1(n4967), .A2(n5077), .ZN(n5187) );
  NAND2_X1 U4014 ( .A1(n7036), .A2(n4792), .ZN(n6254) );
  NAND2_X1 U4015 ( .A1(n5574), .A2(n5573), .ZN(n6264) );
  INV_X1 U4016 ( .A(n6236), .ZN(n6265) );
  AND2_X1 U4017 ( .A1(n5671), .A2(n5670), .ZN(n5900) );
  INV_X1 U4018 ( .A(n6324), .ZN(n6317) );
  NAND2_X1 U4019 ( .A1(n5216), .A2(n6317), .ZN(n6320) );
  INV_X1 U4020 ( .A(n6320), .ZN(n6323) );
  AND2_X1 U4021 ( .A1(n3446), .A2(n6317), .ZN(n6325) );
  NOR2_X2 U4022 ( .A1(n5267), .A2(n6358), .ZN(n6335) );
  NOR2_X2 U4023 ( .A1(n6358), .A2(n5268), .ZN(n6336) );
  INV_X1 U4024 ( .A(n6368), .ZN(n6360) );
  AOI21_X1 U4025 ( .B1(n5264), .B2(n5889), .A(n5263), .ZN(n5265) );
  NAND2_X1 U4026 ( .A1(n5266), .A2(n6365), .ZN(n6368) );
  INV_X1 U4027 ( .A(n6414), .ZN(n6436) );
  OR2_X1 U4028 ( .A1(n4815), .A2(n4814), .ZN(n6464) );
  INV_X1 U4029 ( .A(n6447), .ZN(n6450) );
  INV_X1 U4030 ( .A(n6464), .ZN(n6463) );
  NAND2_X1 U4031 ( .A1(n5504), .A2(n5533), .ZN(n5544) );
  NAND2_X1 U4032 ( .A1(n3251), .A2(n3252), .ZN(n5469) );
  INV_X1 U4033 ( .A(n6496), .ZN(n6484) );
  INV_X1 U4034 ( .A(n5900), .ZN(n5781) );
  NOR2_X1 U4035 ( .A1(n5607), .A2(n5608), .ZN(n4245) );
  INV_X1 U4036 ( .A(n5495), .ZN(n6045) );
  CLKBUF_X1 U4037 ( .A(n6469), .Z(n6470) );
  CLKBUF_X1 U4038 ( .A(n5096), .Z(n5097) );
  NAND2_X1 U4039 ( .A1(n5484), .A2(n6529), .ZN(n4944) );
  CLKBUF_X1 U4040 ( .A(n4895), .Z(n4896) );
  OR2_X1 U4041 ( .A1(n4747), .A2(n6851), .ZN(n5516) );
  INV_X1 U4042 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6769) );
  INV_X1 U4043 ( .A(n3774), .ZN(n6719) );
  NAND2_X1 U4044 ( .A1(STATE2_REG_3__SCAN_IN), .A2(n6891), .ZN(n5753) );
  INV_X1 U4045 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n6070) );
  INV_X1 U4046 ( .A(n5339), .ZN(n5413) );
  AND2_X1 U4047 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6614), .ZN(n6631)
         );
  INV_X1 U4048 ( .A(n6604), .ZN(n6630) );
  OR2_X1 U4049 ( .A1(n6676), .A2(n6675), .ZN(n6716) );
  AND2_X1 U4050 ( .A1(n6720), .A2(n3774), .ZN(n6821) );
  AND2_X1 U4051 ( .A1(n6720), .A2(n6719), .ZN(n6824) );
  INV_X1 U4052 ( .A(n6807), .ZN(n6748) );
  INV_X1 U4053 ( .A(n6819), .ZN(n6756) );
  NAND2_X1 U4054 ( .A1(n5187), .A2(n6719), .ZN(n5444) );
  NAND2_X1 U4055 ( .A1(n4805), .A2(n4804), .ZN(n4806) );
  NAND2_X1 U4056 ( .A1(n5645), .A2(n6496), .ZN(n4240) );
  NAND2_X1 U4057 ( .A1(n4765), .A2(n6496), .ZN(n4772) );
  AOI21_X1 U4058 ( .B1(n5931), .B2(n5989), .A(n4770), .ZN(n4771) );
  AOI21_X1 U4059 ( .B1(n5902), .B2(n6525), .A(n4762), .ZN(n4763) );
  NAND2_X1 U4060 ( .A1(n4765), .A2(n6528), .ZN(n4764) );
  NAND2_X1 U4061 ( .A1(n4761), .A2(n4760), .ZN(n4762) );
  NAND2_X1 U4063 ( .A1(n4072), .A2(n5641), .ZN(n5626) );
  NAND2_X1 U4064 ( .A1(n3191), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5585) );
  AND4_X1 U4065 ( .A1(n3372), .A2(n3371), .A3(n3370), .A4(n3369), .ZN(n3215)
         );
  OAI211_X1 U4066 ( .C1(n3483), .C2(n3518), .A(n3482), .B(n3486), .ZN(n3580)
         );
  XNOR2_X1 U4067 ( .A(n3642), .B(n4948), .ZN(n4938) );
  NAND2_X1 U4068 ( .A1(n3660), .A2(n3658), .ZN(n3679) );
  AND3_X1 U4069 ( .A1(n3245), .A2(n3244), .A3(n3243), .ZN(n3216) );
  AND2_X1 U4070 ( .A1(n5727), .A2(n5726), .ZN(n5724) );
  AND4_X1 U4071 ( .A1(n5234), .A2(n5261), .A3(n3446), .A4(n4611), .ZN(n3217)
         );
  AND4_X1 U4072 ( .A1(n3403), .A2(n3402), .A3(n3401), .A4(n3400), .ZN(n3218)
         );
  AND2_X1 U4073 ( .A1(n4072), .A2(n3261), .ZN(n3219) );
  BUF_X1 U4074 ( .A(n3423), .Z(n3426) );
  NAND2_X1 U4075 ( .A1(n3248), .A2(n3468), .ZN(n3582) );
  AND3_X1 U4076 ( .A1(n3434), .A2(n3433), .A3(n3432), .ZN(n3220) );
  NAND2_X1 U4077 ( .A1(n3641), .A2(n3640), .ZN(n3642) );
  NAND2_X1 U4078 ( .A1(n3675), .A2(n3674), .ZN(n3676) );
  NOR2_X1 U4079 ( .A1(n3211), .A2(n3694), .ZN(n3221) );
  OR2_X1 U4080 ( .A1(n5722), .A2(n5721), .ZN(n5621) );
  OR2_X1 U4081 ( .A1(n5259), .A2(n3483), .ZN(n3468) );
  INV_X1 U4082 ( .A(n3468), .ZN(n3247) );
  NOR2_X1 U4083 ( .A1(n5526), .A2(n5487), .ZN(n3222) );
  NOR2_X1 U4084 ( .A1(n5256), .A2(n5311), .ZN(n5310) );
  NOR2_X1 U4085 ( .A1(n5568), .A2(n5988), .ZN(n5874) );
  XNOR2_X1 U4086 ( .A(n3676), .B(n6521), .ZN(n6468) );
  NAND2_X1 U4087 ( .A1(n3689), .A2(n3688), .ZN(n5397) );
  NAND2_X1 U4088 ( .A1(n3693), .A2(n3692), .ZN(n5493) );
  NAND2_X1 U4089 ( .A1(n3829), .A2(n3828), .ZN(n5256) );
  AND2_X1 U4090 ( .A1(n4603), .A2(n3444), .ZN(n4783) );
  AND2_X1 U4091 ( .A1(n5876), .A2(n3258), .ZN(n3223) );
  INV_X1 U4092 ( .A(n3423), .ZN(n4593) );
  INV_X1 U4093 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n6894) );
  AND2_X1 U4094 ( .A1(n3755), .A2(n3664), .ZN(n3658) );
  INV_X1 U4095 ( .A(n3658), .ZN(n3268) );
  NOR2_X1 U4096 ( .A1(n6050), .A2(n5565), .ZN(n5564) );
  INV_X1 U4097 ( .A(n3262), .ZN(n3261) );
  OR2_X1 U4098 ( .A1(n5627), .A2(n3263), .ZN(n3262) );
  INV_X1 U4099 ( .A(n3781), .ZN(n4773) );
  INV_X1 U4100 ( .A(n4773), .ZN(n4179) );
  XNOR2_X1 U4101 ( .A(n3618), .B(n3571), .ZN(n4894) );
  NAND2_X1 U4102 ( .A1(n6773), .A2(n7000), .ZN(n6776) );
  NAND2_X1 U4103 ( .A1(n3703), .A2(n3702), .ZN(n3224) );
  INV_X1 U4104 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n6164) );
  INV_X1 U4105 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n6128) );
  OR2_X2 U4106 ( .A1(n5710), .A2(n5701), .ZN(n5809) );
  AND2_X2 U4107 ( .A1(n5486), .A2(n5485), .ZN(n5526) );
  NOR2_X2 U4108 ( .A1(n6159), .A2(n5460), .ZN(n5486) );
  NAND2_X1 U4109 ( .A1(n4657), .A2(n4656), .ZN(n6159) );
  NAND4_X4 U4110 ( .A1(n3216), .A2(n3241), .A3(n3176), .A4(n7037), .ZN(n3444)
         );
  NAND2_X1 U4113 ( .A1(n3396), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3236)
         );
  NAND2_X1 U4114 ( .A1(n3475), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3245) );
  INV_X1 U4115 ( .A(n3255), .ZN(n5468) );
  NAND2_X1 U4116 ( .A1(n5543), .A2(n5756), .ZN(n5588) );
  NAND2_X1 U4117 ( .A1(n5853), .A2(n5855), .ZN(n4039) );
  NOR2_X2 U4118 ( .A1(n5860), .A2(n5861), .ZN(n5853) );
  NOR2_X2 U4119 ( .A1(n5807), .A2(n5808), .ZN(n5797) );
  NAND2_X1 U4120 ( .A1(n4939), .A2(n4938), .ZN(n3644) );
  OAI21_X1 U4121 ( .B1(n4882), .B2(n3247), .A(n3270), .ZN(n3505) );
  NAND2_X1 U4122 ( .A1(n5458), .A2(n5459), .ZN(n3691) );
  NAND3_X1 U4123 ( .A1(n4224), .A2(n4226), .A3(n4223), .ZN(n4228) );
  NAND2_X1 U4124 ( .A1(n4224), .A2(n4223), .ZN(n5615) );
  CLKBUF_X1 U4125 ( .A(n5860), .Z(n5875) );
  AND2_X2 U4126 ( .A1(n3292), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3299)
         );
  NAND3_X1 U4127 ( .A1(n3454), .A2(n3453), .A3(n3452), .ZN(n3509) );
  NAND2_X1 U4128 ( .A1(n3421), .A2(n3425), .ZN(n4740) );
  XNOR2_X1 U4129 ( .A(n5611), .B(n5665), .ZN(n5654) );
  NAND2_X1 U4130 ( .A1(n5610), .A2(n5609), .ZN(n5611) );
  AND2_X1 U4131 ( .A1(PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n4213), .ZN(n3283)
         );
  OR2_X1 U4132 ( .A1(INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n5633), .ZN(n3284)
         );
  INV_X1 U4133 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n6118) );
  INV_X1 U4134 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n6170) );
  INV_X1 U4135 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n6144) );
  OR2_X1 U4136 ( .A1(n4780), .A2(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n3285)
         );
  NAND2_X1 U4137 ( .A1(n3268), .A2(n3659), .ZN(n3286) );
  INV_X1 U4138 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n6192) );
  OR2_X1 U4139 ( .A1(n4579), .A2(n4578), .ZN(n3287) );
  OR2_X1 U4140 ( .A1(n3451), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3288)
         );
  NAND2_X1 U4141 ( .A1(n4783), .A2(n3445), .ZN(n3448) );
  OR2_X1 U4142 ( .A1(n4154), .A2(n4153), .ZN(n4161) );
  OR2_X1 U4143 ( .A1(n3704), .A2(n3698), .ZN(n3699) );
  OR2_X1 U4144 ( .A1(n3633), .A2(n3632), .ZN(n3661) );
  NAND2_X1 U4145 ( .A1(n4588), .A2(n3456), .ZN(n3411) );
  INV_X1 U4146 ( .A(n3585), .ZN(n3483) );
  OR2_X1 U4147 ( .A1(n4162), .A2(n4161), .ZN(n4181) );
  AOI22_X1 U4148 ( .A1(n3212), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3399), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3375) );
  NAND2_X1 U4149 ( .A1(n4587), .A2(n3378), .ZN(n3380) );
  AOI22_X1 U4150 ( .A1(n3395), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3209), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3330) );
  NOR2_X1 U4151 ( .A1(n3747), .A2(n3746), .ZN(n3748) );
  AND2_X1 U4152 ( .A1(n4988), .A2(n3444), .ZN(n4708) );
  AND2_X1 U4153 ( .A1(n3390), .A2(n3389), .ZN(n3391) );
  INV_X1 U4154 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3739) );
  OR2_X1 U4155 ( .A1(n3548), .A2(n3547), .ZN(n3610) );
  INV_X1 U4156 ( .A(n6162), .ZN(n4656) );
  NAND2_X1 U4157 ( .A1(n4621), .A2(n4620), .ZN(n4625) );
  NAND2_X1 U4158 ( .A1(n3790), .A2(n3789), .ZN(n3791) );
  NOR2_X1 U4159 ( .A1(n3446), .A2(n6773), .ZN(n3777) );
  NOR2_X1 U4160 ( .A1(n4141), .A2(n5804), .ZN(n4142) );
  AND2_X1 U4161 ( .A1(n4886), .A2(n4742), .ZN(n4745) );
  NAND2_X1 U4162 ( .A1(n3538), .A2(n3537), .ZN(n6573) );
  OR2_X1 U4163 ( .A1(n6537), .A2(n4965), .ZN(n4967) );
  AOI221_X1 U4164 ( .B1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(n3754), .C1(
        n6070), .C2(n3754), .A(n3753), .ZN(n4599) );
  OR2_X1 U4165 ( .A1(n4073), .A2(n5639), .ZN(n4093) );
  INV_X1 U4166 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n6105) );
  NOR2_X1 U4167 ( .A1(n6240), .A2(n4793), .ZN(n6173) );
  AND2_X1 U4168 ( .A1(n3444), .A2(n7022), .ZN(n4787) );
  AND2_X1 U4169 ( .A1(n4661), .A2(n4660), .ZN(n5460) );
  NAND2_X1 U4170 ( .A1(n3446), .A2(n3775), .ZN(n5267) );
  NAND2_X1 U4172 ( .A1(n4024), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n4073)
         );
  NAND2_X1 U4173 ( .A1(n3895), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3900)
         );
  NAND2_X1 U4174 ( .A1(n3774), .A2(n3719), .ZN(n3602) );
  OR2_X1 U4175 ( .A1(n4747), .A2(n4745), .ZN(n5557) );
  OAI21_X1 U4176 ( .B1(n7027), .B2(n5765), .A(n5753), .ZN(n4981) );
  OR2_X1 U4177 ( .A1(n3798), .A2(n5051), .ZN(n5337) );
  OR2_X1 U4178 ( .A1(n3798), .A2(n5052), .ZN(n5076) );
  AND2_X1 U4179 ( .A1(n3210), .A2(n6259), .ZN(n6770) );
  INV_X1 U4180 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n5161) );
  NOR2_X1 U4181 ( .A1(n4967), .A2(n4966), .ZN(n6720) );
  INV_X1 U4182 ( .A(n6834), .ZN(n5422) );
  NAND2_X1 U4183 ( .A1(n3761), .A2(n3760), .ZN(n6891) );
  INV_X1 U4184 ( .A(n4783), .ZN(n6869) );
  INV_X1 U4185 ( .A(n7036), .ZN(n7022) );
  NOR2_X1 U4186 ( .A1(n5821), .A2(n4799), .ZN(n5801) );
  NOR2_X1 U4187 ( .A1(n5862), .A2(n4797), .ZN(n5847) );
  NOR2_X1 U4188 ( .A1(n6950), .A2(n6129), .ZN(n6122) );
  NOR2_X1 U4189 ( .A1(n4789), .A2(n6154), .ZN(n6150) );
  NAND3_X1 U4190 ( .A1(n4788), .A2(n4787), .A3(n4786), .ZN(n6240) );
  OR2_X1 U4191 ( .A1(n6201), .A2(n6200), .ZN(n6246) );
  INV_X1 U4192 ( .A(n5564), .ZN(n6034) );
  AND2_X1 U4193 ( .A1(n5896), .A2(n5895), .ZN(n6324) );
  AOI21_X1 U4194 ( .B1(n5764), .B2(n5763), .A(n6917), .ZN(n6414) );
  INV_X1 U4195 ( .A(n5764), .ZN(n6465) );
  OAI21_X1 U4196 ( .B1(n6490), .B2(n5786), .A(n4769), .ZN(n4770) );
  OAI21_X1 U4197 ( .B1(n6490), .B2(n5839), .A(n4045), .ZN(n4046) );
  NAND2_X1 U4198 ( .A1(n3996), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n4023)
         );
  INV_X1 U4199 ( .A(n5640), .ZN(n6491) );
  AND2_X1 U4200 ( .A1(n6045), .A2(n4756), .ZN(n6011) );
  NOR2_X1 U4201 ( .A1(n5483), .A2(n4944), .ZN(n6036) );
  NAND2_X1 U4202 ( .A1(n5516), .A2(n5557), .ZN(n5484) );
  INV_X1 U4203 ( .A(n6051), .ZN(n6528) );
  NOR2_X1 U4204 ( .A1(n5077), .A2(n6081), .ZN(n6678) );
  OR2_X1 U4205 ( .A1(n5108), .A2(n5107), .ZN(n5427) );
  INV_X1 U4206 ( .A(n5327), .ZN(n5411) );
  INV_X1 U4207 ( .A(n5326), .ZN(n6562) );
  NOR2_X1 U4208 ( .A1(n5076), .A2(n6719), .ZN(n6563) );
  AND2_X1 U4209 ( .A1(n5145), .A2(n3774), .ZN(n6600) );
  INV_X1 U4210 ( .A(n6672), .ZN(n6642) );
  AND2_X1 U4211 ( .A1(n4966), .A2(n3774), .ZN(n6674) );
  INV_X1 U4212 ( .A(n6708), .ZN(n6711) );
  INV_X1 U4213 ( .A(n6716), .ZN(n6763) );
  INV_X1 U4214 ( .A(n6783), .ZN(n6832) );
  AND2_X1 U4215 ( .A1(n3767), .A2(STATE2_REG_0__SCAN_IN), .ZN(n5889) );
  INV_X1 U4216 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n7002) );
  OR2_X1 U4217 ( .A1(n5762), .A2(n6869), .ZN(n4815) );
  INV_X1 U4218 ( .A(n6234), .ZN(n6266) );
  OR2_X1 U4219 ( .A1(n5576), .A2(n5575), .ZN(n6267) );
  NOR2_X1 U4220 ( .A1(n4044), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6216) );
  INV_X1 U4221 ( .A(n6264), .ZN(n6245) );
  INV_X1 U4222 ( .A(n6325), .ZN(n6321) );
  INV_X1 U4223 ( .A(n6140), .ZN(n6349) );
  NAND2_X1 U4224 ( .A1(n6447), .A2(n5265), .ZN(n6365) );
  INV_X1 U4225 ( .A(n6411), .ZN(n6434) );
  OR2_X1 U4226 ( .A1(n4815), .A2(n4812), .ZN(n5764) );
  AOI21_X1 U4227 ( .B1(n5947), .B2(n5989), .A(n4046), .ZN(n4047) );
  OR2_X1 U4228 ( .A1(n4747), .A2(n4615), .ZN(n6051) );
  INV_X1 U4229 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n5603) );
  NAND2_X1 U4230 ( .A1(n5104), .A2(n6719), .ZN(n5433) );
  AOI21_X1 U4231 ( .B1(n5058), .B2(n5057), .A(n6575), .ZN(n5331) );
  INV_X1 U4232 ( .A(n6541), .ZN(n6567) );
  INV_X1 U4233 ( .A(n6563), .ZN(n5441) );
  NAND2_X1 U4234 ( .A1(n5160), .A2(n3774), .ZN(n5416) );
  OR2_X1 U4235 ( .A1(n6676), .A2(n6568), .ZN(n6708) );
  NOR2_X1 U4236 ( .A1(n6728), .A2(n6727), .ZN(n6767) );
  INV_X1 U4237 ( .A(n6774), .ZN(n6830) );
  AND3_X1 U4238 ( .A1(n4975), .A2(n4974), .A3(n6725), .ZN(n5449) );
  INV_X1 U4239 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n7000) );
  INV_X1 U4240 ( .A(n6997), .ZN(n6993) );
  INV_X1 U4241 ( .A(STATE_REG_1__SCAN_IN), .ZN(n6918) );
  INV_X1 U4242 ( .A(n6979), .ZN(n6982) );
  NAND2_X1 U4243 ( .A1(n4772), .A2(n4771), .ZN(U2958) );
  NAND2_X1 U4244 ( .A1(n4764), .A2(n4763), .ZN(U2990) );
  INV_X1 U4245 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3289) );
  AND2_X2 U4246 ( .A1(n3739), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3298)
         );
  NOR2_X4 U4247 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4888) );
  NOR2_X4 U4248 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3300) );
  AND2_X4 U4249 ( .A1(n4888), .A2(n3300), .ZN(n3397) );
  INV_X1 U4250 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3291) );
  AND2_X2 U4251 ( .A1(n3298), .A2(n4880), .ZN(n3395) );
  AND2_X4 U4252 ( .A1(n4880), .A2(n3300), .ZN(n4076) );
  AOI22_X1 U4253 ( .A1(n3395), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n4076), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3295) );
  INV_X1 U4254 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3292) );
  AOI22_X1 U4256 ( .A1(n3212), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3396), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3294) );
  AND2_X2 U4257 ( .A1(n3298), .A2(n4888), .ZN(n3475) );
  AOI22_X1 U4258 ( .A1(n3457), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3399), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3304) );
  AND2_X4 U4259 ( .A1(n3298), .A2(n4887), .ZN(n3386) );
  AOI22_X1 U4260 ( .A1(n3386), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3394), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3302) );
  AND2_X2 U4261 ( .A1(n4880), .A2(n3299), .ZN(n3398) );
  AOI22_X1 U4262 ( .A1(n3398), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3469), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3301) );
  INV_X1 U4263 ( .A(n3406), .ZN(n3326) );
  NAND2_X1 U4264 ( .A1(n3524), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3308)
         );
  NAND2_X1 U4265 ( .A1(n3475), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3307) );
  NAND2_X1 U4266 ( .A1(n3388), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3306)
         );
  NAND2_X1 U4267 ( .A1(n3523), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3305)
         );
  NAND2_X1 U4268 ( .A1(n3212), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3312)
         );
  NAND2_X1 U4269 ( .A1(n3457), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3311) );
  NAND2_X1 U4270 ( .A1(n3399), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3310)
         );
  NAND2_X1 U4271 ( .A1(n3396), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3309)
         );
  NAND2_X1 U4272 ( .A1(n3395), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3316) );
  NAND2_X1 U4273 ( .A1(n4076), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3315) );
  NAND2_X1 U4274 ( .A1(n3386), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3314) );
  NAND2_X1 U4275 ( .A1(n3394), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3313) );
  NAND2_X1 U4276 ( .A1(n3398), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3320) );
  NAND2_X1 U4277 ( .A1(n3349), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3319) );
  NAND2_X1 U4278 ( .A1(n3469), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3318) );
  NAND2_X1 U4279 ( .A1(n3397), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3317) );
  AOI22_X1 U4280 ( .A1(n3457), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n3399), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3329) );
  AOI22_X1 U4281 ( .A1(n3524), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3388), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3328) );
  AOI22_X1 U4282 ( .A1(n3475), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n3523), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3327) );
  AOI22_X1 U4283 ( .A1(n3349), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3398), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3334) );
  AOI22_X1 U4284 ( .A1(n4076), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n3394), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3333) );
  AOI22_X1 U4285 ( .A1(n3213), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3396), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3332) );
  AOI22_X1 U4286 ( .A1(n3397), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n3204), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3331) );
  AND2_X4 U4287 ( .A1(n3336), .A2(n3335), .ZN(n3456) );
  NAND2_X2 U4288 ( .A1(n3410), .A2(n3456), .ZN(n4587) );
  NAND2_X1 U4289 ( .A1(n3395), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3340) );
  NAND2_X1 U4290 ( .A1(n4076), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3339) );
  NAND2_X1 U4291 ( .A1(n4182), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3338) );
  NAND2_X1 U4292 ( .A1(n3394), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3337) );
  NAND2_X1 U4293 ( .A1(n3213), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3344)
         );
  NAND2_X1 U4294 ( .A1(n3834), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3343) );
  NAND2_X1 U4295 ( .A1(n3399), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3342)
         );
  NAND2_X1 U4296 ( .A1(n3396), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3341)
         );
  NAND2_X1 U4297 ( .A1(n3524), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3348)
         );
  NAND2_X1 U4298 ( .A1(n3475), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3347) );
  NAND2_X1 U4299 ( .A1(n3388), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3346)
         );
  NAND2_X1 U4300 ( .A1(n3523), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3345)
         );
  NAND2_X1 U4301 ( .A1(n3398), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3353) );
  NAND2_X1 U4302 ( .A1(n3349), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3352) );
  NAND2_X1 U4303 ( .A1(n3204), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3351) );
  NAND2_X1 U4304 ( .A1(n3397), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3350) );
  NAND2_X1 U4305 ( .A1(n4587), .A2(n4593), .ZN(n3377) );
  AOI22_X1 U4306 ( .A1(n3398), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3397), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3361) );
  AOI22_X1 U4307 ( .A1(n3349), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3475), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3360) );
  AOI22_X1 U4308 ( .A1(n3524), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3388), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3359) );
  AOI22_X1 U4309 ( .A1(n4076), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3394), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3358) );
  NAND4_X1 U4310 ( .A1(n3361), .A2(n3360), .A3(n3359), .A4(n3358), .ZN(n3368)
         );
  AOI22_X1 U4311 ( .A1(n3395), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3208), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3366) );
  AOI22_X1 U4312 ( .A1(n3399), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3396), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3364) );
  AOI22_X1 U4313 ( .A1(n3204), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n3523), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3363) );
  NAND4_X1 U4314 ( .A1(n3366), .A2(n3365), .A3(n3364), .A4(n3363), .ZN(n3367)
         );
  AOI22_X1 U4315 ( .A1(n3524), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3398), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3372) );
  AOI22_X1 U4316 ( .A1(n4182), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4076), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3371) );
  AOI22_X1 U4317 ( .A1(n3397), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3469), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3369) );
  AOI22_X1 U4318 ( .A1(n3475), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3388), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3374) );
  AOI22_X1 U4319 ( .A1(n3349), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3523), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3373) );
  NAND2_X1 U4320 ( .A1(n3427), .A2(n3763), .ZN(n3431) );
  NAND2_X1 U4321 ( .A1(n3410), .A2(n3423), .ZN(n3379) );
  INV_X1 U4322 ( .A(n3378), .ZN(n3775) );
  AOI22_X1 U4323 ( .A1(n3213), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n3457), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3384) );
  AOI22_X1 U4324 ( .A1(n3524), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n3388), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3385) );
  AOI22_X1 U4325 ( .A1(n3349), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3469), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3393) );
  AOI22_X1 U4326 ( .A1(n3213), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3524), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3390) );
  AOI22_X1 U4327 ( .A1(n3475), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n3388), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3389) );
  AOI22_X1 U4328 ( .A1(n3395), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3394), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3403) );
  AOI22_X1 U4329 ( .A1(n3457), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n3396), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3402) );
  AOI22_X1 U4330 ( .A1(n3398), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3397), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3401) );
  AOI22_X1 U4331 ( .A1(n3399), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3523), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3400) );
  AND2_X1 U4332 ( .A1(STATE_REG_2__SCAN_IN), .A2(STATE_REG_1__SCAN_IN), .ZN(
        n6921) );
  INV_X1 U4333 ( .A(n6921), .ZN(n3405) );
  INV_X1 U4334 ( .A(STATE_REG_2__SCAN_IN), .ZN(n6073) );
  NAND2_X1 U4335 ( .A1(n6073), .A2(n6918), .ZN(n3404) );
  NAND2_X1 U4336 ( .A1(n3405), .A2(n3404), .ZN(n4592) );
  INV_X1 U4337 ( .A(n3445), .ZN(n3408) );
  NAND2_X1 U4338 ( .A1(n3763), .A2(n4611), .ZN(n3428) );
  NAND2_X1 U4339 ( .A1(n3407), .A2(n3429), .ZN(n3422) );
  OAI211_X1 U4340 ( .C1(n3408), .C2(n3710), .A(n3428), .B(n3422), .ZN(n3409)
         );
  INV_X1 U4341 ( .A(n3409), .ZN(n3412) );
  INV_X1 U4342 ( .A(n3763), .ZN(n4588) );
  AND2_X1 U4343 ( .A1(n3412), .A2(n3765), .ZN(n3415) );
  NOR2_X2 U4344 ( .A1(n4587), .A2(n5216), .ZN(n3443) );
  INV_X1 U4345 ( .A(n3443), .ZN(n3413) );
  AND2_X4 U4346 ( .A1(n3444), .A2(n3714), .ZN(n3567) );
  NAND2_X1 U4347 ( .A1(n3413), .A2(n3567), .ZN(n3414) );
  NAND2_X1 U4348 ( .A1(n3766), .A2(n7038), .ZN(n4883) );
  NAND3_X1 U4349 ( .A1(n3421), .A2(n3415), .A3(n3435), .ZN(n3416) );
  NAND2_X1 U4350 ( .A1(n3512), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3420) );
  INV_X1 U4351 ( .A(n3767), .ZN(n3417) );
  NAND2_X1 U4352 ( .A1(n7000), .A2(n7002), .ZN(n7008) );
  INV_X1 U4353 ( .A(n4044), .ZN(n3515) );
  MUX2_X1 U4354 ( .A(n3417), .B(n3515), .S(n6769), .Z(n3418) );
  INV_X1 U4355 ( .A(n3418), .ZN(n3419) );
  OAI22_X1 U4356 ( .A1(n3766), .A2(n3422), .B1(n5234), .B2(n3426), .ZN(n3424)
         );
  INV_X1 U4357 ( .A(n3424), .ZN(n3425) );
  INV_X1 U4358 ( .A(n4740), .ZN(n3439) );
  NAND2_X1 U4359 ( .A1(n3428), .A2(n3427), .ZN(n3430) );
  OAI21_X1 U4360 ( .B1(n4733), .B2(n3430), .A(n4812), .ZN(n3434) );
  NAND2_X1 U4361 ( .A1(n3431), .A2(n3567), .ZN(n3433) );
  OR2_X1 U4362 ( .A1(n7008), .A2(n6894), .ZN(n6902) );
  INV_X1 U4363 ( .A(n6902), .ZN(n3432) );
  NAND2_X1 U4364 ( .A1(n5021), .A2(n3220), .ZN(n3437) );
  INV_X1 U4365 ( .A(n3435), .ZN(n3436) );
  NOR2_X1 U4366 ( .A1(n3437), .A2(n3436), .ZN(n3438) );
  NAND2_X1 U4367 ( .A1(n3439), .A2(n3438), .ZN(n3484) );
  INV_X1 U4368 ( .A(n3766), .ZN(n3440) );
  NAND2_X1 U4369 ( .A1(n4586), .A2(n6199), .ZN(n4613) );
  NOR2_X1 U4370 ( .A1(n4734), .A2(n3710), .ZN(n3442) );
  INV_X1 U4371 ( .A(n4612), .ZN(n3447) );
  NAND3_X1 U4372 ( .A1(n4613), .A2(n3448), .A3(n3447), .ZN(n3449) );
  NAND2_X1 U4373 ( .A1(n3449), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3454) );
  INV_X1 U4374 ( .A(n3454), .ZN(n3450) );
  XNOR2_X1 U4375 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6638) );
  NAND2_X1 U4376 ( .A1(n3450), .A2(n3288), .ZN(n3508) );
  NAND2_X1 U4377 ( .A1(n3512), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3453) );
  NAND2_X1 U4378 ( .A1(n3508), .A2(n3509), .ZN(n3455) );
  AOI22_X1 U4379 ( .A1(n3395), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n4191), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3461) );
  AOI22_X1 U4380 ( .A1(n3180), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n3834), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3460) );
  AOI22_X1 U4381 ( .A1(n3209), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4194), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3459) );
  AOI22_X1 U4382 ( .A1(n4196), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4183), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3458) );
  NAND4_X1 U4383 ( .A1(n3461), .A2(n3460), .A3(n3459), .A4(n3458), .ZN(n3467)
         );
  AOI22_X1 U4384 ( .A1(n4193), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n4192), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3465) );
  AOI22_X1 U4385 ( .A1(n4185), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3207), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3464) );
  AOI22_X1 U4386 ( .A1(n4167), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n4186), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3463) );
  INV_X1 U4387 ( .A(n3474), .ZN(n3557) );
  AOI22_X1 U4388 ( .A1(n3524), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3474), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3462) );
  NAND4_X1 U4389 ( .A1(n3465), .A2(n3464), .A3(n3463), .A4(n3462), .ZN(n3466)
         );
  NAND2_X1 U4390 ( .A1(n3749), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3482) );
  AOI22_X1 U4391 ( .A1(n3178), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n3399), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3473) );
  AOI22_X1 U4392 ( .A1(INSTQUEUE_REG_7__7__SCAN_IN), .A2(n3349), .B1(n3398), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3472) );
  AOI22_X1 U4393 ( .A1(n4182), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n4194), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3471) );
  AOI22_X1 U4394 ( .A1(INSTQUEUE_REG_1__7__SCAN_IN), .A2(n4167), .B1(n4186), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3470) );
  NAND4_X1 U4395 ( .A1(n3473), .A2(n3472), .A3(n3471), .A4(n3470), .ZN(n3481)
         );
  AOI22_X1 U4396 ( .A1(n3395), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n4191), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3479) );
  AOI22_X1 U4397 ( .A1(n4195), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n4183), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3478) );
  AOI22_X1 U4398 ( .A1(n3524), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3474), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3477) );
  AOI22_X1 U4399 ( .A1(INSTQUEUE_REG_5__7__SCAN_IN), .A2(n4185), .B1(n3207), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3476) );
  NAND4_X1 U4400 ( .A1(n3479), .A2(n3478), .A3(n3477), .A4(n3476), .ZN(n3480)
         );
  XNOR2_X2 U4401 ( .A(n3485), .B(n3484), .ZN(n3776) );
  INV_X1 U4402 ( .A(n3486), .ZN(n3498) );
  INV_X1 U4403 ( .A(n3683), .ZN(n3487) );
  NOR2_X1 U4404 ( .A1(n5259), .A2(n3487), .ZN(n3680) );
  AOI22_X1 U4405 ( .A1(n4195), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n3399), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3491) );
  AOI22_X1 U4406 ( .A1(n3524), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n3398), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3490) );
  AOI22_X1 U4407 ( .A1(n3945), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n3394), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3489) );
  AOI22_X1 U4408 ( .A1(n4167), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n4186), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3488) );
  NAND4_X1 U4409 ( .A1(n3491), .A2(n3490), .A3(n3489), .A4(n3488), .ZN(n3497)
         );
  AOI22_X1 U4410 ( .A1(n3209), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n4191), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3495) );
  AOI22_X1 U4411 ( .A1(n3180), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n4183), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3494) );
  AOI22_X1 U4412 ( .A1(n4185), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n3474), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3493) );
  AOI22_X1 U4413 ( .A1(n4193), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3207), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3492) );
  NAND4_X1 U4414 ( .A1(n3495), .A2(n3494), .A3(n3493), .A4(n3492), .ZN(n3496)
         );
  INV_X1 U4415 ( .A(n3595), .ZN(n3499) );
  OAI21_X2 U4416 ( .B1(n3776), .B2(STATE2_REG_0__SCAN_IN), .A(n3499), .ZN(
        n3591) );
  NAND2_X1 U4417 ( .A1(n3749), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3504) );
  NAND2_X1 U4418 ( .A1(n3456), .A2(n3683), .ZN(n3500) );
  OAI211_X1 U4419 ( .C1(n3501), .C2(n3444), .A(n3500), .B(
        STATE2_REG_0__SCAN_IN), .ZN(n3502) );
  INV_X1 U4420 ( .A(n3502), .ZN(n3503) );
  NAND2_X1 U4421 ( .A1(n3504), .A2(n3503), .ZN(n3593) );
  AOI21_X2 U4422 ( .B1(n3591), .B2(n3593), .A(n3680), .ZN(n3579) );
  NAND2_X1 U4423 ( .A1(n3505), .A2(n3579), .ZN(n3507) );
  NAND2_X1 U4424 ( .A1(n3510), .A2(n3509), .ZN(n3511) );
  NOR2_X1 U4425 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n6859), .ZN(n5281)
         );
  NAND2_X1 U4426 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5281), .ZN(n6677) );
  NAND2_X1 U4427 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3513) );
  NAND2_X1 U4428 ( .A1(n3513), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3514) );
  NAND2_X1 U4429 ( .A1(n6677), .A2(n3514), .ZN(n4977) );
  NAND2_X1 U4430 ( .A1(n4977), .A2(n3515), .ZN(n3516) );
  OAI21_X1 U4431 ( .B1(n3767), .B2(n5161), .A(n3516), .ZN(n3517) );
  XNOR2_X1 U4432 ( .A(n3535), .B(n3533), .ZN(n4968) );
  NAND2_X1 U4433 ( .A1(n4968), .A2(n6894), .ZN(n3532) );
  AOI22_X1 U4434 ( .A1(n3945), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n4191), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3522) );
  AOI22_X1 U4435 ( .A1(n3180), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n3834), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3521) );
  AOI22_X1 U4436 ( .A1(n3209), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3394), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3520) );
  AOI22_X1 U4437 ( .A1(n4196), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4183), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3519) );
  NAND4_X1 U4438 ( .A1(n3522), .A2(n3521), .A3(n3520), .A4(n3519), .ZN(n3530)
         );
  AOI22_X1 U4439 ( .A1(n3349), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n4192), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3528) );
  AOI22_X1 U4440 ( .A1(n4185), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3207), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3527) );
  AOI22_X1 U4441 ( .A1(n4167), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n4186), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3526) );
  AOI22_X1 U4442 ( .A1(n4184), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3474), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3525) );
  NAND4_X1 U4443 ( .A1(n3528), .A2(n3527), .A3(n3526), .A4(n3525), .ZN(n3529)
         );
  AOI22_X1 U4444 ( .A1(n3755), .A2(n3566), .B1(n3749), .B2(
        INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3531) );
  NAND2_X2 U4445 ( .A1(n3573), .A2(n3572), .ZN(n3609) );
  INV_X1 U4446 ( .A(n3609), .ZN(n3551) );
  INV_X1 U4447 ( .A(n3533), .ZN(n3534) );
  NAND2_X1 U4448 ( .A1(n3512), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3538) );
  NOR3_X1 U4449 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6859), .A3(n5161), 
        .ZN(n6614) );
  NAND3_X1 U4450 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), 
        .ZN(n5192) );
  INV_X1 U4451 ( .A(n5192), .ZN(n5188) );
  AND2_X1 U4452 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5188), .ZN(n6834)
         );
  OAI21_X1 U4453 ( .B1(n6631), .B2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(n5422), 
        .ZN(n6637) );
  OAI22_X1 U4454 ( .A1(n6637), .A2(n4044), .B1(n3767), .B2(n6864), .ZN(n3536)
         );
  INV_X1 U4455 ( .A(n3536), .ZN(n3537) );
  AOI22_X1 U4456 ( .A1(n4076), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n4194), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3542) );
  AOI22_X1 U4457 ( .A1(n4184), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4185), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3541) );
  AOI22_X1 U4458 ( .A1(n4196), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4183), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3540) );
  AOI22_X1 U4459 ( .A1(n4186), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3207), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3539) );
  NAND4_X1 U4460 ( .A1(n3542), .A2(n3541), .A3(n3540), .A4(n3539), .ZN(n3548)
         );
  AOI22_X1 U4461 ( .A1(n3945), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n4182), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3546) );
  AOI22_X1 U4462 ( .A1(n3178), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n3834), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3545) );
  AOI22_X1 U4463 ( .A1(n4193), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3474), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3544) );
  AOI22_X1 U4464 ( .A1(n4192), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3397), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3543) );
  NAND4_X1 U4465 ( .A1(n3546), .A2(n3545), .A3(n3544), .A4(n3543), .ZN(n3547)
         );
  AOI22_X1 U4466 ( .A1(n3755), .A2(n3610), .B1(n3749), .B2(
        INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3549) );
  NAND2_X1 U4467 ( .A1(n3551), .A2(n5042), .ZN(n3621) );
  AOI22_X1 U4468 ( .A1(n3945), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n4191), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3556) );
  AOI22_X1 U4469 ( .A1(n3178), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n3834), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3555) );
  INV_X1 U4470 ( .A(n3394), .ZN(n3552) );
  INV_X2 U4471 ( .A(n3552), .ZN(n4194) );
  AOI22_X1 U4472 ( .A1(n3209), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n4194), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3554) );
  AOI22_X1 U4473 ( .A1(n4196), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4183), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3553) );
  NAND4_X1 U4474 ( .A1(n3556), .A2(n3555), .A3(n3554), .A4(n3553), .ZN(n3563)
         );
  AOI22_X1 U4475 ( .A1(n4193), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n4192), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3561) );
  AOI22_X1 U4476 ( .A1(n4185), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3207), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3560) );
  AOI22_X1 U4477 ( .A1(n4167), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n4186), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3559) );
  AOI22_X1 U4478 ( .A1(n4184), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3474), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3558) );
  NAND4_X1 U4479 ( .A1(n3561), .A2(n3560), .A3(n3559), .A4(n3558), .ZN(n3562)
         );
  NAND2_X1 U4480 ( .A1(n3755), .A2(n3636), .ZN(n3565) );
  NAND2_X1 U4481 ( .A1(n3749), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3564) );
  NAND2_X1 U4482 ( .A1(n3565), .A2(n3564), .ZN(n3622) );
  XNOR2_X1 U4483 ( .A(n3621), .B(n3622), .ZN(n3793) );
  NAND2_X1 U4484 ( .A1(n3793), .A2(n3719), .ZN(n3570) );
  NAND2_X1 U4485 ( .A1(n3585), .A2(n3599), .ZN(n3584) );
  INV_X1 U4486 ( .A(n3566), .ZN(n3575) );
  NAND2_X1 U4487 ( .A1(n3584), .A2(n3575), .ZN(n3612) );
  NAND2_X1 U4488 ( .A1(n3612), .A2(n3610), .ZN(n3638) );
  XNOR2_X1 U4489 ( .A(n3638), .B(n3636), .ZN(n3568) );
  NAND2_X1 U4490 ( .A1(n3568), .A2(n3567), .ZN(n3569) );
  NAND2_X1 U4491 ( .A1(n3570), .A2(n3569), .ZN(n3618) );
  INV_X1 U4492 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n3571) );
  NAND2_X2 U4493 ( .A1(n3574), .A2(n3609), .ZN(n6537) );
  OAI21_X1 U4494 ( .B1(n3575), .B2(n3584), .A(n3612), .ZN(n3577) );
  NAND2_X1 U4495 ( .A1(n5234), .A2(n3427), .ZN(n3598) );
  INV_X1 U4496 ( .A(n3598), .ZN(n3576) );
  AOI21_X1 U4497 ( .B1(n3567), .B2(n3577), .A(n3576), .ZN(n3578) );
  OAI21_X1 U4498 ( .B1(n6537), .B2(n3740), .A(n3578), .ZN(n3605) );
  NAND2_X1 U4499 ( .A1(n3605), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n4912)
         );
  INV_X1 U4500 ( .A(n3579), .ZN(n3581) );
  NAND2_X1 U4501 ( .A1(n3768), .A2(n3719), .ZN(n3590) );
  OAI21_X1 U4502 ( .B1(n3599), .B2(n3585), .A(n3584), .ZN(n3587) );
  INV_X1 U4503 ( .A(n3567), .ZN(n7026) );
  INV_X1 U4504 ( .A(n4734), .ZN(n3586) );
  OAI211_X1 U4505 ( .C1(n3587), .C2(n7026), .A(n3586), .B(n3710), .ZN(n3588)
         );
  INV_X1 U4506 ( .A(n3588), .ZN(n3589) );
  NAND2_X1 U4507 ( .A1(n3590), .A2(n3589), .ZN(n6493) );
  INV_X1 U4508 ( .A(n3591), .ZN(n3592) );
  NAND2_X1 U4509 ( .A1(n3592), .A2(n3593), .ZN(n3597) );
  INV_X1 U4510 ( .A(n3593), .ZN(n3594) );
  NAND2_X1 U4511 ( .A1(n3595), .A2(n3594), .ZN(n3596) );
  OAI21_X1 U4512 ( .B1(n7026), .B2(n3599), .A(n3598), .ZN(n3600) );
  INV_X1 U4513 ( .A(n3600), .ZN(n3601) );
  NAND2_X1 U4514 ( .A1(n3602), .A2(n3601), .ZN(n4849) );
  NAND2_X1 U4515 ( .A1(n4849), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n3603)
         );
  XNOR2_X1 U4516 ( .A(n3603), .B(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n6492)
         );
  NAND2_X1 U4517 ( .A1(n6493), .A2(n6492), .ZN(n6495) );
  INV_X1 U4518 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n6531) );
  OR2_X1 U4519 ( .A1(n3603), .A2(n6531), .ZN(n3604) );
  NAND2_X1 U4520 ( .A1(n4915), .A2(n4912), .ZN(n3608) );
  INV_X1 U4521 ( .A(n3605), .ZN(n3607) );
  INV_X1 U4522 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3606) );
  NAND2_X1 U4523 ( .A1(n3607), .A2(n3606), .ZN(n4913) );
  NAND2_X1 U4524 ( .A1(n3608), .A2(n4913), .ZN(n4905) );
  XNOR2_X2 U4525 ( .A(n3609), .B(n5042), .ZN(n3798) );
  NAND2_X1 U4526 ( .A1(n3798), .A2(n3719), .ZN(n3615) );
  INV_X1 U4527 ( .A(n3610), .ZN(n3611) );
  XNOR2_X1 U4528 ( .A(n3612), .B(n3611), .ZN(n3613) );
  NAND2_X1 U4529 ( .A1(n3613), .A2(n3567), .ZN(n3614) );
  NAND2_X1 U4530 ( .A1(n3616), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n3617)
         );
  OAI21_X2 U4531 ( .B1(n4905), .B2(n4906), .A(n3617), .ZN(n4895) );
  NAND2_X1 U4532 ( .A1(n4894), .A2(n4895), .ZN(n3620) );
  NAND2_X1 U4533 ( .A1(n3618), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n3619)
         );
  NAND2_X1 U4534 ( .A1(n3620), .A2(n3619), .ZN(n4939) );
  INV_X1 U4535 ( .A(n3621), .ZN(n3623) );
  NAND2_X1 U4536 ( .A1(n3623), .A2(n3622), .ZN(n3647) );
  AOI22_X1 U4537 ( .A1(n3945), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n4191), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3627) );
  AOI22_X1 U4538 ( .A1(n3178), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n3834), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3626) );
  AOI22_X1 U4539 ( .A1(n4182), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4194), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3625) );
  AOI22_X1 U4540 ( .A1(n4196), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4183), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3624) );
  NAND4_X1 U4541 ( .A1(n3627), .A2(n3626), .A3(n3625), .A4(n3624), .ZN(n3633)
         );
  AOI22_X1 U4542 ( .A1(n4193), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n4192), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3631) );
  AOI22_X1 U4543 ( .A1(n4185), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3207), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3630) );
  AOI22_X1 U4544 ( .A1(n4167), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n4186), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3629) );
  AOI22_X1 U4545 ( .A1(n4184), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3474), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3628) );
  NAND4_X1 U4546 ( .A1(n3631), .A2(n3630), .A3(n3629), .A4(n3628), .ZN(n3632)
         );
  NAND2_X1 U4547 ( .A1(n3755), .A2(n3661), .ZN(n3635) );
  NAND2_X1 U4548 ( .A1(n3749), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3634) );
  NAND2_X1 U4549 ( .A1(n3635), .A2(n3634), .ZN(n3645) );
  XNOR2_X1 U4550 ( .A(n3647), .B(n3645), .ZN(n3810) );
  NAND2_X1 U4551 ( .A1(n3810), .A2(n3719), .ZN(n3641) );
  INV_X1 U4552 ( .A(n3636), .ZN(n3637) );
  OR2_X1 U4553 ( .A1(n3638), .A2(n3637), .ZN(n3663) );
  XNOR2_X1 U4554 ( .A(n3663), .B(n3661), .ZN(n3639) );
  NAND2_X1 U4555 ( .A1(n3639), .A2(n3567), .ZN(n3640) );
  INV_X1 U4556 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4948) );
  NAND2_X1 U4557 ( .A1(n3642), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n3643)
         );
  NAND2_X1 U4558 ( .A1(n3644), .A2(n3643), .ZN(n5096) );
  AOI22_X1 U4559 ( .A1(n3945), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4191), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3651) );
  AOI22_X1 U4560 ( .A1(n3180), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n3834), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3650) );
  AOI22_X1 U4561 ( .A1(n3209), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4194), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3649) );
  AOI22_X1 U4562 ( .A1(n4196), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4183), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3648) );
  NAND4_X1 U4563 ( .A1(n3651), .A2(n3650), .A3(n3649), .A4(n3648), .ZN(n3657)
         );
  AOI22_X1 U4564 ( .A1(n4193), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n4192), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3655) );
  AOI22_X1 U4565 ( .A1(n4185), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3207), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3654) );
  AOI22_X1 U4566 ( .A1(n4167), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n4186), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3653) );
  AOI22_X1 U4567 ( .A1(n4184), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3474), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3652) );
  NAND4_X1 U4568 ( .A1(n3655), .A2(n3654), .A3(n3653), .A4(n3652), .ZN(n3656)
         );
  NAND2_X1 U4569 ( .A1(n3749), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3659) );
  NAND3_X1 U4570 ( .A1(n3679), .A2(n3719), .A3(n3826), .ZN(n3667) );
  INV_X1 U4571 ( .A(n3661), .ZN(n3662) );
  NOR2_X1 U4572 ( .A1(n3663), .A2(n3662), .ZN(n3665) );
  NAND2_X1 U4573 ( .A1(n3665), .A2(n3664), .ZN(n3685) );
  OAI211_X1 U4574 ( .C1(n3665), .C2(n3664), .A(n3685), .B(n3567), .ZN(n3666)
         );
  NAND2_X1 U4575 ( .A1(n3667), .A2(n3666), .ZN(n3668) );
  INV_X1 U4576 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n4644) );
  XNOR2_X1 U4577 ( .A(n3668), .B(n4644), .ZN(n5095) );
  NAND2_X1 U4578 ( .A1(n5096), .A2(n5095), .ZN(n3670) );
  NAND2_X1 U4579 ( .A1(n3668), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n3669)
         );
  NAND2_X1 U4580 ( .A1(n3670), .A2(n3669), .ZN(n6469) );
  AOI22_X1 U4581 ( .A1(n3755), .A2(n3683), .B1(n3749), .B2(
        INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3671) );
  INV_X1 U4582 ( .A(n3821), .ZN(n3672) );
  NAND2_X1 U4583 ( .A1(n3672), .A2(n3719), .ZN(n3675) );
  XNOR2_X1 U4584 ( .A(n3685), .B(n3683), .ZN(n3673) );
  NAND2_X1 U4585 ( .A1(n3673), .A2(n3567), .ZN(n3674) );
  INV_X1 U4586 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n6521) );
  NAND2_X1 U4587 ( .A1(n6469), .A2(n6468), .ZN(n3678) );
  NAND2_X1 U4588 ( .A1(n3676), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n3677)
         );
  INV_X1 U4589 ( .A(n3680), .ZN(n3681) );
  NAND2_X1 U4590 ( .A1(n3567), .A2(n3683), .ZN(n3684) );
  OR2_X1 U4591 ( .A1(n3685), .A2(n3684), .ZN(n3686) );
  NAND2_X1 U4592 ( .A1(n3704), .A2(n3686), .ZN(n3687) );
  INV_X1 U4593 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n5250) );
  NAND2_X1 U4594 ( .A1(n3687), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n3688)
         );
  INV_X1 U4595 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n5463) );
  INV_X1 U4596 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n5464) );
  OR2_X1 U4597 ( .A1(n3211), .A2(n5464), .ZN(n3690) );
  NAND2_X1 U4598 ( .A1(n3691), .A2(n3690), .ZN(n5476) );
  INV_X1 U4599 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n5496) );
  OR2_X1 U4600 ( .A1(n3211), .A2(n5496), .ZN(n3692) );
  INV_X1 U4601 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n3694) );
  INV_X1 U4602 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n4748) );
  XNOR2_X1 U4603 ( .A(n3704), .B(n4748), .ZN(n5515) );
  NAND2_X1 U4604 ( .A1(n3704), .A2(n4748), .ZN(n3697) );
  NAND2_X1 U4605 ( .A1(n5513), .A2(n3697), .ZN(n5539) );
  NOR2_X1 U4606 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n3698) );
  AND2_X1 U4607 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n6056) );
  INV_X1 U4608 ( .A(n6056), .ZN(n3700) );
  NAND2_X1 U4609 ( .A1(n3211), .A2(n3700), .ZN(n3701) );
  INV_X1 U4610 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n6058) );
  INV_X1 U4611 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n3703) );
  INV_X1 U4612 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n3702) );
  NAND2_X1 U4613 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n6021) );
  INV_X1 U4614 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n6031) );
  XNOR2_X1 U4615 ( .A(n3211), .B(n6031), .ZN(n5980) );
  NAND2_X1 U4616 ( .A1(n3704), .A2(n6031), .ZN(n3705) );
  INV_X1 U4617 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n6017) );
  XNOR2_X1 U4618 ( .A(n3704), .B(n6017), .ZN(n5972) );
  OR2_X1 U4619 ( .A1(n3704), .A2(n6017), .ZN(n3706) );
  NAND2_X1 U4620 ( .A1(n5975), .A2(n3706), .ZN(n5722) );
  INV_X1 U4621 ( .A(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5730) );
  XNOR2_X1 U4622 ( .A(n3211), .B(n5730), .ZN(n5721) );
  NAND2_X1 U4623 ( .A1(n3211), .A2(n5730), .ZN(n3707) );
  NAND2_X1 U4624 ( .A1(n5621), .A2(n3707), .ZN(n5624) );
  NOR2_X1 U4625 ( .A1(n3211), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5622)
         );
  AND2_X1 U4626 ( .A1(n3704), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n3708)
         );
  NOR2_X1 U4627 ( .A1(n5622), .A2(n3708), .ZN(n3709) );
  XNOR2_X1 U4628 ( .A(n5624), .B(n3709), .ZN(n6005) );
  NAND2_X1 U4629 ( .A1(n3755), .A2(n4812), .ZN(n3711) );
  NAND2_X1 U4630 ( .A1(n3711), .A2(n3710), .ZN(n3718) );
  INV_X1 U4631 ( .A(n3718), .ZN(n3723) );
  XNOR2_X1 U4632 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3728) );
  NAND2_X1 U4633 ( .A1(n6769), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3727) );
  XNOR2_X1 U4634 ( .A(n3728), .B(n3727), .ZN(n4596) );
  NAND2_X1 U4635 ( .A1(n4596), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3721) );
  INV_X1 U4636 ( .A(n3755), .ZN(n3732) );
  OAI21_X1 U4637 ( .B1(n6769), .B2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(n3727), 
        .ZN(n3713) );
  NOR2_X1 U4638 ( .A1(n3732), .A2(n3713), .ZN(n3717) );
  OAI21_X1 U4639 ( .B1(n3766), .B2(n3713), .A(n3712), .ZN(n3716) );
  NAND2_X1 U4640 ( .A1(n4999), .A2(n3444), .ZN(n3715) );
  NAND2_X1 U4641 ( .A1(n3715), .A2(n3714), .ZN(n3733) );
  NAND2_X1 U4642 ( .A1(n3716), .A2(n3733), .ZN(n3722) );
  OAI211_X1 U4643 ( .C1(n3718), .C2(n4596), .A(n3717), .B(n3722), .ZN(n3720)
         );
  OAI211_X1 U4644 ( .C1(n3723), .C2(n3721), .A(n3720), .B(n3758), .ZN(n3726)
         );
  INV_X1 U4645 ( .A(n3722), .ZN(n3724) );
  NAND3_X1 U4646 ( .A1(n3724), .A2(n4596), .A3(n3723), .ZN(n3725) );
  NAND2_X1 U4647 ( .A1(n3726), .A2(n3725), .ZN(n3742) );
  INV_X1 U4648 ( .A(n3727), .ZN(n3729) );
  NAND2_X1 U4649 ( .A1(n3729), .A2(n3728), .ZN(n3731) );
  NAND2_X1 U4650 ( .A1(n6859), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3730) );
  NAND2_X1 U4651 ( .A1(n3731), .A2(n3730), .ZN(n3736) );
  XNOR2_X1 U4652 ( .A(n5603), .B(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3737)
         );
  XNOR2_X1 U4653 ( .A(n3736), .B(n3737), .ZN(n4595) );
  INV_X1 U4654 ( .A(n4595), .ZN(n3735) );
  AOI211_X1 U4655 ( .C1(n3742), .C2(n3733), .A(n3732), .B(n3735), .ZN(n3744)
         );
  INV_X1 U4656 ( .A(n3733), .ZN(n3734) );
  AOI21_X1 U4657 ( .B1(n3749), .B2(n3735), .A(n3734), .ZN(n3741) );
  INV_X1 U4658 ( .A(n3736), .ZN(n3738) );
  XNOR2_X1 U4659 ( .A(n3745), .B(n3746), .ZN(n4594) );
  OAI22_X1 U4660 ( .A1(n3742), .A2(n3741), .B1(n4594), .B2(n3740), .ZN(n3743)
         );
  NOR2_X1 U4661 ( .A1(n3744), .A2(n3743), .ZN(n3751) );
  INV_X1 U4662 ( .A(n3745), .ZN(n3747) );
  NAND3_X1 U4663 ( .A1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n3754), .A3(n6070), .ZN(n4597) );
  AOI21_X1 U4664 ( .B1(n4594), .B2(n4597), .A(n3749), .ZN(n3750) );
  OAI22_X1 U4665 ( .A1(n3751), .A2(n3750), .B1(n3758), .B2(n4597), .ZN(n3752)
         );
  AOI21_X1 U4666 ( .B1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n6894), .A(n3752), 
        .ZN(n3757) );
  INV_X1 U4667 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n6536) );
  NOR2_X1 U4668 ( .A1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n6536), .ZN(n3753)
         );
  NAND2_X1 U4669 ( .A1(n4599), .A2(n3755), .ZN(n3756) );
  NAND2_X1 U4670 ( .A1(n3757), .A2(n3756), .ZN(n3761) );
  INV_X1 U4671 ( .A(n3758), .ZN(n3759) );
  NAND2_X1 U4672 ( .A1(n4599), .A2(n3759), .ZN(n3760) );
  NAND2_X1 U4673 ( .A1(n3446), .A2(n4611), .ZN(n3762) );
  NAND2_X1 U4674 ( .A1(n4585), .A2(n5234), .ZN(n3764) );
  AND2_X1 U4675 ( .A1(n3765), .A2(n3764), .ZN(n4609) );
  AND2_X1 U4676 ( .A1(n4609), .A2(n3766), .ZN(n4610) );
  NAND2_X1 U4677 ( .A1(n4966), .A2(n3936), .ZN(n3773) );
  NOR2_X1 U4678 ( .A1(n5267), .A2(n6773), .ZN(n3805) );
  NAND2_X1 U4679 ( .A1(n4214), .A2(EAX_REG_1__SCAN_IN), .ZN(n3770) );
  NAND2_X1 U4680 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n6773), .ZN(n3769)
         );
  NAND2_X1 U4681 ( .A1(n3770), .A2(n3769), .ZN(n3771) );
  AOI21_X1 U4682 ( .B1(n3805), .B2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(n3771), 
        .ZN(n3772) );
  NAND2_X1 U4683 ( .A1(n3773), .A2(n3772), .ZN(n6249) );
  OAI21_X1 U4684 ( .B1(n3774), .B2(n3775), .A(STATE2_REG_2__SCAN_IN), .ZN(
        n4852) );
  INV_X1 U4685 ( .A(n3776), .ZN(n6681) );
  INV_X1 U4686 ( .A(n3936), .ZN(n3820) );
  OR2_X1 U4687 ( .A1(n3776), .A2(n3820), .ZN(n3780) );
  AOI22_X1 U4688 ( .A1(EAX_REG_0__SCAN_IN), .A2(n3777), .B1(
        PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n6773), .ZN(n3779) );
  NAND2_X1 U4689 ( .A1(n3805), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3778) );
  NOR2_X1 U4690 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATEBS16_REG_SCAN_IN), .ZN(
        n3781) );
  NAND2_X1 U4691 ( .A1(n4851), .A2(n4179), .ZN(n3782) );
  NAND2_X1 U4692 ( .A1(n4854), .A2(n3782), .ZN(n6248) );
  NAND2_X1 U4693 ( .A1(n6249), .A2(n6248), .ZN(n6247) );
  NAND2_X1 U4694 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3799) );
  OAI21_X1 U4695 ( .B1(PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .A(n3799), .ZN(n6489) );
  NAND2_X1 U4696 ( .A1(n6489), .A2(n4179), .ZN(n3784) );
  NAND2_X1 U4697 ( .A1(STATEBS16_REG_SCAN_IN), .A2(n6773), .ZN(n3786) );
  AOI22_X1 U4698 ( .A1(PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n4213), .B1(n4214), 
        .B2(EAX_REG_2__SCAN_IN), .ZN(n3783) );
  NAND2_X1 U4699 ( .A1(n3784), .A2(n3783), .ZN(n3785) );
  AOI21_X1 U4700 ( .B1(n3805), .B2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(n3785), 
        .ZN(n3788) );
  NAND2_X1 U4701 ( .A1(n6247), .A2(n3788), .ZN(n5274) );
  OR2_X1 U4702 ( .A1(n6537), .A2(n3820), .ZN(n3787) );
  NAND2_X1 U4703 ( .A1(n3787), .A2(n3786), .ZN(n5273) );
  NAND2_X1 U4704 ( .A1(n5274), .A2(n5273), .ZN(n3792) );
  INV_X1 U4705 ( .A(n6247), .ZN(n3790) );
  INV_X1 U4706 ( .A(n3788), .ZN(n3789) );
  AOI21_X1 U4707 ( .B1(n3800), .B2(n3794), .A(n3811), .ZN(n6217) );
  AOI22_X1 U4708 ( .A1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n3805), .B1(n3777), .B2(EAX_REG_4__SCAN_IN), .ZN(n3796) );
  INV_X1 U4709 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n6081) );
  OAI21_X1 U4710 ( .B1(PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n6081), .A(n6773), 
        .ZN(n3795) );
  AOI22_X1 U4711 ( .A1(n4179), .A2(n6217), .B1(n3796), .B2(n3795), .ZN(n3797)
         );
  AOI21_X1 U4712 ( .B1(n3793), .B2(n3936), .A(n3797), .ZN(n4899) );
  INV_X1 U4713 ( .A(n4899), .ZN(n3808) );
  NAND2_X1 U4714 ( .A1(n3798), .A2(n3936), .ZN(n3807) );
  NAND2_X1 U4715 ( .A1(n4214), .A2(EAX_REG_3__SCAN_IN), .ZN(n3803) );
  INV_X1 U4716 ( .A(n3799), .ZN(n3801) );
  OAI21_X1 U4717 ( .B1(n3801), .B2(PHYADDRPOINTER_REG_3__SCAN_IN), .A(n3800), 
        .ZN(n6226) );
  AOI22_X1 U4718 ( .A1(PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n4213), .B1(n4179), 
        .B2(n6226), .ZN(n3802) );
  NAND2_X1 U4719 ( .A1(n3803), .A2(n3802), .ZN(n3804) );
  AOI21_X1 U4720 ( .B1(n3805), .B2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(n3804), 
        .ZN(n3806) );
  NAND2_X1 U4721 ( .A1(n3807), .A2(n3806), .ZN(n4907) );
  NAND2_X1 U4722 ( .A1(n3810), .A2(n3936), .ZN(n3815) );
  OAI21_X1 U4723 ( .B1(n3811), .B2(PHYADDRPOINTER_REG_5__SCAN_IN), .A(n3822), 
        .ZN(n6477) );
  AOI22_X1 U4724 ( .A1(PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n4213), .B1(n4179), 
        .B2(n6477), .ZN(n3812) );
  INV_X1 U4725 ( .A(n3812), .ZN(n3813) );
  AOI21_X1 U4726 ( .B1(n4214), .B2(EAX_REG_5__SCAN_IN), .A(n3813), .ZN(n3814)
         );
  OAI21_X1 U4727 ( .B1(PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n3816), .A(n3844), 
        .ZN(n6471) );
  AOI22_X1 U4728 ( .A1(n4214), .A2(EAX_REG_7__SCAN_IN), .B1(n3781), .B2(n6471), 
        .ZN(n3817) );
  XNOR2_X1 U4729 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .B(n3822), .ZN(n6195) );
  NAND2_X1 U4730 ( .A1(n3777), .A2(EAX_REG_6__SCAN_IN), .ZN(n3824) );
  OAI21_X1 U4731 ( .B1(PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n6081), .A(n6773), 
        .ZN(n3823) );
  AOI22_X1 U4732 ( .A1(n4179), .A2(n6195), .B1(n3824), .B2(n3823), .ZN(n3825)
         );
  INV_X1 U4733 ( .A(n5099), .ZN(n3827) );
  AOI22_X1 U4734 ( .A1(n3395), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n4191), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3833) );
  AOI22_X1 U4735 ( .A1(n4196), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4185), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3832) );
  AOI22_X1 U4736 ( .A1(n3349), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n4192), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3831) );
  AOI22_X1 U4737 ( .A1(n4167), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n4186), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3830) );
  NAND4_X1 U4738 ( .A1(n3833), .A2(n3832), .A3(n3831), .A4(n3830), .ZN(n3840)
         );
  AOI22_X1 U4739 ( .A1(n3208), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n4194), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3838) );
  AOI22_X1 U4740 ( .A1(n3180), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n3834), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3837) );
  AOI22_X1 U4741 ( .A1(n3524), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n4183), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3836) );
  AOI22_X1 U4742 ( .A1(n3207), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n3474), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3835) );
  NAND4_X1 U4743 ( .A1(n3838), .A2(n3837), .A3(n3836), .A4(n3835), .ZN(n3839)
         );
  OR2_X1 U4744 ( .A1(n3840), .A2(n3839), .ZN(n3843) );
  XNOR2_X1 U4745 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .B(n3844), .ZN(n6171) );
  AOI22_X1 U4746 ( .A1(PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n4213), .B1(n3777), 
        .B2(EAX_REG_8__SCAN_IN), .ZN(n3841) );
  OAI21_X1 U4747 ( .B1(n6171), .B2(n4773), .A(n3841), .ZN(n3842) );
  AOI21_X1 U4748 ( .B1(n3936), .B2(n3843), .A(n3842), .ZN(n5311) );
  AOI21_X1 U4749 ( .B1(n3845), .B2(n6164), .A(n3871), .ZN(n6167) );
  AOI22_X1 U4750 ( .A1(PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n4213), .B1(n3777), 
        .B2(EAX_REG_9__SCAN_IN), .ZN(n3857) );
  AOI22_X1 U4751 ( .A1(n3209), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4191), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3849) );
  AOI22_X1 U4752 ( .A1(n3396), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4194), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3848) );
  AOI22_X1 U4753 ( .A1(n4192), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3397), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3847) );
  AOI22_X1 U4754 ( .A1(n3207), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3474), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3846) );
  NAND4_X1 U4755 ( .A1(n3849), .A2(n3848), .A3(n3847), .A4(n3846), .ZN(n3855)
         );
  AOI22_X1 U4756 ( .A1(n3945), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3834), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3853) );
  AOI22_X1 U4757 ( .A1(n3178), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n4196), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3852) );
  AOI22_X1 U4758 ( .A1(n4184), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n4185), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3851) );
  AOI22_X1 U4759 ( .A1(n4193), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4186), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3850) );
  NAND4_X1 U4760 ( .A1(n3853), .A2(n3852), .A3(n3851), .A4(n3850), .ZN(n3854)
         );
  OAI21_X1 U4761 ( .B1(n3855), .B2(n3854), .A(n3936), .ZN(n3856) );
  OAI211_X1 U4762 ( .C1(n6167), .C2(n4773), .A(n3857), .B(n3856), .ZN(n5399)
         );
  AOI22_X1 U4763 ( .A1(n4195), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n4191), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3861) );
  AOI22_X1 U4764 ( .A1(n4184), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n4185), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3860) );
  AOI22_X1 U4765 ( .A1(n3180), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n4183), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3859) );
  AOI22_X1 U4766 ( .A1(n4192), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3207), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3858) );
  NAND4_X1 U4767 ( .A1(n3861), .A2(n3860), .A3(n3859), .A4(n3858), .ZN(n3867)
         );
  AOI22_X1 U4768 ( .A1(n3945), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n4182), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3865) );
  AOI22_X1 U4769 ( .A1(n4196), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4194), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3864) );
  AOI22_X1 U4770 ( .A1(n4193), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3474), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3863) );
  AOI22_X1 U4771 ( .A1(n4167), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n4186), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3862) );
  NAND4_X1 U4772 ( .A1(n3865), .A2(n3864), .A3(n3863), .A4(n3862), .ZN(n3866)
         );
  OR2_X1 U4773 ( .A1(n3867), .A2(n3866), .ZN(n3870) );
  XOR2_X1 U4774 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .B(n3871), .Z(n6151) );
  AOI22_X1 U4775 ( .A1(PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n4213), .B1(n3777), 
        .B2(EAX_REG_10__SCAN_IN), .ZN(n3868) );
  OAI21_X1 U4776 ( .B1(n6151), .B2(n4773), .A(n3868), .ZN(n3869) );
  AOI21_X1 U4777 ( .B1(n3936), .B2(n3870), .A(n3869), .ZN(n5470) );
  AOI21_X1 U4778 ( .B1(n3872), .B2(n6144), .A(n3895), .ZN(n6147) );
  AOI22_X1 U4779 ( .A1(PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n4213), .B1(n3777), 
        .B2(EAX_REG_11__SCAN_IN), .ZN(n3884) );
  AOI22_X1 U4780 ( .A1(n3945), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4191), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3876) );
  AOI22_X1 U4781 ( .A1(n3209), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4195), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3875) );
  AOI22_X1 U4782 ( .A1(n3178), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n4184), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3874) );
  AOI22_X1 U4783 ( .A1(n4193), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3397), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3873) );
  NAND4_X1 U4784 ( .A1(n3876), .A2(n3875), .A3(n3874), .A4(n3873), .ZN(n3882)
         );
  AOI22_X1 U4785 ( .A1(n3396), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4194), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3880) );
  AOI22_X1 U4786 ( .A1(n4185), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3207), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3879) );
  AOI22_X1 U4787 ( .A1(n4192), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4186), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3878) );
  AOI22_X1 U4788 ( .A1(n4196), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3474), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3877) );
  NAND4_X1 U4789 ( .A1(n3880), .A2(n3879), .A3(n3878), .A4(n3877), .ZN(n3881)
         );
  OAI21_X1 U4790 ( .B1(n3882), .B2(n3881), .A(n3936), .ZN(n3883) );
  OAI211_X1 U4791 ( .C1(n6147), .C2(n4773), .A(n3884), .B(n3883), .ZN(n5478)
         );
  AOI22_X1 U4792 ( .A1(n3209), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n4191), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3888) );
  AOI22_X1 U4793 ( .A1(n4196), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3524), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3887) );
  AOI22_X1 U4794 ( .A1(n4185), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3207), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3886) );
  AOI22_X1 U4795 ( .A1(n4192), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3397), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3885) );
  NAND4_X1 U4796 ( .A1(n3888), .A2(n3887), .A3(n3886), .A4(n3885), .ZN(n3894)
         );
  AOI22_X1 U4797 ( .A1(n3180), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n3457), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3892) );
  AOI22_X1 U4798 ( .A1(n3945), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n4194), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3891) );
  AOI22_X1 U4799 ( .A1(n4183), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3474), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3890) );
  AOI22_X1 U4800 ( .A1(n4193), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n4186), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3889) );
  NAND4_X1 U4801 ( .A1(n3892), .A2(n3891), .A3(n3890), .A4(n3889), .ZN(n3893)
         );
  OR2_X1 U4802 ( .A1(n3894), .A2(n3893), .ZN(n3899) );
  OAI21_X1 U4803 ( .B1(n3895), .B2(PHYADDRPOINTER_REG_12__SCAN_IN), .A(n3900), 
        .ZN(n3896) );
  INV_X1 U4804 ( .A(n3896), .ZN(n6134) );
  AOI22_X1 U4805 ( .A1(PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n4213), .B1(n3777), 
        .B2(EAX_REG_12__SCAN_IN), .ZN(n3897) );
  OAI21_X1 U4806 ( .B1(n6134), .B2(n4773), .A(n3897), .ZN(n3898) );
  AOI21_X1 U4807 ( .B1(n3936), .B2(n3899), .A(n3898), .ZN(n5506) );
  AOI21_X1 U4808 ( .B1(n6128), .B2(n3900), .A(n3923), .ZN(n6132) );
  AOI22_X1 U4809 ( .A1(PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n4213), .B1(n3777), 
        .B2(EAX_REG_13__SCAN_IN), .ZN(n3912) );
  AOI22_X1 U4810 ( .A1(n3945), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n4191), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3904) );
  AOI22_X1 U4811 ( .A1(n3180), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n3457), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3903) );
  AOI22_X1 U4812 ( .A1(n4196), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4185), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3902) );
  AOI22_X1 U4813 ( .A1(n3209), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4194), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3901) );
  NAND4_X1 U4814 ( .A1(n3904), .A2(n3903), .A3(n3902), .A4(n3901), .ZN(n3910)
         );
  AOI22_X1 U4815 ( .A1(n4193), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4192), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3908) );
  AOI22_X1 U4816 ( .A1(n4184), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n4183), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3907) );
  AOI22_X1 U4817 ( .A1(n3207), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3474), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3906) );
  AOI22_X1 U4818 ( .A1(n4167), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n4186), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3905) );
  NAND4_X1 U4819 ( .A1(n3908), .A2(n3907), .A3(n3906), .A4(n3905), .ZN(n3909)
         );
  OAI21_X1 U4820 ( .B1(n3910), .B2(n3909), .A(n3936), .ZN(n3911) );
  OAI211_X1 U4821 ( .C1(n6132), .C2(n4773), .A(n3912), .B(n3911), .ZN(n5533)
         );
  AOI22_X1 U4822 ( .A1(n4195), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n4184), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3916) );
  AOI22_X1 U4823 ( .A1(n4193), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4185), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3915) );
  AOI22_X1 U4824 ( .A1(n3945), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n4194), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3914) );
  AOI22_X1 U4825 ( .A1(n4167), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n4186), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3913) );
  NAND4_X1 U4826 ( .A1(n3916), .A2(n3915), .A3(n3914), .A4(n3913), .ZN(n3922)
         );
  AOI22_X1 U4827 ( .A1(n3209), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4191), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3920) );
  AOI22_X1 U4828 ( .A1(n3178), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n4183), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3919) );
  AOI22_X1 U4829 ( .A1(n4196), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3474), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3918) );
  AOI22_X1 U4830 ( .A1(n4192), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3207), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3917) );
  NAND4_X1 U4831 ( .A1(n3920), .A2(n3919), .A3(n3918), .A4(n3917), .ZN(n3921)
         );
  OR2_X1 U4832 ( .A1(n3922), .A2(n3921), .ZN(n3927) );
  AOI21_X1 U4833 ( .B1(n3924), .B2(n6118), .A(n3950), .ZN(n6120) );
  AOI22_X1 U4834 ( .A1(PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n4213), .B1(n3777), 
        .B2(EAX_REG_14__SCAN_IN), .ZN(n3925) );
  OAI21_X1 U4835 ( .B1(n6120), .B2(n4773), .A(n3925), .ZN(n3926) );
  AOI21_X1 U4836 ( .B1(n3936), .B2(n3927), .A(n3926), .ZN(n5545) );
  XOR2_X1 U4837 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .B(n3950), .Z(n6112) );
  AOI22_X1 U4838 ( .A1(PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n4213), .B1(n4214), 
        .B2(EAX_REG_15__SCAN_IN), .ZN(n3940) );
  AOI22_X1 U4839 ( .A1(INSTQUEUE_REG_7__7__SCAN_IN), .A2(n3945), .B1(n3178), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3931) );
  AOI22_X1 U4840 ( .A1(INSTQUEUE_REG_8__7__SCAN_IN), .A2(n4193), .B1(n4192), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3930) );
  AOI22_X1 U4841 ( .A1(n4185), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3474), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3929) );
  AOI22_X1 U4842 ( .A1(INSTQUEUE_REG_2__7__SCAN_IN), .A2(n4167), .B1(n4186), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3928) );
  NAND4_X1 U4843 ( .A1(n3931), .A2(n3930), .A3(n3929), .A4(n3928), .ZN(n3938)
         );
  AOI22_X1 U4844 ( .A1(n3208), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4191), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3935) );
  AOI22_X1 U4845 ( .A1(n4195), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n4194), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3934) );
  AOI22_X1 U4846 ( .A1(n4196), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4183), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3933) );
  AOI22_X1 U4847 ( .A1(n4184), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n3207), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3932) );
  NAND4_X1 U4848 ( .A1(n3935), .A2(n3934), .A3(n3933), .A4(n3932), .ZN(n3937)
         );
  OAI21_X1 U4849 ( .B1(n3938), .B2(n3937), .A(n3936), .ZN(n3939) );
  OAI211_X1 U4850 ( .C1(n6112), .C2(n4773), .A(n3940), .B(n3939), .ZN(n5756)
         );
  AOI22_X1 U4851 ( .A1(n3208), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n4191), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3944) );
  AOI22_X1 U4852 ( .A1(n4196), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4183), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3943) );
  AOI22_X1 U4853 ( .A1(n4184), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n3207), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3942) );
  AOI22_X1 U4854 ( .A1(n4192), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4186), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3941) );
  NAND4_X1 U4855 ( .A1(n3944), .A2(n3943), .A3(n3942), .A4(n3941), .ZN(n3954)
         );
  AOI22_X1 U4856 ( .A1(n3180), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n3457), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3949) );
  AOI22_X1 U4857 ( .A1(n3945), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n4194), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3948) );
  AOI22_X1 U4858 ( .A1(n4193), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3397), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3947) );
  AOI22_X1 U4859 ( .A1(n4185), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3474), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3946) );
  NAND4_X1 U4860 ( .A1(n3949), .A2(n3948), .A3(n3947), .A4(n3946), .ZN(n3953)
         );
  XNOR2_X1 U4861 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .B(n3955), .ZN(n6108)
         );
  AOI22_X1 U4862 ( .A1(PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n4213), .B1(n3777), 
        .B2(EAX_REG_16__SCAN_IN), .ZN(n3951) );
  OAI21_X1 U4863 ( .B1(n6108), .B2(n4773), .A(n3951), .ZN(n3952) );
  AOI221_X1 U4864 ( .B1(n3954), .B2(n4206), .C1(n3953), .C2(n4206), .A(n3952), 
        .ZN(n5589) );
  XOR2_X1 U4865 ( .A(PHYADDRPOINTER_REG_17__SCAN_IN), .B(n3968), .Z(n5992) );
  AOI22_X1 U4866 ( .A1(EAX_REG_17__SCAN_IN), .A2(n4214), .B1(
        PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n6773), .ZN(n3967) );
  AOI22_X1 U4867 ( .A1(n3209), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4191), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3959) );
  AOI22_X1 U4868 ( .A1(n4193), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4185), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3958) );
  AOI22_X1 U4869 ( .A1(n4184), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n3474), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3957) );
  AOI22_X1 U4870 ( .A1(n4192), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4186), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3956) );
  NAND4_X1 U4871 ( .A1(n3959), .A2(n3958), .A3(n3957), .A4(n3956), .ZN(n3965)
         );
  AOI22_X1 U4872 ( .A1(n3945), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3394), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3963) );
  AOI22_X1 U4873 ( .A1(n3180), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n4195), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3962) );
  AOI22_X1 U4874 ( .A1(n4196), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3396), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3961) );
  AOI22_X1 U4875 ( .A1(n4167), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n3207), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3960) );
  NAND4_X1 U4876 ( .A1(n3963), .A2(n3962), .A3(n3961), .A4(n3960), .ZN(n3964)
         );
  AOI221_X1 U4877 ( .B1(n3965), .B2(n4206), .C1(n3964), .C2(n4206), .A(n3781), 
        .ZN(n3966) );
  AOI22_X1 U4878 ( .A1(n3781), .A2(n5992), .B1(n3967), .B2(n3966), .ZN(n5569)
         );
  OAI21_X1 U4879 ( .B1(n3969), .B2(PHYADDRPOINTER_REG_18__SCAN_IN), .A(n3995), 
        .ZN(n6098) );
  AOI22_X1 U4880 ( .A1(EAX_REG_18__SCAN_IN), .A2(n4214), .B1(
        PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n6773), .ZN(n3981) );
  AOI22_X1 U4881 ( .A1(n3208), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4191), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3973) );
  AOI22_X1 U4882 ( .A1(n4195), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n4194), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3972) );
  AOI22_X1 U4883 ( .A1(n4184), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n4183), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3971) );
  AOI22_X1 U4884 ( .A1(n4192), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3207), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3970) );
  NAND4_X1 U4885 ( .A1(n3973), .A2(n3972), .A3(n3971), .A4(n3970), .ZN(n3979)
         );
  AOI22_X1 U4886 ( .A1(n3945), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3180), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3977) );
  AOI22_X1 U4887 ( .A1(n4193), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4185), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3976) );
  AOI22_X1 U4888 ( .A1(n4196), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3474), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3975) );
  AOI22_X1 U4889 ( .A1(n4167), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n4186), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3974) );
  NAND4_X1 U4890 ( .A1(n3977), .A2(n3976), .A3(n3975), .A4(n3974), .ZN(n3978)
         );
  OAI21_X1 U4891 ( .B1(n3979), .B2(n3978), .A(n4206), .ZN(n3980) );
  NAND3_X1 U4892 ( .A1(n4773), .A2(n3981), .A3(n3980), .ZN(n3982) );
  OAI21_X1 U4893 ( .B1(n4773), .B2(n6098), .A(n3982), .ZN(n5988) );
  XNOR2_X1 U4894 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .B(n3995), .ZN(n5981)
         );
  AOI22_X1 U4895 ( .A1(EAX_REG_19__SCAN_IN), .A2(n4214), .B1(
        PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n6773), .ZN(n3994) );
  AOI22_X1 U4896 ( .A1(n4182), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4191), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3986) );
  AOI22_X1 U4897 ( .A1(n4192), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3207), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3985) );
  AOI22_X1 U4898 ( .A1(n4167), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n4186), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3984) );
  AOI22_X1 U4899 ( .A1(n4195), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3474), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3983) );
  NAND4_X1 U4900 ( .A1(n3986), .A2(n3985), .A3(n3984), .A4(n3983), .ZN(n3992)
         );
  AOI22_X1 U4901 ( .A1(n4196), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4184), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3990) );
  AOI22_X1 U4902 ( .A1(n4193), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4185), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3989) );
  AOI22_X1 U4903 ( .A1(n3945), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3394), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3988) );
  AOI22_X1 U4904 ( .A1(n3178), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3396), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3987) );
  NAND4_X1 U4905 ( .A1(n3990), .A2(n3989), .A3(n3988), .A4(n3987), .ZN(n3991)
         );
  AOI221_X1 U4906 ( .B1(n3992), .B2(n4206), .C1(n3991), .C2(n4206), .A(n3781), 
        .ZN(n3993) );
  AOI22_X1 U4907 ( .A1(n4179), .A2(n5981), .B1(n3994), .B2(n3993), .ZN(n5876)
         );
  INV_X1 U4908 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n5882) );
  OAI21_X1 U4909 ( .B1(n3996), .B2(PHYADDRPOINTER_REG_20__SCAN_IN), .A(n4023), 
        .ZN(n5979) );
  AOI22_X1 U4910 ( .A1(EAX_REG_20__SCAN_IN), .A2(n4214), .B1(
        PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n6773), .ZN(n4008) );
  AOI22_X1 U4911 ( .A1(n3945), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n4194), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n4000) );
  AOI22_X1 U4912 ( .A1(n4193), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n4192), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3999) );
  AOI22_X1 U4913 ( .A1(n4196), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3396), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3998) );
  AOI22_X1 U4914 ( .A1(n3207), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n3474), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3997) );
  NAND4_X1 U4915 ( .A1(n4000), .A2(n3999), .A3(n3998), .A4(n3997), .ZN(n4006)
         );
  AOI22_X1 U4916 ( .A1(n4182), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4076), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4004) );
  AOI22_X1 U4917 ( .A1(n3178), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n4195), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4003) );
  AOI22_X1 U4918 ( .A1(n4184), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n4185), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4002) );
  AOI22_X1 U4919 ( .A1(n4167), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n4186), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n4001) );
  NAND4_X1 U4920 ( .A1(n4004), .A2(n4003), .A3(n4002), .A4(n4001), .ZN(n4005)
         );
  OAI21_X1 U4921 ( .B1(n4006), .B2(n4005), .A(n4206), .ZN(n4007) );
  NAND3_X1 U4922 ( .A1(n4773), .A2(n4008), .A3(n4007), .ZN(n4009) );
  OAI21_X1 U4923 ( .B1(n4773), .B2(n5979), .A(n4009), .ZN(n5861) );
  XNOR2_X1 U4924 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .B(n4023), .ZN(n5967)
         );
  AOI22_X1 U4925 ( .A1(EAX_REG_21__SCAN_IN), .A2(n4214), .B1(
        PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n6773), .ZN(n4021) );
  AOI22_X1 U4926 ( .A1(n4196), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4184), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4013) );
  AOI22_X1 U4927 ( .A1(n4195), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n4183), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4012) );
  AOI22_X1 U4928 ( .A1(n4193), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3207), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4011) );
  AOI22_X1 U4929 ( .A1(n4192), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4186), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4010) );
  NAND4_X1 U4930 ( .A1(n4013), .A2(n4012), .A3(n4011), .A4(n4010), .ZN(n4019)
         );
  AOI22_X1 U4931 ( .A1(n3945), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4191), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4017) );
  AOI22_X1 U4932 ( .A1(n3209), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3394), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n4016) );
  AOI22_X1 U4933 ( .A1(n4185), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n4167), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4015) );
  AOI22_X1 U4934 ( .A1(n3178), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3474), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4014) );
  NAND4_X1 U4935 ( .A1(n4017), .A2(n4016), .A3(n4015), .A4(n4014), .ZN(n4018)
         );
  AOI221_X1 U4936 ( .B1(n4019), .B2(n4206), .C1(n4018), .C2(n4206), .A(n3781), 
        .ZN(n4020) );
  AOI22_X1 U4937 ( .A1(n4179), .A2(n5967), .B1(n4021), .B2(n4020), .ZN(n5855)
         );
  INV_X1 U4938 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n4022) );
  OAI21_X1 U4939 ( .B1(n4024), .B2(PHYADDRPOINTER_REG_22__SCAN_IN), .A(n4073), 
        .ZN(n5839) );
  AOI22_X1 U4940 ( .A1(EAX_REG_22__SCAN_IN), .A2(n4214), .B1(
        PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n6773), .ZN(n4036) );
  AOI22_X1 U4941 ( .A1(n3209), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4076), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4028) );
  AOI22_X1 U4942 ( .A1(n4195), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n4183), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4027) );
  AOI22_X1 U4943 ( .A1(n4196), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3207), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4026) );
  AOI22_X1 U4944 ( .A1(n4192), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4186), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n4025) );
  NAND4_X1 U4945 ( .A1(n4028), .A2(n4027), .A3(n4026), .A4(n4025), .ZN(n4034)
         );
  AOI22_X1 U4946 ( .A1(n3180), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n4184), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4032) );
  AOI22_X1 U4947 ( .A1(n3945), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4194), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n4031) );
  AOI22_X1 U4948 ( .A1(n4193), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4167), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4030) );
  AOI22_X1 U4949 ( .A1(n3475), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3474), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4029) );
  NAND4_X1 U4950 ( .A1(n4032), .A2(n4031), .A3(n4030), .A4(n4029), .ZN(n4033)
         );
  OAI21_X1 U4951 ( .B1(n4034), .B2(n4033), .A(n4206), .ZN(n4035) );
  NAND3_X1 U4952 ( .A1(n4773), .A2(n4036), .A3(n4035), .ZN(n4037) );
  OAI21_X1 U4953 ( .B1(n4773), .B2(n5839), .A(n4037), .ZN(n4038) );
  AND2_X1 U4954 ( .A1(n4039), .A2(n4038), .ZN(n4040) );
  OR2_X1 U4955 ( .A1(n4040), .A2(n4072), .ZN(n5917) );
  NAND3_X1 U4956 ( .A1(n6894), .A2(STATEBS16_REG_SCAN_IN), .A3(
        STATE2_REG_1__SCAN_IN), .ZN(n6907) );
  NAND2_X1 U4957 ( .A1(n4044), .A2(n6776), .ZN(n7023) );
  AND2_X1 U4958 ( .A1(n7023), .A2(n6894), .ZN(n4041) );
  NAND2_X1 U4959 ( .A1(n6894), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4043) );
  NAND2_X1 U4960 ( .A1(n6081), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4042) );
  NAND2_X1 U4961 ( .A1(n4043), .A2(n4042), .ZN(n4850) );
  AOI22_X1 U4962 ( .A1(PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n6491), .B1(n6523), 
        .B2(REIP_REG_22__SCAN_IN), .ZN(n4045) );
  OAI21_X1 U4963 ( .B1(n6005), .B2(n6484), .A(n4047), .ZN(U2964) );
  XNOR2_X1 U4964 ( .A(n4073), .B(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5833)
         );
  AOI22_X1 U4965 ( .A1(EAX_REG_23__SCAN_IN), .A2(n4214), .B1(
        PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n6773), .ZN(n4070) );
  AOI22_X1 U4966 ( .A1(n3209), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4191), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n4051) );
  AOI22_X1 U4967 ( .A1(n4195), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n4194), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n4050) );
  AOI22_X1 U4968 ( .A1(n4185), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3474), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4049) );
  AOI22_X1 U4969 ( .A1(n4167), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n4186), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n4048) );
  NAND4_X1 U4970 ( .A1(n4051), .A2(n4050), .A3(n4049), .A4(n4048), .ZN(n4057)
         );
  AOI22_X1 U4971 ( .A1(n3945), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3178), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4055) );
  AOI22_X1 U4972 ( .A1(n4193), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n4192), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n4054) );
  AOI22_X1 U4973 ( .A1(n4196), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n4183), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4053) );
  AOI22_X1 U4974 ( .A1(n4184), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n3207), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4052) );
  NAND4_X1 U4975 ( .A1(n4055), .A2(n4054), .A3(n4053), .A4(n4052), .ZN(n4056)
         );
  NOR2_X1 U4976 ( .A1(n4057), .A2(n4056), .ZN(n4075) );
  AOI22_X1 U4977 ( .A1(n4196), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4184), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4061) );
  AOI22_X1 U4978 ( .A1(n3180), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n4194), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n4060) );
  AOI22_X1 U4979 ( .A1(n4185), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3207), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4059) );
  AOI22_X1 U4980 ( .A1(INSTQUEUE_REG_3__7__SCAN_IN), .A2(n4167), .B1(n4186), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4058) );
  NAND4_X1 U4981 ( .A1(n4061), .A2(n4060), .A3(n4059), .A4(n4058), .ZN(n4067)
         );
  AOI22_X1 U4982 ( .A1(n3945), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n4191), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4065) );
  AOI22_X1 U4983 ( .A1(n3208), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4195), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4064) );
  AOI22_X1 U4984 ( .A1(n4193), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4192), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n4063) );
  AOI22_X1 U4985 ( .A1(n4183), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3474), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4062) );
  NAND4_X1 U4986 ( .A1(n4065), .A2(n4064), .A3(n4063), .A4(n4062), .ZN(n4066)
         );
  NOR2_X1 U4987 ( .A1(n4067), .A2(n4066), .ZN(n4074) );
  XOR2_X1 U4988 ( .A(n4075), .B(n4074), .Z(n4068) );
  AOI21_X1 U4989 ( .B1(n4206), .B2(n4068), .A(n4179), .ZN(n4069) );
  AND2_X1 U4990 ( .A1(n4070), .A2(n4069), .ZN(n4071) );
  AOI21_X1 U4991 ( .B1(n5833), .B2(n4179), .A(n4071), .ZN(n5641) );
  INV_X1 U4992 ( .A(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5639) );
  XNOR2_X1 U4993 ( .A(n4093), .B(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5826)
         );
  INV_X1 U4994 ( .A(n5826), .ZN(n4092) );
  OR2_X1 U4995 ( .A1(n4075), .A2(n4074), .ZN(n4096) );
  AOI22_X1 U4996 ( .A1(n4076), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n4183), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4080) );
  AOI22_X1 U4997 ( .A1(n3178), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n4195), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n4079) );
  AOI22_X1 U4998 ( .A1(n4185), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4194), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n4078) );
  AOI22_X1 U4999 ( .A1(n4196), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3474), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4077) );
  NAND4_X1 U5000 ( .A1(n4080), .A2(n4079), .A3(n4078), .A4(n4077), .ZN(n4086)
         );
  AOI22_X1 U5001 ( .A1(n4182), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4184), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n4084) );
  AOI22_X1 U5002 ( .A1(n4193), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3207), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4083) );
  AOI22_X1 U5003 ( .A1(n3945), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4167), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4082) );
  AOI22_X1 U5004 ( .A1(n4192), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4186), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n4081) );
  NAND4_X1 U5005 ( .A1(n4084), .A2(n4083), .A3(n4082), .A4(n4081), .ZN(n4085)
         );
  NOR2_X1 U5006 ( .A1(n4086), .A2(n4085), .ZN(n4095) );
  OAI21_X1 U5007 ( .B1(n4095), .B2(n4096), .A(n4206), .ZN(n4087) );
  AOI21_X1 U5008 ( .B1(n4096), .B2(n4095), .A(n4087), .ZN(n4088) );
  INV_X1 U5009 ( .A(n4088), .ZN(n4090) );
  AOI22_X1 U5010 ( .A1(n4214), .A2(EAX_REG_24__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n4213), .ZN(n4089) );
  NAND2_X1 U5011 ( .A1(n4090), .A2(n4089), .ZN(n4091) );
  AOI21_X1 U5012 ( .B1(n4092), .B2(n4179), .A(n4091), .ZN(n5627) );
  INV_X1 U5013 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5630) );
  INV_X1 U5014 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n4389) );
  AOI21_X1 U5015 ( .B1(n4094), .B2(n4389), .A(n4110), .ZN(n5819) );
  AOI22_X1 U5016 ( .A1(EAX_REG_25__SCAN_IN), .A2(n4214), .B1(
        PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n6773), .ZN(n4109) );
  OR2_X1 U5017 ( .A1(n4096), .A2(n4095), .ZN(n4111) );
  AOI22_X1 U5018 ( .A1(n3209), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4191), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4100) );
  AOI22_X1 U5019 ( .A1(n3178), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3457), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n4099) );
  AOI22_X1 U5020 ( .A1(n4196), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4184), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n4098) );
  AOI22_X1 U5021 ( .A1(n4193), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4186), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n4097) );
  NAND4_X1 U5022 ( .A1(n4100), .A2(n4099), .A3(n4098), .A4(n4097), .ZN(n4106)
         );
  AOI22_X1 U5023 ( .A1(n3945), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4194), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n4104) );
  AOI22_X1 U5024 ( .A1(n4192), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3397), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4103) );
  AOI22_X1 U5025 ( .A1(n4185), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3207), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4102) );
  AOI22_X1 U5026 ( .A1(n3396), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n3474), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4101) );
  NAND4_X1 U5027 ( .A1(n4104), .A2(n4103), .A3(n4102), .A4(n4101), .ZN(n4105)
         );
  NOR2_X1 U5028 ( .A1(n4106), .A2(n4105), .ZN(n4112) );
  XOR2_X1 U5029 ( .A(n4111), .B(n4112), .Z(n4107) );
  AOI21_X1 U5030 ( .B1(n4107), .B2(n4206), .A(n3781), .ZN(n4108) );
  AOI22_X1 U5031 ( .A1(n4179), .A2(n5819), .B1(n4109), .B2(n4108), .ZN(n5617)
         );
  OAI21_X1 U5032 ( .B1(n4110), .B2(PHYADDRPOINTER_REG_26__SCAN_IN), .A(n4141), 
        .ZN(n5966) );
  INV_X1 U5033 ( .A(n4206), .ZN(n4175) );
  NOR2_X1 U5034 ( .A1(n4112), .A2(n4111), .ZN(n4137) );
  AOI22_X1 U5035 ( .A1(n3945), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4191), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4116) );
  AOI22_X1 U5036 ( .A1(n3180), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n4195), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n4115) );
  AOI22_X1 U5037 ( .A1(n4182), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4194), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n4114) );
  AOI22_X1 U5038 ( .A1(n4196), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4183), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4113) );
  NAND4_X1 U5039 ( .A1(n4116), .A2(n4115), .A3(n4114), .A4(n4113), .ZN(n4122)
         );
  AOI22_X1 U5040 ( .A1(n4193), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4192), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n4120) );
  AOI22_X1 U5041 ( .A1(n4184), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3474), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4119) );
  INV_X1 U5042 ( .A(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n4568) );
  AOI22_X1 U5043 ( .A1(n4185), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3207), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4118) );
  AOI22_X1 U5044 ( .A1(n4167), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n4186), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n4117) );
  NAND4_X1 U5045 ( .A1(n4120), .A2(n4119), .A3(n4118), .A4(n4117), .ZN(n4121)
         );
  OR2_X1 U5046 ( .A1(n4122), .A2(n4121), .ZN(n4136) );
  XNOR2_X1 U5047 ( .A(n4137), .B(n4136), .ZN(n4124) );
  AOI22_X1 U5048 ( .A1(EAX_REG_26__SCAN_IN), .A2(n4214), .B1(
        PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n6773), .ZN(n4123) );
  OAI21_X1 U5049 ( .B1(n4175), .B2(n4124), .A(n4123), .ZN(n4125) );
  AOI22_X1 U5050 ( .A1(n4179), .A2(n5966), .B1(n4125), .B2(n4773), .ZN(n5808)
         );
  XNOR2_X1 U5051 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .B(n4141), .ZN(n5956)
         );
  AOI22_X1 U5052 ( .A1(n4195), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n4196), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4129) );
  AOI22_X1 U5053 ( .A1(n4193), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3207), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4128) );
  AOI22_X1 U5054 ( .A1(n4192), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3397), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4127) );
  AOI22_X1 U5055 ( .A1(n4184), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n3474), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4126) );
  NAND4_X1 U5056 ( .A1(n4129), .A2(n4128), .A3(n4127), .A4(n4126), .ZN(n4135)
         );
  AOI22_X1 U5057 ( .A1(n3945), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n4191), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4133) );
  AOI22_X1 U5058 ( .A1(n3208), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4194), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n4132) );
  AOI22_X1 U5059 ( .A1(n3180), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n4183), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4131) );
  AOI22_X1 U5060 ( .A1(n4185), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n4186), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4130) );
  NAND4_X1 U5061 ( .A1(n4133), .A2(n4132), .A3(n4131), .A4(n4130), .ZN(n4134)
         );
  NOR2_X1 U5062 ( .A1(n4135), .A2(n4134), .ZN(n4154) );
  NAND2_X1 U5063 ( .A1(n4137), .A2(n4136), .ZN(n4153) );
  XOR2_X1 U5064 ( .A(n4154), .B(n4153), .Z(n4138) );
  AOI22_X1 U5065 ( .A1(n4206), .A2(n4138), .B1(n4214), .B2(EAX_REG_27__SCAN_IN), .ZN(n4140) );
  OAI21_X1 U5066 ( .B1(PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n6081), .A(n6773), 
        .ZN(n4139) );
  AOI22_X1 U5067 ( .A1(n4179), .A2(n5956), .B1(n4140), .B2(n4139), .ZN(n5799)
         );
  INV_X1 U5068 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5804) );
  NAND2_X1 U5069 ( .A1(n4142), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n4159)
         );
  OAI21_X1 U5070 ( .B1(n4142), .B2(PHYADDRPOINTER_REG_28__SCAN_IN), .A(n4159), 
        .ZN(n5786) );
  AOI22_X1 U5071 ( .A1(n4195), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n4191), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4146) );
  AOI22_X1 U5072 ( .A1(n4196), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n4183), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4145) );
  AOI22_X1 U5073 ( .A1(n4193), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3397), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4144) );
  AOI22_X1 U5074 ( .A1(n3475), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3207), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4143) );
  NAND4_X1 U5075 ( .A1(n4146), .A2(n4145), .A3(n4144), .A4(n4143), .ZN(n4152)
         );
  AOI22_X1 U5076 ( .A1(n3945), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3208), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n4150) );
  AOI22_X1 U5077 ( .A1(n3180), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3394), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n4149) );
  AOI22_X1 U5078 ( .A1(n4184), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3474), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4148) );
  AOI22_X1 U5079 ( .A1(n4192), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4186), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4147) );
  NAND4_X1 U5080 ( .A1(n4150), .A2(n4149), .A3(n4148), .A4(n4147), .ZN(n4151)
         );
  NOR2_X1 U5081 ( .A1(n4152), .A2(n4151), .ZN(n4162) );
  XNOR2_X1 U5082 ( .A(n4162), .B(n4161), .ZN(n4156) );
  AOI22_X1 U5083 ( .A1(EAX_REG_28__SCAN_IN), .A2(n4214), .B1(
        PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n6773), .ZN(n4155) );
  OAI21_X1 U5084 ( .B1(n4156), .B2(n4175), .A(n4155), .ZN(n4157) );
  AOI22_X1 U5085 ( .A1(n3781), .A2(n5786), .B1(n4157), .B2(n4773), .ZN(n4766)
         );
  INV_X1 U5086 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4158) );
  NAND2_X1 U5087 ( .A1(n4159), .A2(n4158), .ZN(n4160) );
  NAND2_X1 U5088 ( .A1(n4235), .A2(n4160), .ZN(n5778) );
  AOI22_X1 U5089 ( .A1(n3945), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3209), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n4166) );
  AOI22_X1 U5090 ( .A1(n4195), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4194), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n4165) );
  AOI22_X1 U5091 ( .A1(n3178), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3207), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4164) );
  AOI22_X1 U5092 ( .A1(n4192), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4186), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4163) );
  NAND4_X1 U5093 ( .A1(n4166), .A2(n4165), .A3(n4164), .A4(n4163), .ZN(n4173)
         );
  AOI22_X1 U5094 ( .A1(n4196), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4184), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4171) );
  AOI22_X1 U5095 ( .A1(n4076), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n4183), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4170) );
  AOI22_X1 U5096 ( .A1(n4193), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4167), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4169) );
  AOI22_X1 U5097 ( .A1(n3475), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3474), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4168) );
  NAND4_X1 U5098 ( .A1(n4171), .A2(n4170), .A3(n4169), .A4(n4168), .ZN(n4172)
         );
  NOR2_X1 U5099 ( .A1(n4173), .A2(n4172), .ZN(n4180) );
  XNOR2_X1 U5100 ( .A(n4181), .B(n4180), .ZN(n4176) );
  AOI22_X1 U5101 ( .A1(EAX_REG_29__SCAN_IN), .A2(n4214), .B1(
        PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n6773), .ZN(n4174) );
  OAI211_X1 U5102 ( .C1(n4176), .C2(n4175), .A(n4174), .B(n4773), .ZN(n4177)
         );
  OAI21_X1 U5103 ( .B1(n5778), .B2(n4773), .A(n4177), .ZN(n4178) );
  INV_X1 U5104 ( .A(n4178), .ZN(n4246) );
  INV_X1 U5105 ( .A(n5605), .ZN(n4212) );
  XNOR2_X1 U5106 ( .A(n4235), .B(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5771)
         );
  NAND2_X1 U5107 ( .A1(n5771), .A2(n4179), .ZN(n4210) );
  NOR2_X1 U5108 ( .A1(n4181), .A2(n4180), .ZN(n4204) );
  AOI22_X1 U5109 ( .A1(n3208), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3178), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4190) );
  AOI22_X1 U5110 ( .A1(INSTQUEUE_REG_1__7__SCAN_IN), .A2(n4184), .B1(n4183), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4189) );
  AOI22_X1 U5111 ( .A1(n4185), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3207), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4188) );
  AOI22_X1 U5112 ( .A1(INSTQUEUE_REG_4__7__SCAN_IN), .A2(n4167), .B1(n4186), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4187) );
  NAND4_X1 U5113 ( .A1(n4190), .A2(n4189), .A3(n4188), .A4(n4187), .ZN(n4202)
         );
  AOI22_X1 U5114 ( .A1(n3945), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4191), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4200) );
  AOI22_X1 U5115 ( .A1(INSTQUEUE_REG_10__7__SCAN_IN), .A2(n4193), .B1(n4192), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n4199) );
  AOI22_X1 U5116 ( .A1(n4195), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n4194), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n4198) );
  AOI22_X1 U5117 ( .A1(n4196), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3474), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4197) );
  NAND4_X1 U5118 ( .A1(n4200), .A2(n4199), .A3(n4198), .A4(n4197), .ZN(n4201)
         );
  NOR2_X1 U5119 ( .A1(n4202), .A2(n4201), .ZN(n4203) );
  XNOR2_X1 U5120 ( .A(n4204), .B(n4203), .ZN(n4205) );
  AOI21_X1 U5121 ( .B1(n4206), .B2(n4205), .A(n3781), .ZN(n4208) );
  AOI22_X1 U5122 ( .A1(EAX_REG_30__SCAN_IN), .A2(n4214), .B1(
        PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n6773), .ZN(n4207) );
  NAND2_X1 U5123 ( .A1(n4208), .A2(n4207), .ZN(n4209) );
  NAND2_X1 U5124 ( .A1(n4210), .A2(n4209), .ZN(n5606) );
  INV_X1 U5125 ( .A(n5606), .ZN(n4211) );
  NAND2_X1 U5126 ( .A1(n4212), .A2(n4211), .ZN(n4216) );
  AOI22_X1 U5127 ( .A1(n4214), .A2(EAX_REG_31__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n4213), .ZN(n4215) );
  XNOR2_X2 U5128 ( .A(n4216), .B(n4215), .ZN(n5768) );
  NAND2_X1 U5129 ( .A1(n6017), .A2(n6031), .ZN(n6022) );
  INV_X1 U5130 ( .A(n6022), .ZN(n4219) );
  INV_X1 U5131 ( .A(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n4217) );
  NAND2_X1 U5132 ( .A1(n4217), .A2(n5730), .ZN(n6009) );
  INV_X1 U5133 ( .A(n6009), .ZN(n4218) );
  INV_X1 U5134 ( .A(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5700) );
  INV_X1 U5135 ( .A(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5716) );
  NAND2_X1 U5136 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n6023) );
  NAND2_X1 U5137 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n6010) );
  NAND2_X1 U5138 ( .A1(INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4757) );
  NAND2_X1 U5139 ( .A1(n4222), .A2(n4221), .ZN(n4223) );
  INV_X1 U5140 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n4225) );
  XNOR2_X1 U5141 ( .A(n3704), .B(n4225), .ZN(n5616) );
  INV_X1 U5142 ( .A(n5616), .ZN(n4226) );
  INV_X1 U5143 ( .A(n4228), .ZN(n4227) );
  NAND3_X1 U5144 ( .A1(n4227), .A2(n4229), .A3(n5633), .ZN(n5681) );
  INV_X1 U5145 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5688) );
  INV_X1 U5146 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n4754) );
  NAND2_X1 U5147 ( .A1(n5688), .A2(n4754), .ZN(n4758) );
  INV_X1 U5148 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5673) );
  INV_X1 U5149 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n4229) );
  AND2_X1 U5150 ( .A1(INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5674) );
  INV_X1 U5151 ( .A(n5674), .ZN(n4243) );
  NOR3_X1 U5152 ( .A1(n5962), .A2(n4229), .A3(n4243), .ZN(n4230) );
  INV_X1 U5153 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5665) );
  OR2_X1 U5154 ( .A1(n4230), .A2(n5665), .ZN(n4232) );
  OAI21_X1 U5155 ( .B1(n5633), .B2(n5665), .A(INSTADDRPOINTER_REG_29__SCAN_IN), 
        .ZN(n4231) );
  NAND3_X1 U5156 ( .A1(n4233), .A2(n4232), .A3(n4231), .ZN(n4234) );
  INV_X1 U5157 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4329) );
  INV_X1 U5158 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5769) );
  NAND2_X1 U5159 ( .A1(n5576), .A2(n6498), .ZN(n4237) );
  NAND2_X1 U5160 ( .A1(n6523), .A2(REIP_REG_31__SCAN_IN), .ZN(n5648) );
  OAI211_X1 U5161 ( .C1(n5640), .C2(n4329), .A(n4237), .B(n5648), .ZN(n4238)
         );
  INV_X1 U5162 ( .A(n4238), .ZN(n4239) );
  OAI211_X1 U5163 ( .C1(n5768), .C2(n6476), .A(n4240), .B(n4239), .ZN(U2955)
         );
  NAND2_X1 U5164 ( .A1(n4244), .A2(n4242), .ZN(n4581) );
  NOR2_X2 U5165 ( .A1(n4581), .A2(n4243), .ZN(n5607) );
  NAND2_X1 U5166 ( .A1(n5667), .A2(n6496), .ZN(n4252) );
  NAND2_X1 U5167 ( .A1(n5605), .A2(n4247), .ZN(n5780) );
  INV_X1 U5168 ( .A(n5780), .ZN(n4250) );
  NAND2_X1 U5169 ( .A1(n6523), .A2(REIP_REG_29__SCAN_IN), .ZN(n5676) );
  NAND2_X1 U5170 ( .A1(n6491), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4248)
         );
  OAI211_X1 U5171 ( .C1(n5778), .C2(n6490), .A(n5676), .B(n4248), .ZN(n4249)
         );
  NAND2_X1 U5172 ( .A1(n4252), .A2(n4251), .ZN(n4580) );
  AOI22_X1 U5173 ( .A1(EAX_REG_10__SCAN_IN), .A2(keyinput147), .B1(
        INSTQUEUE_REG_13__4__SCAN_IN), .B2(keyinput164), .ZN(n4253) );
  OAI221_X1 U5174 ( .B1(EAX_REG_10__SCAN_IN), .B2(keyinput147), .C1(
        INSTQUEUE_REG_13__4__SCAN_IN), .C2(keyinput164), .A(n4253), .ZN(n4260)
         );
  AOI22_X1 U5175 ( .A1(BYTEENABLE_REG_0__SCAN_IN), .A2(keyinput233), .B1(
        ADDRESS_REG_25__SCAN_IN), .B2(keyinput230), .ZN(n4254) );
  OAI221_X1 U5176 ( .B1(BYTEENABLE_REG_0__SCAN_IN), .B2(keyinput233), .C1(
        ADDRESS_REG_25__SCAN_IN), .C2(keyinput230), .A(n4254), .ZN(n4259) );
  AOI22_X1 U5177 ( .A1(EBX_REG_17__SCAN_IN), .A2(keyinput232), .B1(
        INSTQUEUE_REG_9__4__SCAN_IN), .B2(keyinput205), .ZN(n4255) );
  OAI221_X1 U5178 ( .B1(EBX_REG_17__SCAN_IN), .B2(keyinput232), .C1(
        INSTQUEUE_REG_9__4__SCAN_IN), .C2(keyinput205), .A(n4255), .ZN(n4258)
         );
  AOI22_X1 U5179 ( .A1(LWORD_REG_1__SCAN_IN), .A2(keyinput201), .B1(
        INSTADDRPOINTER_REG_18__SCAN_IN), .B2(keyinput241), .ZN(n4256) );
  OAI221_X1 U5180 ( .B1(LWORD_REG_1__SCAN_IN), .B2(keyinput201), .C1(
        INSTADDRPOINTER_REG_18__SCAN_IN), .C2(keyinput241), .A(n4256), .ZN(
        n4257) );
  NOR4_X1 U5181 ( .A1(n4260), .A2(n4259), .A3(n4258), .A4(n4257), .ZN(n4288)
         );
  AOI22_X1 U5182 ( .A1(LWORD_REG_15__SCAN_IN), .A2(keyinput228), .B1(
        DATAO_REG_22__SCAN_IN), .B2(keyinput226), .ZN(n4261) );
  OAI221_X1 U5183 ( .B1(LWORD_REG_15__SCAN_IN), .B2(keyinput228), .C1(
        DATAO_REG_22__SCAN_IN), .C2(keyinput226), .A(n4261), .ZN(n4268) );
  AOI22_X1 U5184 ( .A1(REIP_REG_28__SCAN_IN), .A2(keyinput136), .B1(
        EAX_REG_7__SCAN_IN), .B2(keyinput133), .ZN(n4262) );
  OAI221_X1 U5185 ( .B1(REIP_REG_28__SCAN_IN), .B2(keyinput136), .C1(
        EAX_REG_7__SCAN_IN), .C2(keyinput133), .A(n4262), .ZN(n4267) );
  AOI22_X1 U5186 ( .A1(DATAI_9_), .A2(keyinput211), .B1(
        DATAWIDTH_REG_5__SCAN_IN), .B2(keyinput190), .ZN(n4263) );
  OAI221_X1 U5187 ( .B1(DATAI_9_), .B2(keyinput211), .C1(
        DATAWIDTH_REG_5__SCAN_IN), .C2(keyinput190), .A(n4263), .ZN(n4266) );
  AOI22_X1 U5188 ( .A1(PHYADDRPOINTER_REG_29__SCAN_IN), .A2(keyinput166), .B1(
        INSTQUEUE_REG_10__4__SCAN_IN), .B2(keyinput155), .ZN(n4264) );
  OAI221_X1 U5189 ( .B1(PHYADDRPOINTER_REG_29__SCAN_IN), .B2(keyinput166), 
        .C1(INSTQUEUE_REG_10__4__SCAN_IN), .C2(keyinput155), .A(n4264), .ZN(
        n4265) );
  NOR4_X1 U5190 ( .A1(n4268), .A2(n4267), .A3(n4266), .A4(n4265), .ZN(n4287)
         );
  AOI22_X1 U5191 ( .A1(DATAI_24_), .A2(keyinput252), .B1(
        INSTQUEUE_REG_15__0__SCAN_IN), .B2(keyinput134), .ZN(n4269) );
  OAI221_X1 U5192 ( .B1(DATAI_24_), .B2(keyinput252), .C1(
        INSTQUEUE_REG_15__0__SCAN_IN), .C2(keyinput134), .A(n4269), .ZN(n4276)
         );
  AOI22_X1 U5193 ( .A1(DATAI_26_), .A2(keyinput206), .B1(
        INSTQUEUE_REG_13__5__SCAN_IN), .B2(keyinput223), .ZN(n4270) );
  OAI221_X1 U5194 ( .B1(DATAI_26_), .B2(keyinput206), .C1(
        INSTQUEUE_REG_13__5__SCAN_IN), .C2(keyinput223), .A(n4270), .ZN(n4275)
         );
  AOI22_X1 U5195 ( .A1(ADDRESS_REG_18__SCAN_IN), .A2(keyinput188), .B1(
        INSTQUEUE_REG_3__2__SCAN_IN), .B2(keyinput239), .ZN(n4271) );
  OAI221_X1 U5196 ( .B1(ADDRESS_REG_18__SCAN_IN), .B2(keyinput188), .C1(
        INSTQUEUE_REG_3__2__SCAN_IN), .C2(keyinput239), .A(n4271), .ZN(n4274)
         );
  AOI22_X1 U5197 ( .A1(UWORD_REG_4__SCAN_IN), .A2(keyinput183), .B1(
        INSTQUEUE_REG_8__6__SCAN_IN), .B2(keyinput177), .ZN(n4272) );
  OAI221_X1 U5198 ( .B1(UWORD_REG_4__SCAN_IN), .B2(keyinput183), .C1(
        INSTQUEUE_REG_8__6__SCAN_IN), .C2(keyinput177), .A(n4272), .ZN(n4273)
         );
  NOR4_X1 U5199 ( .A1(n4276), .A2(n4275), .A3(n4274), .A4(n4273), .ZN(n4286)
         );
  AOI22_X1 U5200 ( .A1(INSTADDRPOINTER_REG_31__SCAN_IN), .A2(keyinput244), 
        .B1(EAX_REG_13__SCAN_IN), .B2(keyinput197), .ZN(n4277) );
  OAI221_X1 U5201 ( .B1(INSTADDRPOINTER_REG_31__SCAN_IN), .B2(keyinput244), 
        .C1(EAX_REG_13__SCAN_IN), .C2(keyinput197), .A(n4277), .ZN(n4284) );
  AOI22_X1 U5202 ( .A1(INSTADDRPOINTER_REG_8__SCAN_IN), .A2(keyinput231), .B1(
        INSTQUEUE_REG_0__2__SCAN_IN), .B2(keyinput254), .ZN(n4278) );
  OAI221_X1 U5203 ( .B1(INSTADDRPOINTER_REG_8__SCAN_IN), .B2(keyinput231), 
        .C1(INSTQUEUE_REG_0__2__SCAN_IN), .C2(keyinput254), .A(n4278), .ZN(
        n4283) );
  AOI22_X1 U5204 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(keyinput224), .B1(
        INSTQUEUE_REG_11__1__SCAN_IN), .B2(keyinput145), .ZN(n4279) );
  OAI221_X1 U5205 ( .B1(DATAWIDTH_REG_3__SCAN_IN), .B2(keyinput224), .C1(
        INSTQUEUE_REG_11__1__SCAN_IN), .C2(keyinput145), .A(n4279), .ZN(n4282)
         );
  AOI22_X1 U5206 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(keyinput234), .B1(
        INSTQUEUE_REG_1__6__SCAN_IN), .B2(keyinput200), .ZN(n4280) );
  OAI221_X1 U5207 ( .B1(DATAWIDTH_REG_19__SCAN_IN), .B2(keyinput234), .C1(
        INSTQUEUE_REG_1__6__SCAN_IN), .C2(keyinput200), .A(n4280), .ZN(n4281)
         );
  NOR4_X1 U5208 ( .A1(n4284), .A2(n4283), .A3(n4282), .A4(n4281), .ZN(n4285)
         );
  NAND4_X1 U5209 ( .A1(n4288), .A2(n4287), .A3(n4286), .A4(n4285), .ZN(n4411)
         );
  AOI22_X1 U5210 ( .A1(DATAO_REG_2__SCAN_IN), .A2(keyinput236), .B1(
        INSTADDRPOINTER_REG_3__SCAN_IN), .B2(keyinput214), .ZN(n4289) );
  OAI221_X1 U5211 ( .B1(DATAO_REG_2__SCAN_IN), .B2(keyinput236), .C1(
        INSTADDRPOINTER_REG_3__SCAN_IN), .C2(keyinput214), .A(n4289), .ZN(
        n4296) );
  AOI22_X1 U5212 ( .A1(ADDRESS_REG_15__SCAN_IN), .A2(keyinput168), .B1(
        DATAI_29_), .B2(keyinput250), .ZN(n4290) );
  OAI221_X1 U5213 ( .B1(ADDRESS_REG_15__SCAN_IN), .B2(keyinput168), .C1(
        DATAI_29_), .C2(keyinput250), .A(n4290), .ZN(n4295) );
  AOI22_X1 U5214 ( .A1(DATAO_REG_0__SCAN_IN), .A2(keyinput129), .B1(
        PHYADDRPOINTER_REG_12__SCAN_IN), .B2(keyinput237), .ZN(n4291) );
  OAI221_X1 U5215 ( .B1(DATAO_REG_0__SCAN_IN), .B2(keyinput129), .C1(
        PHYADDRPOINTER_REG_12__SCAN_IN), .C2(keyinput237), .A(n4291), .ZN(
        n4294) );
  AOI22_X1 U5216 ( .A1(ADS_N_REG_SCAN_IN), .A2(keyinput159), .B1(
        REIP_REG_12__SCAN_IN), .B2(keyinput135), .ZN(n4292) );
  OAI221_X1 U5217 ( .B1(ADS_N_REG_SCAN_IN), .B2(keyinput159), .C1(
        REIP_REG_12__SCAN_IN), .C2(keyinput135), .A(n4292), .ZN(n4293) );
  NOR4_X1 U5218 ( .A1(n4296), .A2(n4295), .A3(n4294), .A4(n4293), .ZN(n4324)
         );
  AOI22_X1 U5219 ( .A1(ADDRESS_REG_29__SCAN_IN), .A2(keyinput209), .B1(
        INSTQUEUE_REG_2__2__SCAN_IN), .B2(keyinput160), .ZN(n4297) );
  OAI221_X1 U5220 ( .B1(ADDRESS_REG_29__SCAN_IN), .B2(keyinput209), .C1(
        INSTQUEUE_REG_2__2__SCAN_IN), .C2(keyinput160), .A(n4297), .ZN(n4304)
         );
  AOI22_X1 U5221 ( .A1(DATAI_25_), .A2(keyinput215), .B1(EAX_REG_2__SCAN_IN), 
        .B2(keyinput179), .ZN(n4298) );
  OAI221_X1 U5222 ( .B1(DATAI_25_), .B2(keyinput215), .C1(EAX_REG_2__SCAN_IN), 
        .C2(keyinput179), .A(n4298), .ZN(n4303) );
  AOI22_X1 U5223 ( .A1(REIP_REG_9__SCAN_IN), .A2(keyinput151), .B1(
        DATAWIDTH_REG_29__SCAN_IN), .B2(keyinput235), .ZN(n4299) );
  OAI221_X1 U5224 ( .B1(REIP_REG_9__SCAN_IN), .B2(keyinput151), .C1(
        DATAWIDTH_REG_29__SCAN_IN), .C2(keyinput235), .A(n4299), .ZN(n4302) );
  AOI22_X1 U5225 ( .A1(BE_N_REG_1__SCAN_IN), .A2(keyinput240), .B1(
        DATAWIDTH_REG_0__SCAN_IN), .B2(keyinput181), .ZN(n4300) );
  OAI221_X1 U5226 ( .B1(BE_N_REG_1__SCAN_IN), .B2(keyinput240), .C1(
        DATAWIDTH_REG_0__SCAN_IN), .C2(keyinput181), .A(n4300), .ZN(n4301) );
  NOR4_X1 U5227 ( .A1(n4304), .A2(n4303), .A3(n4302), .A4(n4301), .ZN(n4323)
         );
  AOI22_X1 U5228 ( .A1(DATAI_6_), .A2(keyinput149), .B1(DATAO_REG_15__SCAN_IN), 
        .B2(keyinput218), .ZN(n4305) );
  OAI221_X1 U5229 ( .B1(DATAI_6_), .B2(keyinput149), .C1(DATAO_REG_15__SCAN_IN), .C2(keyinput218), .A(n4305), .ZN(n4312) );
  AOI22_X1 U5230 ( .A1(UWORD_REG_10__SCAN_IN), .A2(keyinput163), .B1(
        INSTQUEUE_REG_1__2__SCAN_IN), .B2(keyinput225), .ZN(n4306) );
  OAI221_X1 U5231 ( .B1(UWORD_REG_10__SCAN_IN), .B2(keyinput163), .C1(
        INSTQUEUE_REG_1__2__SCAN_IN), .C2(keyinput225), .A(n4306), .ZN(n4311)
         );
  AOI22_X1 U5232 ( .A1(PHYADDRPOINTER_REG_11__SCAN_IN), .A2(keyinput175), .B1(
        INSTADDRPOINTER_REG_9__SCAN_IN), .B2(keyinput192), .ZN(n4307) );
  OAI221_X1 U5233 ( .B1(PHYADDRPOINTER_REG_11__SCAN_IN), .B2(keyinput175), 
        .C1(INSTADDRPOINTER_REG_9__SCAN_IN), .C2(keyinput192), .A(n4307), .ZN(
        n4310) );
  AOI22_X1 U5234 ( .A1(INSTQUEUE_REG_5__1__SCAN_IN), .A2(keyinput140), .B1(
        INSTQUEUE_REG_12__2__SCAN_IN), .B2(keyinput178), .ZN(n4308) );
  OAI221_X1 U5235 ( .B1(INSTQUEUE_REG_5__1__SCAN_IN), .B2(keyinput140), .C1(
        INSTQUEUE_REG_12__2__SCAN_IN), .C2(keyinput178), .A(n4308), .ZN(n4309)
         );
  NOR4_X1 U5236 ( .A1(n4312), .A2(n4311), .A3(n4310), .A4(n4309), .ZN(n4322)
         );
  AOI22_X1 U5237 ( .A1(BE_N_REG_3__SCAN_IN), .A2(keyinput162), .B1(DATAI_30_), 
        .B2(keyinput167), .ZN(n4313) );
  OAI221_X1 U5238 ( .B1(BE_N_REG_3__SCAN_IN), .B2(keyinput162), .C1(DATAI_30_), 
        .C2(keyinput167), .A(n4313), .ZN(n4320) );
  AOI22_X1 U5239 ( .A1(DATAO_REG_1__SCAN_IN), .A2(keyinput161), .B1(
        INSTQUEUE_REG_15__7__SCAN_IN), .B2(keyinput138), .ZN(n4314) );
  OAI221_X1 U5240 ( .B1(DATAO_REG_1__SCAN_IN), .B2(keyinput161), .C1(
        INSTQUEUE_REG_15__7__SCAN_IN), .C2(keyinput138), .A(n4314), .ZN(n4319)
         );
  AOI22_X1 U5241 ( .A1(REIP_REG_18__SCAN_IN), .A2(keyinput246), .B1(
        INSTQUEUE_REG_9__1__SCAN_IN), .B2(keyinput189), .ZN(n4315) );
  OAI221_X1 U5242 ( .B1(REIP_REG_18__SCAN_IN), .B2(keyinput246), .C1(
        INSTQUEUE_REG_9__1__SCAN_IN), .C2(keyinput189), .A(n4315), .ZN(n4318)
         );
  AOI22_X1 U5243 ( .A1(EBX_REG_8__SCAN_IN), .A2(keyinput165), .B1(
        INSTQUEUE_REG_3__0__SCAN_IN), .B2(keyinput142), .ZN(n4316) );
  OAI221_X1 U5244 ( .B1(EBX_REG_8__SCAN_IN), .B2(keyinput165), .C1(
        INSTQUEUE_REG_3__0__SCAN_IN), .C2(keyinput142), .A(n4316), .ZN(n4317)
         );
  NOR4_X1 U5245 ( .A1(n4320), .A2(n4319), .A3(n4318), .A4(n4317), .ZN(n4321)
         );
  NAND4_X1 U5246 ( .A1(n4324), .A2(n4323), .A3(n4322), .A4(n4321), .ZN(n4410)
         );
  AOI22_X1 U5247 ( .A1(EBX_REG_14__SCAN_IN), .A2(keyinput251), .B1(
        INSTADDRPOINTER_REG_5__SCAN_IN), .B2(keyinput139), .ZN(n4325) );
  OAI221_X1 U5248 ( .B1(EBX_REG_14__SCAN_IN), .B2(keyinput251), .C1(
        INSTADDRPOINTER_REG_5__SCAN_IN), .C2(keyinput139), .A(n4325), .ZN(
        n4334) );
  INV_X1 U5249 ( .A(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n4551) );
  INV_X1 U5250 ( .A(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n4327) );
  AOI22_X1 U5251 ( .A1(n4551), .A2(keyinput182), .B1(n4327), .B2(keyinput153), 
        .ZN(n4326) );
  OAI221_X1 U5252 ( .B1(n4551), .B2(keyinput182), .C1(n4327), .C2(keyinput153), 
        .A(n4326), .ZN(n4333) );
  INV_X1 U5253 ( .A(EAX_REG_14__SCAN_IN), .ZN(n6402) );
  AOI22_X1 U5254 ( .A1(n4329), .A2(keyinput208), .B1(n6402), .B2(keyinput158), 
        .ZN(n4328) );
  OAI221_X1 U5255 ( .B1(n4329), .B2(keyinput208), .C1(n6402), .C2(keyinput158), 
        .A(n4328), .ZN(n4332) );
  INV_X1 U5256 ( .A(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n6755) );
  AOI22_X1 U5257 ( .A1(n6070), .A2(keyinput154), .B1(n6755), .B2(keyinput247), 
        .ZN(n4330) );
  OAI221_X1 U5258 ( .B1(n6070), .B2(keyinput154), .C1(n6755), .C2(keyinput247), 
        .A(n4330), .ZN(n4331) );
  NOR4_X1 U5259 ( .A1(n4334), .A2(n4333), .A3(n4332), .A4(n4331), .ZN(n4365)
         );
  INV_X1 U5260 ( .A(DATAO_REG_18__SCAN_IN), .ZN(n6392) );
  INV_X1 U5261 ( .A(ADDRESS_REG_17__SCAN_IN), .ZN(n6959) );
  AOI22_X1 U5262 ( .A1(n6392), .A2(keyinput227), .B1(keyinput185), .B2(n6959), 
        .ZN(n4335) );
  OAI221_X1 U5263 ( .B1(n6392), .B2(keyinput227), .C1(n6959), .C2(keyinput185), 
        .A(n4335), .ZN(n4343) );
  INV_X1 U5264 ( .A(DATAI_16_), .ZN(n5236) );
  AOI22_X1 U5265 ( .A1(n6164), .A2(keyinput216), .B1(keyinput171), .B2(n5236), 
        .ZN(n4336) );
  OAI221_X1 U5266 ( .B1(n6164), .B2(keyinput216), .C1(n5236), .C2(keyinput171), 
        .A(n4336), .ZN(n4342) );
  INV_X1 U5267 ( .A(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n4517) );
  AOI22_X1 U5268 ( .A1(n4517), .A2(keyinput203), .B1(keyinput213), .B2(n5665), 
        .ZN(n4337) );
  OAI221_X1 U5269 ( .B1(n4517), .B2(keyinput203), .C1(n5665), .C2(keyinput213), 
        .A(n4337), .ZN(n4341) );
  INV_X1 U5270 ( .A(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n6735) );
  XOR2_X1 U5271 ( .A(n6735), .B(keyinput217), .Z(n4339) );
  XNOR2_X1 U5272 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B(keyinput242), .ZN(
        n4338) );
  NAND2_X1 U5273 ( .A1(n4339), .A2(n4338), .ZN(n4340) );
  NOR4_X1 U5274 ( .A1(n4343), .A2(n4342), .A3(n4341), .A4(n4340), .ZN(n4364)
         );
  INV_X1 U5275 ( .A(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4345) );
  INV_X1 U5276 ( .A(ADDRESS_REG_27__SCAN_IN), .ZN(n6977) );
  AOI22_X1 U5277 ( .A1(n4345), .A2(keyinput191), .B1(keyinput148), .B2(n6977), 
        .ZN(n4344) );
  OAI221_X1 U5278 ( .B1(n4345), .B2(keyinput191), .C1(n6977), .C2(keyinput148), 
        .A(n4344), .ZN(n4352) );
  INV_X1 U5279 ( .A(EBX_REG_20__SCAN_IN), .ZN(n5922) );
  INV_X1 U5280 ( .A(EBX_REG_12__SCAN_IN), .ZN(n6296) );
  AOI22_X1 U5281 ( .A1(n5922), .A2(keyinput229), .B1(keyinput255), .B2(n6296), 
        .ZN(n4346) );
  OAI221_X1 U5282 ( .B1(n5922), .B2(keyinput229), .C1(n6296), .C2(keyinput255), 
        .A(n4346), .ZN(n4351) );
  INV_X1 U5283 ( .A(DATAO_REG_8__SCAN_IN), .ZN(n6416) );
  INV_X1 U5284 ( .A(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n4555) );
  AOI22_X1 U5285 ( .A1(n6416), .A2(keyinput176), .B1(n4555), .B2(keyinput198), 
        .ZN(n4347) );
  OAI221_X1 U5286 ( .B1(n6416), .B2(keyinput176), .C1(n4555), .C2(keyinput198), 
        .A(n4347), .ZN(n4350) );
  INV_X1 U5287 ( .A(ADDRESS_REG_23__SCAN_IN), .ZN(n6969) );
  INV_X1 U5288 ( .A(DATAO_REG_24__SCAN_IN), .ZN(n6382) );
  AOI22_X1 U5289 ( .A1(n6969), .A2(keyinput131), .B1(keyinput222), .B2(n6382), 
        .ZN(n4348) );
  OAI221_X1 U5290 ( .B1(n6969), .B2(keyinput131), .C1(n6382), .C2(keyinput222), 
        .A(n4348), .ZN(n4349) );
  NOR4_X1 U5291 ( .A1(n4352), .A2(n4351), .A3(n4350), .A4(n4349), .ZN(n4363)
         );
  INV_X1 U5292 ( .A(UWORD_REG_2__SCAN_IN), .ZN(n6442) );
  INV_X1 U5293 ( .A(DATAO_REG_12__SCAN_IN), .ZN(n6405) );
  AOI22_X1 U5294 ( .A1(n6442), .A2(keyinput202), .B1(keyinput170), .B2(n6405), 
        .ZN(n4353) );
  OAI221_X1 U5295 ( .B1(n6442), .B2(keyinput202), .C1(n6405), .C2(keyinput170), 
        .A(n4353), .ZN(n4361) );
  INV_X1 U5296 ( .A(EBX_REG_16__SCAN_IN), .ZN(n6284) );
  INV_X1 U5297 ( .A(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4355) );
  AOI22_X1 U5298 ( .A1(n6284), .A2(keyinput132), .B1(n4355), .B2(keyinput130), 
        .ZN(n4354) );
  OAI221_X1 U5299 ( .B1(n6284), .B2(keyinput132), .C1(n4355), .C2(keyinput130), 
        .A(n4354), .ZN(n4360) );
  AOI22_X1 U5300 ( .A1(n6118), .A2(keyinput137), .B1(n6128), .B2(keyinput212), 
        .ZN(n4356) );
  OAI221_X1 U5301 ( .B1(n6118), .B2(keyinput137), .C1(n6128), .C2(keyinput212), 
        .A(n4356), .ZN(n4359) );
  INV_X1 U5302 ( .A(REIP_REG_24__SCAN_IN), .ZN(n6968) );
  INV_X1 U5303 ( .A(EAX_REG_5__SCAN_IN), .ZN(n6423) );
  AOI22_X1 U5304 ( .A1(n6968), .A2(keyinput146), .B1(n6423), .B2(keyinput173), 
        .ZN(n4357) );
  OAI221_X1 U5305 ( .B1(n6968), .B2(keyinput146), .C1(n6423), .C2(keyinput173), 
        .A(n4357), .ZN(n4358) );
  NOR4_X1 U5306 ( .A1(n4361), .A2(n4360), .A3(n4359), .A4(n4358), .ZN(n4362)
         );
  NAND4_X1 U5307 ( .A1(n4365), .A2(n4364), .A3(n4363), .A4(n4362), .ZN(n4409)
         );
  INV_X1 U5308 ( .A(DATAI_15_), .ZN(n6339) );
  INV_X1 U5309 ( .A(DATAWIDTH_REG_31__SCAN_IN), .ZN(n6909) );
  AOI22_X1 U5310 ( .A1(n6339), .A2(keyinput150), .B1(keyinput194), .B2(n6909), 
        .ZN(n4366) );
  OAI221_X1 U5311 ( .B1(n6339), .B2(keyinput150), .C1(n6909), .C2(keyinput194), 
        .A(n4366), .ZN(n4374) );
  INV_X1 U5312 ( .A(UWORD_REG_1__SCAN_IN), .ZN(n6440) );
  INV_X1 U5313 ( .A(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n4565) );
  AOI22_X1 U5314 ( .A1(n6440), .A2(keyinput143), .B1(n4565), .B2(keyinput253), 
        .ZN(n4367) );
  OAI221_X1 U5315 ( .B1(n6440), .B2(keyinput143), .C1(n4565), .C2(keyinput253), 
        .A(n4367), .ZN(n4373) );
  INV_X1 U5316 ( .A(DATAO_REG_28__SCAN_IN), .ZN(n6375) );
  AOI22_X1 U5317 ( .A1(n6375), .A2(keyinput220), .B1(n5673), .B2(keyinput207), 
        .ZN(n4368) );
  OAI221_X1 U5318 ( .B1(n6375), .B2(keyinput220), .C1(n5673), .C2(keyinput207), 
        .A(n4368), .ZN(n4372) );
  INV_X1 U5319 ( .A(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4563) );
  XOR2_X1 U5320 ( .A(n4563), .B(keyinput196), .Z(n4370) );
  XNOR2_X1 U5321 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(keyinput128), .ZN(
        n4369) );
  NAND2_X1 U5322 ( .A1(n4370), .A2(n4369), .ZN(n4371) );
  NOR4_X1 U5323 ( .A1(n4374), .A2(n4373), .A3(n4372), .A4(n4371), .ZN(n4407)
         );
  INV_X1 U5324 ( .A(LWORD_REG_10__SCAN_IN), .ZN(n6459) );
  INV_X1 U5325 ( .A(BE_N_REG_0__SCAN_IN), .ZN(n6991) );
  AOI22_X1 U5326 ( .A1(n6459), .A2(keyinput187), .B1(keyinput152), .B2(n6991), 
        .ZN(n4375) );
  OAI221_X1 U5327 ( .B1(n6459), .B2(keyinput187), .C1(n6991), .C2(keyinput152), 
        .A(n4375), .ZN(n4384) );
  INV_X1 U5328 ( .A(LWORD_REG_11__SCAN_IN), .ZN(n6462) );
  INV_X1 U5329 ( .A(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n4569) );
  AOI22_X1 U5330 ( .A1(n6462), .A2(keyinput193), .B1(n4569), .B2(keyinput180), 
        .ZN(n4376) );
  OAI221_X1 U5331 ( .B1(n6462), .B2(keyinput193), .C1(n4569), .C2(keyinput180), 
        .A(n4376), .ZN(n4383) );
  INV_X1 U5332 ( .A(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n6202) );
  INV_X1 U5333 ( .A(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n4378) );
  AOI22_X1 U5334 ( .A1(n6202), .A2(keyinput195), .B1(n4378), .B2(keyinput248), 
        .ZN(n4377) );
  OAI221_X1 U5335 ( .B1(n6202), .B2(keyinput195), .C1(n4378), .C2(keyinput248), 
        .A(n4377), .ZN(n4382) );
  INV_X1 U5336 ( .A(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4457) );
  XOR2_X1 U5337 ( .A(n4457), .B(keyinput144), .Z(n4380) );
  XNOR2_X1 U5338 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(keyinput210), .ZN(
        n4379) );
  NAND2_X1 U5339 ( .A1(n4380), .A2(n4379), .ZN(n4381) );
  NOR4_X1 U5340 ( .A1(n4384), .A2(n4383), .A3(n4382), .A4(n4381), .ZN(n4406)
         );
  INV_X1 U5341 ( .A(REIP_REG_8__SCAN_IN), .ZN(n6941) );
  INV_X1 U5342 ( .A(ADDRESS_REG_5__SCAN_IN), .ZN(n6937) );
  AOI22_X1 U5343 ( .A1(n6941), .A2(keyinput141), .B1(keyinput172), .B2(n6937), 
        .ZN(n4385) );
  OAI221_X1 U5344 ( .B1(n6941), .B2(keyinput141), .C1(n6937), .C2(keyinput172), 
        .A(n4385), .ZN(n4393) );
  INV_X1 U5345 ( .A(ADDRESS_REG_3__SCAN_IN), .ZN(n6932) );
  INV_X1 U5346 ( .A(REIP_REG_31__SCAN_IN), .ZN(n6983) );
  AOI22_X1 U5347 ( .A1(n6932), .A2(keyinput199), .B1(keyinput238), .B2(n6983), 
        .ZN(n4386) );
  OAI221_X1 U5348 ( .B1(n6932), .B2(keyinput199), .C1(n6983), .C2(keyinput238), 
        .A(n4386), .ZN(n4392) );
  INV_X1 U5349 ( .A(EBX_REG_24__SCAN_IN), .ZN(n5913) );
  AOI22_X1 U5350 ( .A1(n6073), .A2(keyinput249), .B1(keyinput156), .B2(n5913), 
        .ZN(n4387) );
  OAI221_X1 U5351 ( .B1(n6073), .B2(keyinput249), .C1(n5913), .C2(keyinput156), 
        .A(n4387), .ZN(n4391) );
  INV_X1 U5352 ( .A(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n4528) );
  AOI22_X1 U5353 ( .A1(n4389), .A2(keyinput184), .B1(n4528), .B2(keyinput221), 
        .ZN(n4388) );
  OAI221_X1 U5354 ( .B1(n4389), .B2(keyinput184), .C1(n4528), .C2(keyinput221), 
        .A(n4388), .ZN(n4390) );
  NOR4_X1 U5355 ( .A1(n4393), .A2(n4392), .A3(n4391), .A4(n4390), .ZN(n4405)
         );
  INV_X1 U5356 ( .A(DATAI_2_), .ZN(n5276) );
  INV_X1 U5357 ( .A(REIP_REG_3__SCAN_IN), .ZN(n6931) );
  AOI22_X1 U5358 ( .A1(n5276), .A2(keyinput169), .B1(keyinput174), .B2(n6931), 
        .ZN(n4394) );
  OAI221_X1 U5359 ( .B1(n5276), .B2(keyinput169), .C1(n6931), .C2(keyinput174), 
        .A(n4394), .ZN(n4403) );
  INV_X1 U5360 ( .A(LWORD_REG_12__SCAN_IN), .ZN(n6407) );
  AOI22_X1 U5361 ( .A1(n6407), .A2(keyinput186), .B1(n4568), .B2(keyinput219), 
        .ZN(n4395) );
  OAI221_X1 U5362 ( .B1(n6407), .B2(keyinput186), .C1(n4568), .C2(keyinput219), 
        .A(n4395), .ZN(n4402) );
  INV_X1 U5363 ( .A(ADDRESS_REG_13__SCAN_IN), .ZN(n6952) );
  AOI22_X1 U5364 ( .A1(n5688), .A2(keyinput245), .B1(keyinput243), .B2(n6952), 
        .ZN(n4396) );
  OAI221_X1 U5365 ( .B1(n5688), .B2(keyinput245), .C1(n6952), .C2(keyinput243), 
        .A(n4396), .ZN(n4401) );
  INV_X1 U5366 ( .A(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n4399) );
  INV_X1 U5367 ( .A(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n4398) );
  AOI22_X1 U5368 ( .A1(n4399), .A2(keyinput204), .B1(n4398), .B2(keyinput157), 
        .ZN(n4397) );
  OAI221_X1 U5369 ( .B1(n4399), .B2(keyinput204), .C1(n4398), .C2(keyinput157), 
        .A(n4397), .ZN(n4400) );
  NOR4_X1 U5370 ( .A1(n4403), .A2(n4402), .A3(n4401), .A4(n4400), .ZN(n4404)
         );
  NAND4_X1 U5371 ( .A1(n4407), .A2(n4406), .A3(n4405), .A4(n4404), .ZN(n4408)
         );
  NOR4_X1 U5372 ( .A1(n4411), .A2(n4410), .A3(n4409), .A4(n4408), .ZN(n4579)
         );
  OAI22_X1 U5373 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(keyinput0), .B1(
        DATAO_REG_22__SCAN_IN), .B2(keyinput98), .ZN(n4412) );
  AOI221_X1 U5374 ( .B1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(keyinput0), .C1(
        keyinput98), .C2(DATAO_REG_22__SCAN_IN), .A(n4412), .ZN(n4419) );
  OAI22_X1 U5375 ( .A1(PHYADDRPOINTER_REG_29__SCAN_IN), .A2(keyinput38), .B1(
        keyinput107), .B2(DATAWIDTH_REG_29__SCAN_IN), .ZN(n4413) );
  AOI221_X1 U5376 ( .B1(PHYADDRPOINTER_REG_29__SCAN_IN), .B2(keyinput38), .C1(
        DATAWIDTH_REG_29__SCAN_IN), .C2(keyinput107), .A(n4413), .ZN(n4418) );
  OAI22_X1 U5377 ( .A1(EAX_REG_7__SCAN_IN), .A2(keyinput5), .B1(keyinput81), 
        .B2(ADDRESS_REG_29__SCAN_IN), .ZN(n4414) );
  AOI221_X1 U5378 ( .B1(EAX_REG_7__SCAN_IN), .B2(keyinput5), .C1(
        ADDRESS_REG_29__SCAN_IN), .C2(keyinput81), .A(n4414), .ZN(n4417) );
  OAI22_X1 U5379 ( .A1(DATAI_6_), .A2(keyinput21), .B1(keyinput28), .B2(
        EBX_REG_24__SCAN_IN), .ZN(n4415) );
  AOI221_X1 U5380 ( .B1(DATAI_6_), .B2(keyinput21), .C1(EBX_REG_24__SCAN_IN), 
        .C2(keyinput28), .A(n4415), .ZN(n4416) );
  NAND4_X1 U5381 ( .A1(n4419), .A2(n4418), .A3(n4417), .A4(n4416), .ZN(n4447)
         );
  OAI22_X1 U5382 ( .A1(INSTADDRPOINTER_REG_31__SCAN_IN), .A2(keyinput116), 
        .B1(DATAWIDTH_REG_0__SCAN_IN), .B2(keyinput53), .ZN(n4420) );
  AOI221_X1 U5383 ( .B1(INSTADDRPOINTER_REG_31__SCAN_IN), .B2(keyinput116), 
        .C1(keyinput53), .C2(DATAWIDTH_REG_0__SCAN_IN), .A(n4420), .ZN(n4427)
         );
  OAI22_X1 U5384 ( .A1(PHYADDRPOINTER_REG_9__SCAN_IN), .A2(keyinput88), .B1(
        DATAO_REG_0__SCAN_IN), .B2(keyinput1), .ZN(n4421) );
  AOI221_X1 U5385 ( .B1(PHYADDRPOINTER_REG_9__SCAN_IN), .B2(keyinput88), .C1(
        keyinput1), .C2(DATAO_REG_0__SCAN_IN), .A(n4421), .ZN(n4426) );
  OAI22_X1 U5386 ( .A1(DATAO_REG_1__SCAN_IN), .A2(keyinput33), .B1(keyinput80), 
        .B2(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4422) );
  AOI221_X1 U5387 ( .B1(DATAO_REG_1__SCAN_IN), .B2(keyinput33), .C1(
        PHYADDRPOINTER_REG_31__SCAN_IN), .C2(keyinput80), .A(n4422), .ZN(n4425) );
  OAI22_X1 U5388 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(keyinput61), .B1(
        keyinput65), .B2(LWORD_REG_11__SCAN_IN), .ZN(n4423) );
  AOI221_X1 U5389 ( .B1(INSTQUEUE_REG_9__1__SCAN_IN), .B2(keyinput61), .C1(
        LWORD_REG_11__SCAN_IN), .C2(keyinput65), .A(n4423), .ZN(n4424) );
  NAND4_X1 U5390 ( .A1(n4427), .A2(n4426), .A3(n4425), .A4(n4424), .ZN(n4446)
         );
  OAI22_X1 U5391 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(keyinput82), .B1(
        keyinput31), .B2(ADS_N_REG_SCAN_IN), .ZN(n4428) );
  AOI221_X1 U5392 ( .B1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(keyinput82), 
        .C1(ADS_N_REG_SCAN_IN), .C2(keyinput31), .A(n4428), .ZN(n4435) );
  OAI22_X1 U5393 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(keyinput113), 
        .B1(DATAO_REG_8__SCAN_IN), .B2(keyinput48), .ZN(n4429) );
  AOI221_X1 U5394 ( .B1(INSTADDRPOINTER_REG_18__SCAN_IN), .B2(keyinput113), 
        .C1(keyinput48), .C2(DATAO_REG_8__SCAN_IN), .A(n4429), .ZN(n4434) );
  OAI22_X1 U5395 ( .A1(INSTQUEUE_REG_12__0__SCAN_IN), .A2(keyinput89), .B1(
        keyinput109), .B2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n4430) );
  AOI221_X1 U5396 ( .B1(INSTQUEUE_REG_12__0__SCAN_IN), .B2(keyinput89), .C1(
        PHYADDRPOINTER_REG_12__SCAN_IN), .C2(keyinput109), .A(n4430), .ZN(
        n4433) );
  OAI22_X1 U5397 ( .A1(DATAI_29_), .A2(keyinput122), .B1(
        ADDRESS_REG_3__SCAN_IN), .B2(keyinput71), .ZN(n4431) );
  AOI221_X1 U5398 ( .B1(DATAI_29_), .B2(keyinput122), .C1(keyinput71), .C2(
        ADDRESS_REG_3__SCAN_IN), .A(n4431), .ZN(n4432) );
  NAND4_X1 U5399 ( .A1(n4435), .A2(n4434), .A3(n4433), .A4(n4432), .ZN(n4445)
         );
  OAI22_X1 U5400 ( .A1(INSTQUEUE_REG_10__4__SCAN_IN), .A2(keyinput27), .B1(
        DATAI_9_), .B2(keyinput83), .ZN(n4436) );
  AOI221_X1 U5401 ( .B1(INSTQUEUE_REG_10__4__SCAN_IN), .B2(keyinput27), .C1(
        keyinput83), .C2(DATAI_9_), .A(n4436), .ZN(n4443) );
  OAI22_X1 U5402 ( .A1(INSTQUEUE_REG_8__1__SCAN_IN), .A2(keyinput76), .B1(
        INSTADDRPOINTER_REG_27__SCAN_IN), .B2(keyinput117), .ZN(n4437) );
  AOI221_X1 U5403 ( .B1(INSTQUEUE_REG_8__1__SCAN_IN), .B2(keyinput76), .C1(
        keyinput117), .C2(INSTADDRPOINTER_REG_27__SCAN_IN), .A(n4437), .ZN(
        n4442) );
  OAI22_X1 U5404 ( .A1(PHYADDRPOINTER_REG_13__SCAN_IN), .A2(keyinput84), .B1(
        keyinput56), .B2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n4438) );
  AOI221_X1 U5405 ( .B1(PHYADDRPOINTER_REG_13__SCAN_IN), .B2(keyinput84), .C1(
        PHYADDRPOINTER_REG_25__SCAN_IN), .C2(keyinput56), .A(n4438), .ZN(n4441) );
  OAI22_X1 U5406 ( .A1(INSTQUEUE_REG_6__7__SCAN_IN), .A2(keyinput2), .B1(
        INSTADDRPOINTER_REG_9__SCAN_IN), .B2(keyinput64), .ZN(n4439) );
  AOI221_X1 U5407 ( .B1(INSTQUEUE_REG_6__7__SCAN_IN), .B2(keyinput2), .C1(
        keyinput64), .C2(INSTADDRPOINTER_REG_9__SCAN_IN), .A(n4439), .ZN(n4440) );
  NAND4_X1 U5408 ( .A1(n4443), .A2(n4442), .A3(n4441), .A4(n4440), .ZN(n4444)
         );
  NOR4_X1 U5409 ( .A1(n4447), .A2(n4446), .A3(n4445), .A4(n4444), .ZN(n4496)
         );
  OAI22_X1 U5410 ( .A1(INSTQUEUE_REG_13__5__SCAN_IN), .A2(keyinput95), .B1(
        BE_N_REG_3__SCAN_IN), .B2(keyinput34), .ZN(n4448) );
  AOI221_X1 U5411 ( .B1(INSTQUEUE_REG_13__5__SCAN_IN), .B2(keyinput95), .C1(
        keyinput34), .C2(BE_N_REG_3__SCAN_IN), .A(n4448), .ZN(n4455) );
  OAI22_X1 U5412 ( .A1(DATAO_REG_24__SCAN_IN), .A2(keyinput94), .B1(keyinput59), .B2(LWORD_REG_10__SCAN_IN), .ZN(n4449) );
  AOI221_X1 U5413 ( .B1(DATAO_REG_24__SCAN_IN), .B2(keyinput94), .C1(
        LWORD_REG_10__SCAN_IN), .C2(keyinput59), .A(n4449), .ZN(n4454) );
  OAI22_X1 U5414 ( .A1(EAX_REG_10__SCAN_IN), .A2(keyinput19), .B1(
        EBX_REG_16__SCAN_IN), .B2(keyinput4), .ZN(n4450) );
  AOI221_X1 U5415 ( .B1(EAX_REG_10__SCAN_IN), .B2(keyinput19), .C1(keyinput4), 
        .C2(EBX_REG_16__SCAN_IN), .A(n4450), .ZN(n4453) );
  OAI22_X1 U5416 ( .A1(INSTQUEUE_REG_2__4__SCAN_IN), .A2(keyinput63), .B1(
        keyinput50), .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n4451) );
  AOI221_X1 U5417 ( .B1(INSTQUEUE_REG_2__4__SCAN_IN), .B2(keyinput63), .C1(
        INSTQUEUE_REG_12__2__SCAN_IN), .C2(keyinput50), .A(n4451), .ZN(n4452)
         );
  NAND4_X1 U5418 ( .A1(n4455), .A2(n4454), .A3(n4453), .A4(n4452), .ZN(n4461)
         );
  INV_X1 U5419 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4953) );
  AOI22_X1 U5420 ( .A1(n4953), .A2(keyinput86), .B1(n4457), .B2(keyinput16), 
        .ZN(n4456) );
  OAI221_X1 U5421 ( .B1(n4953), .B2(keyinput86), .C1(n4457), .C2(keyinput16), 
        .A(n4456), .ZN(n4460) );
  XNOR2_X1 U5422 ( .A(n3289), .B(keyinput114), .ZN(n4459) );
  INV_X1 U5423 ( .A(DATAWIDTH_REG_5__SCAN_IN), .ZN(n6910) );
  XNOR2_X1 U5424 ( .A(n6910), .B(keyinput62), .ZN(n4458) );
  NOR4_X1 U5425 ( .A1(n4461), .A2(n4460), .A3(n4459), .A4(n4458), .ZN(n4495)
         );
  OAI22_X1 U5426 ( .A1(EBX_REG_12__SCAN_IN), .A2(keyinput127), .B1(keyinput58), 
        .B2(LWORD_REG_12__SCAN_IN), .ZN(n4462) );
  AOI221_X1 U5427 ( .B1(EBX_REG_12__SCAN_IN), .B2(keyinput127), .C1(
        LWORD_REG_12__SCAN_IN), .C2(keyinput58), .A(n4462), .ZN(n4469) );
  OAI22_X1 U5428 ( .A1(DATAI_24_), .A2(keyinput124), .B1(
        ADDRESS_REG_17__SCAN_IN), .B2(keyinput57), .ZN(n4463) );
  AOI221_X1 U5429 ( .B1(DATAI_24_), .B2(keyinput124), .C1(keyinput57), .C2(
        ADDRESS_REG_17__SCAN_IN), .A(n4463), .ZN(n4468) );
  OAI22_X1 U5430 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(keyinput106), .B1(
        keyinput24), .B2(BE_N_REG_0__SCAN_IN), .ZN(n4464) );
  AOI221_X1 U5431 ( .B1(DATAWIDTH_REG_19__SCAN_IN), .B2(keyinput106), .C1(
        BE_N_REG_0__SCAN_IN), .C2(keyinput24), .A(n4464), .ZN(n4467) );
  OAI22_X1 U5432 ( .A1(INSTQUEUE_REG_15__7__SCAN_IN), .A2(keyinput10), .B1(
        PHYADDRPOINTER_REG_5__SCAN_IN), .B2(keyinput67), .ZN(n4465) );
  AOI221_X1 U5433 ( .B1(INSTQUEUE_REG_15__7__SCAN_IN), .B2(keyinput10), .C1(
        keyinput67), .C2(PHYADDRPOINTER_REG_5__SCAN_IN), .A(n4465), .ZN(n4466)
         );
  NAND4_X1 U5434 ( .A1(n4469), .A2(n4468), .A3(n4467), .A4(n4466), .ZN(n4474)
         );
  INV_X1 U5435 ( .A(REIP_REG_18__SCAN_IN), .ZN(n6958) );
  AOI22_X1 U5436 ( .A1(n6442), .A2(keyinput74), .B1(n6958), .B2(keyinput118), 
        .ZN(n4470) );
  OAI221_X1 U5437 ( .B1(n6442), .B2(keyinput74), .C1(n6958), .C2(keyinput118), 
        .A(n4470), .ZN(n4473) );
  INV_X1 U5438 ( .A(LWORD_REG_1__SCAN_IN), .ZN(n6430) );
  INV_X1 U5439 ( .A(EBX_REG_17__SCAN_IN), .ZN(n6281) );
  AOI22_X1 U5440 ( .A1(n6430), .A2(keyinput73), .B1(n6281), .B2(keyinput104), 
        .ZN(n4471) );
  OAI221_X1 U5441 ( .B1(n6430), .B2(keyinput73), .C1(n6281), .C2(keyinput104), 
        .A(n4471), .ZN(n4472) );
  NOR3_X1 U5442 ( .A1(n4474), .A2(n4473), .A3(n4472), .ZN(n4494) );
  OAI22_X1 U5443 ( .A1(BYTEENABLE_REG_0__SCAN_IN), .A2(keyinput105), .B1(
        keyinput78), .B2(DATAI_26_), .ZN(n4475) );
  AOI221_X1 U5444 ( .B1(BYTEENABLE_REG_0__SCAN_IN), .B2(keyinput105), .C1(
        DATAI_26_), .C2(keyinput78), .A(n4475), .ZN(n4482) );
  OAI22_X1 U5445 ( .A1(INSTQUEUE_REG_10__5__SCAN_IN), .A2(keyinput25), .B1(
        keyinput90), .B2(DATAO_REG_15__SCAN_IN), .ZN(n4476) );
  AOI221_X1 U5446 ( .B1(INSTQUEUE_REG_10__5__SCAN_IN), .B2(keyinput25), .C1(
        DATAO_REG_15__SCAN_IN), .C2(keyinput90), .A(n4476), .ZN(n4481) );
  OAI22_X1 U5447 ( .A1(INSTQUEUE_REG_8__4__SCAN_IN), .A2(keyinput29), .B1(
        keyinput44), .B2(ADDRESS_REG_5__SCAN_IN), .ZN(n4477) );
  AOI221_X1 U5448 ( .B1(INSTQUEUE_REG_8__4__SCAN_IN), .B2(keyinput29), .C1(
        ADDRESS_REG_5__SCAN_IN), .C2(keyinput44), .A(n4477), .ZN(n4480) );
  OAI22_X1 U5449 ( .A1(PHYADDRPOINTER_REG_14__SCAN_IN), .A2(keyinput9), .B1(
        DATAO_REG_28__SCAN_IN), .B2(keyinput92), .ZN(n4478) );
  AOI221_X1 U5450 ( .B1(PHYADDRPOINTER_REG_14__SCAN_IN), .B2(keyinput9), .C1(
        keyinput92), .C2(DATAO_REG_28__SCAN_IN), .A(n4478), .ZN(n4479) );
  NAND4_X1 U5451 ( .A1(n4482), .A2(n4481), .A3(n4480), .A4(n4479), .ZN(n4492)
         );
  OAI22_X1 U5452 ( .A1(INSTQUEUE_REG_1__6__SCAN_IN), .A2(keyinput72), .B1(
        INSTQUEUE_REG_1__2__SCAN_IN), .B2(keyinput97), .ZN(n4483) );
  AOI221_X1 U5453 ( .B1(INSTQUEUE_REG_1__6__SCAN_IN), .B2(keyinput72), .C1(
        keyinput97), .C2(INSTQUEUE_REG_1__2__SCAN_IN), .A(n4483), .ZN(n4490)
         );
  OAI22_X1 U5454 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(keyinput120), .B1(
        keyinput100), .B2(LWORD_REG_15__SCAN_IN), .ZN(n4484) );
  AOI221_X1 U5455 ( .B1(INSTQUEUE_REG_11__0__SCAN_IN), .B2(keyinput120), .C1(
        LWORD_REG_15__SCAN_IN), .C2(keyinput100), .A(n4484), .ZN(n4489) );
  OAI22_X1 U5456 ( .A1(INSTQUEUE_REG_0__2__SCAN_IN), .A2(keyinput126), .B1(
        INSTQUEUE_REG_2__2__SCAN_IN), .B2(keyinput32), .ZN(n4485) );
  AOI221_X1 U5457 ( .B1(INSTQUEUE_REG_0__2__SCAN_IN), .B2(keyinput126), .C1(
        keyinput32), .C2(INSTQUEUE_REG_2__2__SCAN_IN), .A(n4485), .ZN(n4488)
         );
  OAI22_X1 U5458 ( .A1(INSTQUEUE_REG_3__0__SCAN_IN), .A2(keyinput14), .B1(
        INSTADDRPOINTER_REG_5__SCAN_IN), .B2(keyinput11), .ZN(n4486) );
  AOI221_X1 U5459 ( .B1(INSTQUEUE_REG_3__0__SCAN_IN), .B2(keyinput14), .C1(
        keyinput11), .C2(INSTADDRPOINTER_REG_5__SCAN_IN), .A(n4486), .ZN(n4487) );
  NAND4_X1 U5460 ( .A1(n4490), .A2(n4489), .A3(n4488), .A4(n4487), .ZN(n4491)
         );
  NOR2_X1 U5461 ( .A1(n4492), .A2(n4491), .ZN(n4493) );
  NAND4_X1 U5462 ( .A1(n4496), .A2(n4495), .A3(n4494), .A4(n4493), .ZN(n4540)
         );
  AOI22_X1 U5463 ( .A1(ADDRESS_REG_15__SCAN_IN), .A2(keyinput40), .B1(
        INSTQUEUE_REG_3__2__SCAN_IN), .B2(keyinput111), .ZN(n4497) );
  OAI221_X1 U5464 ( .B1(ADDRESS_REG_15__SCAN_IN), .B2(keyinput40), .C1(
        INSTQUEUE_REG_3__2__SCAN_IN), .C2(keyinput111), .A(n4497), .ZN(n4505)
         );
  INV_X1 U5465 ( .A(REIP_REG_12__SCAN_IN), .ZN(n6948) );
  AOI22_X1 U5466 ( .A1(INSTADDRPOINTER_REG_29__SCAN_IN), .A2(keyinput79), .B1(
        n6948), .B2(keyinput7), .ZN(n4498) );
  OAI221_X1 U5467 ( .B1(INSTADDRPOINTER_REG_29__SCAN_IN), .B2(keyinput79), 
        .C1(n6948), .C2(keyinput7), .A(n4498), .ZN(n4504) );
  INV_X1 U5468 ( .A(DATAO_REG_2__SCAN_IN), .ZN(n6429) );
  AOI22_X1 U5469 ( .A1(n6339), .A2(keyinput22), .B1(n6429), .B2(keyinput108), 
        .ZN(n4499) );
  OAI221_X1 U5470 ( .B1(n6339), .B2(keyinput22), .C1(n6429), .C2(keyinput108), 
        .A(n4499), .ZN(n4503) );
  INV_X1 U5471 ( .A(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n4501) );
  AOI22_X1 U5472 ( .A1(n5250), .A2(keyinput103), .B1(n4501), .B2(keyinput36), 
        .ZN(n4500) );
  OAI221_X1 U5473 ( .B1(n5250), .B2(keyinput103), .C1(n4501), .C2(keyinput36), 
        .A(n4500), .ZN(n4502) );
  NOR4_X1 U5474 ( .A1(n4505), .A2(n4504), .A3(n4503), .A4(n4502), .ZN(n4538)
         );
  INV_X1 U5475 ( .A(EBX_REG_8__SCAN_IN), .ZN(n6304) );
  INV_X1 U5476 ( .A(REIP_REG_9__SCAN_IN), .ZN(n4789) );
  AOI22_X1 U5477 ( .A1(n6304), .A2(keyinput37), .B1(n4789), .B2(keyinput23), 
        .ZN(n4506) );
  OAI221_X1 U5478 ( .B1(n6304), .B2(keyinput37), .C1(n4789), .C2(keyinput23), 
        .A(n4506), .ZN(n4513) );
  AOI22_X1 U5479 ( .A1(n6070), .A2(keyinput26), .B1(keyinput43), .B2(n5236), 
        .ZN(n4507) );
  OAI221_X1 U5480 ( .B1(n6070), .B2(keyinput26), .C1(n5236), .C2(keyinput43), 
        .A(n4507), .ZN(n4512) );
  AOI22_X1 U5481 ( .A1(n6073), .A2(keyinput121), .B1(keyinput30), .B2(n6402), 
        .ZN(n4508) );
  OAI221_X1 U5482 ( .B1(n6073), .B2(keyinput121), .C1(n6402), .C2(keyinput30), 
        .A(n4508), .ZN(n4511) );
  INV_X1 U5483 ( .A(EBX_REG_14__SCAN_IN), .ZN(n6290) );
  AOI22_X1 U5484 ( .A1(n6290), .A2(keyinput123), .B1(n6423), .B2(keyinput45), 
        .ZN(n4509) );
  OAI221_X1 U5485 ( .B1(n6290), .B2(keyinput123), .C1(n6423), .C2(keyinput45), 
        .A(n4509), .ZN(n4510) );
  NOR4_X1 U5486 ( .A1(n4513), .A2(n4512), .A3(n4511), .A4(n4510), .ZN(n4537)
         );
  AOI22_X1 U5487 ( .A1(n6968), .A2(keyinput18), .B1(keyinput110), .B2(n6983), 
        .ZN(n4514) );
  OAI221_X1 U5488 ( .B1(n6968), .B2(keyinput18), .C1(n6983), .C2(keyinput110), 
        .A(n4514), .ZN(n4523) );
  AOI22_X1 U5489 ( .A1(n6909), .A2(keyinput66), .B1(keyinput41), .B2(n5276), 
        .ZN(n4515) );
  OAI221_X1 U5490 ( .B1(n6909), .B2(keyinput66), .C1(n5276), .C2(keyinput41), 
        .A(n4515), .ZN(n4522) );
  AOI22_X1 U5491 ( .A1(n4517), .A2(keyinput75), .B1(n6755), .B2(keyinput119), 
        .ZN(n4516) );
  OAI221_X1 U5492 ( .B1(n4517), .B2(keyinput75), .C1(n6755), .C2(keyinput119), 
        .A(n4516), .ZN(n4521) );
  INV_X1 U5493 ( .A(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n4519) );
  AOI22_X1 U5494 ( .A1(n4519), .A2(keyinput49), .B1(keyinput42), .B2(n6405), 
        .ZN(n4518) );
  OAI221_X1 U5495 ( .B1(n4519), .B2(keyinput49), .C1(n6405), .C2(keyinput42), 
        .A(n4518), .ZN(n4520) );
  NOR4_X1 U5496 ( .A1(n4523), .A2(n4522), .A3(n4521), .A4(n4520), .ZN(n4536)
         );
  INV_X1 U5497 ( .A(REIP_REG_28__SCAN_IN), .ZN(n6978) );
  INV_X1 U5498 ( .A(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n4525) );
  AOI22_X1 U5499 ( .A1(n6978), .A2(keyinput8), .B1(n4525), .B2(keyinput17), 
        .ZN(n4524) );
  OAI221_X1 U5500 ( .B1(n6978), .B2(keyinput8), .C1(n4525), .C2(keyinput17), 
        .A(n4524), .ZN(n4534) );
  INV_X1 U5501 ( .A(DATAI_25_), .ZN(n4527) );
  AOI22_X1 U5502 ( .A1(n4528), .A2(keyinput93), .B1(keyinput87), .B2(n4527), 
        .ZN(n4526) );
  OAI221_X1 U5503 ( .B1(n4528), .B2(keyinput93), .C1(n4527), .C2(keyinput87), 
        .A(n4526), .ZN(n4533) );
  AOI22_X1 U5504 ( .A1(n6952), .A2(keyinput115), .B1(n6440), .B2(keyinput15), 
        .ZN(n4529) );
  OAI221_X1 U5505 ( .B1(n6952), .B2(keyinput115), .C1(n6440), .C2(keyinput15), 
        .A(n4529), .ZN(n4532) );
  INV_X1 U5506 ( .A(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n6842) );
  AOI22_X1 U5507 ( .A1(n6842), .A2(keyinput6), .B1(keyinput46), .B2(n6931), 
        .ZN(n4530) );
  OAI221_X1 U5508 ( .B1(n6842), .B2(keyinput6), .C1(n6931), .C2(keyinput46), 
        .A(n4530), .ZN(n4531) );
  NOR4_X1 U5509 ( .A1(n4534), .A2(n4533), .A3(n4532), .A4(n4531), .ZN(n4535)
         );
  NAND4_X1 U5510 ( .A1(n4538), .A2(n4537), .A3(n4536), .A4(n4535), .ZN(n4539)
         );
  NOR2_X1 U5511 ( .A1(n4540), .A2(n4539), .ZN(n4577) );
  INV_X1 U5512 ( .A(BE_N_REG_1__SCAN_IN), .ZN(n6989) );
  AOI22_X1 U5513 ( .A1(n6989), .A2(keyinput112), .B1(keyinput101), .B2(n5922), 
        .ZN(n4541) );
  OAI221_X1 U5514 ( .B1(n6989), .B2(keyinput112), .C1(n5922), .C2(keyinput101), 
        .A(n4541), .ZN(n4549) );
  INV_X1 U5515 ( .A(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n4543) );
  INV_X1 U5516 ( .A(ADDRESS_REG_25__SCAN_IN), .ZN(n6973) );
  AOI22_X1 U5517 ( .A1(n4543), .A2(keyinput77), .B1(keyinput102), .B2(n6973), 
        .ZN(n4542) );
  OAI221_X1 U5518 ( .B1(n4543), .B2(keyinput77), .C1(n6973), .C2(keyinput102), 
        .A(n4542), .ZN(n4548) );
  INV_X1 U5519 ( .A(UWORD_REG_10__SCAN_IN), .ZN(n6449) );
  AOI22_X1 U5520 ( .A1(n6449), .A2(keyinput35), .B1(keyinput20), .B2(n6977), 
        .ZN(n4544) );
  OAI221_X1 U5521 ( .B1(n6449), .B2(keyinput35), .C1(n6977), .C2(keyinput20), 
        .A(n4544), .ZN(n4547) );
  INV_X1 U5522 ( .A(UWORD_REG_4__SCAN_IN), .ZN(n6445) );
  AOI22_X1 U5523 ( .A1(n6392), .A2(keyinput99), .B1(n6445), .B2(keyinput55), 
        .ZN(n4545) );
  OAI221_X1 U5524 ( .B1(n6392), .B2(keyinput99), .C1(n6445), .C2(keyinput55), 
        .A(n4545), .ZN(n4546) );
  NOR4_X1 U5525 ( .A1(n4549), .A2(n4548), .A3(n4547), .A4(n4546), .ZN(n4576)
         );
  INV_X1 U5526 ( .A(DATAWIDTH_REG_3__SCAN_IN), .ZN(n6911) );
  AOI22_X1 U5527 ( .A1(n6911), .A2(keyinput96), .B1(n4551), .B2(keyinput54), 
        .ZN(n4550) );
  OAI221_X1 U5528 ( .B1(n6911), .B2(keyinput96), .C1(n4551), .C2(keyinput54), 
        .A(n4550), .ZN(n4559) );
  INV_X1 U5529 ( .A(EAX_REG_2__SCAN_IN), .ZN(n6428) );
  AOI22_X1 U5530 ( .A1(n6428), .A2(keyinput51), .B1(keyinput3), .B2(n6969), 
        .ZN(n4552) );
  OAI221_X1 U5531 ( .B1(n6428), .B2(keyinput51), .C1(n6969), .C2(keyinput3), 
        .A(n4552), .ZN(n4558) );
  INV_X1 U5532 ( .A(EAX_REG_13__SCAN_IN), .ZN(n6404) );
  AOI22_X1 U5533 ( .A1(n6404), .A2(keyinput69), .B1(keyinput85), .B2(n5665), 
        .ZN(n4553) );
  OAI221_X1 U5534 ( .B1(n6404), .B2(keyinput69), .C1(n5665), .C2(keyinput85), 
        .A(n4553), .ZN(n4557) );
  AOI22_X1 U5535 ( .A1(n4555), .A2(keyinput70), .B1(keyinput13), .B2(n6941), 
        .ZN(n4554) );
  OAI221_X1 U5536 ( .B1(n4555), .B2(keyinput70), .C1(n6941), .C2(keyinput13), 
        .A(n4554), .ZN(n4556) );
  NOR4_X1 U5537 ( .A1(n4559), .A2(n4558), .A3(n4557), .A4(n4556), .ZN(n4575)
         );
  INV_X1 U5538 ( .A(ADDRESS_REG_18__SCAN_IN), .ZN(n6961) );
  INV_X1 U5539 ( .A(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n4561) );
  AOI22_X1 U5540 ( .A1(n6961), .A2(keyinput60), .B1(n4561), .B2(keyinput12), 
        .ZN(n4560) );
  OAI221_X1 U5541 ( .B1(n6961), .B2(keyinput60), .C1(n4561), .C2(keyinput12), 
        .A(n4560), .ZN(n4573) );
  AOI22_X1 U5542 ( .A1(n4563), .A2(keyinput68), .B1(keyinput47), .B2(n6144), 
        .ZN(n4562) );
  OAI221_X1 U5543 ( .B1(n4563), .B2(keyinput68), .C1(n6144), .C2(keyinput47), 
        .A(n4562), .ZN(n4572) );
  INV_X1 U5544 ( .A(DATAI_30_), .ZN(n4566) );
  AOI22_X1 U5545 ( .A1(n4566), .A2(keyinput39), .B1(n4565), .B2(keyinput125), 
        .ZN(n4564) );
  OAI221_X1 U5546 ( .B1(n4566), .B2(keyinput39), .C1(n4565), .C2(keyinput125), 
        .A(n4564), .ZN(n4571) );
  AOI22_X1 U5547 ( .A1(n4569), .A2(keyinput52), .B1(keyinput91), .B2(n4568), 
        .ZN(n4567) );
  OAI221_X1 U5548 ( .B1(n4569), .B2(keyinput52), .C1(n4568), .C2(keyinput91), 
        .A(n4567), .ZN(n4570) );
  NOR4_X1 U5549 ( .A1(n4573), .A2(n4572), .A3(n4571), .A4(n4570), .ZN(n4574)
         );
  NAND4_X1 U5550 ( .A1(n4577), .A2(n4576), .A3(n4575), .A4(n4574), .ZN(n4578)
         );
  XNOR2_X1 U5551 ( .A(n4580), .B(n3287), .ZN(U2957) );
  INV_X1 U5552 ( .A(n5681), .ZN(n4583) );
  OAI21_X1 U5553 ( .B1(n4583), .B2(INSTADDRPOINTER_REG_27__SCAN_IN), .A(n4582), 
        .ZN(n4584) );
  INV_X1 U5554 ( .A(n4585), .ZN(n6848) );
  NAND2_X1 U5555 ( .A1(n6848), .A2(n4812), .ZN(n4743) );
  NAND2_X1 U5556 ( .A1(n4586), .A2(n5234), .ZN(n6876) );
  NAND2_X1 U5557 ( .A1(n4999), .A2(n3446), .ZN(n5268) );
  AND2_X1 U5558 ( .A1(n5267), .A2(n5268), .ZN(n5266) );
  OR2_X1 U5559 ( .A1(n4587), .A2(n5266), .ZN(n4590) );
  AOI21_X1 U5560 ( .B1(n4588), .B2(n4812), .A(n5234), .ZN(n4589) );
  NAND2_X1 U5561 ( .A1(n4590), .A2(n4589), .ZN(n4738) );
  NAND2_X1 U5562 ( .A1(n4609), .A2(n4738), .ZN(n4591) );
  NAND2_X1 U5563 ( .A1(n6876), .A2(n4591), .ZN(n4873) );
  OR2_X1 U5564 ( .A1(n4592), .A2(STATE_REG_0__SCAN_IN), .ZN(n6917) );
  INV_X1 U5565 ( .A(n6917), .ZN(n4869) );
  AND3_X1 U5566 ( .A1(n4596), .A2(n4595), .A3(n4594), .ZN(n4598) );
  OAI21_X1 U5567 ( .B1(n4599), .B2(n4598), .A(n4597), .ZN(n6877) );
  INV_X1 U5568 ( .A(READY_N), .ZN(n7024) );
  NAND2_X1 U5569 ( .A1(n6877), .A2(n7024), .ZN(n4875) );
  INV_X1 U5570 ( .A(n4875), .ZN(n4600) );
  OAI211_X1 U5571 ( .C1(n3714), .C2(n4869), .A(n4593), .B(n4600), .ZN(n4601)
         );
  OAI211_X1 U5572 ( .C1(n6891), .C2(n4743), .A(n4873), .B(n4601), .ZN(n4602)
         );
  NAND2_X1 U5573 ( .A1(n4602), .A2(n5889), .ZN(n4608) );
  NAND2_X1 U5574 ( .A1(n3714), .A2(n6917), .ZN(n4788) );
  NAND3_X1 U5575 ( .A1(n4603), .A2(n4788), .A3(n7024), .ZN(n4604) );
  NAND3_X1 U5576 ( .A1(n4604), .A2(n3444), .A3(n5267), .ZN(n4605) );
  NAND2_X1 U5577 ( .A1(n4605), .A2(n3426), .ZN(n4606) );
  OR2_X1 U5578 ( .A1(n5762), .A2(n4606), .ZN(n4607) );
  AND2_X1 U5579 ( .A1(n4609), .A2(n6199), .ZN(n5010) );
  NOR2_X1 U5580 ( .A1(n5010), .A2(n4610), .ZN(n6870) );
  NAND2_X1 U5581 ( .A1(n3444), .A2(n4812), .ZN(n4635) );
  AOI22_X1 U5582 ( .A1(n4603), .A2(n6250), .B1(n4612), .B2(n4611), .ZN(n4614)
         );
  AND3_X1 U5583 ( .A1(n6870), .A2(n4614), .A3(n4613), .ZN(n4615) );
  NAND2_X1 U5584 ( .A1(n3177), .A2(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4618)
         );
  NOR2_X1 U5585 ( .A1(n4635), .A2(EBX_REG_1__SCAN_IN), .ZN(n4617) );
  MUX2_X1 U5586 ( .A(n4618), .B(n3177), .S(n4617), .Z(n4621) );
  NAND2_X1 U5587 ( .A1(n4708), .A2(EBX_REG_1__SCAN_IN), .ZN(n4619) );
  AND2_X1 U5588 ( .A1(n4710), .A2(n4619), .ZN(n4620) );
  INV_X1 U5589 ( .A(EBX_REG_0__SCAN_IN), .ZN(n4622) );
  OR2_X1 U5590 ( .A1(n4708), .A2(n4622), .ZN(n4624) );
  NAND2_X1 U5591 ( .A1(n3206), .A2(n4622), .ZN(n4623) );
  NAND2_X1 U5592 ( .A1(n4624), .A2(n4623), .ZN(n4860) );
  XNOR2_X1 U5593 ( .A(n4625), .B(n4860), .ZN(n6251) );
  NAND2_X1 U5594 ( .A1(n6251), .A2(n6250), .ZN(n6252) );
  NAND2_X1 U5595 ( .A1(n6252), .A2(n4625), .ZN(n4920) );
  INV_X1 U5596 ( .A(n4920), .ZN(n4632) );
  NAND2_X1 U5597 ( .A1(n3206), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n4627)
         );
  NOR2_X1 U5598 ( .A1(n4635), .A2(EBX_REG_2__SCAN_IN), .ZN(n4626) );
  MUX2_X1 U5599 ( .A(n4627), .B(n3206), .S(n4626), .Z(n4630) );
  NAND2_X1 U5600 ( .A1(n4708), .A2(EBX_REG_2__SCAN_IN), .ZN(n4628) );
  AND2_X1 U5601 ( .A1(n4710), .A2(n4628), .ZN(n4629) );
  AND2_X1 U5602 ( .A1(n4630), .A2(n4629), .ZN(n4919) );
  NAND2_X1 U5603 ( .A1(n3177), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4633)
         );
  OAI211_X1 U5604 ( .C1(n3205), .C2(EBX_REG_3__SCAN_IN), .A(n4723), .B(n4633), 
        .ZN(n4634) );
  OAI21_X1 U5605 ( .B1(n4713), .B2(EBX_REG_3__SCAN_IN), .A(n4634), .ZN(n4956)
         );
  NAND2_X1 U5606 ( .A1(n3206), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4637)
         );
  NOR2_X1 U5607 ( .A1(n3205), .A2(EBX_REG_4__SCAN_IN), .ZN(n4636) );
  MUX2_X1 U5608 ( .A(n4637), .B(n3206), .S(n4636), .Z(n4640) );
  NAND2_X1 U5609 ( .A1(n4708), .A2(EBX_REG_4__SCAN_IN), .ZN(n4638) );
  AND2_X1 U5610 ( .A1(n4710), .A2(n4638), .ZN(n4639) );
  NAND2_X1 U5611 ( .A1(n4640), .A2(n4639), .ZN(n4927) );
  NAND2_X1 U5612 ( .A1(n3206), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4641)
         );
  OAI211_X1 U5613 ( .C1(n3205), .C2(EBX_REG_5__SCAN_IN), .A(n4723), .B(n4641), 
        .ZN(n4642) );
  OAI21_X1 U5614 ( .B1(n4713), .B2(EBX_REG_5__SCAN_IN), .A(n4642), .ZN(n4940)
         );
  INV_X1 U5615 ( .A(EBX_REG_6__SCAN_IN), .ZN(n6308) );
  NAND2_X1 U5616 ( .A1(n3203), .A2(n6308), .ZN(n4648) );
  NAND2_X1 U5617 ( .A1(n4723), .A2(n4644), .ZN(n4646) );
  NAND2_X1 U5618 ( .A1(n6250), .A2(n6308), .ZN(n4645) );
  NAND3_X1 U5619 ( .A1(n4646), .A2(n3206), .A3(n4645), .ZN(n4647) );
  NAND2_X1 U5620 ( .A1(n3206), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n4649)
         );
  OAI211_X1 U5621 ( .C1(n3205), .C2(EBX_REG_7__SCAN_IN), .A(n4723), .B(n4649), 
        .ZN(n4650) );
  OAI21_X1 U5622 ( .B1(n4713), .B2(EBX_REG_7__SCAN_IN), .A(n4650), .ZN(n6178)
         );
  NOR2_X2 U5623 ( .A1(n6179), .A2(n6178), .ZN(n6180) );
  NAND2_X1 U5624 ( .A1(n4780), .A2(EBX_REG_8__SCAN_IN), .ZN(n4652) );
  NAND2_X1 U5625 ( .A1(n3205), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n4651)
         );
  NAND2_X1 U5626 ( .A1(n4652), .A2(n4651), .ZN(n4653) );
  XNOR2_X1 U5627 ( .A(n4653), .B(n3206), .ZN(n5245) );
  NAND2_X1 U5628 ( .A1(n6180), .A2(n5245), .ZN(n6161) );
  INV_X1 U5629 ( .A(n6161), .ZN(n4657) );
  NAND2_X1 U5630 ( .A1(n3206), .A2(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n4654)
         );
  OAI211_X1 U5631 ( .C1(n3205), .C2(EBX_REG_9__SCAN_IN), .A(n4723), .B(n4654), 
        .ZN(n4655) );
  OAI21_X1 U5632 ( .B1(n4713), .B2(EBX_REG_9__SCAN_IN), .A(n4655), .ZN(n6162)
         );
  INV_X1 U5633 ( .A(EBX_REG_10__SCAN_IN), .ZN(n6299) );
  NAND2_X1 U5634 ( .A1(n3203), .A2(n6299), .ZN(n4661) );
  NAND2_X1 U5635 ( .A1(n4723), .A2(n5464), .ZN(n4659) );
  NAND2_X1 U5636 ( .A1(n6250), .A2(n6299), .ZN(n4658) );
  NAND3_X1 U5637 ( .A1(n4659), .A2(n3206), .A3(n4658), .ZN(n4660) );
  MUX2_X1 U5638 ( .A(n4713), .B(n3177), .S(EBX_REG_11__SCAN_IN), .Z(n4662) );
  INV_X1 U5639 ( .A(n4662), .ZN(n4664) );
  NOR2_X1 U5640 ( .A1(n4780), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n4663)
         );
  NOR2_X1 U5641 ( .A1(n4664), .A2(n4663), .ZN(n5485) );
  NAND2_X1 U5642 ( .A1(n4780), .A2(EBX_REG_12__SCAN_IN), .ZN(n4666) );
  NAND2_X1 U5643 ( .A1(n3205), .A2(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n4665) );
  NAND2_X1 U5644 ( .A1(n4666), .A2(n4665), .ZN(n4667) );
  XNOR2_X1 U5645 ( .A(n4667), .B(n3203), .ZN(n5524) );
  NAND2_X1 U5646 ( .A1(n3206), .A2(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n4668) );
  OAI211_X1 U5647 ( .C1(n3205), .C2(EBX_REG_13__SCAN_IN), .A(n4723), .B(n4668), 
        .ZN(n4669) );
  OAI21_X1 U5648 ( .B1(n4713), .B2(EBX_REG_13__SCAN_IN), .A(n4669), .ZN(n5529)
         );
  NOR2_X1 U5649 ( .A1(n5524), .A2(n5529), .ZN(n4670) );
  NAND2_X1 U5650 ( .A1(n4780), .A2(EBX_REG_14__SCAN_IN), .ZN(n4672) );
  NAND2_X1 U5651 ( .A1(n3205), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n4671) );
  NAND2_X1 U5652 ( .A1(n4672), .A2(n4671), .ZN(n4673) );
  XNOR2_X1 U5653 ( .A(n4673), .B(n3203), .ZN(n5549) );
  NAND2_X1 U5654 ( .A1(n3206), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n4674) );
  OAI211_X1 U5655 ( .C1(n3205), .C2(EBX_REG_15__SCAN_IN), .A(n4723), .B(n4674), 
        .ZN(n4675) );
  OAI21_X1 U5656 ( .B1(n4713), .B2(EBX_REG_15__SCAN_IN), .A(n4675), .ZN(n6059)
         );
  NAND2_X1 U5657 ( .A1(n4780), .A2(EBX_REG_16__SCAN_IN), .ZN(n4677) );
  NAND2_X1 U5658 ( .A1(n3205), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n4676) );
  NAND2_X1 U5659 ( .A1(n4677), .A2(n4676), .ZN(n4678) );
  XNOR2_X1 U5660 ( .A(n4678), .B(n3206), .ZN(n6048) );
  NAND2_X1 U5661 ( .A1(n4780), .A2(EBX_REG_17__SCAN_IN), .ZN(n4680) );
  NAND2_X1 U5662 ( .A1(n3205), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n4679) );
  NAND2_X1 U5663 ( .A1(n4680), .A2(n4679), .ZN(n4681) );
  XNOR2_X1 U5664 ( .A(n4681), .B(n3203), .ZN(n5565) );
  NAND2_X1 U5665 ( .A1(n3206), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n4683) );
  NOR2_X1 U5666 ( .A1(n3205), .A2(EBX_REG_19__SCAN_IN), .ZN(n4682) );
  MUX2_X1 U5667 ( .A(n4683), .B(n3177), .S(n4682), .Z(n4686) );
  NAND2_X1 U5668 ( .A1(n4708), .A2(EBX_REG_19__SCAN_IN), .ZN(n4684) );
  AND2_X1 U5669 ( .A1(n4710), .A2(n4684), .ZN(n4685) );
  NAND2_X1 U5670 ( .A1(n4780), .A2(EBX_REG_18__SCAN_IN), .ZN(n4689) );
  NAND2_X1 U5671 ( .A1(n3205), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n4688) );
  NAND2_X1 U5672 ( .A1(n4689), .A2(n4688), .ZN(n5866) );
  OR2_X1 U5673 ( .A1(n5866), .A2(n3206), .ZN(n5878) );
  NAND2_X1 U5674 ( .A1(n5866), .A2(n3177), .ZN(n5877) );
  OR2_X1 U5675 ( .A1(n4780), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n4691)
         );
  NAND2_X1 U5676 ( .A1(n6250), .A2(n5922), .ZN(n4690) );
  NAND2_X1 U5677 ( .A1(n4691), .A2(n4690), .ZN(n5868) );
  OAI22_X1 U5678 ( .A1(EBX_REG_20__SCAN_IN), .A2(n5878), .B1(n5877), .B2(n5868), .ZN(n4692) );
  INV_X1 U5679 ( .A(n4692), .ZN(n4693) );
  NAND2_X1 U5680 ( .A1(n3177), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n4695) );
  NOR2_X1 U5681 ( .A1(n3205), .A2(EBX_REG_21__SCAN_IN), .ZN(n4694) );
  MUX2_X1 U5682 ( .A(n4695), .B(n3206), .S(n4694), .Z(n4698) );
  NAND2_X1 U5683 ( .A1(n4708), .A2(EBX_REG_21__SCAN_IN), .ZN(n4696) );
  AND2_X1 U5684 ( .A1(n4710), .A2(n4696), .ZN(n4697) );
  NAND2_X1 U5685 ( .A1(n4698), .A2(n4697), .ZN(n5726) );
  MUX2_X1 U5686 ( .A(n4713), .B(n3206), .S(EBX_REG_22__SCAN_IN), .Z(n4699) );
  INV_X1 U5687 ( .A(n4699), .ZN(n4701) );
  NOR2_X1 U5688 ( .A1(n4780), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n4700)
         );
  NOR2_X1 U5689 ( .A1(n4701), .A2(n4700), .ZN(n5842) );
  NAND2_X1 U5690 ( .A1(n4723), .A2(n5716), .ZN(n4703) );
  INV_X1 U5691 ( .A(EBX_REG_23__SCAN_IN), .ZN(n5915) );
  NAND2_X1 U5692 ( .A1(n6250), .A2(n5915), .ZN(n4702) );
  NAND3_X1 U5693 ( .A1(n4703), .A2(n3206), .A3(n4702), .ZN(n4704) );
  OAI21_X1 U5694 ( .B1(n3206), .B2(EBX_REG_23__SCAN_IN), .A(n4704), .ZN(n5711)
         );
  MUX2_X1 U5695 ( .A(n4713), .B(n3206), .S(EBX_REG_24__SCAN_IN), .Z(n4705) );
  NAND2_X1 U5696 ( .A1(n3285), .A2(n4705), .ZN(n5701) );
  NAND2_X1 U5697 ( .A1(n3206), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n4707) );
  NOR2_X1 U5698 ( .A1(n3205), .A2(EBX_REG_25__SCAN_IN), .ZN(n4706) );
  MUX2_X1 U5699 ( .A(n4707), .B(n3206), .S(n4706), .Z(n4712) );
  NAND2_X1 U5700 ( .A1(n4708), .A2(EBX_REG_25__SCAN_IN), .ZN(n4709) );
  AND2_X1 U5701 ( .A1(n4710), .A2(n4709), .ZN(n4711) );
  NAND2_X1 U5702 ( .A1(n4712), .A2(n4711), .ZN(n5811) );
  INV_X1 U5703 ( .A(n4713), .ZN(n4721) );
  INV_X1 U5704 ( .A(EBX_REG_26__SCAN_IN), .ZN(n5908) );
  NAND2_X1 U5705 ( .A1(n4721), .A2(n5908), .ZN(n4716) );
  NAND2_X1 U5706 ( .A1(n3206), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n4714) );
  OAI211_X1 U5707 ( .C1(n3205), .C2(EBX_REG_26__SCAN_IN), .A(n4723), .B(n4714), 
        .ZN(n4715) );
  AND2_X1 U5708 ( .A1(n4716), .A2(n4715), .ZN(n5810) );
  NAND2_X1 U5709 ( .A1(n5811), .A2(n5810), .ZN(n4717) );
  NAND2_X1 U5710 ( .A1(n4723), .A2(n5688), .ZN(n4719) );
  INV_X1 U5711 ( .A(EBX_REG_27__SCAN_IN), .ZN(n5905) );
  NAND2_X1 U5712 ( .A1(n6250), .A2(n5905), .ZN(n4718) );
  NAND3_X1 U5713 ( .A1(n4719), .A2(n3206), .A3(n4718), .ZN(n4720) );
  OAI21_X1 U5714 ( .B1(n3206), .B2(EBX_REG_27__SCAN_IN), .A(n4720), .ZN(n5683)
         );
  AND2_X2 U5715 ( .A1(n5813), .A2(n5683), .ZN(n5685) );
  INV_X1 U5716 ( .A(EBX_REG_28__SCAN_IN), .ZN(n5904) );
  NAND2_X1 U5717 ( .A1(n4721), .A2(n5904), .ZN(n4725) );
  NAND2_X1 U5718 ( .A1(n3206), .A2(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n4722) );
  OAI211_X1 U5719 ( .C1(n3205), .C2(EBX_REG_28__SCAN_IN), .A(n4723), .B(n4722), 
        .ZN(n4724) );
  AND2_X1 U5720 ( .A1(n4725), .A2(n4724), .ZN(n4726) );
  OR2_X1 U5721 ( .A1(n5685), .A2(n4726), .ZN(n4727) );
  NAND2_X1 U5722 ( .A1(n4603), .A2(n3567), .ZN(n6884) );
  INV_X1 U5723 ( .A(n4728), .ZN(n4730) );
  INV_X1 U5724 ( .A(n5267), .ZN(n4729) );
  NAND3_X1 U5725 ( .A1(n4730), .A2(n3456), .A3(n4729), .ZN(n4731) );
  AND2_X1 U5726 ( .A1(n6884), .A2(n4731), .ZN(n4732) );
  NAND2_X1 U5727 ( .A1(INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5999) );
  AOI22_X1 U5728 ( .A1(n4733), .A2(n3203), .B1(n4593), .B2(n5267), .ZN(n4737)
         );
  INV_X1 U5729 ( .A(n4780), .ZN(n4862) );
  OR2_X1 U5730 ( .A1(n3422), .A2(n4593), .ZN(n4872) );
  NAND2_X1 U5731 ( .A1(n4862), .A2(n4872), .ZN(n4735) );
  NAND2_X1 U5732 ( .A1(n4735), .A2(n4734), .ZN(n4736) );
  NAND3_X1 U5733 ( .A1(n4738), .A2(n4737), .A3(n4736), .ZN(n4739) );
  NOR2_X1 U5734 ( .A1(n4740), .A2(n4739), .ZN(n4886) );
  OAI21_X1 U5735 ( .B1(n4883), .B2(n3444), .A(n5021), .ZN(n4741) );
  INV_X1 U5736 ( .A(n4741), .ZN(n4742) );
  INV_X1 U5737 ( .A(n5484), .ZN(n4746) );
  INV_X1 U5738 ( .A(n4743), .ZN(n4744) );
  NAND2_X1 U5739 ( .A1(n4746), .A2(n4929), .ZN(n6530) );
  INV_X1 U5740 ( .A(n4929), .ZN(n5497) );
  NAND2_X1 U5741 ( .A1(n4747), .A2(n3179), .ZN(n4859) );
  INV_X1 U5742 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n5596) );
  NAND2_X1 U5743 ( .A1(n4929), .A2(n5557), .ZN(n5517) );
  NAND2_X1 U5744 ( .A1(n5596), .A2(n5517), .ZN(n4866) );
  NAND2_X1 U5745 ( .A1(n4859), .A2(n4866), .ZN(n6526) );
  NOR2_X1 U5746 ( .A1(n5497), .A2(n6526), .ZN(n5736) );
  NAND2_X1 U5747 ( .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n5522) );
  NOR2_X1 U5748 ( .A1(n4748), .A2(n5522), .ZN(n6046) );
  NAND3_X1 U5749 ( .A1(n6056), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .A3(n6046), .ZN(n5734) );
  NOR3_X1 U5750 ( .A1(n6023), .A2(n6021), .A3(n5734), .ZN(n4756) );
  NOR2_X1 U5751 ( .A1(n5250), .A2(n6521), .ZN(n5462) );
  NAND3_X1 U5752 ( .A1(INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_9__SCAN_IN), .A3(n5462), .ZN(n4749) );
  NAND2_X1 U5753 ( .A1(INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4932) );
  NAND2_X1 U5754 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4930) );
  NOR2_X1 U5755 ( .A1(n4932), .A2(n4930), .ZN(n4943) );
  NAND3_X1 U5756 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_5__SCAN_IN), .A3(n4943), .ZN(n5247) );
  NOR2_X1 U5757 ( .A1(n4749), .A2(n5247), .ZN(n4755) );
  NAND2_X1 U5758 ( .A1(n4755), .A2(n6046), .ZN(n5518) );
  NAND2_X1 U5759 ( .A1(n6056), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n6020) );
  OAI21_X1 U5760 ( .B1(n5596), .B2(n6531), .A(n3606), .ZN(n4931) );
  NAND3_X1 U5761 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .A3(n4931), .ZN(n4947) );
  NOR2_X1 U5762 ( .A1(n4929), .A2(n4947), .ZN(n4950) );
  NAND3_X1 U5763 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_5__SCAN_IN), .A3(n4950), .ZN(n5248) );
  NOR2_X1 U5764 ( .A1(n5736), .A2(n5556), .ZN(n5482) );
  AOI221_X1 U5765 ( .B1(n5518), .B2(n5484), .C1(n6020), .C2(n5484), .A(n5482), 
        .ZN(n5735) );
  OAI21_X1 U5766 ( .B1(n6021), .B2(n6023), .A(n5484), .ZN(n4750) );
  OAI211_X1 U5767 ( .C1(n5736), .C2(n4756), .A(n5735), .B(n4750), .ZN(n6006)
         );
  AND2_X1 U5768 ( .A1(n6530), .A2(n6010), .ZN(n4751) );
  NOR2_X1 U5769 ( .A1(n6006), .A2(n4751), .ZN(n5713) );
  NAND2_X1 U5770 ( .A1(n5596), .A2(n5516), .ZN(n6529) );
  NAND2_X1 U5771 ( .A1(n4944), .A2(n4929), .ZN(n4752) );
  NAND2_X1 U5772 ( .A1(n4752), .A2(n4757), .ZN(n4753) );
  NAND2_X1 U5773 ( .A1(n5713), .A2(n4753), .ZN(n5996) );
  AOI21_X1 U5774 ( .B1(n5999), .B2(n6530), .A(n5996), .ZN(n5687) );
  INV_X1 U5775 ( .A(n4755), .ZN(n5483) );
  INV_X1 U5776 ( .A(n6010), .ZN(n5634) );
  NAND2_X1 U5777 ( .A1(n6011), .A2(n5634), .ZN(n5709) );
  NOR2_X1 U5778 ( .A1(n4757), .A2(n5709), .ZN(n6000) );
  NAND3_X1 U5779 ( .A1(INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_25__SCAN_IN), .A3(n6000), .ZN(n5689) );
  NOR2_X1 U5780 ( .A1(n5674), .A2(n5689), .ZN(n4759) );
  AOI22_X1 U5781 ( .A1(REIP_REG_28__SCAN_IN), .A2(n6523), .B1(n4759), .B2(
        n4758), .ZN(n4760) );
  AND2_X1 U5782 ( .A1(n3195), .A2(n4766), .ZN(n4768) );
  OR2_X1 U5783 ( .A1(n4768), .A2(n4767), .ZN(n5790) );
  AOI22_X1 U5784 ( .A1(PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n6491), .B1(n6523), 
        .B2(REIP_REG_28__SCAN_IN), .ZN(n4769) );
  INV_X1 U5785 ( .A(n5768), .ZN(n4774) );
  NOR3_X1 U5786 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n7002), .A3(n4773), .ZN(
        n6903) );
  NAND2_X1 U5787 ( .A1(n4774), .A2(n6201), .ZN(n4809) );
  OR2_X1 U5788 ( .A1(n4780), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4777)
         );
  INV_X1 U5789 ( .A(EBX_REG_29__SCAN_IN), .ZN(n4775) );
  NAND2_X1 U5790 ( .A1(n6250), .A2(n4775), .ZN(n4776) );
  NAND2_X1 U5791 ( .A1(n4777), .A2(n4776), .ZN(n5655) );
  NAND2_X1 U5792 ( .A1(n5655), .A2(n3177), .ZN(n4779) );
  NAND2_X1 U5793 ( .A1(n3203), .A2(EBX_REG_29__SCAN_IN), .ZN(n4778) );
  NAND2_X1 U5794 ( .A1(n4779), .A2(n4778), .ZN(n5668) );
  OAI22_X1 U5795 ( .A1(n4862), .A2(n5898), .B1(n6250), .B2(n5665), .ZN(n5658)
         );
  NAND2_X1 U5796 ( .A1(n5669), .A2(n3206), .ZN(n5656) );
  AOI22_X1 U5797 ( .A1(n4780), .A2(EBX_REG_31__SCAN_IN), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n3205), .ZN(n4781) );
  XNOR2_X1 U5798 ( .A(n4782), .B(n4781), .ZN(n6274) );
  INV_X1 U5799 ( .A(n6876), .ZN(n4784) );
  NAND2_X1 U5800 ( .A1(n4784), .A2(n6877), .ZN(n6075) );
  INV_X1 U5801 ( .A(n5889), .ZN(n6901) );
  NOR2_X1 U5802 ( .A1(STATEBS16_REG_SCAN_IN), .A2(READY_N), .ZN(n4786) );
  INV_X1 U5803 ( .A(n4786), .ZN(n4803) );
  AND2_X1 U5804 ( .A1(n4787), .A2(n4803), .ZN(n5571) );
  AND2_X1 U5805 ( .A1(n4812), .A2(EBX_REG_31__SCAN_IN), .ZN(n4785) );
  INV_X1 U5806 ( .A(REIP_REG_13__SCAN_IN), .ZN(n6950) );
  INV_X1 U5807 ( .A(REIP_REG_11__SCAN_IN), .ZN(n6945) );
  INV_X1 U5808 ( .A(REIP_REG_6__SCAN_IN), .ZN(n6938) );
  INV_X1 U5809 ( .A(REIP_REG_4__SCAN_IN), .ZN(n6933) );
  NAND3_X1 U5810 ( .A1(REIP_REG_3__SCAN_IN), .A2(REIP_REG_1__SCAN_IN), .A3(
        REIP_REG_2__SCAN_IN), .ZN(n6218) );
  NOR2_X1 U5811 ( .A1(n6933), .A2(n6218), .ZN(n6208) );
  NAND2_X1 U5812 ( .A1(REIP_REG_5__SCAN_IN), .A2(n6208), .ZN(n6184) );
  NOR2_X1 U5813 ( .A1(n6938), .A2(n6184), .ZN(n6187) );
  NAND2_X1 U5814 ( .A1(REIP_REG_7__SCAN_IN), .A2(n6187), .ZN(n4793) );
  NAND2_X1 U5815 ( .A1(REIP_REG_8__SCAN_IN), .A2(n6173), .ZN(n6154) );
  NAND2_X1 U5816 ( .A1(REIP_REG_10__SCAN_IN), .A2(n6150), .ZN(n6142) );
  NAND2_X1 U5817 ( .A1(REIP_REG_12__SCAN_IN), .A2(n6126), .ZN(n6129) );
  NAND3_X1 U5818 ( .A1(REIP_REG_17__SCAN_IN), .A2(REIP_REG_16__SCAN_IN), .A3(
        REIP_REG_15__SCAN_IN), .ZN(n5579) );
  INV_X1 U5819 ( .A(REIP_REG_19__SCAN_IN), .ZN(n6962) );
  NOR3_X1 U5820 ( .A1(n6958), .A2(n5579), .A3(n6962), .ZN(n5863) );
  NAND2_X1 U5821 ( .A1(REIP_REG_20__SCAN_IN), .A2(n5863), .ZN(n4797) );
  NAND4_X1 U5822 ( .A1(REIP_REG_23__SCAN_IN), .A2(REIP_REG_22__SCAN_IN), .A3(
        REIP_REG_21__SCAN_IN), .A4(n5847), .ZN(n5821) );
  NAND3_X1 U5823 ( .A1(REIP_REG_24__SCAN_IN), .A2(REIP_REG_26__SCAN_IN), .A3(
        REIP_REG_25__SCAN_IN), .ZN(n4799) );
  NAND3_X1 U5824 ( .A1(REIP_REG_28__SCAN_IN), .A2(REIP_REG_27__SCAN_IN), .A3(
        n5801), .ZN(n5785) );
  NAND3_X1 U5825 ( .A1(REIP_REG_29__SCAN_IN), .A2(REIP_REG_30__SCAN_IN), .A3(
        n6983), .ZN(n4790) );
  OAI22_X1 U5826 ( .A1(n6274), .A2(n6236), .B1(n5785), .B2(n4790), .ZN(n4807)
         );
  INV_X1 U5827 ( .A(n6240), .ZN(n6256) );
  NAND2_X1 U5828 ( .A1(REIP_REG_29__SCAN_IN), .A2(REIP_REG_30__SCAN_IN), .ZN(
        n4801) );
  INV_X1 U5829 ( .A(REIP_REG_27__SCAN_IN), .ZN(n6972) );
  NOR2_X1 U5830 ( .A1(n6978), .A2(n6972), .ZN(n4800) );
  OR2_X1 U5831 ( .A1(n6523), .A2(n6903), .ZN(n4791) );
  NOR2_X1 U5832 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n7027) );
  AND3_X1 U5833 ( .A1(STATE2_REG_0__SCAN_IN), .A2(STATE2_REG_3__SCAN_IN), .A3(
        n7027), .ZN(n6889) );
  NOR2_X1 U5834 ( .A1(n4791), .A2(n6889), .ZN(n4792) );
  NAND2_X1 U5835 ( .A1(n6254), .A2(n6240), .ZN(n6270) );
  INV_X1 U5836 ( .A(REIP_REG_23__SCAN_IN), .ZN(n6967) );
  NAND2_X1 U5837 ( .A1(REIP_REG_22__SCAN_IN), .A2(REIP_REG_21__SCAN_IN), .ZN(
        n5846) );
  NOR2_X1 U5838 ( .A1(n6967), .A2(n5846), .ZN(n4798) );
  NOR3_X1 U5839 ( .A1(n4802), .A2(n6941), .A3(n4793), .ZN(n6152) );
  NAND4_X1 U5840 ( .A1(REIP_REG_9__SCAN_IN), .A2(REIP_REG_11__SCAN_IN), .A3(
        REIP_REG_10__SCAN_IN), .A4(n6152), .ZN(n4794) );
  NAND2_X1 U5841 ( .A1(n6270), .A2(n4794), .ZN(n6141) );
  INV_X1 U5842 ( .A(REIP_REG_14__SCAN_IN), .ZN(n6951) );
  OR3_X1 U5843 ( .A1(n6948), .A2(n6951), .A3(n6950), .ZN(n4795) );
  NAND2_X1 U5844 ( .A1(n6270), .A2(n4795), .ZN(n4796) );
  NAND2_X1 U5845 ( .A1(n6141), .A2(n4796), .ZN(n6121) );
  AOI21_X1 U5846 ( .B1(n4797), .B2(n6270), .A(n6121), .ZN(n5869) );
  OAI21_X1 U5847 ( .B1(n4798), .B2(n6240), .A(n5869), .ZN(n5836) );
  AOI21_X1 U5848 ( .B1(n4799), .B2(n6270), .A(n5836), .ZN(n5818) );
  OAI21_X1 U5849 ( .B1(n4800), .B2(n6240), .A(n5818), .ZN(n5788) );
  AOI21_X1 U5850 ( .B1(n6256), .B2(n4801), .A(n5788), .ZN(n5773) );
  NOR2_X2 U5851 ( .A1(n4802), .A2(n7000), .ZN(n6234) );
  OR2_X1 U5852 ( .A1(n6917), .A2(n4803), .ZN(n6883) );
  AND3_X1 U5853 ( .A1(n3567), .A2(n7022), .A3(n6883), .ZN(n5572) );
  AOI22_X1 U5854 ( .A1(PHYADDRPOINTER_REG_31__SCAN_IN), .A2(n6234), .B1(
        EBX_REG_31__SCAN_IN), .B2(n5572), .ZN(n4804) );
  NAND2_X1 U5855 ( .A1(n4809), .A2(n4808), .ZN(U2796) );
  NOR2_X1 U5856 ( .A1(n6776), .A2(STATE2_REG_1__SCAN_IN), .ZN(n7033) );
  AOI21_X1 U5857 ( .B1(n4810), .B2(MEMORYFETCH_REG_SCAN_IN), .A(n7033), .ZN(
        n4811) );
  NAND2_X1 U5858 ( .A1(n4815), .A2(n4811), .ZN(U2788) );
  INV_X1 U5859 ( .A(EAX_REG_25__SCAN_IN), .ZN(n6380) );
  NAND2_X1 U5860 ( .A1(n4812), .A2(n7024), .ZN(n4813) );
  NAND2_X1 U5861 ( .A1(n6450), .A2(DATAI_9_), .ZN(n4830) );
  NOR2_X1 U5862 ( .A1(n3567), .A2(n7024), .ZN(n4814) );
  NAND2_X1 U5863 ( .A1(n6464), .A2(UWORD_REG_9__SCAN_IN), .ZN(n4816) );
  OAI211_X1 U5864 ( .C1(n6380), .C2(n5764), .A(n4830), .B(n4816), .ZN(U2933)
         );
  INV_X1 U5865 ( .A(EAX_REG_6__SCAN_IN), .ZN(n6421) );
  NAND2_X1 U5866 ( .A1(n6450), .A2(DATAI_6_), .ZN(n4835) );
  NAND2_X1 U5867 ( .A1(n6464), .A2(LWORD_REG_6__SCAN_IN), .ZN(n4817) );
  OAI211_X1 U5868 ( .C1(n6421), .C2(n5764), .A(n4835), .B(n4817), .ZN(U2945)
         );
  INV_X1 U5869 ( .A(EAX_REG_4__SCAN_IN), .ZN(n6425) );
  INV_X1 U5870 ( .A(DATAI_4_), .ZN(n4818) );
  NOR2_X1 U5871 ( .A1(n6447), .A2(n4818), .ZN(n6443) );
  INV_X1 U5872 ( .A(n6443), .ZN(n4820) );
  NAND2_X1 U5873 ( .A1(n6464), .A2(LWORD_REG_4__SCAN_IN), .ZN(n4819) );
  OAI211_X1 U5874 ( .C1(n6425), .C2(n5764), .A(n4820), .B(n4819), .ZN(U2943)
         );
  INV_X1 U5875 ( .A(EAX_REG_3__SCAN_IN), .ZN(n6427) );
  NAND2_X1 U5876 ( .A1(n6450), .A2(DATAI_3_), .ZN(n4840) );
  NAND2_X1 U5877 ( .A1(n6464), .A2(LWORD_REG_3__SCAN_IN), .ZN(n4821) );
  OAI211_X1 U5878 ( .C1(n6427), .C2(n5764), .A(n4840), .B(n4821), .ZN(U2942)
         );
  INV_X1 U5879 ( .A(EAX_REG_1__SCAN_IN), .ZN(n6432) );
  INV_X1 U5880 ( .A(DATAI_1_), .ZN(n4822) );
  NOR2_X1 U5881 ( .A1(n6447), .A2(n4822), .ZN(n6438) );
  INV_X1 U5882 ( .A(n6438), .ZN(n4824) );
  NAND2_X1 U5883 ( .A1(n6464), .A2(LWORD_REG_1__SCAN_IN), .ZN(n4823) );
  OAI211_X1 U5884 ( .C1(n6432), .C2(n5764), .A(n4824), .B(n4823), .ZN(U2940)
         );
  INV_X1 U5885 ( .A(EAX_REG_0__SCAN_IN), .ZN(n6437) );
  NAND2_X1 U5886 ( .A1(n6450), .A2(DATAI_0_), .ZN(n4842) );
  NAND2_X1 U5887 ( .A1(n6464), .A2(LWORD_REG_0__SCAN_IN), .ZN(n4825) );
  OAI211_X1 U5888 ( .C1(n6437), .C2(n5764), .A(n4842), .B(n4825), .ZN(U2939)
         );
  NAND2_X1 U5889 ( .A1(n6450), .A2(DATAI_5_), .ZN(n4848) );
  NAND2_X1 U5890 ( .A1(n6464), .A2(LWORD_REG_5__SCAN_IN), .ZN(n4826) );
  OAI211_X1 U5891 ( .C1(n6423), .C2(n5764), .A(n4848), .B(n4826), .ZN(U2944)
         );
  NAND2_X1 U5892 ( .A1(n6450), .A2(DATAI_14_), .ZN(n4846) );
  NAND2_X1 U5893 ( .A1(n6464), .A2(LWORD_REG_14__SCAN_IN), .ZN(n4827) );
  OAI211_X1 U5894 ( .C1(n6402), .C2(n5764), .A(n4846), .B(n4827), .ZN(U2953)
         );
  NAND2_X1 U5895 ( .A1(n6450), .A2(DATAI_13_), .ZN(n4832) );
  NAND2_X1 U5896 ( .A1(n6464), .A2(LWORD_REG_13__SCAN_IN), .ZN(n4828) );
  OAI211_X1 U5897 ( .C1(n6404), .C2(n5764), .A(n4832), .B(n4828), .ZN(U2952)
         );
  INV_X1 U5898 ( .A(EAX_REG_9__SCAN_IN), .ZN(n6413) );
  NAND2_X1 U5899 ( .A1(n6464), .A2(LWORD_REG_9__SCAN_IN), .ZN(n4829) );
  OAI211_X1 U5900 ( .C1(n6413), .C2(n5764), .A(n4830), .B(n4829), .ZN(U2948)
         );
  INV_X1 U5901 ( .A(EAX_REG_29__SCAN_IN), .ZN(n6373) );
  NAND2_X1 U5902 ( .A1(n6464), .A2(UWORD_REG_13__SCAN_IN), .ZN(n4831) );
  OAI211_X1 U5903 ( .C1(n6373), .C2(n5764), .A(n4832), .B(n4831), .ZN(U2937)
         );
  INV_X1 U5904 ( .A(EAX_REG_7__SCAN_IN), .ZN(n6418) );
  NAND2_X1 U5905 ( .A1(n6450), .A2(DATAI_7_), .ZN(n4844) );
  NAND2_X1 U5906 ( .A1(n6464), .A2(LWORD_REG_7__SCAN_IN), .ZN(n4833) );
  OAI211_X1 U5907 ( .C1(n6418), .C2(n5764), .A(n4844), .B(n4833), .ZN(U2946)
         );
  INV_X1 U5908 ( .A(EAX_REG_22__SCAN_IN), .ZN(n6386) );
  NAND2_X1 U5909 ( .A1(n6464), .A2(UWORD_REG_6__SCAN_IN), .ZN(n4834) );
  OAI211_X1 U5910 ( .C1(n6386), .C2(n5764), .A(n4835), .B(n4834), .ZN(U2930)
         );
  INV_X1 U5911 ( .A(EAX_REG_27__SCAN_IN), .ZN(n6377) );
  INV_X1 U5912 ( .A(DATAI_11_), .ZN(n4836) );
  NOR2_X1 U5913 ( .A1(n6447), .A2(n4836), .ZN(n6460) );
  INV_X1 U5914 ( .A(n6460), .ZN(n4838) );
  NAND2_X1 U5915 ( .A1(n6464), .A2(UWORD_REG_11__SCAN_IN), .ZN(n4837) );
  OAI211_X1 U5916 ( .C1(n6377), .C2(n5764), .A(n4838), .B(n4837), .ZN(U2935)
         );
  INV_X1 U5917 ( .A(EAX_REG_19__SCAN_IN), .ZN(n6391) );
  NAND2_X1 U5918 ( .A1(n6464), .A2(UWORD_REG_3__SCAN_IN), .ZN(n4839) );
  OAI211_X1 U5919 ( .C1(n6391), .C2(n5764), .A(n4840), .B(n4839), .ZN(U2927)
         );
  INV_X1 U5920 ( .A(EAX_REG_16__SCAN_IN), .ZN(n6398) );
  NAND2_X1 U5921 ( .A1(n6464), .A2(UWORD_REG_0__SCAN_IN), .ZN(n4841) );
  OAI211_X1 U5922 ( .C1(n6398), .C2(n5764), .A(n4842), .B(n4841), .ZN(U2924)
         );
  INV_X1 U5923 ( .A(EAX_REG_23__SCAN_IN), .ZN(n6384) );
  NAND2_X1 U5924 ( .A1(n6464), .A2(UWORD_REG_7__SCAN_IN), .ZN(n4843) );
  OAI211_X1 U5925 ( .C1(n6384), .C2(n5764), .A(n4844), .B(n4843), .ZN(U2931)
         );
  INV_X1 U5926 ( .A(EAX_REG_30__SCAN_IN), .ZN(n6371) );
  NAND2_X1 U5927 ( .A1(n6464), .A2(UWORD_REG_14__SCAN_IN), .ZN(n4845) );
  OAI211_X1 U5928 ( .C1(n6371), .C2(n5764), .A(n4846), .B(n4845), .ZN(U2938)
         );
  INV_X1 U5929 ( .A(EAX_REG_21__SCAN_IN), .ZN(n6388) );
  NAND2_X1 U5930 ( .A1(n6464), .A2(UWORD_REG_5__SCAN_IN), .ZN(n4847) );
  OAI211_X1 U5931 ( .C1(n6388), .C2(n5764), .A(n4848), .B(n4847), .ZN(U2929)
         );
  OAI21_X1 U5932 ( .B1(n4849), .B2(INSTADDRPOINTER_REG_0__SCAN_IN), .A(n3603), 
        .ZN(n4863) );
  OAI21_X1 U5933 ( .B1(n6491), .B2(n4850), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n4856) );
  NAND2_X1 U5934 ( .A1(n4852), .A2(n4851), .ZN(n4853) );
  AND2_X1 U5935 ( .A1(n4854), .A2(n4853), .ZN(n6326) );
  AND2_X1 U5936 ( .A1(n6523), .A2(REIP_REG_0__SCAN_IN), .ZN(n4865) );
  AOI21_X1 U5937 ( .B1(n6326), .B2(n5989), .A(n4865), .ZN(n4855) );
  OAI211_X1 U5938 ( .C1(n4863), .C2(n6484), .A(n4856), .B(n4855), .ZN(U2986)
         );
  INV_X1 U5939 ( .A(LWORD_REG_15__SCAN_IN), .ZN(n4858) );
  AOI22_X1 U5940 ( .A1(n6450), .A2(DATAI_15_), .B1(n6465), .B2(
        EAX_REG_15__SCAN_IN), .ZN(n4857) );
  OAI21_X1 U5941 ( .B1(n6463), .B2(n4858), .A(n4857), .ZN(U2954) );
  AND2_X1 U5942 ( .A1(n5516), .A2(n4859), .ZN(n4868) );
  INV_X1 U5943 ( .A(n4860), .ZN(n4861) );
  AOI21_X1 U5944 ( .B1(n4862), .B2(n5596), .A(n4861), .ZN(n6322) );
  NOR2_X1 U5945 ( .A1(n6051), .A2(n4863), .ZN(n4864) );
  AOI211_X1 U5946 ( .C1(n6322), .C2(n6525), .A(n4865), .B(n4864), .ZN(n4867)
         );
  OAI211_X1 U5947 ( .C1(n4868), .C2(n5596), .A(n4867), .B(n4866), .ZN(U3018)
         );
  OAI21_X1 U5948 ( .B1(n6250), .B2(n4869), .A(n4603), .ZN(n4870) );
  OAI21_X1 U5949 ( .B1(n6851), .B2(n6917), .A(n4870), .ZN(n4871) );
  NAND3_X1 U5950 ( .A1(n6891), .A2(n7024), .A3(n4871), .ZN(n4874) );
  NAND3_X1 U5951 ( .A1(n4874), .A2(n4873), .A3(n4872), .ZN(n4878) );
  NAND2_X1 U5952 ( .A1(n6891), .A2(n5010), .ZN(n4877) );
  OR2_X1 U5953 ( .A1(n4613), .A2(n4875), .ZN(n4876) );
  NAND2_X1 U5954 ( .A1(n4877), .A2(n4876), .ZN(n5264) );
  NOR2_X1 U5955 ( .A1(n6891), .A2(n6872), .ZN(n5890) );
  OR3_X1 U5956 ( .A1(n4878), .A2(n5264), .A3(n5890), .ZN(n6845) );
  NOR2_X1 U5957 ( .A1(n7002), .A2(n6773), .ZN(n5765) );
  NAND2_X1 U5958 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n5765), .ZN(n6998) );
  INV_X1 U5959 ( .A(n6998), .ZN(n4879) );
  AOI22_X1 U5960 ( .A1(n5889), .A2(n6845), .B1(FLUSH_REG_SCAN_IN), .B2(n4879), 
        .ZN(n6072) );
  OAI21_X1 U5961 ( .B1(STATE2_REG_0__SCAN_IN), .B2(n7000), .A(n6072), .ZN(
        n7006) );
  INV_X1 U5962 ( .A(n7006), .ZN(n5601) );
  INV_X1 U5963 ( .A(n5753), .ZN(n5594) );
  INV_X1 U5964 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n4881) );
  AOI22_X1 U5965 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n4881), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n6531), .ZN(n5595) );
  NOR2_X1 U5966 ( .A1(n7002), .A2(n5596), .ZN(n4891) );
  INV_X1 U5967 ( .A(n4882), .ZN(n6259) );
  NAND2_X1 U5968 ( .A1(n4728), .A2(n4883), .ZN(n4884) );
  NOR2_X1 U5969 ( .A1(n4603), .A2(n4884), .ZN(n4885) );
  NAND3_X1 U5970 ( .A1(n4886), .A2(n4885), .A3(n4613), .ZN(n5020) );
  INV_X1 U5971 ( .A(n5020), .ZN(n6847) );
  NOR2_X1 U5972 ( .A1(n6851), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n5026)
         );
  INV_X1 U5973 ( .A(n5026), .ZN(n4890) );
  INV_X1 U5974 ( .A(n4887), .ZN(n5597) );
  INV_X1 U5975 ( .A(n4888), .ZN(n5037) );
  NAND3_X1 U5976 ( .A1(n6848), .A2(n5597), .A3(n5037), .ZN(n4889) );
  OAI211_X1 U5977 ( .C1(n6259), .C2(n6847), .A(n4890), .B(n4889), .ZN(n6854)
         );
  INV_X1 U5978 ( .A(n7008), .ZN(n5600) );
  AOI222_X1 U5979 ( .A1(n5594), .A2(n4880), .B1(n5595), .B2(n4891), .C1(n6854), 
        .C2(n5600), .ZN(n4893) );
  OAI21_X1 U5980 ( .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n5753), .A(n7006), 
        .ZN(n7004) );
  INV_X1 U5981 ( .A(n7004), .ZN(n4892) );
  OAI22_X1 U5982 ( .A1(n5601), .A2(n4893), .B1(n4892), .B2(n3291), .ZN(U3460)
         );
  XNOR2_X1 U5983 ( .A(n4894), .B(n4896), .ZN(n4937) );
  NAND2_X1 U5984 ( .A1(n4898), .A2(n4907), .ZN(n4909) );
  AND2_X1 U5985 ( .A1(n4909), .A2(n4899), .ZN(n4900) );
  NOR2_X1 U5986 ( .A1(n4897), .A2(n4900), .ZN(n6361) );
  INV_X1 U5987 ( .A(n6217), .ZN(n4902) );
  AOI22_X1 U5988 ( .A1(n6491), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .B1(n6523), 
        .B2(REIP_REG_4__SCAN_IN), .ZN(n4901) );
  OAI21_X1 U5989 ( .B1(n6490), .B2(n4902), .A(n4901), .ZN(n4903) );
  AOI21_X1 U5990 ( .B1(n6361), .B2(n5989), .A(n4903), .ZN(n4904) );
  OAI21_X1 U5991 ( .B1(n6484), .B2(n4937), .A(n4904), .ZN(U2982) );
  XNOR2_X1 U5992 ( .A(n4905), .B(n4906), .ZN(n4964) );
  NOR2_X1 U5993 ( .A1(n3179), .A2(n6931), .ZN(n4960) );
  OR2_X1 U5994 ( .A1(n4898), .A2(n4907), .ZN(n4908) );
  NAND2_X1 U5995 ( .A1(n4909), .A2(n4908), .ZN(n6364) );
  OAI22_X1 U5996 ( .A1(n6490), .A2(n6226), .B1(n6476), .B2(n6364), .ZN(n4910)
         );
  AOI211_X1 U5997 ( .C1(n6491), .C2(PHYADDRPOINTER_REG_3__SCAN_IN), .A(n4960), 
        .B(n4910), .ZN(n4911) );
  OAI21_X1 U5998 ( .B1(n4964), .B2(n6484), .A(n4911), .ZN(U2983) );
  NAND2_X1 U5999 ( .A1(n4913), .A2(n4912), .ZN(n4914) );
  XNOR2_X1 U6000 ( .A(n4915), .B(n4914), .ZN(n6485) );
  NOR2_X1 U6001 ( .A1(n6531), .A2(n4944), .ZN(n4917) );
  AOI22_X1 U6002 ( .A1(n4929), .A2(n6526), .B1(n5484), .B2(n4930), .ZN(n4949)
         );
  INV_X1 U6003 ( .A(n4949), .ZN(n4916) );
  MUX2_X1 U6004 ( .A(n4917), .B(n4916), .S(INSTADDRPOINTER_REG_2__SCAN_IN), 
        .Z(n4918) );
  INV_X1 U6005 ( .A(n4918), .ZN(n4926) );
  OAI21_X1 U6006 ( .B1(n5596), .B2(n4930), .A(n4931), .ZN(n4924) );
  NAND2_X1 U6007 ( .A1(n4920), .A2(n4919), .ZN(n4921) );
  NAND2_X1 U6008 ( .A1(n4957), .A2(n4921), .ZN(n6315) );
  INV_X1 U6009 ( .A(REIP_REG_2__SCAN_IN), .ZN(n4922) );
  OAI22_X1 U6010 ( .A1(n6512), .A2(n6315), .B1(n3179), .B2(n4922), .ZN(n4923)
         );
  AOI21_X1 U6011 ( .B1(n5497), .B2(n4924), .A(n4923), .ZN(n4925) );
  OAI211_X1 U6012 ( .C1(n6485), .C2(n6051), .A(n4926), .B(n4925), .ZN(U3016)
         );
  OAI21_X1 U6013 ( .B1(n4929), .B2(n4931), .A(n4949), .ZN(n4955) );
  OR2_X1 U6014 ( .A1(n4958), .A2(n4927), .ZN(n4928) );
  NAND2_X1 U6015 ( .A1(n4941), .A2(n4928), .ZN(n6312) );
  OAI22_X1 U6016 ( .A1(n6512), .A2(n6312), .B1(n6933), .B2(n3179), .ZN(n4935)
         );
  OAI21_X1 U6017 ( .B1(n4930), .B2(n4944), .A(n4929), .ZN(n5128) );
  AND2_X1 U6018 ( .A1(n4931), .A2(n5128), .ZN(n4954) );
  OAI211_X1 U6019 ( .C1(INSTADDRPOINTER_REG_4__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_3__SCAN_IN), .A(n4954), .B(n4932), .ZN(n4933) );
  INV_X1 U6020 ( .A(n4933), .ZN(n4934) );
  AOI211_X1 U6021 ( .C1(INSTADDRPOINTER_REG_4__SCAN_IN), .C2(n4955), .A(n4935), 
        .B(n4934), .ZN(n4936) );
  OAI21_X1 U6022 ( .B1(n6051), .B2(n4937), .A(n4936), .ZN(U3014) );
  XNOR2_X1 U6023 ( .A(n4938), .B(n4939), .ZN(n6478) );
  NAND2_X1 U6024 ( .A1(n4941), .A2(n4940), .ZN(n4942) );
  NAND2_X1 U6025 ( .A1(n5125), .A2(n4942), .ZN(n6309) );
  INV_X1 U6026 ( .A(n6309), .ZN(n6204) );
  INV_X1 U6027 ( .A(REIP_REG_5__SCAN_IN), .ZN(n6935) );
  NOR2_X1 U6028 ( .A1(n3179), .A2(n6935), .ZN(n6480) );
  INV_X1 U6029 ( .A(n4943), .ZN(n4945) );
  NOR3_X1 U6030 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n4945), .A3(n4944), 
        .ZN(n4946) );
  AOI211_X1 U6031 ( .C1(n6525), .C2(n6204), .A(n6480), .B(n4946), .ZN(n4952)
         );
  INV_X1 U6032 ( .A(n6530), .ZN(n5646) );
  NOR2_X1 U6033 ( .A1(n4948), .A2(n4947), .ZN(n5129) );
  OAI21_X1 U6034 ( .B1(n5646), .B2(n5129), .A(n4949), .ZN(n5132) );
  OAI21_X1 U6035 ( .B1(INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n4950), .A(n5132), 
        .ZN(n4951) );
  OAI211_X1 U6036 ( .C1(n6051), .C2(n6478), .A(n4952), .B(n4951), .ZN(U3013)
         );
  AOI22_X1 U6037 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n4955), .B1(n4954), 
        .B2(n4953), .ZN(n4963) );
  AND2_X1 U6038 ( .A1(n4957), .A2(n4956), .ZN(n4959) );
  OR2_X1 U6039 ( .A1(n4959), .A2(n4958), .ZN(n6313) );
  INV_X1 U6040 ( .A(n6313), .ZN(n4961) );
  AOI21_X1 U6041 ( .B1(n6525), .B2(n4961), .A(n4960), .ZN(n4962) );
  OAI211_X1 U6042 ( .C1(n4964), .C2(n6051), .A(n4963), .B(n4962), .ZN(U3015)
         );
  INV_X1 U6043 ( .A(n5042), .ZN(n4965) );
  INV_X1 U6044 ( .A(n5444), .ZN(n6837) );
  OAI21_X1 U6045 ( .B1(n6821), .B2(n6837), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n4970) );
  INV_X1 U6046 ( .A(n6776), .ZN(n6643) );
  AND2_X1 U6047 ( .A1(n4882), .A2(n3210), .ZN(n6607) );
  NAND2_X1 U6048 ( .A1(n6607), .A2(n6636), .ZN(n4976) );
  NAND3_X1 U6049 ( .A1(n4970), .A2(n6643), .A3(n4976), .ZN(n4975) );
  NOR2_X1 U6050 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5192), .ZN(n5442)
         );
  INV_X1 U6051 ( .A(n5442), .ZN(n4972) );
  INV_X1 U6052 ( .A(n6638), .ZN(n5055) );
  NAND2_X1 U6053 ( .A1(n5055), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n5285) );
  AOI21_X1 U6054 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n5285), .A(n6646), .ZN(
        n4971) );
  INV_X1 U6055 ( .A(n4971), .ZN(n5282) );
  AOI21_X1 U6056 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n4972), .A(n5282), .ZN(
        n4974) );
  INV_X1 U6057 ( .A(n4977), .ZN(n4973) );
  NAND2_X1 U6058 ( .A1(n4973), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6725) );
  INV_X1 U6059 ( .A(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4985) );
  NOR2_X2 U6060 ( .A1(n5276), .A2(n6646), .ZN(n6740) );
  OR2_X1 U6061 ( .A1(n4976), .A2(n6776), .ZN(n4979) );
  NAND2_X1 U6062 ( .A1(n4977), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6729) );
  OR2_X1 U6063 ( .A1(n6729), .A2(n5285), .ZN(n4978) );
  NAND2_X1 U6064 ( .A1(n4979), .A2(n4978), .ZN(n5446) );
  INV_X1 U6065 ( .A(DATAI_18_), .ZN(n4980) );
  NOR2_X1 U6066 ( .A1(n6476), .A2(n4980), .ZN(n6791) );
  INV_X1 U6067 ( .A(n6791), .ZN(n6696) );
  NAND2_X1 U6068 ( .A1(n5989), .A2(DATAI_26_), .ZN(n6657) );
  INV_X1 U6069 ( .A(n6657), .ZN(n6792) );
  NOR2_X2 U6070 ( .A1(n5322), .A2(n3426), .ZN(n6790) );
  AOI22_X1 U6071 ( .A1(n6792), .A2(n6821), .B1(n6790), .B2(n5442), .ZN(n4982)
         );
  OAI21_X1 U6072 ( .B1(n6696), .B2(n5444), .A(n4982), .ZN(n4983) );
  AOI21_X1 U6073 ( .B1(n6740), .B2(n5446), .A(n4983), .ZN(n4984) );
  OAI21_X1 U6074 ( .B1(n5449), .B2(n4985), .A(n4984), .ZN(U3134) );
  INV_X1 U6075 ( .A(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4992) );
  INV_X1 U6076 ( .A(DATAI_3_), .ZN(n6363) );
  NOR2_X2 U6077 ( .A1(n6363), .A2(n6646), .ZN(n6744) );
  INV_X1 U6078 ( .A(DATAI_19_), .ZN(n4986) );
  NOR2_X1 U6079 ( .A1(n6476), .A2(n4986), .ZN(n6798) );
  INV_X1 U6080 ( .A(n6798), .ZN(n6588) );
  INV_X1 U6081 ( .A(DATAI_27_), .ZN(n4987) );
  NOR2_X1 U6082 ( .A1(n6476), .A2(n4987), .ZN(n6797) );
  NOR2_X2 U6083 ( .A1(n5322), .A2(n4988), .ZN(n6796) );
  AOI22_X1 U6084 ( .A1(n6797), .A2(n6821), .B1(n6796), .B2(n5442), .ZN(n4989)
         );
  OAI21_X1 U6085 ( .B1(n6588), .B2(n5444), .A(n4989), .ZN(n4990) );
  AOI21_X1 U6086 ( .B1(n6744), .B2(n5446), .A(n4990), .ZN(n4991) );
  OAI21_X1 U6087 ( .B1(n5449), .B2(n4992), .A(n4991), .ZN(U3135) );
  INV_X1 U6088 ( .A(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n4997) );
  NOR2_X2 U6089 ( .A1(n4822), .A2(n6646), .ZN(n6736) );
  INV_X1 U6090 ( .A(DATAI_17_), .ZN(n4993) );
  NOR2_X1 U6091 ( .A1(n6476), .A2(n4993), .ZN(n6786) );
  INV_X1 U6092 ( .A(n6786), .ZN(n6693) );
  NAND2_X1 U6093 ( .A1(n5989), .A2(DATAI_25_), .ZN(n6654) );
  INV_X1 U6094 ( .A(n6654), .ZN(n6785) );
  NOR2_X2 U6095 ( .A1(n5322), .A2(n3714), .ZN(n6784) );
  AOI22_X1 U6096 ( .A1(n6785), .A2(n6821), .B1(n6784), .B2(n5442), .ZN(n4994)
         );
  OAI21_X1 U6097 ( .B1(n6693), .B2(n5444), .A(n4994), .ZN(n4995) );
  AOI21_X1 U6098 ( .B1(n6736), .B2(n5446), .A(n4995), .ZN(n4996) );
  OAI21_X1 U6099 ( .B1(n5449), .B2(n4997), .A(n4996), .ZN(U3133) );
  INV_X1 U6100 ( .A(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n5003) );
  INV_X1 U6101 ( .A(DATAI_5_), .ZN(n5272) );
  NOR2_X2 U6102 ( .A1(n5272), .A2(n6646), .ZN(n6752) );
  INV_X1 U6103 ( .A(DATAI_21_), .ZN(n4998) );
  NOR2_X1 U6104 ( .A1(n6476), .A2(n4998), .ZN(n6810) );
  INV_X1 U6105 ( .A(n6810), .ZN(n6594) );
  NAND2_X1 U6106 ( .A1(n5989), .A2(DATAI_29_), .ZN(n6705) );
  INV_X1 U6107 ( .A(n6705), .ZN(n6809) );
  NOR2_X2 U6108 ( .A1(n5322), .A2(n4999), .ZN(n6808) );
  AOI22_X1 U6109 ( .A1(n6809), .A2(n6821), .B1(n6808), .B2(n5442), .ZN(n5000)
         );
  OAI21_X1 U6110 ( .B1(n6594), .B2(n5444), .A(n5000), .ZN(n5001) );
  AOI21_X1 U6111 ( .B1(n6752), .B2(n5446), .A(n5001), .ZN(n5002) );
  OAI21_X1 U6112 ( .B1(n5449), .B2(n5003), .A(n5002), .ZN(U3137) );
  MUX2_X1 U6113 ( .A(n6845), .B(FLUSH_REG_SCAN_IN), .S(STATE2_REG_1__SCAN_IN), 
        .Z(n5007) );
  INV_X1 U6114 ( .A(n6573), .ZN(n6722) );
  OR2_X1 U6115 ( .A1(n5004), .A2(n6722), .ZN(n5005) );
  XNOR2_X1 U6116 ( .A(n5005), .B(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n6213)
         );
  NOR2_X1 U6117 ( .A1(n4613), .A2(STATE2_REG_1__SCAN_IN), .ZN(n5006) );
  NAND2_X1 U6118 ( .A1(n6213), .A2(n5006), .ZN(n6069) );
  OAI21_X1 U6119 ( .B1(n5007), .B2(n6070), .A(n6069), .ZN(n5038) );
  INV_X1 U6120 ( .A(n6845), .ZN(n6857) );
  NAND2_X1 U6121 ( .A1(n4887), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n5008) );
  NAND2_X1 U6122 ( .A1(n5008), .A2(n3739), .ZN(n5009) );
  NAND2_X1 U6123 ( .A1(n3557), .A2(n5009), .ZN(n5752) );
  NAND2_X1 U6124 ( .A1(n6636), .A2(n5020), .ZN(n5019) );
  INV_X1 U6125 ( .A(n5010), .ZN(n5011) );
  NAND2_X1 U6126 ( .A1(n6872), .A2(n5011), .ZN(n5023) );
  NAND2_X1 U6127 ( .A1(n5597), .A2(n5603), .ZN(n5014) );
  NAND2_X1 U6128 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n5012) );
  NOR2_X1 U6129 ( .A1(n6851), .A2(n5012), .ZN(n5013) );
  AOI21_X1 U6130 ( .B1(n5023), .B2(n5014), .A(n5013), .ZN(n5017) );
  NAND2_X1 U6131 ( .A1(n4887), .A2(n6851), .ZN(n5015) );
  AOI21_X1 U6132 ( .B1(n5015), .B2(n5603), .A(n5026), .ZN(n5016) );
  MUX2_X1 U6133 ( .A(n5017), .B(n5016), .S(INSTQUEUERD_ADDR_REG_3__SCAN_IN), 
        .Z(n5018) );
  OAI211_X1 U6134 ( .C1(n5021), .C2(n5752), .A(n5019), .B(n5018), .ZN(n6844)
         );
  NAND2_X1 U6135 ( .A1(n3210), .A2(n5020), .ZN(n5030) );
  INV_X1 U6136 ( .A(n5021), .ZN(n5024) );
  XNOR2_X1 U6137 ( .A(n4887), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n5022)
         );
  MUX2_X1 U6138 ( .A(n5024), .B(n5023), .S(n5022), .Z(n5028) );
  NOR2_X1 U6139 ( .A1(n6851), .A2(n3291), .ZN(n5025) );
  MUX2_X1 U6140 ( .A(n5026), .B(n5025), .S(n5603), .Z(n5027) );
  NOR2_X1 U6141 ( .A1(n5028), .A2(n5027), .ZN(n5029) );
  NAND2_X1 U6142 ( .A1(n5030), .A2(n5029), .ZN(n6846) );
  NAND3_X1 U6143 ( .A1(n6844), .A2(n7002), .A3(n6846), .ZN(n5035) );
  INV_X1 U6144 ( .A(FLUSH_REG_SCAN_IN), .ZN(n6083) );
  NAND2_X1 U6145 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6083), .ZN(n5031) );
  OAI21_X1 U6146 ( .B1(n6845), .B2(STATE2_REG_1__SCAN_IN), .A(n5031), .ZN(
        n5033) );
  NAND2_X1 U6147 ( .A1(n5033), .A2(n5032), .ZN(n5034) );
  OAI21_X1 U6148 ( .B1(n6857), .B2(n5035), .A(n5034), .ZN(n5036) );
  NOR2_X1 U6149 ( .A1(n5038), .A2(n5036), .ZN(n6880) );
  NOR2_X1 U6150 ( .A1(n5038), .A2(n5037), .ZN(n5039) );
  NOR2_X1 U6151 ( .A1(n6880), .A2(n5039), .ZN(n5048) );
  NOR2_X1 U6152 ( .A1(n5048), .A2(FLUSH_REG_SCAN_IN), .ZN(n5040) );
  OAI21_X1 U6153 ( .B1(n5040), .B2(n6998), .A(n6646), .ZN(n6535) );
  INV_X1 U6154 ( .A(n6720), .ZN(n5041) );
  NOR2_X1 U6155 ( .A1(n5041), .A2(n6081), .ZN(n6768) );
  NAND2_X1 U6156 ( .A1(n3798), .A2(n6537), .ZN(n6676) );
  INV_X1 U6157 ( .A(n6676), .ZN(n6679) );
  NOR2_X1 U6158 ( .A1(n6768), .A2(n6679), .ZN(n6538) );
  NOR2_X1 U6159 ( .A1(n6537), .A2(n5042), .ZN(n6615) );
  NAND2_X1 U6160 ( .A1(n6678), .A2(n6615), .ZN(n6605) );
  AOI21_X1 U6161 ( .B1(n6538), .B2(n6605), .A(n6776), .ZN(n5045) );
  INV_X1 U6162 ( .A(n3798), .ZN(n5043) );
  OR2_X1 U6163 ( .A1(n6776), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5186) );
  INV_X1 U6164 ( .A(n6636), .ZN(n6731) );
  AND2_X1 U6165 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n7000), .ZN(n5748) );
  OAI22_X1 U6166 ( .A1(n5043), .A2(n5186), .B1(n6731), .B2(n5748), .ZN(n5044)
         );
  OAI21_X1 U6167 ( .B1(n5045), .B2(n5044), .A(n6535), .ZN(n5046) );
  OAI21_X1 U6168 ( .B1(n6535), .B2(n6864), .A(n5046), .ZN(U3462) );
  INV_X1 U6169 ( .A(n5765), .ZN(n5047) );
  NOR2_X1 U6170 ( .A1(n5048), .A2(n5047), .ZN(n6890) );
  OAI22_X1 U6171 ( .A1(n6719), .A2(n6776), .B1(n3776), .B2(n5748), .ZN(n5049)
         );
  OAI21_X1 U6172 ( .B1(n6890), .B2(n5049), .A(n6535), .ZN(n5050) );
  OAI21_X1 U6173 ( .B1(n6535), .B2(n6769), .A(n5050), .ZN(U3465) );
  NAND2_X1 U6174 ( .A1(n5077), .A2(n6537), .ZN(n5051) );
  NAND2_X1 U6175 ( .A1(n5104), .A2(n3774), .ZN(n5327) );
  NAND2_X1 U6176 ( .A1(n6537), .A2(n3768), .ZN(n5052) );
  INV_X1 U6177 ( .A(n5076), .ZN(n5053) );
  NAND2_X1 U6178 ( .A1(n5053), .A2(n6719), .ZN(n5326) );
  INV_X1 U6179 ( .A(n5186), .ZN(n6723) );
  AOI21_X1 U6180 ( .B1(n5327), .B2(n5326), .A(n6723), .ZN(n5054) );
  OR2_X1 U6181 ( .A1(n3210), .A2(n6259), .ZN(n5279) );
  NOR2_X1 U6182 ( .A1(n5279), .A2(n6636), .ZN(n6540) );
  OAI21_X1 U6183 ( .B1(n5054), .B2(n6540), .A(n7000), .ZN(n5058) );
  NAND2_X1 U6184 ( .A1(n5281), .A2(n6864), .ZN(n6543) );
  NOR2_X1 U6185 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6543), .ZN(n5323)
         );
  INV_X1 U6186 ( .A(n5323), .ZN(n5057) );
  NAND2_X1 U6187 ( .A1(n5055), .A2(n6864), .ZN(n6571) );
  AOI21_X1 U6188 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6571), .A(n6646), .ZN(
        n5056) );
  INV_X1 U6189 ( .A(n5056), .ZN(n6575) );
  INV_X1 U6190 ( .A(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n5063) );
  INV_X1 U6191 ( .A(n6540), .ZN(n5059) );
  OAI22_X1 U6192 ( .A1(n5059), .A2(n6776), .B1(n6725), .B2(n6571), .ZN(n5324)
         );
  AOI22_X1 U6193 ( .A1(n6752), .A2(n5324), .B1(n6808), .B2(n5323), .ZN(n5062)
         );
  OAI22_X1 U6194 ( .A1(n6705), .A2(n5327), .B1(n5326), .B2(n6594), .ZN(n5060)
         );
  INV_X1 U6195 ( .A(n5060), .ZN(n5061) );
  OAI211_X1 U6196 ( .C1(n5331), .C2(n5063), .A(n5062), .B(n5061), .ZN(U3041)
         );
  INV_X1 U6197 ( .A(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n5067) );
  AOI22_X1 U6198 ( .A1(n6744), .A2(n5324), .B1(n6796), .B2(n5323), .ZN(n5066)
         );
  INV_X1 U6199 ( .A(n6797), .ZN(n6699) );
  OAI22_X1 U6200 ( .A1(n6699), .A2(n5327), .B1(n5326), .B2(n6588), .ZN(n5064)
         );
  INV_X1 U6201 ( .A(n5064), .ZN(n5065) );
  OAI211_X1 U6202 ( .C1(n5331), .C2(n5067), .A(n5066), .B(n5065), .ZN(U3039)
         );
  INV_X1 U6203 ( .A(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n5071) );
  AOI22_X1 U6204 ( .A1(n6740), .A2(n5324), .B1(n6790), .B2(n5323), .ZN(n5070)
         );
  OAI22_X1 U6205 ( .A1(n6657), .A2(n5327), .B1(n5326), .B2(n6696), .ZN(n5068)
         );
  INV_X1 U6206 ( .A(n5068), .ZN(n5069) );
  OAI211_X1 U6207 ( .C1(n5331), .C2(n5071), .A(n5070), .B(n5069), .ZN(U3038)
         );
  INV_X1 U6208 ( .A(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n5075) );
  AOI22_X1 U6209 ( .A1(n6736), .A2(n5324), .B1(n6784), .B2(n5323), .ZN(n5074)
         );
  OAI22_X1 U6210 ( .A1(n6654), .A2(n5327), .B1(n5326), .B2(n6693), .ZN(n5072)
         );
  INV_X1 U6211 ( .A(n5072), .ZN(n5073) );
  OAI211_X1 U6212 ( .C1(n5331), .C2(n5075), .A(n5074), .B(n5073), .ZN(U3037)
         );
  NAND2_X1 U6213 ( .A1(n6770), .A2(n6643), .ZN(n6732) );
  NAND2_X1 U6214 ( .A1(n6637), .A2(n6638), .ZN(n5109) );
  OAI22_X1 U6215 ( .A1(n6732), .A2(n6636), .B1(n5109), .B2(n6729), .ZN(n5437)
         );
  INV_X1 U6216 ( .A(n6784), .ZN(n5204) );
  NAND3_X1 U6217 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n6859), .A3(n6864), .ZN(n5142) );
  NOR2_X1 U6218 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5142), .ZN(n5080)
         );
  INV_X1 U6219 ( .A(n5080), .ZN(n5434) );
  NAND2_X1 U6220 ( .A1(n5145), .A2(n6719), .ZN(n5452) );
  OAI22_X1 U6221 ( .A1(n5204), .A2(n5434), .B1(n5452), .B2(n6693), .ZN(n5078)
         );
  AOI21_X1 U6222 ( .B1(n6736), .B2(n5437), .A(n5078), .ZN(n5085) );
  INV_X1 U6223 ( .A(n6770), .ZN(n6721) );
  AOI21_X1 U6224 ( .B1(n5145), .B2(STATEBS16_REG_SCAN_IN), .A(n6776), .ZN(
        n5141) );
  NAND2_X1 U6225 ( .A1(n6563), .A2(n5186), .ZN(n5079) );
  OAI211_X1 U6226 ( .C1(n6573), .C2(n6721), .A(n5141), .B(n5079), .ZN(n5083)
         );
  AOI21_X1 U6227 ( .B1(n5109), .B2(STATE2_REG_2__SCAN_IN), .A(n6646), .ZN(
        n5106) );
  OAI21_X1 U6228 ( .B1(n7000), .B2(n5080), .A(n5106), .ZN(n5081) );
  INV_X1 U6229 ( .A(n5081), .ZN(n5082) );
  NAND3_X1 U6230 ( .A1(n5083), .A2(n5082), .A3(n6725), .ZN(n5438) );
  NAND2_X1 U6231 ( .A1(n5438), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n5084) );
  OAI211_X1 U6232 ( .C1(n5441), .C2(n6654), .A(n5085), .B(n5084), .ZN(U3053)
         );
  INV_X1 U6233 ( .A(n6808), .ZN(n5209) );
  OAI22_X1 U6234 ( .A1(n5209), .A2(n5434), .B1(n5452), .B2(n6594), .ZN(n5086)
         );
  AOI21_X1 U6235 ( .B1(n6752), .B2(n5437), .A(n5086), .ZN(n5088) );
  NAND2_X1 U6236 ( .A1(n5438), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n5087) );
  OAI211_X1 U6237 ( .C1(n5441), .C2(n6705), .A(n5088), .B(n5087), .ZN(U3057)
         );
  INV_X1 U6238 ( .A(n6790), .ZN(n5199) );
  OAI22_X1 U6239 ( .A1(n5199), .A2(n5434), .B1(n5452), .B2(n6696), .ZN(n5089)
         );
  AOI21_X1 U6240 ( .B1(n6740), .B2(n5437), .A(n5089), .ZN(n5091) );
  NAND2_X1 U6241 ( .A1(n5438), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n5090) );
  OAI211_X1 U6242 ( .C1(n5441), .C2(n6657), .A(n5091), .B(n5090), .ZN(U3054)
         );
  INV_X1 U6243 ( .A(n6796), .ZN(n5194) );
  OAI22_X1 U6244 ( .A1(n5194), .A2(n5434), .B1(n5452), .B2(n6588), .ZN(n5092)
         );
  AOI21_X1 U6245 ( .B1(n6744), .B2(n5437), .A(n5092), .ZN(n5094) );
  NAND2_X1 U6246 ( .A1(n5438), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n5093) );
  OAI211_X1 U6247 ( .C1(n5441), .C2(n6699), .A(n5094), .B(n5093), .ZN(U3055)
         );
  XNOR2_X1 U6248 ( .A(n5095), .B(n5097), .ZN(n5134) );
  OR2_X1 U6249 ( .A1(n5270), .A2(n5099), .ZN(n5255) );
  NAND2_X1 U6250 ( .A1(n5270), .A2(n5099), .ZN(n5100) );
  AND2_X1 U6251 ( .A1(n5255), .A2(n5100), .ZN(n6306) );
  NAND2_X1 U6252 ( .A1(n6498), .A2(n6195), .ZN(n5101) );
  NAND2_X1 U6253 ( .A1(n6523), .A2(REIP_REG_6__SCAN_IN), .ZN(n5127) );
  OAI211_X1 U6254 ( .C1(n5640), .C2(n6192), .A(n5101), .B(n5127), .ZN(n5102)
         );
  AOI21_X1 U6255 ( .B1(n6306), .B2(n5989), .A(n5102), .ZN(n5103) );
  OAI21_X1 U6256 ( .B1(n5134), .B2(n6484), .A(n5103), .ZN(U2980) );
  NAND2_X1 U6257 ( .A1(n5187), .A2(n3774), .ZN(n6835) );
  AOI21_X1 U6258 ( .B1(n5433), .B2(n6835), .A(n6081), .ZN(n5105) );
  OR2_X1 U6259 ( .A1(n3210), .A2(n4882), .ZN(n6645) );
  NOR2_X1 U6260 ( .A1(n6645), .A2(n6636), .ZN(n5338) );
  NOR3_X1 U6261 ( .A1(n5105), .A2(n5338), .A3(n6776), .ZN(n5108) );
  NAND3_X1 U6262 ( .A1(n5161), .A2(n6859), .A3(n6864), .ZN(n5341) );
  NOR2_X1 U6263 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5341), .ZN(n5111)
         );
  OAI211_X1 U6264 ( .C1(n7000), .C2(n5111), .A(n6729), .B(n5106), .ZN(n5107)
         );
  NAND2_X1 U6265 ( .A1(n5427), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n5114) );
  INV_X1 U6266 ( .A(n5338), .ZN(n5110) );
  OAI22_X1 U6267 ( .A1(n5110), .A2(n6776), .B1(n6725), .B2(n5109), .ZN(n5430)
         );
  INV_X1 U6268 ( .A(n5111), .ZN(n5428) );
  OAI22_X1 U6269 ( .A1(n5194), .A2(n5428), .B1(n6699), .B2(n6835), .ZN(n5112)
         );
  AOI21_X1 U6270 ( .B1(n6744), .B2(n5430), .A(n5112), .ZN(n5113) );
  OAI211_X1 U6271 ( .C1(n5433), .C2(n6588), .A(n5114), .B(n5113), .ZN(U3023)
         );
  NAND2_X1 U6272 ( .A1(n5427), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n5117) );
  OAI22_X1 U6273 ( .A1(n5199), .A2(n5428), .B1(n6657), .B2(n6835), .ZN(n5115)
         );
  AOI21_X1 U6274 ( .B1(n6740), .B2(n5430), .A(n5115), .ZN(n5116) );
  OAI211_X1 U6275 ( .C1(n5433), .C2(n6696), .A(n5117), .B(n5116), .ZN(U3022)
         );
  NAND2_X1 U6276 ( .A1(n5427), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n5120) );
  OAI22_X1 U6277 ( .A1(n5209), .A2(n5428), .B1(n6705), .B2(n6835), .ZN(n5118)
         );
  AOI21_X1 U6278 ( .B1(n6752), .B2(n5430), .A(n5118), .ZN(n5119) );
  OAI211_X1 U6279 ( .C1(n5433), .C2(n6594), .A(n5120), .B(n5119), .ZN(U3025)
         );
  NAND2_X1 U6280 ( .A1(n5427), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n5123) );
  OAI22_X1 U6281 ( .A1(n5204), .A2(n5428), .B1(n6654), .B2(n6835), .ZN(n5121)
         );
  AOI21_X1 U6282 ( .B1(n6736), .B2(n5430), .A(n5121), .ZN(n5122) );
  OAI211_X1 U6283 ( .C1(n5433), .C2(n6693), .A(n5123), .B(n5122), .ZN(U3021)
         );
  NAND2_X1 U6284 ( .A1(n5125), .A2(n5124), .ZN(n5126) );
  NAND2_X1 U6285 ( .A1(n6179), .A2(n5126), .ZN(n6307) );
  OAI21_X1 U6286 ( .B1(n6512), .B2(n6307), .A(n5127), .ZN(n5131) );
  NAND2_X1 U6287 ( .A1(n5129), .A2(n5128), .ZN(n5244) );
  NOR2_X1 U6288 ( .A1(n5244), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n5130)
         );
  AOI211_X1 U6289 ( .C1(n5132), .C2(INSTADDRPOINTER_REG_6__SCAN_IN), .A(n5131), 
        .B(n5130), .ZN(n5133) );
  OAI21_X1 U6290 ( .B1(n6051), .B2(n5134), .A(n5133), .ZN(U3012) );
  INV_X1 U6291 ( .A(n6646), .ZN(n5321) );
  NAND2_X1 U6292 ( .A1(DATAI_6_), .A2(n5321), .ZN(n6819) );
  NOR2_X2 U6293 ( .A1(n5322), .A2(n5261), .ZN(n6814) );
  AOI22_X1 U6294 ( .A1(n6756), .A2(n5324), .B1(n6814), .B2(n5323), .ZN(n5138)
         );
  NOR2_X1 U6295 ( .A1(n6476), .A2(n4566), .ZN(n6815) );
  INV_X1 U6296 ( .A(n6815), .ZN(n6709) );
  INV_X1 U6297 ( .A(DATAI_22_), .ZN(n5135) );
  NOR2_X1 U6298 ( .A1(n6476), .A2(n5135), .ZN(n6816) );
  INV_X1 U6299 ( .A(n6816), .ZN(n6597) );
  OAI22_X1 U6300 ( .A1(n6709), .A2(n5327), .B1(n5326), .B2(n6597), .ZN(n5136)
         );
  INV_X1 U6301 ( .A(n5136), .ZN(n5137) );
  OAI211_X1 U6302 ( .C1(n5331), .C2(n4563), .A(n5138), .B(n5137), .ZN(U3042)
         );
  NOR2_X1 U6303 ( .A1(n3776), .A2(n6573), .ZN(n6606) );
  NOR2_X1 U6304 ( .A1(n6769), .A2(n5142), .ZN(n5450) );
  AOI21_X1 U6305 ( .B1(n6770), .B2(n6606), .A(n5450), .ZN(n5143) );
  INV_X1 U6306 ( .A(n5142), .ZN(n5139) );
  OAI21_X1 U6307 ( .B1(n6643), .B2(n5139), .A(n6780), .ZN(n5140) );
  AOI21_X1 U6308 ( .B1(n5141), .B2(n5143), .A(n5140), .ZN(n5457) );
  INV_X1 U6309 ( .A(n5141), .ZN(n5144) );
  OAI22_X1 U6310 ( .A1(n5144), .A2(n5143), .B1(n5142), .B2(n6773), .ZN(n5454)
         );
  AOI22_X1 U6311 ( .A1(n6600), .A2(n6810), .B1(n6808), .B2(n5450), .ZN(n5146)
         );
  OAI21_X1 U6312 ( .B1(n6705), .B2(n5452), .A(n5146), .ZN(n5147) );
  AOI21_X1 U6313 ( .B1(n5454), .B2(n6752), .A(n5147), .ZN(n5148) );
  OAI21_X1 U6314 ( .B1(n5457), .B2(n4457), .A(n5148), .ZN(U3065) );
  AOI22_X1 U6315 ( .A1(n6600), .A2(n6786), .B1(n6784), .B2(n5450), .ZN(n5149)
         );
  OAI21_X1 U6316 ( .B1(n6654), .B2(n5452), .A(n5149), .ZN(n5150) );
  AOI21_X1 U6317 ( .B1(n5454), .B2(n6736), .A(n5150), .ZN(n5151) );
  OAI21_X1 U6318 ( .B1(n5457), .B2(n4561), .A(n5151), .ZN(U3061) );
  INV_X1 U6319 ( .A(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n5155) );
  AOI22_X1 U6320 ( .A1(n6600), .A2(n6798), .B1(n6796), .B2(n5450), .ZN(n5152)
         );
  OAI21_X1 U6321 ( .B1(n6699), .B2(n5452), .A(n5152), .ZN(n5153) );
  AOI21_X1 U6322 ( .B1(n5454), .B2(n6744), .A(n5153), .ZN(n5154) );
  OAI21_X1 U6323 ( .B1(n5457), .B2(n5155), .A(n5154), .ZN(U3063) );
  INV_X1 U6324 ( .A(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n5159) );
  AOI22_X1 U6325 ( .A1(n6600), .A2(n6791), .B1(n6790), .B2(n5450), .ZN(n5156)
         );
  OAI21_X1 U6326 ( .B1(n6657), .B2(n5452), .A(n5156), .ZN(n5157) );
  AOI21_X1 U6327 ( .B1(n5454), .B2(n6740), .A(n5157), .ZN(n5158) );
  OAI21_X1 U6328 ( .B1(n5457), .B2(n5159), .A(n5158), .ZN(U3062) );
  INV_X1 U6329 ( .A(n5167), .ZN(n5160) );
  OAI21_X1 U6330 ( .B1(n5167), .B2(n6081), .A(n6643), .ZN(n5166) );
  AND2_X1 U6331 ( .A1(n6636), .A2(n6681), .ZN(n6771) );
  INV_X1 U6332 ( .A(n6645), .ZN(n5162) );
  NAND3_X1 U6333 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n5161), .A3(n6859), .ZN(n6641) );
  NOR2_X1 U6334 ( .A1(n6769), .A2(n6641), .ZN(n5377) );
  AOI21_X1 U6335 ( .B1(n6771), .B2(n5162), .A(n5377), .ZN(n5165) );
  INV_X1 U6336 ( .A(n5165), .ZN(n5164) );
  NAND2_X1 U6337 ( .A1(n6776), .A2(n6641), .ZN(n5163) );
  OAI211_X1 U6338 ( .C1(n5166), .C2(n5164), .A(n6780), .B(n5163), .ZN(n5376)
         );
  OAI22_X1 U6339 ( .A1(n5166), .A2(n5165), .B1(n6773), .B2(n6641), .ZN(n5375)
         );
  AOI22_X1 U6340 ( .A1(INSTQUEUE_REG_9__3__SCAN_IN), .A2(n5376), .B1(n6744), 
        .B2(n5375), .ZN(n5169) );
  NOR2_X2 U6341 ( .A1(n5167), .A2(n3774), .ZN(n6668) );
  AOI22_X1 U6342 ( .A1(n6668), .A2(n6797), .B1(n5377), .B2(n6796), .ZN(n5168)
         );
  OAI211_X1 U6343 ( .C1(n5416), .C2(n6588), .A(n5169), .B(n5168), .ZN(U3095)
         );
  AOI22_X1 U6344 ( .A1(INSTQUEUE_REG_9__6__SCAN_IN), .A2(n5376), .B1(n6756), 
        .B2(n5375), .ZN(n5171) );
  AOI22_X1 U6345 ( .A1(n6668), .A2(n6815), .B1(n5377), .B2(n6814), .ZN(n5170)
         );
  OAI211_X1 U6346 ( .C1(n5416), .C2(n6597), .A(n5171), .B(n5170), .ZN(U3098)
         );
  AOI22_X1 U6347 ( .A1(INSTQUEUE_REG_9__2__SCAN_IN), .A2(n5376), .B1(n6740), 
        .B2(n5375), .ZN(n5173) );
  AOI22_X1 U6348 ( .A1(n6668), .A2(n6792), .B1(n5377), .B2(n6790), .ZN(n5172)
         );
  OAI211_X1 U6349 ( .C1(n5416), .C2(n6696), .A(n5173), .B(n5172), .ZN(U3094)
         );
  AOI22_X1 U6350 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(n5376), .B1(n6736), 
        .B2(n5375), .ZN(n5175) );
  AOI22_X1 U6351 ( .A1(n6668), .A2(n6785), .B1(n5377), .B2(n6784), .ZN(n5174)
         );
  OAI211_X1 U6352 ( .C1(n5416), .C2(n6693), .A(n5175), .B(n5174), .ZN(U3093)
         );
  AOI22_X1 U6353 ( .A1(INSTQUEUE_REG_9__5__SCAN_IN), .A2(n5376), .B1(n6752), 
        .B2(n5375), .ZN(n5177) );
  AOI22_X1 U6354 ( .A1(n6668), .A2(n6809), .B1(n5377), .B2(n6808), .ZN(n5176)
         );
  OAI211_X1 U6355 ( .C1(n5416), .C2(n6594), .A(n5177), .B(n5176), .ZN(U3097)
         );
  INV_X1 U6356 ( .A(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n5181) );
  AOI22_X1 U6357 ( .A1(n6815), .A2(n6821), .B1(n6814), .B2(n5442), .ZN(n5178)
         );
  OAI21_X1 U6358 ( .B1(n6597), .B2(n5444), .A(n5178), .ZN(n5179) );
  AOI21_X1 U6359 ( .B1(n6756), .B2(n5446), .A(n5179), .ZN(n5180) );
  OAI21_X1 U6360 ( .B1(n5449), .B2(n5181), .A(n5180), .ZN(U3138) );
  INV_X1 U6361 ( .A(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n5185) );
  AOI22_X1 U6362 ( .A1(n6600), .A2(n6816), .B1(n6814), .B2(n5450), .ZN(n5182)
         );
  OAI21_X1 U6363 ( .B1(n6709), .B2(n5452), .A(n5182), .ZN(n5183) );
  AOI21_X1 U6364 ( .B1(n5454), .B2(n6756), .A(n5183), .ZN(n5184) );
  OAI21_X1 U6365 ( .B1(n5457), .B2(n5185), .A(n5184), .ZN(U3066) );
  OAI21_X1 U6366 ( .B1(n5187), .B2(n6476), .A(n5186), .ZN(n5191) );
  AOI21_X1 U6367 ( .B1(n6771), .B2(n6607), .A(n6834), .ZN(n5193) );
  INV_X1 U6368 ( .A(n6780), .ZN(n5190) );
  NOR2_X1 U6369 ( .A1(n6643), .A2(n5188), .ZN(n5189) );
  AOI211_X2 U6370 ( .C1(n5191), .C2(n5193), .A(n5190), .B(n5189), .ZN(n6843)
         );
  INV_X1 U6371 ( .A(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n5198) );
  OAI22_X1 U6372 ( .A1(n5193), .A2(n6776), .B1(n5192), .B2(n6773), .ZN(n6831)
         );
  NOR2_X1 U6373 ( .A1(n5444), .A2(n6699), .ZN(n5196) );
  OAI22_X1 U6374 ( .A1(n5194), .A2(n5422), .B1(n6588), .B2(n6835), .ZN(n5195)
         );
  AOI211_X1 U6375 ( .C1(n6744), .C2(n6831), .A(n5196), .B(n5195), .ZN(n5197)
         );
  OAI21_X1 U6376 ( .B1(n6843), .B2(n5198), .A(n5197), .ZN(U3143) );
  INV_X1 U6377 ( .A(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n5203) );
  NOR2_X1 U6378 ( .A1(n5444), .A2(n6657), .ZN(n5201) );
  OAI22_X1 U6379 ( .A1(n5199), .A2(n5422), .B1(n6696), .B2(n6835), .ZN(n5200)
         );
  AOI211_X1 U6380 ( .C1(n6740), .C2(n6831), .A(n5201), .B(n5200), .ZN(n5202)
         );
  OAI21_X1 U6381 ( .B1(n6843), .B2(n5203), .A(n5202), .ZN(U3142) );
  INV_X1 U6382 ( .A(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n5208) );
  NOR2_X1 U6383 ( .A1(n5444), .A2(n6654), .ZN(n5206) );
  OAI22_X1 U6384 ( .A1(n5204), .A2(n5422), .B1(n6693), .B2(n6835), .ZN(n5205)
         );
  AOI211_X1 U6385 ( .C1(n6736), .C2(n6831), .A(n5206), .B(n5205), .ZN(n5207)
         );
  OAI21_X1 U6386 ( .B1(n6843), .B2(n5208), .A(n5207), .ZN(U3141) );
  INV_X1 U6387 ( .A(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n5213) );
  NOR2_X1 U6388 ( .A1(n5444), .A2(n6705), .ZN(n5211) );
  OAI22_X1 U6389 ( .A1(n5209), .A2(n5422), .B1(n6594), .B2(n6835), .ZN(n5210)
         );
  AOI211_X1 U6390 ( .C1(n6752), .C2(n6831), .A(n5211), .B(n5210), .ZN(n5212)
         );
  OAI21_X1 U6391 ( .B1(n6843), .B2(n5213), .A(n5212), .ZN(U3145) );
  INV_X1 U6392 ( .A(DATAI_23_), .ZN(n5214) );
  NOR2_X1 U6393 ( .A1(n6476), .A2(n5214), .ZN(n6820) );
  INV_X1 U6394 ( .A(n6820), .ZN(n6717) );
  INV_X1 U6395 ( .A(DATAI_7_), .ZN(n5269) );
  NOR2_X2 U6396 ( .A1(n5269), .A2(n6646), .ZN(n6762) );
  AOI22_X1 U6397 ( .A1(INSTQUEUE_REG_9__7__SCAN_IN), .A2(n5376), .B1(n6762), 
        .B2(n5375), .ZN(n5218) );
  INV_X1 U6398 ( .A(DATAI_31_), .ZN(n5215) );
  NOR2_X1 U6399 ( .A1(n6476), .A2(n5215), .ZN(n6825) );
  NOR2_X2 U6400 ( .A1(n5322), .A2(n5216), .ZN(n6823) );
  AOI22_X1 U6401 ( .A1(n6668), .A2(n6825), .B1(n5377), .B2(n6823), .ZN(n5217)
         );
  OAI211_X1 U6402 ( .C1(n5416), .C2(n6717), .A(n5218), .B(n5217), .ZN(U3099)
         );
  INV_X1 U6403 ( .A(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n5222) );
  AOI22_X1 U6404 ( .A1(n6762), .A2(n5324), .B1(n6823), .B2(n5323), .ZN(n5221)
         );
  INV_X1 U6405 ( .A(n6825), .ZN(n6673) );
  OAI22_X1 U6406 ( .A1(n6673), .A2(n5327), .B1(n5326), .B2(n6717), .ZN(n5219)
         );
  INV_X1 U6407 ( .A(n5219), .ZN(n5220) );
  OAI211_X1 U6408 ( .C1(n5331), .C2(n5222), .A(n5221), .B(n5220), .ZN(U3043)
         );
  INV_X1 U6409 ( .A(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n5226) );
  NOR2_X1 U6410 ( .A1(n5444), .A2(n6709), .ZN(n5224) );
  INV_X1 U6411 ( .A(n6814), .ZN(n5230) );
  OAI22_X1 U6412 ( .A1(n5230), .A2(n5422), .B1(n6597), .B2(n6835), .ZN(n5223)
         );
  AOI211_X1 U6413 ( .C1(n6756), .C2(n6831), .A(n5224), .B(n5223), .ZN(n5225)
         );
  OAI21_X1 U6414 ( .B1(n6843), .B2(n5226), .A(n5225), .ZN(U3146) );
  NAND2_X1 U6415 ( .A1(n5427), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n5229) );
  OAI22_X1 U6416 ( .A1(n5230), .A2(n5428), .B1(n6709), .B2(n6835), .ZN(n5227)
         );
  AOI21_X1 U6417 ( .B1(n6756), .B2(n5430), .A(n5227), .ZN(n5228) );
  OAI211_X1 U6418 ( .C1(n5433), .C2(n6597), .A(n5229), .B(n5228), .ZN(U3026)
         );
  OAI22_X1 U6419 ( .A1(n5230), .A2(n5434), .B1(n5452), .B2(n6597), .ZN(n5231)
         );
  AOI21_X1 U6420 ( .B1(n6756), .B2(n5437), .A(n5231), .ZN(n5233) );
  NAND2_X1 U6421 ( .A1(n5438), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n5232) );
  OAI211_X1 U6422 ( .C1(n5441), .C2(n6709), .A(n5233), .B(n5232), .ZN(U3058)
         );
  INV_X1 U6423 ( .A(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n5239) );
  NAND2_X1 U6424 ( .A1(DATAI_0_), .A2(n5321), .ZN(n6783) );
  NOR2_X2 U6425 ( .A1(n5322), .A2(n5234), .ZN(n6833) );
  AOI22_X1 U6426 ( .A1(n6832), .A2(n5324), .B1(n6833), .B2(n5323), .ZN(n5238)
         );
  INV_X1 U6427 ( .A(DATAI_24_), .ZN(n5235) );
  NOR2_X1 U6428 ( .A1(n6476), .A2(n5235), .ZN(n6836) );
  AOI22_X1 U6429 ( .A1(n6836), .A2(n5411), .B1(n6562), .B2(n6839), .ZN(n5237)
         );
  OAI211_X1 U6430 ( .C1(n5331), .C2(n5239), .A(n5238), .B(n5237), .ZN(U3036)
         );
  INV_X1 U6431 ( .A(n6839), .ZN(n6581) );
  AOI22_X1 U6432 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n5376), .B1(n6832), 
        .B2(n5375), .ZN(n5241) );
  AOI22_X1 U6433 ( .A1(n6668), .A2(n6836), .B1(n6833), .B2(n5377), .ZN(n5240)
         );
  OAI211_X1 U6434 ( .C1(n5416), .C2(n6581), .A(n5241), .B(n5240), .ZN(U3092)
         );
  XNOR2_X1 U6435 ( .A(n5242), .B(n5243), .ZN(n5316) );
  AOI21_X1 U6436 ( .B1(n5250), .B2(n6521), .A(n5462), .ZN(n5253) );
  NOR2_X1 U6437 ( .A1(n4644), .A2(n5244), .ZN(n6513) );
  OR2_X1 U6438 ( .A1(n6180), .A2(n5245), .ZN(n5246) );
  NAND2_X1 U6439 ( .A1(n6161), .A2(n5246), .ZN(n6303) );
  NAND2_X1 U6440 ( .A1(n6523), .A2(REIP_REG_8__SCAN_IN), .ZN(n5312) );
  OAI21_X1 U6441 ( .B1(n6512), .B2(n6303), .A(n5312), .ZN(n5252) );
  INV_X1 U6442 ( .A(n5736), .ZN(n5249) );
  AOI22_X1 U6443 ( .A1(n5249), .A2(n5248), .B1(n5484), .B2(n5247), .ZN(n6522)
         );
  NOR2_X1 U6444 ( .A1(n6522), .A2(n5250), .ZN(n5251) );
  AOI211_X1 U6445 ( .C1(n5253), .C2(n6513), .A(n5252), .B(n5251), .ZN(n5254)
         );
  OAI21_X1 U6446 ( .B1(n6051), .B2(n5316), .A(n5254), .ZN(U3010) );
  INV_X1 U6447 ( .A(n5255), .ZN(n5258) );
  OAI21_X1 U6448 ( .B1(n5258), .B2(n5257), .A(n5256), .ZN(n6475) );
  INV_X1 U6449 ( .A(n5259), .ZN(n5260) );
  NAND3_X1 U6450 ( .A1(n5260), .A2(n4214), .A3(n7002), .ZN(n5891) );
  OR2_X1 U6451 ( .A1(n5891), .A2(n5261), .ZN(n5262) );
  NOR2_X1 U6452 ( .A1(n5262), .A2(n4728), .ZN(n5263) );
  NOR2_X2 U6453 ( .A1(n6335), .A2(n6336), .ZN(n6366) );
  OAI222_X1 U6454 ( .A1(n6475), .A2(n6368), .B1(n5269), .B2(n6366), .C1(n6418), 
        .C2(n6365), .ZN(U2884) );
  OAI21_X1 U6455 ( .B1(n4897), .B2(n5271), .A(n5270), .ZN(n6482) );
  OAI222_X1 U6456 ( .A1(n6482), .A2(n6368), .B1(n5272), .B2(n6366), .C1(n6423), 
        .C2(n6365), .ZN(U2886) );
  NOR2_X1 U6457 ( .A1(n5274), .A2(n5273), .ZN(n5275) );
  OR2_X1 U6458 ( .A1(n4898), .A2(n5275), .ZN(n6483) );
  OAI222_X1 U6459 ( .A1(n6483), .A2(n6368), .B1(n5276), .B2(n6366), .C1(n6428), 
        .C2(n6365), .ZN(U2889) );
  INV_X1 U6460 ( .A(n5416), .ZN(n5277) );
  NAND2_X1 U6461 ( .A1(n4966), .A2(n6719), .ZN(n6568) );
  OAI21_X1 U6462 ( .B1(n5277), .B2(n6711), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n5278) );
  NAND2_X1 U6463 ( .A1(n5278), .A2(n6643), .ZN(n5286) );
  INV_X1 U6464 ( .A(n5286), .ZN(n5284) );
  INV_X1 U6465 ( .A(n5279), .ZN(n5280) );
  NAND2_X1 U6466 ( .A1(n5280), .A2(n6636), .ZN(n6680) );
  NAND2_X1 U6467 ( .A1(n5281), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6685) );
  NOR2_X1 U6468 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6685), .ZN(n5414)
         );
  OAI21_X1 U6469 ( .B1(n7000), .B2(n5414), .A(n6729), .ZN(n5283) );
  AOI211_X2 U6470 ( .C1(n5284), .C2(n6680), .A(n5283), .B(n5282), .ZN(n5421)
         );
  INV_X1 U6471 ( .A(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n5290) );
  OAI22_X1 U6472 ( .A1(n5286), .A2(n6680), .B1(n5285), .B2(n6725), .ZN(n5418)
         );
  AOI22_X1 U6473 ( .A1(n6786), .A2(n6711), .B1(n6784), .B2(n5414), .ZN(n5287)
         );
  OAI21_X1 U6474 ( .B1(n5416), .B2(n6654), .A(n5287), .ZN(n5288) );
  AOI21_X1 U6475 ( .B1(n5418), .B2(n6736), .A(n5288), .ZN(n5289) );
  OAI21_X1 U6476 ( .B1(n5421), .B2(n5290), .A(n5289), .ZN(U3101) );
  INV_X1 U6477 ( .A(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n5294) );
  AOI22_X1 U6478 ( .A1(n6816), .A2(n6711), .B1(n6814), .B2(n5414), .ZN(n5291)
         );
  OAI21_X1 U6479 ( .B1(n5416), .B2(n6709), .A(n5291), .ZN(n5292) );
  AOI21_X1 U6480 ( .B1(n5418), .B2(n6756), .A(n5292), .ZN(n5293) );
  OAI21_X1 U6481 ( .B1(n5421), .B2(n5294), .A(n5293), .ZN(U3106) );
  AOI22_X1 U6482 ( .A1(n6810), .A2(n6711), .B1(n6808), .B2(n5414), .ZN(n5295)
         );
  OAI21_X1 U6483 ( .B1(n5416), .B2(n6705), .A(n5295), .ZN(n5296) );
  AOI21_X1 U6484 ( .B1(n5418), .B2(n6752), .A(n5296), .ZN(n5297) );
  OAI21_X1 U6485 ( .B1(n5421), .B2(n4327), .A(n5297), .ZN(U3105) );
  INV_X1 U6486 ( .A(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n5301) );
  AOI22_X1 U6487 ( .A1(n6791), .A2(n6711), .B1(n6790), .B2(n5414), .ZN(n5298)
         );
  OAI21_X1 U6488 ( .B1(n5416), .B2(n6657), .A(n5298), .ZN(n5299) );
  AOI21_X1 U6489 ( .B1(n5418), .B2(n6740), .A(n5299), .ZN(n5300) );
  OAI21_X1 U6490 ( .B1(n5421), .B2(n5301), .A(n5300), .ZN(U3102) );
  INV_X1 U6491 ( .A(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n5305) );
  AOI22_X1 U6492 ( .A1(n6798), .A2(n6711), .B1(n6796), .B2(n5414), .ZN(n5302)
         );
  OAI21_X1 U6493 ( .B1(n5416), .B2(n6699), .A(n5302), .ZN(n5303) );
  AOI21_X1 U6494 ( .B1(n5418), .B2(n6744), .A(n5303), .ZN(n5304) );
  OAI21_X1 U6495 ( .B1(n5421), .B2(n5305), .A(n5304), .ZN(U3103) );
  INV_X1 U6496 ( .A(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n5309) );
  AOI22_X1 U6497 ( .A1(n6823), .A2(n5442), .B1(n6821), .B2(n6825), .ZN(n5306)
         );
  OAI21_X1 U6498 ( .B1(n6717), .B2(n5444), .A(n5306), .ZN(n5307) );
  AOI21_X1 U6499 ( .B1(n6762), .B2(n5446), .A(n5307), .ZN(n5308) );
  OAI21_X1 U6500 ( .B1(n5449), .B2(n5309), .A(n5308), .ZN(U3139) );
  AOI21_X1 U6501 ( .B1(n5311), .B2(n5256), .A(n5310), .ZN(n6302) );
  NAND2_X1 U6502 ( .A1(n6302), .A2(n5989), .ZN(n5315) );
  OAI21_X1 U6503 ( .B1(n5640), .B2(n6170), .A(n5312), .ZN(n5313) );
  AOI21_X1 U6504 ( .B1(n6498), .B2(n6171), .A(n5313), .ZN(n5314) );
  OAI211_X1 U6505 ( .C1(n6484), .C2(n5316), .A(n5315), .B(n5314), .ZN(U2978)
         );
  INV_X1 U6506 ( .A(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n5320) );
  AOI22_X1 U6507 ( .A1(n6820), .A2(n6711), .B1(n6823), .B2(n5414), .ZN(n5317)
         );
  OAI21_X1 U6508 ( .B1(n5416), .B2(n6673), .A(n5317), .ZN(n5318) );
  AOI21_X1 U6509 ( .B1(n5418), .B2(n6762), .A(n5318), .ZN(n5319) );
  OAI21_X1 U6510 ( .B1(n5421), .B2(n5320), .A(n5319), .ZN(U3107) );
  NAND2_X1 U6511 ( .A1(DATAI_4_), .A2(n5321), .ZN(n6807) );
  NOR2_X2 U6512 ( .A1(n5322), .A2(n3456), .ZN(n6802) );
  AOI22_X1 U6513 ( .A1(n6748), .A2(n5324), .B1(n6802), .B2(n5323), .ZN(n5330)
         );
  NAND2_X1 U6514 ( .A1(n5989), .A2(DATAI_28_), .ZN(n6702) );
  INV_X1 U6515 ( .A(DATAI_20_), .ZN(n5325) );
  NOR2_X1 U6516 ( .A1(n6476), .A2(n5325), .ZN(n6804) );
  INV_X1 U6517 ( .A(n6804), .ZN(n6591) );
  OAI22_X1 U6518 ( .A1(n6702), .A2(n5327), .B1(n5326), .B2(n6591), .ZN(n5328)
         );
  INV_X1 U6519 ( .A(n5328), .ZN(n5329) );
  OAI211_X1 U6520 ( .C1(n5331), .C2(n4345), .A(n5330), .B(n5329), .ZN(U3040)
         );
  INV_X1 U6521 ( .A(n5449), .ZN(n5335) );
  AOI22_X1 U6522 ( .A1(n6833), .A2(n5442), .B1(n6821), .B2(n6836), .ZN(n5333)
         );
  NAND2_X1 U6523 ( .A1(n6832), .A2(n5446), .ZN(n5332) );
  OAI211_X1 U6524 ( .C1(n5444), .C2(n6581), .A(n5333), .B(n5332), .ZN(n5334)
         );
  AOI21_X1 U6525 ( .B1(n5335), .B2(INSTQUEUE_REG_14__0__SCAN_IN), .A(n5334), 
        .ZN(n5336) );
  INV_X1 U6526 ( .A(n5336), .ZN(U3132) );
  AOI21_X1 U6527 ( .B1(n5337), .B2(n6643), .A(n6723), .ZN(n5340) );
  NOR2_X1 U6528 ( .A1(n6769), .A2(n5341), .ZN(n5408) );
  AOI21_X1 U6529 ( .B1(n5338), .B2(n6681), .A(n5408), .ZN(n5343) );
  OAI22_X1 U6530 ( .A1(n5340), .A2(n5343), .B1(n5341), .B2(n6773), .ZN(n5339)
         );
  INV_X1 U6531 ( .A(n6744), .ZN(n6801) );
  INV_X1 U6532 ( .A(n5340), .ZN(n5342) );
  AOI22_X1 U6533 ( .A1(n5343), .A2(n5342), .B1(n5341), .B2(n6776), .ZN(n5344)
         );
  NAND2_X1 U6534 ( .A1(n6780), .A2(n5344), .ZN(n5407) );
  AOI22_X1 U6535 ( .A1(n6796), .A2(n5408), .B1(INSTQUEUE_REG_1__3__SCAN_IN), 
        .B2(n5407), .ZN(n5345) );
  OAI21_X1 U6536 ( .B1(n6699), .B2(n5433), .A(n5345), .ZN(n5346) );
  AOI21_X1 U6537 ( .B1(n6798), .B2(n5411), .A(n5346), .ZN(n5347) );
  OAI21_X1 U6538 ( .B1(n5413), .B2(n6801), .A(n5347), .ZN(U3031) );
  INV_X1 U6539 ( .A(n6762), .ZN(n6829) );
  AOI22_X1 U6540 ( .A1(n6823), .A2(n5408), .B1(INSTQUEUE_REG_1__7__SCAN_IN), 
        .B2(n5407), .ZN(n5348) );
  OAI21_X1 U6541 ( .B1(n6673), .B2(n5433), .A(n5348), .ZN(n5349) );
  AOI21_X1 U6542 ( .B1(n6820), .B2(n5411), .A(n5349), .ZN(n5350) );
  OAI21_X1 U6543 ( .B1(n5413), .B2(n6829), .A(n5350), .ZN(U3035) );
  INV_X1 U6544 ( .A(n6740), .ZN(n6795) );
  AOI22_X1 U6545 ( .A1(n6790), .A2(n5408), .B1(INSTQUEUE_REG_1__2__SCAN_IN), 
        .B2(n5407), .ZN(n5351) );
  OAI21_X1 U6546 ( .B1(n6657), .B2(n5433), .A(n5351), .ZN(n5352) );
  AOI21_X1 U6547 ( .B1(n6791), .B2(n5411), .A(n5352), .ZN(n5353) );
  OAI21_X1 U6548 ( .B1(n5413), .B2(n6795), .A(n5353), .ZN(U3030) );
  INV_X1 U6549 ( .A(n6736), .ZN(n6789) );
  AOI22_X1 U6550 ( .A1(n6784), .A2(n5408), .B1(INSTQUEUE_REG_1__1__SCAN_IN), 
        .B2(n5407), .ZN(n5354) );
  OAI21_X1 U6551 ( .B1(n6654), .B2(n5433), .A(n5354), .ZN(n5355) );
  AOI21_X1 U6552 ( .B1(n6786), .B2(n5411), .A(n5355), .ZN(n5356) );
  OAI21_X1 U6553 ( .B1(n5413), .B2(n6789), .A(n5356), .ZN(U3029) );
  INV_X1 U6554 ( .A(n6752), .ZN(n6813) );
  AOI22_X1 U6555 ( .A1(n6808), .A2(n5408), .B1(INSTQUEUE_REG_1__5__SCAN_IN), 
        .B2(n5407), .ZN(n5357) );
  OAI21_X1 U6556 ( .B1(n6705), .B2(n5433), .A(n5357), .ZN(n5358) );
  AOI21_X1 U6557 ( .B1(n6810), .B2(n5411), .A(n5358), .ZN(n5359) );
  OAI21_X1 U6558 ( .B1(n5413), .B2(n6813), .A(n5359), .ZN(U3033) );
  INV_X1 U6559 ( .A(n6823), .ZN(n5367) );
  OAI22_X1 U6560 ( .A1(n5367), .A2(n5434), .B1(n6717), .B2(n5452), .ZN(n5360)
         );
  AOI21_X1 U6561 ( .B1(n6762), .B2(n5437), .A(n5360), .ZN(n5362) );
  NAND2_X1 U6562 ( .A1(n5438), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n5361) );
  OAI211_X1 U6563 ( .C1(n5441), .C2(n6673), .A(n5362), .B(n5361), .ZN(U3059)
         );
  INV_X1 U6564 ( .A(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n5366) );
  NOR2_X1 U6565 ( .A1(n5444), .A2(n6673), .ZN(n5364) );
  OAI22_X1 U6566 ( .A1(n5367), .A2(n5422), .B1(n6717), .B2(n6835), .ZN(n5363)
         );
  AOI211_X1 U6567 ( .C1(n6762), .C2(n6831), .A(n5364), .B(n5363), .ZN(n5365)
         );
  OAI21_X1 U6568 ( .B1(n6843), .B2(n5366), .A(n5365), .ZN(U3147) );
  NAND2_X1 U6569 ( .A1(n5427), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n5370) );
  OAI22_X1 U6570 ( .A1(n5367), .A2(n5428), .B1(n6673), .B2(n6835), .ZN(n5368)
         );
  AOI21_X1 U6571 ( .B1(n6762), .B2(n5430), .A(n5368), .ZN(n5369) );
  OAI211_X1 U6572 ( .C1(n5433), .C2(n6717), .A(n5370), .B(n5369), .ZN(U3027)
         );
  INV_X1 U6573 ( .A(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n5374) );
  AOI22_X1 U6574 ( .A1(n6600), .A2(n6820), .B1(n6823), .B2(n5450), .ZN(n5371)
         );
  OAI21_X1 U6575 ( .B1(n6673), .B2(n5452), .A(n5371), .ZN(n5372) );
  AOI21_X1 U6576 ( .B1(n5454), .B2(n6762), .A(n5372), .ZN(n5373) );
  OAI21_X1 U6577 ( .B1(n5457), .B2(n5374), .A(n5373), .ZN(U3067) );
  AOI22_X1 U6578 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n5376), .B1(n6748), 
        .B2(n5375), .ZN(n5379) );
  INV_X1 U6579 ( .A(n6702), .ZN(n6803) );
  AOI22_X1 U6580 ( .A1(n6668), .A2(n6803), .B1(n5377), .B2(n6802), .ZN(n5378)
         );
  OAI211_X1 U6581 ( .C1(n5416), .C2(n6591), .A(n5379), .B(n5378), .ZN(U3096)
         );
  INV_X1 U6582 ( .A(n6836), .ZN(n6690) );
  AOI22_X1 U6583 ( .A1(n6833), .A2(n5408), .B1(INSTQUEUE_REG_1__0__SCAN_IN), 
        .B2(n5407), .ZN(n5380) );
  OAI21_X1 U6584 ( .B1(n6690), .B2(n5433), .A(n5380), .ZN(n5381) );
  AOI21_X1 U6585 ( .B1(n6839), .B2(n5411), .A(n5381), .ZN(n5382) );
  OAI21_X1 U6586 ( .B1(n5413), .B2(n6783), .A(n5382), .ZN(U3028) );
  AOI22_X1 U6587 ( .A1(n6814), .A2(n5408), .B1(INSTQUEUE_REG_1__6__SCAN_IN), 
        .B2(n5407), .ZN(n5383) );
  OAI21_X1 U6588 ( .B1(n6709), .B2(n5433), .A(n5383), .ZN(n5384) );
  AOI21_X1 U6589 ( .B1(n6816), .B2(n5411), .A(n5384), .ZN(n5385) );
  OAI21_X1 U6590 ( .B1(n5413), .B2(n6819), .A(n5385), .ZN(U3034) );
  NAND2_X1 U6591 ( .A1(n5427), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n5388) );
  INV_X1 U6592 ( .A(n6833), .ZN(n5389) );
  OAI22_X1 U6593 ( .A1(n5389), .A2(n5428), .B1(n6690), .B2(n6835), .ZN(n5386)
         );
  AOI21_X1 U6594 ( .B1(n6832), .B2(n5430), .A(n5386), .ZN(n5387) );
  OAI211_X1 U6595 ( .C1(n5433), .C2(n6581), .A(n5388), .B(n5387), .ZN(U3020)
         );
  OAI22_X1 U6596 ( .A1(n5389), .A2(n5434), .B1(n6581), .B2(n5452), .ZN(n5390)
         );
  AOI21_X1 U6597 ( .B1(n6832), .B2(n5437), .A(n5390), .ZN(n5392) );
  NAND2_X1 U6598 ( .A1(n5438), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n5391) );
  OAI211_X1 U6599 ( .C1(n5441), .C2(n6690), .A(n5392), .B(n5391), .ZN(U3052)
         );
  INV_X1 U6600 ( .A(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n5396) );
  AOI22_X1 U6601 ( .A1(n6839), .A2(n6711), .B1(n6833), .B2(n5414), .ZN(n5393)
         );
  OAI21_X1 U6602 ( .B1(n5416), .B2(n6690), .A(n5393), .ZN(n5394) );
  AOI21_X1 U6603 ( .B1(n5418), .B2(n6832), .A(n5394), .ZN(n5395) );
  OAI21_X1 U6604 ( .B1(n5421), .B2(n5396), .A(n5395), .ZN(U3100) );
  XNOR2_X1 U6605 ( .A(n5397), .B(n5398), .ZN(n6505) );
  XOR2_X1 U6606 ( .A(n5310), .B(n5399), .Z(n6352) );
  NAND2_X1 U6607 ( .A1(n6352), .A2(n5989), .ZN(n5402) );
  NAND2_X1 U6608 ( .A1(n6216), .A2(REIP_REG_9__SCAN_IN), .ZN(n6502) );
  OAI21_X1 U6609 ( .B1(n5640), .B2(n6164), .A(n6502), .ZN(n5400) );
  AOI21_X1 U6610 ( .B1(n6498), .B2(n6167), .A(n5400), .ZN(n5401) );
  OAI211_X1 U6611 ( .C1(n6505), .C2(n6484), .A(n5402), .B(n5401), .ZN(U2977)
         );
  INV_X1 U6612 ( .A(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n5406) );
  AOI22_X1 U6613 ( .A1(n6600), .A2(n6839), .B1(n6833), .B2(n5450), .ZN(n5403)
         );
  OAI21_X1 U6614 ( .B1(n6690), .B2(n5452), .A(n5403), .ZN(n5404) );
  AOI21_X1 U6615 ( .B1(n5454), .B2(n6832), .A(n5404), .ZN(n5405) );
  OAI21_X1 U6616 ( .B1(n5457), .B2(n5406), .A(n5405), .ZN(U3060) );
  AOI22_X1 U6617 ( .A1(n6802), .A2(n5408), .B1(INSTQUEUE_REG_1__4__SCAN_IN), 
        .B2(n5407), .ZN(n5409) );
  OAI21_X1 U6618 ( .B1(n6702), .B2(n5433), .A(n5409), .ZN(n5410) );
  AOI21_X1 U6619 ( .B1(n6804), .B2(n5411), .A(n5410), .ZN(n5412) );
  OAI21_X1 U6620 ( .B1(n5413), .B2(n6807), .A(n5412), .ZN(U3032) );
  INV_X1 U6621 ( .A(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n5420) );
  AOI22_X1 U6622 ( .A1(n6804), .A2(n6711), .B1(n6802), .B2(n5414), .ZN(n5415)
         );
  OAI21_X1 U6623 ( .B1(n5416), .B2(n6702), .A(n5415), .ZN(n5417) );
  AOI21_X1 U6624 ( .B1(n5418), .B2(n6748), .A(n5417), .ZN(n5419) );
  OAI21_X1 U6625 ( .B1(n5421), .B2(n5420), .A(n5419), .ZN(U3104) );
  INV_X1 U6626 ( .A(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n5426) );
  NOR2_X1 U6627 ( .A1(n5444), .A2(n6702), .ZN(n5424) );
  INV_X1 U6628 ( .A(n6802), .ZN(n5435) );
  OAI22_X1 U6629 ( .A1(n5435), .A2(n5422), .B1(n6591), .B2(n6835), .ZN(n5423)
         );
  AOI211_X1 U6630 ( .C1(n6748), .C2(n6831), .A(n5424), .B(n5423), .ZN(n5425)
         );
  OAI21_X1 U6631 ( .B1(n6843), .B2(n5426), .A(n5425), .ZN(U3144) );
  NAND2_X1 U6632 ( .A1(n5427), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n5432) );
  OAI22_X1 U6633 ( .A1(n5435), .A2(n5428), .B1(n6702), .B2(n6835), .ZN(n5429)
         );
  AOI21_X1 U6634 ( .B1(n6748), .B2(n5430), .A(n5429), .ZN(n5431) );
  OAI211_X1 U6635 ( .C1(n5433), .C2(n6591), .A(n5432), .B(n5431), .ZN(U3024)
         );
  OAI22_X1 U6636 ( .A1(n5435), .A2(n5434), .B1(n5452), .B2(n6591), .ZN(n5436)
         );
  AOI21_X1 U6637 ( .B1(n6748), .B2(n5437), .A(n5436), .ZN(n5440) );
  NAND2_X1 U6638 ( .A1(n5438), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n5439) );
  OAI211_X1 U6639 ( .C1(n5441), .C2(n6702), .A(n5440), .B(n5439), .ZN(U3056)
         );
  INV_X1 U6640 ( .A(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n5448) );
  AOI22_X1 U6641 ( .A1(n6803), .A2(n6821), .B1(n6802), .B2(n5442), .ZN(n5443)
         );
  OAI21_X1 U6642 ( .B1(n6591), .B2(n5444), .A(n5443), .ZN(n5445) );
  AOI21_X1 U6643 ( .B1(n6748), .B2(n5446), .A(n5445), .ZN(n5447) );
  OAI21_X1 U6644 ( .B1(n5449), .B2(n5448), .A(n5447), .ZN(U3136) );
  INV_X1 U6645 ( .A(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n5456) );
  AOI22_X1 U6646 ( .A1(n6600), .A2(n6804), .B1(n6802), .B2(n5450), .ZN(n5451)
         );
  OAI21_X1 U6647 ( .B1(n6702), .B2(n5452), .A(n5451), .ZN(n5453) );
  AOI21_X1 U6648 ( .B1(n5454), .B2(n6748), .A(n5453), .ZN(n5455) );
  OAI21_X1 U6649 ( .B1(n5457), .B2(n5456), .A(n5455), .ZN(U3064) );
  XNOR2_X1 U6650 ( .A(n5458), .B(n5459), .ZN(n5475) );
  OAI21_X1 U6651 ( .B1(n5646), .B2(n5462), .A(n6522), .ZN(n6506) );
  AND2_X1 U6652 ( .A1(n6159), .A2(n5460), .ZN(n5461) );
  OR2_X1 U6653 ( .A1(n5461), .A2(n5486), .ZN(n6298) );
  INV_X1 U6654 ( .A(REIP_REG_10__SCAN_IN), .ZN(n6943) );
  OAI22_X1 U6655 ( .A1(n6512), .A2(n6298), .B1(n6943), .B2(n3179), .ZN(n5466)
         );
  NAND2_X1 U6656 ( .A1(n5462), .A2(n6513), .ZN(n6510) );
  AOI221_X1 U6657 ( .B1(INSTADDRPOINTER_REG_10__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_9__SCAN_IN), .C1(n5464), .C2(n5463), .A(n6510), 
        .ZN(n5465) );
  AOI211_X1 U6658 ( .C1(INSTADDRPOINTER_REG_10__SCAN_IN), .C2(n6506), .A(n5466), .B(n5465), .ZN(n5467) );
  OAI21_X1 U6659 ( .B1(n5475), .B2(n6051), .A(n5467), .ZN(U3008) );
  AOI21_X1 U6660 ( .B1(n5470), .B2(n5469), .A(n5468), .ZN(n6149) );
  NAND2_X1 U6661 ( .A1(n6149), .A2(n5989), .ZN(n5474) );
  INV_X1 U6662 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n5471) );
  OAI22_X1 U6663 ( .A1(n5640), .A2(n5471), .B1(n3179), .B2(n6943), .ZN(n5472)
         );
  AOI21_X1 U6664 ( .B1(n6498), .B2(n6151), .A(n5472), .ZN(n5473) );
  OAI211_X1 U6665 ( .C1(n5475), .C2(n6484), .A(n5474), .B(n5473), .ZN(U2976)
         );
  XNOR2_X1 U6666 ( .A(n5476), .B(n5477), .ZN(n5492) );
  XOR2_X1 U6667 ( .A(n5468), .B(n5478), .Z(n6140) );
  NAND2_X1 U6668 ( .A1(n6140), .A2(n5989), .ZN(n5481) );
  NAND2_X1 U6669 ( .A1(n6216), .A2(REIP_REG_11__SCAN_IN), .ZN(n5488) );
  OAI21_X1 U6670 ( .B1(n5640), .B2(n6144), .A(n5488), .ZN(n5479) );
  AOI21_X1 U6671 ( .B1(n6498), .B2(n6147), .A(n5479), .ZN(n5480) );
  OAI211_X1 U6672 ( .C1(n5492), .C2(n6484), .A(n5481), .B(n5480), .ZN(U2975)
         );
  AOI21_X1 U6673 ( .B1(n5484), .B2(n5483), .A(n5482), .ZN(n5521) );
  INV_X1 U6674 ( .A(n5521), .ZN(n6043) );
  AOI22_X1 U6675 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n6043), .B1(n6045), .B2(n5496), .ZN(n5491) );
  NOR2_X1 U6676 ( .A1(n5486), .A2(n5485), .ZN(n5487) );
  INV_X1 U6677 ( .A(n5488), .ZN(n5489) );
  AOI21_X1 U6678 ( .B1(n6525), .B2(n3222), .A(n5489), .ZN(n5490) );
  OAI211_X1 U6679 ( .C1(n5492), .C2(n6051), .A(n5491), .B(n5490), .ZN(U3007)
         );
  XNOR2_X1 U6680 ( .A(n5493), .B(n5494), .ZN(n5511) );
  XNOR2_X1 U6681 ( .A(n5526), .B(n5524), .ZN(n6294) );
  NOR2_X1 U6682 ( .A1(n3179), .A2(n6948), .ZN(n5502) );
  NOR2_X1 U6683 ( .A1(n5495), .A2(n5496), .ZN(n5500) );
  AOI221_X1 U6684 ( .B1(n5497), .B2(n5496), .C1(n6036), .C2(n5496), .A(n6043), 
        .ZN(n5498) );
  INV_X1 U6685 ( .A(n5498), .ZN(n5499) );
  MUX2_X1 U6686 ( .A(n5500), .B(n5499), .S(INSTADDRPOINTER_REG_12__SCAN_IN), 
        .Z(n5501) );
  AOI211_X1 U6687 ( .C1(n6525), .C2(n6294), .A(n5502), .B(n5501), .ZN(n5503)
         );
  OAI21_X1 U6688 ( .B1(n5511), .B2(n6051), .A(n5503), .ZN(U3006) );
  AOI21_X1 U6689 ( .B1(n5506), .B2(n5505), .A(n5504), .ZN(n6345) );
  NAND2_X1 U6690 ( .A1(n6345), .A2(n5989), .ZN(n5510) );
  INV_X1 U6691 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n5507) );
  OAI22_X1 U6692 ( .A1(n5640), .A2(n5507), .B1(n3179), .B2(n6948), .ZN(n5508)
         );
  AOI21_X1 U6693 ( .B1(n6498), .B2(n6134), .A(n5508), .ZN(n5509) );
  OAI211_X1 U6694 ( .C1(n5511), .C2(n6484), .A(n5510), .B(n5509), .ZN(U2974)
         );
  INV_X1 U6695 ( .A(n5513), .ZN(n5514) );
  AOI21_X1 U6696 ( .B1(n5515), .B2(n3185), .A(n5514), .ZN(n5538) );
  INV_X1 U6697 ( .A(n5516), .ZN(n5519) );
  AOI22_X1 U6698 ( .A1(n5519), .A2(n5518), .B1(n5517), .B2(n5522), .ZN(n5520)
         );
  NAND2_X1 U6699 ( .A1(n5521), .A2(n5520), .ZN(n5560) );
  NOR2_X1 U6700 ( .A1(INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n5522), .ZN(n5523)
         );
  AOI22_X1 U6701 ( .A1(INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n5560), .B1(n5523), .B2(n6045), .ZN(n5532) );
  INV_X1 U6702 ( .A(n5524), .ZN(n5525) );
  NAND2_X1 U6703 ( .A1(n5526), .A2(n5525), .ZN(n5528) );
  INV_X1 U6704 ( .A(n5550), .ZN(n5527) );
  AOI21_X1 U6705 ( .B1(n5529), .B2(n5528), .A(n5527), .ZN(n6291) );
  NAND2_X1 U6706 ( .A1(n6216), .A2(REIP_REG_13__SCAN_IN), .ZN(n5534) );
  INV_X1 U6707 ( .A(n5534), .ZN(n5530) );
  AOI21_X1 U6708 ( .B1(n6291), .B2(n6525), .A(n5530), .ZN(n5531) );
  OAI211_X1 U6709 ( .C1(n5538), .C2(n6051), .A(n5532), .B(n5531), .ZN(U3005)
         );
  XOR2_X1 U6710 ( .A(n5504), .B(n5533), .Z(n6292) );
  NAND2_X1 U6711 ( .A1(n6292), .A2(n5989), .ZN(n5537) );
  OAI21_X1 U6712 ( .B1(n5640), .B2(n6128), .A(n5534), .ZN(n5535) );
  AOI21_X1 U6713 ( .B1(n6498), .B2(n6132), .A(n5535), .ZN(n5536) );
  OAI211_X1 U6714 ( .C1(n5538), .C2(n6484), .A(n5537), .B(n5536), .ZN(U2973)
         );
  INV_X1 U6715 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5554) );
  NAND2_X1 U6716 ( .A1(n5633), .A2(n5554), .ZN(n5758) );
  NAND2_X1 U6717 ( .A1(n3704), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5541) );
  NAND2_X1 U6718 ( .A1(n5758), .A2(n5541), .ZN(n5540) );
  MUX2_X1 U6719 ( .A(n5758), .B(n5540), .S(n5539), .Z(n5542) );
  OR2_X1 U6720 ( .A1(n5539), .A2(n5541), .ZN(n5757) );
  NAND2_X1 U6721 ( .A1(n5542), .A2(n5757), .ZN(n5563) );
  AOI21_X1 U6722 ( .B1(n5545), .B2(n5544), .A(n5543), .ZN(n6288) );
  NAND2_X1 U6723 ( .A1(n6498), .A2(n6120), .ZN(n5546) );
  NAND2_X1 U6724 ( .A1(n6216), .A2(REIP_REG_14__SCAN_IN), .ZN(n5552) );
  OAI211_X1 U6725 ( .C1(n5640), .C2(n6118), .A(n5546), .B(n5552), .ZN(n5547)
         );
  AOI21_X1 U6726 ( .B1(n6288), .B2(n5989), .A(n5547), .ZN(n5548) );
  OAI21_X1 U6727 ( .B1(n6484), .B2(n5563), .A(n5548), .ZN(U2972) );
  NAND2_X1 U6728 ( .A1(n6046), .A2(n6045), .ZN(n6047) );
  INV_X1 U6729 ( .A(n6047), .ZN(n5555) );
  NAND2_X1 U6730 ( .A1(n5550), .A2(n5549), .ZN(n5551) );
  NAND2_X1 U6731 ( .A1(n6060), .A2(n5551), .ZN(n6289) );
  OAI21_X1 U6732 ( .B1(n6289), .B2(n6512), .A(n5552), .ZN(n5553) );
  AOI21_X1 U6733 ( .B1(n5555), .B2(n5554), .A(n5553), .ZN(n5562) );
  INV_X1 U6734 ( .A(n5556), .ZN(n5558) );
  AOI21_X1 U6735 ( .B1(n5558), .B2(n5557), .A(INSTADDRPOINTER_REG_13__SCAN_IN), 
        .ZN(n5559) );
  OAI21_X1 U6736 ( .B1(n5560), .B2(n5559), .A(INSTADDRPOINTER_REG_14__SCAN_IN), 
        .ZN(n5561) );
  OAI211_X1 U6737 ( .C1(n5563), .C2(n6051), .A(n5562), .B(n5561), .ZN(U3004)
         );
  NAND2_X1 U6738 ( .A1(n6050), .A2(n5565), .ZN(n5566) );
  NAND2_X1 U6739 ( .A1(n6034), .A2(n5566), .ZN(n6280) );
  OAI21_X1 U6740 ( .B1(n5569), .B2(n5567), .A(n5568), .ZN(n6282) );
  INV_X1 U6741 ( .A(n6282), .ZN(n6331) );
  INV_X1 U6742 ( .A(EBX_REG_31__SCAN_IN), .ZN(n5570) );
  NAND2_X1 U6743 ( .A1(n5571), .A2(n5570), .ZN(n5574) );
  INV_X1 U6744 ( .A(n5572), .ZN(n5573) );
  INV_X1 U6745 ( .A(n6903), .ZN(n5575) );
  AOI22_X1 U6746 ( .A1(PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n6234), .B1(n5992), 
        .B2(n6261), .ZN(n5577) );
  OAI211_X1 U6747 ( .C1(n6245), .C2(n6281), .A(n5577), .B(n3179), .ZN(n5578)
         );
  AOI21_X1 U6748 ( .B1(n6201), .B2(n6331), .A(n5578), .ZN(n5584) );
  INV_X1 U6749 ( .A(REIP_REG_16__SCAN_IN), .ZN(n6955) );
  INV_X1 U6750 ( .A(REIP_REG_15__SCAN_IN), .ZN(n6953) );
  NOR3_X1 U6751 ( .A1(n5862), .A2(n6955), .A3(n6953), .ZN(n5884) );
  INV_X1 U6752 ( .A(n5579), .ZN(n5580) );
  NOR2_X1 U6753 ( .A1(n6240), .A2(n5580), .ZN(n5581) );
  NOR2_X1 U6754 ( .A1(n6121), .A2(n5581), .ZN(n6099) );
  INV_X1 U6755 ( .A(n6099), .ZN(n5582) );
  OAI21_X1 U6756 ( .B1(n5884), .B2(REIP_REG_17__SCAN_IN), .A(n5582), .ZN(n5583) );
  OAI211_X1 U6757 ( .C1(n6236), .C2(n6280), .A(n5584), .B(n5583), .ZN(U2810)
         );
  NAND2_X1 U6758 ( .A1(n5585), .A2(n5586), .ZN(n5587) );
  XNOR2_X1 U6759 ( .A(n5587), .B(n3211), .ZN(n6052) );
  AOI21_X1 U6760 ( .B1(n5589), .B2(n5588), .A(n5567), .ZN(n6334) );
  INV_X1 U6761 ( .A(n6108), .ZN(n5591) );
  AOI22_X1 U6762 ( .A1(n6491), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .B1(n6523), 
        .B2(REIP_REG_16__SCAN_IN), .ZN(n5590) );
  OAI21_X1 U6763 ( .B1(n6490), .B2(n5591), .A(n5590), .ZN(n5592) );
  AOI21_X1 U6764 ( .B1(n6334), .B2(n5989), .A(n5592), .ZN(n5593) );
  OAI21_X1 U6765 ( .B1(n6484), .B2(n6052), .A(n5593), .ZN(U2970) );
  AOI21_X1 U6766 ( .B1(n5597), .B2(n5594), .A(n5601), .ZN(n5604) );
  NOR3_X1 U6767 ( .A1(n7002), .A2(n5596), .A3(n5595), .ZN(n5599) );
  NOR3_X1 U6768 ( .A1(n5597), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n5753), 
        .ZN(n5598) );
  AOI211_X1 U6769 ( .C1(n6846), .C2(n5600), .A(n5599), .B(n5598), .ZN(n5602)
         );
  OAI22_X1 U6770 ( .A1(n5604), .A2(n5603), .B1(n5602), .B2(n5601), .ZN(U3459)
         );
  NAND2_X1 U6771 ( .A1(n5607), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5610) );
  NAND2_X1 U6772 ( .A1(n5608), .A2(n5673), .ZN(n5609) );
  NAND2_X1 U6773 ( .A1(n5771), .A2(n6498), .ZN(n5612) );
  NAND2_X1 U6774 ( .A1(n6216), .A2(REIP_REG_30__SCAN_IN), .ZN(n5660) );
  OAI211_X1 U6775 ( .C1(n5640), .C2(n5769), .A(n5612), .B(n5660), .ZN(n5613)
         );
  AOI21_X1 U6776 ( .B1(n5654), .B2(n6496), .A(n5613), .ZN(n5614) );
  OAI21_X1 U6777 ( .B1(n5927), .B2(n6476), .A(n5614), .ZN(U2956) );
  AOI21_X1 U6778 ( .B1(n5616), .B2(n5615), .A(n4227), .ZN(n5699) );
  XOR2_X1 U6779 ( .A(n5617), .B(n3219), .Z(n5938) );
  NAND2_X1 U6780 ( .A1(n5938), .A2(n5989), .ZN(n5620) );
  NAND2_X1 U6781 ( .A1(n6523), .A2(REIP_REG_25__SCAN_IN), .ZN(n5694) );
  OAI21_X1 U6782 ( .B1(n5640), .B2(n4389), .A(n5694), .ZN(n5618) );
  AOI21_X1 U6783 ( .B1(n5819), .B2(n6498), .A(n5618), .ZN(n5619) );
  OAI211_X1 U6784 ( .C1(n5699), .C2(n6484), .A(n5620), .B(n5619), .ZN(U2961)
         );
  INV_X1 U6785 ( .A(n5621), .ZN(n5720) );
  NAND2_X1 U6786 ( .A1(n5720), .A2(n5622), .ZN(n5636) );
  NAND3_X1 U6787 ( .A1(n3704), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5623) );
  OAI22_X1 U6788 ( .A1(n5636), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .B1(n5624), .B2(n5623), .ZN(n5625) );
  XNOR2_X1 U6789 ( .A(n5625), .B(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5708)
         );
  INV_X1 U6790 ( .A(n5627), .ZN(n5628) );
  XNOR2_X1 U6791 ( .A(n5626), .B(n5628), .ZN(n5941) );
  NAND2_X1 U6792 ( .A1(n6498), .A2(n5826), .ZN(n5629) );
  NAND2_X1 U6793 ( .A1(n6216), .A2(REIP_REG_24__SCAN_IN), .ZN(n5704) );
  OAI211_X1 U6794 ( .C1(n5640), .C2(n5630), .A(n5629), .B(n5704), .ZN(n5631)
         );
  AOI21_X1 U6795 ( .B1(n5941), .B2(n5989), .A(n5631), .ZN(n5632) );
  OAI21_X1 U6796 ( .B1(n5708), .B2(n6484), .A(n5632), .ZN(U2962) );
  NOR2_X1 U6797 ( .A1(n5585), .A2(n5633), .ZN(n5739) );
  NAND2_X1 U6798 ( .A1(n5739), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5985) );
  INV_X1 U6799 ( .A(n6023), .ZN(n5635) );
  NAND3_X1 U6800 ( .A1(n5635), .A2(n5634), .A3(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5637) );
  OAI21_X1 U6801 ( .B1(n5985), .B2(n5637), .A(n5636), .ZN(n5638) );
  XNOR2_X1 U6802 ( .A(n5638), .B(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5719)
         );
  NAND2_X1 U6803 ( .A1(n6523), .A2(REIP_REG_23__SCAN_IN), .ZN(n5712) );
  OAI21_X1 U6804 ( .B1(n5640), .B2(n5639), .A(n5712), .ZN(n5643) );
  OAI21_X1 U6805 ( .B1(n4072), .B2(n5641), .A(n5626), .ZN(n5946) );
  NOR2_X1 U6806 ( .A1(n5946), .A2(n6476), .ZN(n5642) );
  AOI211_X1 U6807 ( .C1(n5833), .C2(n6498), .A(n5643), .B(n5642), .ZN(n5644)
         );
  OAI21_X1 U6808 ( .B1(n5719), .B2(n6484), .A(n5644), .ZN(U2963) );
  INV_X1 U6809 ( .A(n5645), .ZN(n5653) );
  OAI21_X1 U6810 ( .B1(n5674), .B2(n5646), .A(n5687), .ZN(n5678) );
  AOI21_X1 U6811 ( .B1(n5673), .B2(n6530), .A(n5678), .ZN(n5666) );
  OAI21_X1 U6812 ( .B1(INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n5646), .A(n5666), 
        .ZN(n5651) );
  INV_X1 U6813 ( .A(n5689), .ZN(n5672) );
  AND2_X1 U6814 ( .A1(INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n5672), .ZN(n5647)
         );
  NAND2_X1 U6815 ( .A1(n5674), .A2(n5647), .ZN(n5661) );
  OR3_X1 U6816 ( .A1(n5661), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .A3(n5665), 
        .ZN(n5649) );
  OAI211_X1 U6817 ( .C1(n6274), .C2(n6512), .A(n5649), .B(n5648), .ZN(n5650)
         );
  AOI21_X1 U6818 ( .B1(INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n5651), .A(n5650), 
        .ZN(n5652) );
  OAI21_X1 U6819 ( .B1(n5653), .B2(n6051), .A(n5652), .ZN(U2987) );
  NAND2_X1 U6820 ( .A1(n5654), .A2(n6528), .ZN(n5664) );
  INV_X1 U6821 ( .A(n5655), .ZN(n5657) );
  OAI21_X1 U6822 ( .B1(n5657), .B2(n5669), .A(n5656), .ZN(n5659) );
  XNOR2_X1 U6823 ( .A(n5659), .B(n5658), .ZN(n5897) );
  OAI21_X1 U6824 ( .B1(INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n5661), .A(n5660), 
        .ZN(n5662) );
  AOI21_X1 U6825 ( .B1(n5897), .B2(n6525), .A(n5662), .ZN(n5663) );
  OAI211_X1 U6826 ( .C1(n5666), .C2(n5665), .A(n5664), .B(n5663), .ZN(U2988)
         );
  INV_X1 U6827 ( .A(n5667), .ZN(n5680) );
  NAND2_X1 U6828 ( .A1(n5669), .A2(n5668), .ZN(n5670) );
  NAND3_X1 U6829 ( .A1(n5674), .A2(n5673), .A3(n5672), .ZN(n5675) );
  OAI211_X1 U6830 ( .C1(n5781), .C2(n6512), .A(n5676), .B(n5675), .ZN(n5677)
         );
  AOI21_X1 U6831 ( .B1(INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n5678), .A(n5677), 
        .ZN(n5679) );
  OAI21_X1 U6832 ( .B1(n5680), .B2(n6051), .A(n5679), .ZN(U2989) );
  NAND2_X1 U6833 ( .A1(n4581), .A2(n5681), .ZN(n5682) );
  XNOR2_X1 U6834 ( .A(n5682), .B(n5688), .ZN(n5957) );
  INV_X1 U6835 ( .A(n5957), .ZN(n5693) );
  NOR2_X1 U6836 ( .A1(n5813), .A2(n5683), .ZN(n5684) );
  OR2_X1 U6837 ( .A1(n5685), .A2(n5684), .ZN(n5906) );
  INV_X1 U6838 ( .A(n5906), .ZN(n5691) );
  NAND2_X1 U6839 ( .A1(n6523), .A2(REIP_REG_27__SCAN_IN), .ZN(n5686) );
  OAI221_X1 U6840 ( .B1(INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n5689), .C1(
        n5688), .C2(n5687), .A(n5686), .ZN(n5690) );
  AOI21_X1 U6841 ( .B1(n5691), .B2(n6525), .A(n5690), .ZN(n5692) );
  OAI21_X1 U6842 ( .B1(n5693), .B2(n6051), .A(n5692), .ZN(U2991) );
  INV_X1 U6843 ( .A(n6000), .ZN(n5696) );
  XNOR2_X1 U6844 ( .A(n5809), .B(n5811), .ZN(n5909) );
  NAND2_X1 U6845 ( .A1(n5909), .A2(n6525), .ZN(n5695) );
  OAI211_X1 U6846 ( .C1(INSTADDRPOINTER_REG_25__SCAN_IN), .C2(n5696), .A(n5695), .B(n5694), .ZN(n5697) );
  AOI21_X1 U6847 ( .B1(INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n5996), .A(n5697), 
        .ZN(n5698) );
  OAI21_X1 U6848 ( .B1(n5699), .B2(n6051), .A(n5698), .ZN(U2993) );
  OAI21_X1 U6849 ( .B1(n5709), .B2(n5716), .A(n5700), .ZN(n5706) );
  INV_X1 U6850 ( .A(n5710), .ZN(n5703) );
  INV_X1 U6851 ( .A(n5701), .ZN(n5702) );
  OAI21_X1 U6852 ( .B1(n5703), .B2(n5702), .A(n5809), .ZN(n5912) );
  OAI21_X1 U6853 ( .B1(n5912), .B2(n6512), .A(n5704), .ZN(n5705) );
  AOI21_X1 U6854 ( .B1(n5996), .B2(n5706), .A(n5705), .ZN(n5707) );
  OAI21_X1 U6855 ( .B1(n5708), .B2(n6051), .A(n5707), .ZN(U2994) );
  INV_X1 U6856 ( .A(n5709), .ZN(n5717) );
  OAI21_X1 U6857 ( .B1(n5844), .B2(n5711), .A(n5710), .ZN(n5916) );
  OAI21_X1 U6858 ( .B1(n5916), .B2(n6512), .A(n5712), .ZN(n5715) );
  NOR2_X1 U6859 ( .A1(n5713), .A2(n5716), .ZN(n5714) );
  AOI211_X1 U6860 ( .C1(n5717), .C2(n5716), .A(n5715), .B(n5714), .ZN(n5718)
         );
  OAI21_X1 U6861 ( .B1(n5719), .B2(n6051), .A(n5718), .ZN(U2995) );
  NAND2_X1 U6862 ( .A1(n5722), .A2(n5721), .ZN(n5723) );
  NAND2_X1 U6863 ( .A1(n5621), .A2(n5723), .ZN(n5968) );
  INV_X1 U6864 ( .A(n5968), .ZN(n5733) );
  INV_X1 U6865 ( .A(n5724), .ZN(n5725) );
  OAI21_X1 U6866 ( .B1(n5727), .B2(n5726), .A(n5725), .ZN(n5921) );
  INV_X1 U6867 ( .A(REIP_REG_21__SCAN_IN), .ZN(n5728) );
  OAI22_X1 U6868 ( .A1(n5921), .A2(n6512), .B1(n3179), .B2(n5728), .ZN(n5729)
         );
  AOI21_X1 U6869 ( .B1(n6011), .B2(n5730), .A(n5729), .ZN(n5732) );
  NAND2_X1 U6870 ( .A1(n6006), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5731) );
  OAI211_X1 U6871 ( .C1(n5733), .C2(n6051), .A(n5732), .B(n5731), .ZN(U2997)
         );
  NOR2_X1 U6872 ( .A1(n3703), .A2(n5734), .ZN(n6038) );
  OAI21_X1 U6873 ( .B1(n5736), .B2(n6038), .A(n5735), .ZN(n6037) );
  INV_X1 U6874 ( .A(n6037), .ZN(n5745) );
  NOR2_X1 U6875 ( .A1(n6020), .A2(n6047), .ZN(n5743) );
  NAND3_X1 U6876 ( .A1(n5737), .A2(n5633), .A3(n6058), .ZN(n5986) );
  INV_X1 U6877 ( .A(n5986), .ZN(n5738) );
  NOR2_X1 U6878 ( .A1(n5739), .A2(n5738), .ZN(n5740) );
  XNOR2_X1 U6879 ( .A(n5740), .B(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5993)
         );
  AOI22_X1 U6880 ( .A1(n6528), .A2(n5993), .B1(n6523), .B2(
        REIP_REG_17__SCAN_IN), .ZN(n5741) );
  OAI21_X1 U6881 ( .B1(n6280), .B2(n6512), .A(n5741), .ZN(n5742) );
  AOI21_X1 U6882 ( .B1(n5743), .B2(n3703), .A(n5742), .ZN(n5744) );
  OAI21_X1 U6883 ( .B1(n5745), .B2(n3703), .A(n5744), .ZN(U3001) );
  OAI21_X1 U6884 ( .B1(n3768), .B2(STATEBS16_REG_SCAN_IN), .A(n6643), .ZN(
        n5746) );
  OAI22_X1 U6885 ( .A1(n6678), .A2(n5746), .B1(n6259), .B2(n5748), .ZN(n5747)
         );
  MUX2_X1 U6886 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n5747), .S(n6535), 
        .Z(U3464) );
  XOR2_X1 U6887 ( .A(n6537), .B(n6678), .Z(n5750) );
  INV_X1 U6888 ( .A(n3210), .ZN(n5749) );
  OAI22_X1 U6889 ( .A1(n5750), .A2(n6776), .B1(n5749), .B2(n5748), .ZN(n5751)
         );
  MUX2_X1 U6890 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n5751), .S(n6535), 
        .Z(U3463) );
  INV_X1 U6891 ( .A(n6844), .ZN(n5754) );
  OAI22_X1 U6892 ( .A1(n5754), .A2(n7008), .B1(n5753), .B2(n5752), .ZN(n5755)
         );
  MUX2_X1 U6893 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n5755), .S(n7006), 
        .Z(U3456) );
  OAI21_X1 U6894 ( .B1(n5543), .B2(n5756), .A(n5588), .ZN(n6340) );
  AOI22_X1 U6895 ( .A1(PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n6491), .B1(n6523), 
        .B2(REIP_REG_15__SCAN_IN), .ZN(n5761) );
  OAI21_X1 U6896 ( .B1(n5513), .B2(n5758), .A(n5757), .ZN(n5759) );
  XOR2_X1 U6897 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .B(n5759), .Z(n6066) );
  AOI22_X1 U6898 ( .A1(n6496), .A2(n6066), .B1(n6498), .B2(n6112), .ZN(n5760)
         );
  OAI211_X1 U6899 ( .C1(n6476), .C2(n6340), .A(n5761), .B(n5760), .ZN(U2971)
         );
  OR2_X1 U6900 ( .A1(n5762), .A2(n6851), .ZN(n5763) );
  NAND2_X1 U6901 ( .A1(n6894), .A2(n5765), .ZN(n6431) );
  NOR2_X4 U6902 ( .A1(n6414), .A2(n6419), .ZN(n6411) );
  AND2_X1 U6903 ( .A1(n6411), .A2(DATAO_REG_31__SCAN_IN), .ZN(U2892) );
  NAND2_X1 U6904 ( .A1(n6365), .A2(n5216), .ZN(n5767) );
  AOI22_X1 U6905 ( .A1(EAX_REG_31__SCAN_IN), .A2(n6358), .B1(DATAI_31_), .B2(
        n6335), .ZN(n5766) );
  OAI21_X1 U6906 ( .B1(n5768), .B2(n5767), .A(n5766), .ZN(U2860) );
  INV_X1 U6907 ( .A(REIP_REG_30__SCAN_IN), .ZN(n6985) );
  INV_X1 U6908 ( .A(EBX_REG_30__SCAN_IN), .ZN(n5898) );
  OAI22_X1 U6909 ( .A1(n6245), .A2(n5898), .B1(n5769), .B2(n6266), .ZN(n5770)
         );
  AOI21_X1 U6910 ( .B1(n6261), .B2(n5771), .A(n5770), .ZN(n5772) );
  OAI21_X1 U6911 ( .B1(n5773), .B2(n6985), .A(n5772), .ZN(n5774) );
  AOI21_X1 U6912 ( .B1(n6265), .B2(n5897), .A(n5774), .ZN(n5776) );
  INV_X1 U6913 ( .A(REIP_REG_29__SCAN_IN), .ZN(n6981) );
  OR3_X1 U6914 ( .A1(n6981), .A2(n5785), .A3(REIP_REG_30__SCAN_IN), .ZN(n5775)
         );
  OAI211_X1 U6915 ( .C1(n6185), .C2(n5927), .A(n5776), .B(n5775), .ZN(U2797)
         );
  AOI22_X1 U6916 ( .A1(PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n6234), .B1(
        REIP_REG_29__SCAN_IN), .B2(n5788), .ZN(n5777) );
  OAI21_X1 U6917 ( .B1(n5778), .B2(n6267), .A(n5777), .ZN(n5779) );
  AOI21_X1 U6918 ( .B1(EBX_REG_29__SCAN_IN), .B2(n6264), .A(n5779), .ZN(n5784)
         );
  INV_X1 U6919 ( .A(n5782), .ZN(n5783) );
  OAI211_X1 U6920 ( .C1(REIP_REG_29__SCAN_IN), .C2(n5785), .A(n5784), .B(n5783), .ZN(U2798) );
  INV_X1 U6921 ( .A(n5786), .ZN(n5787) );
  AOI22_X1 U6922 ( .A1(PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n6234), .B1(n5787), 
        .B2(n6261), .ZN(n5795) );
  AOI22_X1 U6923 ( .A1(REIP_REG_28__SCAN_IN), .A2(n5788), .B1(
        EBX_REG_28__SCAN_IN), .B2(n6264), .ZN(n5794) );
  INV_X1 U6924 ( .A(n5902), .ZN(n5789) );
  OAI22_X1 U6925 ( .A1(n5790), .A2(n6185), .B1(n6236), .B2(n5789), .ZN(n5791)
         );
  INV_X1 U6926 ( .A(n5791), .ZN(n5793) );
  NAND3_X1 U6927 ( .A1(REIP_REG_27__SCAN_IN), .A2(n5801), .A3(n6978), .ZN(
        n5792) );
  NAND4_X1 U6928 ( .A1(n5795), .A2(n5794), .A3(n5793), .A4(n5792), .ZN(U2799)
         );
  OAI22_X1 U6929 ( .A1(n5818), .A2(n6972), .B1(n6245), .B2(n5905), .ZN(n5796)
         );
  AOI21_X1 U6930 ( .B1(n5956), .B2(n6261), .A(n5796), .ZN(n5803) );
  OAI21_X1 U6931 ( .B1(n5799), .B2(n5798), .A(n3195), .ZN(n5960) );
  OAI22_X1 U6932 ( .A1(n5960), .A2(n6185), .B1(n6236), .B2(n5906), .ZN(n5800)
         );
  AOI21_X1 U6933 ( .B1(n5801), .B2(n6972), .A(n5800), .ZN(n5802) );
  OAI211_X1 U6934 ( .C1(n5804), .C2(n6266), .A(n5803), .B(n5802), .ZN(U2800)
         );
  NOR2_X1 U6935 ( .A1(n6968), .A2(n5821), .ZN(n5820) );
  AOI21_X1 U6936 ( .B1(REIP_REG_25__SCAN_IN), .B2(n5820), .A(
        REIP_REG_26__SCAN_IN), .ZN(n5817) );
  INV_X1 U6937 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n5805) );
  OAI22_X1 U6938 ( .A1(n5805), .A2(n6266), .B1(n5966), .B2(n6267), .ZN(n5806)
         );
  AOI21_X1 U6939 ( .B1(EBX_REG_26__SCAN_IN), .B2(n6264), .A(n5806), .ZN(n5816)
         );
  AOI21_X1 U6940 ( .B1(n5808), .B2(n5807), .A(n5798), .ZN(n5963) );
  INV_X1 U6941 ( .A(n5809), .ZN(n5812) );
  AOI21_X1 U6942 ( .B1(n5812), .B2(n5811), .A(n5810), .ZN(n5814) );
  NOR2_X1 U6943 ( .A1(n5814), .A2(n5813), .ZN(n5998) );
  AOI22_X1 U6944 ( .A1(n5963), .A2(n6201), .B1(n6265), .B2(n5998), .ZN(n5815)
         );
  OAI211_X1 U6945 ( .C1(n5818), .C2(n5817), .A(n5816), .B(n5815), .ZN(U2801)
         );
  AOI22_X1 U6946 ( .A1(PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n6234), .B1(
        EBX_REG_25__SCAN_IN), .B2(n6264), .ZN(n5825) );
  AOI22_X1 U6947 ( .A1(n5909), .A2(n6265), .B1(n5819), .B2(n6261), .ZN(n5824)
         );
  INV_X1 U6948 ( .A(REIP_REG_25__SCAN_IN), .ZN(n6971) );
  AOI22_X1 U6949 ( .A1(n5938), .A2(n6201), .B1(n5820), .B2(n6971), .ZN(n5823)
         );
  NOR2_X1 U6950 ( .A1(REIP_REG_24__SCAN_IN), .A2(n5821), .ZN(n5828) );
  OAI21_X1 U6951 ( .B1(n5828), .B2(n5836), .A(REIP_REG_25__SCAN_IN), .ZN(n5822) );
  NAND4_X1 U6952 ( .A1(n5825), .A2(n5824), .A3(n5823), .A4(n5822), .ZN(U2802)
         );
  AOI22_X1 U6953 ( .A1(PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n6234), .B1(
        EBX_REG_24__SCAN_IN), .B2(n6264), .ZN(n5832) );
  AOI22_X1 U6954 ( .A1(n5826), .A2(n6261), .B1(REIP_REG_24__SCAN_IN), .B2(
        n5836), .ZN(n5831) );
  INV_X1 U6955 ( .A(n5912), .ZN(n5827) );
  AOI22_X1 U6956 ( .A1(n5941), .A2(n6201), .B1(n6265), .B2(n5827), .ZN(n5830)
         );
  INV_X1 U6957 ( .A(n5828), .ZN(n5829) );
  NAND4_X1 U6958 ( .A1(n5832), .A2(n5831), .A3(n5830), .A4(n5829), .ZN(U2803)
         );
  AOI22_X1 U6959 ( .A1(PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n6234), .B1(n5833), 
        .B2(n6261), .ZN(n5838) );
  INV_X1 U6960 ( .A(n5847), .ZN(n5859) );
  OAI21_X1 U6961 ( .B1(n5859), .B2(n5846), .A(n6967), .ZN(n5835) );
  OAI22_X1 U6962 ( .A1(n5946), .A2(n6185), .B1(n6236), .B2(n5916), .ZN(n5834)
         );
  AOI21_X1 U6963 ( .B1(n5836), .B2(n5835), .A(n5834), .ZN(n5837) );
  OAI211_X1 U6964 ( .C1(n6245), .C2(n5915), .A(n5838), .B(n5837), .ZN(U2804)
         );
  AOI22_X1 U6965 ( .A1(PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n6234), .B1(
        EBX_REG_22__SCAN_IN), .B2(n6264), .ZN(n5851) );
  INV_X1 U6966 ( .A(n5839), .ZN(n5841) );
  INV_X1 U6967 ( .A(n5869), .ZN(n5840) );
  AOI22_X1 U6968 ( .A1(n5841), .A2(n6261), .B1(REIP_REG_22__SCAN_IN), .B2(
        n5840), .ZN(n5850) );
  NOR2_X1 U6969 ( .A1(n5724), .A2(n5842), .ZN(n5843) );
  OR2_X1 U6970 ( .A1(n5844), .A2(n5843), .ZN(n5918) );
  OAI22_X1 U6971 ( .A1(n5917), .A2(n6185), .B1(n6236), .B2(n5918), .ZN(n5845)
         );
  INV_X1 U6972 ( .A(n5845), .ZN(n5849) );
  OAI211_X1 U6973 ( .C1(REIP_REG_22__SCAN_IN), .C2(REIP_REG_21__SCAN_IN), .A(
        n5847), .B(n5846), .ZN(n5848) );
  NAND4_X1 U6974 ( .A1(n5851), .A2(n5850), .A3(n5849), .A4(n5848), .ZN(U2805)
         );
  AOI22_X1 U6975 ( .A1(n5967), .A2(n6261), .B1(EBX_REG_21__SCAN_IN), .B2(n6264), .ZN(n5852) );
  OAI21_X1 U6976 ( .B1(n5869), .B2(n5728), .A(n5852), .ZN(n5857) );
  OAI21_X1 U6977 ( .B1(n5855), .B2(n5854), .A(n4039), .ZN(n5971) );
  OAI22_X1 U6978 ( .A1(n5971), .A2(n6185), .B1(n6236), .B2(n5921), .ZN(n5856)
         );
  AOI211_X1 U6979 ( .C1(PHYADDRPOINTER_REG_21__SCAN_IN), .C2(n6234), .A(n5857), 
        .B(n5856), .ZN(n5858) );
  OAI21_X1 U6980 ( .B1(REIP_REG_21__SCAN_IN), .B2(n5859), .A(n5858), .ZN(U2806) );
  AOI22_X1 U6981 ( .A1(PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n6234), .B1(
        EBX_REG_20__SCAN_IN), .B2(n6264), .ZN(n5873) );
  AOI21_X1 U6982 ( .B1(n5861), .B2(n5875), .A(n5854), .ZN(n5976) );
  INV_X1 U6983 ( .A(n5862), .ZN(n6115) );
  AOI21_X1 U6984 ( .B1(n6115), .B2(n5863), .A(REIP_REG_20__SCAN_IN), .ZN(n5870) );
  MUX2_X1 U6985 ( .A(n5866), .B(n3203), .S(n5864), .Z(n5867) );
  XOR2_X1 U6986 ( .A(n5868), .B(n5867), .Z(n6016) );
  OAI22_X1 U6987 ( .A1(n5870), .A2(n5869), .B1(n6016), .B2(n6236), .ZN(n5871)
         );
  AOI21_X1 U6988 ( .B1(n5976), .B2(n6201), .A(n5871), .ZN(n5872) );
  OAI211_X1 U6989 ( .C1(n5979), .C2(n6267), .A(n5873), .B(n5872), .ZN(U2807)
         );
  OAI21_X1 U6990 ( .B1(n5876), .B2(n5874), .A(n5875), .ZN(n5984) );
  NAND2_X1 U6991 ( .A1(n5878), .A2(n5877), .ZN(n6033) );
  NAND2_X1 U6992 ( .A1(n5564), .A2(n6033), .ZN(n5879) );
  XOR2_X1 U6993 ( .A(n5880), .B(n5879), .Z(n6027) );
  AOI22_X1 U6994 ( .A1(n5981), .A2(n6261), .B1(EBX_REG_19__SCAN_IN), .B2(n6264), .ZN(n5881) );
  OAI211_X1 U6995 ( .C1(n6266), .C2(n5882), .A(n5881), .B(n3179), .ZN(n5883)
         );
  AOI21_X1 U6996 ( .B1(n6265), .B2(n6027), .A(n5883), .ZN(n5888) );
  NOR2_X1 U6997 ( .A1(n6958), .A2(n6962), .ZN(n5885) );
  NAND2_X1 U6998 ( .A1(REIP_REG_17__SCAN_IN), .A2(n5884), .ZN(n6104) );
  OAI22_X1 U6999 ( .A1(n5885), .A2(n6104), .B1(n6099), .B2(n6962), .ZN(n5886)
         );
  OAI21_X1 U7000 ( .B1(REIP_REG_18__SCAN_IN), .B2(REIP_REG_19__SCAN_IN), .A(
        n5886), .ZN(n5887) );
  OAI211_X1 U7001 ( .C1(n5984), .C2(n6185), .A(n5888), .B(n5887), .ZN(U2808)
         );
  NAND2_X1 U7002 ( .A1(n5890), .A2(n5889), .ZN(n5896) );
  INV_X1 U7003 ( .A(n5891), .ZN(n5894) );
  INV_X1 U7004 ( .A(n3410), .ZN(n5893) );
  NAND4_X1 U7005 ( .A1(n5894), .A2(n6250), .A3(n5893), .A4(n5892), .ZN(n5895)
         );
  INV_X1 U7006 ( .A(n5897), .ZN(n5899) );
  OAI222_X1 U7007 ( .A1(n6321), .A2(n5927), .B1(n6320), .B2(n5899), .C1(n5898), 
        .C2(n6317), .ZN(U2829) );
  AOI22_X1 U7008 ( .A1(EBX_REG_29__SCAN_IN), .A2(n6324), .B1(n5900), .B2(n6323), .ZN(n5901) );
  OAI21_X1 U7009 ( .B1(n5930), .B2(n6321), .A(n5901), .ZN(U2830) );
  AOI22_X1 U7010 ( .A1(n5931), .A2(n6325), .B1(n5902), .B2(n6323), .ZN(n5903)
         );
  OAI21_X1 U7011 ( .B1(n5904), .B2(n6317), .A(n5903), .ZN(U2831) );
  OAI222_X1 U7012 ( .A1(n6320), .A2(n5906), .B1(n6317), .B2(n5905), .C1(n6321), 
        .C2(n5960), .ZN(U2832) );
  AOI22_X1 U7013 ( .A1(n5963), .A2(n6325), .B1(n5998), .B2(n6323), .ZN(n5907)
         );
  OAI21_X1 U7014 ( .B1(n5908), .B2(n6317), .A(n5907), .ZN(U2833) );
  INV_X1 U7015 ( .A(n5938), .ZN(n5911) );
  AOI22_X1 U7016 ( .A1(EBX_REG_25__SCAN_IN), .A2(n6324), .B1(n5909), .B2(n6323), .ZN(n5910) );
  OAI21_X1 U7017 ( .B1(n5911), .B2(n6321), .A(n5910), .ZN(U2834) );
  INV_X1 U7018 ( .A(n5941), .ZN(n5914) );
  OAI222_X1 U7019 ( .A1(n6321), .A2(n5914), .B1(n6317), .B2(n5913), .C1(n5912), 
        .C2(n6320), .ZN(U2835) );
  OAI222_X1 U7020 ( .A1(n6320), .A2(n5916), .B1(n6317), .B2(n5915), .C1(n6321), 
        .C2(n5946), .ZN(U2836) );
  INV_X1 U7021 ( .A(n5917), .ZN(n5947) );
  INV_X1 U7022 ( .A(n5918), .ZN(n6008) );
  AOI22_X1 U7023 ( .A1(EBX_REG_22__SCAN_IN), .A2(n6324), .B1(n6008), .B2(n6323), .ZN(n5919) );
  OAI21_X1 U7024 ( .B1(n5917), .B2(n6321), .A(n5919), .ZN(U2837) );
  INV_X1 U7025 ( .A(EBX_REG_21__SCAN_IN), .ZN(n5920) );
  OAI222_X1 U7026 ( .A1(n6320), .A2(n5921), .B1(n6317), .B2(n5920), .C1(n6321), 
        .C2(n5971), .ZN(U2838) );
  INV_X1 U7027 ( .A(n5976), .ZN(n5923) );
  OAI222_X1 U7028 ( .A1(n6321), .A2(n5923), .B1(n6320), .B2(n6016), .C1(n5922), 
        .C2(n6317), .ZN(U2839) );
  AOI22_X1 U7029 ( .A1(EBX_REG_19__SCAN_IN), .A2(n6324), .B1(n6323), .B2(n6027), .ZN(n5924) );
  OAI21_X1 U7030 ( .B1(n6321), .B2(n5984), .A(n5924), .ZN(U2840) );
  AOI22_X1 U7031 ( .A1(DATAI_30_), .A2(n6335), .B1(DATAI_14_), .B2(n6336), 
        .ZN(n5926) );
  NAND2_X1 U7032 ( .A1(EAX_REG_30__SCAN_IN), .A2(n6358), .ZN(n5925) );
  OAI211_X1 U7033 ( .C1(n5927), .C2(n6368), .A(n5926), .B(n5925), .ZN(U2861)
         );
  AOI22_X1 U7034 ( .A1(DATAI_29_), .A2(n6335), .B1(n6336), .B2(DATAI_13_), 
        .ZN(n5929) );
  NAND2_X1 U7035 ( .A1(EAX_REG_29__SCAN_IN), .A2(n6358), .ZN(n5928) );
  OAI211_X1 U7036 ( .C1(n6368), .C2(n5930), .A(n5929), .B(n5928), .ZN(U2862)
         );
  AOI22_X1 U7037 ( .A1(n5931), .A2(n6360), .B1(n6335), .B2(DATAI_28_), .ZN(
        n5933) );
  AOI22_X1 U7038 ( .A1(EAX_REG_28__SCAN_IN), .A2(n6358), .B1(n6336), .B2(
        DATAI_12_), .ZN(n5932) );
  NAND2_X1 U7039 ( .A1(n5933), .A2(n5932), .ZN(U2863) );
  AOI22_X1 U7040 ( .A1(EAX_REG_27__SCAN_IN), .A2(n6358), .B1(n6335), .B2(
        DATAI_27_), .ZN(n5935) );
  NAND2_X1 U7041 ( .A1(n6336), .A2(DATAI_11_), .ZN(n5934) );
  OAI211_X1 U7042 ( .C1(n6368), .C2(n5960), .A(n5935), .B(n5934), .ZN(U2864)
         );
  AOI22_X1 U7043 ( .A1(DATAI_26_), .A2(n6335), .B1(n5963), .B2(n6360), .ZN(
        n5937) );
  AOI22_X1 U7044 ( .A1(EAX_REG_26__SCAN_IN), .A2(n6358), .B1(n6336), .B2(
        DATAI_10_), .ZN(n5936) );
  NAND2_X1 U7045 ( .A1(n5937), .A2(n5936), .ZN(U2865) );
  AOI22_X1 U7046 ( .A1(DATAI_25_), .A2(n6335), .B1(n5938), .B2(n6360), .ZN(
        n5940) );
  AOI22_X1 U7047 ( .A1(EAX_REG_25__SCAN_IN), .A2(n6358), .B1(DATAI_9_), .B2(
        n6336), .ZN(n5939) );
  NAND2_X1 U7048 ( .A1(n5940), .A2(n5939), .ZN(U2866) );
  AOI22_X1 U7049 ( .A1(DATAI_24_), .A2(n6335), .B1(n5941), .B2(n6360), .ZN(
        n5943) );
  AOI22_X1 U7050 ( .A1(EAX_REG_24__SCAN_IN), .A2(n6358), .B1(n6336), .B2(
        DATAI_8_), .ZN(n5942) );
  NAND2_X1 U7051 ( .A1(n5943), .A2(n5942), .ZN(U2867) );
  AOI22_X1 U7052 ( .A1(n6335), .A2(DATAI_23_), .B1(n6336), .B2(DATAI_7_), .ZN(
        n5945) );
  NAND2_X1 U7053 ( .A1(EAX_REG_23__SCAN_IN), .A2(n6358), .ZN(n5944) );
  OAI211_X1 U7054 ( .C1(n6368), .C2(n5946), .A(n5945), .B(n5944), .ZN(U2868)
         );
  AOI22_X1 U7055 ( .A1(n5947), .A2(n6360), .B1(n6335), .B2(DATAI_22_), .ZN(
        n5949) );
  AOI22_X1 U7056 ( .A1(EAX_REG_22__SCAN_IN), .A2(n6358), .B1(DATAI_6_), .B2(
        n6336), .ZN(n5948) );
  NAND2_X1 U7057 ( .A1(n5949), .A2(n5948), .ZN(U2869) );
  AOI22_X1 U7058 ( .A1(n6335), .A2(DATAI_21_), .B1(n6336), .B2(DATAI_5_), .ZN(
        n5951) );
  NAND2_X1 U7059 ( .A1(EAX_REG_21__SCAN_IN), .A2(n6358), .ZN(n5950) );
  OAI211_X1 U7060 ( .C1(n6368), .C2(n5971), .A(n5951), .B(n5950), .ZN(U2870)
         );
  AOI22_X1 U7061 ( .A1(n5976), .A2(n6360), .B1(n6335), .B2(DATAI_20_), .ZN(
        n5953) );
  AOI22_X1 U7062 ( .A1(EAX_REG_20__SCAN_IN), .A2(n6358), .B1(n6336), .B2(
        DATAI_4_), .ZN(n5952) );
  NAND2_X1 U7063 ( .A1(n5953), .A2(n5952), .ZN(U2871) );
  AOI22_X1 U7064 ( .A1(EAX_REG_19__SCAN_IN), .A2(n6358), .B1(n6335), .B2(
        DATAI_19_), .ZN(n5955) );
  NAND2_X1 U7065 ( .A1(n6336), .A2(DATAI_3_), .ZN(n5954) );
  OAI211_X1 U7066 ( .C1(n5984), .C2(n6368), .A(n5955), .B(n5954), .ZN(U2872)
         );
  AOI22_X1 U7067 ( .A1(PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n6491), .B1(n6523), 
        .B2(REIP_REG_27__SCAN_IN), .ZN(n5959) );
  AOI22_X1 U7068 ( .A1(n6496), .A2(n5957), .B1(n6498), .B2(n5956), .ZN(n5958)
         );
  OAI211_X1 U7069 ( .C1(n6476), .C2(n5960), .A(n5959), .B(n5958), .ZN(U2959)
         );
  AOI22_X1 U7070 ( .A1(PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n6491), .B1(n6523), 
        .B2(REIP_REG_26__SCAN_IN), .ZN(n5965) );
  XNOR2_X1 U7071 ( .A(n3704), .B(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5961)
         );
  XNOR2_X1 U7072 ( .A(n5962), .B(n5961), .ZN(n5997) );
  AOI22_X1 U7073 ( .A1(n5963), .A2(n5989), .B1(n6496), .B2(n5997), .ZN(n5964)
         );
  OAI211_X1 U7074 ( .C1(n6490), .C2(n5966), .A(n5965), .B(n5964), .ZN(U2960)
         );
  AOI22_X1 U7075 ( .A1(PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n6491), .B1(n6523), 
        .B2(REIP_REG_21__SCAN_IN), .ZN(n5970) );
  AOI22_X1 U7076 ( .A1(n5968), .A2(n6496), .B1(n6498), .B2(n5967), .ZN(n5969)
         );
  OAI211_X1 U7077 ( .C1(n6476), .C2(n5971), .A(n5970), .B(n5969), .ZN(U2965)
         );
  AOI22_X1 U7078 ( .A1(PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n6491), .B1(n6523), 
        .B2(REIP_REG_20__SCAN_IN), .ZN(n5978) );
  NAND2_X1 U7079 ( .A1(n5973), .A2(n5972), .ZN(n5974) );
  AND2_X1 U7080 ( .A1(n5975), .A2(n5974), .ZN(n6019) );
  AOI22_X1 U7081 ( .A1(n5976), .A2(n5989), .B1(n6496), .B2(n6019), .ZN(n5977)
         );
  OAI211_X1 U7082 ( .C1(n6490), .C2(n5979), .A(n5978), .B(n5977), .ZN(U2966)
         );
  AOI22_X1 U7083 ( .A1(PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n6491), .B1(n6523), 
        .B2(REIP_REG_19__SCAN_IN), .ZN(n5983) );
  XNOR2_X1 U7084 ( .A(n4222), .B(n5980), .ZN(n6028) );
  AOI22_X1 U7085 ( .A1(n6028), .A2(n6496), .B1(n6498), .B2(n5981), .ZN(n5982)
         );
  OAI211_X1 U7086 ( .C1(n6476), .C2(n5984), .A(n5983), .B(n5982), .ZN(U2967)
         );
  AOI22_X1 U7087 ( .A1(PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n6491), .B1(n6523), 
        .B2(REIP_REG_18__SCAN_IN), .ZN(n5991) );
  OAI21_X1 U7088 ( .B1(INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n5986), .A(n5985), 
        .ZN(n5987) );
  XOR2_X1 U7089 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .B(n5987), .Z(n6035) );
  AOI21_X1 U7090 ( .B1(n5988), .B2(n5568), .A(n5874), .ZN(n6328) );
  AOI22_X1 U7091 ( .A1(n6496), .A2(n6035), .B1(n5989), .B2(n6328), .ZN(n5990)
         );
  OAI211_X1 U7092 ( .C1(n6490), .C2(n6098), .A(n5991), .B(n5990), .ZN(U2968)
         );
  AOI22_X1 U7093 ( .A1(PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n6491), .B1(n6523), 
        .B2(REIP_REG_17__SCAN_IN), .ZN(n5995) );
  AOI22_X1 U7094 ( .A1(n6496), .A2(n5993), .B1(n6498), .B2(n5992), .ZN(n5994)
         );
  OAI211_X1 U7095 ( .C1(n6476), .C2(n6282), .A(n5995), .B(n5994), .ZN(U2969)
         );
  AOI22_X1 U7096 ( .A1(n5997), .A2(n6528), .B1(INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n5996), .ZN(n6004) );
  NAND2_X1 U7097 ( .A1(n6523), .A2(REIP_REG_26__SCAN_IN), .ZN(n6003) );
  NAND2_X1 U7098 ( .A1(n5998), .A2(n6525), .ZN(n6002) );
  OAI211_X1 U7099 ( .C1(INSTADDRPOINTER_REG_26__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_25__SCAN_IN), .A(n6000), .B(n5999), .ZN(n6001) );
  NAND4_X1 U7100 ( .A1(n6004), .A2(n6003), .A3(n6002), .A4(n6001), .ZN(U2992)
         );
  INV_X1 U7101 ( .A(n6005), .ZN(n6007) );
  AOI22_X1 U7102 ( .A1(n6007), .A2(n6528), .B1(INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n6006), .ZN(n6015) );
  NAND2_X1 U7103 ( .A1(n6523), .A2(REIP_REG_22__SCAN_IN), .ZN(n6014) );
  NAND2_X1 U7104 ( .A1(n6008), .A2(n6525), .ZN(n6013) );
  NAND3_X1 U7105 ( .A1(n6011), .A2(n6010), .A3(n6009), .ZN(n6012) );
  NAND4_X1 U7106 ( .A1(n6015), .A2(n6014), .A3(n6013), .A4(n6012), .ZN(U2996)
         );
  INV_X1 U7107 ( .A(REIP_REG_20__SCAN_IN), .ZN(n6960) );
  AOI21_X1 U7108 ( .B1(n6021), .B2(n6530), .A(n6037), .ZN(n6032) );
  OAI22_X1 U7109 ( .A1(n6032), .A2(n6017), .B1(n6016), .B2(n6512), .ZN(n6018)
         );
  AOI21_X1 U7110 ( .B1(n6019), .B2(n6528), .A(n6018), .ZN(n6025) );
  NOR3_X1 U7111 ( .A1(n6021), .A2(n6020), .A3(n6047), .ZN(n6026) );
  NAND3_X1 U7112 ( .A1(n6026), .A2(n6023), .A3(n6022), .ZN(n6024) );
  OAI211_X1 U7113 ( .C1(n6960), .C2(n3179), .A(n6025), .B(n6024), .ZN(U2998)
         );
  AOI22_X1 U7114 ( .A1(REIP_REG_19__SCAN_IN), .A2(n6523), .B1(n6026), .B2(
        n6031), .ZN(n6030) );
  AOI22_X1 U7115 ( .A1(n6028), .A2(n6528), .B1(n6525), .B2(n6027), .ZN(n6029)
         );
  OAI211_X1 U7116 ( .C1(n6032), .C2(n6031), .A(n6030), .B(n6029), .ZN(U2999)
         );
  XNOR2_X1 U7117 ( .A(n6034), .B(n6033), .ZN(n6277) );
  AOI22_X1 U7118 ( .A1(n6035), .A2(n6528), .B1(n6525), .B2(n6277), .ZN(n6042)
         );
  NAND2_X1 U7119 ( .A1(n6523), .A2(REIP_REG_18__SCAN_IN), .ZN(n6041) );
  OAI221_X1 U7120 ( .B1(n6037), .B2(n6036), .C1(n6037), .C2(n3703), .A(
        INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n6040) );
  NAND3_X1 U7121 ( .A1(n6038), .A2(n3702), .A3(n6045), .ZN(n6039) );
  NAND4_X1 U7122 ( .A1(n6042), .A2(n6041), .A3(n6040), .A4(n6039), .ZN(U3000)
         );
  NAND2_X1 U7123 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n6046), .ZN(n6044) );
  AOI21_X1 U7124 ( .B1(n6044), .B2(n6530), .A(n6043), .ZN(n6064) );
  INV_X1 U7125 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n6063) );
  NAND4_X1 U7126 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n6046), .A3(n6063), .A4(n6045), .ZN(n6067) );
  NOR2_X1 U7127 ( .A1(INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n6047), .ZN(n6055)
         );
  NOR2_X1 U7128 ( .A1(n3179), .A2(n6955), .ZN(n6054) );
  OR2_X1 U7129 ( .A1(n6061), .A2(n6048), .ZN(n6049) );
  NAND2_X1 U7130 ( .A1(n6050), .A2(n6049), .ZN(n6283) );
  OAI22_X1 U7131 ( .A1(n6052), .A2(n6051), .B1(n6512), .B2(n6283), .ZN(n6053)
         );
  AOI211_X1 U7132 ( .C1(n6056), .C2(n6055), .A(n6054), .B(n6053), .ZN(n6057)
         );
  OAI221_X1 U7133 ( .B1(n6058), .B2(n6064), .C1(n6058), .C2(n6067), .A(n6057), 
        .ZN(U3002) );
  AND2_X1 U7134 ( .A1(n6060), .A2(n6059), .ZN(n6062) );
  OR2_X1 U7135 ( .A1(n6062), .A2(n6061), .ZN(n6286) );
  OAI22_X1 U7136 ( .A1(n6064), .A2(n6063), .B1(n6512), .B2(n6286), .ZN(n6065)
         );
  AOI21_X1 U7137 ( .B1(n6528), .B2(n6066), .A(n6065), .ZN(n6068) );
  OAI211_X1 U7138 ( .C1(n6953), .C2(n3179), .A(n6068), .B(n6067), .ZN(U3003)
         );
  OR2_X1 U7139 ( .A1(n6069), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6071) );
  OAI22_X1 U7140 ( .A1(n6072), .A2(n6071), .B1(n6070), .B2(n7006), .ZN(U3455)
         );
  INV_X1 U7141 ( .A(STATE_REG_0__SCAN_IN), .ZN(n6919) );
  AOI21_X1 U7142 ( .B1(STATE_REG_1__SCAN_IN), .B2(n6073), .A(n6919), .ZN(n6079) );
  INV_X1 U7143 ( .A(ADS_N_REG_SCAN_IN), .ZN(n6074) );
  NOR2_X2 U7144 ( .A1(STATE_REG_0__SCAN_IN), .A2(n6918), .ZN(n7032) );
  AOI21_X1 U7145 ( .B1(n6079), .B2(n6074), .A(n7032), .ZN(U2789) );
  INV_X1 U7146 ( .A(n6075), .ZN(n6076) );
  OAI22_X1 U7147 ( .A1(n6891), .A2(n6199), .B1(n4783), .B2(n6076), .ZN(n6082)
         );
  OAI21_X1 U7148 ( .B1(n6082), .B2(n6901), .A(CODEFETCH_REG_SCAN_IN), .ZN(
        n6077) );
  OAI21_X1 U7149 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6902), .A(n6077), .ZN(
        U2790) );
  INV_X2 U7150 ( .A(n7032), .ZN(n7019) );
  NOR2_X1 U7151 ( .A1(STATE_REG_2__SCAN_IN), .A2(STATE_REG_0__SCAN_IN), .ZN(
        n6080) );
  OAI21_X1 U7152 ( .B1(D_C_N_REG_SCAN_IN), .B2(n6080), .A(n7019), .ZN(n6078)
         );
  OAI21_X1 U7153 ( .B1(CODEFETCH_REG_SCAN_IN), .B2(n7019), .A(n6078), .ZN(
        U2791) );
  NOR2_X1 U7154 ( .A1(n7032), .A2(n6079), .ZN(n6997) );
  OAI21_X1 U7155 ( .B1(BS16_N), .B2(n6080), .A(n6997), .ZN(n6995) );
  OAI21_X1 U7156 ( .B1(n6997), .B2(n6081), .A(n6995), .ZN(U2792) );
  NAND2_X1 U7157 ( .A1(n7026), .A2(n3422), .ZN(n7035) );
  AOI21_X1 U7158 ( .B1(n7035), .B2(n6917), .A(READY_N), .ZN(n7025) );
  NOR2_X1 U7159 ( .A1(n6082), .A2(n7025), .ZN(n6866) );
  NOR2_X1 U7160 ( .A1(n6866), .A2(n6901), .ZN(n7020) );
  OAI21_X1 U7161 ( .B1(n7020), .B2(n6083), .A(n6484), .ZN(U2793) );
  NOR4_X1 U7162 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(
        DATAWIDTH_REG_18__SCAN_IN), .A3(DATAWIDTH_REG_20__SCAN_IN), .A4(
        DATAWIDTH_REG_21__SCAN_IN), .ZN(n6087) );
  NOR4_X1 U7163 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(
        DATAWIDTH_REG_14__SCAN_IN), .A3(DATAWIDTH_REG_15__SCAN_IN), .A4(
        DATAWIDTH_REG_16__SCAN_IN), .ZN(n6086) );
  NOR4_X1 U7164 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(
        DATAWIDTH_REG_27__SCAN_IN), .A3(DATAWIDTH_REG_28__SCAN_IN), .A4(
        DATAWIDTH_REG_30__SCAN_IN), .ZN(n6085) );
  NOR4_X1 U7165 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(
        DATAWIDTH_REG_23__SCAN_IN), .A3(DATAWIDTH_REG_24__SCAN_IN), .A4(
        DATAWIDTH_REG_25__SCAN_IN), .ZN(n6084) );
  NAND4_X1 U7166 ( .A1(n6087), .A2(n6086), .A3(n6085), .A4(n6084), .ZN(n6093)
         );
  NOR4_X1 U7167 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(DATAWIDTH_REG_3__SCAN_IN), 
        .A3(DATAWIDTH_REG_31__SCAN_IN), .A4(DATAWIDTH_REG_2__SCAN_IN), .ZN(
        n6091) );
  AOI211_X1 U7168 ( .C1(DATAWIDTH_REG_0__SCAN_IN), .C2(
        DATAWIDTH_REG_1__SCAN_IN), .A(DATAWIDTH_REG_19__SCAN_IN), .B(
        DATAWIDTH_REG_29__SCAN_IN), .ZN(n6090) );
  NOR4_X1 U7169 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(DATAWIDTH_REG_10__SCAN_IN), .A3(DATAWIDTH_REG_11__SCAN_IN), .A4(DATAWIDTH_REG_12__SCAN_IN), .ZN(n6089)
         );
  NOR4_X1 U7170 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(DATAWIDTH_REG_6__SCAN_IN), 
        .A3(DATAWIDTH_REG_7__SCAN_IN), .A4(DATAWIDTH_REG_8__SCAN_IN), .ZN(
        n6088) );
  NAND4_X1 U7171 ( .A1(n6091), .A2(n6090), .A3(n6089), .A4(n6088), .ZN(n6092)
         );
  NOR2_X1 U7172 ( .A1(n6093), .A2(n6092), .ZN(n7013) );
  INV_X1 U7173 ( .A(BYTEENABLE_REG_1__SCAN_IN), .ZN(n6990) );
  NOR3_X1 U7174 ( .A1(DATAWIDTH_REG_0__SCAN_IN), .A2(REIP_REG_0__SCAN_IN), 
        .A3(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6095) );
  OAI21_X1 U7175 ( .B1(REIP_REG_1__SCAN_IN), .B2(n6095), .A(n7013), .ZN(n6094)
         );
  OAI21_X1 U7176 ( .B1(n7013), .B2(n6990), .A(n6094), .ZN(U2794) );
  INV_X1 U7177 ( .A(REIP_REG_1__SCAN_IN), .ZN(n7015) );
  INV_X1 U7178 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6996) );
  AOI21_X1 U7179 ( .B1(n7015), .B2(n6996), .A(n6095), .ZN(n6096) );
  INV_X1 U7180 ( .A(BYTEENABLE_REG_3__SCAN_IN), .ZN(n6988) );
  INV_X1 U7181 ( .A(n7013), .ZN(n7016) );
  AOI22_X1 U7182 ( .A1(n7013), .A2(n6096), .B1(n6988), .B2(n7016), .ZN(U2795)
         );
  INV_X1 U7183 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n6097) );
  OAI21_X1 U7184 ( .B1(n6266), .B2(n6097), .A(n3179), .ZN(n6101) );
  OAI22_X1 U7185 ( .A1(n6099), .A2(n6958), .B1(n6098), .B2(n6267), .ZN(n6100)
         );
  AOI211_X1 U7186 ( .C1(EBX_REG_18__SCAN_IN), .C2(n6264), .A(n6101), .B(n6100), 
        .ZN(n6103) );
  AOI22_X1 U7187 ( .A1(n6328), .A2(n6201), .B1(n6265), .B2(n6277), .ZN(n6102)
         );
  OAI211_X1 U7188 ( .C1(REIP_REG_18__SCAN_IN), .C2(n6104), .A(n6103), .B(n6102), .ZN(U2809) );
  INV_X1 U7189 ( .A(n6334), .ZN(n6285) );
  OAI21_X1 U7190 ( .B1(n6266), .B2(n6105), .A(n3179), .ZN(n6107) );
  OAI22_X1 U7191 ( .A1(n6245), .A2(n6284), .B1(n6236), .B2(n6283), .ZN(n6106)
         );
  AOI211_X1 U7192 ( .C1(n6108), .C2(n6261), .A(n6107), .B(n6106), .ZN(n6111)
         );
  XNOR2_X1 U7193 ( .A(REIP_REG_16__SCAN_IN), .B(n6953), .ZN(n6109) );
  AOI22_X1 U7194 ( .A1(REIP_REG_16__SCAN_IN), .A2(n6121), .B1(n6115), .B2(
        n6109), .ZN(n6110) );
  OAI211_X1 U7195 ( .C1(n6185), .C2(n6285), .A(n6111), .B(n6110), .ZN(U2811)
         );
  AOI22_X1 U7196 ( .A1(n6112), .A2(n6261), .B1(EBX_REG_15__SCAN_IN), .B2(n6264), .ZN(n6117) );
  AOI22_X1 U7197 ( .A1(PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n6234), .B1(
        REIP_REG_15__SCAN_IN), .B2(n6121), .ZN(n6113) );
  OAI211_X1 U7198 ( .C1(n6236), .C2(n6286), .A(n6113), .B(n3179), .ZN(n6114)
         );
  AOI21_X1 U7199 ( .B1(n6115), .B2(n6953), .A(n6114), .ZN(n6116) );
  OAI211_X1 U7200 ( .C1(n6185), .C2(n6340), .A(n6117), .B(n6116), .ZN(U2812)
         );
  OAI22_X1 U7201 ( .A1(n6236), .A2(n6289), .B1(n6118), .B2(n6266), .ZN(n6119)
         );
  AOI21_X1 U7202 ( .B1(EBX_REG_14__SCAN_IN), .B2(n6264), .A(n6119), .ZN(n6125)
         );
  AOI22_X1 U7203 ( .A1(n6120), .A2(n6261), .B1(n6201), .B2(n6288), .ZN(n6124)
         );
  OAI21_X1 U7204 ( .B1(REIP_REG_14__SCAN_IN), .B2(n6122), .A(n6121), .ZN(n6123) );
  NAND4_X1 U7205 ( .A1(n6125), .A2(n6124), .A3(n3179), .A4(n6123), .ZN(U2813)
         );
  NAND2_X1 U7206 ( .A1(n6126), .A2(n6948), .ZN(n6138) );
  AOI22_X1 U7207 ( .A1(n6265), .A2(n6291), .B1(n6264), .B2(EBX_REG_13__SCAN_IN), .ZN(n6127) );
  OAI211_X1 U7208 ( .C1(n6266), .C2(n6128), .A(n6127), .B(n3179), .ZN(n6131)
         );
  INV_X1 U7209 ( .A(n6292), .ZN(n6344) );
  OAI22_X1 U7210 ( .A1(REIP_REG_13__SCAN_IN), .A2(n6129), .B1(n6344), .B2(
        n6185), .ZN(n6130) );
  AOI211_X1 U7211 ( .C1(n6132), .C2(n6261), .A(n6131), .B(n6130), .ZN(n6133)
         );
  OAI221_X1 U7212 ( .B1(n6950), .B2(n6141), .C1(n6950), .C2(n6138), .A(n6133), 
        .ZN(U2814) );
  OAI22_X1 U7213 ( .A1(n6245), .A2(n6296), .B1(n6948), .B2(n6141), .ZN(n6137)
         );
  AOI22_X1 U7214 ( .A1(n6261), .A2(n6134), .B1(n6265), .B2(n6294), .ZN(n6135)
         );
  OAI211_X1 U7215 ( .C1(n6266), .C2(n5507), .A(n6135), .B(n3179), .ZN(n6136)
         );
  AOI211_X1 U7216 ( .C1(n6201), .C2(n6345), .A(n6137), .B(n6136), .ZN(n6139)
         );
  NAND2_X1 U7217 ( .A1(n6139), .A2(n6138), .ZN(U2815) );
  AOI21_X1 U7218 ( .B1(n6945), .B2(n6142), .A(n6141), .ZN(n6146) );
  AOI22_X1 U7219 ( .A1(n6265), .A2(n3222), .B1(n6264), .B2(EBX_REG_11__SCAN_IN), .ZN(n6143) );
  OAI211_X1 U7220 ( .C1(n6266), .C2(n6144), .A(n6143), .B(n3179), .ZN(n6145)
         );
  AOI211_X1 U7221 ( .C1(n6261), .C2(n6147), .A(n6146), .B(n6145), .ZN(n6148)
         );
  OAI21_X1 U7222 ( .B1(n6185), .B2(n6349), .A(n6148), .ZN(U2816) );
  INV_X1 U7223 ( .A(n6149), .ZN(n6351) );
  AOI22_X1 U7224 ( .A1(n6151), .A2(n6261), .B1(n6150), .B2(n6943), .ZN(n6158)
         );
  INV_X1 U7225 ( .A(n6270), .ZN(n6153) );
  NOR2_X1 U7226 ( .A1(n6153), .A2(n6152), .ZN(n6172) );
  NOR2_X1 U7227 ( .A1(REIP_REG_9__SCAN_IN), .A2(n6154), .ZN(n6166) );
  AOI22_X1 U7228 ( .A1(PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n6234), .B1(
        EBX_REG_10__SCAN_IN), .B2(n6264), .ZN(n6155) );
  OAI211_X1 U7229 ( .C1(n6236), .C2(n6298), .A(n6155), .B(n3179), .ZN(n6156)
         );
  AOI221_X1 U7230 ( .B1(n6172), .B2(REIP_REG_10__SCAN_IN), .C1(n6166), .C2(
        REIP_REG_10__SCAN_IN), .A(n6156), .ZN(n6157) );
  OAI211_X1 U7231 ( .C1(n6185), .C2(n6351), .A(n6158), .B(n6157), .ZN(U2817)
         );
  INV_X1 U7232 ( .A(n6159), .ZN(n6160) );
  AOI21_X1 U7233 ( .B1(n6162), .B2(n6161), .A(n6160), .ZN(n6504) );
  AOI22_X1 U7234 ( .A1(n6265), .A2(n6504), .B1(n6264), .B2(EBX_REG_9__SCAN_IN), 
        .ZN(n6163) );
  OAI211_X1 U7235 ( .C1(n6266), .C2(n6164), .A(n6163), .B(n3179), .ZN(n6165)
         );
  AOI211_X1 U7236 ( .C1(n6172), .C2(REIP_REG_9__SCAN_IN), .A(n6166), .B(n6165), 
        .ZN(n6169) );
  AOI22_X1 U7237 ( .A1(n6167), .A2(n6261), .B1(n6201), .B2(n6352), .ZN(n6168)
         );
  NAND2_X1 U7238 ( .A1(n6169), .A2(n6168), .ZN(U2818) );
  OAI22_X1 U7239 ( .A1(n6236), .A2(n6303), .B1(n6170), .B2(n6266), .ZN(n6177)
         );
  AOI22_X1 U7240 ( .A1(n6171), .A2(n6261), .B1(n6201), .B2(n6302), .ZN(n6175)
         );
  OAI21_X1 U7241 ( .B1(REIP_REG_8__SCAN_IN), .B2(n6173), .A(n6172), .ZN(n6174)
         );
  OAI211_X1 U7242 ( .C1(n6245), .C2(n6304), .A(n6175), .B(n6174), .ZN(n6176)
         );
  OR3_X1 U7243 ( .A1(n6216), .A2(n6177), .A3(n6176), .ZN(U2819) );
  AOI21_X1 U7244 ( .B1(n6234), .B2(PHYADDRPOINTER_REG_7__SCAN_IN), .A(n6216), 
        .ZN(n6191) );
  AND2_X1 U7245 ( .A1(n6179), .A2(n6178), .ZN(n6181) );
  OR2_X1 U7246 ( .A1(n6181), .A2(n6180), .ZN(n6511) );
  INV_X1 U7247 ( .A(n6511), .ZN(n6182) );
  AOI22_X1 U7248 ( .A1(n6265), .A2(n6182), .B1(n6264), .B2(EBX_REG_7__SCAN_IN), 
        .ZN(n6190) );
  INV_X1 U7249 ( .A(n6184), .ZN(n6183) );
  OAI21_X1 U7250 ( .B1(n6183), .B2(n6240), .A(n6254), .ZN(n6209) );
  NOR3_X1 U7251 ( .A1(n6240), .A2(REIP_REG_6__SCAN_IN), .A3(n6184), .ZN(n6194)
         );
  OAI22_X1 U7252 ( .A1(n6471), .A2(n6267), .B1(n6185), .B2(n6475), .ZN(n6186)
         );
  AOI221_X1 U7253 ( .B1(n6209), .B2(REIP_REG_7__SCAN_IN), .C1(n6194), .C2(
        REIP_REG_7__SCAN_IN), .A(n6186), .ZN(n6189) );
  INV_X1 U7254 ( .A(REIP_REG_7__SCAN_IN), .ZN(n6936) );
  NAND3_X1 U7255 ( .A1(n6256), .A2(n6936), .A3(n6187), .ZN(n6188) );
  NAND4_X1 U7256 ( .A1(n6191), .A2(n6190), .A3(n6189), .A4(n6188), .ZN(U2820)
         );
  AOI22_X1 U7257 ( .A1(EBX_REG_6__SCAN_IN), .A2(n6264), .B1(
        REIP_REG_6__SCAN_IN), .B2(n6209), .ZN(n6198) );
  OAI22_X1 U7258 ( .A1(n6236), .A2(n6307), .B1(n6192), .B2(n6266), .ZN(n6193)
         );
  NOR3_X1 U7259 ( .A1(n6216), .A2(n6194), .A3(n6193), .ZN(n6197) );
  AOI22_X1 U7260 ( .A1(n6195), .A2(n6261), .B1(n6201), .B2(n6306), .ZN(n6196)
         );
  NAND3_X1 U7261 ( .A1(n6198), .A2(n6197), .A3(n6196), .ZN(U2821) );
  INV_X1 U7262 ( .A(EBX_REG_5__SCAN_IN), .ZN(n6310) );
  AND2_X1 U7263 ( .A1(n6199), .A2(n7022), .ZN(n6200) );
  INV_X1 U7264 ( .A(n6482), .ZN(n6207) );
  OAI21_X1 U7265 ( .B1(n6266), .B2(n6202), .A(n3179), .ZN(n6203) );
  AOI21_X1 U7266 ( .B1(n6204), .B2(n6265), .A(n6203), .ZN(n6205) );
  OAI21_X1 U7267 ( .B1(n6267), .B2(n6477), .A(n6205), .ZN(n6206) );
  AOI21_X1 U7268 ( .B1(n6246), .B2(n6207), .A(n6206), .ZN(n6212) );
  AND2_X1 U7269 ( .A1(n6256), .A2(n6208), .ZN(n6210) );
  OAI21_X1 U7270 ( .B1(REIP_REG_5__SCAN_IN), .B2(n6210), .A(n6209), .ZN(n6211)
         );
  OAI211_X1 U7271 ( .C1(n6245), .C2(n6310), .A(n6212), .B(n6211), .ZN(U2822)
         );
  NAND2_X1 U7272 ( .A1(n6256), .A2(n6218), .ZN(n6232) );
  NAND2_X1 U7273 ( .A1(n6254), .A2(n6232), .ZN(n6229) );
  AOI22_X1 U7274 ( .A1(EBX_REG_4__SCAN_IN), .A2(n6264), .B1(
        REIP_REG_4__SCAN_IN), .B2(n6229), .ZN(n6222) );
  INV_X1 U7275 ( .A(n6213), .ZN(n6214) );
  NOR2_X1 U7276 ( .A1(n3422), .A2(n7036), .ZN(n6269) );
  INV_X1 U7277 ( .A(n6269), .ZN(n6258) );
  OAI22_X1 U7278 ( .A1(n6236), .A2(n6312), .B1(n6214), .B2(n6258), .ZN(n6215)
         );
  AOI211_X1 U7279 ( .C1(n6234), .C2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n6216), 
        .B(n6215), .ZN(n6221) );
  AOI22_X1 U7280 ( .A1(n6217), .A2(n6261), .B1(n6361), .B2(n6246), .ZN(n6220)
         );
  OR3_X1 U7281 ( .A1(n6240), .A2(REIP_REG_4__SCAN_IN), .A3(n6218), .ZN(n6219)
         );
  NAND4_X1 U7282 ( .A1(n6222), .A2(n6221), .A3(n6220), .A4(n6219), .ZN(U2823)
         );
  NAND2_X1 U7283 ( .A1(REIP_REG_2__SCAN_IN), .A2(REIP_REG_1__SCAN_IN), .ZN(
        n6233) );
  INV_X1 U7284 ( .A(n6364), .ZN(n6228) );
  AOI22_X1 U7285 ( .A1(n6636), .A2(n6269), .B1(PHYADDRPOINTER_REG_3__SCAN_IN), 
        .B2(n6234), .ZN(n6223) );
  OAI21_X1 U7286 ( .B1(n6236), .B2(n6313), .A(n6223), .ZN(n6224) );
  AOI21_X1 U7287 ( .B1(EBX_REG_3__SCAN_IN), .B2(n6264), .A(n6224), .ZN(n6225)
         );
  OAI21_X1 U7288 ( .B1(n6267), .B2(n6226), .A(n6225), .ZN(n6227) );
  AOI21_X1 U7289 ( .B1(n6228), .B2(n6246), .A(n6227), .ZN(n6231) );
  NAND2_X1 U7290 ( .A1(REIP_REG_3__SCAN_IN), .A2(n6229), .ZN(n6230) );
  OAI211_X1 U7291 ( .C1(n6233), .C2(n6232), .A(n6231), .B(n6230), .ZN(U2824)
         );
  INV_X1 U7292 ( .A(EBX_REG_2__SCAN_IN), .ZN(n6316) );
  INV_X1 U7293 ( .A(n6483), .ZN(n6239) );
  AOI22_X1 U7294 ( .A1(n3210), .A2(n6269), .B1(n6234), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n6235) );
  OAI21_X1 U7295 ( .B1(n6236), .B2(n6315), .A(n6235), .ZN(n6238) );
  NOR2_X1 U7296 ( .A1(n6267), .A2(n6489), .ZN(n6237) );
  AOI211_X1 U7297 ( .C1(n6239), .C2(n6246), .A(n6238), .B(n6237), .ZN(n6244)
         );
  NOR2_X1 U7298 ( .A1(n6240), .A2(n7015), .ZN(n6242) );
  NAND3_X1 U7299 ( .A1(n6254), .A2(REIP_REG_2__SCAN_IN), .A3(
        REIP_REG_1__SCAN_IN), .ZN(n6241) );
  OAI211_X1 U7300 ( .C1(REIP_REG_2__SCAN_IN), .C2(n6242), .A(n6270), .B(n6241), 
        .ZN(n6243) );
  OAI211_X1 U7301 ( .C1(n6245), .C2(n6316), .A(n6244), .B(n6243), .ZN(U2825)
         );
  INV_X1 U7302 ( .A(n6246), .ZN(n6273) );
  OAI21_X1 U7303 ( .B1(n6249), .B2(n6248), .A(n6247), .ZN(n6501) );
  OR2_X1 U7304 ( .A1(n6251), .A2(n6250), .ZN(n6253) );
  AND2_X1 U7305 ( .A1(n6253), .A2(n6252), .ZN(n6319) );
  INV_X1 U7306 ( .A(n6319), .ZN(n6524) );
  INV_X1 U7307 ( .A(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n6497) );
  OAI22_X1 U7308 ( .A1(n6497), .A2(n6266), .B1(n6254), .B2(n7015), .ZN(n6255)
         );
  AOI21_X1 U7309 ( .B1(n6256), .B2(n7015), .A(n6255), .ZN(n6257) );
  OAI21_X1 U7310 ( .B1(n6259), .B2(n6258), .A(n6257), .ZN(n6260) );
  AOI21_X1 U7311 ( .B1(n6265), .B2(n6524), .A(n6260), .ZN(n6263) );
  AOI22_X1 U7312 ( .A1(EBX_REG_1__SCAN_IN), .A2(n6264), .B1(n6261), .B2(n6497), 
        .ZN(n6262) );
  OAI211_X1 U7313 ( .C1(n6273), .C2(n6501), .A(n6263), .B(n6262), .ZN(U2826)
         );
  INV_X1 U7314 ( .A(n6326), .ZN(n6369) );
  AOI22_X1 U7315 ( .A1(n6265), .A2(n6322), .B1(n6264), .B2(EBX_REG_0__SCAN_IN), 
        .ZN(n6272) );
  NAND2_X1 U7316 ( .A1(n6267), .A2(n6266), .ZN(n6268) );
  AOI222_X1 U7317 ( .A1(REIP_REG_0__SCAN_IN), .A2(n6270), .B1(n6681), .B2(
        n6269), .C1(n6268), .C2(PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n6271) );
  OAI211_X1 U7318 ( .C1(n6273), .C2(n6369), .A(n6272), .B(n6271), .ZN(U2827)
         );
  INV_X1 U7319 ( .A(n6274), .ZN(n6275) );
  AOI22_X1 U7320 ( .A1(n6275), .A2(n6323), .B1(EBX_REG_31__SCAN_IN), .B2(n6324), .ZN(n6276) );
  INV_X1 U7321 ( .A(n6276), .ZN(U2828) );
  INV_X1 U7322 ( .A(n6328), .ZN(n6279) );
  AOI22_X1 U7323 ( .A1(EBX_REG_18__SCAN_IN), .A2(n6324), .B1(n6277), .B2(n6323), .ZN(n6278) );
  OAI21_X1 U7324 ( .B1(n6279), .B2(n6321), .A(n6278), .ZN(U2841) );
  OAI222_X1 U7325 ( .A1(n6282), .A2(n6321), .B1(n6317), .B2(n6281), .C1(n6320), 
        .C2(n6280), .ZN(U2842) );
  OAI222_X1 U7326 ( .A1(n6285), .A2(n6321), .B1(n6317), .B2(n6284), .C1(n6320), 
        .C2(n6283), .ZN(U2843) );
  INV_X1 U7327 ( .A(EBX_REG_15__SCAN_IN), .ZN(n6287) );
  OAI222_X1 U7328 ( .A1(n6340), .A2(n6321), .B1(n6317), .B2(n6287), .C1(n6320), 
        .C2(n6286), .ZN(U2844) );
  INV_X1 U7329 ( .A(n6288), .ZN(n6342) );
  OAI222_X1 U7330 ( .A1(n6342), .A2(n6321), .B1(n6317), .B2(n6290), .C1(n6320), 
        .C2(n6289), .ZN(U2845) );
  AOI222_X1 U7331 ( .A1(n6292), .A2(n6325), .B1(n6324), .B2(
        EBX_REG_13__SCAN_IN), .C1(n6323), .C2(n6291), .ZN(n6293) );
  INV_X1 U7332 ( .A(n6293), .ZN(U2846) );
  AOI22_X1 U7333 ( .A1(n6325), .A2(n6345), .B1(n6323), .B2(n6294), .ZN(n6295)
         );
  OAI21_X1 U7334 ( .B1(n6296), .B2(n6317), .A(n6295), .ZN(U2847) );
  AOI22_X1 U7335 ( .A1(EBX_REG_11__SCAN_IN), .A2(n6324), .B1(n6323), .B2(n3222), .ZN(n6297) );
  OAI21_X1 U7336 ( .B1(n6321), .B2(n6349), .A(n6297), .ZN(U2848) );
  OAI222_X1 U7337 ( .A1(n6351), .A2(n6321), .B1(n6317), .B2(n6299), .C1(n6320), 
        .C2(n6298), .ZN(U2849) );
  INV_X1 U7338 ( .A(EBX_REG_9__SCAN_IN), .ZN(n6301) );
  AOI22_X1 U7339 ( .A1(n6325), .A2(n6352), .B1(n6323), .B2(n6504), .ZN(n6300)
         );
  OAI21_X1 U7340 ( .B1(n6301), .B2(n6317), .A(n6300), .ZN(U2850) );
  INV_X1 U7341 ( .A(n6302), .ZN(n6355) );
  OAI222_X1 U7342 ( .A1(n6355), .A2(n6321), .B1(n6317), .B2(n6304), .C1(n6320), 
        .C2(n6303), .ZN(U2851) );
  INV_X1 U7343 ( .A(EBX_REG_7__SCAN_IN), .ZN(n6305) );
  OAI222_X1 U7344 ( .A1(n6475), .A2(n6321), .B1(n6317), .B2(n6305), .C1(n6320), 
        .C2(n6511), .ZN(U2852) );
  INV_X1 U7345 ( .A(n6306), .ZN(n6357) );
  OAI222_X1 U7346 ( .A1(n6357), .A2(n6321), .B1(n6317), .B2(n6308), .C1(n6320), 
        .C2(n6307), .ZN(U2853) );
  OAI222_X1 U7347 ( .A1(n6482), .A2(n6321), .B1(n6317), .B2(n6310), .C1(n6320), 
        .C2(n6309), .ZN(U2854) );
  AOI22_X1 U7348 ( .A1(EBX_REG_4__SCAN_IN), .A2(n6324), .B1(n6325), .B2(n6361), 
        .ZN(n6311) );
  OAI21_X1 U7349 ( .B1(n6320), .B2(n6312), .A(n6311), .ZN(U2855) );
  INV_X1 U7350 ( .A(EBX_REG_3__SCAN_IN), .ZN(n6314) );
  OAI222_X1 U7351 ( .A1(n6364), .A2(n6321), .B1(n6317), .B2(n6314), .C1(n6320), 
        .C2(n6313), .ZN(U2856) );
  OAI222_X1 U7352 ( .A1(n6483), .A2(n6321), .B1(n6317), .B2(n6316), .C1(n6320), 
        .C2(n6315), .ZN(U2857) );
  INV_X1 U7353 ( .A(EBX_REG_1__SCAN_IN), .ZN(n6318) );
  OAI222_X1 U7354 ( .A1(n6501), .A2(n6321), .B1(n6320), .B2(n6319), .C1(n6318), 
        .C2(n6317), .ZN(U2858) );
  AOI222_X1 U7355 ( .A1(n6326), .A2(n6325), .B1(n6324), .B2(EBX_REG_0__SCAN_IN), .C1(n6323), .C2(n6322), .ZN(n6327) );
  INV_X1 U7356 ( .A(n6327), .ZN(U2859) );
  AOI22_X1 U7357 ( .A1(n6335), .A2(DATAI_18_), .B1(n6328), .B2(n6360), .ZN(
        n6330) );
  AOI22_X1 U7358 ( .A1(EAX_REG_18__SCAN_IN), .A2(n6358), .B1(DATAI_2_), .B2(
        n6336), .ZN(n6329) );
  NAND2_X1 U7359 ( .A1(n6330), .A2(n6329), .ZN(U2873) );
  AOI22_X1 U7360 ( .A1(n6335), .A2(DATAI_17_), .B1(n6360), .B2(n6331), .ZN(
        n6333) );
  AOI22_X1 U7361 ( .A1(EAX_REG_17__SCAN_IN), .A2(n6358), .B1(n6336), .B2(
        DATAI_1_), .ZN(n6332) );
  NAND2_X1 U7362 ( .A1(n6333), .A2(n6332), .ZN(U2874) );
  AOI22_X1 U7363 ( .A1(DATAI_16_), .A2(n6335), .B1(n6360), .B2(n6334), .ZN(
        n6338) );
  AOI22_X1 U7364 ( .A1(EAX_REG_16__SCAN_IN), .A2(n6358), .B1(n6336), .B2(
        DATAI_0_), .ZN(n6337) );
  NAND2_X1 U7365 ( .A1(n6338), .A2(n6337), .ZN(U2875) );
  INV_X1 U7366 ( .A(EAX_REG_15__SCAN_IN), .ZN(n6400) );
  OAI222_X1 U7367 ( .A1(n6340), .A2(n6368), .B1(n6339), .B2(n6366), .C1(n6400), 
        .C2(n6365), .ZN(U2876) );
  INV_X1 U7368 ( .A(DATAI_14_), .ZN(n6341) );
  OAI222_X1 U7369 ( .A1(n6342), .A2(n6368), .B1(n6341), .B2(n6366), .C1(n6402), 
        .C2(n6365), .ZN(U2877) );
  INV_X1 U7370 ( .A(DATAI_13_), .ZN(n6343) );
  OAI222_X1 U7371 ( .A1(n6344), .A2(n6368), .B1(n6343), .B2(n6366), .C1(n6404), 
        .C2(n6365), .ZN(U2878) );
  INV_X1 U7372 ( .A(n6345), .ZN(n6347) );
  INV_X1 U7373 ( .A(n6366), .ZN(n6359) );
  AOI22_X1 U7374 ( .A1(EAX_REG_12__SCAN_IN), .A2(n6358), .B1(DATAI_12_), .B2(
        n6359), .ZN(n6346) );
  OAI21_X1 U7375 ( .B1(n6368), .B2(n6347), .A(n6346), .ZN(U2879) );
  AOI22_X1 U7376 ( .A1(EAX_REG_11__SCAN_IN), .A2(n6358), .B1(DATAI_11_), .B2(
        n6359), .ZN(n6348) );
  OAI21_X1 U7377 ( .B1(n6368), .B2(n6349), .A(n6348), .ZN(U2880) );
  INV_X1 U7378 ( .A(DATAI_10_), .ZN(n6350) );
  INV_X1 U7379 ( .A(EAX_REG_10__SCAN_IN), .ZN(n6410) );
  OAI222_X1 U7380 ( .A1(n6351), .A2(n6368), .B1(n6350), .B2(n6366), .C1(n6410), 
        .C2(n6365), .ZN(U2881) );
  AOI222_X1 U7381 ( .A1(n6352), .A2(n6360), .B1(DATAI_9_), .B2(n6359), .C1(
        EAX_REG_9__SCAN_IN), .C2(n6358), .ZN(n6353) );
  INV_X1 U7382 ( .A(n6353), .ZN(U2882) );
  AOI22_X1 U7383 ( .A1(EAX_REG_8__SCAN_IN), .A2(n6358), .B1(DATAI_8_), .B2(
        n6359), .ZN(n6354) );
  OAI21_X1 U7384 ( .B1(n6368), .B2(n6355), .A(n6354), .ZN(U2883) );
  INV_X1 U7385 ( .A(DATAI_6_), .ZN(n6356) );
  OAI222_X1 U7386 ( .A1(n6357), .A2(n6368), .B1(n6356), .B2(n6366), .C1(n6421), 
        .C2(n6365), .ZN(U2885) );
  AOI222_X1 U7387 ( .A1(n6361), .A2(n6360), .B1(DATAI_4_), .B2(n6359), .C1(
        EAX_REG_4__SCAN_IN), .C2(n6358), .ZN(n6362) );
  INV_X1 U7388 ( .A(n6362), .ZN(U2887) );
  OAI222_X1 U7389 ( .A1(n6364), .A2(n6368), .B1(n6363), .B2(n6366), .C1(n6427), 
        .C2(n6365), .ZN(U2888) );
  OAI222_X1 U7390 ( .A1(n6501), .A2(n6368), .B1(n4822), .B2(n6366), .C1(n6432), 
        .C2(n6365), .ZN(U2890) );
  INV_X1 U7391 ( .A(DATAI_0_), .ZN(n6367) );
  OAI222_X1 U7392 ( .A1(n6369), .A2(n6368), .B1(n6367), .B2(n6366), .C1(n6437), 
        .C2(n6365), .ZN(U2891) );
  NAND2_X1 U7393 ( .A1(n6414), .A2(n3444), .ZN(n6397) );
  AOI22_X1 U7394 ( .A1(n6419), .A2(UWORD_REG_14__SCAN_IN), .B1(n6411), .B2(
        DATAO_REG_30__SCAN_IN), .ZN(n6370) );
  OAI21_X1 U7395 ( .B1(n6371), .B2(n6397), .A(n6370), .ZN(U2893) );
  AOI22_X1 U7396 ( .A1(n6419), .A2(UWORD_REG_13__SCAN_IN), .B1(n6411), .B2(
        DATAO_REG_29__SCAN_IN), .ZN(n6372) );
  OAI21_X1 U7397 ( .B1(n6373), .B2(n6397), .A(n6372), .ZN(U2894) );
  INV_X1 U7398 ( .A(n6397), .ZN(n6394) );
  AOI22_X1 U7399 ( .A1(EAX_REG_28__SCAN_IN), .A2(n6394), .B1(n6419), .B2(
        UWORD_REG_12__SCAN_IN), .ZN(n6374) );
  OAI21_X1 U7400 ( .B1(n6375), .B2(n6434), .A(n6374), .ZN(U2895) );
  AOI22_X1 U7401 ( .A1(n6419), .A2(UWORD_REG_11__SCAN_IN), .B1(n6411), .B2(
        DATAO_REG_27__SCAN_IN), .ZN(n6376) );
  OAI21_X1 U7402 ( .B1(n6377), .B2(n6397), .A(n6376), .ZN(U2896) );
  AOI22_X1 U7403 ( .A1(EAX_REG_26__SCAN_IN), .A2(n6394), .B1(n6411), .B2(
        DATAO_REG_26__SCAN_IN), .ZN(n6378) );
  OAI21_X1 U7404 ( .B1(n6449), .B2(n6431), .A(n6378), .ZN(U2897) );
  AOI22_X1 U7405 ( .A1(n6419), .A2(UWORD_REG_9__SCAN_IN), .B1(n6411), .B2(
        DATAO_REG_25__SCAN_IN), .ZN(n6379) );
  OAI21_X1 U7406 ( .B1(n6380), .B2(n6397), .A(n6379), .ZN(U2898) );
  AOI22_X1 U7407 ( .A1(EAX_REG_24__SCAN_IN), .A2(n6394), .B1(n6419), .B2(
        UWORD_REG_8__SCAN_IN), .ZN(n6381) );
  OAI21_X1 U7408 ( .B1(n6382), .B2(n6434), .A(n6381), .ZN(U2899) );
  AOI22_X1 U7409 ( .A1(n6419), .A2(UWORD_REG_7__SCAN_IN), .B1(n6411), .B2(
        DATAO_REG_23__SCAN_IN), .ZN(n6383) );
  OAI21_X1 U7410 ( .B1(n6384), .B2(n6397), .A(n6383), .ZN(U2900) );
  AOI22_X1 U7411 ( .A1(DATAO_REG_22__SCAN_IN), .A2(n6411), .B1(n6419), .B2(
        UWORD_REG_6__SCAN_IN), .ZN(n6385) );
  OAI21_X1 U7412 ( .B1(n6386), .B2(n6397), .A(n6385), .ZN(U2901) );
  AOI22_X1 U7413 ( .A1(n6419), .A2(UWORD_REG_5__SCAN_IN), .B1(n6411), .B2(
        DATAO_REG_21__SCAN_IN), .ZN(n6387) );
  OAI21_X1 U7414 ( .B1(n6388), .B2(n6397), .A(n6387), .ZN(U2902) );
  AOI22_X1 U7415 ( .A1(EAX_REG_20__SCAN_IN), .A2(n6394), .B1(n6411), .B2(
        DATAO_REG_20__SCAN_IN), .ZN(n6389) );
  OAI21_X1 U7416 ( .B1(n6445), .B2(n6431), .A(n6389), .ZN(U2903) );
  AOI22_X1 U7417 ( .A1(n6419), .A2(UWORD_REG_3__SCAN_IN), .B1(n6411), .B2(
        DATAO_REG_19__SCAN_IN), .ZN(n6390) );
  OAI21_X1 U7418 ( .B1(n6391), .B2(n6397), .A(n6390), .ZN(U2904) );
  INV_X1 U7419 ( .A(EAX_REG_18__SCAN_IN), .ZN(n6393) );
  OAI222_X1 U7420 ( .A1(n6431), .A2(n6442), .B1(n6397), .B2(n6393), .C1(n6392), 
        .C2(n6434), .ZN(U2905) );
  AOI22_X1 U7421 ( .A1(EAX_REG_17__SCAN_IN), .A2(n6394), .B1(n6411), .B2(
        DATAO_REG_17__SCAN_IN), .ZN(n6395) );
  OAI21_X1 U7422 ( .B1(n6440), .B2(n6431), .A(n6395), .ZN(U2906) );
  AOI22_X1 U7423 ( .A1(n6419), .A2(UWORD_REG_0__SCAN_IN), .B1(n6411), .B2(
        DATAO_REG_16__SCAN_IN), .ZN(n6396) );
  OAI21_X1 U7424 ( .B1(n6398), .B2(n6397), .A(n6396), .ZN(U2907) );
  AOI22_X1 U7425 ( .A1(LWORD_REG_15__SCAN_IN), .A2(n6419), .B1(
        DATAO_REG_15__SCAN_IN), .B2(n6411), .ZN(n6399) );
  OAI21_X1 U7426 ( .B1(n6400), .B2(n6436), .A(n6399), .ZN(U2908) );
  AOI22_X1 U7427 ( .A1(n6419), .A2(LWORD_REG_14__SCAN_IN), .B1(n6411), .B2(
        DATAO_REG_14__SCAN_IN), .ZN(n6401) );
  OAI21_X1 U7428 ( .B1(n6402), .B2(n6436), .A(n6401), .ZN(U2909) );
  AOI22_X1 U7429 ( .A1(n6419), .A2(LWORD_REG_13__SCAN_IN), .B1(n6411), .B2(
        DATAO_REG_13__SCAN_IN), .ZN(n6403) );
  OAI21_X1 U7430 ( .B1(n6404), .B2(n6436), .A(n6403), .ZN(U2910) );
  INV_X1 U7431 ( .A(EAX_REG_12__SCAN_IN), .ZN(n6406) );
  OAI222_X1 U7432 ( .A1(n6431), .A2(n6407), .B1(n6436), .B2(n6406), .C1(n6405), 
        .C2(n6434), .ZN(U2911) );
  AOI22_X1 U7433 ( .A1(EAX_REG_11__SCAN_IN), .A2(n6414), .B1(n6411), .B2(
        DATAO_REG_11__SCAN_IN), .ZN(n6408) );
  OAI21_X1 U7434 ( .B1(n6462), .B2(n6431), .A(n6408), .ZN(U2912) );
  AOI22_X1 U7435 ( .A1(LWORD_REG_10__SCAN_IN), .A2(n6419), .B1(n6411), .B2(
        DATAO_REG_10__SCAN_IN), .ZN(n6409) );
  OAI21_X1 U7436 ( .B1(n6410), .B2(n6436), .A(n6409), .ZN(U2913) );
  AOI22_X1 U7437 ( .A1(n6419), .A2(LWORD_REG_9__SCAN_IN), .B1(n6411), .B2(
        DATAO_REG_9__SCAN_IN), .ZN(n6412) );
  OAI21_X1 U7438 ( .B1(n6413), .B2(n6436), .A(n6412), .ZN(U2914) );
  AOI22_X1 U7439 ( .A1(EAX_REG_8__SCAN_IN), .A2(n6414), .B1(n6419), .B2(
        LWORD_REG_8__SCAN_IN), .ZN(n6415) );
  OAI21_X1 U7440 ( .B1(n6416), .B2(n6434), .A(n6415), .ZN(U2915) );
  AOI22_X1 U7441 ( .A1(n6419), .A2(LWORD_REG_7__SCAN_IN), .B1(n6411), .B2(
        DATAO_REG_7__SCAN_IN), .ZN(n6417) );
  OAI21_X1 U7442 ( .B1(n6418), .B2(n6436), .A(n6417), .ZN(U2916) );
  AOI22_X1 U7443 ( .A1(n6419), .A2(LWORD_REG_6__SCAN_IN), .B1(n6411), .B2(
        DATAO_REG_6__SCAN_IN), .ZN(n6420) );
  OAI21_X1 U7444 ( .B1(n6421), .B2(n6436), .A(n6420), .ZN(U2917) );
  AOI22_X1 U7445 ( .A1(n6419), .A2(LWORD_REG_5__SCAN_IN), .B1(n6411), .B2(
        DATAO_REG_5__SCAN_IN), .ZN(n6422) );
  OAI21_X1 U7446 ( .B1(n6423), .B2(n6436), .A(n6422), .ZN(U2918) );
  AOI22_X1 U7447 ( .A1(n6419), .A2(LWORD_REG_4__SCAN_IN), .B1(n6411), .B2(
        DATAO_REG_4__SCAN_IN), .ZN(n6424) );
  OAI21_X1 U7448 ( .B1(n6425), .B2(n6436), .A(n6424), .ZN(U2919) );
  AOI22_X1 U7449 ( .A1(n6419), .A2(LWORD_REG_3__SCAN_IN), .B1(n6411), .B2(
        DATAO_REG_3__SCAN_IN), .ZN(n6426) );
  OAI21_X1 U7450 ( .B1(n6427), .B2(n6436), .A(n6426), .ZN(U2920) );
  INV_X1 U7451 ( .A(LWORD_REG_2__SCAN_IN), .ZN(n6454) );
  OAI222_X1 U7452 ( .A1(n6434), .A2(n6429), .B1(n6436), .B2(n6428), .C1(n6431), 
        .C2(n6454), .ZN(U2921) );
  INV_X1 U7453 ( .A(DATAO_REG_1__SCAN_IN), .ZN(n6433) );
  OAI222_X1 U7454 ( .A1(n6434), .A2(n6433), .B1(n6436), .B2(n6432), .C1(n6431), 
        .C2(n6430), .ZN(U2922) );
  AOI22_X1 U7455 ( .A1(DATAO_REG_0__SCAN_IN), .A2(n6411), .B1(n6419), .B2(
        LWORD_REG_0__SCAN_IN), .ZN(n6435) );
  OAI21_X1 U7456 ( .B1(n6437), .B2(n6436), .A(n6435), .ZN(U2923) );
  AOI21_X1 U7457 ( .B1(n6465), .B2(EAX_REG_17__SCAN_IN), .A(n6438), .ZN(n6439)
         );
  OAI21_X1 U7458 ( .B1(n6463), .B2(n6440), .A(n6439), .ZN(U2925) );
  NOR2_X1 U7459 ( .A1(n6447), .A2(n5276), .ZN(n6452) );
  AOI21_X1 U7460 ( .B1(n6465), .B2(EAX_REG_18__SCAN_IN), .A(n6452), .ZN(n6441)
         );
  OAI21_X1 U7461 ( .B1(n6463), .B2(n6442), .A(n6441), .ZN(U2926) );
  AOI21_X1 U7462 ( .B1(n6465), .B2(EAX_REG_20__SCAN_IN), .A(n6443), .ZN(n6444)
         );
  OAI21_X1 U7463 ( .B1(n6463), .B2(n6445), .A(n6444), .ZN(U2928) );
  AOI22_X1 U7464 ( .A1(n6465), .A2(EAX_REG_24__SCAN_IN), .B1(n6464), .B2(
        UWORD_REG_8__SCAN_IN), .ZN(n6446) );
  NAND2_X1 U7465 ( .A1(n6450), .A2(DATAI_8_), .ZN(n6455) );
  NAND2_X1 U7466 ( .A1(n6446), .A2(n6455), .ZN(U2932) );
  NOR2_X1 U7467 ( .A1(n6447), .A2(n6350), .ZN(n6457) );
  AOI21_X1 U7468 ( .B1(n6465), .B2(EAX_REG_26__SCAN_IN), .A(n6457), .ZN(n6448)
         );
  OAI21_X1 U7469 ( .B1(n6463), .B2(n6449), .A(n6448), .ZN(U2934) );
  AOI22_X1 U7470 ( .A1(n6465), .A2(EAX_REG_28__SCAN_IN), .B1(n6464), .B2(
        UWORD_REG_12__SCAN_IN), .ZN(n6451) );
  NAND2_X1 U7471 ( .A1(n6450), .A2(DATAI_12_), .ZN(n6466) );
  NAND2_X1 U7472 ( .A1(n6451), .A2(n6466), .ZN(U2936) );
  AOI21_X1 U7473 ( .B1(n6465), .B2(EAX_REG_2__SCAN_IN), .A(n6452), .ZN(n6453)
         );
  OAI21_X1 U7474 ( .B1(n6463), .B2(n6454), .A(n6453), .ZN(U2941) );
  AOI22_X1 U7475 ( .A1(n6465), .A2(EAX_REG_8__SCAN_IN), .B1(n6464), .B2(
        LWORD_REG_8__SCAN_IN), .ZN(n6456) );
  NAND2_X1 U7476 ( .A1(n6456), .A2(n6455), .ZN(U2947) );
  AOI21_X1 U7477 ( .B1(n6465), .B2(EAX_REG_10__SCAN_IN), .A(n6457), .ZN(n6458)
         );
  OAI21_X1 U7478 ( .B1(n6463), .B2(n6459), .A(n6458), .ZN(U2949) );
  AOI21_X1 U7479 ( .B1(n6465), .B2(EAX_REG_11__SCAN_IN), .A(n6460), .ZN(n6461)
         );
  OAI21_X1 U7480 ( .B1(n6463), .B2(n6462), .A(n6461), .ZN(U2950) );
  AOI22_X1 U7481 ( .A1(n6465), .A2(EAX_REG_12__SCAN_IN), .B1(n6464), .B2(
        LWORD_REG_12__SCAN_IN), .ZN(n6467) );
  NAND2_X1 U7482 ( .A1(n6467), .A2(n6466), .ZN(U2951) );
  NOR2_X1 U7483 ( .A1(n3179), .A2(n6936), .ZN(n6514) );
  XOR2_X1 U7484 ( .A(n6468), .B(n6470), .Z(n6519) );
  INV_X1 U7485 ( .A(n6519), .ZN(n6472) );
  OAI22_X1 U7486 ( .A1(n6472), .A2(n6484), .B1(n6471), .B2(n6490), .ZN(n6473)
         );
  AOI211_X1 U7487 ( .C1(n6491), .C2(PHYADDRPOINTER_REG_7__SCAN_IN), .A(n6514), 
        .B(n6473), .ZN(n6474) );
  OAI21_X1 U7488 ( .B1(n6476), .B2(n6475), .A(n6474), .ZN(U2979) );
  OAI22_X1 U7489 ( .A1(n6478), .A2(n6484), .B1(n6477), .B2(n6490), .ZN(n6479)
         );
  AOI211_X1 U7490 ( .C1(n6491), .C2(PHYADDRPOINTER_REG_5__SCAN_IN), .A(n6480), 
        .B(n6479), .ZN(n6481) );
  OAI21_X1 U7491 ( .B1(n6476), .B2(n6482), .A(n6481), .ZN(U2981) );
  AOI22_X1 U7492 ( .A1(PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n6491), .B1(n6523), 
        .B2(REIP_REG_2__SCAN_IN), .ZN(n6488) );
  OAI22_X1 U7493 ( .A1(n6485), .A2(n6484), .B1(n6483), .B2(n6476), .ZN(n6486)
         );
  INV_X1 U7494 ( .A(n6486), .ZN(n6487) );
  OAI211_X1 U7495 ( .C1(n6490), .C2(n6489), .A(n6488), .B(n6487), .ZN(U2984)
         );
  AOI22_X1 U7496 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n6491), .B1(n6523), 
        .B2(REIP_REG_1__SCAN_IN), .ZN(n6500) );
  OR2_X1 U7497 ( .A1(n6493), .A2(n6492), .ZN(n6494) );
  AND2_X1 U7498 ( .A1(n6495), .A2(n6494), .ZN(n6527) );
  AOI22_X1 U7499 ( .A1(n6498), .A2(n6497), .B1(n6527), .B2(n6496), .ZN(n6499)
         );
  OAI211_X1 U7500 ( .C1(n6476), .C2(n6501), .A(n6500), .B(n6499), .ZN(U2985)
         );
  INV_X1 U7501 ( .A(n6502), .ZN(n6503) );
  AOI21_X1 U7502 ( .B1(n6525), .B2(n6504), .A(n6503), .ZN(n6509) );
  INV_X1 U7503 ( .A(n6505), .ZN(n6507) );
  AOI22_X1 U7504 ( .A1(n6507), .A2(n6528), .B1(INSTADDRPOINTER_REG_9__SCAN_IN), 
        .B2(n6506), .ZN(n6508) );
  OAI211_X1 U7505 ( .C1(INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n6510), .A(n6509), 
        .B(n6508), .ZN(U3009) );
  NOR2_X1 U7506 ( .A1(n6512), .A2(n6511), .ZN(n6518) );
  INV_X1 U7507 ( .A(n6513), .ZN(n6516) );
  INV_X1 U7508 ( .A(n6514), .ZN(n6515) );
  OAI21_X1 U7509 ( .B1(INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n6516), .A(n6515), 
        .ZN(n6517) );
  AOI211_X1 U7510 ( .C1(n6519), .C2(n6528), .A(n6518), .B(n6517), .ZN(n6520)
         );
  OAI21_X1 U7511 ( .B1(n6522), .B2(n6521), .A(n6520), .ZN(U3011) );
  AOI22_X1 U7512 ( .A1(n6525), .A2(n6524), .B1(n6523), .B2(REIP_REG_1__SCAN_IN), .ZN(n6534) );
  AOI22_X1 U7513 ( .A1(n6528), .A2(n6527), .B1(INSTADDRPOINTER_REG_1__SCAN_IN), 
        .B2(n6526), .ZN(n6533) );
  NAND3_X1 U7514 ( .A1(n6531), .A2(n6530), .A3(n6529), .ZN(n6532) );
  NAND3_X1 U7515 ( .A1(n6534), .A2(n6533), .A3(n6532), .ZN(U3017) );
  NOR2_X1 U7516 ( .A1(n6536), .A2(n6535), .ZN(U3019) );
  NAND3_X1 U7517 ( .A1(n6538), .A2(n6678), .A3(n6537), .ZN(n6539) );
  NAND2_X1 U7518 ( .A1(n6539), .A2(n6643), .ZN(n6546) );
  NOR2_X1 U7519 ( .A1(n6677), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6561)
         );
  AOI21_X1 U7520 ( .B1(n6540), .B2(n6681), .A(n6561), .ZN(n6542) );
  OAI22_X1 U7521 ( .A1(n6546), .A2(n6542), .B1(n6543), .B2(n6773), .ZN(n6541)
         );
  AOI22_X1 U7522 ( .A1(n6562), .A2(n6836), .B1(n6833), .B2(n6561), .ZN(n6548)
         );
  INV_X1 U7523 ( .A(n6542), .ZN(n6545) );
  NAND2_X1 U7524 ( .A1(n6543), .A2(n6776), .ZN(n6544) );
  OAI211_X1 U7525 ( .C1(n6546), .C2(n6545), .A(n6780), .B(n6544), .ZN(n6564)
         );
  AOI22_X1 U7526 ( .A1(INSTQUEUE_REG_3__0__SCAN_IN), .A2(n6564), .B1(n6839), 
        .B2(n6563), .ZN(n6547) );
  OAI211_X1 U7527 ( .C1(n6567), .C2(n6783), .A(n6548), .B(n6547), .ZN(U3044)
         );
  AOI22_X1 U7528 ( .A1(n6562), .A2(n6785), .B1(n6784), .B2(n6561), .ZN(n6550)
         );
  AOI22_X1 U7529 ( .A1(INSTQUEUE_REG_3__1__SCAN_IN), .A2(n6564), .B1(n6786), 
        .B2(n6563), .ZN(n6549) );
  OAI211_X1 U7530 ( .C1(n6567), .C2(n6789), .A(n6550), .B(n6549), .ZN(U3045)
         );
  AOI22_X1 U7531 ( .A1(n6562), .A2(n6792), .B1(n6790), .B2(n6561), .ZN(n6552)
         );
  AOI22_X1 U7532 ( .A1(INSTQUEUE_REG_3__2__SCAN_IN), .A2(n6564), .B1(n6791), 
        .B2(n6563), .ZN(n6551) );
  OAI211_X1 U7533 ( .C1(n6567), .C2(n6795), .A(n6552), .B(n6551), .ZN(U3046)
         );
  AOI22_X1 U7534 ( .A1(n6562), .A2(n6797), .B1(n6796), .B2(n6561), .ZN(n6554)
         );
  AOI22_X1 U7535 ( .A1(INSTQUEUE_REG_3__3__SCAN_IN), .A2(n6564), .B1(n6798), 
        .B2(n6563), .ZN(n6553) );
  OAI211_X1 U7536 ( .C1(n6567), .C2(n6801), .A(n6554), .B(n6553), .ZN(U3047)
         );
  AOI22_X1 U7537 ( .A1(n6562), .A2(n6803), .B1(n6802), .B2(n6561), .ZN(n6556)
         );
  AOI22_X1 U7538 ( .A1(INSTQUEUE_REG_3__4__SCAN_IN), .A2(n6564), .B1(n6804), 
        .B2(n6563), .ZN(n6555) );
  OAI211_X1 U7539 ( .C1(n6567), .C2(n6807), .A(n6556), .B(n6555), .ZN(U3048)
         );
  AOI22_X1 U7540 ( .A1(n6562), .A2(n6809), .B1(n6808), .B2(n6561), .ZN(n6558)
         );
  AOI22_X1 U7541 ( .A1(INSTQUEUE_REG_3__5__SCAN_IN), .A2(n6564), .B1(n6810), 
        .B2(n6563), .ZN(n6557) );
  OAI211_X1 U7542 ( .C1(n6567), .C2(n6813), .A(n6558), .B(n6557), .ZN(U3049)
         );
  AOI22_X1 U7543 ( .A1(n6562), .A2(n6815), .B1(n6814), .B2(n6561), .ZN(n6560)
         );
  AOI22_X1 U7544 ( .A1(INSTQUEUE_REG_3__6__SCAN_IN), .A2(n6564), .B1(n6816), 
        .B2(n6563), .ZN(n6559) );
  OAI211_X1 U7545 ( .C1(n6567), .C2(n6819), .A(n6560), .B(n6559), .ZN(U3050)
         );
  AOI22_X1 U7546 ( .A1(n6562), .A2(n6825), .B1(n6823), .B2(n6561), .ZN(n6566)
         );
  AOI22_X1 U7547 ( .A1(INSTQUEUE_REG_3__7__SCAN_IN), .A2(n6564), .B1(n6820), 
        .B2(n6563), .ZN(n6565) );
  OAI211_X1 U7548 ( .C1(n6567), .C2(n6829), .A(n6566), .B(n6565), .ZN(U3051)
         );
  INV_X1 U7549 ( .A(n6568), .ZN(n6569) );
  NAND2_X1 U7550 ( .A1(n6615), .A2(n6569), .ZN(n6604) );
  NAND3_X1 U7551 ( .A1(n6731), .A2(n6643), .A3(n6607), .ZN(n6570) );
  OAI21_X1 U7552 ( .B1(n6729), .B2(n6571), .A(n6570), .ZN(n6599) );
  NAND2_X1 U7553 ( .A1(n6769), .A2(n6614), .ZN(n6576) );
  INV_X1 U7554 ( .A(n6576), .ZN(n6598) );
  AOI22_X1 U7555 ( .A1(n6832), .A2(n6599), .B1(n6833), .B2(n6598), .ZN(n6580)
         );
  NOR3_X1 U7556 ( .A1(n6600), .A2(n6630), .A3(n6776), .ZN(n6574) );
  INV_X1 U7557 ( .A(n6607), .ZN(n6572) );
  OAI22_X1 U7558 ( .A1(n6574), .A2(n6723), .B1(n6573), .B2(n6572), .ZN(n6578)
         );
  AOI21_X1 U7559 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n6576), .A(n6575), .ZN(
        n6577) );
  NAND3_X1 U7560 ( .A1(n6578), .A2(n6577), .A3(n6725), .ZN(n6601) );
  AOI22_X1 U7561 ( .A1(n6601), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n6836), 
        .B2(n6600), .ZN(n6579) );
  OAI211_X1 U7562 ( .C1(n6581), .C2(n6604), .A(n6580), .B(n6579), .ZN(U3068)
         );
  AOI22_X1 U7563 ( .A1(n6736), .A2(n6599), .B1(n6784), .B2(n6598), .ZN(n6583)
         );
  AOI22_X1 U7564 ( .A1(n6601), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n6785), 
        .B2(n6600), .ZN(n6582) );
  OAI211_X1 U7565 ( .C1(n6693), .C2(n6604), .A(n6583), .B(n6582), .ZN(U3069)
         );
  AOI22_X1 U7566 ( .A1(n6740), .A2(n6599), .B1(n6790), .B2(n6598), .ZN(n6585)
         );
  AOI22_X1 U7567 ( .A1(n6601), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n6792), 
        .B2(n6600), .ZN(n6584) );
  OAI211_X1 U7568 ( .C1(n6696), .C2(n6604), .A(n6585), .B(n6584), .ZN(U3070)
         );
  AOI22_X1 U7569 ( .A1(n6744), .A2(n6599), .B1(n6796), .B2(n6598), .ZN(n6587)
         );
  AOI22_X1 U7570 ( .A1(n6601), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n6797), 
        .B2(n6600), .ZN(n6586) );
  OAI211_X1 U7571 ( .C1(n6588), .C2(n6604), .A(n6587), .B(n6586), .ZN(U3071)
         );
  AOI22_X1 U7572 ( .A1(n6748), .A2(n6599), .B1(n6802), .B2(n6598), .ZN(n6590)
         );
  AOI22_X1 U7573 ( .A1(n6601), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n6803), 
        .B2(n6600), .ZN(n6589) );
  OAI211_X1 U7574 ( .C1(n6591), .C2(n6604), .A(n6590), .B(n6589), .ZN(U3072)
         );
  AOI22_X1 U7575 ( .A1(n6752), .A2(n6599), .B1(n6808), .B2(n6598), .ZN(n6593)
         );
  AOI22_X1 U7576 ( .A1(n6601), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n6809), 
        .B2(n6600), .ZN(n6592) );
  OAI211_X1 U7577 ( .C1(n6594), .C2(n6604), .A(n6593), .B(n6592), .ZN(U3073)
         );
  AOI22_X1 U7578 ( .A1(n6756), .A2(n6599), .B1(n6814), .B2(n6598), .ZN(n6596)
         );
  AOI22_X1 U7579 ( .A1(n6601), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n6815), 
        .B2(n6600), .ZN(n6595) );
  OAI211_X1 U7580 ( .C1(n6597), .C2(n6604), .A(n6596), .B(n6595), .ZN(U3074)
         );
  AOI22_X1 U7581 ( .A1(n6762), .A2(n6599), .B1(n6823), .B2(n6598), .ZN(n6603)
         );
  AOI22_X1 U7582 ( .A1(n6601), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n6825), 
        .B2(n6600), .ZN(n6602) );
  OAI211_X1 U7583 ( .C1(n6717), .C2(n6604), .A(n6603), .B(n6602), .ZN(U3075)
         );
  AND2_X1 U7584 ( .A1(n6605), .A2(n6643), .ZN(n6612) );
  NAND2_X1 U7585 ( .A1(n6607), .A2(n6606), .ZN(n6609) );
  INV_X1 U7586 ( .A(n6631), .ZN(n6608) );
  NAND2_X1 U7587 ( .A1(n6609), .A2(n6608), .ZN(n6610) );
  AOI22_X1 U7588 ( .A1(n6612), .A2(n6610), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n6614), .ZN(n6635) );
  AOI22_X1 U7589 ( .A1(n6631), .A2(n6833), .B1(n6836), .B2(n6630), .ZN(n6617)
         );
  INV_X1 U7590 ( .A(n6610), .ZN(n6611) );
  NAND2_X1 U7591 ( .A1(n6612), .A2(n6611), .ZN(n6613) );
  OAI211_X1 U7592 ( .C1(n6643), .C2(n6614), .A(n6613), .B(n6780), .ZN(n6632)
         );
  NAND2_X1 U7593 ( .A1(n6615), .A2(n6674), .ZN(n6672) );
  AOI22_X1 U7594 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n6632), .B1(n6839), 
        .B2(n6642), .ZN(n6616) );
  OAI211_X1 U7595 ( .C1(n6635), .C2(n6783), .A(n6617), .B(n6616), .ZN(U3076)
         );
  AOI22_X1 U7596 ( .A1(n6631), .A2(n6784), .B1(n6630), .B2(n6785), .ZN(n6619)
         );
  AOI22_X1 U7597 ( .A1(INSTQUEUE_REG_7__1__SCAN_IN), .A2(n6632), .B1(n6786), 
        .B2(n6642), .ZN(n6618) );
  OAI211_X1 U7598 ( .C1(n6635), .C2(n6789), .A(n6619), .B(n6618), .ZN(U3077)
         );
  AOI22_X1 U7599 ( .A1(n6631), .A2(n6790), .B1(n6630), .B2(n6792), .ZN(n6621)
         );
  AOI22_X1 U7600 ( .A1(INSTQUEUE_REG_7__2__SCAN_IN), .A2(n6632), .B1(n6791), 
        .B2(n6642), .ZN(n6620) );
  OAI211_X1 U7601 ( .C1(n6635), .C2(n6795), .A(n6621), .B(n6620), .ZN(U3078)
         );
  AOI22_X1 U7602 ( .A1(n6631), .A2(n6796), .B1(n6642), .B2(n6798), .ZN(n6623)
         );
  AOI22_X1 U7603 ( .A1(INSTQUEUE_REG_7__3__SCAN_IN), .A2(n6632), .B1(n6797), 
        .B2(n6630), .ZN(n6622) );
  OAI211_X1 U7604 ( .C1(n6635), .C2(n6801), .A(n6623), .B(n6622), .ZN(U3079)
         );
  AOI22_X1 U7605 ( .A1(n6631), .A2(n6802), .B1(n6630), .B2(n6803), .ZN(n6625)
         );
  AOI22_X1 U7606 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n6632), .B1(n6804), 
        .B2(n6642), .ZN(n6624) );
  OAI211_X1 U7607 ( .C1(n6635), .C2(n6807), .A(n6625), .B(n6624), .ZN(U3080)
         );
  AOI22_X1 U7608 ( .A1(n6631), .A2(n6808), .B1(n6630), .B2(n6809), .ZN(n6627)
         );
  AOI22_X1 U7609 ( .A1(INSTQUEUE_REG_7__5__SCAN_IN), .A2(n6632), .B1(n6810), 
        .B2(n6642), .ZN(n6626) );
  OAI211_X1 U7610 ( .C1(n6635), .C2(n6813), .A(n6627), .B(n6626), .ZN(U3081)
         );
  AOI22_X1 U7611 ( .A1(n6631), .A2(n6814), .B1(n6642), .B2(n6816), .ZN(n6629)
         );
  AOI22_X1 U7612 ( .A1(INSTQUEUE_REG_7__6__SCAN_IN), .A2(n6632), .B1(n6815), 
        .B2(n6630), .ZN(n6628) );
  OAI211_X1 U7613 ( .C1(n6635), .C2(n6819), .A(n6629), .B(n6628), .ZN(U3082)
         );
  AOI22_X1 U7614 ( .A1(n6631), .A2(n6823), .B1(n6825), .B2(n6630), .ZN(n6634)
         );
  AOI22_X1 U7615 ( .A1(INSTQUEUE_REG_7__7__SCAN_IN), .A2(n6632), .B1(n6820), 
        .B2(n6642), .ZN(n6633) );
  OAI211_X1 U7616 ( .C1(n6635), .C2(n6829), .A(n6634), .B(n6633), .ZN(U3083)
         );
  NAND2_X1 U7617 ( .A1(n6636), .A2(n6643), .ZN(n6640) );
  INV_X1 U7618 ( .A(n6637), .ZN(n6639) );
  NAND2_X1 U7619 ( .A1(n6639), .A2(n6638), .ZN(n6730) );
  OAI22_X1 U7620 ( .A1(n6640), .A2(n6645), .B1(n6725), .B2(n6730), .ZN(n6667)
         );
  NOR2_X1 U7621 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6641), .ZN(n6666)
         );
  AOI22_X1 U7622 ( .A1(n6832), .A2(n6667), .B1(n6833), .B2(n6666), .ZN(n6651)
         );
  OAI21_X1 U7623 ( .B1(n6668), .B2(n6642), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n6644) );
  OAI211_X1 U7624 ( .C1(n6731), .C2(n6645), .A(n6644), .B(n6643), .ZN(n6649)
         );
  AOI21_X1 U7625 ( .B1(n6730), .B2(STATE2_REG_2__SCAN_IN), .A(n6646), .ZN(
        n6718) );
  OAI211_X1 U7626 ( .C1(n7000), .C2(n6666), .A(n6729), .B(n6718), .ZN(n6647)
         );
  INV_X1 U7627 ( .A(n6647), .ZN(n6648) );
  NAND2_X1 U7628 ( .A1(n6649), .A2(n6648), .ZN(n6669) );
  AOI22_X1 U7629 ( .A1(n6669), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n6839), 
        .B2(n6668), .ZN(n6650) );
  OAI211_X1 U7630 ( .C1(n6690), .C2(n6672), .A(n6651), .B(n6650), .ZN(U3084)
         );
  AOI22_X1 U7631 ( .A1(n6736), .A2(n6667), .B1(n6784), .B2(n6666), .ZN(n6653)
         );
  AOI22_X1 U7632 ( .A1(n6669), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n6668), 
        .B2(n6786), .ZN(n6652) );
  OAI211_X1 U7633 ( .C1(n6654), .C2(n6672), .A(n6653), .B(n6652), .ZN(U3085)
         );
  AOI22_X1 U7634 ( .A1(n6740), .A2(n6667), .B1(n6790), .B2(n6666), .ZN(n6656)
         );
  AOI22_X1 U7635 ( .A1(n6669), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n6668), 
        .B2(n6791), .ZN(n6655) );
  OAI211_X1 U7636 ( .C1(n6657), .C2(n6672), .A(n6656), .B(n6655), .ZN(U3086)
         );
  AOI22_X1 U7637 ( .A1(n6744), .A2(n6667), .B1(n6796), .B2(n6666), .ZN(n6659)
         );
  AOI22_X1 U7638 ( .A1(n6669), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n6668), 
        .B2(n6798), .ZN(n6658) );
  OAI211_X1 U7639 ( .C1(n6699), .C2(n6672), .A(n6659), .B(n6658), .ZN(U3087)
         );
  AOI22_X1 U7640 ( .A1(n6748), .A2(n6667), .B1(n6802), .B2(n6666), .ZN(n6661)
         );
  AOI22_X1 U7641 ( .A1(n6669), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n6668), 
        .B2(n6804), .ZN(n6660) );
  OAI211_X1 U7642 ( .C1(n6702), .C2(n6672), .A(n6661), .B(n6660), .ZN(U3088)
         );
  AOI22_X1 U7643 ( .A1(n6752), .A2(n6667), .B1(n6808), .B2(n6666), .ZN(n6663)
         );
  AOI22_X1 U7644 ( .A1(n6669), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n6668), 
        .B2(n6810), .ZN(n6662) );
  OAI211_X1 U7645 ( .C1(n6705), .C2(n6672), .A(n6663), .B(n6662), .ZN(U3089)
         );
  AOI22_X1 U7646 ( .A1(n6756), .A2(n6667), .B1(n6814), .B2(n6666), .ZN(n6665)
         );
  AOI22_X1 U7647 ( .A1(n6669), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n6668), 
        .B2(n6816), .ZN(n6664) );
  OAI211_X1 U7648 ( .C1(n6709), .C2(n6672), .A(n6665), .B(n6664), .ZN(U3090)
         );
  AOI22_X1 U7649 ( .A1(n6762), .A2(n6667), .B1(n6823), .B2(n6666), .ZN(n6671)
         );
  AOI22_X1 U7650 ( .A1(n6669), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n6668), 
        .B2(n6820), .ZN(n6670) );
  OAI211_X1 U7651 ( .C1(n6673), .C2(n6672), .A(n6671), .B(n6670), .ZN(U3091)
         );
  INV_X1 U7652 ( .A(n6674), .ZN(n6675) );
  NOR2_X1 U7653 ( .A1(n6677), .A2(n6864), .ZN(n6710) );
  AOI22_X1 U7654 ( .A1(n6839), .A2(n6763), .B1(n6833), .B2(n6710), .ZN(n6689)
         );
  AOI21_X1 U7655 ( .B1(n6679), .B2(n6678), .A(n6776), .ZN(n6684) );
  INV_X1 U7656 ( .A(n6680), .ZN(n6682) );
  AOI21_X1 U7657 ( .B1(n6682), .B2(n6681), .A(n6710), .ZN(n6686) );
  AOI22_X1 U7658 ( .A1(n6684), .A2(n6686), .B1(n6685), .B2(n6776), .ZN(n6683)
         );
  NAND2_X1 U7659 ( .A1(n6780), .A2(n6683), .ZN(n6713) );
  INV_X1 U7660 ( .A(n6684), .ZN(n6687) );
  OAI22_X1 U7661 ( .A1(n6687), .A2(n6686), .B1(n6685), .B2(n6773), .ZN(n6712)
         );
  AOI22_X1 U7662 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n6713), .B1(n6832), 
        .B2(n6712), .ZN(n6688) );
  OAI211_X1 U7663 ( .C1(n6690), .C2(n6708), .A(n6689), .B(n6688), .ZN(U3108)
         );
  AOI22_X1 U7664 ( .A1(n6711), .A2(n6785), .B1(n6784), .B2(n6710), .ZN(n6692)
         );
  AOI22_X1 U7665 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(n6713), .B1(n6736), 
        .B2(n6712), .ZN(n6691) );
  OAI211_X1 U7666 ( .C1(n6693), .C2(n6716), .A(n6692), .B(n6691), .ZN(U3109)
         );
  AOI22_X1 U7667 ( .A1(n6711), .A2(n6792), .B1(n6790), .B2(n6710), .ZN(n6695)
         );
  AOI22_X1 U7668 ( .A1(INSTQUEUE_REG_11__2__SCAN_IN), .A2(n6713), .B1(n6740), 
        .B2(n6712), .ZN(n6694) );
  OAI211_X1 U7669 ( .C1(n6696), .C2(n6716), .A(n6695), .B(n6694), .ZN(U3110)
         );
  AOI22_X1 U7670 ( .A1(n6763), .A2(n6798), .B1(n6796), .B2(n6710), .ZN(n6698)
         );
  AOI22_X1 U7671 ( .A1(INSTQUEUE_REG_11__3__SCAN_IN), .A2(n6713), .B1(n6744), 
        .B2(n6712), .ZN(n6697) );
  OAI211_X1 U7672 ( .C1(n6699), .C2(n6708), .A(n6698), .B(n6697), .ZN(U3111)
         );
  AOI22_X1 U7673 ( .A1(n6763), .A2(n6804), .B1(n6802), .B2(n6710), .ZN(n6701)
         );
  AOI22_X1 U7674 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n6713), .B1(n6748), 
        .B2(n6712), .ZN(n6700) );
  OAI211_X1 U7675 ( .C1(n6702), .C2(n6708), .A(n6701), .B(n6700), .ZN(U3112)
         );
  AOI22_X1 U7676 ( .A1(n6763), .A2(n6810), .B1(n6808), .B2(n6710), .ZN(n6704)
         );
  AOI22_X1 U7677 ( .A1(INSTQUEUE_REG_11__5__SCAN_IN), .A2(n6713), .B1(n6752), 
        .B2(n6712), .ZN(n6703) );
  OAI211_X1 U7678 ( .C1(n6705), .C2(n6708), .A(n6704), .B(n6703), .ZN(U3113)
         );
  AOI22_X1 U7679 ( .A1(n6763), .A2(n6816), .B1(n6814), .B2(n6710), .ZN(n6707)
         );
  AOI22_X1 U7680 ( .A1(INSTQUEUE_REG_11__6__SCAN_IN), .A2(n6713), .B1(n6756), 
        .B2(n6712), .ZN(n6706) );
  OAI211_X1 U7681 ( .C1(n6709), .C2(n6708), .A(n6707), .B(n6706), .ZN(U3114)
         );
  AOI22_X1 U7682 ( .A1(n6825), .A2(n6711), .B1(n6823), .B2(n6710), .ZN(n6715)
         );
  AOI22_X1 U7683 ( .A1(INSTQUEUE_REG_11__7__SCAN_IN), .A2(n6713), .B1(n6762), 
        .B2(n6712), .ZN(n6714) );
  OAI211_X1 U7684 ( .C1(n6717), .C2(n6716), .A(n6715), .B(n6714), .ZN(U3115)
         );
  INV_X1 U7685 ( .A(n6718), .ZN(n6728) );
  NAND3_X1 U7686 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n6859), .ZN(n6775) );
  NOR2_X1 U7687 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6775), .ZN(n6760)
         );
  NOR3_X1 U7688 ( .A1(n6763), .A2(n6824), .A3(n6776), .ZN(n6724) );
  OAI22_X1 U7689 ( .A1(n6724), .A2(n6723), .B1(n6722), .B2(n6721), .ZN(n6726)
         );
  OAI211_X1 U7690 ( .C1(n6760), .C2(n7000), .A(n6726), .B(n6725), .ZN(n6727)
         );
  OAI22_X1 U7691 ( .A1(n6732), .A2(n6731), .B1(n6730), .B2(n6729), .ZN(n6761)
         );
  AOI22_X1 U7692 ( .A1(n6832), .A2(n6761), .B1(n6833), .B2(n6760), .ZN(n6734)
         );
  AOI22_X1 U7693 ( .A1(n6836), .A2(n6763), .B1(n6824), .B2(n6839), .ZN(n6733)
         );
  OAI211_X1 U7694 ( .C1(n6767), .C2(n6735), .A(n6734), .B(n6733), .ZN(U3116)
         );
  INV_X1 U7695 ( .A(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n6739) );
  AOI22_X1 U7696 ( .A1(n6736), .A2(n6761), .B1(n6784), .B2(n6760), .ZN(n6738)
         );
  AOI22_X1 U7697 ( .A1(n6785), .A2(n6763), .B1(n6824), .B2(n6786), .ZN(n6737)
         );
  OAI211_X1 U7698 ( .C1(n6767), .C2(n6739), .A(n6738), .B(n6737), .ZN(U3117)
         );
  INV_X1 U7699 ( .A(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n6743) );
  AOI22_X1 U7700 ( .A1(n6740), .A2(n6761), .B1(n6790), .B2(n6760), .ZN(n6742)
         );
  AOI22_X1 U7701 ( .A1(n6792), .A2(n6763), .B1(n6824), .B2(n6791), .ZN(n6741)
         );
  OAI211_X1 U7702 ( .C1(n6767), .C2(n6743), .A(n6742), .B(n6741), .ZN(U3118)
         );
  INV_X1 U7703 ( .A(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n6747) );
  AOI22_X1 U7704 ( .A1(n6744), .A2(n6761), .B1(n6796), .B2(n6760), .ZN(n6746)
         );
  AOI22_X1 U7705 ( .A1(n6797), .A2(n6763), .B1(n6824), .B2(n6798), .ZN(n6745)
         );
  OAI211_X1 U7706 ( .C1(n6767), .C2(n6747), .A(n6746), .B(n6745), .ZN(U3119)
         );
  INV_X1 U7707 ( .A(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n6751) );
  AOI22_X1 U7708 ( .A1(n6748), .A2(n6761), .B1(n6802), .B2(n6760), .ZN(n6750)
         );
  AOI22_X1 U7709 ( .A1(n6803), .A2(n6763), .B1(n6824), .B2(n6804), .ZN(n6749)
         );
  OAI211_X1 U7710 ( .C1(n6767), .C2(n6751), .A(n6750), .B(n6749), .ZN(U3120)
         );
  AOI22_X1 U7711 ( .A1(n6752), .A2(n6761), .B1(n6808), .B2(n6760), .ZN(n6754)
         );
  AOI22_X1 U7712 ( .A1(n6809), .A2(n6763), .B1(n6824), .B2(n6810), .ZN(n6753)
         );
  OAI211_X1 U7713 ( .C1(n6767), .C2(n6755), .A(n6754), .B(n6753), .ZN(U3121)
         );
  INV_X1 U7714 ( .A(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n6759) );
  AOI22_X1 U7715 ( .A1(n6756), .A2(n6761), .B1(n6814), .B2(n6760), .ZN(n6758)
         );
  AOI22_X1 U7716 ( .A1(n6815), .A2(n6763), .B1(n6824), .B2(n6816), .ZN(n6757)
         );
  OAI211_X1 U7717 ( .C1(n6767), .C2(n6759), .A(n6758), .B(n6757), .ZN(U3122)
         );
  INV_X1 U7718 ( .A(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n6766) );
  AOI22_X1 U7719 ( .A1(n6762), .A2(n6761), .B1(n6823), .B2(n6760), .ZN(n6765)
         );
  AOI22_X1 U7720 ( .A1(n6825), .A2(n6763), .B1(n6824), .B2(n6820), .ZN(n6764)
         );
  OAI211_X1 U7721 ( .C1(n6767), .C2(n6766), .A(n6765), .B(n6764), .ZN(U3123)
         );
  NOR2_X1 U7722 ( .A1(n6768), .A2(n6776), .ZN(n6777) );
  INV_X1 U7723 ( .A(n6777), .ZN(n6772) );
  NOR2_X1 U7724 ( .A1(n6769), .A2(n6775), .ZN(n6822) );
  AOI21_X1 U7725 ( .B1(n6771), .B2(n6770), .A(n6822), .ZN(n6778) );
  OAI22_X1 U7726 ( .A1(n6773), .A2(n6775), .B1(n6772), .B2(n6778), .ZN(n6774)
         );
  AOI22_X1 U7727 ( .A1(n6833), .A2(n6822), .B1(n6824), .B2(n6836), .ZN(n6782)
         );
  AOI22_X1 U7728 ( .A1(n6778), .A2(n6777), .B1(n6776), .B2(n6775), .ZN(n6779)
         );
  NAND2_X1 U7729 ( .A1(n6780), .A2(n6779), .ZN(n6826) );
  AOI22_X1 U7730 ( .A1(n6826), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n6839), 
        .B2(n6821), .ZN(n6781) );
  OAI211_X1 U7731 ( .C1(n6830), .C2(n6783), .A(n6782), .B(n6781), .ZN(U3124)
         );
  AOI22_X1 U7732 ( .A1(n6785), .A2(n6824), .B1(n6784), .B2(n6822), .ZN(n6788)
         );
  AOI22_X1 U7733 ( .A1(n6826), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n6786), 
        .B2(n6821), .ZN(n6787) );
  OAI211_X1 U7734 ( .C1(n6830), .C2(n6789), .A(n6788), .B(n6787), .ZN(U3125)
         );
  AOI22_X1 U7735 ( .A1(n6791), .A2(n6821), .B1(n6790), .B2(n6822), .ZN(n6794)
         );
  AOI22_X1 U7736 ( .A1(n6826), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n6792), 
        .B2(n6824), .ZN(n6793) );
  OAI211_X1 U7737 ( .C1(n6830), .C2(n6795), .A(n6794), .B(n6793), .ZN(U3126)
         );
  AOI22_X1 U7738 ( .A1(n6797), .A2(n6824), .B1(n6796), .B2(n6822), .ZN(n6800)
         );
  AOI22_X1 U7739 ( .A1(n6826), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n6798), 
        .B2(n6821), .ZN(n6799) );
  OAI211_X1 U7740 ( .C1(n6830), .C2(n6801), .A(n6800), .B(n6799), .ZN(U3127)
         );
  AOI22_X1 U7741 ( .A1(n6803), .A2(n6824), .B1(n6802), .B2(n6822), .ZN(n6806)
         );
  AOI22_X1 U7742 ( .A1(n6826), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n6804), 
        .B2(n6821), .ZN(n6805) );
  OAI211_X1 U7743 ( .C1(n6830), .C2(n6807), .A(n6806), .B(n6805), .ZN(U3128)
         );
  AOI22_X1 U7744 ( .A1(n6809), .A2(n6824), .B1(n6808), .B2(n6822), .ZN(n6812)
         );
  AOI22_X1 U7745 ( .A1(n6826), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n6810), 
        .B2(n6821), .ZN(n6811) );
  OAI211_X1 U7746 ( .C1(n6830), .C2(n6813), .A(n6812), .B(n6811), .ZN(U3129)
         );
  AOI22_X1 U7747 ( .A1(n6815), .A2(n6824), .B1(n6814), .B2(n6822), .ZN(n6818)
         );
  AOI22_X1 U7748 ( .A1(n6826), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n6816), 
        .B2(n6821), .ZN(n6817) );
  OAI211_X1 U7749 ( .C1(n6830), .C2(n6819), .A(n6818), .B(n6817), .ZN(U3130)
         );
  AOI22_X1 U7750 ( .A1(n6823), .A2(n6822), .B1(n6821), .B2(n6820), .ZN(n6828)
         );
  AOI22_X1 U7751 ( .A1(n6826), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n6825), 
        .B2(n6824), .ZN(n6827) );
  OAI211_X1 U7752 ( .C1(n6830), .C2(n6829), .A(n6828), .B(n6827), .ZN(U3131)
         );
  AOI22_X1 U7753 ( .A1(n6834), .A2(n6833), .B1(n6832), .B2(n6831), .ZN(n6841)
         );
  INV_X1 U7754 ( .A(n6835), .ZN(n6838) );
  AOI22_X1 U7755 ( .A1(n6839), .A2(n6838), .B1(n6837), .B2(n6836), .ZN(n6840)
         );
  OAI211_X1 U7756 ( .C1(n6843), .C2(n6842), .A(n6841), .B(n6840), .ZN(U3140)
         );
  AND2_X1 U7757 ( .A1(n6845), .A2(n6844), .ZN(n6865) );
  NAND2_X1 U7758 ( .A1(n6845), .A2(n6846), .ZN(n6862) );
  OR2_X1 U7759 ( .A1(n3776), .A2(n6847), .ZN(n6850) );
  NAND2_X1 U7760 ( .A1(n6848), .A2(n3289), .ZN(n6849) );
  NAND2_X1 U7761 ( .A1(n6850), .A2(n6849), .ZN(n7001) );
  INV_X1 U7762 ( .A(n6851), .ZN(n6852) );
  NAND2_X1 U7763 ( .A1(n6852), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n7009) );
  NAND2_X1 U7764 ( .A1(n7009), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6853) );
  NOR2_X1 U7765 ( .A1(n7001), .A2(n6853), .ZN(n6855) );
  INV_X1 U7766 ( .A(n6855), .ZN(n6860) );
  INV_X1 U7767 ( .A(n6854), .ZN(n6856) );
  OAI22_X1 U7768 ( .A1(n6857), .A2(n6856), .B1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n6855), .ZN(n6858) );
  OAI21_X1 U7769 ( .B1(n6860), .B2(n6859), .A(n6858), .ZN(n6861) );
  AOI222_X1 U7770 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n6862), .B1(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n6861), .C1(n6862), .C2(n6861), 
        .ZN(n6863) );
  AOI222_X1 U7771 ( .A1(n6865), .A2(n6864), .B1(n6865), .B2(n6863), .C1(n6864), 
        .C2(n6863), .ZN(n6868) );
  OAI21_X1 U7772 ( .B1(FLUSH_REG_SCAN_IN), .B2(MORE_REG_SCAN_IN), .A(n6866), 
        .ZN(n6867) );
  OAI21_X1 U7773 ( .B1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(n6868), .A(n6867), 
        .ZN(n6882) );
  AND2_X1 U7774 ( .A1(n6870), .A2(n6869), .ZN(n6871) );
  OR2_X1 U7775 ( .A1(n6891), .A2(n6871), .ZN(n6875) );
  INV_X1 U7776 ( .A(n6872), .ZN(n6873) );
  NAND2_X1 U7777 ( .A1(n6891), .A2(n6873), .ZN(n6874) );
  OAI211_X1 U7778 ( .C1(n6877), .C2(n6876), .A(n6875), .B(n6874), .ZN(n7021)
         );
  NOR2_X1 U7779 ( .A1(n7021), .A2(n6878), .ZN(n6879) );
  NAND2_X1 U7780 ( .A1(n6880), .A2(n6879), .ZN(n6881) );
  NOR2_X1 U7781 ( .A1(n6882), .A2(n6881), .ZN(n6899) );
  OR2_X1 U7782 ( .A1(n6884), .A2(n6883), .ZN(n6888) );
  AOI21_X1 U7783 ( .B1(STATE2_REG_1__SCAN_IN), .B2(READY_N), .A(
        STATE2_REG_0__SCAN_IN), .ZN(n6885) );
  INV_X1 U7784 ( .A(n6885), .ZN(n6886) );
  AND2_X1 U7785 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n6886), .ZN(n6887) );
  AND2_X1 U7786 ( .A1(n6888), .A2(n6887), .ZN(n6892) );
  OAI221_X1 U7787 ( .B1(n6894), .B2(n6899), .C1(n6894), .C2(n7002), .A(n6892), 
        .ZN(n6999) );
  OAI21_X1 U7788 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n7024), .A(n6999), .ZN(
        n6900) );
  AOI221_X1 U7789 ( .B1(n6890), .B2(STATE2_REG_0__SCAN_IN), .C1(n6900), .C2(
        STATE2_REG_0__SCAN_IN), .A(n6889), .ZN(n6898) );
  INV_X1 U7790 ( .A(n6891), .ZN(n6896) );
  NAND2_X1 U7791 ( .A1(STATE2_REG_3__SCAN_IN), .A2(n7027), .ZN(n6895) );
  INV_X1 U7792 ( .A(n6892), .ZN(n6893) );
  OAI211_X1 U7793 ( .C1(n6896), .C2(n6895), .A(n6894), .B(n6893), .ZN(n6897)
         );
  OAI211_X1 U7794 ( .C1(n6899), .C2(n6901), .A(n6898), .B(n6897), .ZN(U3148)
         );
  OAI211_X1 U7795 ( .C1(STATE2_REG_0__SCAN_IN), .C2(STATE2_REG_2__SCAN_IN), 
        .A(STATE2_REG_1__SCAN_IN), .B(n6900), .ZN(n6906) );
  OAI21_X1 U7796 ( .B1(READY_N), .B2(n6902), .A(n6901), .ZN(n6904) );
  AOI21_X1 U7797 ( .B1(n6904), .B2(n6999), .A(n6903), .ZN(n6905) );
  NAND2_X1 U7798 ( .A1(n6906), .A2(n6905), .ZN(U3149) );
  OAI221_X1 U7799 ( .B1(STATE2_REG_2__SCAN_IN), .B2(STATE2_REG_0__SCAN_IN), 
        .C1(STATE2_REG_2__SCAN_IN), .C2(n7024), .A(n6998), .ZN(n6908) );
  OAI21_X1 U7800 ( .B1(n7027), .B2(n6908), .A(n6907), .ZN(U3150) );
  NOR2_X1 U7801 ( .A1(n6997), .A2(n6909), .ZN(U3151) );
  AND2_X1 U7802 ( .A1(DATAWIDTH_REG_30__SCAN_IN), .A2(n6993), .ZN(U3152) );
  AND2_X1 U7803 ( .A1(n6993), .A2(DATAWIDTH_REG_29__SCAN_IN), .ZN(U3153) );
  AND2_X1 U7804 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(n6993), .ZN(U3154) );
  AND2_X1 U7805 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(n6993), .ZN(U3155) );
  AND2_X1 U7806 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(n6993), .ZN(U3156) );
  AND2_X1 U7807 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(n6993), .ZN(U3157) );
  AND2_X1 U7808 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(n6993), .ZN(U3158) );
  AND2_X1 U7809 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(n6993), .ZN(U3159) );
  AND2_X1 U7810 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(n6993), .ZN(U3160) );
  AND2_X1 U7811 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(n6993), .ZN(U3161) );
  AND2_X1 U7812 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(n6993), .ZN(U3162) );
  AND2_X1 U7813 ( .A1(n6993), .A2(DATAWIDTH_REG_19__SCAN_IN), .ZN(U3163) );
  AND2_X1 U7814 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(n6993), .ZN(U3164) );
  AND2_X1 U7815 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(n6993), .ZN(U3165) );
  AND2_X1 U7816 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(n6993), .ZN(U3166) );
  AND2_X1 U7817 ( .A1(DATAWIDTH_REG_15__SCAN_IN), .A2(n6993), .ZN(U3167) );
  AND2_X1 U7818 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(n6993), .ZN(U3168) );
  AND2_X1 U7819 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(n6993), .ZN(U3169) );
  AND2_X1 U7820 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(n6993), .ZN(U3170) );
  AND2_X1 U7821 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(n6993), .ZN(U3171) );
  AND2_X1 U7822 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(n6993), .ZN(U3172) );
  AND2_X1 U7823 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(n6993), .ZN(U3173) );
  AND2_X1 U7824 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(n6993), .ZN(U3174) );
  AND2_X1 U7825 ( .A1(DATAWIDTH_REG_7__SCAN_IN), .A2(n6993), .ZN(U3175) );
  AND2_X1 U7826 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(n6993), .ZN(U3176) );
  NOR2_X1 U7827 ( .A1(n6997), .A2(n6910), .ZN(U3177) );
  AND2_X1 U7828 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(n6993), .ZN(U3178) );
  NOR2_X1 U7829 ( .A1(n6997), .A2(n6911), .ZN(U3179) );
  AND2_X1 U7830 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(n6993), .ZN(U3180) );
  AOI22_X1 U7831 ( .A1(STATE_REG_1__SCAN_IN), .A2(READY_N), .B1(
        STATE_REG_2__SCAN_IN), .B2(HOLD), .ZN(n6925) );
  AND2_X1 U7832 ( .A1(STATE_REG_1__SCAN_IN), .A2(HOLD), .ZN(n6915) );
  INV_X1 U7833 ( .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6913) );
  INV_X1 U7834 ( .A(NA_N), .ZN(n6922) );
  AOI211_X1 U7835 ( .C1(STATE_REG_2__SCAN_IN), .C2(n6922), .A(
        STATE_REG_0__SCAN_IN), .B(n6921), .ZN(n6927) );
  AOI221_X1 U7836 ( .B1(n6915), .B2(n7019), .C1(n6913), .C2(n7019), .A(n6927), 
        .ZN(n6912) );
  OAI21_X1 U7837 ( .B1(n6921), .B2(n6925), .A(n6912), .ZN(U3181) );
  NOR2_X1 U7838 ( .A1(n6919), .A2(n6913), .ZN(n6923) );
  NAND2_X1 U7839 ( .A1(STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n6914) );
  OAI21_X1 U7840 ( .B1(n6923), .B2(n6915), .A(n6914), .ZN(n6916) );
  OAI211_X1 U7841 ( .C1(n7024), .C2(n6918), .A(n6917), .B(n6916), .ZN(U3182)
         );
  AOI221_X1 U7842 ( .B1(NA_N), .B2(STATE_REG_1__SCAN_IN), .C1(n7024), .C2(
        STATE_REG_1__SCAN_IN), .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6920) );
  AOI221_X1 U7843 ( .B1(STATE_REG_2__SCAN_IN), .B2(HOLD), .C1(n6920), .C2(HOLD), .A(n6919), .ZN(n6926) );
  AOI21_X1 U7844 ( .B1(n6923), .B2(n6922), .A(n6921), .ZN(n6924) );
  OAI22_X1 U7845 ( .A1(n6927), .A2(n6926), .B1(n6925), .B2(n6924), .ZN(U3183)
         );
  NAND2_X1 U7846 ( .A1(STATE_REG_2__SCAN_IN), .A2(n7032), .ZN(n6986) );
  NOR2_X1 U7847 ( .A1(STATE_REG_2__SCAN_IN), .A2(n7019), .ZN(n6979) );
  AOI22_X1 U7848 ( .A1(REIP_REG_2__SCAN_IN), .A2(n6979), .B1(
        ADDRESS_REG_0__SCAN_IN), .B2(n7019), .ZN(n6928) );
  OAI21_X1 U7849 ( .B1(n7015), .B2(n6986), .A(n6928), .ZN(U3184) );
  INV_X1 U7850 ( .A(n6986), .ZN(n6975) );
  AOI22_X1 U7851 ( .A1(REIP_REG_2__SCAN_IN), .A2(n6975), .B1(
        ADDRESS_REG_1__SCAN_IN), .B2(n7019), .ZN(n6929) );
  OAI21_X1 U7852 ( .B1(n6931), .B2(n6982), .A(n6929), .ZN(U3185) );
  AOI22_X1 U7853 ( .A1(REIP_REG_4__SCAN_IN), .A2(n6979), .B1(
        ADDRESS_REG_2__SCAN_IN), .B2(n7019), .ZN(n6930) );
  OAI21_X1 U7854 ( .B1(n6931), .B2(n6986), .A(n6930), .ZN(U3186) );
  OAI222_X1 U7855 ( .A1(n6986), .A2(n6933), .B1(n6932), .B2(n7032), .C1(n6935), 
        .C2(n6982), .ZN(U3187) );
  AOI22_X1 U7856 ( .A1(REIP_REG_6__SCAN_IN), .A2(n6979), .B1(
        ADDRESS_REG_4__SCAN_IN), .B2(n7019), .ZN(n6934) );
  OAI21_X1 U7857 ( .B1(n6935), .B2(n6986), .A(n6934), .ZN(U3188) );
  OAI222_X1 U7858 ( .A1(n6986), .A2(n6938), .B1(n6937), .B2(n7032), .C1(n6936), 
        .C2(n6982), .ZN(U3189) );
  AOI22_X1 U7859 ( .A1(REIP_REG_7__SCAN_IN), .A2(n6975), .B1(
        ADDRESS_REG_6__SCAN_IN), .B2(n7019), .ZN(n6939) );
  OAI21_X1 U7860 ( .B1(n6941), .B2(n6982), .A(n6939), .ZN(U3190) );
  AOI22_X1 U7861 ( .A1(REIP_REG_9__SCAN_IN), .A2(n6979), .B1(
        ADDRESS_REG_7__SCAN_IN), .B2(n7019), .ZN(n6940) );
  OAI21_X1 U7862 ( .B1(n6941), .B2(n6986), .A(n6940), .ZN(U3191) );
  AOI22_X1 U7863 ( .A1(REIP_REG_9__SCAN_IN), .A2(n6975), .B1(
        ADDRESS_REG_8__SCAN_IN), .B2(n7019), .ZN(n6942) );
  OAI21_X1 U7864 ( .B1(n6943), .B2(n6982), .A(n6942), .ZN(U3192) );
  AOI22_X1 U7865 ( .A1(REIP_REG_10__SCAN_IN), .A2(n6975), .B1(
        ADDRESS_REG_9__SCAN_IN), .B2(n7019), .ZN(n6944) );
  OAI21_X1 U7866 ( .B1(n6945), .B2(n6982), .A(n6944), .ZN(U3193) );
  AOI22_X1 U7867 ( .A1(REIP_REG_11__SCAN_IN), .A2(n6975), .B1(
        ADDRESS_REG_10__SCAN_IN), .B2(n7019), .ZN(n6946) );
  OAI21_X1 U7868 ( .B1(n6948), .B2(n6982), .A(n6946), .ZN(U3194) );
  AOI22_X1 U7869 ( .A1(REIP_REG_13__SCAN_IN), .A2(n6979), .B1(
        ADDRESS_REG_11__SCAN_IN), .B2(n7019), .ZN(n6947) );
  OAI21_X1 U7870 ( .B1(n6948), .B2(n6986), .A(n6947), .ZN(U3195) );
  AOI22_X1 U7871 ( .A1(REIP_REG_14__SCAN_IN), .A2(n6979), .B1(
        ADDRESS_REG_12__SCAN_IN), .B2(n7019), .ZN(n6949) );
  OAI21_X1 U7872 ( .B1(n6950), .B2(n6986), .A(n6949), .ZN(U3196) );
  OAI222_X1 U7873 ( .A1(n6982), .A2(n6953), .B1(n6952), .B2(n7032), .C1(n6951), 
        .C2(n6986), .ZN(U3197) );
  AOI22_X1 U7874 ( .A1(REIP_REG_15__SCAN_IN), .A2(n6975), .B1(
        ADDRESS_REG_14__SCAN_IN), .B2(n7019), .ZN(n6954) );
  OAI21_X1 U7875 ( .B1(n6955), .B2(n6982), .A(n6954), .ZN(U3198) );
  AOI222_X1 U7876 ( .A1(n6975), .A2(REIP_REG_16__SCAN_IN), .B1(
        ADDRESS_REG_15__SCAN_IN), .B2(n7019), .C1(REIP_REG_17__SCAN_IN), .C2(
        n6979), .ZN(n6956) );
  INV_X1 U7877 ( .A(n6956), .ZN(U3199) );
  AOI22_X1 U7878 ( .A1(REIP_REG_17__SCAN_IN), .A2(n6975), .B1(
        ADDRESS_REG_16__SCAN_IN), .B2(n7019), .ZN(n6957) );
  OAI21_X1 U7879 ( .B1(n6958), .B2(n6982), .A(n6957), .ZN(U3200) );
  OAI222_X1 U7880 ( .A1(n6982), .A2(n6962), .B1(n6959), .B2(n7032), .C1(n6958), 
        .C2(n6986), .ZN(U3201) );
  OAI222_X1 U7881 ( .A1(n6986), .A2(n6962), .B1(n6961), .B2(n7032), .C1(n6960), 
        .C2(n6982), .ZN(U3202) );
  AOI22_X1 U7882 ( .A1(REIP_REG_20__SCAN_IN), .A2(n6975), .B1(
        ADDRESS_REG_19__SCAN_IN), .B2(n7019), .ZN(n6963) );
  OAI21_X1 U7883 ( .B1(n5728), .B2(n6982), .A(n6963), .ZN(U3203) );
  AOI22_X1 U7884 ( .A1(REIP_REG_22__SCAN_IN), .A2(n6979), .B1(
        ADDRESS_REG_20__SCAN_IN), .B2(n7019), .ZN(n6964) );
  OAI21_X1 U7885 ( .B1(n5728), .B2(n6986), .A(n6964), .ZN(U3204) );
  AOI22_X1 U7886 ( .A1(REIP_REG_22__SCAN_IN), .A2(n6975), .B1(
        ADDRESS_REG_21__SCAN_IN), .B2(n7019), .ZN(n6965) );
  OAI21_X1 U7887 ( .B1(n6967), .B2(n6982), .A(n6965), .ZN(U3205) );
  AOI22_X1 U7888 ( .A1(REIP_REG_24__SCAN_IN), .A2(n6979), .B1(
        ADDRESS_REG_22__SCAN_IN), .B2(n7019), .ZN(n6966) );
  OAI21_X1 U7889 ( .B1(n6967), .B2(n6986), .A(n6966), .ZN(U3206) );
  OAI222_X1 U7890 ( .A1(n6982), .A2(n6971), .B1(n6969), .B2(n7032), .C1(n6968), 
        .C2(n6986), .ZN(U3207) );
  AOI22_X1 U7891 ( .A1(REIP_REG_26__SCAN_IN), .A2(n6979), .B1(
        ADDRESS_REG_24__SCAN_IN), .B2(n7019), .ZN(n6970) );
  OAI21_X1 U7892 ( .B1(n6971), .B2(n6986), .A(n6970), .ZN(U3208) );
  INV_X1 U7893 ( .A(REIP_REG_26__SCAN_IN), .ZN(n6974) );
  OAI222_X1 U7894 ( .A1(n6986), .A2(n6974), .B1(n6973), .B2(n7032), .C1(n6972), 
        .C2(n6982), .ZN(U3209) );
  AOI22_X1 U7895 ( .A1(REIP_REG_27__SCAN_IN), .A2(n6975), .B1(
        ADDRESS_REG_26__SCAN_IN), .B2(n7019), .ZN(n6976) );
  OAI21_X1 U7896 ( .B1(n6978), .B2(n6982), .A(n6976), .ZN(U3210) );
  OAI222_X1 U7897 ( .A1(n6986), .A2(n6978), .B1(n6977), .B2(n7032), .C1(n6981), 
        .C2(n6982), .ZN(U3211) );
  AOI22_X1 U7898 ( .A1(REIP_REG_30__SCAN_IN), .A2(n6979), .B1(
        ADDRESS_REG_28__SCAN_IN), .B2(n7019), .ZN(n6980) );
  OAI21_X1 U7899 ( .B1(n6981), .B2(n6986), .A(n6980), .ZN(U3212) );
  INV_X1 U7900 ( .A(ADDRESS_REG_29__SCAN_IN), .ZN(n6984) );
  OAI222_X1 U7901 ( .A1(n6986), .A2(n6985), .B1(n6984), .B2(n7032), .C1(n6983), 
        .C2(n6982), .ZN(U3213) );
  INV_X1 U7902 ( .A(BE_N_REG_3__SCAN_IN), .ZN(n6987) );
  AOI22_X1 U7903 ( .A1(n7032), .A2(n6988), .B1(n6987), .B2(n7019), .ZN(U3445)
         );
  MUX2_X1 U7904 ( .A(BE_N_REG_2__SCAN_IN), .B(BYTEENABLE_REG_2__SCAN_IN), .S(
        n7032), .Z(U3446) );
  AOI22_X1 U7905 ( .A1(n7032), .A2(n6990), .B1(n6989), .B2(n7019), .ZN(U3447)
         );
  INV_X1 U7906 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n7017) );
  AOI22_X1 U7907 ( .A1(n7032), .A2(n7017), .B1(n6991), .B2(n7019), .ZN(U3448)
         );
  INV_X1 U7908 ( .A(DATAWIDTH_REG_0__SCAN_IN), .ZN(n6994) );
  INV_X1 U7909 ( .A(n6995), .ZN(n6992) );
  AOI21_X1 U7910 ( .B1(n6994), .B2(n6993), .A(n6992), .ZN(U3451) );
  OAI21_X1 U7911 ( .B1(n6997), .B2(n6996), .A(n6995), .ZN(U3452) );
  OAI221_X1 U7912 ( .B1(n7000), .B2(STATE2_REG_0__SCAN_IN), .C1(n7000), .C2(
        n6999), .A(n6998), .ZN(U3453) );
  INV_X1 U7913 ( .A(n7001), .ZN(n7003) );
  OAI22_X1 U7914 ( .A1(n7003), .A2(n7008), .B1(INSTADDRPOINTER_REG_0__SCAN_IN), 
        .B2(n7002), .ZN(n7005) );
  OAI22_X1 U7915 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n7006), .B1(n7005), .B2(n7004), .ZN(n7007) );
  OAI21_X1 U7916 ( .B1(n7009), .B2(n7008), .A(n7007), .ZN(U3461) );
  AOI21_X1 U7917 ( .B1(REIP_REG_0__SCAN_IN), .B2(DATAWIDTH_REG_0__SCAN_IN), 
        .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n7010) );
  AOI22_X1 U7918 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_0__SCAN_IN), .B1(
        n7010), .B2(n7015), .ZN(n7012) );
  INV_X1 U7919 ( .A(BYTEENABLE_REG_2__SCAN_IN), .ZN(n7011) );
  AOI22_X1 U7920 ( .A1(n7013), .A2(n7012), .B1(n7011), .B2(n7016), .ZN(U3468)
         );
  NOR2_X1 U7921 ( .A1(n7016), .A2(REIP_REG_0__SCAN_IN), .ZN(n7014) );
  AOI22_X1 U7922 ( .A1(n7017), .A2(n7016), .B1(n7015), .B2(n7014), .ZN(U3469)
         );
  NAND2_X1 U7923 ( .A1(n7019), .A2(W_R_N_REG_SCAN_IN), .ZN(n7018) );
  OAI21_X1 U7924 ( .B1(n7019), .B2(READREQUEST_REG_SCAN_IN), .A(n7018), .ZN(
        U3470) );
  MUX2_X1 U7925 ( .A(MORE_REG_SCAN_IN), .B(n7021), .S(n7020), .Z(U3471) );
  AOI211_X1 U7926 ( .C1(n6419), .C2(n7024), .A(n7023), .B(n7022), .ZN(n7031)
         );
  OAI211_X1 U7927 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n7026), .A(n7025), .B(
        STATE2_REG_2__SCAN_IN), .ZN(n7028) );
  AOI21_X1 U7928 ( .B1(STATE2_REG_0__SCAN_IN), .B2(n7028), .A(n7027), .ZN(
        n7030) );
  NAND2_X1 U7929 ( .A1(n7031), .A2(REQUESTPENDING_REG_SCAN_IN), .ZN(n7029) );
  OAI21_X1 U7930 ( .B1(n7031), .B2(n7030), .A(n7029), .ZN(U3472) );
  MUX2_X1 U7931 ( .A(M_IO_N_REG_SCAN_IN), .B(MEMORYFETCH_REG_SCAN_IN), .S(
        n7032), .Z(U3473) );
  OAI21_X1 U7932 ( .B1(n7033), .B2(READREQUEST_REG_SCAN_IN), .A(n7036), .ZN(
        n7034) );
  OAI21_X1 U7933 ( .B1(n7036), .B2(n7035), .A(n7034), .ZN(U3474) );
  CLKBUF_X1 U3648 ( .A(n3777), .Z(n4214) );
  AND2_X2 U3739 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4887) );
  CLKBUF_X2 U3745 ( .A(n3429), .Z(n4812) );
  AND4_X1 U4062 ( .A1(n3237), .A2(n3236), .A3(n3235), .A4(n3232), .ZN(n7037)
         );
  AND2_X1 U4111 ( .A1(n3427), .A2(n3429), .ZN(n7038) );
endmodule

